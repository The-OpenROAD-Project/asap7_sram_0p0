VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_64x4x32_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_64x4x32_6t122 0 0 ;
  SIZE 9.612 BY 43.2 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1010 1.1720 9.5090 1.2200 ;
        RECT 0.1010 2.2520 9.5090 2.3000 ;
        RECT 0.1010 3.3320 9.5090 3.3800 ;
        RECT 0.1010 4.4120 9.5090 4.4600 ;
        RECT 0.1010 5.4920 9.5090 5.5400 ;
        RECT 0.1010 6.5720 9.5090 6.6200 ;
        RECT 0.1010 7.6520 9.5090 7.7000 ;
        RECT 0.1010 8.7320 9.5090 8.7800 ;
        RECT 0.1010 9.8120 9.5090 9.8600 ;
        RECT 0.1010 10.8920 9.5090 10.9400 ;
        RECT 0.1010 11.9720 9.5090 12.0200 ;
        RECT 0.1010 13.0520 9.5090 13.1000 ;
        RECT 0.1010 14.1320 9.5090 14.1800 ;
        RECT 0.1010 15.2120 9.5090 15.2600 ;
        RECT 0.1010 16.2920 9.5090 16.3400 ;
        RECT 0.1010 17.3720 9.5090 17.4200 ;
        RECT 0.1080 17.8590 9.5040 18.0750 ;
        RECT 5.6100 17.5790 5.8730 17.6030 ;
        RECT 5.7410 21.3630 5.8530 21.3870 ;
        RECT 3.9420 21.0270 5.6700 21.2430 ;
        RECT 3.9420 24.1950 5.6700 24.4110 ;
        RECT 0.1010 26.5790 9.5090 26.6270 ;
        RECT 0.1010 27.6590 9.5090 27.7070 ;
        RECT 0.1010 28.7390 9.5090 28.7870 ;
        RECT 0.1010 29.8190 9.5090 29.8670 ;
        RECT 0.1010 30.8990 9.5090 30.9470 ;
        RECT 0.1010 31.9790 9.5090 32.0270 ;
        RECT 0.1010 33.0590 9.5090 33.1070 ;
        RECT 0.1010 34.1390 9.5090 34.1870 ;
        RECT 0.1010 35.2190 9.5090 35.2670 ;
        RECT 0.1010 36.2990 9.5090 36.3470 ;
        RECT 0.1010 37.3790 9.5090 37.4270 ;
        RECT 0.1010 38.4590 9.5090 38.5070 ;
        RECT 0.1010 39.5390 9.5090 39.5870 ;
        RECT 0.1010 40.6190 9.5090 40.6670 ;
        RECT 0.1010 41.6990 9.5090 41.7470 ;
        RECT 0.1010 42.7790 9.5090 42.8270 ;
      LAYER M3  ;
        RECT 9.4770 0.2165 9.4950 1.3765 ;
        RECT 5.8230 0.2170 5.8410 1.3760 ;
        RECT 4.4190 0.2530 4.5090 1.3670 ;
        RECT 3.7710 0.2170 3.7890 1.3760 ;
        RECT 0.1170 0.2165 0.1350 1.3765 ;
        RECT 9.4770 1.2965 9.4950 2.4565 ;
        RECT 5.8230 1.2970 5.8410 2.4560 ;
        RECT 4.4190 1.3330 4.5090 2.4470 ;
        RECT 3.7710 1.2970 3.7890 2.4560 ;
        RECT 0.1170 1.2965 0.1350 2.4565 ;
        RECT 9.4770 2.3765 9.4950 3.5365 ;
        RECT 5.8230 2.3770 5.8410 3.5360 ;
        RECT 4.4190 2.4130 4.5090 3.5270 ;
        RECT 3.7710 2.3770 3.7890 3.5360 ;
        RECT 0.1170 2.3765 0.1350 3.5365 ;
        RECT 9.4770 3.4565 9.4950 4.6165 ;
        RECT 5.8230 3.4570 5.8410 4.6160 ;
        RECT 4.4190 3.4930 4.5090 4.6070 ;
        RECT 3.7710 3.4570 3.7890 4.6160 ;
        RECT 0.1170 3.4565 0.1350 4.6165 ;
        RECT 9.4770 4.5365 9.4950 5.6965 ;
        RECT 5.8230 4.5370 5.8410 5.6960 ;
        RECT 4.4190 4.5730 4.5090 5.6870 ;
        RECT 3.7710 4.5370 3.7890 5.6960 ;
        RECT 0.1170 4.5365 0.1350 5.6965 ;
        RECT 9.4770 5.6165 9.4950 6.7765 ;
        RECT 5.8230 5.6170 5.8410 6.7760 ;
        RECT 4.4190 5.6530 4.5090 6.7670 ;
        RECT 3.7710 5.6170 3.7890 6.7760 ;
        RECT 0.1170 5.6165 0.1350 6.7765 ;
        RECT 9.4770 6.6965 9.4950 7.8565 ;
        RECT 5.8230 6.6970 5.8410 7.8560 ;
        RECT 4.4190 6.7330 4.5090 7.8470 ;
        RECT 3.7710 6.6970 3.7890 7.8560 ;
        RECT 0.1170 6.6965 0.1350 7.8565 ;
        RECT 9.4770 7.7765 9.4950 8.9365 ;
        RECT 5.8230 7.7770 5.8410 8.9360 ;
        RECT 4.4190 7.8130 4.5090 8.9270 ;
        RECT 3.7710 7.7770 3.7890 8.9360 ;
        RECT 0.1170 7.7765 0.1350 8.9365 ;
        RECT 9.4770 8.8565 9.4950 10.0165 ;
        RECT 5.8230 8.8570 5.8410 10.0160 ;
        RECT 4.4190 8.8930 4.5090 10.0070 ;
        RECT 3.7710 8.8570 3.7890 10.0160 ;
        RECT 0.1170 8.8565 0.1350 10.0165 ;
        RECT 9.4770 9.9365 9.4950 11.0965 ;
        RECT 5.8230 9.9370 5.8410 11.0960 ;
        RECT 4.4190 9.9730 4.5090 11.0870 ;
        RECT 3.7710 9.9370 3.7890 11.0960 ;
        RECT 0.1170 9.9365 0.1350 11.0965 ;
        RECT 9.4770 11.0165 9.4950 12.1765 ;
        RECT 5.8230 11.0170 5.8410 12.1760 ;
        RECT 4.4190 11.0530 4.5090 12.1670 ;
        RECT 3.7710 11.0170 3.7890 12.1760 ;
        RECT 0.1170 11.0165 0.1350 12.1765 ;
        RECT 9.4770 12.0965 9.4950 13.2565 ;
        RECT 5.8230 12.0970 5.8410 13.2560 ;
        RECT 4.4190 12.1330 4.5090 13.2470 ;
        RECT 3.7710 12.0970 3.7890 13.2560 ;
        RECT 0.1170 12.0965 0.1350 13.2565 ;
        RECT 9.4770 13.1765 9.4950 14.3365 ;
        RECT 5.8230 13.1770 5.8410 14.3360 ;
        RECT 4.4190 13.2130 4.5090 14.3270 ;
        RECT 3.7710 13.1770 3.7890 14.3360 ;
        RECT 0.1170 13.1765 0.1350 14.3365 ;
        RECT 9.4770 14.2565 9.4950 15.4165 ;
        RECT 5.8230 14.2570 5.8410 15.4160 ;
        RECT 4.4190 14.2930 4.5090 15.4070 ;
        RECT 3.7710 14.2570 3.7890 15.4160 ;
        RECT 0.1170 14.2565 0.1350 15.4165 ;
        RECT 9.4770 15.3365 9.4950 16.4965 ;
        RECT 5.8230 15.3370 5.8410 16.4960 ;
        RECT 4.4190 15.3730 4.5090 16.4870 ;
        RECT 3.7710 15.3370 3.7890 16.4960 ;
        RECT 0.1170 15.3365 0.1350 16.4965 ;
        RECT 9.4770 16.4165 9.4950 17.5765 ;
        RECT 5.8230 16.4170 5.8410 17.5760 ;
        RECT 4.4190 16.4530 4.5090 17.5670 ;
        RECT 3.7710 16.4170 3.7890 17.5760 ;
        RECT 0.1170 16.4165 0.1350 17.5765 ;
        RECT 9.4770 17.4965 9.4950 25.7035 ;
        RECT 5.8230 17.5760 5.8410 17.6675 ;
        RECT 5.8230 21.3160 5.8410 25.6760 ;
        RECT 4.4550 17.8200 4.6890 25.4030 ;
        RECT 4.4190 25.3170 4.5090 25.8520 ;
        RECT 4.4190 17.5400 4.5090 18.0750 ;
        RECT 0.1170 17.4965 0.1350 25.7035 ;
        RECT 9.4770 25.6235 9.4950 26.7835 ;
        RECT 5.8230 25.6240 5.8410 26.7830 ;
        RECT 4.4190 25.6600 4.5090 26.7740 ;
        RECT 3.7710 25.6240 3.7890 26.7830 ;
        RECT 0.1170 25.6235 0.1350 26.7835 ;
        RECT 9.4770 26.7035 9.4950 27.8635 ;
        RECT 5.8230 26.7040 5.8410 27.8630 ;
        RECT 4.4190 26.7400 4.5090 27.8540 ;
        RECT 3.7710 26.7040 3.7890 27.8630 ;
        RECT 0.1170 26.7035 0.1350 27.8635 ;
        RECT 9.4770 27.7835 9.4950 28.9435 ;
        RECT 5.8230 27.7840 5.8410 28.9430 ;
        RECT 4.4190 27.8200 4.5090 28.9340 ;
        RECT 3.7710 27.7840 3.7890 28.9430 ;
        RECT 0.1170 27.7835 0.1350 28.9435 ;
        RECT 9.4770 28.8635 9.4950 30.0235 ;
        RECT 5.8230 28.8640 5.8410 30.0230 ;
        RECT 4.4190 28.9000 4.5090 30.0140 ;
        RECT 3.7710 28.8640 3.7890 30.0230 ;
        RECT 0.1170 28.8635 0.1350 30.0235 ;
        RECT 9.4770 29.9435 9.4950 31.1035 ;
        RECT 5.8230 29.9440 5.8410 31.1030 ;
        RECT 4.4190 29.9800 4.5090 31.0940 ;
        RECT 3.7710 29.9440 3.7890 31.1030 ;
        RECT 0.1170 29.9435 0.1350 31.1035 ;
        RECT 9.4770 31.0235 9.4950 32.1835 ;
        RECT 5.8230 31.0240 5.8410 32.1830 ;
        RECT 4.4190 31.0600 4.5090 32.1740 ;
        RECT 3.7710 31.0240 3.7890 32.1830 ;
        RECT 0.1170 31.0235 0.1350 32.1835 ;
        RECT 9.4770 32.1035 9.4950 33.2635 ;
        RECT 5.8230 32.1040 5.8410 33.2630 ;
        RECT 4.4190 32.1400 4.5090 33.2540 ;
        RECT 3.7710 32.1040 3.7890 33.2630 ;
        RECT 0.1170 32.1035 0.1350 33.2635 ;
        RECT 9.4770 33.1835 9.4950 34.3435 ;
        RECT 5.8230 33.1840 5.8410 34.3430 ;
        RECT 4.4190 33.2200 4.5090 34.3340 ;
        RECT 3.7710 33.1840 3.7890 34.3430 ;
        RECT 0.1170 33.1835 0.1350 34.3435 ;
        RECT 9.4770 34.2635 9.4950 35.4235 ;
        RECT 5.8230 34.2640 5.8410 35.4230 ;
        RECT 4.4190 34.3000 4.5090 35.4140 ;
        RECT 3.7710 34.2640 3.7890 35.4230 ;
        RECT 0.1170 34.2635 0.1350 35.4235 ;
        RECT 9.4770 35.3435 9.4950 36.5035 ;
        RECT 5.8230 35.3440 5.8410 36.5030 ;
        RECT 4.4190 35.3800 4.5090 36.4940 ;
        RECT 3.7710 35.3440 3.7890 36.5030 ;
        RECT 0.1170 35.3435 0.1350 36.5035 ;
        RECT 9.4770 36.4235 9.4950 37.5835 ;
        RECT 5.8230 36.4240 5.8410 37.5830 ;
        RECT 4.4190 36.4600 4.5090 37.5740 ;
        RECT 3.7710 36.4240 3.7890 37.5830 ;
        RECT 0.1170 36.4235 0.1350 37.5835 ;
        RECT 9.4770 37.5035 9.4950 38.6635 ;
        RECT 5.8230 37.5040 5.8410 38.6630 ;
        RECT 4.4190 37.5400 4.5090 38.6540 ;
        RECT 3.7710 37.5040 3.7890 38.6630 ;
        RECT 0.1170 37.5035 0.1350 38.6635 ;
        RECT 9.4770 38.5835 9.4950 39.7435 ;
        RECT 5.8230 38.5840 5.8410 39.7430 ;
        RECT 4.4190 38.6200 4.5090 39.7340 ;
        RECT 3.7710 38.5840 3.7890 39.7430 ;
        RECT 0.1170 38.5835 0.1350 39.7435 ;
        RECT 9.4770 39.6635 9.4950 40.8235 ;
        RECT 5.8230 39.6640 5.8410 40.8230 ;
        RECT 4.4190 39.7000 4.5090 40.8140 ;
        RECT 3.7710 39.6640 3.7890 40.8230 ;
        RECT 0.1170 39.6635 0.1350 40.8235 ;
        RECT 9.4770 40.7435 9.4950 41.9035 ;
        RECT 5.8230 40.7440 5.8410 41.9030 ;
        RECT 4.4190 40.7800 4.5090 41.8940 ;
        RECT 3.7710 40.7440 3.7890 41.9030 ;
        RECT 0.1170 40.7435 0.1350 41.9035 ;
        RECT 9.4770 41.8235 9.4950 42.9835 ;
        RECT 5.8230 41.8240 5.8410 42.9830 ;
        RECT 4.4190 41.8600 4.5090 42.9740 ;
        RECT 3.7710 41.8240 3.7890 42.9830 ;
        RECT 0.1170 41.8235 0.1350 42.9835 ;
      LAYER V3  ;
        RECT 0.1170 1.1720 0.1350 1.2200 ;
        RECT 3.7710 1.1720 3.7890 1.2200 ;
        RECT 4.4190 1.1720 4.5090 1.2200 ;
        RECT 5.8230 1.1720 5.8410 1.2200 ;
        RECT 9.4770 1.1720 9.4950 1.2200 ;
        RECT 0.1170 2.2520 0.1350 2.3000 ;
        RECT 3.7710 2.2520 3.7890 2.3000 ;
        RECT 4.4190 2.2520 4.5090 2.3000 ;
        RECT 5.8230 2.2520 5.8410 2.3000 ;
        RECT 9.4770 2.2520 9.4950 2.3000 ;
        RECT 0.1170 3.3320 0.1350 3.3800 ;
        RECT 3.7710 3.3320 3.7890 3.3800 ;
        RECT 4.4190 3.3320 4.5090 3.3800 ;
        RECT 5.8230 3.3320 5.8410 3.3800 ;
        RECT 9.4770 3.3320 9.4950 3.3800 ;
        RECT 0.1170 4.4120 0.1350 4.4600 ;
        RECT 3.7710 4.4120 3.7890 4.4600 ;
        RECT 4.4190 4.4120 4.5090 4.4600 ;
        RECT 5.8230 4.4120 5.8410 4.4600 ;
        RECT 9.4770 4.4120 9.4950 4.4600 ;
        RECT 0.1170 5.4920 0.1350 5.5400 ;
        RECT 3.7710 5.4920 3.7890 5.5400 ;
        RECT 4.4190 5.4920 4.5090 5.5400 ;
        RECT 5.8230 5.4920 5.8410 5.5400 ;
        RECT 9.4770 5.4920 9.4950 5.5400 ;
        RECT 0.1170 6.5720 0.1350 6.6200 ;
        RECT 3.7710 6.5720 3.7890 6.6200 ;
        RECT 4.4190 6.5720 4.5090 6.6200 ;
        RECT 5.8230 6.5720 5.8410 6.6200 ;
        RECT 9.4770 6.5720 9.4950 6.6200 ;
        RECT 0.1170 7.6520 0.1350 7.7000 ;
        RECT 3.7710 7.6520 3.7890 7.7000 ;
        RECT 4.4190 7.6520 4.5090 7.7000 ;
        RECT 5.8230 7.6520 5.8410 7.7000 ;
        RECT 9.4770 7.6520 9.4950 7.7000 ;
        RECT 0.1170 8.7320 0.1350 8.7800 ;
        RECT 3.7710 8.7320 3.7890 8.7800 ;
        RECT 4.4190 8.7320 4.5090 8.7800 ;
        RECT 5.8230 8.7320 5.8410 8.7800 ;
        RECT 9.4770 8.7320 9.4950 8.7800 ;
        RECT 0.1170 9.8120 0.1350 9.8600 ;
        RECT 3.7710 9.8120 3.7890 9.8600 ;
        RECT 4.4190 9.8120 4.5090 9.8600 ;
        RECT 5.8230 9.8120 5.8410 9.8600 ;
        RECT 9.4770 9.8120 9.4950 9.8600 ;
        RECT 0.1170 10.8920 0.1350 10.9400 ;
        RECT 3.7710 10.8920 3.7890 10.9400 ;
        RECT 4.4190 10.8920 4.5090 10.9400 ;
        RECT 5.8230 10.8920 5.8410 10.9400 ;
        RECT 9.4770 10.8920 9.4950 10.9400 ;
        RECT 0.1170 11.9720 0.1350 12.0200 ;
        RECT 3.7710 11.9720 3.7890 12.0200 ;
        RECT 4.4190 11.9720 4.5090 12.0200 ;
        RECT 5.8230 11.9720 5.8410 12.0200 ;
        RECT 9.4770 11.9720 9.4950 12.0200 ;
        RECT 0.1170 13.0520 0.1350 13.1000 ;
        RECT 3.7710 13.0520 3.7890 13.1000 ;
        RECT 4.4190 13.0520 4.5090 13.1000 ;
        RECT 5.8230 13.0520 5.8410 13.1000 ;
        RECT 9.4770 13.0520 9.4950 13.1000 ;
        RECT 0.1170 14.1320 0.1350 14.1800 ;
        RECT 3.7710 14.1320 3.7890 14.1800 ;
        RECT 4.4190 14.1320 4.5090 14.1800 ;
        RECT 5.8230 14.1320 5.8410 14.1800 ;
        RECT 9.4770 14.1320 9.4950 14.1800 ;
        RECT 0.1170 15.2120 0.1350 15.2600 ;
        RECT 3.7710 15.2120 3.7890 15.2600 ;
        RECT 4.4190 15.2120 4.5090 15.2600 ;
        RECT 5.8230 15.2120 5.8410 15.2600 ;
        RECT 9.4770 15.2120 9.4950 15.2600 ;
        RECT 0.1170 16.2920 0.1350 16.3400 ;
        RECT 3.7710 16.2920 3.7890 16.3400 ;
        RECT 4.4190 16.2920 4.5090 16.3400 ;
        RECT 5.8230 16.2920 5.8410 16.3400 ;
        RECT 9.4770 16.2920 9.4950 16.3400 ;
        RECT 0.1170 17.3720 0.1350 17.4200 ;
        RECT 3.7710 17.3720 3.7890 17.4200 ;
        RECT 4.4190 17.3720 4.5090 17.4200 ;
        RECT 5.8230 17.3720 5.8410 17.4200 ;
        RECT 9.4770 17.3720 9.4950 17.4200 ;
        RECT 0.1170 17.8590 0.1350 18.0750 ;
        RECT 4.4590 24.1950 4.4770 24.4110 ;
        RECT 4.4590 21.0270 4.4770 21.2430 ;
        RECT 4.4590 17.8590 4.4770 18.0750 ;
        RECT 4.5110 24.1950 4.5290 24.4110 ;
        RECT 4.5110 21.0270 4.5290 21.2430 ;
        RECT 4.5110 17.8590 4.5290 18.0750 ;
        RECT 4.5630 24.1950 4.5810 24.4110 ;
        RECT 4.5630 21.0270 4.5810 21.2430 ;
        RECT 4.5630 17.8590 4.5810 18.0750 ;
        RECT 4.6150 24.1950 4.6330 24.4110 ;
        RECT 4.6150 21.0270 4.6330 21.2430 ;
        RECT 4.6150 17.8590 4.6330 18.0750 ;
        RECT 4.6670 24.1950 4.6850 24.4110 ;
        RECT 4.6670 21.0270 4.6850 21.2430 ;
        RECT 4.6670 17.8590 4.6850 18.0750 ;
        RECT 5.8230 21.3630 5.8410 21.3870 ;
        RECT 5.8230 17.5790 5.8410 17.6030 ;
        RECT 0.1170 26.5790 0.1350 26.6270 ;
        RECT 3.7710 26.5790 3.7890 26.6270 ;
        RECT 4.4190 26.5790 4.5090 26.6270 ;
        RECT 5.8230 26.5790 5.8410 26.6270 ;
        RECT 9.4770 26.5790 9.4950 26.6270 ;
        RECT 0.1170 27.6590 0.1350 27.7070 ;
        RECT 3.7710 27.6590 3.7890 27.7070 ;
        RECT 4.4190 27.6590 4.5090 27.7070 ;
        RECT 5.8230 27.6590 5.8410 27.7070 ;
        RECT 9.4770 27.6590 9.4950 27.7070 ;
        RECT 0.1170 28.7390 0.1350 28.7870 ;
        RECT 3.7710 28.7390 3.7890 28.7870 ;
        RECT 4.4190 28.7390 4.5090 28.7870 ;
        RECT 5.8230 28.7390 5.8410 28.7870 ;
        RECT 9.4770 28.7390 9.4950 28.7870 ;
        RECT 0.1170 29.8190 0.1350 29.8670 ;
        RECT 3.7710 29.8190 3.7890 29.8670 ;
        RECT 4.4190 29.8190 4.5090 29.8670 ;
        RECT 5.8230 29.8190 5.8410 29.8670 ;
        RECT 9.4770 29.8190 9.4950 29.8670 ;
        RECT 0.1170 30.8990 0.1350 30.9470 ;
        RECT 3.7710 30.8990 3.7890 30.9470 ;
        RECT 4.4190 30.8990 4.5090 30.9470 ;
        RECT 5.8230 30.8990 5.8410 30.9470 ;
        RECT 9.4770 30.8990 9.4950 30.9470 ;
        RECT 0.1170 31.9790 0.1350 32.0270 ;
        RECT 3.7710 31.9790 3.7890 32.0270 ;
        RECT 4.4190 31.9790 4.5090 32.0270 ;
        RECT 5.8230 31.9790 5.8410 32.0270 ;
        RECT 9.4770 31.9790 9.4950 32.0270 ;
        RECT 0.1170 33.0590 0.1350 33.1070 ;
        RECT 3.7710 33.0590 3.7890 33.1070 ;
        RECT 4.4190 33.0590 4.5090 33.1070 ;
        RECT 5.8230 33.0590 5.8410 33.1070 ;
        RECT 9.4770 33.0590 9.4950 33.1070 ;
        RECT 0.1170 34.1390 0.1350 34.1870 ;
        RECT 3.7710 34.1390 3.7890 34.1870 ;
        RECT 4.4190 34.1390 4.5090 34.1870 ;
        RECT 5.8230 34.1390 5.8410 34.1870 ;
        RECT 9.4770 34.1390 9.4950 34.1870 ;
        RECT 0.1170 35.2190 0.1350 35.2670 ;
        RECT 3.7710 35.2190 3.7890 35.2670 ;
        RECT 4.4190 35.2190 4.5090 35.2670 ;
        RECT 5.8230 35.2190 5.8410 35.2670 ;
        RECT 9.4770 35.2190 9.4950 35.2670 ;
        RECT 0.1170 36.2990 0.1350 36.3470 ;
        RECT 3.7710 36.2990 3.7890 36.3470 ;
        RECT 4.4190 36.2990 4.5090 36.3470 ;
        RECT 5.8230 36.2990 5.8410 36.3470 ;
        RECT 9.4770 36.2990 9.4950 36.3470 ;
        RECT 0.1170 37.3790 0.1350 37.4270 ;
        RECT 3.7710 37.3790 3.7890 37.4270 ;
        RECT 4.4190 37.3790 4.5090 37.4270 ;
        RECT 5.8230 37.3790 5.8410 37.4270 ;
        RECT 9.4770 37.3790 9.4950 37.4270 ;
        RECT 0.1170 38.4590 0.1350 38.5070 ;
        RECT 3.7710 38.4590 3.7890 38.5070 ;
        RECT 4.4190 38.4590 4.5090 38.5070 ;
        RECT 5.8230 38.4590 5.8410 38.5070 ;
        RECT 9.4770 38.4590 9.4950 38.5070 ;
        RECT 0.1170 39.5390 0.1350 39.5870 ;
        RECT 3.7710 39.5390 3.7890 39.5870 ;
        RECT 4.4190 39.5390 4.5090 39.5870 ;
        RECT 5.8230 39.5390 5.8410 39.5870 ;
        RECT 9.4770 39.5390 9.4950 39.5870 ;
        RECT 0.1170 40.6190 0.1350 40.6670 ;
        RECT 3.7710 40.6190 3.7890 40.6670 ;
        RECT 4.4190 40.6190 4.5090 40.6670 ;
        RECT 5.8230 40.6190 5.8410 40.6670 ;
        RECT 9.4770 40.6190 9.4950 40.6670 ;
        RECT 0.1170 41.6990 0.1350 41.7470 ;
        RECT 3.7710 41.6990 3.7890 41.7470 ;
        RECT 4.4190 41.6990 4.5090 41.7470 ;
        RECT 5.8230 41.6990 5.8410 41.7470 ;
        RECT 9.4770 41.6990 9.4950 41.7470 ;
        RECT 0.1170 42.7790 0.1350 42.8270 ;
        RECT 3.7710 42.7790 3.7890 42.8270 ;
        RECT 4.4190 42.7790 4.5090 42.8270 ;
        RECT 5.8230 42.7790 5.8410 42.8270 ;
        RECT 9.4770 42.7790 9.4950 42.8270 ;
      LAYER M5  ;
        RECT 5.7590 17.5610 5.7830 21.4050 ;
      LAYER V4  ;
        RECT 5.7590 21.3630 5.7830 21.3870 ;
        RECT 5.7590 17.5790 5.7830 17.6030 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1010 1.0760 9.5040 1.1240 ;
        RECT 0.1010 2.1560 9.5040 2.2040 ;
        RECT 0.1010 3.2360 9.5040 3.2840 ;
        RECT 0.1010 4.3160 9.5040 4.3640 ;
        RECT 0.1010 5.3960 9.5040 5.4440 ;
        RECT 0.1010 6.4760 9.5040 6.5240 ;
        RECT 0.1010 7.5560 9.5040 7.6040 ;
        RECT 0.1010 8.6360 9.5040 8.6840 ;
        RECT 0.1010 9.7160 9.5040 9.7640 ;
        RECT 0.1010 10.7960 9.5040 10.8440 ;
        RECT 0.1010 11.8760 9.5040 11.9240 ;
        RECT 0.1010 12.9560 9.5040 13.0040 ;
        RECT 0.1010 14.0360 9.5040 14.0840 ;
        RECT 0.1010 15.1160 9.5040 15.1640 ;
        RECT 0.1010 16.1960 9.5040 16.2440 ;
        RECT 0.1010 17.2760 9.5040 17.3240 ;
        RECT 0.1080 18.2910 9.5040 18.5070 ;
        RECT 3.9420 21.4590 5.6700 21.6750 ;
        RECT 3.9420 24.6270 5.6700 24.8430 ;
        RECT 0.1010 26.4830 9.5040 26.5310 ;
        RECT 0.1010 27.5630 9.5040 27.6110 ;
        RECT 0.1010 28.6430 9.5040 28.6910 ;
        RECT 0.1010 29.7230 9.5040 29.7710 ;
        RECT 0.1010 30.8030 9.5040 30.8510 ;
        RECT 0.1010 31.8830 9.5040 31.9310 ;
        RECT 0.1010 32.9630 9.5040 33.0110 ;
        RECT 0.1010 34.0430 9.5040 34.0910 ;
        RECT 0.1010 35.1230 9.5040 35.1710 ;
        RECT 0.1010 36.2030 9.5040 36.2510 ;
        RECT 0.1010 37.2830 9.5040 37.3310 ;
        RECT 0.1010 38.3630 9.5040 38.4110 ;
        RECT 0.1010 39.4430 9.5040 39.4910 ;
        RECT 0.1010 40.5230 9.5040 40.5710 ;
        RECT 0.1010 41.6030 9.5040 41.6510 ;
        RECT 0.1010 42.6830 9.5040 42.7310 ;
      LAYER M3  ;
        RECT 9.4410 0.2165 9.4590 1.3765 ;
        RECT 5.8770 0.2165 5.8950 1.3765 ;
        RECT 5.1120 0.2530 5.1480 1.3670 ;
        RECT 4.9590 0.2530 4.9860 1.3670 ;
        RECT 3.7170 0.2165 3.7350 1.3765 ;
        RECT 0.1530 0.2165 0.1710 1.3765 ;
        RECT 9.4410 1.2965 9.4590 2.4565 ;
        RECT 5.8770 1.2965 5.8950 2.4565 ;
        RECT 5.1120 1.3330 5.1480 2.4470 ;
        RECT 4.9590 1.3330 4.9860 2.4470 ;
        RECT 3.7170 1.2965 3.7350 2.4565 ;
        RECT 0.1530 1.2965 0.1710 2.4565 ;
        RECT 9.4410 2.3765 9.4590 3.5365 ;
        RECT 5.8770 2.3765 5.8950 3.5365 ;
        RECT 5.1120 2.4130 5.1480 3.5270 ;
        RECT 4.9590 2.4130 4.9860 3.5270 ;
        RECT 3.7170 2.3765 3.7350 3.5365 ;
        RECT 0.1530 2.3765 0.1710 3.5365 ;
        RECT 9.4410 3.4565 9.4590 4.6165 ;
        RECT 5.8770 3.4565 5.8950 4.6165 ;
        RECT 5.1120 3.4930 5.1480 4.6070 ;
        RECT 4.9590 3.4930 4.9860 4.6070 ;
        RECT 3.7170 3.4565 3.7350 4.6165 ;
        RECT 0.1530 3.4565 0.1710 4.6165 ;
        RECT 9.4410 4.5365 9.4590 5.6965 ;
        RECT 5.8770 4.5365 5.8950 5.6965 ;
        RECT 5.1120 4.5730 5.1480 5.6870 ;
        RECT 4.9590 4.5730 4.9860 5.6870 ;
        RECT 3.7170 4.5365 3.7350 5.6965 ;
        RECT 0.1530 4.5365 0.1710 5.6965 ;
        RECT 9.4410 5.6165 9.4590 6.7765 ;
        RECT 5.8770 5.6165 5.8950 6.7765 ;
        RECT 5.1120 5.6530 5.1480 6.7670 ;
        RECT 4.9590 5.6530 4.9860 6.7670 ;
        RECT 3.7170 5.6165 3.7350 6.7765 ;
        RECT 0.1530 5.6165 0.1710 6.7765 ;
        RECT 9.4410 6.6965 9.4590 7.8565 ;
        RECT 5.8770 6.6965 5.8950 7.8565 ;
        RECT 5.1120 6.7330 5.1480 7.8470 ;
        RECT 4.9590 6.7330 4.9860 7.8470 ;
        RECT 3.7170 6.6965 3.7350 7.8565 ;
        RECT 0.1530 6.6965 0.1710 7.8565 ;
        RECT 9.4410 7.7765 9.4590 8.9365 ;
        RECT 5.8770 7.7765 5.8950 8.9365 ;
        RECT 5.1120 7.8130 5.1480 8.9270 ;
        RECT 4.9590 7.8130 4.9860 8.9270 ;
        RECT 3.7170 7.7765 3.7350 8.9365 ;
        RECT 0.1530 7.7765 0.1710 8.9365 ;
        RECT 9.4410 8.8565 9.4590 10.0165 ;
        RECT 5.8770 8.8565 5.8950 10.0165 ;
        RECT 5.1120 8.8930 5.1480 10.0070 ;
        RECT 4.9590 8.8930 4.9860 10.0070 ;
        RECT 3.7170 8.8565 3.7350 10.0165 ;
        RECT 0.1530 8.8565 0.1710 10.0165 ;
        RECT 9.4410 9.9365 9.4590 11.0965 ;
        RECT 5.8770 9.9365 5.8950 11.0965 ;
        RECT 5.1120 9.9730 5.1480 11.0870 ;
        RECT 4.9590 9.9730 4.9860 11.0870 ;
        RECT 3.7170 9.9365 3.7350 11.0965 ;
        RECT 0.1530 9.9365 0.1710 11.0965 ;
        RECT 9.4410 11.0165 9.4590 12.1765 ;
        RECT 5.8770 11.0165 5.8950 12.1765 ;
        RECT 5.1120 11.0530 5.1480 12.1670 ;
        RECT 4.9590 11.0530 4.9860 12.1670 ;
        RECT 3.7170 11.0165 3.7350 12.1765 ;
        RECT 0.1530 11.0165 0.1710 12.1765 ;
        RECT 9.4410 12.0965 9.4590 13.2565 ;
        RECT 5.8770 12.0965 5.8950 13.2565 ;
        RECT 5.1120 12.1330 5.1480 13.2470 ;
        RECT 4.9590 12.1330 4.9860 13.2470 ;
        RECT 3.7170 12.0965 3.7350 13.2565 ;
        RECT 0.1530 12.0965 0.1710 13.2565 ;
        RECT 9.4410 13.1765 9.4590 14.3365 ;
        RECT 5.8770 13.1765 5.8950 14.3365 ;
        RECT 5.1120 13.2130 5.1480 14.3270 ;
        RECT 4.9590 13.2130 4.9860 14.3270 ;
        RECT 3.7170 13.1765 3.7350 14.3365 ;
        RECT 0.1530 13.1765 0.1710 14.3365 ;
        RECT 9.4410 14.2565 9.4590 15.4165 ;
        RECT 5.8770 14.2565 5.8950 15.4165 ;
        RECT 5.1120 14.2930 5.1480 15.4070 ;
        RECT 4.9590 14.2930 4.9860 15.4070 ;
        RECT 3.7170 14.2565 3.7350 15.4165 ;
        RECT 0.1530 14.2565 0.1710 15.4165 ;
        RECT 9.4410 15.3365 9.4590 16.4965 ;
        RECT 5.8770 15.3365 5.8950 16.4965 ;
        RECT 5.1120 15.3730 5.1480 16.4870 ;
        RECT 4.9590 15.3730 4.9860 16.4870 ;
        RECT 3.7170 15.3365 3.7350 16.4965 ;
        RECT 0.1530 15.3365 0.1710 16.4965 ;
        RECT 9.4410 16.4165 9.4590 17.5765 ;
        RECT 5.8770 16.4165 5.8950 17.5765 ;
        RECT 5.1120 16.4530 5.1480 17.5670 ;
        RECT 4.9590 16.4530 4.9860 17.5670 ;
        RECT 3.7170 16.4165 3.7350 17.5765 ;
        RECT 0.1530 16.4165 0.1710 17.5765 ;
        RECT 9.4410 17.4965 9.4590 25.7035 ;
        RECT 5.8770 17.4965 5.8950 25.7035 ;
        RECT 4.9230 17.7200 5.1570 25.4030 ;
        RECT 5.1120 17.5400 5.1480 25.6770 ;
        RECT 4.9590 17.5400 4.9860 25.6740 ;
        RECT 3.7170 17.4965 3.7350 25.7035 ;
        RECT 0.1530 17.4965 0.1710 25.7035 ;
        RECT 9.4410 25.6235 9.4590 26.7835 ;
        RECT 5.8770 25.6235 5.8950 26.7835 ;
        RECT 5.1120 25.6600 5.1480 26.7740 ;
        RECT 4.9590 25.6600 4.9860 26.7740 ;
        RECT 3.7170 25.6235 3.7350 26.7835 ;
        RECT 0.1530 25.6235 0.1710 26.7835 ;
        RECT 9.4410 26.7035 9.4590 27.8635 ;
        RECT 5.8770 26.7035 5.8950 27.8635 ;
        RECT 5.1120 26.7400 5.1480 27.8540 ;
        RECT 4.9590 26.7400 4.9860 27.8540 ;
        RECT 3.7170 26.7035 3.7350 27.8635 ;
        RECT 0.1530 26.7035 0.1710 27.8635 ;
        RECT 9.4410 27.7835 9.4590 28.9435 ;
        RECT 5.8770 27.7835 5.8950 28.9435 ;
        RECT 5.1120 27.8200 5.1480 28.9340 ;
        RECT 4.9590 27.8200 4.9860 28.9340 ;
        RECT 3.7170 27.7835 3.7350 28.9435 ;
        RECT 0.1530 27.7835 0.1710 28.9435 ;
        RECT 9.4410 28.8635 9.4590 30.0235 ;
        RECT 5.8770 28.8635 5.8950 30.0235 ;
        RECT 5.1120 28.9000 5.1480 30.0140 ;
        RECT 4.9590 28.9000 4.9860 30.0140 ;
        RECT 3.7170 28.8635 3.7350 30.0235 ;
        RECT 0.1530 28.8635 0.1710 30.0235 ;
        RECT 9.4410 29.9435 9.4590 31.1035 ;
        RECT 5.8770 29.9435 5.8950 31.1035 ;
        RECT 5.1120 29.9800 5.1480 31.0940 ;
        RECT 4.9590 29.9800 4.9860 31.0940 ;
        RECT 3.7170 29.9435 3.7350 31.1035 ;
        RECT 0.1530 29.9435 0.1710 31.1035 ;
        RECT 9.4410 31.0235 9.4590 32.1835 ;
        RECT 5.8770 31.0235 5.8950 32.1835 ;
        RECT 5.1120 31.0600 5.1480 32.1740 ;
        RECT 4.9590 31.0600 4.9860 32.1740 ;
        RECT 3.7170 31.0235 3.7350 32.1835 ;
        RECT 0.1530 31.0235 0.1710 32.1835 ;
        RECT 9.4410 32.1035 9.4590 33.2635 ;
        RECT 5.8770 32.1035 5.8950 33.2635 ;
        RECT 5.1120 32.1400 5.1480 33.2540 ;
        RECT 4.9590 32.1400 4.9860 33.2540 ;
        RECT 3.7170 32.1035 3.7350 33.2635 ;
        RECT 0.1530 32.1035 0.1710 33.2635 ;
        RECT 9.4410 33.1835 9.4590 34.3435 ;
        RECT 5.8770 33.1835 5.8950 34.3435 ;
        RECT 5.1120 33.2200 5.1480 34.3340 ;
        RECT 4.9590 33.2200 4.9860 34.3340 ;
        RECT 3.7170 33.1835 3.7350 34.3435 ;
        RECT 0.1530 33.1835 0.1710 34.3435 ;
        RECT 9.4410 34.2635 9.4590 35.4235 ;
        RECT 5.8770 34.2635 5.8950 35.4235 ;
        RECT 5.1120 34.3000 5.1480 35.4140 ;
        RECT 4.9590 34.3000 4.9860 35.4140 ;
        RECT 3.7170 34.2635 3.7350 35.4235 ;
        RECT 0.1530 34.2635 0.1710 35.4235 ;
        RECT 9.4410 35.3435 9.4590 36.5035 ;
        RECT 5.8770 35.3435 5.8950 36.5035 ;
        RECT 5.1120 35.3800 5.1480 36.4940 ;
        RECT 4.9590 35.3800 4.9860 36.4940 ;
        RECT 3.7170 35.3435 3.7350 36.5035 ;
        RECT 0.1530 35.3435 0.1710 36.5035 ;
        RECT 9.4410 36.4235 9.4590 37.5835 ;
        RECT 5.8770 36.4235 5.8950 37.5835 ;
        RECT 5.1120 36.4600 5.1480 37.5740 ;
        RECT 4.9590 36.4600 4.9860 37.5740 ;
        RECT 3.7170 36.4235 3.7350 37.5835 ;
        RECT 0.1530 36.4235 0.1710 37.5835 ;
        RECT 9.4410 37.5035 9.4590 38.6635 ;
        RECT 5.8770 37.5035 5.8950 38.6635 ;
        RECT 5.1120 37.5400 5.1480 38.6540 ;
        RECT 4.9590 37.5400 4.9860 38.6540 ;
        RECT 3.7170 37.5035 3.7350 38.6635 ;
        RECT 0.1530 37.5035 0.1710 38.6635 ;
        RECT 9.4410 38.5835 9.4590 39.7435 ;
        RECT 5.8770 38.5835 5.8950 39.7435 ;
        RECT 5.1120 38.6200 5.1480 39.7340 ;
        RECT 4.9590 38.6200 4.9860 39.7340 ;
        RECT 3.7170 38.5835 3.7350 39.7435 ;
        RECT 0.1530 38.5835 0.1710 39.7435 ;
        RECT 9.4410 39.6635 9.4590 40.8235 ;
        RECT 5.8770 39.6635 5.8950 40.8235 ;
        RECT 5.1120 39.7000 5.1480 40.8140 ;
        RECT 4.9590 39.7000 4.9860 40.8140 ;
        RECT 3.7170 39.6635 3.7350 40.8235 ;
        RECT 0.1530 39.6635 0.1710 40.8235 ;
        RECT 9.4410 40.7435 9.4590 41.9035 ;
        RECT 5.8770 40.7435 5.8950 41.9035 ;
        RECT 5.1120 40.7800 5.1480 41.8940 ;
        RECT 4.9590 40.7800 4.9860 41.8940 ;
        RECT 3.7170 40.7435 3.7350 41.9035 ;
        RECT 0.1530 40.7435 0.1710 41.9035 ;
        RECT 9.4410 41.8235 9.4590 42.9835 ;
        RECT 5.8770 41.8235 5.8950 42.9835 ;
        RECT 5.1120 41.8600 5.1480 42.9740 ;
        RECT 4.9590 41.8600 4.9860 42.9740 ;
        RECT 3.7170 41.8235 3.7350 42.9835 ;
        RECT 0.1530 41.8235 0.1710 42.9835 ;
      LAYER V3  ;
        RECT 0.1530 1.0760 0.1710 1.1240 ;
        RECT 3.7170 1.0760 3.7350 1.1240 ;
        RECT 4.9590 1.0760 4.9860 1.1240 ;
        RECT 5.1120 1.0760 5.1480 1.1240 ;
        RECT 5.8770 1.0760 5.8950 1.1240 ;
        RECT 9.4410 1.0760 9.4590 1.1240 ;
        RECT 0.1530 2.1560 0.1710 2.2040 ;
        RECT 3.7170 2.1560 3.7350 2.2040 ;
        RECT 4.9590 2.1560 4.9860 2.2040 ;
        RECT 5.1120 2.1560 5.1480 2.2040 ;
        RECT 5.8770 2.1560 5.8950 2.2040 ;
        RECT 9.4410 2.1560 9.4590 2.2040 ;
        RECT 0.1530 3.2360 0.1710 3.2840 ;
        RECT 3.7170 3.2360 3.7350 3.2840 ;
        RECT 4.9590 3.2360 4.9860 3.2840 ;
        RECT 5.1120 3.2360 5.1480 3.2840 ;
        RECT 5.8770 3.2360 5.8950 3.2840 ;
        RECT 9.4410 3.2360 9.4590 3.2840 ;
        RECT 0.1530 4.3160 0.1710 4.3640 ;
        RECT 3.7170 4.3160 3.7350 4.3640 ;
        RECT 4.9590 4.3160 4.9860 4.3640 ;
        RECT 5.1120 4.3160 5.1480 4.3640 ;
        RECT 5.8770 4.3160 5.8950 4.3640 ;
        RECT 9.4410 4.3160 9.4590 4.3640 ;
        RECT 0.1530 5.3960 0.1710 5.4440 ;
        RECT 3.7170 5.3960 3.7350 5.4440 ;
        RECT 4.9590 5.3960 4.9860 5.4440 ;
        RECT 5.1120 5.3960 5.1480 5.4440 ;
        RECT 5.8770 5.3960 5.8950 5.4440 ;
        RECT 9.4410 5.3960 9.4590 5.4440 ;
        RECT 0.1530 6.4760 0.1710 6.5240 ;
        RECT 3.7170 6.4760 3.7350 6.5240 ;
        RECT 4.9590 6.4760 4.9860 6.5240 ;
        RECT 5.1120 6.4760 5.1480 6.5240 ;
        RECT 5.8770 6.4760 5.8950 6.5240 ;
        RECT 9.4410 6.4760 9.4590 6.5240 ;
        RECT 0.1530 7.5560 0.1710 7.6040 ;
        RECT 3.7170 7.5560 3.7350 7.6040 ;
        RECT 4.9590 7.5560 4.9860 7.6040 ;
        RECT 5.1120 7.5560 5.1480 7.6040 ;
        RECT 5.8770 7.5560 5.8950 7.6040 ;
        RECT 9.4410 7.5560 9.4590 7.6040 ;
        RECT 0.1530 8.6360 0.1710 8.6840 ;
        RECT 3.7170 8.6360 3.7350 8.6840 ;
        RECT 4.9590 8.6360 4.9860 8.6840 ;
        RECT 5.1120 8.6360 5.1480 8.6840 ;
        RECT 5.8770 8.6360 5.8950 8.6840 ;
        RECT 9.4410 8.6360 9.4590 8.6840 ;
        RECT 0.1530 9.7160 0.1710 9.7640 ;
        RECT 3.7170 9.7160 3.7350 9.7640 ;
        RECT 4.9590 9.7160 4.9860 9.7640 ;
        RECT 5.1120 9.7160 5.1480 9.7640 ;
        RECT 5.8770 9.7160 5.8950 9.7640 ;
        RECT 9.4410 9.7160 9.4590 9.7640 ;
        RECT 0.1530 10.7960 0.1710 10.8440 ;
        RECT 3.7170 10.7960 3.7350 10.8440 ;
        RECT 4.9590 10.7960 4.9860 10.8440 ;
        RECT 5.1120 10.7960 5.1480 10.8440 ;
        RECT 5.8770 10.7960 5.8950 10.8440 ;
        RECT 9.4410 10.7960 9.4590 10.8440 ;
        RECT 0.1530 11.8760 0.1710 11.9240 ;
        RECT 3.7170 11.8760 3.7350 11.9240 ;
        RECT 4.9590 11.8760 4.9860 11.9240 ;
        RECT 5.1120 11.8760 5.1480 11.9240 ;
        RECT 5.8770 11.8760 5.8950 11.9240 ;
        RECT 9.4410 11.8760 9.4590 11.9240 ;
        RECT 0.1530 12.9560 0.1710 13.0040 ;
        RECT 3.7170 12.9560 3.7350 13.0040 ;
        RECT 4.9590 12.9560 4.9860 13.0040 ;
        RECT 5.1120 12.9560 5.1480 13.0040 ;
        RECT 5.8770 12.9560 5.8950 13.0040 ;
        RECT 9.4410 12.9560 9.4590 13.0040 ;
        RECT 0.1530 14.0360 0.1710 14.0840 ;
        RECT 3.7170 14.0360 3.7350 14.0840 ;
        RECT 4.9590 14.0360 4.9860 14.0840 ;
        RECT 5.1120 14.0360 5.1480 14.0840 ;
        RECT 5.8770 14.0360 5.8950 14.0840 ;
        RECT 9.4410 14.0360 9.4590 14.0840 ;
        RECT 0.1530 15.1160 0.1710 15.1640 ;
        RECT 3.7170 15.1160 3.7350 15.1640 ;
        RECT 4.9590 15.1160 4.9860 15.1640 ;
        RECT 5.1120 15.1160 5.1480 15.1640 ;
        RECT 5.8770 15.1160 5.8950 15.1640 ;
        RECT 9.4410 15.1160 9.4590 15.1640 ;
        RECT 0.1530 16.1960 0.1710 16.2440 ;
        RECT 3.7170 16.1960 3.7350 16.2440 ;
        RECT 4.9590 16.1960 4.9860 16.2440 ;
        RECT 5.1120 16.1960 5.1480 16.2440 ;
        RECT 5.8770 16.1960 5.8950 16.2440 ;
        RECT 9.4410 16.1960 9.4590 16.2440 ;
        RECT 0.1530 17.2760 0.1710 17.3240 ;
        RECT 3.7170 17.2760 3.7350 17.3240 ;
        RECT 4.9590 17.2760 4.9860 17.3240 ;
        RECT 5.1120 17.2760 5.1480 17.3240 ;
        RECT 5.8770 17.2760 5.8950 17.3240 ;
        RECT 9.4410 17.2760 9.4590 17.3240 ;
        RECT 0.1530 18.2910 0.1710 18.5070 ;
        RECT 4.9270 24.6270 4.9450 24.8430 ;
        RECT 4.9270 21.4590 4.9450 21.6750 ;
        RECT 4.9270 18.2910 4.9450 18.5070 ;
        RECT 4.9790 24.6270 4.9970 24.8430 ;
        RECT 4.9790 21.4590 4.9970 21.6750 ;
        RECT 4.9790 18.2910 4.9970 18.5070 ;
        RECT 5.0310 24.6270 5.0490 24.8430 ;
        RECT 5.0310 21.4590 5.0490 21.6750 ;
        RECT 5.0310 18.2910 5.0490 18.5070 ;
        RECT 5.0830 24.6270 5.1010 24.8430 ;
        RECT 5.0830 21.4590 5.1010 21.6750 ;
        RECT 5.0830 18.2910 5.1010 18.5070 ;
        RECT 5.1350 24.6270 5.1530 24.8430 ;
        RECT 5.1350 21.4590 5.1530 21.6750 ;
        RECT 5.1350 18.2910 5.1530 18.5070 ;
        RECT 0.1530 26.4830 0.1710 26.5310 ;
        RECT 3.7170 26.4830 3.7350 26.5310 ;
        RECT 4.9590 26.4830 4.9860 26.5310 ;
        RECT 5.1120 26.4830 5.1480 26.5310 ;
        RECT 5.8770 26.4830 5.8950 26.5310 ;
        RECT 9.4410 26.4830 9.4590 26.5310 ;
        RECT 0.1530 27.5630 0.1710 27.6110 ;
        RECT 3.7170 27.5630 3.7350 27.6110 ;
        RECT 4.9590 27.5630 4.9860 27.6110 ;
        RECT 5.1120 27.5630 5.1480 27.6110 ;
        RECT 5.8770 27.5630 5.8950 27.6110 ;
        RECT 9.4410 27.5630 9.4590 27.6110 ;
        RECT 0.1530 28.6430 0.1710 28.6910 ;
        RECT 3.7170 28.6430 3.7350 28.6910 ;
        RECT 4.9590 28.6430 4.9860 28.6910 ;
        RECT 5.1120 28.6430 5.1480 28.6910 ;
        RECT 5.8770 28.6430 5.8950 28.6910 ;
        RECT 9.4410 28.6430 9.4590 28.6910 ;
        RECT 0.1530 29.7230 0.1710 29.7710 ;
        RECT 3.7170 29.7230 3.7350 29.7710 ;
        RECT 4.9590 29.7230 4.9860 29.7710 ;
        RECT 5.1120 29.7230 5.1480 29.7710 ;
        RECT 5.8770 29.7230 5.8950 29.7710 ;
        RECT 9.4410 29.7230 9.4590 29.7710 ;
        RECT 0.1530 30.8030 0.1710 30.8510 ;
        RECT 3.7170 30.8030 3.7350 30.8510 ;
        RECT 4.9590 30.8030 4.9860 30.8510 ;
        RECT 5.1120 30.8030 5.1480 30.8510 ;
        RECT 5.8770 30.8030 5.8950 30.8510 ;
        RECT 9.4410 30.8030 9.4590 30.8510 ;
        RECT 0.1530 31.8830 0.1710 31.9310 ;
        RECT 3.7170 31.8830 3.7350 31.9310 ;
        RECT 4.9590 31.8830 4.9860 31.9310 ;
        RECT 5.1120 31.8830 5.1480 31.9310 ;
        RECT 5.8770 31.8830 5.8950 31.9310 ;
        RECT 9.4410 31.8830 9.4590 31.9310 ;
        RECT 0.1530 32.9630 0.1710 33.0110 ;
        RECT 3.7170 32.9630 3.7350 33.0110 ;
        RECT 4.9590 32.9630 4.9860 33.0110 ;
        RECT 5.1120 32.9630 5.1480 33.0110 ;
        RECT 5.8770 32.9630 5.8950 33.0110 ;
        RECT 9.4410 32.9630 9.4590 33.0110 ;
        RECT 0.1530 34.0430 0.1710 34.0910 ;
        RECT 3.7170 34.0430 3.7350 34.0910 ;
        RECT 4.9590 34.0430 4.9860 34.0910 ;
        RECT 5.1120 34.0430 5.1480 34.0910 ;
        RECT 5.8770 34.0430 5.8950 34.0910 ;
        RECT 9.4410 34.0430 9.4590 34.0910 ;
        RECT 0.1530 35.1230 0.1710 35.1710 ;
        RECT 3.7170 35.1230 3.7350 35.1710 ;
        RECT 4.9590 35.1230 4.9860 35.1710 ;
        RECT 5.1120 35.1230 5.1480 35.1710 ;
        RECT 5.8770 35.1230 5.8950 35.1710 ;
        RECT 9.4410 35.1230 9.4590 35.1710 ;
        RECT 0.1530 36.2030 0.1710 36.2510 ;
        RECT 3.7170 36.2030 3.7350 36.2510 ;
        RECT 4.9590 36.2030 4.9860 36.2510 ;
        RECT 5.1120 36.2030 5.1480 36.2510 ;
        RECT 5.8770 36.2030 5.8950 36.2510 ;
        RECT 9.4410 36.2030 9.4590 36.2510 ;
        RECT 0.1530 37.2830 0.1710 37.3310 ;
        RECT 3.7170 37.2830 3.7350 37.3310 ;
        RECT 4.9590 37.2830 4.9860 37.3310 ;
        RECT 5.1120 37.2830 5.1480 37.3310 ;
        RECT 5.8770 37.2830 5.8950 37.3310 ;
        RECT 9.4410 37.2830 9.4590 37.3310 ;
        RECT 0.1530 38.3630 0.1710 38.4110 ;
        RECT 3.7170 38.3630 3.7350 38.4110 ;
        RECT 4.9590 38.3630 4.9860 38.4110 ;
        RECT 5.1120 38.3630 5.1480 38.4110 ;
        RECT 5.8770 38.3630 5.8950 38.4110 ;
        RECT 9.4410 38.3630 9.4590 38.4110 ;
        RECT 0.1530 39.4430 0.1710 39.4910 ;
        RECT 3.7170 39.4430 3.7350 39.4910 ;
        RECT 4.9590 39.4430 4.9860 39.4910 ;
        RECT 5.1120 39.4430 5.1480 39.4910 ;
        RECT 5.8770 39.4430 5.8950 39.4910 ;
        RECT 9.4410 39.4430 9.4590 39.4910 ;
        RECT 0.1530 40.5230 0.1710 40.5710 ;
        RECT 3.7170 40.5230 3.7350 40.5710 ;
        RECT 4.9590 40.5230 4.9860 40.5710 ;
        RECT 5.1120 40.5230 5.1480 40.5710 ;
        RECT 5.8770 40.5230 5.8950 40.5710 ;
        RECT 9.4410 40.5230 9.4590 40.5710 ;
        RECT 0.1530 41.6030 0.1710 41.6510 ;
        RECT 3.7170 41.6030 3.7350 41.6510 ;
        RECT 4.9590 41.6030 4.9860 41.6510 ;
        RECT 5.1120 41.6030 5.1480 41.6510 ;
        RECT 5.8770 41.6030 5.8950 41.6510 ;
        RECT 9.4410 41.6030 9.4590 41.6510 ;
        RECT 0.1530 42.6830 0.1710 42.7310 ;
        RECT 3.7170 42.6830 3.7350 42.7310 ;
        RECT 4.9590 42.6830 4.9860 42.7310 ;
        RECT 5.1120 42.6830 5.1480 42.7310 ;
        RECT 5.8770 42.6830 5.8950 42.7310 ;
        RECT 9.4410 42.6830 9.4590 42.7310 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.3350 18.7630 7.3530 18.8000 ;
      LAYER M4  ;
        RECT 7.2830 18.7710 7.3670 18.7950 ;
      LAYER M5  ;
        RECT 7.3320 17.8200 7.3560 21.0600 ;
      LAYER V3  ;
        RECT 7.3350 18.7710 7.3530 18.7950 ;
      LAYER V4  ;
        RECT 7.3320 18.7710 7.3560 18.7950 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.1190 18.7660 7.1370 18.8030 ;
      LAYER M4  ;
        RECT 7.0670 18.7710 7.1510 18.7950 ;
      LAYER M5  ;
        RECT 7.1160 17.8200 7.1400 21.0600 ;
      LAYER V3  ;
        RECT 7.1190 18.7710 7.1370 18.7950 ;
      LAYER V4  ;
        RECT 7.1160 18.7710 7.1400 18.7950 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.9030 18.1870 6.9210 18.2240 ;
      LAYER M4  ;
        RECT 6.8510 18.1950 6.9350 18.2190 ;
      LAYER M5  ;
        RECT 6.9000 17.8200 6.9240 21.0600 ;
      LAYER V3  ;
        RECT 6.9030 18.1950 6.9210 18.2190 ;
      LAYER V4  ;
        RECT 6.9000 18.1950 6.9240 18.2190 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.6870 18.4270 6.7050 18.6080 ;
      LAYER M4  ;
        RECT 6.6350 18.5790 6.7190 18.6030 ;
      LAYER M5  ;
        RECT 6.6840 17.8200 6.7080 21.0600 ;
      LAYER V3  ;
        RECT 6.6870 18.5790 6.7050 18.6030 ;
      LAYER V4  ;
        RECT 6.6840 18.5790 6.7080 18.6030 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.4710 18.1900 6.4890 18.2570 ;
      LAYER M4  ;
        RECT 6.4190 18.1950 6.5030 18.2190 ;
      LAYER M5  ;
        RECT 6.4680 17.8200 6.4920 21.0600 ;
      LAYER V3  ;
        RECT 6.4710 18.1950 6.4890 18.2190 ;
      LAYER V4  ;
        RECT 6.4680 18.1950 6.4920 18.2190 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.2550 17.9230 6.2730 18.1760 ;
      LAYER M4  ;
        RECT 6.2030 18.1470 6.2870 18.1710 ;
      LAYER M5  ;
        RECT 6.2520 17.8200 6.2760 21.0600 ;
      LAYER V3  ;
        RECT 6.2550 18.1470 6.2730 18.1710 ;
      LAYER V4  ;
        RECT 6.2520 18.1470 6.2760 18.1710 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.0390 18.9580 6.0570 18.9950 ;
      LAYER M4  ;
        RECT 5.9870 18.9630 6.0710 18.9870 ;
      LAYER M5  ;
        RECT 6.0360 17.8200 6.0600 21.0600 ;
      LAYER V3  ;
        RECT 6.0390 18.9630 6.0570 18.9870 ;
      LAYER V4  ;
        RECT 6.0360 18.9630 6.0600 18.9870 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 5.1750 18.1900 5.1930 18.2570 ;
      LAYER M4  ;
        RECT 4.8910 18.1950 5.2040 18.2190 ;
      LAYER M5  ;
        RECT 4.9020 17.8200 4.9260 21.0600 ;
      LAYER V3  ;
        RECT 5.1750 18.1950 5.1930 18.2190 ;
      LAYER V4  ;
        RECT 4.9020 18.1950 4.9260 18.2190 ;
    END
  END ADDRESS[7]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 4.7790 17.9230 4.7970 18.1760 ;
      LAYER M4  ;
        RECT 4.5670 18.1470 4.8080 18.1710 ;
      LAYER M5  ;
        RECT 4.5780 17.8200 4.6020 21.0600 ;
      LAYER V3  ;
        RECT 4.7790 18.1470 4.7970 18.1710 ;
      LAYER V4  ;
        RECT 4.5780 18.1470 4.6020 18.1710 ;
    END
  END banksel
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.9870 18.1900 4.0050 18.2570 ;
      LAYER M4  ;
        RECT 3.9350 18.1950 4.0190 18.2190 ;
      LAYER M5  ;
        RECT 3.9840 17.8200 4.0080 21.0600 ;
      LAYER V3  ;
        RECT 3.9870 18.1950 4.0050 18.2190 ;
      LAYER V4  ;
        RECT 3.9840 18.1950 4.0080 18.2190 ;
    END
  END write
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.7710 19.0540 3.7890 19.1030 ;
      LAYER M4  ;
        RECT 3.7190 19.0590 3.8030 19.0830 ;
      LAYER M5  ;
        RECT 3.7680 17.8200 3.7920 21.0600 ;
      LAYER V3  ;
        RECT 3.7710 19.0590 3.7890 19.0830 ;
      LAYER V4  ;
        RECT 3.7680 19.0590 3.7920 19.0830 ;
    END
  END clk
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.8070 17.9230 3.8250 18.1760 ;
      LAYER M4  ;
        RECT 3.5410 18.1470 3.8360 18.1710 ;
      LAYER M5  ;
        RECT 3.5520 17.8200 3.5760 21.0600 ;
      LAYER V3  ;
        RECT 3.8070 18.1470 3.8250 18.1710 ;
      LAYER V4  ;
        RECT 3.5520 18.1470 3.5760 18.1710 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.3390 18.7630 3.3570 18.8000 ;
      LAYER M4  ;
        RECT 3.2870 18.7710 3.3710 18.7950 ;
      LAYER M5  ;
        RECT 3.3360 17.8200 3.3600 21.0600 ;
      LAYER V3  ;
        RECT 3.3390 18.7710 3.3570 18.7950 ;
      LAYER V4  ;
        RECT 3.3360 18.7710 3.3600 18.7950 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.1230 18.1900 3.1410 18.4190 ;
      LAYER M4  ;
        RECT 3.0710 18.1950 3.1550 18.2190 ;
      LAYER M5  ;
        RECT 3.1200 17.8200 3.1440 21.0600 ;
      LAYER V3  ;
        RECT 3.1230 18.1950 3.1410 18.2190 ;
      LAYER V4  ;
        RECT 3.1200 18.1950 3.1440 18.2190 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.9070 17.9230 2.9250 18.1760 ;
      LAYER M4  ;
        RECT 2.8550 18.1470 2.9390 18.1710 ;
      LAYER M5  ;
        RECT 2.9040 17.8200 2.9280 21.0600 ;
      LAYER V3  ;
        RECT 2.9070 18.1470 2.9250 18.1710 ;
      LAYER V4  ;
        RECT 2.9040 18.1470 2.9280 18.1710 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.6910 18.1870 2.7090 18.2240 ;
      LAYER M4  ;
        RECT 2.6390 18.1950 2.7230 18.2190 ;
      LAYER M5  ;
        RECT 2.6880 17.8200 2.7120 21.0600 ;
      LAYER V3  ;
        RECT 2.6910 18.1950 2.7090 18.2190 ;
      LAYER V4  ;
        RECT 2.6880 18.1950 2.7120 18.2190 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.4750 18.7630 2.4930 18.8000 ;
      LAYER M4  ;
        RECT 2.4230 18.7710 2.5070 18.7950 ;
      LAYER M5  ;
        RECT 2.4720 17.8200 2.4960 21.0600 ;
      LAYER V3  ;
        RECT 2.4750 18.7710 2.4930 18.7950 ;
      LAYER V4  ;
        RECT 2.4720 18.7710 2.4960 18.7950 ;
    END
  END sdel[4]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 0.4280 5.1360 0.4520 ;
      LAYER M3  ;
        RECT 5.0760 0.3775 5.0940 0.6170 ;
      LAYER V3  ;
        RECT 5.0760 0.4280 5.0940 0.4520 ;
    END
  END dataout[0]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 0.3320 5.2040 0.3560 ;
      LAYER M3  ;
        RECT 4.8510 0.2700 4.8690 0.6750 ;
      LAYER V3  ;
        RECT 4.8510 0.3320 4.8690 0.3560 ;
    END
  END wd[0]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 1.5080 5.1360 1.5320 ;
      LAYER M3  ;
        RECT 5.0760 1.4575 5.0940 1.6970 ;
      LAYER V3  ;
        RECT 5.0760 1.5080 5.0940 1.5320 ;
    END
  END dataout[1]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 1.4120 5.2040 1.4360 ;
      LAYER M3  ;
        RECT 4.8510 1.3500 4.8690 1.7550 ;
      LAYER V3  ;
        RECT 4.8510 1.4120 4.8690 1.4360 ;
    END
  END wd[1]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 2.5880 5.1360 2.6120 ;
      LAYER M3  ;
        RECT 5.0760 2.5375 5.0940 2.7770 ;
      LAYER V3  ;
        RECT 5.0760 2.5880 5.0940 2.6120 ;
    END
  END dataout[2]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 2.4920 5.2040 2.5160 ;
      LAYER M3  ;
        RECT 4.8510 2.4300 4.8690 2.8350 ;
      LAYER V3  ;
        RECT 4.8510 2.4920 4.8690 2.5160 ;
    END
  END wd[2]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 3.6680 5.1360 3.6920 ;
      LAYER M3  ;
        RECT 5.0760 3.6175 5.0940 3.8570 ;
      LAYER V3  ;
        RECT 5.0760 3.6680 5.0940 3.6920 ;
    END
  END dataout[3]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 3.5720 5.2040 3.5960 ;
      LAYER M3  ;
        RECT 4.8510 3.5100 4.8690 3.9150 ;
      LAYER V3  ;
        RECT 4.8510 3.5720 4.8690 3.5960 ;
    END
  END wd[3]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 4.7480 5.1360 4.7720 ;
      LAYER M3  ;
        RECT 5.0760 4.6975 5.0940 4.9370 ;
      LAYER V3  ;
        RECT 5.0760 4.7480 5.0940 4.7720 ;
    END
  END dataout[4]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 4.6520 5.2040 4.6760 ;
      LAYER M3  ;
        RECT 4.8510 4.5900 4.8690 4.9950 ;
      LAYER V3  ;
        RECT 4.8510 4.6520 4.8690 4.6760 ;
    END
  END wd[4]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 5.8280 5.1360 5.8520 ;
      LAYER M3  ;
        RECT 5.0760 5.7775 5.0940 6.0170 ;
      LAYER V3  ;
        RECT 5.0760 5.8280 5.0940 5.8520 ;
    END
  END dataout[5]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 5.7320 5.2040 5.7560 ;
      LAYER M3  ;
        RECT 4.8510 5.6700 4.8690 6.0750 ;
      LAYER V3  ;
        RECT 4.8510 5.7320 4.8690 5.7560 ;
    END
  END wd[5]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 6.9080 5.1360 6.9320 ;
      LAYER M3  ;
        RECT 5.0760 6.8575 5.0940 7.0970 ;
      LAYER V3  ;
        RECT 5.0760 6.9080 5.0940 6.9320 ;
    END
  END dataout[6]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 6.8120 5.2040 6.8360 ;
      LAYER M3  ;
        RECT 4.8510 6.7500 4.8690 7.1550 ;
      LAYER V3  ;
        RECT 4.8510 6.8120 4.8690 6.8360 ;
    END
  END wd[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 7.9880 5.1360 8.0120 ;
      LAYER M3  ;
        RECT 5.0760 7.9375 5.0940 8.1770 ;
      LAYER V3  ;
        RECT 5.0760 7.9880 5.0940 8.0120 ;
    END
  END dataout[7]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 7.8920 5.2040 7.9160 ;
      LAYER M3  ;
        RECT 4.8510 7.8300 4.8690 8.2350 ;
      LAYER V3  ;
        RECT 4.8510 7.8920 4.8690 7.9160 ;
    END
  END wd[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 9.0680 5.1360 9.0920 ;
      LAYER M3  ;
        RECT 5.0760 9.0175 5.0940 9.2570 ;
      LAYER V3  ;
        RECT 5.0760 9.0680 5.0940 9.0920 ;
    END
  END dataout[8]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 8.9720 5.2040 8.9960 ;
      LAYER M3  ;
        RECT 4.8510 8.9100 4.8690 9.3150 ;
      LAYER V3  ;
        RECT 4.8510 8.9720 4.8690 8.9960 ;
    END
  END wd[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 10.1480 5.1360 10.1720 ;
      LAYER M3  ;
        RECT 5.0760 10.0975 5.0940 10.3370 ;
      LAYER V3  ;
        RECT 5.0760 10.1480 5.0940 10.1720 ;
    END
  END dataout[9]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 10.0520 5.2040 10.0760 ;
      LAYER M3  ;
        RECT 4.8510 9.9900 4.8690 10.3950 ;
      LAYER V3  ;
        RECT 4.8510 10.0520 4.8690 10.0760 ;
    END
  END wd[9]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 11.2280 5.1360 11.2520 ;
      LAYER M3  ;
        RECT 5.0760 11.1775 5.0940 11.4170 ;
      LAYER V3  ;
        RECT 5.0760 11.2280 5.0940 11.2520 ;
    END
  END dataout[10]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 11.1320 5.2040 11.1560 ;
      LAYER M3  ;
        RECT 4.8510 11.0700 4.8690 11.4750 ;
      LAYER V3  ;
        RECT 4.8510 11.1320 4.8690 11.1560 ;
    END
  END wd[10]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 12.3080 5.1360 12.3320 ;
      LAYER M3  ;
        RECT 5.0760 12.2575 5.0940 12.4970 ;
      LAYER V3  ;
        RECT 5.0760 12.3080 5.0940 12.3320 ;
    END
  END dataout[11]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 12.2120 5.2040 12.2360 ;
      LAYER M3  ;
        RECT 4.8510 12.1500 4.8690 12.5550 ;
      LAYER V3  ;
        RECT 4.8510 12.2120 4.8690 12.2360 ;
    END
  END wd[11]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 13.3880 5.1360 13.4120 ;
      LAYER M3  ;
        RECT 5.0760 13.3375 5.0940 13.5770 ;
      LAYER V3  ;
        RECT 5.0760 13.3880 5.0940 13.4120 ;
    END
  END dataout[12]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 13.2920 5.2040 13.3160 ;
      LAYER M3  ;
        RECT 4.8510 13.2300 4.8690 13.6350 ;
      LAYER V3  ;
        RECT 4.8510 13.2920 4.8690 13.3160 ;
    END
  END wd[12]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 14.4680 5.1360 14.4920 ;
      LAYER M3  ;
        RECT 5.0760 14.4175 5.0940 14.6570 ;
      LAYER V3  ;
        RECT 5.0760 14.4680 5.0940 14.4920 ;
    END
  END dataout[13]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 14.3720 5.2040 14.3960 ;
      LAYER M3  ;
        RECT 4.8510 14.3100 4.8690 14.7150 ;
      LAYER V3  ;
        RECT 4.8510 14.3720 4.8690 14.3960 ;
    END
  END wd[13]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 15.5480 5.1360 15.5720 ;
      LAYER M3  ;
        RECT 5.0760 15.4975 5.0940 15.7370 ;
      LAYER V3  ;
        RECT 5.0760 15.5480 5.0940 15.5720 ;
    END
  END dataout[14]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 15.4520 5.2040 15.4760 ;
      LAYER M3  ;
        RECT 4.8510 15.3900 4.8690 15.7950 ;
      LAYER V3  ;
        RECT 4.8510 15.4520 4.8690 15.4760 ;
    END
  END wd[14]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 16.6280 5.1360 16.6520 ;
      LAYER M3  ;
        RECT 5.0760 16.5775 5.0940 16.8170 ;
      LAYER V3  ;
        RECT 5.0760 16.6280 5.0940 16.6520 ;
    END
  END dataout[15]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 16.5320 5.2040 16.5560 ;
      LAYER M3  ;
        RECT 4.8510 16.4700 4.8690 16.8750 ;
      LAYER V3  ;
        RECT 4.8510 16.5320 4.8690 16.5560 ;
    END
  END wd[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 25.8350 5.1360 25.8590 ;
      LAYER M3  ;
        RECT 5.0760 25.7845 5.0940 26.0240 ;
      LAYER V3  ;
        RECT 5.0760 25.8350 5.0940 25.8590 ;
    END
  END dataout[16]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 25.7390 5.2040 25.7630 ;
      LAYER M3  ;
        RECT 4.8510 25.6770 4.8690 26.0820 ;
      LAYER V3  ;
        RECT 4.8510 25.7390 4.8690 25.7630 ;
    END
  END wd[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 26.9150 5.1360 26.9390 ;
      LAYER M3  ;
        RECT 5.0760 26.8645 5.0940 27.1040 ;
      LAYER V3  ;
        RECT 5.0760 26.9150 5.0940 26.9390 ;
    END
  END dataout[17]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 26.8190 5.2040 26.8430 ;
      LAYER M3  ;
        RECT 4.8510 26.7570 4.8690 27.1620 ;
      LAYER V3  ;
        RECT 4.8510 26.8190 4.8690 26.8430 ;
    END
  END wd[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 27.9950 5.1360 28.0190 ;
      LAYER M3  ;
        RECT 5.0760 27.9445 5.0940 28.1840 ;
      LAYER V3  ;
        RECT 5.0760 27.9950 5.0940 28.0190 ;
    END
  END dataout[18]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 27.8990 5.2040 27.9230 ;
      LAYER M3  ;
        RECT 4.8510 27.8370 4.8690 28.2420 ;
      LAYER V3  ;
        RECT 4.8510 27.8990 4.8690 27.9230 ;
    END
  END wd[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 29.0750 5.1360 29.0990 ;
      LAYER M3  ;
        RECT 5.0760 29.0245 5.0940 29.2640 ;
      LAYER V3  ;
        RECT 5.0760 29.0750 5.0940 29.0990 ;
    END
  END dataout[19]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 28.9790 5.2040 29.0030 ;
      LAYER M3  ;
        RECT 4.8510 28.9170 4.8690 29.3220 ;
      LAYER V3  ;
        RECT 4.8510 28.9790 4.8690 29.0030 ;
    END
  END wd[19]
  PIN dataout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 30.1550 5.1360 30.1790 ;
      LAYER M3  ;
        RECT 5.0760 30.1045 5.0940 30.3440 ;
      LAYER V3  ;
        RECT 5.0760 30.1550 5.0940 30.1790 ;
    END
  END dataout[20]
  PIN wd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 30.0590 5.2040 30.0830 ;
      LAYER M3  ;
        RECT 4.8510 29.9970 4.8690 30.4020 ;
      LAYER V3  ;
        RECT 4.8510 30.0590 4.8690 30.0830 ;
    END
  END wd[20]
  PIN dataout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 31.2350 5.1360 31.2590 ;
      LAYER M3  ;
        RECT 5.0760 31.1845 5.0940 31.4240 ;
      LAYER V3  ;
        RECT 5.0760 31.2350 5.0940 31.2590 ;
    END
  END dataout[21]
  PIN wd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 31.1390 5.2040 31.1630 ;
      LAYER M3  ;
        RECT 4.8510 31.0770 4.8690 31.4820 ;
      LAYER V3  ;
        RECT 4.8510 31.1390 4.8690 31.1630 ;
    END
  END wd[21]
  PIN dataout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 32.3150 5.1360 32.3390 ;
      LAYER M3  ;
        RECT 5.0760 32.2645 5.0940 32.5040 ;
      LAYER V3  ;
        RECT 5.0760 32.3150 5.0940 32.3390 ;
    END
  END dataout[22]
  PIN wd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 32.2190 5.2040 32.2430 ;
      LAYER M3  ;
        RECT 4.8510 32.1570 4.8690 32.5620 ;
      LAYER V3  ;
        RECT 4.8510 32.2190 4.8690 32.2430 ;
    END
  END wd[22]
  PIN dataout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 33.3950 5.1360 33.4190 ;
      LAYER M3  ;
        RECT 5.0760 33.3445 5.0940 33.5840 ;
      LAYER V3  ;
        RECT 5.0760 33.3950 5.0940 33.4190 ;
    END
  END dataout[23]
  PIN wd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 33.2990 5.2040 33.3230 ;
      LAYER M3  ;
        RECT 4.8510 33.2370 4.8690 33.6420 ;
      LAYER V3  ;
        RECT 4.8510 33.2990 4.8690 33.3230 ;
    END
  END wd[23]
  PIN dataout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 34.4750 5.1360 34.4990 ;
      LAYER M3  ;
        RECT 5.0760 34.4245 5.0940 34.6640 ;
      LAYER V3  ;
        RECT 5.0760 34.4750 5.0940 34.4990 ;
    END
  END dataout[24]
  PIN wd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 34.3790 5.2040 34.4030 ;
      LAYER M3  ;
        RECT 4.8510 34.3170 4.8690 34.7220 ;
      LAYER V3  ;
        RECT 4.8510 34.3790 4.8690 34.4030 ;
    END
  END wd[24]
  PIN dataout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 35.5550 5.1360 35.5790 ;
      LAYER M3  ;
        RECT 5.0760 35.5045 5.0940 35.7440 ;
      LAYER V3  ;
        RECT 5.0760 35.5550 5.0940 35.5790 ;
    END
  END dataout[25]
  PIN wd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 35.4590 5.2040 35.4830 ;
      LAYER M3  ;
        RECT 4.8510 35.3970 4.8690 35.8020 ;
      LAYER V3  ;
        RECT 4.8510 35.4590 4.8690 35.4830 ;
    END
  END wd[25]
  PIN dataout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 36.6350 5.1360 36.6590 ;
      LAYER M3  ;
        RECT 5.0760 36.5845 5.0940 36.8240 ;
      LAYER V3  ;
        RECT 5.0760 36.6350 5.0940 36.6590 ;
    END
  END dataout[26]
  PIN wd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 36.5390 5.2040 36.5630 ;
      LAYER M3  ;
        RECT 4.8510 36.4770 4.8690 36.8820 ;
      LAYER V3  ;
        RECT 4.8510 36.5390 4.8690 36.5630 ;
    END
  END wd[26]
  PIN dataout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 37.7150 5.1360 37.7390 ;
      LAYER M3  ;
        RECT 5.0760 37.6645 5.0940 37.9040 ;
      LAYER V3  ;
        RECT 5.0760 37.7150 5.0940 37.7390 ;
    END
  END dataout[27]
  PIN wd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 37.6190 5.2040 37.6430 ;
      LAYER M3  ;
        RECT 4.8510 37.5570 4.8690 37.9620 ;
      LAYER V3  ;
        RECT 4.8510 37.6190 4.8690 37.6430 ;
    END
  END wd[27]
  PIN dataout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 38.7950 5.1360 38.8190 ;
      LAYER M3  ;
        RECT 5.0760 38.7445 5.0940 38.9840 ;
      LAYER V3  ;
        RECT 5.0760 38.7950 5.0940 38.8190 ;
    END
  END dataout[28]
  PIN wd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 38.6990 5.2040 38.7230 ;
      LAYER M3  ;
        RECT 4.8510 38.6370 4.8690 39.0420 ;
      LAYER V3  ;
        RECT 4.8510 38.6990 4.8690 38.7230 ;
    END
  END wd[28]
  PIN dataout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 39.8750 5.1360 39.8990 ;
      LAYER M3  ;
        RECT 5.0760 39.8245 5.0940 40.0640 ;
      LAYER V3  ;
        RECT 5.0760 39.8750 5.0940 39.8990 ;
    END
  END dataout[29]
  PIN wd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 39.7790 5.2040 39.8030 ;
      LAYER M3  ;
        RECT 4.8510 39.7170 4.8690 40.1220 ;
      LAYER V3  ;
        RECT 4.8510 39.7790 4.8690 39.8030 ;
    END
  END wd[29]
  PIN dataout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 40.9550 5.1360 40.9790 ;
      LAYER M3  ;
        RECT 5.0760 40.9045 5.0940 41.1440 ;
      LAYER V3  ;
        RECT 5.0760 40.9550 5.0940 40.9790 ;
    END
  END dataout[30]
  PIN wd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 40.8590 5.2040 40.8830 ;
      LAYER M3  ;
        RECT 4.8510 40.7970 4.8690 41.2020 ;
      LAYER V3  ;
        RECT 4.8510 40.8590 4.8690 40.8830 ;
    END
  END wd[30]
  PIN dataout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 42.0350 5.1360 42.0590 ;
      LAYER M3  ;
        RECT 5.0760 41.9845 5.0940 42.2240 ;
      LAYER V3  ;
        RECT 5.0760 42.0350 5.0940 42.0590 ;
    END
  END dataout[31]
  PIN wd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 41.9390 5.2040 41.9630 ;
      LAYER M3  ;
        RECT 4.8510 41.8770 4.8690 42.2820 ;
      LAYER V3  ;
        RECT 4.8510 41.9390 4.8690 41.9630 ;
    END
  END wd[31]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5230 9.6120 26.1765 ;
        RECT 0.0000 25.6635 9.6120 26.7570 ;
        RECT 0.0000 26.7435 9.6120 27.8370 ;
        RECT 0.0000 27.8235 9.6120 28.9170 ;
        RECT 0.0000 28.9035 9.6120 29.9970 ;
        RECT 0.0000 29.9835 9.6120 31.0770 ;
        RECT 0.0000 31.0635 9.6120 32.1570 ;
        RECT 0.0000 32.1435 9.6120 33.2370 ;
        RECT 0.0000 33.2235 9.6120 34.3170 ;
        RECT 0.0000 34.3035 9.6120 35.3970 ;
        RECT 0.0000 35.3835 9.6120 36.4770 ;
        RECT 0.0000 36.4635 9.6120 37.5570 ;
        RECT 0.0000 37.5435 9.6120 38.6370 ;
        RECT 0.0000 38.6235 9.6120 39.7170 ;
        RECT 0.0000 39.7035 9.6120 40.7970 ;
        RECT 0.0000 40.7835 9.6120 41.8770 ;
        RECT 0.0000 41.8635 9.6120 42.9570 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5230 9.6120 26.1765 ;
        RECT 0.0000 25.6635 9.6120 26.7570 ;
        RECT 0.0000 26.7435 9.6120 27.8370 ;
        RECT 0.0000 27.8235 9.6120 28.9170 ;
        RECT 0.0000 28.9035 9.6120 29.9970 ;
        RECT 0.0000 29.9835 9.6120 31.0770 ;
        RECT 0.0000 31.0635 9.6120 32.1570 ;
        RECT 0.0000 32.1435 9.6120 33.2370 ;
        RECT 0.0000 33.2235 9.6120 34.3170 ;
        RECT 0.0000 34.3035 9.6120 35.3970 ;
        RECT 0.0000 35.3835 9.6120 36.4770 ;
        RECT 0.0000 36.4635 9.6120 37.5570 ;
        RECT 0.0000 37.5435 9.6120 38.6370 ;
        RECT 0.0000 38.6235 9.6120 39.7170 ;
        RECT 0.0000 39.7035 9.6120 40.7970 ;
        RECT 0.0000 40.7835 9.6120 41.8770 ;
        RECT 0.0000 41.8635 9.6120 42.9570 ;
  LAYER V1  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5230 9.6120 26.1765 ;
        RECT 0.0000 25.6635 9.6120 26.7570 ;
        RECT 0.0000 26.7435 9.6120 27.8370 ;
        RECT 0.0000 27.8235 9.6120 28.9170 ;
        RECT 0.0000 28.9035 9.6120 29.9970 ;
        RECT 0.0000 29.9835 9.6120 31.0770 ;
        RECT 0.0000 31.0635 9.6120 32.1570 ;
        RECT 0.0000 32.1435 9.6120 33.2370 ;
        RECT 0.0000 33.2235 9.6120 34.3170 ;
        RECT 0.0000 34.3035 9.6120 35.3970 ;
        RECT 0.0000 35.3835 9.6120 36.4770 ;
        RECT 0.0000 36.4635 9.6120 37.5570 ;
        RECT 0.0000 37.5435 9.6120 38.6370 ;
        RECT 0.0000 38.6235 9.6120 39.7170 ;
        RECT 0.0000 39.7035 9.6120 40.7970 ;
        RECT 0.0000 40.7835 9.6120 41.8770 ;
        RECT 0.0000 41.8635 9.6120 42.9570 ;
  LAYER V2  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5230 9.6120 26.1765 ;
        RECT 0.0000 25.6635 9.6120 26.7570 ;
        RECT 0.0000 26.7435 9.6120 27.8370 ;
        RECT 0.0000 27.8235 9.6120 28.9170 ;
        RECT 0.0000 28.9035 9.6120 29.9970 ;
        RECT 0.0000 29.9835 9.6120 31.0770 ;
        RECT 0.0000 31.0635 9.6120 32.1570 ;
        RECT 0.0000 32.1435 9.6120 33.2370 ;
        RECT 0.0000 33.2235 9.6120 34.3170 ;
        RECT 0.0000 34.3035 9.6120 35.3970 ;
        RECT 0.0000 35.3835 9.6120 36.4770 ;
        RECT 0.0000 36.4635 9.6120 37.5570 ;
        RECT 0.0000 37.5435 9.6120 38.6370 ;
        RECT 0.0000 38.6235 9.6120 39.7170 ;
        RECT 0.0000 39.7035 9.6120 40.7970 ;
        RECT 0.0000 40.7835 9.6120 41.8770 ;
        RECT 0.0000 41.8635 9.6120 42.9570 ;
  LAYER M3  ;
      RECT 5.2380 0.3450 5.2560 1.2805 ;
      RECT 5.2020 0.3450 5.2200 1.2805 ;
      RECT 5.1660 0.9220 5.1840 1.2445 ;
      RECT 5.0490 1.1190 5.0670 1.2285 ;
      RECT 5.0400 0.3775 5.0580 0.6170 ;
      RECT 5.0040 0.9585 5.0220 1.1120 ;
      RECT 4.9230 0.9840 4.9410 1.2420 ;
      RECT 4.3830 0.3450 4.4010 1.2805 ;
      RECT 4.3470 0.3450 4.3650 1.2805 ;
      RECT 4.3110 0.5260 4.3290 1.0940 ;
      RECT 5.2380 1.4250 5.2560 2.3605 ;
      RECT 5.2020 1.4250 5.2200 2.3605 ;
      RECT 5.1660 2.0020 5.1840 2.3245 ;
      RECT 5.0490 2.1990 5.0670 2.3085 ;
      RECT 5.0400 1.4575 5.0580 1.6970 ;
      RECT 5.0040 2.0385 5.0220 2.1920 ;
      RECT 4.9230 2.0640 4.9410 2.3220 ;
      RECT 4.3830 1.4250 4.4010 2.3605 ;
      RECT 4.3470 1.4250 4.3650 2.3605 ;
      RECT 4.3110 1.6060 4.3290 2.1740 ;
      RECT 5.2380 2.5050 5.2560 3.4405 ;
      RECT 5.2020 2.5050 5.2200 3.4405 ;
      RECT 5.1660 3.0820 5.1840 3.4045 ;
      RECT 5.0490 3.2790 5.0670 3.3885 ;
      RECT 5.0400 2.5375 5.0580 2.7770 ;
      RECT 5.0040 3.1185 5.0220 3.2720 ;
      RECT 4.9230 3.1440 4.9410 3.4020 ;
      RECT 4.3830 2.5050 4.4010 3.4405 ;
      RECT 4.3470 2.5050 4.3650 3.4405 ;
      RECT 4.3110 2.6860 4.3290 3.2540 ;
      RECT 5.2380 3.5850 5.2560 4.5205 ;
      RECT 5.2020 3.5850 5.2200 4.5205 ;
      RECT 5.1660 4.1620 5.1840 4.4845 ;
      RECT 5.0490 4.3590 5.0670 4.4685 ;
      RECT 5.0400 3.6175 5.0580 3.8570 ;
      RECT 5.0040 4.1985 5.0220 4.3520 ;
      RECT 4.9230 4.2240 4.9410 4.4820 ;
      RECT 4.3830 3.5850 4.4010 4.5205 ;
      RECT 4.3470 3.5850 4.3650 4.5205 ;
      RECT 4.3110 3.7660 4.3290 4.3340 ;
      RECT 5.2380 4.6650 5.2560 5.6005 ;
      RECT 5.2020 4.6650 5.2200 5.6005 ;
      RECT 5.1660 5.2420 5.1840 5.5645 ;
      RECT 5.0490 5.4390 5.0670 5.5485 ;
      RECT 5.0400 4.6975 5.0580 4.9370 ;
      RECT 5.0040 5.2785 5.0220 5.4320 ;
      RECT 4.9230 5.3040 4.9410 5.5620 ;
      RECT 4.3830 4.6650 4.4010 5.6005 ;
      RECT 4.3470 4.6650 4.3650 5.6005 ;
      RECT 4.3110 4.8460 4.3290 5.4140 ;
      RECT 5.2380 5.7450 5.2560 6.6805 ;
      RECT 5.2020 5.7450 5.2200 6.6805 ;
      RECT 5.1660 6.3220 5.1840 6.6445 ;
      RECT 5.0490 6.5190 5.0670 6.6285 ;
      RECT 5.0400 5.7775 5.0580 6.0170 ;
      RECT 5.0040 6.3585 5.0220 6.5120 ;
      RECT 4.9230 6.3840 4.9410 6.6420 ;
      RECT 4.3830 5.7450 4.4010 6.6805 ;
      RECT 4.3470 5.7450 4.3650 6.6805 ;
      RECT 4.3110 5.9260 4.3290 6.4940 ;
      RECT 5.2380 6.8250 5.2560 7.7605 ;
      RECT 5.2020 6.8250 5.2200 7.7605 ;
      RECT 5.1660 7.4020 5.1840 7.7245 ;
      RECT 5.0490 7.5990 5.0670 7.7085 ;
      RECT 5.0400 6.8575 5.0580 7.0970 ;
      RECT 5.0040 7.4385 5.0220 7.5920 ;
      RECT 4.9230 7.4640 4.9410 7.7220 ;
      RECT 4.3830 6.8250 4.4010 7.7605 ;
      RECT 4.3470 6.8250 4.3650 7.7605 ;
      RECT 4.3110 7.0060 4.3290 7.5740 ;
      RECT 5.2380 7.9050 5.2560 8.8405 ;
      RECT 5.2020 7.9050 5.2200 8.8405 ;
      RECT 5.1660 8.4820 5.1840 8.8045 ;
      RECT 5.0490 8.6790 5.0670 8.7885 ;
      RECT 5.0400 7.9375 5.0580 8.1770 ;
      RECT 5.0040 8.5185 5.0220 8.6720 ;
      RECT 4.9230 8.5440 4.9410 8.8020 ;
      RECT 4.3830 7.9050 4.4010 8.8405 ;
      RECT 4.3470 7.9050 4.3650 8.8405 ;
      RECT 4.3110 8.0860 4.3290 8.6540 ;
      RECT 5.2380 8.9850 5.2560 9.9205 ;
      RECT 5.2020 8.9850 5.2200 9.9205 ;
      RECT 5.1660 9.5620 5.1840 9.8845 ;
      RECT 5.0490 9.7590 5.0670 9.8685 ;
      RECT 5.0400 9.0175 5.0580 9.2570 ;
      RECT 5.0040 9.5985 5.0220 9.7520 ;
      RECT 4.9230 9.6240 4.9410 9.8820 ;
      RECT 4.3830 8.9850 4.4010 9.9205 ;
      RECT 4.3470 8.9850 4.3650 9.9205 ;
      RECT 4.3110 9.1660 4.3290 9.7340 ;
      RECT 5.2380 10.0650 5.2560 11.0005 ;
      RECT 5.2020 10.0650 5.2200 11.0005 ;
      RECT 5.1660 10.6420 5.1840 10.9645 ;
      RECT 5.0490 10.8390 5.0670 10.9485 ;
      RECT 5.0400 10.0975 5.0580 10.3370 ;
      RECT 5.0040 10.6785 5.0220 10.8320 ;
      RECT 4.9230 10.7040 4.9410 10.9620 ;
      RECT 4.3830 10.0650 4.4010 11.0005 ;
      RECT 4.3470 10.0650 4.3650 11.0005 ;
      RECT 4.3110 10.2460 4.3290 10.8140 ;
      RECT 5.2380 11.1450 5.2560 12.0805 ;
      RECT 5.2020 11.1450 5.2200 12.0805 ;
      RECT 5.1660 11.7220 5.1840 12.0445 ;
      RECT 5.0490 11.9190 5.0670 12.0285 ;
      RECT 5.0400 11.1775 5.0580 11.4170 ;
      RECT 5.0040 11.7585 5.0220 11.9120 ;
      RECT 4.9230 11.7840 4.9410 12.0420 ;
      RECT 4.3830 11.1450 4.4010 12.0805 ;
      RECT 4.3470 11.1450 4.3650 12.0805 ;
      RECT 4.3110 11.3260 4.3290 11.8940 ;
      RECT 5.2380 12.2250 5.2560 13.1605 ;
      RECT 5.2020 12.2250 5.2200 13.1605 ;
      RECT 5.1660 12.8020 5.1840 13.1245 ;
      RECT 5.0490 12.9990 5.0670 13.1085 ;
      RECT 5.0400 12.2575 5.0580 12.4970 ;
      RECT 5.0040 12.8385 5.0220 12.9920 ;
      RECT 4.9230 12.8640 4.9410 13.1220 ;
      RECT 4.3830 12.2250 4.4010 13.1605 ;
      RECT 4.3470 12.2250 4.3650 13.1605 ;
      RECT 4.3110 12.4060 4.3290 12.9740 ;
      RECT 5.2380 13.3050 5.2560 14.2405 ;
      RECT 5.2020 13.3050 5.2200 14.2405 ;
      RECT 5.1660 13.8820 5.1840 14.2045 ;
      RECT 5.0490 14.0790 5.0670 14.1885 ;
      RECT 5.0400 13.3375 5.0580 13.5770 ;
      RECT 5.0040 13.9185 5.0220 14.0720 ;
      RECT 4.9230 13.9440 4.9410 14.2020 ;
      RECT 4.3830 13.3050 4.4010 14.2405 ;
      RECT 4.3470 13.3050 4.3650 14.2405 ;
      RECT 4.3110 13.4860 4.3290 14.0540 ;
      RECT 5.2380 14.3850 5.2560 15.3205 ;
      RECT 5.2020 14.3850 5.2200 15.3205 ;
      RECT 5.1660 14.9620 5.1840 15.2845 ;
      RECT 5.0490 15.1590 5.0670 15.2685 ;
      RECT 5.0400 14.4175 5.0580 14.6570 ;
      RECT 5.0040 14.9985 5.0220 15.1520 ;
      RECT 4.9230 15.0240 4.9410 15.2820 ;
      RECT 4.3830 14.3850 4.4010 15.3205 ;
      RECT 4.3470 14.3850 4.3650 15.3205 ;
      RECT 4.3110 14.5660 4.3290 15.1340 ;
      RECT 5.2380 15.4650 5.2560 16.4005 ;
      RECT 5.2020 15.4650 5.2200 16.4005 ;
      RECT 5.1660 16.0420 5.1840 16.3645 ;
      RECT 5.0490 16.2390 5.0670 16.3485 ;
      RECT 5.0400 15.4975 5.0580 15.7370 ;
      RECT 5.0040 16.0785 5.0220 16.2320 ;
      RECT 4.9230 16.1040 4.9410 16.3620 ;
      RECT 4.3830 15.4650 4.4010 16.4005 ;
      RECT 4.3470 15.4650 4.3650 16.4005 ;
      RECT 4.3110 15.6460 4.3290 16.2140 ;
      RECT 5.2380 16.5450 5.2560 17.4805 ;
      RECT 5.2020 16.5450 5.2200 17.4805 ;
      RECT 5.1660 17.1220 5.1840 17.4445 ;
      RECT 5.0490 17.3190 5.0670 17.4285 ;
      RECT 5.0400 16.5775 5.0580 16.8170 ;
      RECT 5.0040 17.1585 5.0220 17.3120 ;
      RECT 4.9230 17.1840 4.9410 17.4420 ;
      RECT 4.3830 16.5450 4.4010 17.4805 ;
      RECT 4.3470 16.5450 4.3650 17.4805 ;
      RECT 4.3110 16.7260 4.3290 17.2940 ;
      RECT 9.4050 21.3160 9.4230 25.6715 ;
      RECT 9.3690 20.0010 9.3870 20.0700 ;
      RECT 9.3690 21.8090 9.3870 22.2735 ;
      RECT 9.3330 17.4965 9.3510 25.7035 ;
      RECT 9.2970 21.2660 9.3150 22.0385 ;
      RECT 9.2970 22.0897 9.3150 22.5810 ;
      RECT 9.2970 22.6310 9.3150 23.0025 ;
      RECT 9.2970 23.0655 9.3150 23.8770 ;
      RECT 9.2610 21.3515 9.2790 21.9935 ;
      RECT 9.2610 22.6710 9.2790 23.2030 ;
      RECT 9.2250 17.4965 9.2430 17.8465 ;
      RECT 9.1170 17.4965 9.1350 17.8465 ;
      RECT 9.0090 17.4965 9.0270 17.8465 ;
      RECT 8.9010 17.4965 8.9190 17.8465 ;
      RECT 8.7930 17.4965 8.8110 17.8465 ;
      RECT 8.6850 17.4965 8.7030 17.8465 ;
      RECT 8.5770 17.4965 8.5950 17.8465 ;
      RECT 8.4690 17.4965 8.4870 17.8465 ;
      RECT 8.3610 17.4965 8.3790 17.8465 ;
      RECT 8.2530 17.4965 8.2710 17.8465 ;
      RECT 8.1450 17.4965 8.1630 17.8465 ;
      RECT 8.0370 17.4965 8.0550 17.8465 ;
      RECT 7.9290 17.4965 7.9470 17.8465 ;
      RECT 7.8210 17.4965 7.8390 17.8465 ;
      RECT 7.7130 17.4965 7.7310 17.8465 ;
      RECT 7.6050 17.4965 7.6230 17.8465 ;
      RECT 7.4970 17.4965 7.5150 17.8465 ;
      RECT 7.3890 17.4965 7.4070 17.8465 ;
      RECT 7.2810 17.4965 7.2990 17.8465 ;
      RECT 7.1730 17.4965 7.1910 17.8465 ;
      RECT 7.0650 17.4965 7.0830 17.8465 ;
      RECT 6.9570 17.4965 6.9750 17.8465 ;
      RECT 6.8490 17.4965 6.8670 17.8465 ;
      RECT 6.7410 17.4965 6.7590 17.8465 ;
      RECT 6.6330 17.4965 6.6510 17.8465 ;
      RECT 6.5250 17.4965 6.5430 17.8465 ;
      RECT 6.4170 17.4965 6.4350 17.8465 ;
      RECT 6.3090 17.4965 6.3270 17.8465 ;
      RECT 6.2010 17.4965 6.2190 17.8465 ;
      RECT 6.0930 17.4965 6.1110 17.8465 ;
      RECT 6.0570 21.2850 6.0750 21.9897 ;
      RECT 6.0570 22.7320 6.0750 23.9130 ;
      RECT 6.0390 18.1570 6.0570 18.8330 ;
      RECT 6.0390 19.5790 6.0570 19.8770 ;
      RECT 6.0210 21.3485 6.0390 22.0385 ;
      RECT 6.0210 22.0895 6.0390 23.0810 ;
      RECT 6.0210 23.1110 6.0390 23.8950 ;
      RECT 5.9850 17.4965 6.0030 25.7035 ;
      RECT 5.9490 21.6210 5.9670 21.7040 ;
      RECT 5.9310 18.2650 5.9490 18.8960 ;
      RECT 5.9310 19.3090 5.9490 19.4990 ;
      RECT 5.9310 20.1910 5.9490 20.2400 ;
      RECT 5.9130 21.3160 5.9310 25.6760 ;
      RECT 5.8230 17.8870 5.8410 18.6890 ;
      RECT 5.8230 19.2370 5.8410 19.8050 ;
      RECT 5.7870 19.3090 5.8050 19.6790 ;
      RECT 5.7510 18.6610 5.7690 18.7970 ;
      RECT 5.7510 19.6510 5.7690 19.8770 ;
      RECT 5.7510 20.8930 5.7690 20.9570 ;
      RECT 5.7150 18.7630 5.7330 18.8000 ;
      RECT 5.7150 20.3890 5.7330 20.4320 ;
      RECT 5.7150 20.9230 5.7330 20.9600 ;
      RECT 5.6790 19.0750 5.6970 19.5710 ;
      RECT 5.6790 19.6150 5.6970 19.8050 ;
      RECT 5.6790 20.5750 5.6970 20.8850 ;
      RECT 5.6430 22.8550 5.6610 23.5850 ;
      RECT 5.6430 23.9350 5.6610 24.6650 ;
      RECT 5.3190 18.6970 5.3370 18.9950 ;
      RECT 5.3190 19.8850 5.3370 19.9490 ;
      RECT 5.3190 20.1550 5.3370 20.6150 ;
      RECT 5.3190 21.3550 5.3370 21.3920 ;
      RECT 5.3190 23.3950 5.3370 23.6930 ;
      RECT 5.2830 18.7690 5.3010 19.2740 ;
      RECT 5.2830 19.5430 5.3010 20.3450 ;
      RECT 5.2830 21.3880 5.3010 21.6590 ;
      RECT 5.2830 21.7390 5.3010 21.9650 ;
      RECT 5.2470 18.6970 5.2650 19.3730 ;
      RECT 5.2470 19.4710 5.2650 19.8050 ;
      RECT 5.2470 20.0110 5.2650 20.1470 ;
      RECT 5.2470 20.6950 5.2650 21.4970 ;
      RECT 5.2470 21.9310 5.2650 21.9680 ;
      RECT 5.2470 24.0970 5.2650 24.4310 ;
      RECT 5.2110 18.9310 5.2290 19.0670 ;
      RECT 5.2110 20.8210 5.2290 21.8030 ;
      RECT 5.2110 22.2430 5.2290 22.5410 ;
      RECT 5.2110 23.9350 5.2290 24.1970 ;
      RECT 5.1750 17.9950 5.1930 18.1490 ;
      RECT 5.1750 18.8050 5.1930 20.5910 ;
      RECT 5.1750 21.6310 5.1930 23.9630 ;
      RECT 5.1750 24.1690 5.1930 25.2770 ;
      RECT 4.8870 18.2650 4.9050 18.5270 ;
      RECT 4.8870 18.6610 4.9050 18.7250 ;
      RECT 4.8870 18.8050 4.9050 19.0310 ;
      RECT 4.8870 19.0750 4.9050 19.2650 ;
      RECT 4.8870 19.3450 4.9050 21.9650 ;
      RECT 4.8870 22.0090 4.9050 23.3150 ;
      RECT 4.8870 24.4030 4.9050 24.6650 ;
      RECT 4.8510 19.2640 4.8690 19.5350 ;
      RECT 4.8510 19.6150 4.8690 20.4530 ;
      RECT 4.8510 20.6230 4.8690 21.4610 ;
      RECT 4.8510 21.5050 4.8690 22.7750 ;
      RECT 4.8510 22.9810 4.8690 23.1530 ;
      RECT 4.8510 23.8630 4.8690 24.9350 ;
      RECT 4.8150 19.3450 4.8330 19.6160 ;
      RECT 4.8150 19.7710 4.8330 19.8080 ;
      RECT 4.8150 20.5510 4.8330 21.5330 ;
      RECT 4.8150 21.7750 4.8330 22.2350 ;
      RECT 4.8150 22.5850 4.8330 23.3240 ;
      RECT 4.7790 18.4630 4.7970 19.5350 ;
      RECT 4.7790 21.1270 4.7970 21.3440 ;
      RECT 4.7790 22.5130 4.7970 22.8110 ;
      RECT 4.7430 19.1110 4.7610 19.5710 ;
      RECT 4.7430 20.6950 4.7610 20.8850 ;
      RECT 4.7430 20.9260 4.7610 20.9630 ;
      RECT 4.7430 21.1990 4.7610 21.5330 ;
      RECT 4.7430 21.6670 4.7610 23.0090 ;
      RECT 4.7430 23.1160 4.7610 24.2330 ;
      RECT 4.7070 18.5350 4.7250 18.7250 ;
      RECT 4.7070 18.9310 4.7250 19.0670 ;
      RECT 4.7070 19.3450 4.7250 22.5050 ;
      RECT 4.7070 22.5850 4.7250 23.0450 ;
      RECT 4.7070 23.6650 4.7250 24.1250 ;
      RECT 4.7070 24.9790 4.7250 25.2050 ;
      RECT 4.6710 17.5230 4.6890 17.6770 ;
      RECT 4.6710 25.5340 4.6890 25.6880 ;
      RECT 4.6350 17.5230 4.6530 17.5730 ;
      RECT 4.5630 17.5230 4.5810 17.5945 ;
      RECT 4.5630 25.6035 4.5810 25.7035 ;
      RECT 4.4190 19.0390 4.4370 19.2290 ;
      RECT 4.4190 19.7770 4.4370 20.1470 ;
      RECT 4.4190 21.7390 4.4370 21.9650 ;
      RECT 4.4190 22.2790 4.4370 23.4230 ;
      RECT 4.4190 24.2050 4.4370 24.6650 ;
      RECT 4.4190 25.2430 4.4370 25.2800 ;
      RECT 4.3830 17.9950 4.4010 18.4910 ;
      RECT 4.3830 22.0750 4.4010 22.1120 ;
      RECT 4.3830 23.1520 4.4010 23.9630 ;
      RECT 4.3470 18.4630 4.3650 18.7250 ;
      RECT 4.3470 19.0030 4.3650 19.3370 ;
      RECT 4.3470 19.5430 4.3650 19.6430 ;
      RECT 4.3470 20.4250 4.3650 23.1890 ;
      RECT 4.3470 23.3230 4.3650 23.5490 ;
      RECT 4.3110 18.1210 4.3290 19.2650 ;
      RECT 4.3110 22.8550 4.3290 23.0450 ;
      RECT 4.3110 23.6590 4.3290 23.6960 ;
      RECT 4.3110 23.9350 4.3290 24.7370 ;
      RECT 4.2750 19.0750 4.2930 20.0750 ;
      RECT 4.2750 23.5150 4.2930 23.5520 ;
      RECT 4.2390 18.2650 4.2570 18.2930 ;
      RECT 3.9150 18.6610 3.9330 19.0670 ;
      RECT 3.8430 18.6970 3.8610 19.3010 ;
      RECT 3.8070 18.5350 3.8250 18.5990 ;
      RECT 3.7710 17.5760 3.7890 17.6270 ;
      RECT 3.7710 20.6950 3.7890 20.8850 ;
      RECT 3.7710 21.3160 3.7890 25.6760 ;
      RECT 3.6810 21.3160 3.6990 25.6760 ;
      RECT 3.6630 17.9950 3.6810 18.1850 ;
      RECT 3.6630 18.7690 3.6810 21.0290 ;
      RECT 3.6450 21.6210 3.6630 21.7040 ;
      RECT 3.6090 17.4965 3.6270 25.7035 ;
      RECT 3.5730 21.3485 3.5910 22.0385 ;
      RECT 3.5730 22.0895 3.5910 23.0810 ;
      RECT 3.5730 23.1110 3.5910 23.8950 ;
      RECT 3.5550 17.9950 3.5730 18.4910 ;
      RECT 3.5550 19.2730 3.5730 19.8410 ;
      RECT 3.5550 20.1550 3.5730 20.8850 ;
      RECT 3.5370 21.2850 3.5550 21.9897 ;
      RECT 3.5370 22.7320 3.5550 23.9130 ;
      RECT 3.5010 17.4965 3.5190 17.8465 ;
      RECT 3.3930 17.4965 3.4110 17.8465 ;
      RECT 3.2850 17.4965 3.3030 17.8465 ;
      RECT 3.1770 17.4965 3.1950 17.8465 ;
      RECT 3.0690 17.4965 3.0870 17.8465 ;
      RECT 2.9610 17.4965 2.9790 17.8465 ;
      RECT 2.8530 17.4965 2.8710 17.8465 ;
      RECT 2.7450 17.4965 2.7630 17.8465 ;
      RECT 2.6370 17.4965 2.6550 17.8465 ;
      RECT 2.5290 17.4965 2.5470 17.8465 ;
      RECT 2.4210 17.4965 2.4390 17.8465 ;
      RECT 2.3130 17.4965 2.3310 17.8465 ;
      RECT 2.2050 17.4965 2.2230 17.8465 ;
      RECT 2.0970 17.4965 2.1150 17.8465 ;
      RECT 1.9890 17.4965 2.0070 17.8465 ;
      RECT 1.8810 17.4965 1.8990 17.8465 ;
      RECT 1.7730 17.4965 1.7910 17.8465 ;
      RECT 1.6650 17.4965 1.6830 17.8465 ;
      RECT 1.5570 17.4965 1.5750 17.8465 ;
      RECT 1.4490 17.4965 1.4670 17.8465 ;
      RECT 1.3410 17.4965 1.3590 17.8465 ;
      RECT 1.2330 17.4965 1.2510 17.8465 ;
      RECT 1.1250 17.4965 1.1430 17.8465 ;
      RECT 1.0170 17.4965 1.0350 17.8465 ;
      RECT 0.9090 17.4965 0.9270 17.8465 ;
      RECT 0.8010 17.4965 0.8190 17.8465 ;
      RECT 0.6930 17.4965 0.7110 17.8465 ;
      RECT 0.5850 17.4965 0.6030 17.8465 ;
      RECT 0.4770 17.4965 0.4950 17.8465 ;
      RECT 0.3690 17.4965 0.3870 17.8465 ;
      RECT 0.3330 21.3515 0.3510 21.9935 ;
      RECT 0.3330 22.6710 0.3510 23.2030 ;
      RECT 0.3150 18.5350 0.3330 18.7610 ;
      RECT 0.2970 21.2660 0.3150 22.0385 ;
      RECT 0.2970 22.0897 0.3150 22.5810 ;
      RECT 0.2970 22.6310 0.3150 23.0025 ;
      RECT 0.2970 23.0655 0.3150 23.8770 ;
      RECT 0.2610 17.4965 0.2790 25.7035 ;
      RECT 0.2250 20.0010 0.2430 20.0700 ;
      RECT 0.2250 21.8090 0.2430 22.2735 ;
      RECT 0.1890 21.3160 0.2070 25.6715 ;
        RECT 5.2380 25.7520 5.2560 26.6875 ;
        RECT 5.2020 25.7520 5.2200 26.6875 ;
        RECT 5.1660 26.3290 5.1840 26.6515 ;
        RECT 5.0490 26.5260 5.0670 26.6355 ;
        RECT 5.0400 25.7845 5.0580 26.0240 ;
        RECT 5.0040 26.3655 5.0220 26.5190 ;
        RECT 4.9230 26.3910 4.9410 26.6490 ;
        RECT 4.3830 25.7520 4.4010 26.6875 ;
        RECT 4.3470 25.7520 4.3650 26.6875 ;
        RECT 4.3110 25.9330 4.3290 26.5010 ;
        RECT 5.2380 26.8320 5.2560 27.7675 ;
        RECT 5.2020 26.8320 5.2200 27.7675 ;
        RECT 5.1660 27.4090 5.1840 27.7315 ;
        RECT 5.0490 27.6060 5.0670 27.7155 ;
        RECT 5.0400 26.8645 5.0580 27.1040 ;
        RECT 5.0040 27.4455 5.0220 27.5990 ;
        RECT 4.9230 27.4710 4.9410 27.7290 ;
        RECT 4.3830 26.8320 4.4010 27.7675 ;
        RECT 4.3470 26.8320 4.3650 27.7675 ;
        RECT 4.3110 27.0130 4.3290 27.5810 ;
        RECT 5.2380 27.9120 5.2560 28.8475 ;
        RECT 5.2020 27.9120 5.2200 28.8475 ;
        RECT 5.1660 28.4890 5.1840 28.8115 ;
        RECT 5.0490 28.6860 5.0670 28.7955 ;
        RECT 5.0400 27.9445 5.0580 28.1840 ;
        RECT 5.0040 28.5255 5.0220 28.6790 ;
        RECT 4.9230 28.5510 4.9410 28.8090 ;
        RECT 4.3830 27.9120 4.4010 28.8475 ;
        RECT 4.3470 27.9120 4.3650 28.8475 ;
        RECT 4.3110 28.0930 4.3290 28.6610 ;
        RECT 5.2380 28.9920 5.2560 29.9275 ;
        RECT 5.2020 28.9920 5.2200 29.9275 ;
        RECT 5.1660 29.5690 5.1840 29.8915 ;
        RECT 5.0490 29.7660 5.0670 29.8755 ;
        RECT 5.0400 29.0245 5.0580 29.2640 ;
        RECT 5.0040 29.6055 5.0220 29.7590 ;
        RECT 4.9230 29.6310 4.9410 29.8890 ;
        RECT 4.3830 28.9920 4.4010 29.9275 ;
        RECT 4.3470 28.9920 4.3650 29.9275 ;
        RECT 4.3110 29.1730 4.3290 29.7410 ;
        RECT 5.2380 30.0720 5.2560 31.0075 ;
        RECT 5.2020 30.0720 5.2200 31.0075 ;
        RECT 5.1660 30.6490 5.1840 30.9715 ;
        RECT 5.0490 30.8460 5.0670 30.9555 ;
        RECT 5.0400 30.1045 5.0580 30.3440 ;
        RECT 5.0040 30.6855 5.0220 30.8390 ;
        RECT 4.9230 30.7110 4.9410 30.9690 ;
        RECT 4.3830 30.0720 4.4010 31.0075 ;
        RECT 4.3470 30.0720 4.3650 31.0075 ;
        RECT 4.3110 30.2530 4.3290 30.8210 ;
        RECT 5.2380 31.1520 5.2560 32.0875 ;
        RECT 5.2020 31.1520 5.2200 32.0875 ;
        RECT 5.1660 31.7290 5.1840 32.0515 ;
        RECT 5.0490 31.9260 5.0670 32.0355 ;
        RECT 5.0400 31.1845 5.0580 31.4240 ;
        RECT 5.0040 31.7655 5.0220 31.9190 ;
        RECT 4.9230 31.7910 4.9410 32.0490 ;
        RECT 4.3830 31.1520 4.4010 32.0875 ;
        RECT 4.3470 31.1520 4.3650 32.0875 ;
        RECT 4.3110 31.3330 4.3290 31.9010 ;
        RECT 5.2380 32.2320 5.2560 33.1675 ;
        RECT 5.2020 32.2320 5.2200 33.1675 ;
        RECT 5.1660 32.8090 5.1840 33.1315 ;
        RECT 5.0490 33.0060 5.0670 33.1155 ;
        RECT 5.0400 32.2645 5.0580 32.5040 ;
        RECT 5.0040 32.8455 5.0220 32.9990 ;
        RECT 4.9230 32.8710 4.9410 33.1290 ;
        RECT 4.3830 32.2320 4.4010 33.1675 ;
        RECT 4.3470 32.2320 4.3650 33.1675 ;
        RECT 4.3110 32.4130 4.3290 32.9810 ;
        RECT 5.2380 33.3120 5.2560 34.2475 ;
        RECT 5.2020 33.3120 5.2200 34.2475 ;
        RECT 5.1660 33.8890 5.1840 34.2115 ;
        RECT 5.0490 34.0860 5.0670 34.1955 ;
        RECT 5.0400 33.3445 5.0580 33.5840 ;
        RECT 5.0040 33.9255 5.0220 34.0790 ;
        RECT 4.9230 33.9510 4.9410 34.2090 ;
        RECT 4.3830 33.3120 4.4010 34.2475 ;
        RECT 4.3470 33.3120 4.3650 34.2475 ;
        RECT 4.3110 33.4930 4.3290 34.0610 ;
        RECT 5.2380 34.3920 5.2560 35.3275 ;
        RECT 5.2020 34.3920 5.2200 35.3275 ;
        RECT 5.1660 34.9690 5.1840 35.2915 ;
        RECT 5.0490 35.1660 5.0670 35.2755 ;
        RECT 5.0400 34.4245 5.0580 34.6640 ;
        RECT 5.0040 35.0055 5.0220 35.1590 ;
        RECT 4.9230 35.0310 4.9410 35.2890 ;
        RECT 4.3830 34.3920 4.4010 35.3275 ;
        RECT 4.3470 34.3920 4.3650 35.3275 ;
        RECT 4.3110 34.5730 4.3290 35.1410 ;
        RECT 5.2380 35.4720 5.2560 36.4075 ;
        RECT 5.2020 35.4720 5.2200 36.4075 ;
        RECT 5.1660 36.0490 5.1840 36.3715 ;
        RECT 5.0490 36.2460 5.0670 36.3555 ;
        RECT 5.0400 35.5045 5.0580 35.7440 ;
        RECT 5.0040 36.0855 5.0220 36.2390 ;
        RECT 4.9230 36.1110 4.9410 36.3690 ;
        RECT 4.3830 35.4720 4.4010 36.4075 ;
        RECT 4.3470 35.4720 4.3650 36.4075 ;
        RECT 4.3110 35.6530 4.3290 36.2210 ;
        RECT 5.2380 36.5520 5.2560 37.4875 ;
        RECT 5.2020 36.5520 5.2200 37.4875 ;
        RECT 5.1660 37.1290 5.1840 37.4515 ;
        RECT 5.0490 37.3260 5.0670 37.4355 ;
        RECT 5.0400 36.5845 5.0580 36.8240 ;
        RECT 5.0040 37.1655 5.0220 37.3190 ;
        RECT 4.9230 37.1910 4.9410 37.4490 ;
        RECT 4.3830 36.5520 4.4010 37.4875 ;
        RECT 4.3470 36.5520 4.3650 37.4875 ;
        RECT 4.3110 36.7330 4.3290 37.3010 ;
        RECT 5.2380 37.6320 5.2560 38.5675 ;
        RECT 5.2020 37.6320 5.2200 38.5675 ;
        RECT 5.1660 38.2090 5.1840 38.5315 ;
        RECT 5.0490 38.4060 5.0670 38.5155 ;
        RECT 5.0400 37.6645 5.0580 37.9040 ;
        RECT 5.0040 38.2455 5.0220 38.3990 ;
        RECT 4.9230 38.2710 4.9410 38.5290 ;
        RECT 4.3830 37.6320 4.4010 38.5675 ;
        RECT 4.3470 37.6320 4.3650 38.5675 ;
        RECT 4.3110 37.8130 4.3290 38.3810 ;
        RECT 5.2380 38.7120 5.2560 39.6475 ;
        RECT 5.2020 38.7120 5.2200 39.6475 ;
        RECT 5.1660 39.2890 5.1840 39.6115 ;
        RECT 5.0490 39.4860 5.0670 39.5955 ;
        RECT 5.0400 38.7445 5.0580 38.9840 ;
        RECT 5.0040 39.3255 5.0220 39.4790 ;
        RECT 4.9230 39.3510 4.9410 39.6090 ;
        RECT 4.3830 38.7120 4.4010 39.6475 ;
        RECT 4.3470 38.7120 4.3650 39.6475 ;
        RECT 4.3110 38.8930 4.3290 39.4610 ;
        RECT 5.2380 39.7920 5.2560 40.7275 ;
        RECT 5.2020 39.7920 5.2200 40.7275 ;
        RECT 5.1660 40.3690 5.1840 40.6915 ;
        RECT 5.0490 40.5660 5.0670 40.6755 ;
        RECT 5.0400 39.8245 5.0580 40.0640 ;
        RECT 5.0040 40.4055 5.0220 40.5590 ;
        RECT 4.9230 40.4310 4.9410 40.6890 ;
        RECT 4.3830 39.7920 4.4010 40.7275 ;
        RECT 4.3470 39.7920 4.3650 40.7275 ;
        RECT 4.3110 39.9730 4.3290 40.5410 ;
        RECT 5.2380 40.8720 5.2560 41.8075 ;
        RECT 5.2020 40.8720 5.2200 41.8075 ;
        RECT 5.1660 41.4490 5.1840 41.7715 ;
        RECT 5.0490 41.6460 5.0670 41.7555 ;
        RECT 5.0400 40.9045 5.0580 41.1440 ;
        RECT 5.0040 41.4855 5.0220 41.6390 ;
        RECT 4.9230 41.5110 4.9410 41.7690 ;
        RECT 4.3830 40.8720 4.4010 41.8075 ;
        RECT 4.3470 40.8720 4.3650 41.8075 ;
        RECT 4.3110 41.0530 4.3290 41.6210 ;
        RECT 5.2380 41.9520 5.2560 42.8875 ;
        RECT 5.2020 41.9520 5.2200 42.8875 ;
        RECT 5.1660 42.5290 5.1840 42.8515 ;
        RECT 5.0490 42.7260 5.0670 42.8355 ;
        RECT 5.0400 41.9845 5.0580 42.2240 ;
        RECT 5.0040 42.5655 5.0220 42.7190 ;
        RECT 4.9230 42.5910 4.9410 42.8490 ;
        RECT 4.3830 41.9520 4.4010 42.8875 ;
        RECT 4.3470 41.9520 4.3650 42.8875 ;
        RECT 4.3110 42.1330 4.3290 42.7010 ;
  LAYER M3 SPACING 0.018  ;
      RECT 5.1800 0.2565 5.3080 1.3500 ;
      RECT 5.1660 0.9220 5.3080 1.2445 ;
      RECT 5.0180 0.6490 5.0800 1.3500 ;
      RECT 5.0040 0.9585 5.0800 1.1120 ;
      RECT 5.0180 0.2565 5.0440 1.3500 ;
      RECT 5.0180 0.3775 5.0580 0.6170 ;
      RECT 5.0180 0.2565 5.0800 0.3455 ;
      RECT 4.7210 0.7070 4.9270 1.3500 ;
      RECT 4.9010 0.2565 4.9270 1.3500 ;
      RECT 4.7210 0.9840 4.9410 1.2420 ;
      RECT 4.7210 0.2565 4.8190 1.3500 ;
      RECT 4.3040 0.2565 4.3870 1.3500 ;
      RECT 4.3040 0.3450 4.4010 1.2805 ;
      RECT 9.5270 0.2565 9.6120 1.3500 ;
      RECT 9.3830 0.2565 9.4090 1.3500 ;
      RECT 9.2750 0.2565 9.3010 1.3500 ;
      RECT 9.1670 0.2565 9.1930 1.3500 ;
      RECT 9.0590 0.2565 9.0850 1.3500 ;
      RECT 8.9510 0.2565 8.9770 1.3500 ;
      RECT 8.8430 0.2565 8.8690 1.3500 ;
      RECT 8.7350 0.2565 8.7610 1.3500 ;
      RECT 8.6270 0.2565 8.6530 1.3500 ;
      RECT 8.5190 0.2565 8.5450 1.3500 ;
      RECT 8.4110 0.2565 8.4370 1.3500 ;
      RECT 8.3030 0.2565 8.3290 1.3500 ;
      RECT 8.1950 0.2565 8.2210 1.3500 ;
      RECT 8.0870 0.2565 8.1130 1.3500 ;
      RECT 7.9790 0.2565 8.0050 1.3500 ;
      RECT 7.8710 0.2565 7.8970 1.3500 ;
      RECT 7.7630 0.2565 7.7890 1.3500 ;
      RECT 7.6550 0.2565 7.6810 1.3500 ;
      RECT 7.5470 0.2565 7.5730 1.3500 ;
      RECT 7.4390 0.2565 7.4650 1.3500 ;
      RECT 7.3310 0.2565 7.3570 1.3500 ;
      RECT 7.2230 0.2565 7.2490 1.3500 ;
      RECT 7.1150 0.2565 7.1410 1.3500 ;
      RECT 7.0070 0.2565 7.0330 1.3500 ;
      RECT 6.8990 0.2565 6.9250 1.3500 ;
      RECT 6.7910 0.2565 6.8170 1.3500 ;
      RECT 6.6830 0.2565 6.7090 1.3500 ;
      RECT 6.5750 0.2565 6.6010 1.3500 ;
      RECT 6.4670 0.2565 6.4930 1.3500 ;
      RECT 6.3590 0.2565 6.3850 1.3500 ;
      RECT 6.2510 0.2565 6.2770 1.3500 ;
      RECT 6.1430 0.2565 6.1690 1.3500 ;
      RECT 6.0350 0.2565 6.0610 1.3500 ;
      RECT 5.9270 0.2565 5.9530 1.3500 ;
      RECT 5.7140 0.2565 5.7910 1.3500 ;
      RECT 3.8210 0.2565 3.8980 1.3500 ;
      RECT 3.6590 0.2565 3.6850 1.3500 ;
      RECT 3.5510 0.2565 3.5770 1.3500 ;
      RECT 3.4430 0.2565 3.4690 1.3500 ;
      RECT 3.3350 0.2565 3.3610 1.3500 ;
      RECT 3.2270 0.2565 3.2530 1.3500 ;
      RECT 3.1190 0.2565 3.1450 1.3500 ;
      RECT 3.0110 0.2565 3.0370 1.3500 ;
      RECT 2.9030 0.2565 2.9290 1.3500 ;
      RECT 2.7950 0.2565 2.8210 1.3500 ;
      RECT 2.6870 0.2565 2.7130 1.3500 ;
      RECT 2.5790 0.2565 2.6050 1.3500 ;
      RECT 2.4710 0.2565 2.4970 1.3500 ;
      RECT 2.3630 0.2565 2.3890 1.3500 ;
      RECT 2.2550 0.2565 2.2810 1.3500 ;
      RECT 2.1470 0.2565 2.1730 1.3500 ;
      RECT 2.0390 0.2565 2.0650 1.3500 ;
      RECT 1.9310 0.2565 1.9570 1.3500 ;
      RECT 1.8230 0.2565 1.8490 1.3500 ;
      RECT 1.7150 0.2565 1.7410 1.3500 ;
      RECT 1.6070 0.2565 1.6330 1.3500 ;
      RECT 1.4990 0.2565 1.5250 1.3500 ;
      RECT 1.3910 0.2565 1.4170 1.3500 ;
      RECT 1.2830 0.2565 1.3090 1.3500 ;
      RECT 1.1750 0.2565 1.2010 1.3500 ;
      RECT 1.0670 0.2565 1.0930 1.3500 ;
      RECT 0.9590 0.2565 0.9850 1.3500 ;
      RECT 0.8510 0.2565 0.8770 1.3500 ;
      RECT 0.7430 0.2565 0.7690 1.3500 ;
      RECT 0.6350 0.2565 0.6610 1.3500 ;
      RECT 0.5270 0.2565 0.5530 1.3500 ;
      RECT 0.4190 0.2565 0.4450 1.3500 ;
      RECT 0.3110 0.2565 0.3370 1.3500 ;
      RECT 0.2030 0.2565 0.2290 1.3500 ;
      RECT 0.0000 0.2565 0.0850 1.3500 ;
      RECT 5.1800 1.3365 5.3080 2.4300 ;
      RECT 5.1660 2.0020 5.3080 2.3245 ;
      RECT 5.0180 1.7290 5.0800 2.4300 ;
      RECT 5.0040 2.0385 5.0800 2.1920 ;
      RECT 5.0180 1.3365 5.0440 2.4300 ;
      RECT 5.0180 1.4575 5.0580 1.6970 ;
      RECT 5.0180 1.3365 5.0800 1.4255 ;
      RECT 4.7210 1.7870 4.9270 2.4300 ;
      RECT 4.9010 1.3365 4.9270 2.4300 ;
      RECT 4.7210 2.0640 4.9410 2.3220 ;
      RECT 4.7210 1.3365 4.8190 2.4300 ;
      RECT 4.3040 1.3365 4.3870 2.4300 ;
      RECT 4.3040 1.4250 4.4010 2.3605 ;
      RECT 9.5270 1.3365 9.6120 2.4300 ;
      RECT 9.3830 1.3365 9.4090 2.4300 ;
      RECT 9.2750 1.3365 9.3010 2.4300 ;
      RECT 9.1670 1.3365 9.1930 2.4300 ;
      RECT 9.0590 1.3365 9.0850 2.4300 ;
      RECT 8.9510 1.3365 8.9770 2.4300 ;
      RECT 8.8430 1.3365 8.8690 2.4300 ;
      RECT 8.7350 1.3365 8.7610 2.4300 ;
      RECT 8.6270 1.3365 8.6530 2.4300 ;
      RECT 8.5190 1.3365 8.5450 2.4300 ;
      RECT 8.4110 1.3365 8.4370 2.4300 ;
      RECT 8.3030 1.3365 8.3290 2.4300 ;
      RECT 8.1950 1.3365 8.2210 2.4300 ;
      RECT 8.0870 1.3365 8.1130 2.4300 ;
      RECT 7.9790 1.3365 8.0050 2.4300 ;
      RECT 7.8710 1.3365 7.8970 2.4300 ;
      RECT 7.7630 1.3365 7.7890 2.4300 ;
      RECT 7.6550 1.3365 7.6810 2.4300 ;
      RECT 7.5470 1.3365 7.5730 2.4300 ;
      RECT 7.4390 1.3365 7.4650 2.4300 ;
      RECT 7.3310 1.3365 7.3570 2.4300 ;
      RECT 7.2230 1.3365 7.2490 2.4300 ;
      RECT 7.1150 1.3365 7.1410 2.4300 ;
      RECT 7.0070 1.3365 7.0330 2.4300 ;
      RECT 6.8990 1.3365 6.9250 2.4300 ;
      RECT 6.7910 1.3365 6.8170 2.4300 ;
      RECT 6.6830 1.3365 6.7090 2.4300 ;
      RECT 6.5750 1.3365 6.6010 2.4300 ;
      RECT 6.4670 1.3365 6.4930 2.4300 ;
      RECT 6.3590 1.3365 6.3850 2.4300 ;
      RECT 6.2510 1.3365 6.2770 2.4300 ;
      RECT 6.1430 1.3365 6.1690 2.4300 ;
      RECT 6.0350 1.3365 6.0610 2.4300 ;
      RECT 5.9270 1.3365 5.9530 2.4300 ;
      RECT 5.7140 1.3365 5.7910 2.4300 ;
      RECT 3.8210 1.3365 3.8980 2.4300 ;
      RECT 3.6590 1.3365 3.6850 2.4300 ;
      RECT 3.5510 1.3365 3.5770 2.4300 ;
      RECT 3.4430 1.3365 3.4690 2.4300 ;
      RECT 3.3350 1.3365 3.3610 2.4300 ;
      RECT 3.2270 1.3365 3.2530 2.4300 ;
      RECT 3.1190 1.3365 3.1450 2.4300 ;
      RECT 3.0110 1.3365 3.0370 2.4300 ;
      RECT 2.9030 1.3365 2.9290 2.4300 ;
      RECT 2.7950 1.3365 2.8210 2.4300 ;
      RECT 2.6870 1.3365 2.7130 2.4300 ;
      RECT 2.5790 1.3365 2.6050 2.4300 ;
      RECT 2.4710 1.3365 2.4970 2.4300 ;
      RECT 2.3630 1.3365 2.3890 2.4300 ;
      RECT 2.2550 1.3365 2.2810 2.4300 ;
      RECT 2.1470 1.3365 2.1730 2.4300 ;
      RECT 2.0390 1.3365 2.0650 2.4300 ;
      RECT 1.9310 1.3365 1.9570 2.4300 ;
      RECT 1.8230 1.3365 1.8490 2.4300 ;
      RECT 1.7150 1.3365 1.7410 2.4300 ;
      RECT 1.6070 1.3365 1.6330 2.4300 ;
      RECT 1.4990 1.3365 1.5250 2.4300 ;
      RECT 1.3910 1.3365 1.4170 2.4300 ;
      RECT 1.2830 1.3365 1.3090 2.4300 ;
      RECT 1.1750 1.3365 1.2010 2.4300 ;
      RECT 1.0670 1.3365 1.0930 2.4300 ;
      RECT 0.9590 1.3365 0.9850 2.4300 ;
      RECT 0.8510 1.3365 0.8770 2.4300 ;
      RECT 0.7430 1.3365 0.7690 2.4300 ;
      RECT 0.6350 1.3365 0.6610 2.4300 ;
      RECT 0.5270 1.3365 0.5530 2.4300 ;
      RECT 0.4190 1.3365 0.4450 2.4300 ;
      RECT 0.3110 1.3365 0.3370 2.4300 ;
      RECT 0.2030 1.3365 0.2290 2.4300 ;
      RECT 0.0000 1.3365 0.0850 2.4300 ;
      RECT 5.1800 2.4165 5.3080 3.5100 ;
      RECT 5.1660 3.0820 5.3080 3.4045 ;
      RECT 5.0180 2.8090 5.0800 3.5100 ;
      RECT 5.0040 3.1185 5.0800 3.2720 ;
      RECT 5.0180 2.4165 5.0440 3.5100 ;
      RECT 5.0180 2.5375 5.0580 2.7770 ;
      RECT 5.0180 2.4165 5.0800 2.5055 ;
      RECT 4.7210 2.8670 4.9270 3.5100 ;
      RECT 4.9010 2.4165 4.9270 3.5100 ;
      RECT 4.7210 3.1440 4.9410 3.4020 ;
      RECT 4.7210 2.4165 4.8190 3.5100 ;
      RECT 4.3040 2.4165 4.3870 3.5100 ;
      RECT 4.3040 2.5050 4.4010 3.4405 ;
      RECT 9.5270 2.4165 9.6120 3.5100 ;
      RECT 9.3830 2.4165 9.4090 3.5100 ;
      RECT 9.2750 2.4165 9.3010 3.5100 ;
      RECT 9.1670 2.4165 9.1930 3.5100 ;
      RECT 9.0590 2.4165 9.0850 3.5100 ;
      RECT 8.9510 2.4165 8.9770 3.5100 ;
      RECT 8.8430 2.4165 8.8690 3.5100 ;
      RECT 8.7350 2.4165 8.7610 3.5100 ;
      RECT 8.6270 2.4165 8.6530 3.5100 ;
      RECT 8.5190 2.4165 8.5450 3.5100 ;
      RECT 8.4110 2.4165 8.4370 3.5100 ;
      RECT 8.3030 2.4165 8.3290 3.5100 ;
      RECT 8.1950 2.4165 8.2210 3.5100 ;
      RECT 8.0870 2.4165 8.1130 3.5100 ;
      RECT 7.9790 2.4165 8.0050 3.5100 ;
      RECT 7.8710 2.4165 7.8970 3.5100 ;
      RECT 7.7630 2.4165 7.7890 3.5100 ;
      RECT 7.6550 2.4165 7.6810 3.5100 ;
      RECT 7.5470 2.4165 7.5730 3.5100 ;
      RECT 7.4390 2.4165 7.4650 3.5100 ;
      RECT 7.3310 2.4165 7.3570 3.5100 ;
      RECT 7.2230 2.4165 7.2490 3.5100 ;
      RECT 7.1150 2.4165 7.1410 3.5100 ;
      RECT 7.0070 2.4165 7.0330 3.5100 ;
      RECT 6.8990 2.4165 6.9250 3.5100 ;
      RECT 6.7910 2.4165 6.8170 3.5100 ;
      RECT 6.6830 2.4165 6.7090 3.5100 ;
      RECT 6.5750 2.4165 6.6010 3.5100 ;
      RECT 6.4670 2.4165 6.4930 3.5100 ;
      RECT 6.3590 2.4165 6.3850 3.5100 ;
      RECT 6.2510 2.4165 6.2770 3.5100 ;
      RECT 6.1430 2.4165 6.1690 3.5100 ;
      RECT 6.0350 2.4165 6.0610 3.5100 ;
      RECT 5.9270 2.4165 5.9530 3.5100 ;
      RECT 5.7140 2.4165 5.7910 3.5100 ;
      RECT 3.8210 2.4165 3.8980 3.5100 ;
      RECT 3.6590 2.4165 3.6850 3.5100 ;
      RECT 3.5510 2.4165 3.5770 3.5100 ;
      RECT 3.4430 2.4165 3.4690 3.5100 ;
      RECT 3.3350 2.4165 3.3610 3.5100 ;
      RECT 3.2270 2.4165 3.2530 3.5100 ;
      RECT 3.1190 2.4165 3.1450 3.5100 ;
      RECT 3.0110 2.4165 3.0370 3.5100 ;
      RECT 2.9030 2.4165 2.9290 3.5100 ;
      RECT 2.7950 2.4165 2.8210 3.5100 ;
      RECT 2.6870 2.4165 2.7130 3.5100 ;
      RECT 2.5790 2.4165 2.6050 3.5100 ;
      RECT 2.4710 2.4165 2.4970 3.5100 ;
      RECT 2.3630 2.4165 2.3890 3.5100 ;
      RECT 2.2550 2.4165 2.2810 3.5100 ;
      RECT 2.1470 2.4165 2.1730 3.5100 ;
      RECT 2.0390 2.4165 2.0650 3.5100 ;
      RECT 1.9310 2.4165 1.9570 3.5100 ;
      RECT 1.8230 2.4165 1.8490 3.5100 ;
      RECT 1.7150 2.4165 1.7410 3.5100 ;
      RECT 1.6070 2.4165 1.6330 3.5100 ;
      RECT 1.4990 2.4165 1.5250 3.5100 ;
      RECT 1.3910 2.4165 1.4170 3.5100 ;
      RECT 1.2830 2.4165 1.3090 3.5100 ;
      RECT 1.1750 2.4165 1.2010 3.5100 ;
      RECT 1.0670 2.4165 1.0930 3.5100 ;
      RECT 0.9590 2.4165 0.9850 3.5100 ;
      RECT 0.8510 2.4165 0.8770 3.5100 ;
      RECT 0.7430 2.4165 0.7690 3.5100 ;
      RECT 0.6350 2.4165 0.6610 3.5100 ;
      RECT 0.5270 2.4165 0.5530 3.5100 ;
      RECT 0.4190 2.4165 0.4450 3.5100 ;
      RECT 0.3110 2.4165 0.3370 3.5100 ;
      RECT 0.2030 2.4165 0.2290 3.5100 ;
      RECT 0.0000 2.4165 0.0850 3.5100 ;
      RECT 5.1800 3.4965 5.3080 4.5900 ;
      RECT 5.1660 4.1620 5.3080 4.4845 ;
      RECT 5.0180 3.8890 5.0800 4.5900 ;
      RECT 5.0040 4.1985 5.0800 4.3520 ;
      RECT 5.0180 3.4965 5.0440 4.5900 ;
      RECT 5.0180 3.6175 5.0580 3.8570 ;
      RECT 5.0180 3.4965 5.0800 3.5855 ;
      RECT 4.7210 3.9470 4.9270 4.5900 ;
      RECT 4.9010 3.4965 4.9270 4.5900 ;
      RECT 4.7210 4.2240 4.9410 4.4820 ;
      RECT 4.7210 3.4965 4.8190 4.5900 ;
      RECT 4.3040 3.4965 4.3870 4.5900 ;
      RECT 4.3040 3.5850 4.4010 4.5205 ;
      RECT 9.5270 3.4965 9.6120 4.5900 ;
      RECT 9.3830 3.4965 9.4090 4.5900 ;
      RECT 9.2750 3.4965 9.3010 4.5900 ;
      RECT 9.1670 3.4965 9.1930 4.5900 ;
      RECT 9.0590 3.4965 9.0850 4.5900 ;
      RECT 8.9510 3.4965 8.9770 4.5900 ;
      RECT 8.8430 3.4965 8.8690 4.5900 ;
      RECT 8.7350 3.4965 8.7610 4.5900 ;
      RECT 8.6270 3.4965 8.6530 4.5900 ;
      RECT 8.5190 3.4965 8.5450 4.5900 ;
      RECT 8.4110 3.4965 8.4370 4.5900 ;
      RECT 8.3030 3.4965 8.3290 4.5900 ;
      RECT 8.1950 3.4965 8.2210 4.5900 ;
      RECT 8.0870 3.4965 8.1130 4.5900 ;
      RECT 7.9790 3.4965 8.0050 4.5900 ;
      RECT 7.8710 3.4965 7.8970 4.5900 ;
      RECT 7.7630 3.4965 7.7890 4.5900 ;
      RECT 7.6550 3.4965 7.6810 4.5900 ;
      RECT 7.5470 3.4965 7.5730 4.5900 ;
      RECT 7.4390 3.4965 7.4650 4.5900 ;
      RECT 7.3310 3.4965 7.3570 4.5900 ;
      RECT 7.2230 3.4965 7.2490 4.5900 ;
      RECT 7.1150 3.4965 7.1410 4.5900 ;
      RECT 7.0070 3.4965 7.0330 4.5900 ;
      RECT 6.8990 3.4965 6.9250 4.5900 ;
      RECT 6.7910 3.4965 6.8170 4.5900 ;
      RECT 6.6830 3.4965 6.7090 4.5900 ;
      RECT 6.5750 3.4965 6.6010 4.5900 ;
      RECT 6.4670 3.4965 6.4930 4.5900 ;
      RECT 6.3590 3.4965 6.3850 4.5900 ;
      RECT 6.2510 3.4965 6.2770 4.5900 ;
      RECT 6.1430 3.4965 6.1690 4.5900 ;
      RECT 6.0350 3.4965 6.0610 4.5900 ;
      RECT 5.9270 3.4965 5.9530 4.5900 ;
      RECT 5.7140 3.4965 5.7910 4.5900 ;
      RECT 3.8210 3.4965 3.8980 4.5900 ;
      RECT 3.6590 3.4965 3.6850 4.5900 ;
      RECT 3.5510 3.4965 3.5770 4.5900 ;
      RECT 3.4430 3.4965 3.4690 4.5900 ;
      RECT 3.3350 3.4965 3.3610 4.5900 ;
      RECT 3.2270 3.4965 3.2530 4.5900 ;
      RECT 3.1190 3.4965 3.1450 4.5900 ;
      RECT 3.0110 3.4965 3.0370 4.5900 ;
      RECT 2.9030 3.4965 2.9290 4.5900 ;
      RECT 2.7950 3.4965 2.8210 4.5900 ;
      RECT 2.6870 3.4965 2.7130 4.5900 ;
      RECT 2.5790 3.4965 2.6050 4.5900 ;
      RECT 2.4710 3.4965 2.4970 4.5900 ;
      RECT 2.3630 3.4965 2.3890 4.5900 ;
      RECT 2.2550 3.4965 2.2810 4.5900 ;
      RECT 2.1470 3.4965 2.1730 4.5900 ;
      RECT 2.0390 3.4965 2.0650 4.5900 ;
      RECT 1.9310 3.4965 1.9570 4.5900 ;
      RECT 1.8230 3.4965 1.8490 4.5900 ;
      RECT 1.7150 3.4965 1.7410 4.5900 ;
      RECT 1.6070 3.4965 1.6330 4.5900 ;
      RECT 1.4990 3.4965 1.5250 4.5900 ;
      RECT 1.3910 3.4965 1.4170 4.5900 ;
      RECT 1.2830 3.4965 1.3090 4.5900 ;
      RECT 1.1750 3.4965 1.2010 4.5900 ;
      RECT 1.0670 3.4965 1.0930 4.5900 ;
      RECT 0.9590 3.4965 0.9850 4.5900 ;
      RECT 0.8510 3.4965 0.8770 4.5900 ;
      RECT 0.7430 3.4965 0.7690 4.5900 ;
      RECT 0.6350 3.4965 0.6610 4.5900 ;
      RECT 0.5270 3.4965 0.5530 4.5900 ;
      RECT 0.4190 3.4965 0.4450 4.5900 ;
      RECT 0.3110 3.4965 0.3370 4.5900 ;
      RECT 0.2030 3.4965 0.2290 4.5900 ;
      RECT 0.0000 3.4965 0.0850 4.5900 ;
      RECT 5.1800 4.5765 5.3080 5.6700 ;
      RECT 5.1660 5.2420 5.3080 5.5645 ;
      RECT 5.0180 4.9690 5.0800 5.6700 ;
      RECT 5.0040 5.2785 5.0800 5.4320 ;
      RECT 5.0180 4.5765 5.0440 5.6700 ;
      RECT 5.0180 4.6975 5.0580 4.9370 ;
      RECT 5.0180 4.5765 5.0800 4.6655 ;
      RECT 4.7210 5.0270 4.9270 5.6700 ;
      RECT 4.9010 4.5765 4.9270 5.6700 ;
      RECT 4.7210 5.3040 4.9410 5.5620 ;
      RECT 4.7210 4.5765 4.8190 5.6700 ;
      RECT 4.3040 4.5765 4.3870 5.6700 ;
      RECT 4.3040 4.6650 4.4010 5.6005 ;
      RECT 9.5270 4.5765 9.6120 5.6700 ;
      RECT 9.3830 4.5765 9.4090 5.6700 ;
      RECT 9.2750 4.5765 9.3010 5.6700 ;
      RECT 9.1670 4.5765 9.1930 5.6700 ;
      RECT 9.0590 4.5765 9.0850 5.6700 ;
      RECT 8.9510 4.5765 8.9770 5.6700 ;
      RECT 8.8430 4.5765 8.8690 5.6700 ;
      RECT 8.7350 4.5765 8.7610 5.6700 ;
      RECT 8.6270 4.5765 8.6530 5.6700 ;
      RECT 8.5190 4.5765 8.5450 5.6700 ;
      RECT 8.4110 4.5765 8.4370 5.6700 ;
      RECT 8.3030 4.5765 8.3290 5.6700 ;
      RECT 8.1950 4.5765 8.2210 5.6700 ;
      RECT 8.0870 4.5765 8.1130 5.6700 ;
      RECT 7.9790 4.5765 8.0050 5.6700 ;
      RECT 7.8710 4.5765 7.8970 5.6700 ;
      RECT 7.7630 4.5765 7.7890 5.6700 ;
      RECT 7.6550 4.5765 7.6810 5.6700 ;
      RECT 7.5470 4.5765 7.5730 5.6700 ;
      RECT 7.4390 4.5765 7.4650 5.6700 ;
      RECT 7.3310 4.5765 7.3570 5.6700 ;
      RECT 7.2230 4.5765 7.2490 5.6700 ;
      RECT 7.1150 4.5765 7.1410 5.6700 ;
      RECT 7.0070 4.5765 7.0330 5.6700 ;
      RECT 6.8990 4.5765 6.9250 5.6700 ;
      RECT 6.7910 4.5765 6.8170 5.6700 ;
      RECT 6.6830 4.5765 6.7090 5.6700 ;
      RECT 6.5750 4.5765 6.6010 5.6700 ;
      RECT 6.4670 4.5765 6.4930 5.6700 ;
      RECT 6.3590 4.5765 6.3850 5.6700 ;
      RECT 6.2510 4.5765 6.2770 5.6700 ;
      RECT 6.1430 4.5765 6.1690 5.6700 ;
      RECT 6.0350 4.5765 6.0610 5.6700 ;
      RECT 5.9270 4.5765 5.9530 5.6700 ;
      RECT 5.7140 4.5765 5.7910 5.6700 ;
      RECT 3.8210 4.5765 3.8980 5.6700 ;
      RECT 3.6590 4.5765 3.6850 5.6700 ;
      RECT 3.5510 4.5765 3.5770 5.6700 ;
      RECT 3.4430 4.5765 3.4690 5.6700 ;
      RECT 3.3350 4.5765 3.3610 5.6700 ;
      RECT 3.2270 4.5765 3.2530 5.6700 ;
      RECT 3.1190 4.5765 3.1450 5.6700 ;
      RECT 3.0110 4.5765 3.0370 5.6700 ;
      RECT 2.9030 4.5765 2.9290 5.6700 ;
      RECT 2.7950 4.5765 2.8210 5.6700 ;
      RECT 2.6870 4.5765 2.7130 5.6700 ;
      RECT 2.5790 4.5765 2.6050 5.6700 ;
      RECT 2.4710 4.5765 2.4970 5.6700 ;
      RECT 2.3630 4.5765 2.3890 5.6700 ;
      RECT 2.2550 4.5765 2.2810 5.6700 ;
      RECT 2.1470 4.5765 2.1730 5.6700 ;
      RECT 2.0390 4.5765 2.0650 5.6700 ;
      RECT 1.9310 4.5765 1.9570 5.6700 ;
      RECT 1.8230 4.5765 1.8490 5.6700 ;
      RECT 1.7150 4.5765 1.7410 5.6700 ;
      RECT 1.6070 4.5765 1.6330 5.6700 ;
      RECT 1.4990 4.5765 1.5250 5.6700 ;
      RECT 1.3910 4.5765 1.4170 5.6700 ;
      RECT 1.2830 4.5765 1.3090 5.6700 ;
      RECT 1.1750 4.5765 1.2010 5.6700 ;
      RECT 1.0670 4.5765 1.0930 5.6700 ;
      RECT 0.9590 4.5765 0.9850 5.6700 ;
      RECT 0.8510 4.5765 0.8770 5.6700 ;
      RECT 0.7430 4.5765 0.7690 5.6700 ;
      RECT 0.6350 4.5765 0.6610 5.6700 ;
      RECT 0.5270 4.5765 0.5530 5.6700 ;
      RECT 0.4190 4.5765 0.4450 5.6700 ;
      RECT 0.3110 4.5765 0.3370 5.6700 ;
      RECT 0.2030 4.5765 0.2290 5.6700 ;
      RECT 0.0000 4.5765 0.0850 5.6700 ;
      RECT 5.1800 5.6565 5.3080 6.7500 ;
      RECT 5.1660 6.3220 5.3080 6.6445 ;
      RECT 5.0180 6.0490 5.0800 6.7500 ;
      RECT 5.0040 6.3585 5.0800 6.5120 ;
      RECT 5.0180 5.6565 5.0440 6.7500 ;
      RECT 5.0180 5.7775 5.0580 6.0170 ;
      RECT 5.0180 5.6565 5.0800 5.7455 ;
      RECT 4.7210 6.1070 4.9270 6.7500 ;
      RECT 4.9010 5.6565 4.9270 6.7500 ;
      RECT 4.7210 6.3840 4.9410 6.6420 ;
      RECT 4.7210 5.6565 4.8190 6.7500 ;
      RECT 4.3040 5.6565 4.3870 6.7500 ;
      RECT 4.3040 5.7450 4.4010 6.6805 ;
      RECT 9.5270 5.6565 9.6120 6.7500 ;
      RECT 9.3830 5.6565 9.4090 6.7500 ;
      RECT 9.2750 5.6565 9.3010 6.7500 ;
      RECT 9.1670 5.6565 9.1930 6.7500 ;
      RECT 9.0590 5.6565 9.0850 6.7500 ;
      RECT 8.9510 5.6565 8.9770 6.7500 ;
      RECT 8.8430 5.6565 8.8690 6.7500 ;
      RECT 8.7350 5.6565 8.7610 6.7500 ;
      RECT 8.6270 5.6565 8.6530 6.7500 ;
      RECT 8.5190 5.6565 8.5450 6.7500 ;
      RECT 8.4110 5.6565 8.4370 6.7500 ;
      RECT 8.3030 5.6565 8.3290 6.7500 ;
      RECT 8.1950 5.6565 8.2210 6.7500 ;
      RECT 8.0870 5.6565 8.1130 6.7500 ;
      RECT 7.9790 5.6565 8.0050 6.7500 ;
      RECT 7.8710 5.6565 7.8970 6.7500 ;
      RECT 7.7630 5.6565 7.7890 6.7500 ;
      RECT 7.6550 5.6565 7.6810 6.7500 ;
      RECT 7.5470 5.6565 7.5730 6.7500 ;
      RECT 7.4390 5.6565 7.4650 6.7500 ;
      RECT 7.3310 5.6565 7.3570 6.7500 ;
      RECT 7.2230 5.6565 7.2490 6.7500 ;
      RECT 7.1150 5.6565 7.1410 6.7500 ;
      RECT 7.0070 5.6565 7.0330 6.7500 ;
      RECT 6.8990 5.6565 6.9250 6.7500 ;
      RECT 6.7910 5.6565 6.8170 6.7500 ;
      RECT 6.6830 5.6565 6.7090 6.7500 ;
      RECT 6.5750 5.6565 6.6010 6.7500 ;
      RECT 6.4670 5.6565 6.4930 6.7500 ;
      RECT 6.3590 5.6565 6.3850 6.7500 ;
      RECT 6.2510 5.6565 6.2770 6.7500 ;
      RECT 6.1430 5.6565 6.1690 6.7500 ;
      RECT 6.0350 5.6565 6.0610 6.7500 ;
      RECT 5.9270 5.6565 5.9530 6.7500 ;
      RECT 5.7140 5.6565 5.7910 6.7500 ;
      RECT 3.8210 5.6565 3.8980 6.7500 ;
      RECT 3.6590 5.6565 3.6850 6.7500 ;
      RECT 3.5510 5.6565 3.5770 6.7500 ;
      RECT 3.4430 5.6565 3.4690 6.7500 ;
      RECT 3.3350 5.6565 3.3610 6.7500 ;
      RECT 3.2270 5.6565 3.2530 6.7500 ;
      RECT 3.1190 5.6565 3.1450 6.7500 ;
      RECT 3.0110 5.6565 3.0370 6.7500 ;
      RECT 2.9030 5.6565 2.9290 6.7500 ;
      RECT 2.7950 5.6565 2.8210 6.7500 ;
      RECT 2.6870 5.6565 2.7130 6.7500 ;
      RECT 2.5790 5.6565 2.6050 6.7500 ;
      RECT 2.4710 5.6565 2.4970 6.7500 ;
      RECT 2.3630 5.6565 2.3890 6.7500 ;
      RECT 2.2550 5.6565 2.2810 6.7500 ;
      RECT 2.1470 5.6565 2.1730 6.7500 ;
      RECT 2.0390 5.6565 2.0650 6.7500 ;
      RECT 1.9310 5.6565 1.9570 6.7500 ;
      RECT 1.8230 5.6565 1.8490 6.7500 ;
      RECT 1.7150 5.6565 1.7410 6.7500 ;
      RECT 1.6070 5.6565 1.6330 6.7500 ;
      RECT 1.4990 5.6565 1.5250 6.7500 ;
      RECT 1.3910 5.6565 1.4170 6.7500 ;
      RECT 1.2830 5.6565 1.3090 6.7500 ;
      RECT 1.1750 5.6565 1.2010 6.7500 ;
      RECT 1.0670 5.6565 1.0930 6.7500 ;
      RECT 0.9590 5.6565 0.9850 6.7500 ;
      RECT 0.8510 5.6565 0.8770 6.7500 ;
      RECT 0.7430 5.6565 0.7690 6.7500 ;
      RECT 0.6350 5.6565 0.6610 6.7500 ;
      RECT 0.5270 5.6565 0.5530 6.7500 ;
      RECT 0.4190 5.6565 0.4450 6.7500 ;
      RECT 0.3110 5.6565 0.3370 6.7500 ;
      RECT 0.2030 5.6565 0.2290 6.7500 ;
      RECT 0.0000 5.6565 0.0850 6.7500 ;
      RECT 5.1800 6.7365 5.3080 7.8300 ;
      RECT 5.1660 7.4020 5.3080 7.7245 ;
      RECT 5.0180 7.1290 5.0800 7.8300 ;
      RECT 5.0040 7.4385 5.0800 7.5920 ;
      RECT 5.0180 6.7365 5.0440 7.8300 ;
      RECT 5.0180 6.8575 5.0580 7.0970 ;
      RECT 5.0180 6.7365 5.0800 6.8255 ;
      RECT 4.7210 7.1870 4.9270 7.8300 ;
      RECT 4.9010 6.7365 4.9270 7.8300 ;
      RECT 4.7210 7.4640 4.9410 7.7220 ;
      RECT 4.7210 6.7365 4.8190 7.8300 ;
      RECT 4.3040 6.7365 4.3870 7.8300 ;
      RECT 4.3040 6.8250 4.4010 7.7605 ;
      RECT 9.5270 6.7365 9.6120 7.8300 ;
      RECT 9.3830 6.7365 9.4090 7.8300 ;
      RECT 9.2750 6.7365 9.3010 7.8300 ;
      RECT 9.1670 6.7365 9.1930 7.8300 ;
      RECT 9.0590 6.7365 9.0850 7.8300 ;
      RECT 8.9510 6.7365 8.9770 7.8300 ;
      RECT 8.8430 6.7365 8.8690 7.8300 ;
      RECT 8.7350 6.7365 8.7610 7.8300 ;
      RECT 8.6270 6.7365 8.6530 7.8300 ;
      RECT 8.5190 6.7365 8.5450 7.8300 ;
      RECT 8.4110 6.7365 8.4370 7.8300 ;
      RECT 8.3030 6.7365 8.3290 7.8300 ;
      RECT 8.1950 6.7365 8.2210 7.8300 ;
      RECT 8.0870 6.7365 8.1130 7.8300 ;
      RECT 7.9790 6.7365 8.0050 7.8300 ;
      RECT 7.8710 6.7365 7.8970 7.8300 ;
      RECT 7.7630 6.7365 7.7890 7.8300 ;
      RECT 7.6550 6.7365 7.6810 7.8300 ;
      RECT 7.5470 6.7365 7.5730 7.8300 ;
      RECT 7.4390 6.7365 7.4650 7.8300 ;
      RECT 7.3310 6.7365 7.3570 7.8300 ;
      RECT 7.2230 6.7365 7.2490 7.8300 ;
      RECT 7.1150 6.7365 7.1410 7.8300 ;
      RECT 7.0070 6.7365 7.0330 7.8300 ;
      RECT 6.8990 6.7365 6.9250 7.8300 ;
      RECT 6.7910 6.7365 6.8170 7.8300 ;
      RECT 6.6830 6.7365 6.7090 7.8300 ;
      RECT 6.5750 6.7365 6.6010 7.8300 ;
      RECT 6.4670 6.7365 6.4930 7.8300 ;
      RECT 6.3590 6.7365 6.3850 7.8300 ;
      RECT 6.2510 6.7365 6.2770 7.8300 ;
      RECT 6.1430 6.7365 6.1690 7.8300 ;
      RECT 6.0350 6.7365 6.0610 7.8300 ;
      RECT 5.9270 6.7365 5.9530 7.8300 ;
      RECT 5.7140 6.7365 5.7910 7.8300 ;
      RECT 3.8210 6.7365 3.8980 7.8300 ;
      RECT 3.6590 6.7365 3.6850 7.8300 ;
      RECT 3.5510 6.7365 3.5770 7.8300 ;
      RECT 3.4430 6.7365 3.4690 7.8300 ;
      RECT 3.3350 6.7365 3.3610 7.8300 ;
      RECT 3.2270 6.7365 3.2530 7.8300 ;
      RECT 3.1190 6.7365 3.1450 7.8300 ;
      RECT 3.0110 6.7365 3.0370 7.8300 ;
      RECT 2.9030 6.7365 2.9290 7.8300 ;
      RECT 2.7950 6.7365 2.8210 7.8300 ;
      RECT 2.6870 6.7365 2.7130 7.8300 ;
      RECT 2.5790 6.7365 2.6050 7.8300 ;
      RECT 2.4710 6.7365 2.4970 7.8300 ;
      RECT 2.3630 6.7365 2.3890 7.8300 ;
      RECT 2.2550 6.7365 2.2810 7.8300 ;
      RECT 2.1470 6.7365 2.1730 7.8300 ;
      RECT 2.0390 6.7365 2.0650 7.8300 ;
      RECT 1.9310 6.7365 1.9570 7.8300 ;
      RECT 1.8230 6.7365 1.8490 7.8300 ;
      RECT 1.7150 6.7365 1.7410 7.8300 ;
      RECT 1.6070 6.7365 1.6330 7.8300 ;
      RECT 1.4990 6.7365 1.5250 7.8300 ;
      RECT 1.3910 6.7365 1.4170 7.8300 ;
      RECT 1.2830 6.7365 1.3090 7.8300 ;
      RECT 1.1750 6.7365 1.2010 7.8300 ;
      RECT 1.0670 6.7365 1.0930 7.8300 ;
      RECT 0.9590 6.7365 0.9850 7.8300 ;
      RECT 0.8510 6.7365 0.8770 7.8300 ;
      RECT 0.7430 6.7365 0.7690 7.8300 ;
      RECT 0.6350 6.7365 0.6610 7.8300 ;
      RECT 0.5270 6.7365 0.5530 7.8300 ;
      RECT 0.4190 6.7365 0.4450 7.8300 ;
      RECT 0.3110 6.7365 0.3370 7.8300 ;
      RECT 0.2030 6.7365 0.2290 7.8300 ;
      RECT 0.0000 6.7365 0.0850 7.8300 ;
      RECT 5.1800 7.8165 5.3080 8.9100 ;
      RECT 5.1660 8.4820 5.3080 8.8045 ;
      RECT 5.0180 8.2090 5.0800 8.9100 ;
      RECT 5.0040 8.5185 5.0800 8.6720 ;
      RECT 5.0180 7.8165 5.0440 8.9100 ;
      RECT 5.0180 7.9375 5.0580 8.1770 ;
      RECT 5.0180 7.8165 5.0800 7.9055 ;
      RECT 4.7210 8.2670 4.9270 8.9100 ;
      RECT 4.9010 7.8165 4.9270 8.9100 ;
      RECT 4.7210 8.5440 4.9410 8.8020 ;
      RECT 4.7210 7.8165 4.8190 8.9100 ;
      RECT 4.3040 7.8165 4.3870 8.9100 ;
      RECT 4.3040 7.9050 4.4010 8.8405 ;
      RECT 9.5270 7.8165 9.6120 8.9100 ;
      RECT 9.3830 7.8165 9.4090 8.9100 ;
      RECT 9.2750 7.8165 9.3010 8.9100 ;
      RECT 9.1670 7.8165 9.1930 8.9100 ;
      RECT 9.0590 7.8165 9.0850 8.9100 ;
      RECT 8.9510 7.8165 8.9770 8.9100 ;
      RECT 8.8430 7.8165 8.8690 8.9100 ;
      RECT 8.7350 7.8165 8.7610 8.9100 ;
      RECT 8.6270 7.8165 8.6530 8.9100 ;
      RECT 8.5190 7.8165 8.5450 8.9100 ;
      RECT 8.4110 7.8165 8.4370 8.9100 ;
      RECT 8.3030 7.8165 8.3290 8.9100 ;
      RECT 8.1950 7.8165 8.2210 8.9100 ;
      RECT 8.0870 7.8165 8.1130 8.9100 ;
      RECT 7.9790 7.8165 8.0050 8.9100 ;
      RECT 7.8710 7.8165 7.8970 8.9100 ;
      RECT 7.7630 7.8165 7.7890 8.9100 ;
      RECT 7.6550 7.8165 7.6810 8.9100 ;
      RECT 7.5470 7.8165 7.5730 8.9100 ;
      RECT 7.4390 7.8165 7.4650 8.9100 ;
      RECT 7.3310 7.8165 7.3570 8.9100 ;
      RECT 7.2230 7.8165 7.2490 8.9100 ;
      RECT 7.1150 7.8165 7.1410 8.9100 ;
      RECT 7.0070 7.8165 7.0330 8.9100 ;
      RECT 6.8990 7.8165 6.9250 8.9100 ;
      RECT 6.7910 7.8165 6.8170 8.9100 ;
      RECT 6.6830 7.8165 6.7090 8.9100 ;
      RECT 6.5750 7.8165 6.6010 8.9100 ;
      RECT 6.4670 7.8165 6.4930 8.9100 ;
      RECT 6.3590 7.8165 6.3850 8.9100 ;
      RECT 6.2510 7.8165 6.2770 8.9100 ;
      RECT 6.1430 7.8165 6.1690 8.9100 ;
      RECT 6.0350 7.8165 6.0610 8.9100 ;
      RECT 5.9270 7.8165 5.9530 8.9100 ;
      RECT 5.7140 7.8165 5.7910 8.9100 ;
      RECT 3.8210 7.8165 3.8980 8.9100 ;
      RECT 3.6590 7.8165 3.6850 8.9100 ;
      RECT 3.5510 7.8165 3.5770 8.9100 ;
      RECT 3.4430 7.8165 3.4690 8.9100 ;
      RECT 3.3350 7.8165 3.3610 8.9100 ;
      RECT 3.2270 7.8165 3.2530 8.9100 ;
      RECT 3.1190 7.8165 3.1450 8.9100 ;
      RECT 3.0110 7.8165 3.0370 8.9100 ;
      RECT 2.9030 7.8165 2.9290 8.9100 ;
      RECT 2.7950 7.8165 2.8210 8.9100 ;
      RECT 2.6870 7.8165 2.7130 8.9100 ;
      RECT 2.5790 7.8165 2.6050 8.9100 ;
      RECT 2.4710 7.8165 2.4970 8.9100 ;
      RECT 2.3630 7.8165 2.3890 8.9100 ;
      RECT 2.2550 7.8165 2.2810 8.9100 ;
      RECT 2.1470 7.8165 2.1730 8.9100 ;
      RECT 2.0390 7.8165 2.0650 8.9100 ;
      RECT 1.9310 7.8165 1.9570 8.9100 ;
      RECT 1.8230 7.8165 1.8490 8.9100 ;
      RECT 1.7150 7.8165 1.7410 8.9100 ;
      RECT 1.6070 7.8165 1.6330 8.9100 ;
      RECT 1.4990 7.8165 1.5250 8.9100 ;
      RECT 1.3910 7.8165 1.4170 8.9100 ;
      RECT 1.2830 7.8165 1.3090 8.9100 ;
      RECT 1.1750 7.8165 1.2010 8.9100 ;
      RECT 1.0670 7.8165 1.0930 8.9100 ;
      RECT 0.9590 7.8165 0.9850 8.9100 ;
      RECT 0.8510 7.8165 0.8770 8.9100 ;
      RECT 0.7430 7.8165 0.7690 8.9100 ;
      RECT 0.6350 7.8165 0.6610 8.9100 ;
      RECT 0.5270 7.8165 0.5530 8.9100 ;
      RECT 0.4190 7.8165 0.4450 8.9100 ;
      RECT 0.3110 7.8165 0.3370 8.9100 ;
      RECT 0.2030 7.8165 0.2290 8.9100 ;
      RECT 0.0000 7.8165 0.0850 8.9100 ;
      RECT 5.1800 8.8965 5.3080 9.9900 ;
      RECT 5.1660 9.5620 5.3080 9.8845 ;
      RECT 5.0180 9.2890 5.0800 9.9900 ;
      RECT 5.0040 9.5985 5.0800 9.7520 ;
      RECT 5.0180 8.8965 5.0440 9.9900 ;
      RECT 5.0180 9.0175 5.0580 9.2570 ;
      RECT 5.0180 8.8965 5.0800 8.9855 ;
      RECT 4.7210 9.3470 4.9270 9.9900 ;
      RECT 4.9010 8.8965 4.9270 9.9900 ;
      RECT 4.7210 9.6240 4.9410 9.8820 ;
      RECT 4.7210 8.8965 4.8190 9.9900 ;
      RECT 4.3040 8.8965 4.3870 9.9900 ;
      RECT 4.3040 8.9850 4.4010 9.9205 ;
      RECT 9.5270 8.8965 9.6120 9.9900 ;
      RECT 9.3830 8.8965 9.4090 9.9900 ;
      RECT 9.2750 8.8965 9.3010 9.9900 ;
      RECT 9.1670 8.8965 9.1930 9.9900 ;
      RECT 9.0590 8.8965 9.0850 9.9900 ;
      RECT 8.9510 8.8965 8.9770 9.9900 ;
      RECT 8.8430 8.8965 8.8690 9.9900 ;
      RECT 8.7350 8.8965 8.7610 9.9900 ;
      RECT 8.6270 8.8965 8.6530 9.9900 ;
      RECT 8.5190 8.8965 8.5450 9.9900 ;
      RECT 8.4110 8.8965 8.4370 9.9900 ;
      RECT 8.3030 8.8965 8.3290 9.9900 ;
      RECT 8.1950 8.8965 8.2210 9.9900 ;
      RECT 8.0870 8.8965 8.1130 9.9900 ;
      RECT 7.9790 8.8965 8.0050 9.9900 ;
      RECT 7.8710 8.8965 7.8970 9.9900 ;
      RECT 7.7630 8.8965 7.7890 9.9900 ;
      RECT 7.6550 8.8965 7.6810 9.9900 ;
      RECT 7.5470 8.8965 7.5730 9.9900 ;
      RECT 7.4390 8.8965 7.4650 9.9900 ;
      RECT 7.3310 8.8965 7.3570 9.9900 ;
      RECT 7.2230 8.8965 7.2490 9.9900 ;
      RECT 7.1150 8.8965 7.1410 9.9900 ;
      RECT 7.0070 8.8965 7.0330 9.9900 ;
      RECT 6.8990 8.8965 6.9250 9.9900 ;
      RECT 6.7910 8.8965 6.8170 9.9900 ;
      RECT 6.6830 8.8965 6.7090 9.9900 ;
      RECT 6.5750 8.8965 6.6010 9.9900 ;
      RECT 6.4670 8.8965 6.4930 9.9900 ;
      RECT 6.3590 8.8965 6.3850 9.9900 ;
      RECT 6.2510 8.8965 6.2770 9.9900 ;
      RECT 6.1430 8.8965 6.1690 9.9900 ;
      RECT 6.0350 8.8965 6.0610 9.9900 ;
      RECT 5.9270 8.8965 5.9530 9.9900 ;
      RECT 5.7140 8.8965 5.7910 9.9900 ;
      RECT 3.8210 8.8965 3.8980 9.9900 ;
      RECT 3.6590 8.8965 3.6850 9.9900 ;
      RECT 3.5510 8.8965 3.5770 9.9900 ;
      RECT 3.4430 8.8965 3.4690 9.9900 ;
      RECT 3.3350 8.8965 3.3610 9.9900 ;
      RECT 3.2270 8.8965 3.2530 9.9900 ;
      RECT 3.1190 8.8965 3.1450 9.9900 ;
      RECT 3.0110 8.8965 3.0370 9.9900 ;
      RECT 2.9030 8.8965 2.9290 9.9900 ;
      RECT 2.7950 8.8965 2.8210 9.9900 ;
      RECT 2.6870 8.8965 2.7130 9.9900 ;
      RECT 2.5790 8.8965 2.6050 9.9900 ;
      RECT 2.4710 8.8965 2.4970 9.9900 ;
      RECT 2.3630 8.8965 2.3890 9.9900 ;
      RECT 2.2550 8.8965 2.2810 9.9900 ;
      RECT 2.1470 8.8965 2.1730 9.9900 ;
      RECT 2.0390 8.8965 2.0650 9.9900 ;
      RECT 1.9310 8.8965 1.9570 9.9900 ;
      RECT 1.8230 8.8965 1.8490 9.9900 ;
      RECT 1.7150 8.8965 1.7410 9.9900 ;
      RECT 1.6070 8.8965 1.6330 9.9900 ;
      RECT 1.4990 8.8965 1.5250 9.9900 ;
      RECT 1.3910 8.8965 1.4170 9.9900 ;
      RECT 1.2830 8.8965 1.3090 9.9900 ;
      RECT 1.1750 8.8965 1.2010 9.9900 ;
      RECT 1.0670 8.8965 1.0930 9.9900 ;
      RECT 0.9590 8.8965 0.9850 9.9900 ;
      RECT 0.8510 8.8965 0.8770 9.9900 ;
      RECT 0.7430 8.8965 0.7690 9.9900 ;
      RECT 0.6350 8.8965 0.6610 9.9900 ;
      RECT 0.5270 8.8965 0.5530 9.9900 ;
      RECT 0.4190 8.8965 0.4450 9.9900 ;
      RECT 0.3110 8.8965 0.3370 9.9900 ;
      RECT 0.2030 8.8965 0.2290 9.9900 ;
      RECT 0.0000 8.8965 0.0850 9.9900 ;
      RECT 5.1800 9.9765 5.3080 11.0700 ;
      RECT 5.1660 10.6420 5.3080 10.9645 ;
      RECT 5.0180 10.3690 5.0800 11.0700 ;
      RECT 5.0040 10.6785 5.0800 10.8320 ;
      RECT 5.0180 9.9765 5.0440 11.0700 ;
      RECT 5.0180 10.0975 5.0580 10.3370 ;
      RECT 5.0180 9.9765 5.0800 10.0655 ;
      RECT 4.7210 10.4270 4.9270 11.0700 ;
      RECT 4.9010 9.9765 4.9270 11.0700 ;
      RECT 4.7210 10.7040 4.9410 10.9620 ;
      RECT 4.7210 9.9765 4.8190 11.0700 ;
      RECT 4.3040 9.9765 4.3870 11.0700 ;
      RECT 4.3040 10.0650 4.4010 11.0005 ;
      RECT 9.5270 9.9765 9.6120 11.0700 ;
      RECT 9.3830 9.9765 9.4090 11.0700 ;
      RECT 9.2750 9.9765 9.3010 11.0700 ;
      RECT 9.1670 9.9765 9.1930 11.0700 ;
      RECT 9.0590 9.9765 9.0850 11.0700 ;
      RECT 8.9510 9.9765 8.9770 11.0700 ;
      RECT 8.8430 9.9765 8.8690 11.0700 ;
      RECT 8.7350 9.9765 8.7610 11.0700 ;
      RECT 8.6270 9.9765 8.6530 11.0700 ;
      RECT 8.5190 9.9765 8.5450 11.0700 ;
      RECT 8.4110 9.9765 8.4370 11.0700 ;
      RECT 8.3030 9.9765 8.3290 11.0700 ;
      RECT 8.1950 9.9765 8.2210 11.0700 ;
      RECT 8.0870 9.9765 8.1130 11.0700 ;
      RECT 7.9790 9.9765 8.0050 11.0700 ;
      RECT 7.8710 9.9765 7.8970 11.0700 ;
      RECT 7.7630 9.9765 7.7890 11.0700 ;
      RECT 7.6550 9.9765 7.6810 11.0700 ;
      RECT 7.5470 9.9765 7.5730 11.0700 ;
      RECT 7.4390 9.9765 7.4650 11.0700 ;
      RECT 7.3310 9.9765 7.3570 11.0700 ;
      RECT 7.2230 9.9765 7.2490 11.0700 ;
      RECT 7.1150 9.9765 7.1410 11.0700 ;
      RECT 7.0070 9.9765 7.0330 11.0700 ;
      RECT 6.8990 9.9765 6.9250 11.0700 ;
      RECT 6.7910 9.9765 6.8170 11.0700 ;
      RECT 6.6830 9.9765 6.7090 11.0700 ;
      RECT 6.5750 9.9765 6.6010 11.0700 ;
      RECT 6.4670 9.9765 6.4930 11.0700 ;
      RECT 6.3590 9.9765 6.3850 11.0700 ;
      RECT 6.2510 9.9765 6.2770 11.0700 ;
      RECT 6.1430 9.9765 6.1690 11.0700 ;
      RECT 6.0350 9.9765 6.0610 11.0700 ;
      RECT 5.9270 9.9765 5.9530 11.0700 ;
      RECT 5.7140 9.9765 5.7910 11.0700 ;
      RECT 3.8210 9.9765 3.8980 11.0700 ;
      RECT 3.6590 9.9765 3.6850 11.0700 ;
      RECT 3.5510 9.9765 3.5770 11.0700 ;
      RECT 3.4430 9.9765 3.4690 11.0700 ;
      RECT 3.3350 9.9765 3.3610 11.0700 ;
      RECT 3.2270 9.9765 3.2530 11.0700 ;
      RECT 3.1190 9.9765 3.1450 11.0700 ;
      RECT 3.0110 9.9765 3.0370 11.0700 ;
      RECT 2.9030 9.9765 2.9290 11.0700 ;
      RECT 2.7950 9.9765 2.8210 11.0700 ;
      RECT 2.6870 9.9765 2.7130 11.0700 ;
      RECT 2.5790 9.9765 2.6050 11.0700 ;
      RECT 2.4710 9.9765 2.4970 11.0700 ;
      RECT 2.3630 9.9765 2.3890 11.0700 ;
      RECT 2.2550 9.9765 2.2810 11.0700 ;
      RECT 2.1470 9.9765 2.1730 11.0700 ;
      RECT 2.0390 9.9765 2.0650 11.0700 ;
      RECT 1.9310 9.9765 1.9570 11.0700 ;
      RECT 1.8230 9.9765 1.8490 11.0700 ;
      RECT 1.7150 9.9765 1.7410 11.0700 ;
      RECT 1.6070 9.9765 1.6330 11.0700 ;
      RECT 1.4990 9.9765 1.5250 11.0700 ;
      RECT 1.3910 9.9765 1.4170 11.0700 ;
      RECT 1.2830 9.9765 1.3090 11.0700 ;
      RECT 1.1750 9.9765 1.2010 11.0700 ;
      RECT 1.0670 9.9765 1.0930 11.0700 ;
      RECT 0.9590 9.9765 0.9850 11.0700 ;
      RECT 0.8510 9.9765 0.8770 11.0700 ;
      RECT 0.7430 9.9765 0.7690 11.0700 ;
      RECT 0.6350 9.9765 0.6610 11.0700 ;
      RECT 0.5270 9.9765 0.5530 11.0700 ;
      RECT 0.4190 9.9765 0.4450 11.0700 ;
      RECT 0.3110 9.9765 0.3370 11.0700 ;
      RECT 0.2030 9.9765 0.2290 11.0700 ;
      RECT 0.0000 9.9765 0.0850 11.0700 ;
      RECT 5.1800 11.0565 5.3080 12.1500 ;
      RECT 5.1660 11.7220 5.3080 12.0445 ;
      RECT 5.0180 11.4490 5.0800 12.1500 ;
      RECT 5.0040 11.7585 5.0800 11.9120 ;
      RECT 5.0180 11.0565 5.0440 12.1500 ;
      RECT 5.0180 11.1775 5.0580 11.4170 ;
      RECT 5.0180 11.0565 5.0800 11.1455 ;
      RECT 4.7210 11.5070 4.9270 12.1500 ;
      RECT 4.9010 11.0565 4.9270 12.1500 ;
      RECT 4.7210 11.7840 4.9410 12.0420 ;
      RECT 4.7210 11.0565 4.8190 12.1500 ;
      RECT 4.3040 11.0565 4.3870 12.1500 ;
      RECT 4.3040 11.1450 4.4010 12.0805 ;
      RECT 9.5270 11.0565 9.6120 12.1500 ;
      RECT 9.3830 11.0565 9.4090 12.1500 ;
      RECT 9.2750 11.0565 9.3010 12.1500 ;
      RECT 9.1670 11.0565 9.1930 12.1500 ;
      RECT 9.0590 11.0565 9.0850 12.1500 ;
      RECT 8.9510 11.0565 8.9770 12.1500 ;
      RECT 8.8430 11.0565 8.8690 12.1500 ;
      RECT 8.7350 11.0565 8.7610 12.1500 ;
      RECT 8.6270 11.0565 8.6530 12.1500 ;
      RECT 8.5190 11.0565 8.5450 12.1500 ;
      RECT 8.4110 11.0565 8.4370 12.1500 ;
      RECT 8.3030 11.0565 8.3290 12.1500 ;
      RECT 8.1950 11.0565 8.2210 12.1500 ;
      RECT 8.0870 11.0565 8.1130 12.1500 ;
      RECT 7.9790 11.0565 8.0050 12.1500 ;
      RECT 7.8710 11.0565 7.8970 12.1500 ;
      RECT 7.7630 11.0565 7.7890 12.1500 ;
      RECT 7.6550 11.0565 7.6810 12.1500 ;
      RECT 7.5470 11.0565 7.5730 12.1500 ;
      RECT 7.4390 11.0565 7.4650 12.1500 ;
      RECT 7.3310 11.0565 7.3570 12.1500 ;
      RECT 7.2230 11.0565 7.2490 12.1500 ;
      RECT 7.1150 11.0565 7.1410 12.1500 ;
      RECT 7.0070 11.0565 7.0330 12.1500 ;
      RECT 6.8990 11.0565 6.9250 12.1500 ;
      RECT 6.7910 11.0565 6.8170 12.1500 ;
      RECT 6.6830 11.0565 6.7090 12.1500 ;
      RECT 6.5750 11.0565 6.6010 12.1500 ;
      RECT 6.4670 11.0565 6.4930 12.1500 ;
      RECT 6.3590 11.0565 6.3850 12.1500 ;
      RECT 6.2510 11.0565 6.2770 12.1500 ;
      RECT 6.1430 11.0565 6.1690 12.1500 ;
      RECT 6.0350 11.0565 6.0610 12.1500 ;
      RECT 5.9270 11.0565 5.9530 12.1500 ;
      RECT 5.7140 11.0565 5.7910 12.1500 ;
      RECT 3.8210 11.0565 3.8980 12.1500 ;
      RECT 3.6590 11.0565 3.6850 12.1500 ;
      RECT 3.5510 11.0565 3.5770 12.1500 ;
      RECT 3.4430 11.0565 3.4690 12.1500 ;
      RECT 3.3350 11.0565 3.3610 12.1500 ;
      RECT 3.2270 11.0565 3.2530 12.1500 ;
      RECT 3.1190 11.0565 3.1450 12.1500 ;
      RECT 3.0110 11.0565 3.0370 12.1500 ;
      RECT 2.9030 11.0565 2.9290 12.1500 ;
      RECT 2.7950 11.0565 2.8210 12.1500 ;
      RECT 2.6870 11.0565 2.7130 12.1500 ;
      RECT 2.5790 11.0565 2.6050 12.1500 ;
      RECT 2.4710 11.0565 2.4970 12.1500 ;
      RECT 2.3630 11.0565 2.3890 12.1500 ;
      RECT 2.2550 11.0565 2.2810 12.1500 ;
      RECT 2.1470 11.0565 2.1730 12.1500 ;
      RECT 2.0390 11.0565 2.0650 12.1500 ;
      RECT 1.9310 11.0565 1.9570 12.1500 ;
      RECT 1.8230 11.0565 1.8490 12.1500 ;
      RECT 1.7150 11.0565 1.7410 12.1500 ;
      RECT 1.6070 11.0565 1.6330 12.1500 ;
      RECT 1.4990 11.0565 1.5250 12.1500 ;
      RECT 1.3910 11.0565 1.4170 12.1500 ;
      RECT 1.2830 11.0565 1.3090 12.1500 ;
      RECT 1.1750 11.0565 1.2010 12.1500 ;
      RECT 1.0670 11.0565 1.0930 12.1500 ;
      RECT 0.9590 11.0565 0.9850 12.1500 ;
      RECT 0.8510 11.0565 0.8770 12.1500 ;
      RECT 0.7430 11.0565 0.7690 12.1500 ;
      RECT 0.6350 11.0565 0.6610 12.1500 ;
      RECT 0.5270 11.0565 0.5530 12.1500 ;
      RECT 0.4190 11.0565 0.4450 12.1500 ;
      RECT 0.3110 11.0565 0.3370 12.1500 ;
      RECT 0.2030 11.0565 0.2290 12.1500 ;
      RECT 0.0000 11.0565 0.0850 12.1500 ;
      RECT 5.1800 12.1365 5.3080 13.2300 ;
      RECT 5.1660 12.8020 5.3080 13.1245 ;
      RECT 5.0180 12.5290 5.0800 13.2300 ;
      RECT 5.0040 12.8385 5.0800 12.9920 ;
      RECT 5.0180 12.1365 5.0440 13.2300 ;
      RECT 5.0180 12.2575 5.0580 12.4970 ;
      RECT 5.0180 12.1365 5.0800 12.2255 ;
      RECT 4.7210 12.5870 4.9270 13.2300 ;
      RECT 4.9010 12.1365 4.9270 13.2300 ;
      RECT 4.7210 12.8640 4.9410 13.1220 ;
      RECT 4.7210 12.1365 4.8190 13.2300 ;
      RECT 4.3040 12.1365 4.3870 13.2300 ;
      RECT 4.3040 12.2250 4.4010 13.1605 ;
      RECT 9.5270 12.1365 9.6120 13.2300 ;
      RECT 9.3830 12.1365 9.4090 13.2300 ;
      RECT 9.2750 12.1365 9.3010 13.2300 ;
      RECT 9.1670 12.1365 9.1930 13.2300 ;
      RECT 9.0590 12.1365 9.0850 13.2300 ;
      RECT 8.9510 12.1365 8.9770 13.2300 ;
      RECT 8.8430 12.1365 8.8690 13.2300 ;
      RECT 8.7350 12.1365 8.7610 13.2300 ;
      RECT 8.6270 12.1365 8.6530 13.2300 ;
      RECT 8.5190 12.1365 8.5450 13.2300 ;
      RECT 8.4110 12.1365 8.4370 13.2300 ;
      RECT 8.3030 12.1365 8.3290 13.2300 ;
      RECT 8.1950 12.1365 8.2210 13.2300 ;
      RECT 8.0870 12.1365 8.1130 13.2300 ;
      RECT 7.9790 12.1365 8.0050 13.2300 ;
      RECT 7.8710 12.1365 7.8970 13.2300 ;
      RECT 7.7630 12.1365 7.7890 13.2300 ;
      RECT 7.6550 12.1365 7.6810 13.2300 ;
      RECT 7.5470 12.1365 7.5730 13.2300 ;
      RECT 7.4390 12.1365 7.4650 13.2300 ;
      RECT 7.3310 12.1365 7.3570 13.2300 ;
      RECT 7.2230 12.1365 7.2490 13.2300 ;
      RECT 7.1150 12.1365 7.1410 13.2300 ;
      RECT 7.0070 12.1365 7.0330 13.2300 ;
      RECT 6.8990 12.1365 6.9250 13.2300 ;
      RECT 6.7910 12.1365 6.8170 13.2300 ;
      RECT 6.6830 12.1365 6.7090 13.2300 ;
      RECT 6.5750 12.1365 6.6010 13.2300 ;
      RECT 6.4670 12.1365 6.4930 13.2300 ;
      RECT 6.3590 12.1365 6.3850 13.2300 ;
      RECT 6.2510 12.1365 6.2770 13.2300 ;
      RECT 6.1430 12.1365 6.1690 13.2300 ;
      RECT 6.0350 12.1365 6.0610 13.2300 ;
      RECT 5.9270 12.1365 5.9530 13.2300 ;
      RECT 5.7140 12.1365 5.7910 13.2300 ;
      RECT 3.8210 12.1365 3.8980 13.2300 ;
      RECT 3.6590 12.1365 3.6850 13.2300 ;
      RECT 3.5510 12.1365 3.5770 13.2300 ;
      RECT 3.4430 12.1365 3.4690 13.2300 ;
      RECT 3.3350 12.1365 3.3610 13.2300 ;
      RECT 3.2270 12.1365 3.2530 13.2300 ;
      RECT 3.1190 12.1365 3.1450 13.2300 ;
      RECT 3.0110 12.1365 3.0370 13.2300 ;
      RECT 2.9030 12.1365 2.9290 13.2300 ;
      RECT 2.7950 12.1365 2.8210 13.2300 ;
      RECT 2.6870 12.1365 2.7130 13.2300 ;
      RECT 2.5790 12.1365 2.6050 13.2300 ;
      RECT 2.4710 12.1365 2.4970 13.2300 ;
      RECT 2.3630 12.1365 2.3890 13.2300 ;
      RECT 2.2550 12.1365 2.2810 13.2300 ;
      RECT 2.1470 12.1365 2.1730 13.2300 ;
      RECT 2.0390 12.1365 2.0650 13.2300 ;
      RECT 1.9310 12.1365 1.9570 13.2300 ;
      RECT 1.8230 12.1365 1.8490 13.2300 ;
      RECT 1.7150 12.1365 1.7410 13.2300 ;
      RECT 1.6070 12.1365 1.6330 13.2300 ;
      RECT 1.4990 12.1365 1.5250 13.2300 ;
      RECT 1.3910 12.1365 1.4170 13.2300 ;
      RECT 1.2830 12.1365 1.3090 13.2300 ;
      RECT 1.1750 12.1365 1.2010 13.2300 ;
      RECT 1.0670 12.1365 1.0930 13.2300 ;
      RECT 0.9590 12.1365 0.9850 13.2300 ;
      RECT 0.8510 12.1365 0.8770 13.2300 ;
      RECT 0.7430 12.1365 0.7690 13.2300 ;
      RECT 0.6350 12.1365 0.6610 13.2300 ;
      RECT 0.5270 12.1365 0.5530 13.2300 ;
      RECT 0.4190 12.1365 0.4450 13.2300 ;
      RECT 0.3110 12.1365 0.3370 13.2300 ;
      RECT 0.2030 12.1365 0.2290 13.2300 ;
      RECT 0.0000 12.1365 0.0850 13.2300 ;
      RECT 5.1800 13.2165 5.3080 14.3100 ;
      RECT 5.1660 13.8820 5.3080 14.2045 ;
      RECT 5.0180 13.6090 5.0800 14.3100 ;
      RECT 5.0040 13.9185 5.0800 14.0720 ;
      RECT 5.0180 13.2165 5.0440 14.3100 ;
      RECT 5.0180 13.3375 5.0580 13.5770 ;
      RECT 5.0180 13.2165 5.0800 13.3055 ;
      RECT 4.7210 13.6670 4.9270 14.3100 ;
      RECT 4.9010 13.2165 4.9270 14.3100 ;
      RECT 4.7210 13.9440 4.9410 14.2020 ;
      RECT 4.7210 13.2165 4.8190 14.3100 ;
      RECT 4.3040 13.2165 4.3870 14.3100 ;
      RECT 4.3040 13.3050 4.4010 14.2405 ;
      RECT 9.5270 13.2165 9.6120 14.3100 ;
      RECT 9.3830 13.2165 9.4090 14.3100 ;
      RECT 9.2750 13.2165 9.3010 14.3100 ;
      RECT 9.1670 13.2165 9.1930 14.3100 ;
      RECT 9.0590 13.2165 9.0850 14.3100 ;
      RECT 8.9510 13.2165 8.9770 14.3100 ;
      RECT 8.8430 13.2165 8.8690 14.3100 ;
      RECT 8.7350 13.2165 8.7610 14.3100 ;
      RECT 8.6270 13.2165 8.6530 14.3100 ;
      RECT 8.5190 13.2165 8.5450 14.3100 ;
      RECT 8.4110 13.2165 8.4370 14.3100 ;
      RECT 8.3030 13.2165 8.3290 14.3100 ;
      RECT 8.1950 13.2165 8.2210 14.3100 ;
      RECT 8.0870 13.2165 8.1130 14.3100 ;
      RECT 7.9790 13.2165 8.0050 14.3100 ;
      RECT 7.8710 13.2165 7.8970 14.3100 ;
      RECT 7.7630 13.2165 7.7890 14.3100 ;
      RECT 7.6550 13.2165 7.6810 14.3100 ;
      RECT 7.5470 13.2165 7.5730 14.3100 ;
      RECT 7.4390 13.2165 7.4650 14.3100 ;
      RECT 7.3310 13.2165 7.3570 14.3100 ;
      RECT 7.2230 13.2165 7.2490 14.3100 ;
      RECT 7.1150 13.2165 7.1410 14.3100 ;
      RECT 7.0070 13.2165 7.0330 14.3100 ;
      RECT 6.8990 13.2165 6.9250 14.3100 ;
      RECT 6.7910 13.2165 6.8170 14.3100 ;
      RECT 6.6830 13.2165 6.7090 14.3100 ;
      RECT 6.5750 13.2165 6.6010 14.3100 ;
      RECT 6.4670 13.2165 6.4930 14.3100 ;
      RECT 6.3590 13.2165 6.3850 14.3100 ;
      RECT 6.2510 13.2165 6.2770 14.3100 ;
      RECT 6.1430 13.2165 6.1690 14.3100 ;
      RECT 6.0350 13.2165 6.0610 14.3100 ;
      RECT 5.9270 13.2165 5.9530 14.3100 ;
      RECT 5.7140 13.2165 5.7910 14.3100 ;
      RECT 3.8210 13.2165 3.8980 14.3100 ;
      RECT 3.6590 13.2165 3.6850 14.3100 ;
      RECT 3.5510 13.2165 3.5770 14.3100 ;
      RECT 3.4430 13.2165 3.4690 14.3100 ;
      RECT 3.3350 13.2165 3.3610 14.3100 ;
      RECT 3.2270 13.2165 3.2530 14.3100 ;
      RECT 3.1190 13.2165 3.1450 14.3100 ;
      RECT 3.0110 13.2165 3.0370 14.3100 ;
      RECT 2.9030 13.2165 2.9290 14.3100 ;
      RECT 2.7950 13.2165 2.8210 14.3100 ;
      RECT 2.6870 13.2165 2.7130 14.3100 ;
      RECT 2.5790 13.2165 2.6050 14.3100 ;
      RECT 2.4710 13.2165 2.4970 14.3100 ;
      RECT 2.3630 13.2165 2.3890 14.3100 ;
      RECT 2.2550 13.2165 2.2810 14.3100 ;
      RECT 2.1470 13.2165 2.1730 14.3100 ;
      RECT 2.0390 13.2165 2.0650 14.3100 ;
      RECT 1.9310 13.2165 1.9570 14.3100 ;
      RECT 1.8230 13.2165 1.8490 14.3100 ;
      RECT 1.7150 13.2165 1.7410 14.3100 ;
      RECT 1.6070 13.2165 1.6330 14.3100 ;
      RECT 1.4990 13.2165 1.5250 14.3100 ;
      RECT 1.3910 13.2165 1.4170 14.3100 ;
      RECT 1.2830 13.2165 1.3090 14.3100 ;
      RECT 1.1750 13.2165 1.2010 14.3100 ;
      RECT 1.0670 13.2165 1.0930 14.3100 ;
      RECT 0.9590 13.2165 0.9850 14.3100 ;
      RECT 0.8510 13.2165 0.8770 14.3100 ;
      RECT 0.7430 13.2165 0.7690 14.3100 ;
      RECT 0.6350 13.2165 0.6610 14.3100 ;
      RECT 0.5270 13.2165 0.5530 14.3100 ;
      RECT 0.4190 13.2165 0.4450 14.3100 ;
      RECT 0.3110 13.2165 0.3370 14.3100 ;
      RECT 0.2030 13.2165 0.2290 14.3100 ;
      RECT 0.0000 13.2165 0.0850 14.3100 ;
      RECT 5.1800 14.2965 5.3080 15.3900 ;
      RECT 5.1660 14.9620 5.3080 15.2845 ;
      RECT 5.0180 14.6890 5.0800 15.3900 ;
      RECT 5.0040 14.9985 5.0800 15.1520 ;
      RECT 5.0180 14.2965 5.0440 15.3900 ;
      RECT 5.0180 14.4175 5.0580 14.6570 ;
      RECT 5.0180 14.2965 5.0800 14.3855 ;
      RECT 4.7210 14.7470 4.9270 15.3900 ;
      RECT 4.9010 14.2965 4.9270 15.3900 ;
      RECT 4.7210 15.0240 4.9410 15.2820 ;
      RECT 4.7210 14.2965 4.8190 15.3900 ;
      RECT 4.3040 14.2965 4.3870 15.3900 ;
      RECT 4.3040 14.3850 4.4010 15.3205 ;
      RECT 9.5270 14.2965 9.6120 15.3900 ;
      RECT 9.3830 14.2965 9.4090 15.3900 ;
      RECT 9.2750 14.2965 9.3010 15.3900 ;
      RECT 9.1670 14.2965 9.1930 15.3900 ;
      RECT 9.0590 14.2965 9.0850 15.3900 ;
      RECT 8.9510 14.2965 8.9770 15.3900 ;
      RECT 8.8430 14.2965 8.8690 15.3900 ;
      RECT 8.7350 14.2965 8.7610 15.3900 ;
      RECT 8.6270 14.2965 8.6530 15.3900 ;
      RECT 8.5190 14.2965 8.5450 15.3900 ;
      RECT 8.4110 14.2965 8.4370 15.3900 ;
      RECT 8.3030 14.2965 8.3290 15.3900 ;
      RECT 8.1950 14.2965 8.2210 15.3900 ;
      RECT 8.0870 14.2965 8.1130 15.3900 ;
      RECT 7.9790 14.2965 8.0050 15.3900 ;
      RECT 7.8710 14.2965 7.8970 15.3900 ;
      RECT 7.7630 14.2965 7.7890 15.3900 ;
      RECT 7.6550 14.2965 7.6810 15.3900 ;
      RECT 7.5470 14.2965 7.5730 15.3900 ;
      RECT 7.4390 14.2965 7.4650 15.3900 ;
      RECT 7.3310 14.2965 7.3570 15.3900 ;
      RECT 7.2230 14.2965 7.2490 15.3900 ;
      RECT 7.1150 14.2965 7.1410 15.3900 ;
      RECT 7.0070 14.2965 7.0330 15.3900 ;
      RECT 6.8990 14.2965 6.9250 15.3900 ;
      RECT 6.7910 14.2965 6.8170 15.3900 ;
      RECT 6.6830 14.2965 6.7090 15.3900 ;
      RECT 6.5750 14.2965 6.6010 15.3900 ;
      RECT 6.4670 14.2965 6.4930 15.3900 ;
      RECT 6.3590 14.2965 6.3850 15.3900 ;
      RECT 6.2510 14.2965 6.2770 15.3900 ;
      RECT 6.1430 14.2965 6.1690 15.3900 ;
      RECT 6.0350 14.2965 6.0610 15.3900 ;
      RECT 5.9270 14.2965 5.9530 15.3900 ;
      RECT 5.7140 14.2965 5.7910 15.3900 ;
      RECT 3.8210 14.2965 3.8980 15.3900 ;
      RECT 3.6590 14.2965 3.6850 15.3900 ;
      RECT 3.5510 14.2965 3.5770 15.3900 ;
      RECT 3.4430 14.2965 3.4690 15.3900 ;
      RECT 3.3350 14.2965 3.3610 15.3900 ;
      RECT 3.2270 14.2965 3.2530 15.3900 ;
      RECT 3.1190 14.2965 3.1450 15.3900 ;
      RECT 3.0110 14.2965 3.0370 15.3900 ;
      RECT 2.9030 14.2965 2.9290 15.3900 ;
      RECT 2.7950 14.2965 2.8210 15.3900 ;
      RECT 2.6870 14.2965 2.7130 15.3900 ;
      RECT 2.5790 14.2965 2.6050 15.3900 ;
      RECT 2.4710 14.2965 2.4970 15.3900 ;
      RECT 2.3630 14.2965 2.3890 15.3900 ;
      RECT 2.2550 14.2965 2.2810 15.3900 ;
      RECT 2.1470 14.2965 2.1730 15.3900 ;
      RECT 2.0390 14.2965 2.0650 15.3900 ;
      RECT 1.9310 14.2965 1.9570 15.3900 ;
      RECT 1.8230 14.2965 1.8490 15.3900 ;
      RECT 1.7150 14.2965 1.7410 15.3900 ;
      RECT 1.6070 14.2965 1.6330 15.3900 ;
      RECT 1.4990 14.2965 1.5250 15.3900 ;
      RECT 1.3910 14.2965 1.4170 15.3900 ;
      RECT 1.2830 14.2965 1.3090 15.3900 ;
      RECT 1.1750 14.2965 1.2010 15.3900 ;
      RECT 1.0670 14.2965 1.0930 15.3900 ;
      RECT 0.9590 14.2965 0.9850 15.3900 ;
      RECT 0.8510 14.2965 0.8770 15.3900 ;
      RECT 0.7430 14.2965 0.7690 15.3900 ;
      RECT 0.6350 14.2965 0.6610 15.3900 ;
      RECT 0.5270 14.2965 0.5530 15.3900 ;
      RECT 0.4190 14.2965 0.4450 15.3900 ;
      RECT 0.3110 14.2965 0.3370 15.3900 ;
      RECT 0.2030 14.2965 0.2290 15.3900 ;
      RECT 0.0000 14.2965 0.0850 15.3900 ;
      RECT 5.1800 15.3765 5.3080 16.4700 ;
      RECT 5.1660 16.0420 5.3080 16.3645 ;
      RECT 5.0180 15.7690 5.0800 16.4700 ;
      RECT 5.0040 16.0785 5.0800 16.2320 ;
      RECT 5.0180 15.3765 5.0440 16.4700 ;
      RECT 5.0180 15.4975 5.0580 15.7370 ;
      RECT 5.0180 15.3765 5.0800 15.4655 ;
      RECT 4.7210 15.8270 4.9270 16.4700 ;
      RECT 4.9010 15.3765 4.9270 16.4700 ;
      RECT 4.7210 16.1040 4.9410 16.3620 ;
      RECT 4.7210 15.3765 4.8190 16.4700 ;
      RECT 4.3040 15.3765 4.3870 16.4700 ;
      RECT 4.3040 15.4650 4.4010 16.4005 ;
      RECT 9.5270 15.3765 9.6120 16.4700 ;
      RECT 9.3830 15.3765 9.4090 16.4700 ;
      RECT 9.2750 15.3765 9.3010 16.4700 ;
      RECT 9.1670 15.3765 9.1930 16.4700 ;
      RECT 9.0590 15.3765 9.0850 16.4700 ;
      RECT 8.9510 15.3765 8.9770 16.4700 ;
      RECT 8.8430 15.3765 8.8690 16.4700 ;
      RECT 8.7350 15.3765 8.7610 16.4700 ;
      RECT 8.6270 15.3765 8.6530 16.4700 ;
      RECT 8.5190 15.3765 8.5450 16.4700 ;
      RECT 8.4110 15.3765 8.4370 16.4700 ;
      RECT 8.3030 15.3765 8.3290 16.4700 ;
      RECT 8.1950 15.3765 8.2210 16.4700 ;
      RECT 8.0870 15.3765 8.1130 16.4700 ;
      RECT 7.9790 15.3765 8.0050 16.4700 ;
      RECT 7.8710 15.3765 7.8970 16.4700 ;
      RECT 7.7630 15.3765 7.7890 16.4700 ;
      RECT 7.6550 15.3765 7.6810 16.4700 ;
      RECT 7.5470 15.3765 7.5730 16.4700 ;
      RECT 7.4390 15.3765 7.4650 16.4700 ;
      RECT 7.3310 15.3765 7.3570 16.4700 ;
      RECT 7.2230 15.3765 7.2490 16.4700 ;
      RECT 7.1150 15.3765 7.1410 16.4700 ;
      RECT 7.0070 15.3765 7.0330 16.4700 ;
      RECT 6.8990 15.3765 6.9250 16.4700 ;
      RECT 6.7910 15.3765 6.8170 16.4700 ;
      RECT 6.6830 15.3765 6.7090 16.4700 ;
      RECT 6.5750 15.3765 6.6010 16.4700 ;
      RECT 6.4670 15.3765 6.4930 16.4700 ;
      RECT 6.3590 15.3765 6.3850 16.4700 ;
      RECT 6.2510 15.3765 6.2770 16.4700 ;
      RECT 6.1430 15.3765 6.1690 16.4700 ;
      RECT 6.0350 15.3765 6.0610 16.4700 ;
      RECT 5.9270 15.3765 5.9530 16.4700 ;
      RECT 5.7140 15.3765 5.7910 16.4700 ;
      RECT 3.8210 15.3765 3.8980 16.4700 ;
      RECT 3.6590 15.3765 3.6850 16.4700 ;
      RECT 3.5510 15.3765 3.5770 16.4700 ;
      RECT 3.4430 15.3765 3.4690 16.4700 ;
      RECT 3.3350 15.3765 3.3610 16.4700 ;
      RECT 3.2270 15.3765 3.2530 16.4700 ;
      RECT 3.1190 15.3765 3.1450 16.4700 ;
      RECT 3.0110 15.3765 3.0370 16.4700 ;
      RECT 2.9030 15.3765 2.9290 16.4700 ;
      RECT 2.7950 15.3765 2.8210 16.4700 ;
      RECT 2.6870 15.3765 2.7130 16.4700 ;
      RECT 2.5790 15.3765 2.6050 16.4700 ;
      RECT 2.4710 15.3765 2.4970 16.4700 ;
      RECT 2.3630 15.3765 2.3890 16.4700 ;
      RECT 2.2550 15.3765 2.2810 16.4700 ;
      RECT 2.1470 15.3765 2.1730 16.4700 ;
      RECT 2.0390 15.3765 2.0650 16.4700 ;
      RECT 1.9310 15.3765 1.9570 16.4700 ;
      RECT 1.8230 15.3765 1.8490 16.4700 ;
      RECT 1.7150 15.3765 1.7410 16.4700 ;
      RECT 1.6070 15.3765 1.6330 16.4700 ;
      RECT 1.4990 15.3765 1.5250 16.4700 ;
      RECT 1.3910 15.3765 1.4170 16.4700 ;
      RECT 1.2830 15.3765 1.3090 16.4700 ;
      RECT 1.1750 15.3765 1.2010 16.4700 ;
      RECT 1.0670 15.3765 1.0930 16.4700 ;
      RECT 0.9590 15.3765 0.9850 16.4700 ;
      RECT 0.8510 15.3765 0.8770 16.4700 ;
      RECT 0.7430 15.3765 0.7690 16.4700 ;
      RECT 0.6350 15.3765 0.6610 16.4700 ;
      RECT 0.5270 15.3765 0.5530 16.4700 ;
      RECT 0.4190 15.3765 0.4450 16.4700 ;
      RECT 0.3110 15.3765 0.3370 16.4700 ;
      RECT 0.2030 15.3765 0.2290 16.4700 ;
      RECT 0.0000 15.3765 0.0850 16.4700 ;
      RECT 5.1800 16.4565 5.3080 17.5500 ;
      RECT 5.1660 17.1220 5.3080 17.4445 ;
      RECT 5.0180 16.8490 5.0800 17.5500 ;
      RECT 5.0040 17.1585 5.0800 17.3120 ;
      RECT 5.0180 16.4565 5.0440 17.5500 ;
      RECT 5.0180 16.5775 5.0580 16.8170 ;
      RECT 5.0180 16.4565 5.0800 16.5455 ;
      RECT 4.7210 16.9070 4.9270 17.5500 ;
      RECT 4.9010 16.4565 4.9270 17.5500 ;
      RECT 4.7210 17.1840 4.9410 17.4420 ;
      RECT 4.7210 16.4565 4.8190 17.5500 ;
      RECT 4.3040 16.4565 4.3870 17.5500 ;
      RECT 4.3040 16.5450 4.4010 17.4805 ;
      RECT 9.5270 16.4565 9.6120 17.5500 ;
      RECT 9.3830 16.4565 9.4090 17.5500 ;
      RECT 9.2750 16.4565 9.3010 17.5500 ;
      RECT 9.1670 16.4565 9.1930 17.5500 ;
      RECT 9.0590 16.4565 9.0850 17.5500 ;
      RECT 8.9510 16.4565 8.9770 17.5500 ;
      RECT 8.8430 16.4565 8.8690 17.5500 ;
      RECT 8.7350 16.4565 8.7610 17.5500 ;
      RECT 8.6270 16.4565 8.6530 17.5500 ;
      RECT 8.5190 16.4565 8.5450 17.5500 ;
      RECT 8.4110 16.4565 8.4370 17.5500 ;
      RECT 8.3030 16.4565 8.3290 17.5500 ;
      RECT 8.1950 16.4565 8.2210 17.5500 ;
      RECT 8.0870 16.4565 8.1130 17.5500 ;
      RECT 7.9790 16.4565 8.0050 17.5500 ;
      RECT 7.8710 16.4565 7.8970 17.5500 ;
      RECT 7.7630 16.4565 7.7890 17.5500 ;
      RECT 7.6550 16.4565 7.6810 17.5500 ;
      RECT 7.5470 16.4565 7.5730 17.5500 ;
      RECT 7.4390 16.4565 7.4650 17.5500 ;
      RECT 7.3310 16.4565 7.3570 17.5500 ;
      RECT 7.2230 16.4565 7.2490 17.5500 ;
      RECT 7.1150 16.4565 7.1410 17.5500 ;
      RECT 7.0070 16.4565 7.0330 17.5500 ;
      RECT 6.8990 16.4565 6.9250 17.5500 ;
      RECT 6.7910 16.4565 6.8170 17.5500 ;
      RECT 6.6830 16.4565 6.7090 17.5500 ;
      RECT 6.5750 16.4565 6.6010 17.5500 ;
      RECT 6.4670 16.4565 6.4930 17.5500 ;
      RECT 6.3590 16.4565 6.3850 17.5500 ;
      RECT 6.2510 16.4565 6.2770 17.5500 ;
      RECT 6.1430 16.4565 6.1690 17.5500 ;
      RECT 6.0350 16.4565 6.0610 17.5500 ;
      RECT 5.9270 16.4565 5.9530 17.5500 ;
      RECT 5.7140 16.4565 5.7910 17.5500 ;
      RECT 3.8210 16.4565 3.8980 17.5500 ;
      RECT 3.6590 16.4565 3.6850 17.5500 ;
      RECT 3.5510 16.4565 3.5770 17.5500 ;
      RECT 3.4430 16.4565 3.4690 17.5500 ;
      RECT 3.3350 16.4565 3.3610 17.5500 ;
      RECT 3.2270 16.4565 3.2530 17.5500 ;
      RECT 3.1190 16.4565 3.1450 17.5500 ;
      RECT 3.0110 16.4565 3.0370 17.5500 ;
      RECT 2.9030 16.4565 2.9290 17.5500 ;
      RECT 2.7950 16.4565 2.8210 17.5500 ;
      RECT 2.6870 16.4565 2.7130 17.5500 ;
      RECT 2.5790 16.4565 2.6050 17.5500 ;
      RECT 2.4710 16.4565 2.4970 17.5500 ;
      RECT 2.3630 16.4565 2.3890 17.5500 ;
      RECT 2.2550 16.4565 2.2810 17.5500 ;
      RECT 2.1470 16.4565 2.1730 17.5500 ;
      RECT 2.0390 16.4565 2.0650 17.5500 ;
      RECT 1.9310 16.4565 1.9570 17.5500 ;
      RECT 1.8230 16.4565 1.8490 17.5500 ;
      RECT 1.7150 16.4565 1.7410 17.5500 ;
      RECT 1.6070 16.4565 1.6330 17.5500 ;
      RECT 1.4990 16.4565 1.5250 17.5500 ;
      RECT 1.3910 16.4565 1.4170 17.5500 ;
      RECT 1.2830 16.4565 1.3090 17.5500 ;
      RECT 1.1750 16.4565 1.2010 17.5500 ;
      RECT 1.0670 16.4565 1.0930 17.5500 ;
      RECT 0.9590 16.4565 0.9850 17.5500 ;
      RECT 0.8510 16.4565 0.8770 17.5500 ;
      RECT 0.7430 16.4565 0.7690 17.5500 ;
      RECT 0.6350 16.4565 0.6610 17.5500 ;
      RECT 0.5270 16.4565 0.5530 17.5500 ;
      RECT 0.4190 16.4565 0.4450 17.5500 ;
      RECT 0.3110 16.4565 0.3370 17.5500 ;
      RECT 0.2030 16.4565 0.2290 17.5500 ;
      RECT 0.0000 16.4565 0.0850 17.5500 ;
      RECT 0.0000 25.8840 9.6120 26.1765 ;
      RECT 9.5270 17.5230 9.6120 26.1765 ;
      RECT 4.5410 25.7355 9.6120 26.1765 ;
      RECT 0.0000 25.7355 4.3870 26.1765 ;
      RECT 5.9270 19.0270 9.4090 26.1765 ;
      RECT 7.3850 17.5230 9.4090 26.1765 ;
      RECT 4.5410 25.7090 5.8450 26.1765 ;
      RECT 5.1800 25.7080 5.8450 26.1765 ;
      RECT 3.7670 19.1350 4.3870 26.1765 ;
      RECT 3.8210 18.2890 4.3870 26.1765 ;
      RECT 0.2030 18.8320 3.6850 26.1765 ;
      RECT 3.3890 17.5230 3.6850 26.1765 ;
      RECT 0.0000 17.5230 0.0850 26.1765 ;
      RECT 4.5410 25.7060 5.0800 26.1765 ;
      RECT 5.0180 25.4350 5.0800 26.1765 ;
      RECT 5.1800 25.4350 5.7910 26.1765 ;
      RECT 4.5410 25.4350 4.9270 26.1765 ;
      RECT 5.9130 21.3160 9.4090 25.6760 ;
      RECT 0.2030 21.3160 3.6990 25.6760 ;
      RECT 5.9130 21.3160 9.4230 25.6715 ;
      RECT 0.1890 21.3160 3.6990 25.6715 ;
      RECT 5.1890 18.2890 5.7910 26.1765 ;
      RECT 4.7210 18.2080 4.8910 26.1765 ;
      RECT 4.8290 17.5230 4.8910 26.1765 ;
      RECT 4.0370 18.1070 4.4230 25.2850 ;
      RECT 3.7670 25.2430 4.4370 25.2800 ;
      RECT 5.1750 24.1690 5.7910 25.2770 ;
      RECT 4.7070 24.9790 4.8910 25.2050 ;
      RECT 4.7210 24.4030 4.9050 24.6650 ;
      RECT 3.7670 24.2050 4.4370 24.6650 ;
      RECT 4.7070 23.6650 4.8910 24.1250 ;
      RECT 5.1750 21.6310 5.7910 23.9630 ;
      RECT 3.7670 22.2790 4.4370 23.4230 ;
      RECT 4.7210 22.0090 4.9050 23.3150 ;
      RECT 4.7070 22.5850 4.9050 23.0450 ;
      RECT 4.7070 19.3450 4.8910 22.5050 ;
      RECT 4.7070 19.3450 4.9050 21.9650 ;
      RECT 3.7670 21.7390 4.4370 21.9650 ;
      RECT 5.2250 17.6995 5.8450 21.2840 ;
      RECT 5.1750 18.8050 5.8450 20.5910 ;
      RECT 3.7670 19.7770 4.4370 20.1470 ;
      RECT 4.7210 19.0750 4.9050 19.2650 ;
      RECT 3.8210 19.0390 4.4370 19.2290 ;
      RECT 4.7070 18.9310 4.8910 19.0670 ;
      RECT 4.7210 18.8050 4.9050 19.0310 ;
      RECT 6.0890 18.8350 9.4090 26.1765 ;
      RECT 7.1690 18.8320 9.4090 26.1765 ;
      RECT 5.9270 17.5230 6.0070 26.1765 ;
      RECT 3.7670 18.2080 3.9550 19.0220 ;
      RECT 5.9270 17.5230 6.2230 18.9260 ;
      RECT 5.9270 18.6400 7.0870 18.9260 ;
      RECT 7.1690 17.5230 7.3030 26.1765 ;
      RECT 2.5250 18.4510 3.3070 26.1765 ;
      RECT 0.2030 17.5230 2.4430 26.1765 ;
      RECT 5.9270 18.6400 7.3030 18.7340 ;
      RECT 6.9530 17.5230 9.4090 18.7310 ;
      RECT 3.1730 17.5230 3.6850 18.7310 ;
      RECT 4.7070 18.6610 4.9050 18.7250 ;
      RECT 4.7070 18.5350 4.8910 18.7250 ;
      RECT 6.7370 18.2560 9.4090 18.7310 ;
      RECT 5.9270 18.2890 6.6550 18.9260 ;
      RECT 4.7210 18.2650 4.9050 18.5270 ;
      RECT 0.2030 18.2560 3.0910 18.7310 ;
      RECT 2.9570 17.5230 3.0910 26.1765 ;
      RECT 6.5210 17.5230 6.8710 18.3950 ;
      RECT 5.9270 18.2080 6.4390 18.9260 ;
      RECT 6.3050 17.5230 6.4390 26.1765 ;
      RECT 2.7410 18.2080 3.0910 26.1765 ;
      RECT 0.2030 17.5230 2.6590 18.7310 ;
      RECT 4.7210 17.5230 4.7470 26.1765 ;
      RECT 3.8570 17.5230 3.9550 26.1765 ;
      RECT 2.7410 17.5230 2.8750 26.1765 ;
      RECT 6.3050 17.5230 6.8710 18.1580 ;
      RECT 5.1890 17.5230 5.7910 18.1580 ;
      RECT 3.8570 17.5230 4.3870 18.1580 ;
      RECT 2.9570 17.5230 3.6850 18.1580 ;
      RECT 6.3050 17.5230 9.4090 18.1550 ;
      RECT 0.2030 17.5230 2.8750 18.1550 ;
      RECT 5.1750 17.9950 5.8450 18.1490 ;
      RECT 3.8570 17.9950 4.4010 18.1580 ;
      RECT 5.9270 17.5230 9.4090 17.8910 ;
      RECT 4.7210 17.5230 4.8910 17.8910 ;
      RECT 3.7670 17.5230 4.3870 17.8910 ;
      RECT 0.2030 17.5230 3.6850 17.8910 ;
      RECT 4.5410 17.5230 4.8910 17.7880 ;
      RECT 5.1800 17.5230 5.7910 17.6880 ;
      RECT 4.5410 17.5230 4.9270 17.6880 ;
      RECT 5.1800 17.5230 5.8450 17.5440 ;
      RECT 6.3090 17.4965 6.3270 26.1765 ;
      RECT 6.2010 17.4965 6.2190 26.1765 ;
      RECT 2.9610 17.4965 2.9790 26.1765 ;
      RECT 2.8530 17.4965 2.8710 26.1765 ;
      RECT 5.0180 17.5230 5.0800 17.6880 ;
        RECT 5.1800 25.6635 5.3080 26.7570 ;
        RECT 5.1660 26.3290 5.3080 26.6515 ;
        RECT 5.0180 26.0560 5.0800 26.7570 ;
        RECT 5.0040 26.3655 5.0800 26.5190 ;
        RECT 5.0180 25.6635 5.0440 26.7570 ;
        RECT 5.0180 25.7845 5.0580 26.0240 ;
        RECT 5.0180 25.6635 5.0800 25.7525 ;
        RECT 4.7210 26.1140 4.9270 26.7570 ;
        RECT 4.9010 25.6635 4.9270 26.7570 ;
        RECT 4.7210 26.3910 4.9410 26.6490 ;
        RECT 4.7210 25.6635 4.8190 26.7570 ;
        RECT 4.3040 25.6635 4.3870 26.7570 ;
        RECT 4.3040 25.7520 4.4010 26.6875 ;
        RECT 9.5270 25.6635 9.6120 26.7570 ;
        RECT 9.3830 25.6635 9.4090 26.7570 ;
        RECT 9.2750 25.6635 9.3010 26.7570 ;
        RECT 9.1670 25.6635 9.1930 26.7570 ;
        RECT 9.0590 25.6635 9.0850 26.7570 ;
        RECT 8.9510 25.6635 8.9770 26.7570 ;
        RECT 8.8430 25.6635 8.8690 26.7570 ;
        RECT 8.7350 25.6635 8.7610 26.7570 ;
        RECT 8.6270 25.6635 8.6530 26.7570 ;
        RECT 8.5190 25.6635 8.5450 26.7570 ;
        RECT 8.4110 25.6635 8.4370 26.7570 ;
        RECT 8.3030 25.6635 8.3290 26.7570 ;
        RECT 8.1950 25.6635 8.2210 26.7570 ;
        RECT 8.0870 25.6635 8.1130 26.7570 ;
        RECT 7.9790 25.6635 8.0050 26.7570 ;
        RECT 7.8710 25.6635 7.8970 26.7570 ;
        RECT 7.7630 25.6635 7.7890 26.7570 ;
        RECT 7.6550 25.6635 7.6810 26.7570 ;
        RECT 7.5470 25.6635 7.5730 26.7570 ;
        RECT 7.4390 25.6635 7.4650 26.7570 ;
        RECT 7.3310 25.6635 7.3570 26.7570 ;
        RECT 7.2230 25.6635 7.2490 26.7570 ;
        RECT 7.1150 25.6635 7.1410 26.7570 ;
        RECT 7.0070 25.6635 7.0330 26.7570 ;
        RECT 6.8990 25.6635 6.9250 26.7570 ;
        RECT 6.7910 25.6635 6.8170 26.7570 ;
        RECT 6.6830 25.6635 6.7090 26.7570 ;
        RECT 6.5750 25.6635 6.6010 26.7570 ;
        RECT 6.4670 25.6635 6.4930 26.7570 ;
        RECT 6.3590 25.6635 6.3850 26.7570 ;
        RECT 6.2510 25.6635 6.2770 26.7570 ;
        RECT 6.1430 25.6635 6.1690 26.7570 ;
        RECT 6.0350 25.6635 6.0610 26.7570 ;
        RECT 5.9270 25.6635 5.9530 26.7570 ;
        RECT 5.7140 25.6635 5.7910 26.7570 ;
        RECT 3.8210 25.6635 3.8980 26.7570 ;
        RECT 3.6590 25.6635 3.6850 26.7570 ;
        RECT 3.5510 25.6635 3.5770 26.7570 ;
        RECT 3.4430 25.6635 3.4690 26.7570 ;
        RECT 3.3350 25.6635 3.3610 26.7570 ;
        RECT 3.2270 25.6635 3.2530 26.7570 ;
        RECT 3.1190 25.6635 3.1450 26.7570 ;
        RECT 3.0110 25.6635 3.0370 26.7570 ;
        RECT 2.9030 25.6635 2.9290 26.7570 ;
        RECT 2.7950 25.6635 2.8210 26.7570 ;
        RECT 2.6870 25.6635 2.7130 26.7570 ;
        RECT 2.5790 25.6635 2.6050 26.7570 ;
        RECT 2.4710 25.6635 2.4970 26.7570 ;
        RECT 2.3630 25.6635 2.3890 26.7570 ;
        RECT 2.2550 25.6635 2.2810 26.7570 ;
        RECT 2.1470 25.6635 2.1730 26.7570 ;
        RECT 2.0390 25.6635 2.0650 26.7570 ;
        RECT 1.9310 25.6635 1.9570 26.7570 ;
        RECT 1.8230 25.6635 1.8490 26.7570 ;
        RECT 1.7150 25.6635 1.7410 26.7570 ;
        RECT 1.6070 25.6635 1.6330 26.7570 ;
        RECT 1.4990 25.6635 1.5250 26.7570 ;
        RECT 1.3910 25.6635 1.4170 26.7570 ;
        RECT 1.2830 25.6635 1.3090 26.7570 ;
        RECT 1.1750 25.6635 1.2010 26.7570 ;
        RECT 1.0670 25.6635 1.0930 26.7570 ;
        RECT 0.9590 25.6635 0.9850 26.7570 ;
        RECT 0.8510 25.6635 0.8770 26.7570 ;
        RECT 0.7430 25.6635 0.7690 26.7570 ;
        RECT 0.6350 25.6635 0.6610 26.7570 ;
        RECT 0.5270 25.6635 0.5530 26.7570 ;
        RECT 0.4190 25.6635 0.4450 26.7570 ;
        RECT 0.3110 25.6635 0.3370 26.7570 ;
        RECT 0.2030 25.6635 0.2290 26.7570 ;
        RECT 0.0000 25.6635 0.0850 26.7570 ;
        RECT 5.1800 26.7435 5.3080 27.8370 ;
        RECT 5.1660 27.4090 5.3080 27.7315 ;
        RECT 5.0180 27.1360 5.0800 27.8370 ;
        RECT 5.0040 27.4455 5.0800 27.5990 ;
        RECT 5.0180 26.7435 5.0440 27.8370 ;
        RECT 5.0180 26.8645 5.0580 27.1040 ;
        RECT 5.0180 26.7435 5.0800 26.8325 ;
        RECT 4.7210 27.1940 4.9270 27.8370 ;
        RECT 4.9010 26.7435 4.9270 27.8370 ;
        RECT 4.7210 27.4710 4.9410 27.7290 ;
        RECT 4.7210 26.7435 4.8190 27.8370 ;
        RECT 4.3040 26.7435 4.3870 27.8370 ;
        RECT 4.3040 26.8320 4.4010 27.7675 ;
        RECT 9.5270 26.7435 9.6120 27.8370 ;
        RECT 9.3830 26.7435 9.4090 27.8370 ;
        RECT 9.2750 26.7435 9.3010 27.8370 ;
        RECT 9.1670 26.7435 9.1930 27.8370 ;
        RECT 9.0590 26.7435 9.0850 27.8370 ;
        RECT 8.9510 26.7435 8.9770 27.8370 ;
        RECT 8.8430 26.7435 8.8690 27.8370 ;
        RECT 8.7350 26.7435 8.7610 27.8370 ;
        RECT 8.6270 26.7435 8.6530 27.8370 ;
        RECT 8.5190 26.7435 8.5450 27.8370 ;
        RECT 8.4110 26.7435 8.4370 27.8370 ;
        RECT 8.3030 26.7435 8.3290 27.8370 ;
        RECT 8.1950 26.7435 8.2210 27.8370 ;
        RECT 8.0870 26.7435 8.1130 27.8370 ;
        RECT 7.9790 26.7435 8.0050 27.8370 ;
        RECT 7.8710 26.7435 7.8970 27.8370 ;
        RECT 7.7630 26.7435 7.7890 27.8370 ;
        RECT 7.6550 26.7435 7.6810 27.8370 ;
        RECT 7.5470 26.7435 7.5730 27.8370 ;
        RECT 7.4390 26.7435 7.4650 27.8370 ;
        RECT 7.3310 26.7435 7.3570 27.8370 ;
        RECT 7.2230 26.7435 7.2490 27.8370 ;
        RECT 7.1150 26.7435 7.1410 27.8370 ;
        RECT 7.0070 26.7435 7.0330 27.8370 ;
        RECT 6.8990 26.7435 6.9250 27.8370 ;
        RECT 6.7910 26.7435 6.8170 27.8370 ;
        RECT 6.6830 26.7435 6.7090 27.8370 ;
        RECT 6.5750 26.7435 6.6010 27.8370 ;
        RECT 6.4670 26.7435 6.4930 27.8370 ;
        RECT 6.3590 26.7435 6.3850 27.8370 ;
        RECT 6.2510 26.7435 6.2770 27.8370 ;
        RECT 6.1430 26.7435 6.1690 27.8370 ;
        RECT 6.0350 26.7435 6.0610 27.8370 ;
        RECT 5.9270 26.7435 5.9530 27.8370 ;
        RECT 5.7140 26.7435 5.7910 27.8370 ;
        RECT 3.8210 26.7435 3.8980 27.8370 ;
        RECT 3.6590 26.7435 3.6850 27.8370 ;
        RECT 3.5510 26.7435 3.5770 27.8370 ;
        RECT 3.4430 26.7435 3.4690 27.8370 ;
        RECT 3.3350 26.7435 3.3610 27.8370 ;
        RECT 3.2270 26.7435 3.2530 27.8370 ;
        RECT 3.1190 26.7435 3.1450 27.8370 ;
        RECT 3.0110 26.7435 3.0370 27.8370 ;
        RECT 2.9030 26.7435 2.9290 27.8370 ;
        RECT 2.7950 26.7435 2.8210 27.8370 ;
        RECT 2.6870 26.7435 2.7130 27.8370 ;
        RECT 2.5790 26.7435 2.6050 27.8370 ;
        RECT 2.4710 26.7435 2.4970 27.8370 ;
        RECT 2.3630 26.7435 2.3890 27.8370 ;
        RECT 2.2550 26.7435 2.2810 27.8370 ;
        RECT 2.1470 26.7435 2.1730 27.8370 ;
        RECT 2.0390 26.7435 2.0650 27.8370 ;
        RECT 1.9310 26.7435 1.9570 27.8370 ;
        RECT 1.8230 26.7435 1.8490 27.8370 ;
        RECT 1.7150 26.7435 1.7410 27.8370 ;
        RECT 1.6070 26.7435 1.6330 27.8370 ;
        RECT 1.4990 26.7435 1.5250 27.8370 ;
        RECT 1.3910 26.7435 1.4170 27.8370 ;
        RECT 1.2830 26.7435 1.3090 27.8370 ;
        RECT 1.1750 26.7435 1.2010 27.8370 ;
        RECT 1.0670 26.7435 1.0930 27.8370 ;
        RECT 0.9590 26.7435 0.9850 27.8370 ;
        RECT 0.8510 26.7435 0.8770 27.8370 ;
        RECT 0.7430 26.7435 0.7690 27.8370 ;
        RECT 0.6350 26.7435 0.6610 27.8370 ;
        RECT 0.5270 26.7435 0.5530 27.8370 ;
        RECT 0.4190 26.7435 0.4450 27.8370 ;
        RECT 0.3110 26.7435 0.3370 27.8370 ;
        RECT 0.2030 26.7435 0.2290 27.8370 ;
        RECT 0.0000 26.7435 0.0850 27.8370 ;
        RECT 5.1800 27.8235 5.3080 28.9170 ;
        RECT 5.1660 28.4890 5.3080 28.8115 ;
        RECT 5.0180 28.2160 5.0800 28.9170 ;
        RECT 5.0040 28.5255 5.0800 28.6790 ;
        RECT 5.0180 27.8235 5.0440 28.9170 ;
        RECT 5.0180 27.9445 5.0580 28.1840 ;
        RECT 5.0180 27.8235 5.0800 27.9125 ;
        RECT 4.7210 28.2740 4.9270 28.9170 ;
        RECT 4.9010 27.8235 4.9270 28.9170 ;
        RECT 4.7210 28.5510 4.9410 28.8090 ;
        RECT 4.7210 27.8235 4.8190 28.9170 ;
        RECT 4.3040 27.8235 4.3870 28.9170 ;
        RECT 4.3040 27.9120 4.4010 28.8475 ;
        RECT 9.5270 27.8235 9.6120 28.9170 ;
        RECT 9.3830 27.8235 9.4090 28.9170 ;
        RECT 9.2750 27.8235 9.3010 28.9170 ;
        RECT 9.1670 27.8235 9.1930 28.9170 ;
        RECT 9.0590 27.8235 9.0850 28.9170 ;
        RECT 8.9510 27.8235 8.9770 28.9170 ;
        RECT 8.8430 27.8235 8.8690 28.9170 ;
        RECT 8.7350 27.8235 8.7610 28.9170 ;
        RECT 8.6270 27.8235 8.6530 28.9170 ;
        RECT 8.5190 27.8235 8.5450 28.9170 ;
        RECT 8.4110 27.8235 8.4370 28.9170 ;
        RECT 8.3030 27.8235 8.3290 28.9170 ;
        RECT 8.1950 27.8235 8.2210 28.9170 ;
        RECT 8.0870 27.8235 8.1130 28.9170 ;
        RECT 7.9790 27.8235 8.0050 28.9170 ;
        RECT 7.8710 27.8235 7.8970 28.9170 ;
        RECT 7.7630 27.8235 7.7890 28.9170 ;
        RECT 7.6550 27.8235 7.6810 28.9170 ;
        RECT 7.5470 27.8235 7.5730 28.9170 ;
        RECT 7.4390 27.8235 7.4650 28.9170 ;
        RECT 7.3310 27.8235 7.3570 28.9170 ;
        RECT 7.2230 27.8235 7.2490 28.9170 ;
        RECT 7.1150 27.8235 7.1410 28.9170 ;
        RECT 7.0070 27.8235 7.0330 28.9170 ;
        RECT 6.8990 27.8235 6.9250 28.9170 ;
        RECT 6.7910 27.8235 6.8170 28.9170 ;
        RECT 6.6830 27.8235 6.7090 28.9170 ;
        RECT 6.5750 27.8235 6.6010 28.9170 ;
        RECT 6.4670 27.8235 6.4930 28.9170 ;
        RECT 6.3590 27.8235 6.3850 28.9170 ;
        RECT 6.2510 27.8235 6.2770 28.9170 ;
        RECT 6.1430 27.8235 6.1690 28.9170 ;
        RECT 6.0350 27.8235 6.0610 28.9170 ;
        RECT 5.9270 27.8235 5.9530 28.9170 ;
        RECT 5.7140 27.8235 5.7910 28.9170 ;
        RECT 3.8210 27.8235 3.8980 28.9170 ;
        RECT 3.6590 27.8235 3.6850 28.9170 ;
        RECT 3.5510 27.8235 3.5770 28.9170 ;
        RECT 3.4430 27.8235 3.4690 28.9170 ;
        RECT 3.3350 27.8235 3.3610 28.9170 ;
        RECT 3.2270 27.8235 3.2530 28.9170 ;
        RECT 3.1190 27.8235 3.1450 28.9170 ;
        RECT 3.0110 27.8235 3.0370 28.9170 ;
        RECT 2.9030 27.8235 2.9290 28.9170 ;
        RECT 2.7950 27.8235 2.8210 28.9170 ;
        RECT 2.6870 27.8235 2.7130 28.9170 ;
        RECT 2.5790 27.8235 2.6050 28.9170 ;
        RECT 2.4710 27.8235 2.4970 28.9170 ;
        RECT 2.3630 27.8235 2.3890 28.9170 ;
        RECT 2.2550 27.8235 2.2810 28.9170 ;
        RECT 2.1470 27.8235 2.1730 28.9170 ;
        RECT 2.0390 27.8235 2.0650 28.9170 ;
        RECT 1.9310 27.8235 1.9570 28.9170 ;
        RECT 1.8230 27.8235 1.8490 28.9170 ;
        RECT 1.7150 27.8235 1.7410 28.9170 ;
        RECT 1.6070 27.8235 1.6330 28.9170 ;
        RECT 1.4990 27.8235 1.5250 28.9170 ;
        RECT 1.3910 27.8235 1.4170 28.9170 ;
        RECT 1.2830 27.8235 1.3090 28.9170 ;
        RECT 1.1750 27.8235 1.2010 28.9170 ;
        RECT 1.0670 27.8235 1.0930 28.9170 ;
        RECT 0.9590 27.8235 0.9850 28.9170 ;
        RECT 0.8510 27.8235 0.8770 28.9170 ;
        RECT 0.7430 27.8235 0.7690 28.9170 ;
        RECT 0.6350 27.8235 0.6610 28.9170 ;
        RECT 0.5270 27.8235 0.5530 28.9170 ;
        RECT 0.4190 27.8235 0.4450 28.9170 ;
        RECT 0.3110 27.8235 0.3370 28.9170 ;
        RECT 0.2030 27.8235 0.2290 28.9170 ;
        RECT 0.0000 27.8235 0.0850 28.9170 ;
        RECT 5.1800 28.9035 5.3080 29.9970 ;
        RECT 5.1660 29.5690 5.3080 29.8915 ;
        RECT 5.0180 29.2960 5.0800 29.9970 ;
        RECT 5.0040 29.6055 5.0800 29.7590 ;
        RECT 5.0180 28.9035 5.0440 29.9970 ;
        RECT 5.0180 29.0245 5.0580 29.2640 ;
        RECT 5.0180 28.9035 5.0800 28.9925 ;
        RECT 4.7210 29.3540 4.9270 29.9970 ;
        RECT 4.9010 28.9035 4.9270 29.9970 ;
        RECT 4.7210 29.6310 4.9410 29.8890 ;
        RECT 4.7210 28.9035 4.8190 29.9970 ;
        RECT 4.3040 28.9035 4.3870 29.9970 ;
        RECT 4.3040 28.9920 4.4010 29.9275 ;
        RECT 9.5270 28.9035 9.6120 29.9970 ;
        RECT 9.3830 28.9035 9.4090 29.9970 ;
        RECT 9.2750 28.9035 9.3010 29.9970 ;
        RECT 9.1670 28.9035 9.1930 29.9970 ;
        RECT 9.0590 28.9035 9.0850 29.9970 ;
        RECT 8.9510 28.9035 8.9770 29.9970 ;
        RECT 8.8430 28.9035 8.8690 29.9970 ;
        RECT 8.7350 28.9035 8.7610 29.9970 ;
        RECT 8.6270 28.9035 8.6530 29.9970 ;
        RECT 8.5190 28.9035 8.5450 29.9970 ;
        RECT 8.4110 28.9035 8.4370 29.9970 ;
        RECT 8.3030 28.9035 8.3290 29.9970 ;
        RECT 8.1950 28.9035 8.2210 29.9970 ;
        RECT 8.0870 28.9035 8.1130 29.9970 ;
        RECT 7.9790 28.9035 8.0050 29.9970 ;
        RECT 7.8710 28.9035 7.8970 29.9970 ;
        RECT 7.7630 28.9035 7.7890 29.9970 ;
        RECT 7.6550 28.9035 7.6810 29.9970 ;
        RECT 7.5470 28.9035 7.5730 29.9970 ;
        RECT 7.4390 28.9035 7.4650 29.9970 ;
        RECT 7.3310 28.9035 7.3570 29.9970 ;
        RECT 7.2230 28.9035 7.2490 29.9970 ;
        RECT 7.1150 28.9035 7.1410 29.9970 ;
        RECT 7.0070 28.9035 7.0330 29.9970 ;
        RECT 6.8990 28.9035 6.9250 29.9970 ;
        RECT 6.7910 28.9035 6.8170 29.9970 ;
        RECT 6.6830 28.9035 6.7090 29.9970 ;
        RECT 6.5750 28.9035 6.6010 29.9970 ;
        RECT 6.4670 28.9035 6.4930 29.9970 ;
        RECT 6.3590 28.9035 6.3850 29.9970 ;
        RECT 6.2510 28.9035 6.2770 29.9970 ;
        RECT 6.1430 28.9035 6.1690 29.9970 ;
        RECT 6.0350 28.9035 6.0610 29.9970 ;
        RECT 5.9270 28.9035 5.9530 29.9970 ;
        RECT 5.7140 28.9035 5.7910 29.9970 ;
        RECT 3.8210 28.9035 3.8980 29.9970 ;
        RECT 3.6590 28.9035 3.6850 29.9970 ;
        RECT 3.5510 28.9035 3.5770 29.9970 ;
        RECT 3.4430 28.9035 3.4690 29.9970 ;
        RECT 3.3350 28.9035 3.3610 29.9970 ;
        RECT 3.2270 28.9035 3.2530 29.9970 ;
        RECT 3.1190 28.9035 3.1450 29.9970 ;
        RECT 3.0110 28.9035 3.0370 29.9970 ;
        RECT 2.9030 28.9035 2.9290 29.9970 ;
        RECT 2.7950 28.9035 2.8210 29.9970 ;
        RECT 2.6870 28.9035 2.7130 29.9970 ;
        RECT 2.5790 28.9035 2.6050 29.9970 ;
        RECT 2.4710 28.9035 2.4970 29.9970 ;
        RECT 2.3630 28.9035 2.3890 29.9970 ;
        RECT 2.2550 28.9035 2.2810 29.9970 ;
        RECT 2.1470 28.9035 2.1730 29.9970 ;
        RECT 2.0390 28.9035 2.0650 29.9970 ;
        RECT 1.9310 28.9035 1.9570 29.9970 ;
        RECT 1.8230 28.9035 1.8490 29.9970 ;
        RECT 1.7150 28.9035 1.7410 29.9970 ;
        RECT 1.6070 28.9035 1.6330 29.9970 ;
        RECT 1.4990 28.9035 1.5250 29.9970 ;
        RECT 1.3910 28.9035 1.4170 29.9970 ;
        RECT 1.2830 28.9035 1.3090 29.9970 ;
        RECT 1.1750 28.9035 1.2010 29.9970 ;
        RECT 1.0670 28.9035 1.0930 29.9970 ;
        RECT 0.9590 28.9035 0.9850 29.9970 ;
        RECT 0.8510 28.9035 0.8770 29.9970 ;
        RECT 0.7430 28.9035 0.7690 29.9970 ;
        RECT 0.6350 28.9035 0.6610 29.9970 ;
        RECT 0.5270 28.9035 0.5530 29.9970 ;
        RECT 0.4190 28.9035 0.4450 29.9970 ;
        RECT 0.3110 28.9035 0.3370 29.9970 ;
        RECT 0.2030 28.9035 0.2290 29.9970 ;
        RECT 0.0000 28.9035 0.0850 29.9970 ;
        RECT 5.1800 29.9835 5.3080 31.0770 ;
        RECT 5.1660 30.6490 5.3080 30.9715 ;
        RECT 5.0180 30.3760 5.0800 31.0770 ;
        RECT 5.0040 30.6855 5.0800 30.8390 ;
        RECT 5.0180 29.9835 5.0440 31.0770 ;
        RECT 5.0180 30.1045 5.0580 30.3440 ;
        RECT 5.0180 29.9835 5.0800 30.0725 ;
        RECT 4.7210 30.4340 4.9270 31.0770 ;
        RECT 4.9010 29.9835 4.9270 31.0770 ;
        RECT 4.7210 30.7110 4.9410 30.9690 ;
        RECT 4.7210 29.9835 4.8190 31.0770 ;
        RECT 4.3040 29.9835 4.3870 31.0770 ;
        RECT 4.3040 30.0720 4.4010 31.0075 ;
        RECT 9.5270 29.9835 9.6120 31.0770 ;
        RECT 9.3830 29.9835 9.4090 31.0770 ;
        RECT 9.2750 29.9835 9.3010 31.0770 ;
        RECT 9.1670 29.9835 9.1930 31.0770 ;
        RECT 9.0590 29.9835 9.0850 31.0770 ;
        RECT 8.9510 29.9835 8.9770 31.0770 ;
        RECT 8.8430 29.9835 8.8690 31.0770 ;
        RECT 8.7350 29.9835 8.7610 31.0770 ;
        RECT 8.6270 29.9835 8.6530 31.0770 ;
        RECT 8.5190 29.9835 8.5450 31.0770 ;
        RECT 8.4110 29.9835 8.4370 31.0770 ;
        RECT 8.3030 29.9835 8.3290 31.0770 ;
        RECT 8.1950 29.9835 8.2210 31.0770 ;
        RECT 8.0870 29.9835 8.1130 31.0770 ;
        RECT 7.9790 29.9835 8.0050 31.0770 ;
        RECT 7.8710 29.9835 7.8970 31.0770 ;
        RECT 7.7630 29.9835 7.7890 31.0770 ;
        RECT 7.6550 29.9835 7.6810 31.0770 ;
        RECT 7.5470 29.9835 7.5730 31.0770 ;
        RECT 7.4390 29.9835 7.4650 31.0770 ;
        RECT 7.3310 29.9835 7.3570 31.0770 ;
        RECT 7.2230 29.9835 7.2490 31.0770 ;
        RECT 7.1150 29.9835 7.1410 31.0770 ;
        RECT 7.0070 29.9835 7.0330 31.0770 ;
        RECT 6.8990 29.9835 6.9250 31.0770 ;
        RECT 6.7910 29.9835 6.8170 31.0770 ;
        RECT 6.6830 29.9835 6.7090 31.0770 ;
        RECT 6.5750 29.9835 6.6010 31.0770 ;
        RECT 6.4670 29.9835 6.4930 31.0770 ;
        RECT 6.3590 29.9835 6.3850 31.0770 ;
        RECT 6.2510 29.9835 6.2770 31.0770 ;
        RECT 6.1430 29.9835 6.1690 31.0770 ;
        RECT 6.0350 29.9835 6.0610 31.0770 ;
        RECT 5.9270 29.9835 5.9530 31.0770 ;
        RECT 5.7140 29.9835 5.7910 31.0770 ;
        RECT 3.8210 29.9835 3.8980 31.0770 ;
        RECT 3.6590 29.9835 3.6850 31.0770 ;
        RECT 3.5510 29.9835 3.5770 31.0770 ;
        RECT 3.4430 29.9835 3.4690 31.0770 ;
        RECT 3.3350 29.9835 3.3610 31.0770 ;
        RECT 3.2270 29.9835 3.2530 31.0770 ;
        RECT 3.1190 29.9835 3.1450 31.0770 ;
        RECT 3.0110 29.9835 3.0370 31.0770 ;
        RECT 2.9030 29.9835 2.9290 31.0770 ;
        RECT 2.7950 29.9835 2.8210 31.0770 ;
        RECT 2.6870 29.9835 2.7130 31.0770 ;
        RECT 2.5790 29.9835 2.6050 31.0770 ;
        RECT 2.4710 29.9835 2.4970 31.0770 ;
        RECT 2.3630 29.9835 2.3890 31.0770 ;
        RECT 2.2550 29.9835 2.2810 31.0770 ;
        RECT 2.1470 29.9835 2.1730 31.0770 ;
        RECT 2.0390 29.9835 2.0650 31.0770 ;
        RECT 1.9310 29.9835 1.9570 31.0770 ;
        RECT 1.8230 29.9835 1.8490 31.0770 ;
        RECT 1.7150 29.9835 1.7410 31.0770 ;
        RECT 1.6070 29.9835 1.6330 31.0770 ;
        RECT 1.4990 29.9835 1.5250 31.0770 ;
        RECT 1.3910 29.9835 1.4170 31.0770 ;
        RECT 1.2830 29.9835 1.3090 31.0770 ;
        RECT 1.1750 29.9835 1.2010 31.0770 ;
        RECT 1.0670 29.9835 1.0930 31.0770 ;
        RECT 0.9590 29.9835 0.9850 31.0770 ;
        RECT 0.8510 29.9835 0.8770 31.0770 ;
        RECT 0.7430 29.9835 0.7690 31.0770 ;
        RECT 0.6350 29.9835 0.6610 31.0770 ;
        RECT 0.5270 29.9835 0.5530 31.0770 ;
        RECT 0.4190 29.9835 0.4450 31.0770 ;
        RECT 0.3110 29.9835 0.3370 31.0770 ;
        RECT 0.2030 29.9835 0.2290 31.0770 ;
        RECT 0.0000 29.9835 0.0850 31.0770 ;
        RECT 5.1800 31.0635 5.3080 32.1570 ;
        RECT 5.1660 31.7290 5.3080 32.0515 ;
        RECT 5.0180 31.4560 5.0800 32.1570 ;
        RECT 5.0040 31.7655 5.0800 31.9190 ;
        RECT 5.0180 31.0635 5.0440 32.1570 ;
        RECT 5.0180 31.1845 5.0580 31.4240 ;
        RECT 5.0180 31.0635 5.0800 31.1525 ;
        RECT 4.7210 31.5140 4.9270 32.1570 ;
        RECT 4.9010 31.0635 4.9270 32.1570 ;
        RECT 4.7210 31.7910 4.9410 32.0490 ;
        RECT 4.7210 31.0635 4.8190 32.1570 ;
        RECT 4.3040 31.0635 4.3870 32.1570 ;
        RECT 4.3040 31.1520 4.4010 32.0875 ;
        RECT 9.5270 31.0635 9.6120 32.1570 ;
        RECT 9.3830 31.0635 9.4090 32.1570 ;
        RECT 9.2750 31.0635 9.3010 32.1570 ;
        RECT 9.1670 31.0635 9.1930 32.1570 ;
        RECT 9.0590 31.0635 9.0850 32.1570 ;
        RECT 8.9510 31.0635 8.9770 32.1570 ;
        RECT 8.8430 31.0635 8.8690 32.1570 ;
        RECT 8.7350 31.0635 8.7610 32.1570 ;
        RECT 8.6270 31.0635 8.6530 32.1570 ;
        RECT 8.5190 31.0635 8.5450 32.1570 ;
        RECT 8.4110 31.0635 8.4370 32.1570 ;
        RECT 8.3030 31.0635 8.3290 32.1570 ;
        RECT 8.1950 31.0635 8.2210 32.1570 ;
        RECT 8.0870 31.0635 8.1130 32.1570 ;
        RECT 7.9790 31.0635 8.0050 32.1570 ;
        RECT 7.8710 31.0635 7.8970 32.1570 ;
        RECT 7.7630 31.0635 7.7890 32.1570 ;
        RECT 7.6550 31.0635 7.6810 32.1570 ;
        RECT 7.5470 31.0635 7.5730 32.1570 ;
        RECT 7.4390 31.0635 7.4650 32.1570 ;
        RECT 7.3310 31.0635 7.3570 32.1570 ;
        RECT 7.2230 31.0635 7.2490 32.1570 ;
        RECT 7.1150 31.0635 7.1410 32.1570 ;
        RECT 7.0070 31.0635 7.0330 32.1570 ;
        RECT 6.8990 31.0635 6.9250 32.1570 ;
        RECT 6.7910 31.0635 6.8170 32.1570 ;
        RECT 6.6830 31.0635 6.7090 32.1570 ;
        RECT 6.5750 31.0635 6.6010 32.1570 ;
        RECT 6.4670 31.0635 6.4930 32.1570 ;
        RECT 6.3590 31.0635 6.3850 32.1570 ;
        RECT 6.2510 31.0635 6.2770 32.1570 ;
        RECT 6.1430 31.0635 6.1690 32.1570 ;
        RECT 6.0350 31.0635 6.0610 32.1570 ;
        RECT 5.9270 31.0635 5.9530 32.1570 ;
        RECT 5.7140 31.0635 5.7910 32.1570 ;
        RECT 3.8210 31.0635 3.8980 32.1570 ;
        RECT 3.6590 31.0635 3.6850 32.1570 ;
        RECT 3.5510 31.0635 3.5770 32.1570 ;
        RECT 3.4430 31.0635 3.4690 32.1570 ;
        RECT 3.3350 31.0635 3.3610 32.1570 ;
        RECT 3.2270 31.0635 3.2530 32.1570 ;
        RECT 3.1190 31.0635 3.1450 32.1570 ;
        RECT 3.0110 31.0635 3.0370 32.1570 ;
        RECT 2.9030 31.0635 2.9290 32.1570 ;
        RECT 2.7950 31.0635 2.8210 32.1570 ;
        RECT 2.6870 31.0635 2.7130 32.1570 ;
        RECT 2.5790 31.0635 2.6050 32.1570 ;
        RECT 2.4710 31.0635 2.4970 32.1570 ;
        RECT 2.3630 31.0635 2.3890 32.1570 ;
        RECT 2.2550 31.0635 2.2810 32.1570 ;
        RECT 2.1470 31.0635 2.1730 32.1570 ;
        RECT 2.0390 31.0635 2.0650 32.1570 ;
        RECT 1.9310 31.0635 1.9570 32.1570 ;
        RECT 1.8230 31.0635 1.8490 32.1570 ;
        RECT 1.7150 31.0635 1.7410 32.1570 ;
        RECT 1.6070 31.0635 1.6330 32.1570 ;
        RECT 1.4990 31.0635 1.5250 32.1570 ;
        RECT 1.3910 31.0635 1.4170 32.1570 ;
        RECT 1.2830 31.0635 1.3090 32.1570 ;
        RECT 1.1750 31.0635 1.2010 32.1570 ;
        RECT 1.0670 31.0635 1.0930 32.1570 ;
        RECT 0.9590 31.0635 0.9850 32.1570 ;
        RECT 0.8510 31.0635 0.8770 32.1570 ;
        RECT 0.7430 31.0635 0.7690 32.1570 ;
        RECT 0.6350 31.0635 0.6610 32.1570 ;
        RECT 0.5270 31.0635 0.5530 32.1570 ;
        RECT 0.4190 31.0635 0.4450 32.1570 ;
        RECT 0.3110 31.0635 0.3370 32.1570 ;
        RECT 0.2030 31.0635 0.2290 32.1570 ;
        RECT 0.0000 31.0635 0.0850 32.1570 ;
        RECT 5.1800 32.1435 5.3080 33.2370 ;
        RECT 5.1660 32.8090 5.3080 33.1315 ;
        RECT 5.0180 32.5360 5.0800 33.2370 ;
        RECT 5.0040 32.8455 5.0800 32.9990 ;
        RECT 5.0180 32.1435 5.0440 33.2370 ;
        RECT 5.0180 32.2645 5.0580 32.5040 ;
        RECT 5.0180 32.1435 5.0800 32.2325 ;
        RECT 4.7210 32.5940 4.9270 33.2370 ;
        RECT 4.9010 32.1435 4.9270 33.2370 ;
        RECT 4.7210 32.8710 4.9410 33.1290 ;
        RECT 4.7210 32.1435 4.8190 33.2370 ;
        RECT 4.3040 32.1435 4.3870 33.2370 ;
        RECT 4.3040 32.2320 4.4010 33.1675 ;
        RECT 9.5270 32.1435 9.6120 33.2370 ;
        RECT 9.3830 32.1435 9.4090 33.2370 ;
        RECT 9.2750 32.1435 9.3010 33.2370 ;
        RECT 9.1670 32.1435 9.1930 33.2370 ;
        RECT 9.0590 32.1435 9.0850 33.2370 ;
        RECT 8.9510 32.1435 8.9770 33.2370 ;
        RECT 8.8430 32.1435 8.8690 33.2370 ;
        RECT 8.7350 32.1435 8.7610 33.2370 ;
        RECT 8.6270 32.1435 8.6530 33.2370 ;
        RECT 8.5190 32.1435 8.5450 33.2370 ;
        RECT 8.4110 32.1435 8.4370 33.2370 ;
        RECT 8.3030 32.1435 8.3290 33.2370 ;
        RECT 8.1950 32.1435 8.2210 33.2370 ;
        RECT 8.0870 32.1435 8.1130 33.2370 ;
        RECT 7.9790 32.1435 8.0050 33.2370 ;
        RECT 7.8710 32.1435 7.8970 33.2370 ;
        RECT 7.7630 32.1435 7.7890 33.2370 ;
        RECT 7.6550 32.1435 7.6810 33.2370 ;
        RECT 7.5470 32.1435 7.5730 33.2370 ;
        RECT 7.4390 32.1435 7.4650 33.2370 ;
        RECT 7.3310 32.1435 7.3570 33.2370 ;
        RECT 7.2230 32.1435 7.2490 33.2370 ;
        RECT 7.1150 32.1435 7.1410 33.2370 ;
        RECT 7.0070 32.1435 7.0330 33.2370 ;
        RECT 6.8990 32.1435 6.9250 33.2370 ;
        RECT 6.7910 32.1435 6.8170 33.2370 ;
        RECT 6.6830 32.1435 6.7090 33.2370 ;
        RECT 6.5750 32.1435 6.6010 33.2370 ;
        RECT 6.4670 32.1435 6.4930 33.2370 ;
        RECT 6.3590 32.1435 6.3850 33.2370 ;
        RECT 6.2510 32.1435 6.2770 33.2370 ;
        RECT 6.1430 32.1435 6.1690 33.2370 ;
        RECT 6.0350 32.1435 6.0610 33.2370 ;
        RECT 5.9270 32.1435 5.9530 33.2370 ;
        RECT 5.7140 32.1435 5.7910 33.2370 ;
        RECT 3.8210 32.1435 3.8980 33.2370 ;
        RECT 3.6590 32.1435 3.6850 33.2370 ;
        RECT 3.5510 32.1435 3.5770 33.2370 ;
        RECT 3.4430 32.1435 3.4690 33.2370 ;
        RECT 3.3350 32.1435 3.3610 33.2370 ;
        RECT 3.2270 32.1435 3.2530 33.2370 ;
        RECT 3.1190 32.1435 3.1450 33.2370 ;
        RECT 3.0110 32.1435 3.0370 33.2370 ;
        RECT 2.9030 32.1435 2.9290 33.2370 ;
        RECT 2.7950 32.1435 2.8210 33.2370 ;
        RECT 2.6870 32.1435 2.7130 33.2370 ;
        RECT 2.5790 32.1435 2.6050 33.2370 ;
        RECT 2.4710 32.1435 2.4970 33.2370 ;
        RECT 2.3630 32.1435 2.3890 33.2370 ;
        RECT 2.2550 32.1435 2.2810 33.2370 ;
        RECT 2.1470 32.1435 2.1730 33.2370 ;
        RECT 2.0390 32.1435 2.0650 33.2370 ;
        RECT 1.9310 32.1435 1.9570 33.2370 ;
        RECT 1.8230 32.1435 1.8490 33.2370 ;
        RECT 1.7150 32.1435 1.7410 33.2370 ;
        RECT 1.6070 32.1435 1.6330 33.2370 ;
        RECT 1.4990 32.1435 1.5250 33.2370 ;
        RECT 1.3910 32.1435 1.4170 33.2370 ;
        RECT 1.2830 32.1435 1.3090 33.2370 ;
        RECT 1.1750 32.1435 1.2010 33.2370 ;
        RECT 1.0670 32.1435 1.0930 33.2370 ;
        RECT 0.9590 32.1435 0.9850 33.2370 ;
        RECT 0.8510 32.1435 0.8770 33.2370 ;
        RECT 0.7430 32.1435 0.7690 33.2370 ;
        RECT 0.6350 32.1435 0.6610 33.2370 ;
        RECT 0.5270 32.1435 0.5530 33.2370 ;
        RECT 0.4190 32.1435 0.4450 33.2370 ;
        RECT 0.3110 32.1435 0.3370 33.2370 ;
        RECT 0.2030 32.1435 0.2290 33.2370 ;
        RECT 0.0000 32.1435 0.0850 33.2370 ;
        RECT 5.1800 33.2235 5.3080 34.3170 ;
        RECT 5.1660 33.8890 5.3080 34.2115 ;
        RECT 5.0180 33.6160 5.0800 34.3170 ;
        RECT 5.0040 33.9255 5.0800 34.0790 ;
        RECT 5.0180 33.2235 5.0440 34.3170 ;
        RECT 5.0180 33.3445 5.0580 33.5840 ;
        RECT 5.0180 33.2235 5.0800 33.3125 ;
        RECT 4.7210 33.6740 4.9270 34.3170 ;
        RECT 4.9010 33.2235 4.9270 34.3170 ;
        RECT 4.7210 33.9510 4.9410 34.2090 ;
        RECT 4.7210 33.2235 4.8190 34.3170 ;
        RECT 4.3040 33.2235 4.3870 34.3170 ;
        RECT 4.3040 33.3120 4.4010 34.2475 ;
        RECT 9.5270 33.2235 9.6120 34.3170 ;
        RECT 9.3830 33.2235 9.4090 34.3170 ;
        RECT 9.2750 33.2235 9.3010 34.3170 ;
        RECT 9.1670 33.2235 9.1930 34.3170 ;
        RECT 9.0590 33.2235 9.0850 34.3170 ;
        RECT 8.9510 33.2235 8.9770 34.3170 ;
        RECT 8.8430 33.2235 8.8690 34.3170 ;
        RECT 8.7350 33.2235 8.7610 34.3170 ;
        RECT 8.6270 33.2235 8.6530 34.3170 ;
        RECT 8.5190 33.2235 8.5450 34.3170 ;
        RECT 8.4110 33.2235 8.4370 34.3170 ;
        RECT 8.3030 33.2235 8.3290 34.3170 ;
        RECT 8.1950 33.2235 8.2210 34.3170 ;
        RECT 8.0870 33.2235 8.1130 34.3170 ;
        RECT 7.9790 33.2235 8.0050 34.3170 ;
        RECT 7.8710 33.2235 7.8970 34.3170 ;
        RECT 7.7630 33.2235 7.7890 34.3170 ;
        RECT 7.6550 33.2235 7.6810 34.3170 ;
        RECT 7.5470 33.2235 7.5730 34.3170 ;
        RECT 7.4390 33.2235 7.4650 34.3170 ;
        RECT 7.3310 33.2235 7.3570 34.3170 ;
        RECT 7.2230 33.2235 7.2490 34.3170 ;
        RECT 7.1150 33.2235 7.1410 34.3170 ;
        RECT 7.0070 33.2235 7.0330 34.3170 ;
        RECT 6.8990 33.2235 6.9250 34.3170 ;
        RECT 6.7910 33.2235 6.8170 34.3170 ;
        RECT 6.6830 33.2235 6.7090 34.3170 ;
        RECT 6.5750 33.2235 6.6010 34.3170 ;
        RECT 6.4670 33.2235 6.4930 34.3170 ;
        RECT 6.3590 33.2235 6.3850 34.3170 ;
        RECT 6.2510 33.2235 6.2770 34.3170 ;
        RECT 6.1430 33.2235 6.1690 34.3170 ;
        RECT 6.0350 33.2235 6.0610 34.3170 ;
        RECT 5.9270 33.2235 5.9530 34.3170 ;
        RECT 5.7140 33.2235 5.7910 34.3170 ;
        RECT 3.8210 33.2235 3.8980 34.3170 ;
        RECT 3.6590 33.2235 3.6850 34.3170 ;
        RECT 3.5510 33.2235 3.5770 34.3170 ;
        RECT 3.4430 33.2235 3.4690 34.3170 ;
        RECT 3.3350 33.2235 3.3610 34.3170 ;
        RECT 3.2270 33.2235 3.2530 34.3170 ;
        RECT 3.1190 33.2235 3.1450 34.3170 ;
        RECT 3.0110 33.2235 3.0370 34.3170 ;
        RECT 2.9030 33.2235 2.9290 34.3170 ;
        RECT 2.7950 33.2235 2.8210 34.3170 ;
        RECT 2.6870 33.2235 2.7130 34.3170 ;
        RECT 2.5790 33.2235 2.6050 34.3170 ;
        RECT 2.4710 33.2235 2.4970 34.3170 ;
        RECT 2.3630 33.2235 2.3890 34.3170 ;
        RECT 2.2550 33.2235 2.2810 34.3170 ;
        RECT 2.1470 33.2235 2.1730 34.3170 ;
        RECT 2.0390 33.2235 2.0650 34.3170 ;
        RECT 1.9310 33.2235 1.9570 34.3170 ;
        RECT 1.8230 33.2235 1.8490 34.3170 ;
        RECT 1.7150 33.2235 1.7410 34.3170 ;
        RECT 1.6070 33.2235 1.6330 34.3170 ;
        RECT 1.4990 33.2235 1.5250 34.3170 ;
        RECT 1.3910 33.2235 1.4170 34.3170 ;
        RECT 1.2830 33.2235 1.3090 34.3170 ;
        RECT 1.1750 33.2235 1.2010 34.3170 ;
        RECT 1.0670 33.2235 1.0930 34.3170 ;
        RECT 0.9590 33.2235 0.9850 34.3170 ;
        RECT 0.8510 33.2235 0.8770 34.3170 ;
        RECT 0.7430 33.2235 0.7690 34.3170 ;
        RECT 0.6350 33.2235 0.6610 34.3170 ;
        RECT 0.5270 33.2235 0.5530 34.3170 ;
        RECT 0.4190 33.2235 0.4450 34.3170 ;
        RECT 0.3110 33.2235 0.3370 34.3170 ;
        RECT 0.2030 33.2235 0.2290 34.3170 ;
        RECT 0.0000 33.2235 0.0850 34.3170 ;
        RECT 5.1800 34.3035 5.3080 35.3970 ;
        RECT 5.1660 34.9690 5.3080 35.2915 ;
        RECT 5.0180 34.6960 5.0800 35.3970 ;
        RECT 5.0040 35.0055 5.0800 35.1590 ;
        RECT 5.0180 34.3035 5.0440 35.3970 ;
        RECT 5.0180 34.4245 5.0580 34.6640 ;
        RECT 5.0180 34.3035 5.0800 34.3925 ;
        RECT 4.7210 34.7540 4.9270 35.3970 ;
        RECT 4.9010 34.3035 4.9270 35.3970 ;
        RECT 4.7210 35.0310 4.9410 35.2890 ;
        RECT 4.7210 34.3035 4.8190 35.3970 ;
        RECT 4.3040 34.3035 4.3870 35.3970 ;
        RECT 4.3040 34.3920 4.4010 35.3275 ;
        RECT 9.5270 34.3035 9.6120 35.3970 ;
        RECT 9.3830 34.3035 9.4090 35.3970 ;
        RECT 9.2750 34.3035 9.3010 35.3970 ;
        RECT 9.1670 34.3035 9.1930 35.3970 ;
        RECT 9.0590 34.3035 9.0850 35.3970 ;
        RECT 8.9510 34.3035 8.9770 35.3970 ;
        RECT 8.8430 34.3035 8.8690 35.3970 ;
        RECT 8.7350 34.3035 8.7610 35.3970 ;
        RECT 8.6270 34.3035 8.6530 35.3970 ;
        RECT 8.5190 34.3035 8.5450 35.3970 ;
        RECT 8.4110 34.3035 8.4370 35.3970 ;
        RECT 8.3030 34.3035 8.3290 35.3970 ;
        RECT 8.1950 34.3035 8.2210 35.3970 ;
        RECT 8.0870 34.3035 8.1130 35.3970 ;
        RECT 7.9790 34.3035 8.0050 35.3970 ;
        RECT 7.8710 34.3035 7.8970 35.3970 ;
        RECT 7.7630 34.3035 7.7890 35.3970 ;
        RECT 7.6550 34.3035 7.6810 35.3970 ;
        RECT 7.5470 34.3035 7.5730 35.3970 ;
        RECT 7.4390 34.3035 7.4650 35.3970 ;
        RECT 7.3310 34.3035 7.3570 35.3970 ;
        RECT 7.2230 34.3035 7.2490 35.3970 ;
        RECT 7.1150 34.3035 7.1410 35.3970 ;
        RECT 7.0070 34.3035 7.0330 35.3970 ;
        RECT 6.8990 34.3035 6.9250 35.3970 ;
        RECT 6.7910 34.3035 6.8170 35.3970 ;
        RECT 6.6830 34.3035 6.7090 35.3970 ;
        RECT 6.5750 34.3035 6.6010 35.3970 ;
        RECT 6.4670 34.3035 6.4930 35.3970 ;
        RECT 6.3590 34.3035 6.3850 35.3970 ;
        RECT 6.2510 34.3035 6.2770 35.3970 ;
        RECT 6.1430 34.3035 6.1690 35.3970 ;
        RECT 6.0350 34.3035 6.0610 35.3970 ;
        RECT 5.9270 34.3035 5.9530 35.3970 ;
        RECT 5.7140 34.3035 5.7910 35.3970 ;
        RECT 3.8210 34.3035 3.8980 35.3970 ;
        RECT 3.6590 34.3035 3.6850 35.3970 ;
        RECT 3.5510 34.3035 3.5770 35.3970 ;
        RECT 3.4430 34.3035 3.4690 35.3970 ;
        RECT 3.3350 34.3035 3.3610 35.3970 ;
        RECT 3.2270 34.3035 3.2530 35.3970 ;
        RECT 3.1190 34.3035 3.1450 35.3970 ;
        RECT 3.0110 34.3035 3.0370 35.3970 ;
        RECT 2.9030 34.3035 2.9290 35.3970 ;
        RECT 2.7950 34.3035 2.8210 35.3970 ;
        RECT 2.6870 34.3035 2.7130 35.3970 ;
        RECT 2.5790 34.3035 2.6050 35.3970 ;
        RECT 2.4710 34.3035 2.4970 35.3970 ;
        RECT 2.3630 34.3035 2.3890 35.3970 ;
        RECT 2.2550 34.3035 2.2810 35.3970 ;
        RECT 2.1470 34.3035 2.1730 35.3970 ;
        RECT 2.0390 34.3035 2.0650 35.3970 ;
        RECT 1.9310 34.3035 1.9570 35.3970 ;
        RECT 1.8230 34.3035 1.8490 35.3970 ;
        RECT 1.7150 34.3035 1.7410 35.3970 ;
        RECT 1.6070 34.3035 1.6330 35.3970 ;
        RECT 1.4990 34.3035 1.5250 35.3970 ;
        RECT 1.3910 34.3035 1.4170 35.3970 ;
        RECT 1.2830 34.3035 1.3090 35.3970 ;
        RECT 1.1750 34.3035 1.2010 35.3970 ;
        RECT 1.0670 34.3035 1.0930 35.3970 ;
        RECT 0.9590 34.3035 0.9850 35.3970 ;
        RECT 0.8510 34.3035 0.8770 35.3970 ;
        RECT 0.7430 34.3035 0.7690 35.3970 ;
        RECT 0.6350 34.3035 0.6610 35.3970 ;
        RECT 0.5270 34.3035 0.5530 35.3970 ;
        RECT 0.4190 34.3035 0.4450 35.3970 ;
        RECT 0.3110 34.3035 0.3370 35.3970 ;
        RECT 0.2030 34.3035 0.2290 35.3970 ;
        RECT 0.0000 34.3035 0.0850 35.3970 ;
        RECT 5.1800 35.3835 5.3080 36.4770 ;
        RECT 5.1660 36.0490 5.3080 36.3715 ;
        RECT 5.0180 35.7760 5.0800 36.4770 ;
        RECT 5.0040 36.0855 5.0800 36.2390 ;
        RECT 5.0180 35.3835 5.0440 36.4770 ;
        RECT 5.0180 35.5045 5.0580 35.7440 ;
        RECT 5.0180 35.3835 5.0800 35.4725 ;
        RECT 4.7210 35.8340 4.9270 36.4770 ;
        RECT 4.9010 35.3835 4.9270 36.4770 ;
        RECT 4.7210 36.1110 4.9410 36.3690 ;
        RECT 4.7210 35.3835 4.8190 36.4770 ;
        RECT 4.3040 35.3835 4.3870 36.4770 ;
        RECT 4.3040 35.4720 4.4010 36.4075 ;
        RECT 9.5270 35.3835 9.6120 36.4770 ;
        RECT 9.3830 35.3835 9.4090 36.4770 ;
        RECT 9.2750 35.3835 9.3010 36.4770 ;
        RECT 9.1670 35.3835 9.1930 36.4770 ;
        RECT 9.0590 35.3835 9.0850 36.4770 ;
        RECT 8.9510 35.3835 8.9770 36.4770 ;
        RECT 8.8430 35.3835 8.8690 36.4770 ;
        RECT 8.7350 35.3835 8.7610 36.4770 ;
        RECT 8.6270 35.3835 8.6530 36.4770 ;
        RECT 8.5190 35.3835 8.5450 36.4770 ;
        RECT 8.4110 35.3835 8.4370 36.4770 ;
        RECT 8.3030 35.3835 8.3290 36.4770 ;
        RECT 8.1950 35.3835 8.2210 36.4770 ;
        RECT 8.0870 35.3835 8.1130 36.4770 ;
        RECT 7.9790 35.3835 8.0050 36.4770 ;
        RECT 7.8710 35.3835 7.8970 36.4770 ;
        RECT 7.7630 35.3835 7.7890 36.4770 ;
        RECT 7.6550 35.3835 7.6810 36.4770 ;
        RECT 7.5470 35.3835 7.5730 36.4770 ;
        RECT 7.4390 35.3835 7.4650 36.4770 ;
        RECT 7.3310 35.3835 7.3570 36.4770 ;
        RECT 7.2230 35.3835 7.2490 36.4770 ;
        RECT 7.1150 35.3835 7.1410 36.4770 ;
        RECT 7.0070 35.3835 7.0330 36.4770 ;
        RECT 6.8990 35.3835 6.9250 36.4770 ;
        RECT 6.7910 35.3835 6.8170 36.4770 ;
        RECT 6.6830 35.3835 6.7090 36.4770 ;
        RECT 6.5750 35.3835 6.6010 36.4770 ;
        RECT 6.4670 35.3835 6.4930 36.4770 ;
        RECT 6.3590 35.3835 6.3850 36.4770 ;
        RECT 6.2510 35.3835 6.2770 36.4770 ;
        RECT 6.1430 35.3835 6.1690 36.4770 ;
        RECT 6.0350 35.3835 6.0610 36.4770 ;
        RECT 5.9270 35.3835 5.9530 36.4770 ;
        RECT 5.7140 35.3835 5.7910 36.4770 ;
        RECT 3.8210 35.3835 3.8980 36.4770 ;
        RECT 3.6590 35.3835 3.6850 36.4770 ;
        RECT 3.5510 35.3835 3.5770 36.4770 ;
        RECT 3.4430 35.3835 3.4690 36.4770 ;
        RECT 3.3350 35.3835 3.3610 36.4770 ;
        RECT 3.2270 35.3835 3.2530 36.4770 ;
        RECT 3.1190 35.3835 3.1450 36.4770 ;
        RECT 3.0110 35.3835 3.0370 36.4770 ;
        RECT 2.9030 35.3835 2.9290 36.4770 ;
        RECT 2.7950 35.3835 2.8210 36.4770 ;
        RECT 2.6870 35.3835 2.7130 36.4770 ;
        RECT 2.5790 35.3835 2.6050 36.4770 ;
        RECT 2.4710 35.3835 2.4970 36.4770 ;
        RECT 2.3630 35.3835 2.3890 36.4770 ;
        RECT 2.2550 35.3835 2.2810 36.4770 ;
        RECT 2.1470 35.3835 2.1730 36.4770 ;
        RECT 2.0390 35.3835 2.0650 36.4770 ;
        RECT 1.9310 35.3835 1.9570 36.4770 ;
        RECT 1.8230 35.3835 1.8490 36.4770 ;
        RECT 1.7150 35.3835 1.7410 36.4770 ;
        RECT 1.6070 35.3835 1.6330 36.4770 ;
        RECT 1.4990 35.3835 1.5250 36.4770 ;
        RECT 1.3910 35.3835 1.4170 36.4770 ;
        RECT 1.2830 35.3835 1.3090 36.4770 ;
        RECT 1.1750 35.3835 1.2010 36.4770 ;
        RECT 1.0670 35.3835 1.0930 36.4770 ;
        RECT 0.9590 35.3835 0.9850 36.4770 ;
        RECT 0.8510 35.3835 0.8770 36.4770 ;
        RECT 0.7430 35.3835 0.7690 36.4770 ;
        RECT 0.6350 35.3835 0.6610 36.4770 ;
        RECT 0.5270 35.3835 0.5530 36.4770 ;
        RECT 0.4190 35.3835 0.4450 36.4770 ;
        RECT 0.3110 35.3835 0.3370 36.4770 ;
        RECT 0.2030 35.3835 0.2290 36.4770 ;
        RECT 0.0000 35.3835 0.0850 36.4770 ;
        RECT 5.1800 36.4635 5.3080 37.5570 ;
        RECT 5.1660 37.1290 5.3080 37.4515 ;
        RECT 5.0180 36.8560 5.0800 37.5570 ;
        RECT 5.0040 37.1655 5.0800 37.3190 ;
        RECT 5.0180 36.4635 5.0440 37.5570 ;
        RECT 5.0180 36.5845 5.0580 36.8240 ;
        RECT 5.0180 36.4635 5.0800 36.5525 ;
        RECT 4.7210 36.9140 4.9270 37.5570 ;
        RECT 4.9010 36.4635 4.9270 37.5570 ;
        RECT 4.7210 37.1910 4.9410 37.4490 ;
        RECT 4.7210 36.4635 4.8190 37.5570 ;
        RECT 4.3040 36.4635 4.3870 37.5570 ;
        RECT 4.3040 36.5520 4.4010 37.4875 ;
        RECT 9.5270 36.4635 9.6120 37.5570 ;
        RECT 9.3830 36.4635 9.4090 37.5570 ;
        RECT 9.2750 36.4635 9.3010 37.5570 ;
        RECT 9.1670 36.4635 9.1930 37.5570 ;
        RECT 9.0590 36.4635 9.0850 37.5570 ;
        RECT 8.9510 36.4635 8.9770 37.5570 ;
        RECT 8.8430 36.4635 8.8690 37.5570 ;
        RECT 8.7350 36.4635 8.7610 37.5570 ;
        RECT 8.6270 36.4635 8.6530 37.5570 ;
        RECT 8.5190 36.4635 8.5450 37.5570 ;
        RECT 8.4110 36.4635 8.4370 37.5570 ;
        RECT 8.3030 36.4635 8.3290 37.5570 ;
        RECT 8.1950 36.4635 8.2210 37.5570 ;
        RECT 8.0870 36.4635 8.1130 37.5570 ;
        RECT 7.9790 36.4635 8.0050 37.5570 ;
        RECT 7.8710 36.4635 7.8970 37.5570 ;
        RECT 7.7630 36.4635 7.7890 37.5570 ;
        RECT 7.6550 36.4635 7.6810 37.5570 ;
        RECT 7.5470 36.4635 7.5730 37.5570 ;
        RECT 7.4390 36.4635 7.4650 37.5570 ;
        RECT 7.3310 36.4635 7.3570 37.5570 ;
        RECT 7.2230 36.4635 7.2490 37.5570 ;
        RECT 7.1150 36.4635 7.1410 37.5570 ;
        RECT 7.0070 36.4635 7.0330 37.5570 ;
        RECT 6.8990 36.4635 6.9250 37.5570 ;
        RECT 6.7910 36.4635 6.8170 37.5570 ;
        RECT 6.6830 36.4635 6.7090 37.5570 ;
        RECT 6.5750 36.4635 6.6010 37.5570 ;
        RECT 6.4670 36.4635 6.4930 37.5570 ;
        RECT 6.3590 36.4635 6.3850 37.5570 ;
        RECT 6.2510 36.4635 6.2770 37.5570 ;
        RECT 6.1430 36.4635 6.1690 37.5570 ;
        RECT 6.0350 36.4635 6.0610 37.5570 ;
        RECT 5.9270 36.4635 5.9530 37.5570 ;
        RECT 5.7140 36.4635 5.7910 37.5570 ;
        RECT 3.8210 36.4635 3.8980 37.5570 ;
        RECT 3.6590 36.4635 3.6850 37.5570 ;
        RECT 3.5510 36.4635 3.5770 37.5570 ;
        RECT 3.4430 36.4635 3.4690 37.5570 ;
        RECT 3.3350 36.4635 3.3610 37.5570 ;
        RECT 3.2270 36.4635 3.2530 37.5570 ;
        RECT 3.1190 36.4635 3.1450 37.5570 ;
        RECT 3.0110 36.4635 3.0370 37.5570 ;
        RECT 2.9030 36.4635 2.9290 37.5570 ;
        RECT 2.7950 36.4635 2.8210 37.5570 ;
        RECT 2.6870 36.4635 2.7130 37.5570 ;
        RECT 2.5790 36.4635 2.6050 37.5570 ;
        RECT 2.4710 36.4635 2.4970 37.5570 ;
        RECT 2.3630 36.4635 2.3890 37.5570 ;
        RECT 2.2550 36.4635 2.2810 37.5570 ;
        RECT 2.1470 36.4635 2.1730 37.5570 ;
        RECT 2.0390 36.4635 2.0650 37.5570 ;
        RECT 1.9310 36.4635 1.9570 37.5570 ;
        RECT 1.8230 36.4635 1.8490 37.5570 ;
        RECT 1.7150 36.4635 1.7410 37.5570 ;
        RECT 1.6070 36.4635 1.6330 37.5570 ;
        RECT 1.4990 36.4635 1.5250 37.5570 ;
        RECT 1.3910 36.4635 1.4170 37.5570 ;
        RECT 1.2830 36.4635 1.3090 37.5570 ;
        RECT 1.1750 36.4635 1.2010 37.5570 ;
        RECT 1.0670 36.4635 1.0930 37.5570 ;
        RECT 0.9590 36.4635 0.9850 37.5570 ;
        RECT 0.8510 36.4635 0.8770 37.5570 ;
        RECT 0.7430 36.4635 0.7690 37.5570 ;
        RECT 0.6350 36.4635 0.6610 37.5570 ;
        RECT 0.5270 36.4635 0.5530 37.5570 ;
        RECT 0.4190 36.4635 0.4450 37.5570 ;
        RECT 0.3110 36.4635 0.3370 37.5570 ;
        RECT 0.2030 36.4635 0.2290 37.5570 ;
        RECT 0.0000 36.4635 0.0850 37.5570 ;
        RECT 5.1800 37.5435 5.3080 38.6370 ;
        RECT 5.1660 38.2090 5.3080 38.5315 ;
        RECT 5.0180 37.9360 5.0800 38.6370 ;
        RECT 5.0040 38.2455 5.0800 38.3990 ;
        RECT 5.0180 37.5435 5.0440 38.6370 ;
        RECT 5.0180 37.6645 5.0580 37.9040 ;
        RECT 5.0180 37.5435 5.0800 37.6325 ;
        RECT 4.7210 37.9940 4.9270 38.6370 ;
        RECT 4.9010 37.5435 4.9270 38.6370 ;
        RECT 4.7210 38.2710 4.9410 38.5290 ;
        RECT 4.7210 37.5435 4.8190 38.6370 ;
        RECT 4.3040 37.5435 4.3870 38.6370 ;
        RECT 4.3040 37.6320 4.4010 38.5675 ;
        RECT 9.5270 37.5435 9.6120 38.6370 ;
        RECT 9.3830 37.5435 9.4090 38.6370 ;
        RECT 9.2750 37.5435 9.3010 38.6370 ;
        RECT 9.1670 37.5435 9.1930 38.6370 ;
        RECT 9.0590 37.5435 9.0850 38.6370 ;
        RECT 8.9510 37.5435 8.9770 38.6370 ;
        RECT 8.8430 37.5435 8.8690 38.6370 ;
        RECT 8.7350 37.5435 8.7610 38.6370 ;
        RECT 8.6270 37.5435 8.6530 38.6370 ;
        RECT 8.5190 37.5435 8.5450 38.6370 ;
        RECT 8.4110 37.5435 8.4370 38.6370 ;
        RECT 8.3030 37.5435 8.3290 38.6370 ;
        RECT 8.1950 37.5435 8.2210 38.6370 ;
        RECT 8.0870 37.5435 8.1130 38.6370 ;
        RECT 7.9790 37.5435 8.0050 38.6370 ;
        RECT 7.8710 37.5435 7.8970 38.6370 ;
        RECT 7.7630 37.5435 7.7890 38.6370 ;
        RECT 7.6550 37.5435 7.6810 38.6370 ;
        RECT 7.5470 37.5435 7.5730 38.6370 ;
        RECT 7.4390 37.5435 7.4650 38.6370 ;
        RECT 7.3310 37.5435 7.3570 38.6370 ;
        RECT 7.2230 37.5435 7.2490 38.6370 ;
        RECT 7.1150 37.5435 7.1410 38.6370 ;
        RECT 7.0070 37.5435 7.0330 38.6370 ;
        RECT 6.8990 37.5435 6.9250 38.6370 ;
        RECT 6.7910 37.5435 6.8170 38.6370 ;
        RECT 6.6830 37.5435 6.7090 38.6370 ;
        RECT 6.5750 37.5435 6.6010 38.6370 ;
        RECT 6.4670 37.5435 6.4930 38.6370 ;
        RECT 6.3590 37.5435 6.3850 38.6370 ;
        RECT 6.2510 37.5435 6.2770 38.6370 ;
        RECT 6.1430 37.5435 6.1690 38.6370 ;
        RECT 6.0350 37.5435 6.0610 38.6370 ;
        RECT 5.9270 37.5435 5.9530 38.6370 ;
        RECT 5.7140 37.5435 5.7910 38.6370 ;
        RECT 3.8210 37.5435 3.8980 38.6370 ;
        RECT 3.6590 37.5435 3.6850 38.6370 ;
        RECT 3.5510 37.5435 3.5770 38.6370 ;
        RECT 3.4430 37.5435 3.4690 38.6370 ;
        RECT 3.3350 37.5435 3.3610 38.6370 ;
        RECT 3.2270 37.5435 3.2530 38.6370 ;
        RECT 3.1190 37.5435 3.1450 38.6370 ;
        RECT 3.0110 37.5435 3.0370 38.6370 ;
        RECT 2.9030 37.5435 2.9290 38.6370 ;
        RECT 2.7950 37.5435 2.8210 38.6370 ;
        RECT 2.6870 37.5435 2.7130 38.6370 ;
        RECT 2.5790 37.5435 2.6050 38.6370 ;
        RECT 2.4710 37.5435 2.4970 38.6370 ;
        RECT 2.3630 37.5435 2.3890 38.6370 ;
        RECT 2.2550 37.5435 2.2810 38.6370 ;
        RECT 2.1470 37.5435 2.1730 38.6370 ;
        RECT 2.0390 37.5435 2.0650 38.6370 ;
        RECT 1.9310 37.5435 1.9570 38.6370 ;
        RECT 1.8230 37.5435 1.8490 38.6370 ;
        RECT 1.7150 37.5435 1.7410 38.6370 ;
        RECT 1.6070 37.5435 1.6330 38.6370 ;
        RECT 1.4990 37.5435 1.5250 38.6370 ;
        RECT 1.3910 37.5435 1.4170 38.6370 ;
        RECT 1.2830 37.5435 1.3090 38.6370 ;
        RECT 1.1750 37.5435 1.2010 38.6370 ;
        RECT 1.0670 37.5435 1.0930 38.6370 ;
        RECT 0.9590 37.5435 0.9850 38.6370 ;
        RECT 0.8510 37.5435 0.8770 38.6370 ;
        RECT 0.7430 37.5435 0.7690 38.6370 ;
        RECT 0.6350 37.5435 0.6610 38.6370 ;
        RECT 0.5270 37.5435 0.5530 38.6370 ;
        RECT 0.4190 37.5435 0.4450 38.6370 ;
        RECT 0.3110 37.5435 0.3370 38.6370 ;
        RECT 0.2030 37.5435 0.2290 38.6370 ;
        RECT 0.0000 37.5435 0.0850 38.6370 ;
        RECT 5.1800 38.6235 5.3080 39.7170 ;
        RECT 5.1660 39.2890 5.3080 39.6115 ;
        RECT 5.0180 39.0160 5.0800 39.7170 ;
        RECT 5.0040 39.3255 5.0800 39.4790 ;
        RECT 5.0180 38.6235 5.0440 39.7170 ;
        RECT 5.0180 38.7445 5.0580 38.9840 ;
        RECT 5.0180 38.6235 5.0800 38.7125 ;
        RECT 4.7210 39.0740 4.9270 39.7170 ;
        RECT 4.9010 38.6235 4.9270 39.7170 ;
        RECT 4.7210 39.3510 4.9410 39.6090 ;
        RECT 4.7210 38.6235 4.8190 39.7170 ;
        RECT 4.3040 38.6235 4.3870 39.7170 ;
        RECT 4.3040 38.7120 4.4010 39.6475 ;
        RECT 9.5270 38.6235 9.6120 39.7170 ;
        RECT 9.3830 38.6235 9.4090 39.7170 ;
        RECT 9.2750 38.6235 9.3010 39.7170 ;
        RECT 9.1670 38.6235 9.1930 39.7170 ;
        RECT 9.0590 38.6235 9.0850 39.7170 ;
        RECT 8.9510 38.6235 8.9770 39.7170 ;
        RECT 8.8430 38.6235 8.8690 39.7170 ;
        RECT 8.7350 38.6235 8.7610 39.7170 ;
        RECT 8.6270 38.6235 8.6530 39.7170 ;
        RECT 8.5190 38.6235 8.5450 39.7170 ;
        RECT 8.4110 38.6235 8.4370 39.7170 ;
        RECT 8.3030 38.6235 8.3290 39.7170 ;
        RECT 8.1950 38.6235 8.2210 39.7170 ;
        RECT 8.0870 38.6235 8.1130 39.7170 ;
        RECT 7.9790 38.6235 8.0050 39.7170 ;
        RECT 7.8710 38.6235 7.8970 39.7170 ;
        RECT 7.7630 38.6235 7.7890 39.7170 ;
        RECT 7.6550 38.6235 7.6810 39.7170 ;
        RECT 7.5470 38.6235 7.5730 39.7170 ;
        RECT 7.4390 38.6235 7.4650 39.7170 ;
        RECT 7.3310 38.6235 7.3570 39.7170 ;
        RECT 7.2230 38.6235 7.2490 39.7170 ;
        RECT 7.1150 38.6235 7.1410 39.7170 ;
        RECT 7.0070 38.6235 7.0330 39.7170 ;
        RECT 6.8990 38.6235 6.9250 39.7170 ;
        RECT 6.7910 38.6235 6.8170 39.7170 ;
        RECT 6.6830 38.6235 6.7090 39.7170 ;
        RECT 6.5750 38.6235 6.6010 39.7170 ;
        RECT 6.4670 38.6235 6.4930 39.7170 ;
        RECT 6.3590 38.6235 6.3850 39.7170 ;
        RECT 6.2510 38.6235 6.2770 39.7170 ;
        RECT 6.1430 38.6235 6.1690 39.7170 ;
        RECT 6.0350 38.6235 6.0610 39.7170 ;
        RECT 5.9270 38.6235 5.9530 39.7170 ;
        RECT 5.7140 38.6235 5.7910 39.7170 ;
        RECT 3.8210 38.6235 3.8980 39.7170 ;
        RECT 3.6590 38.6235 3.6850 39.7170 ;
        RECT 3.5510 38.6235 3.5770 39.7170 ;
        RECT 3.4430 38.6235 3.4690 39.7170 ;
        RECT 3.3350 38.6235 3.3610 39.7170 ;
        RECT 3.2270 38.6235 3.2530 39.7170 ;
        RECT 3.1190 38.6235 3.1450 39.7170 ;
        RECT 3.0110 38.6235 3.0370 39.7170 ;
        RECT 2.9030 38.6235 2.9290 39.7170 ;
        RECT 2.7950 38.6235 2.8210 39.7170 ;
        RECT 2.6870 38.6235 2.7130 39.7170 ;
        RECT 2.5790 38.6235 2.6050 39.7170 ;
        RECT 2.4710 38.6235 2.4970 39.7170 ;
        RECT 2.3630 38.6235 2.3890 39.7170 ;
        RECT 2.2550 38.6235 2.2810 39.7170 ;
        RECT 2.1470 38.6235 2.1730 39.7170 ;
        RECT 2.0390 38.6235 2.0650 39.7170 ;
        RECT 1.9310 38.6235 1.9570 39.7170 ;
        RECT 1.8230 38.6235 1.8490 39.7170 ;
        RECT 1.7150 38.6235 1.7410 39.7170 ;
        RECT 1.6070 38.6235 1.6330 39.7170 ;
        RECT 1.4990 38.6235 1.5250 39.7170 ;
        RECT 1.3910 38.6235 1.4170 39.7170 ;
        RECT 1.2830 38.6235 1.3090 39.7170 ;
        RECT 1.1750 38.6235 1.2010 39.7170 ;
        RECT 1.0670 38.6235 1.0930 39.7170 ;
        RECT 0.9590 38.6235 0.9850 39.7170 ;
        RECT 0.8510 38.6235 0.8770 39.7170 ;
        RECT 0.7430 38.6235 0.7690 39.7170 ;
        RECT 0.6350 38.6235 0.6610 39.7170 ;
        RECT 0.5270 38.6235 0.5530 39.7170 ;
        RECT 0.4190 38.6235 0.4450 39.7170 ;
        RECT 0.3110 38.6235 0.3370 39.7170 ;
        RECT 0.2030 38.6235 0.2290 39.7170 ;
        RECT 0.0000 38.6235 0.0850 39.7170 ;
        RECT 5.1800 39.7035 5.3080 40.7970 ;
        RECT 5.1660 40.3690 5.3080 40.6915 ;
        RECT 5.0180 40.0960 5.0800 40.7970 ;
        RECT 5.0040 40.4055 5.0800 40.5590 ;
        RECT 5.0180 39.7035 5.0440 40.7970 ;
        RECT 5.0180 39.8245 5.0580 40.0640 ;
        RECT 5.0180 39.7035 5.0800 39.7925 ;
        RECT 4.7210 40.1540 4.9270 40.7970 ;
        RECT 4.9010 39.7035 4.9270 40.7970 ;
        RECT 4.7210 40.4310 4.9410 40.6890 ;
        RECT 4.7210 39.7035 4.8190 40.7970 ;
        RECT 4.3040 39.7035 4.3870 40.7970 ;
        RECT 4.3040 39.7920 4.4010 40.7275 ;
        RECT 9.5270 39.7035 9.6120 40.7970 ;
        RECT 9.3830 39.7035 9.4090 40.7970 ;
        RECT 9.2750 39.7035 9.3010 40.7970 ;
        RECT 9.1670 39.7035 9.1930 40.7970 ;
        RECT 9.0590 39.7035 9.0850 40.7970 ;
        RECT 8.9510 39.7035 8.9770 40.7970 ;
        RECT 8.8430 39.7035 8.8690 40.7970 ;
        RECT 8.7350 39.7035 8.7610 40.7970 ;
        RECT 8.6270 39.7035 8.6530 40.7970 ;
        RECT 8.5190 39.7035 8.5450 40.7970 ;
        RECT 8.4110 39.7035 8.4370 40.7970 ;
        RECT 8.3030 39.7035 8.3290 40.7970 ;
        RECT 8.1950 39.7035 8.2210 40.7970 ;
        RECT 8.0870 39.7035 8.1130 40.7970 ;
        RECT 7.9790 39.7035 8.0050 40.7970 ;
        RECT 7.8710 39.7035 7.8970 40.7970 ;
        RECT 7.7630 39.7035 7.7890 40.7970 ;
        RECT 7.6550 39.7035 7.6810 40.7970 ;
        RECT 7.5470 39.7035 7.5730 40.7970 ;
        RECT 7.4390 39.7035 7.4650 40.7970 ;
        RECT 7.3310 39.7035 7.3570 40.7970 ;
        RECT 7.2230 39.7035 7.2490 40.7970 ;
        RECT 7.1150 39.7035 7.1410 40.7970 ;
        RECT 7.0070 39.7035 7.0330 40.7970 ;
        RECT 6.8990 39.7035 6.9250 40.7970 ;
        RECT 6.7910 39.7035 6.8170 40.7970 ;
        RECT 6.6830 39.7035 6.7090 40.7970 ;
        RECT 6.5750 39.7035 6.6010 40.7970 ;
        RECT 6.4670 39.7035 6.4930 40.7970 ;
        RECT 6.3590 39.7035 6.3850 40.7970 ;
        RECT 6.2510 39.7035 6.2770 40.7970 ;
        RECT 6.1430 39.7035 6.1690 40.7970 ;
        RECT 6.0350 39.7035 6.0610 40.7970 ;
        RECT 5.9270 39.7035 5.9530 40.7970 ;
        RECT 5.7140 39.7035 5.7910 40.7970 ;
        RECT 3.8210 39.7035 3.8980 40.7970 ;
        RECT 3.6590 39.7035 3.6850 40.7970 ;
        RECT 3.5510 39.7035 3.5770 40.7970 ;
        RECT 3.4430 39.7035 3.4690 40.7970 ;
        RECT 3.3350 39.7035 3.3610 40.7970 ;
        RECT 3.2270 39.7035 3.2530 40.7970 ;
        RECT 3.1190 39.7035 3.1450 40.7970 ;
        RECT 3.0110 39.7035 3.0370 40.7970 ;
        RECT 2.9030 39.7035 2.9290 40.7970 ;
        RECT 2.7950 39.7035 2.8210 40.7970 ;
        RECT 2.6870 39.7035 2.7130 40.7970 ;
        RECT 2.5790 39.7035 2.6050 40.7970 ;
        RECT 2.4710 39.7035 2.4970 40.7970 ;
        RECT 2.3630 39.7035 2.3890 40.7970 ;
        RECT 2.2550 39.7035 2.2810 40.7970 ;
        RECT 2.1470 39.7035 2.1730 40.7970 ;
        RECT 2.0390 39.7035 2.0650 40.7970 ;
        RECT 1.9310 39.7035 1.9570 40.7970 ;
        RECT 1.8230 39.7035 1.8490 40.7970 ;
        RECT 1.7150 39.7035 1.7410 40.7970 ;
        RECT 1.6070 39.7035 1.6330 40.7970 ;
        RECT 1.4990 39.7035 1.5250 40.7970 ;
        RECT 1.3910 39.7035 1.4170 40.7970 ;
        RECT 1.2830 39.7035 1.3090 40.7970 ;
        RECT 1.1750 39.7035 1.2010 40.7970 ;
        RECT 1.0670 39.7035 1.0930 40.7970 ;
        RECT 0.9590 39.7035 0.9850 40.7970 ;
        RECT 0.8510 39.7035 0.8770 40.7970 ;
        RECT 0.7430 39.7035 0.7690 40.7970 ;
        RECT 0.6350 39.7035 0.6610 40.7970 ;
        RECT 0.5270 39.7035 0.5530 40.7970 ;
        RECT 0.4190 39.7035 0.4450 40.7970 ;
        RECT 0.3110 39.7035 0.3370 40.7970 ;
        RECT 0.2030 39.7035 0.2290 40.7970 ;
        RECT 0.0000 39.7035 0.0850 40.7970 ;
        RECT 5.1800 40.7835 5.3080 41.8770 ;
        RECT 5.1660 41.4490 5.3080 41.7715 ;
        RECT 5.0180 41.1760 5.0800 41.8770 ;
        RECT 5.0040 41.4855 5.0800 41.6390 ;
        RECT 5.0180 40.7835 5.0440 41.8770 ;
        RECT 5.0180 40.9045 5.0580 41.1440 ;
        RECT 5.0180 40.7835 5.0800 40.8725 ;
        RECT 4.7210 41.2340 4.9270 41.8770 ;
        RECT 4.9010 40.7835 4.9270 41.8770 ;
        RECT 4.7210 41.5110 4.9410 41.7690 ;
        RECT 4.7210 40.7835 4.8190 41.8770 ;
        RECT 4.3040 40.7835 4.3870 41.8770 ;
        RECT 4.3040 40.8720 4.4010 41.8075 ;
        RECT 9.5270 40.7835 9.6120 41.8770 ;
        RECT 9.3830 40.7835 9.4090 41.8770 ;
        RECT 9.2750 40.7835 9.3010 41.8770 ;
        RECT 9.1670 40.7835 9.1930 41.8770 ;
        RECT 9.0590 40.7835 9.0850 41.8770 ;
        RECT 8.9510 40.7835 8.9770 41.8770 ;
        RECT 8.8430 40.7835 8.8690 41.8770 ;
        RECT 8.7350 40.7835 8.7610 41.8770 ;
        RECT 8.6270 40.7835 8.6530 41.8770 ;
        RECT 8.5190 40.7835 8.5450 41.8770 ;
        RECT 8.4110 40.7835 8.4370 41.8770 ;
        RECT 8.3030 40.7835 8.3290 41.8770 ;
        RECT 8.1950 40.7835 8.2210 41.8770 ;
        RECT 8.0870 40.7835 8.1130 41.8770 ;
        RECT 7.9790 40.7835 8.0050 41.8770 ;
        RECT 7.8710 40.7835 7.8970 41.8770 ;
        RECT 7.7630 40.7835 7.7890 41.8770 ;
        RECT 7.6550 40.7835 7.6810 41.8770 ;
        RECT 7.5470 40.7835 7.5730 41.8770 ;
        RECT 7.4390 40.7835 7.4650 41.8770 ;
        RECT 7.3310 40.7835 7.3570 41.8770 ;
        RECT 7.2230 40.7835 7.2490 41.8770 ;
        RECT 7.1150 40.7835 7.1410 41.8770 ;
        RECT 7.0070 40.7835 7.0330 41.8770 ;
        RECT 6.8990 40.7835 6.9250 41.8770 ;
        RECT 6.7910 40.7835 6.8170 41.8770 ;
        RECT 6.6830 40.7835 6.7090 41.8770 ;
        RECT 6.5750 40.7835 6.6010 41.8770 ;
        RECT 6.4670 40.7835 6.4930 41.8770 ;
        RECT 6.3590 40.7835 6.3850 41.8770 ;
        RECT 6.2510 40.7835 6.2770 41.8770 ;
        RECT 6.1430 40.7835 6.1690 41.8770 ;
        RECT 6.0350 40.7835 6.0610 41.8770 ;
        RECT 5.9270 40.7835 5.9530 41.8770 ;
        RECT 5.7140 40.7835 5.7910 41.8770 ;
        RECT 3.8210 40.7835 3.8980 41.8770 ;
        RECT 3.6590 40.7835 3.6850 41.8770 ;
        RECT 3.5510 40.7835 3.5770 41.8770 ;
        RECT 3.4430 40.7835 3.4690 41.8770 ;
        RECT 3.3350 40.7835 3.3610 41.8770 ;
        RECT 3.2270 40.7835 3.2530 41.8770 ;
        RECT 3.1190 40.7835 3.1450 41.8770 ;
        RECT 3.0110 40.7835 3.0370 41.8770 ;
        RECT 2.9030 40.7835 2.9290 41.8770 ;
        RECT 2.7950 40.7835 2.8210 41.8770 ;
        RECT 2.6870 40.7835 2.7130 41.8770 ;
        RECT 2.5790 40.7835 2.6050 41.8770 ;
        RECT 2.4710 40.7835 2.4970 41.8770 ;
        RECT 2.3630 40.7835 2.3890 41.8770 ;
        RECT 2.2550 40.7835 2.2810 41.8770 ;
        RECT 2.1470 40.7835 2.1730 41.8770 ;
        RECT 2.0390 40.7835 2.0650 41.8770 ;
        RECT 1.9310 40.7835 1.9570 41.8770 ;
        RECT 1.8230 40.7835 1.8490 41.8770 ;
        RECT 1.7150 40.7835 1.7410 41.8770 ;
        RECT 1.6070 40.7835 1.6330 41.8770 ;
        RECT 1.4990 40.7835 1.5250 41.8770 ;
        RECT 1.3910 40.7835 1.4170 41.8770 ;
        RECT 1.2830 40.7835 1.3090 41.8770 ;
        RECT 1.1750 40.7835 1.2010 41.8770 ;
        RECT 1.0670 40.7835 1.0930 41.8770 ;
        RECT 0.9590 40.7835 0.9850 41.8770 ;
        RECT 0.8510 40.7835 0.8770 41.8770 ;
        RECT 0.7430 40.7835 0.7690 41.8770 ;
        RECT 0.6350 40.7835 0.6610 41.8770 ;
        RECT 0.5270 40.7835 0.5530 41.8770 ;
        RECT 0.4190 40.7835 0.4450 41.8770 ;
        RECT 0.3110 40.7835 0.3370 41.8770 ;
        RECT 0.2030 40.7835 0.2290 41.8770 ;
        RECT 0.0000 40.7835 0.0850 41.8770 ;
        RECT 5.1800 41.8635 5.3080 42.9570 ;
        RECT 5.1660 42.5290 5.3080 42.8515 ;
        RECT 5.0180 42.2560 5.0800 42.9570 ;
        RECT 5.0040 42.5655 5.0800 42.7190 ;
        RECT 5.0180 41.8635 5.0440 42.9570 ;
        RECT 5.0180 41.9845 5.0580 42.2240 ;
        RECT 5.0180 41.8635 5.0800 41.9525 ;
        RECT 4.7210 42.3140 4.9270 42.9570 ;
        RECT 4.9010 41.8635 4.9270 42.9570 ;
        RECT 4.7210 42.5910 4.9410 42.8490 ;
        RECT 4.7210 41.8635 4.8190 42.9570 ;
        RECT 4.3040 41.8635 4.3870 42.9570 ;
        RECT 4.3040 41.9520 4.4010 42.8875 ;
        RECT 9.5270 41.8635 9.6120 42.9570 ;
        RECT 9.3830 41.8635 9.4090 42.9570 ;
        RECT 9.2750 41.8635 9.3010 42.9570 ;
        RECT 9.1670 41.8635 9.1930 42.9570 ;
        RECT 9.0590 41.8635 9.0850 42.9570 ;
        RECT 8.9510 41.8635 8.9770 42.9570 ;
        RECT 8.8430 41.8635 8.8690 42.9570 ;
        RECT 8.7350 41.8635 8.7610 42.9570 ;
        RECT 8.6270 41.8635 8.6530 42.9570 ;
        RECT 8.5190 41.8635 8.5450 42.9570 ;
        RECT 8.4110 41.8635 8.4370 42.9570 ;
        RECT 8.3030 41.8635 8.3290 42.9570 ;
        RECT 8.1950 41.8635 8.2210 42.9570 ;
        RECT 8.0870 41.8635 8.1130 42.9570 ;
        RECT 7.9790 41.8635 8.0050 42.9570 ;
        RECT 7.8710 41.8635 7.8970 42.9570 ;
        RECT 7.7630 41.8635 7.7890 42.9570 ;
        RECT 7.6550 41.8635 7.6810 42.9570 ;
        RECT 7.5470 41.8635 7.5730 42.9570 ;
        RECT 7.4390 41.8635 7.4650 42.9570 ;
        RECT 7.3310 41.8635 7.3570 42.9570 ;
        RECT 7.2230 41.8635 7.2490 42.9570 ;
        RECT 7.1150 41.8635 7.1410 42.9570 ;
        RECT 7.0070 41.8635 7.0330 42.9570 ;
        RECT 6.8990 41.8635 6.9250 42.9570 ;
        RECT 6.7910 41.8635 6.8170 42.9570 ;
        RECT 6.6830 41.8635 6.7090 42.9570 ;
        RECT 6.5750 41.8635 6.6010 42.9570 ;
        RECT 6.4670 41.8635 6.4930 42.9570 ;
        RECT 6.3590 41.8635 6.3850 42.9570 ;
        RECT 6.2510 41.8635 6.2770 42.9570 ;
        RECT 6.1430 41.8635 6.1690 42.9570 ;
        RECT 6.0350 41.8635 6.0610 42.9570 ;
        RECT 5.9270 41.8635 5.9530 42.9570 ;
        RECT 5.7140 41.8635 5.7910 42.9570 ;
        RECT 3.8210 41.8635 3.8980 42.9570 ;
        RECT 3.6590 41.8635 3.6850 42.9570 ;
        RECT 3.5510 41.8635 3.5770 42.9570 ;
        RECT 3.4430 41.8635 3.4690 42.9570 ;
        RECT 3.3350 41.8635 3.3610 42.9570 ;
        RECT 3.2270 41.8635 3.2530 42.9570 ;
        RECT 3.1190 41.8635 3.1450 42.9570 ;
        RECT 3.0110 41.8635 3.0370 42.9570 ;
        RECT 2.9030 41.8635 2.9290 42.9570 ;
        RECT 2.7950 41.8635 2.8210 42.9570 ;
        RECT 2.6870 41.8635 2.7130 42.9570 ;
        RECT 2.5790 41.8635 2.6050 42.9570 ;
        RECT 2.4710 41.8635 2.4970 42.9570 ;
        RECT 2.3630 41.8635 2.3890 42.9570 ;
        RECT 2.2550 41.8635 2.2810 42.9570 ;
        RECT 2.1470 41.8635 2.1730 42.9570 ;
        RECT 2.0390 41.8635 2.0650 42.9570 ;
        RECT 1.9310 41.8635 1.9570 42.9570 ;
        RECT 1.8230 41.8635 1.8490 42.9570 ;
        RECT 1.7150 41.8635 1.7410 42.9570 ;
        RECT 1.6070 41.8635 1.6330 42.9570 ;
        RECT 1.4990 41.8635 1.5250 42.9570 ;
        RECT 1.3910 41.8635 1.4170 42.9570 ;
        RECT 1.2830 41.8635 1.3090 42.9570 ;
        RECT 1.1750 41.8635 1.2010 42.9570 ;
        RECT 1.0670 41.8635 1.0930 42.9570 ;
        RECT 0.9590 41.8635 0.9850 42.9570 ;
        RECT 0.8510 41.8635 0.8770 42.9570 ;
        RECT 0.7430 41.8635 0.7690 42.9570 ;
        RECT 0.6350 41.8635 0.6610 42.9570 ;
        RECT 0.5270 41.8635 0.5530 42.9570 ;
        RECT 0.4190 41.8635 0.4450 42.9570 ;
        RECT 0.3110 41.8635 0.3370 42.9570 ;
        RECT 0.2030 41.8635 0.2290 42.9570 ;
        RECT 0.0000 41.8635 0.0850 42.9570 ;
  LAYER V3  ;
      RECT 0.0000 1.2200 9.6120 1.3500 ;
      RECT 9.4950 0.2565 9.6120 1.3500 ;
      RECT 5.8410 1.1240 9.4770 1.3500 ;
      RECT 4.5090 1.1240 5.8230 1.3500 ;
      RECT 3.7890 0.2565 4.4190 1.3500 ;
      RECT 0.1350 1.1240 3.7710 1.3500 ;
      RECT 0.0000 0.2565 0.1170 1.3500 ;
      RECT 9.4590 0.2565 9.6120 1.1720 ;
      RECT 5.8950 0.2565 9.4410 1.3500 ;
      RECT 5.1480 0.2565 5.8770 1.1720 ;
      RECT 4.9860 0.4520 5.1120 1.3500 ;
      RECT 3.7350 0.3560 4.9590 1.1720 ;
      RECT 0.1710 0.2565 3.7170 1.3500 ;
      RECT 0.0000 0.2565 0.1530 1.1720 ;
      RECT 5.0940 0.2565 9.6120 1.0760 ;
      RECT 0.0000 0.3560 5.0760 1.0760 ;
      RECT 4.8690 0.2565 9.6120 0.4280 ;
      RECT 0.0000 0.2565 4.8510 1.0760 ;
      RECT 0.0000 0.2565 9.6120 0.3320 ;
      RECT 0.0000 2.3000 9.6120 2.4300 ;
      RECT 9.4950 1.3365 9.6120 2.4300 ;
      RECT 5.8410 2.2040 9.4770 2.4300 ;
      RECT 4.5090 2.2040 5.8230 2.4300 ;
      RECT 3.7890 1.3365 4.4190 2.4300 ;
      RECT 0.1350 2.2040 3.7710 2.4300 ;
      RECT 0.0000 1.3365 0.1170 2.4300 ;
      RECT 9.4590 1.3365 9.6120 2.2520 ;
      RECT 5.8950 1.3365 9.4410 2.4300 ;
      RECT 5.1480 1.3365 5.8770 2.2520 ;
      RECT 4.9860 1.5320 5.1120 2.4300 ;
      RECT 3.7350 1.4360 4.9590 2.2520 ;
      RECT 0.1710 1.3365 3.7170 2.4300 ;
      RECT 0.0000 1.3365 0.1530 2.2520 ;
      RECT 5.0940 1.3365 9.6120 2.1560 ;
      RECT 0.0000 1.4360 5.0760 2.1560 ;
      RECT 4.8690 1.3365 9.6120 1.5080 ;
      RECT 0.0000 1.3365 4.8510 2.1560 ;
      RECT 0.0000 1.3365 9.6120 1.4120 ;
      RECT 0.0000 3.3800 9.6120 3.5100 ;
      RECT 9.4950 2.4165 9.6120 3.5100 ;
      RECT 5.8410 3.2840 9.4770 3.5100 ;
      RECT 4.5090 3.2840 5.8230 3.5100 ;
      RECT 3.7890 2.4165 4.4190 3.5100 ;
      RECT 0.1350 3.2840 3.7710 3.5100 ;
      RECT 0.0000 2.4165 0.1170 3.5100 ;
      RECT 9.4590 2.4165 9.6120 3.3320 ;
      RECT 5.8950 2.4165 9.4410 3.5100 ;
      RECT 5.1480 2.4165 5.8770 3.3320 ;
      RECT 4.9860 2.6120 5.1120 3.5100 ;
      RECT 3.7350 2.5160 4.9590 3.3320 ;
      RECT 0.1710 2.4165 3.7170 3.5100 ;
      RECT 0.0000 2.4165 0.1530 3.3320 ;
      RECT 5.0940 2.4165 9.6120 3.2360 ;
      RECT 0.0000 2.5160 5.0760 3.2360 ;
      RECT 4.8690 2.4165 9.6120 2.5880 ;
      RECT 0.0000 2.4165 4.8510 3.2360 ;
      RECT 0.0000 2.4165 9.6120 2.4920 ;
      RECT 0.0000 4.4600 9.6120 4.5900 ;
      RECT 9.4950 3.4965 9.6120 4.5900 ;
      RECT 5.8410 4.3640 9.4770 4.5900 ;
      RECT 4.5090 4.3640 5.8230 4.5900 ;
      RECT 3.7890 3.4965 4.4190 4.5900 ;
      RECT 0.1350 4.3640 3.7710 4.5900 ;
      RECT 0.0000 3.4965 0.1170 4.5900 ;
      RECT 9.4590 3.4965 9.6120 4.4120 ;
      RECT 5.8950 3.4965 9.4410 4.5900 ;
      RECT 5.1480 3.4965 5.8770 4.4120 ;
      RECT 4.9860 3.6920 5.1120 4.5900 ;
      RECT 3.7350 3.5960 4.9590 4.4120 ;
      RECT 0.1710 3.4965 3.7170 4.5900 ;
      RECT 0.0000 3.4965 0.1530 4.4120 ;
      RECT 5.0940 3.4965 9.6120 4.3160 ;
      RECT 0.0000 3.5960 5.0760 4.3160 ;
      RECT 4.8690 3.4965 9.6120 3.6680 ;
      RECT 0.0000 3.4965 4.8510 4.3160 ;
      RECT 0.0000 3.4965 9.6120 3.5720 ;
      RECT 0.0000 5.5400 9.6120 5.6700 ;
      RECT 9.4950 4.5765 9.6120 5.6700 ;
      RECT 5.8410 5.4440 9.4770 5.6700 ;
      RECT 4.5090 5.4440 5.8230 5.6700 ;
      RECT 3.7890 4.5765 4.4190 5.6700 ;
      RECT 0.1350 5.4440 3.7710 5.6700 ;
      RECT 0.0000 4.5765 0.1170 5.6700 ;
      RECT 9.4590 4.5765 9.6120 5.4920 ;
      RECT 5.8950 4.5765 9.4410 5.6700 ;
      RECT 5.1480 4.5765 5.8770 5.4920 ;
      RECT 4.9860 4.7720 5.1120 5.6700 ;
      RECT 3.7350 4.6760 4.9590 5.4920 ;
      RECT 0.1710 4.5765 3.7170 5.6700 ;
      RECT 0.0000 4.5765 0.1530 5.4920 ;
      RECT 5.0940 4.5765 9.6120 5.3960 ;
      RECT 0.0000 4.6760 5.0760 5.3960 ;
      RECT 4.8690 4.5765 9.6120 4.7480 ;
      RECT 0.0000 4.5765 4.8510 5.3960 ;
      RECT 0.0000 4.5765 9.6120 4.6520 ;
      RECT 0.0000 6.6200 9.6120 6.7500 ;
      RECT 9.4950 5.6565 9.6120 6.7500 ;
      RECT 5.8410 6.5240 9.4770 6.7500 ;
      RECT 4.5090 6.5240 5.8230 6.7500 ;
      RECT 3.7890 5.6565 4.4190 6.7500 ;
      RECT 0.1350 6.5240 3.7710 6.7500 ;
      RECT 0.0000 5.6565 0.1170 6.7500 ;
      RECT 9.4590 5.6565 9.6120 6.5720 ;
      RECT 5.8950 5.6565 9.4410 6.7500 ;
      RECT 5.1480 5.6565 5.8770 6.5720 ;
      RECT 4.9860 5.8520 5.1120 6.7500 ;
      RECT 3.7350 5.7560 4.9590 6.5720 ;
      RECT 0.1710 5.6565 3.7170 6.7500 ;
      RECT 0.0000 5.6565 0.1530 6.5720 ;
      RECT 5.0940 5.6565 9.6120 6.4760 ;
      RECT 0.0000 5.7560 5.0760 6.4760 ;
      RECT 4.8690 5.6565 9.6120 5.8280 ;
      RECT 0.0000 5.6565 4.8510 6.4760 ;
      RECT 0.0000 5.6565 9.6120 5.7320 ;
      RECT 0.0000 7.7000 9.6120 7.8300 ;
      RECT 9.4950 6.7365 9.6120 7.8300 ;
      RECT 5.8410 7.6040 9.4770 7.8300 ;
      RECT 4.5090 7.6040 5.8230 7.8300 ;
      RECT 3.7890 6.7365 4.4190 7.8300 ;
      RECT 0.1350 7.6040 3.7710 7.8300 ;
      RECT 0.0000 6.7365 0.1170 7.8300 ;
      RECT 9.4590 6.7365 9.6120 7.6520 ;
      RECT 5.8950 6.7365 9.4410 7.8300 ;
      RECT 5.1480 6.7365 5.8770 7.6520 ;
      RECT 4.9860 6.9320 5.1120 7.8300 ;
      RECT 3.7350 6.8360 4.9590 7.6520 ;
      RECT 0.1710 6.7365 3.7170 7.8300 ;
      RECT 0.0000 6.7365 0.1530 7.6520 ;
      RECT 5.0940 6.7365 9.6120 7.5560 ;
      RECT 0.0000 6.8360 5.0760 7.5560 ;
      RECT 4.8690 6.7365 9.6120 6.9080 ;
      RECT 0.0000 6.7365 4.8510 7.5560 ;
      RECT 0.0000 6.7365 9.6120 6.8120 ;
      RECT 0.0000 8.7800 9.6120 8.9100 ;
      RECT 9.4950 7.8165 9.6120 8.9100 ;
      RECT 5.8410 8.6840 9.4770 8.9100 ;
      RECT 4.5090 8.6840 5.8230 8.9100 ;
      RECT 3.7890 7.8165 4.4190 8.9100 ;
      RECT 0.1350 8.6840 3.7710 8.9100 ;
      RECT 0.0000 7.8165 0.1170 8.9100 ;
      RECT 9.4590 7.8165 9.6120 8.7320 ;
      RECT 5.8950 7.8165 9.4410 8.9100 ;
      RECT 5.1480 7.8165 5.8770 8.7320 ;
      RECT 4.9860 8.0120 5.1120 8.9100 ;
      RECT 3.7350 7.9160 4.9590 8.7320 ;
      RECT 0.1710 7.8165 3.7170 8.9100 ;
      RECT 0.0000 7.8165 0.1530 8.7320 ;
      RECT 5.0940 7.8165 9.6120 8.6360 ;
      RECT 0.0000 7.9160 5.0760 8.6360 ;
      RECT 4.8690 7.8165 9.6120 7.9880 ;
      RECT 0.0000 7.8165 4.8510 8.6360 ;
      RECT 0.0000 7.8165 9.6120 7.8920 ;
      RECT 0.0000 9.8600 9.6120 9.9900 ;
      RECT 9.4950 8.8965 9.6120 9.9900 ;
      RECT 5.8410 9.7640 9.4770 9.9900 ;
      RECT 4.5090 9.7640 5.8230 9.9900 ;
      RECT 3.7890 8.8965 4.4190 9.9900 ;
      RECT 0.1350 9.7640 3.7710 9.9900 ;
      RECT 0.0000 8.8965 0.1170 9.9900 ;
      RECT 9.4590 8.8965 9.6120 9.8120 ;
      RECT 5.8950 8.8965 9.4410 9.9900 ;
      RECT 5.1480 8.8965 5.8770 9.8120 ;
      RECT 4.9860 9.0920 5.1120 9.9900 ;
      RECT 3.7350 8.9960 4.9590 9.8120 ;
      RECT 0.1710 8.8965 3.7170 9.9900 ;
      RECT 0.0000 8.8965 0.1530 9.8120 ;
      RECT 5.0940 8.8965 9.6120 9.7160 ;
      RECT 0.0000 8.9960 5.0760 9.7160 ;
      RECT 4.8690 8.8965 9.6120 9.0680 ;
      RECT 0.0000 8.8965 4.8510 9.7160 ;
      RECT 0.0000 8.8965 9.6120 8.9720 ;
      RECT 0.0000 10.9400 9.6120 11.0700 ;
      RECT 9.4950 9.9765 9.6120 11.0700 ;
      RECT 5.8410 10.8440 9.4770 11.0700 ;
      RECT 4.5090 10.8440 5.8230 11.0700 ;
      RECT 3.7890 9.9765 4.4190 11.0700 ;
      RECT 0.1350 10.8440 3.7710 11.0700 ;
      RECT 0.0000 9.9765 0.1170 11.0700 ;
      RECT 9.4590 9.9765 9.6120 10.8920 ;
      RECT 5.8950 9.9765 9.4410 11.0700 ;
      RECT 5.1480 9.9765 5.8770 10.8920 ;
      RECT 4.9860 10.1720 5.1120 11.0700 ;
      RECT 3.7350 10.0760 4.9590 10.8920 ;
      RECT 0.1710 9.9765 3.7170 11.0700 ;
      RECT 0.0000 9.9765 0.1530 10.8920 ;
      RECT 5.0940 9.9765 9.6120 10.7960 ;
      RECT 0.0000 10.0760 5.0760 10.7960 ;
      RECT 4.8690 9.9765 9.6120 10.1480 ;
      RECT 0.0000 9.9765 4.8510 10.7960 ;
      RECT 0.0000 9.9765 9.6120 10.0520 ;
      RECT 0.0000 12.0200 9.6120 12.1500 ;
      RECT 9.4950 11.0565 9.6120 12.1500 ;
      RECT 5.8410 11.9240 9.4770 12.1500 ;
      RECT 4.5090 11.9240 5.8230 12.1500 ;
      RECT 3.7890 11.0565 4.4190 12.1500 ;
      RECT 0.1350 11.9240 3.7710 12.1500 ;
      RECT 0.0000 11.0565 0.1170 12.1500 ;
      RECT 9.4590 11.0565 9.6120 11.9720 ;
      RECT 5.8950 11.0565 9.4410 12.1500 ;
      RECT 5.1480 11.0565 5.8770 11.9720 ;
      RECT 4.9860 11.2520 5.1120 12.1500 ;
      RECT 3.7350 11.1560 4.9590 11.9720 ;
      RECT 0.1710 11.0565 3.7170 12.1500 ;
      RECT 0.0000 11.0565 0.1530 11.9720 ;
      RECT 5.0940 11.0565 9.6120 11.8760 ;
      RECT 0.0000 11.1560 5.0760 11.8760 ;
      RECT 4.8690 11.0565 9.6120 11.2280 ;
      RECT 0.0000 11.0565 4.8510 11.8760 ;
      RECT 0.0000 11.0565 9.6120 11.1320 ;
      RECT 0.0000 13.1000 9.6120 13.2300 ;
      RECT 9.4950 12.1365 9.6120 13.2300 ;
      RECT 5.8410 13.0040 9.4770 13.2300 ;
      RECT 4.5090 13.0040 5.8230 13.2300 ;
      RECT 3.7890 12.1365 4.4190 13.2300 ;
      RECT 0.1350 13.0040 3.7710 13.2300 ;
      RECT 0.0000 12.1365 0.1170 13.2300 ;
      RECT 9.4590 12.1365 9.6120 13.0520 ;
      RECT 5.8950 12.1365 9.4410 13.2300 ;
      RECT 5.1480 12.1365 5.8770 13.0520 ;
      RECT 4.9860 12.3320 5.1120 13.2300 ;
      RECT 3.7350 12.2360 4.9590 13.0520 ;
      RECT 0.1710 12.1365 3.7170 13.2300 ;
      RECT 0.0000 12.1365 0.1530 13.0520 ;
      RECT 5.0940 12.1365 9.6120 12.9560 ;
      RECT 0.0000 12.2360 5.0760 12.9560 ;
      RECT 4.8690 12.1365 9.6120 12.3080 ;
      RECT 0.0000 12.1365 4.8510 12.9560 ;
      RECT 0.0000 12.1365 9.6120 12.2120 ;
      RECT 0.0000 14.1800 9.6120 14.3100 ;
      RECT 9.4950 13.2165 9.6120 14.3100 ;
      RECT 5.8410 14.0840 9.4770 14.3100 ;
      RECT 4.5090 14.0840 5.8230 14.3100 ;
      RECT 3.7890 13.2165 4.4190 14.3100 ;
      RECT 0.1350 14.0840 3.7710 14.3100 ;
      RECT 0.0000 13.2165 0.1170 14.3100 ;
      RECT 9.4590 13.2165 9.6120 14.1320 ;
      RECT 5.8950 13.2165 9.4410 14.3100 ;
      RECT 5.1480 13.2165 5.8770 14.1320 ;
      RECT 4.9860 13.4120 5.1120 14.3100 ;
      RECT 3.7350 13.3160 4.9590 14.1320 ;
      RECT 0.1710 13.2165 3.7170 14.3100 ;
      RECT 0.0000 13.2165 0.1530 14.1320 ;
      RECT 5.0940 13.2165 9.6120 14.0360 ;
      RECT 0.0000 13.3160 5.0760 14.0360 ;
      RECT 4.8690 13.2165 9.6120 13.3880 ;
      RECT 0.0000 13.2165 4.8510 14.0360 ;
      RECT 0.0000 13.2165 9.6120 13.2920 ;
      RECT 0.0000 15.2600 9.6120 15.3900 ;
      RECT 9.4950 14.2965 9.6120 15.3900 ;
      RECT 5.8410 15.1640 9.4770 15.3900 ;
      RECT 4.5090 15.1640 5.8230 15.3900 ;
      RECT 3.7890 14.2965 4.4190 15.3900 ;
      RECT 0.1350 15.1640 3.7710 15.3900 ;
      RECT 0.0000 14.2965 0.1170 15.3900 ;
      RECT 9.4590 14.2965 9.6120 15.2120 ;
      RECT 5.8950 14.2965 9.4410 15.3900 ;
      RECT 5.1480 14.2965 5.8770 15.2120 ;
      RECT 4.9860 14.4920 5.1120 15.3900 ;
      RECT 3.7350 14.3960 4.9590 15.2120 ;
      RECT 0.1710 14.2965 3.7170 15.3900 ;
      RECT 0.0000 14.2965 0.1530 15.2120 ;
      RECT 5.0940 14.2965 9.6120 15.1160 ;
      RECT 0.0000 14.3960 5.0760 15.1160 ;
      RECT 4.8690 14.2965 9.6120 14.4680 ;
      RECT 0.0000 14.2965 4.8510 15.1160 ;
      RECT 0.0000 14.2965 9.6120 14.3720 ;
      RECT 0.0000 16.3400 9.6120 16.4700 ;
      RECT 9.4950 15.3765 9.6120 16.4700 ;
      RECT 5.8410 16.2440 9.4770 16.4700 ;
      RECT 4.5090 16.2440 5.8230 16.4700 ;
      RECT 3.7890 15.3765 4.4190 16.4700 ;
      RECT 0.1350 16.2440 3.7710 16.4700 ;
      RECT 0.0000 15.3765 0.1170 16.4700 ;
      RECT 9.4590 15.3765 9.6120 16.2920 ;
      RECT 5.8950 15.3765 9.4410 16.4700 ;
      RECT 5.1480 15.3765 5.8770 16.2920 ;
      RECT 4.9860 15.5720 5.1120 16.4700 ;
      RECT 3.7350 15.4760 4.9590 16.2920 ;
      RECT 0.1710 15.3765 3.7170 16.4700 ;
      RECT 0.0000 15.3765 0.1530 16.2920 ;
      RECT 5.0940 15.3765 9.6120 16.1960 ;
      RECT 0.0000 15.4760 5.0760 16.1960 ;
      RECT 4.8690 15.3765 9.6120 15.5480 ;
      RECT 0.0000 15.3765 4.8510 16.1960 ;
      RECT 0.0000 15.3765 9.6120 15.4520 ;
      RECT 0.0000 17.4200 9.6120 17.5500 ;
      RECT 9.4950 16.4565 9.6120 17.5500 ;
      RECT 5.8410 17.3240 9.4770 17.5500 ;
      RECT 4.5090 17.3240 5.8230 17.5500 ;
      RECT 3.7890 16.4565 4.4190 17.5500 ;
      RECT 0.1350 17.3240 3.7710 17.5500 ;
      RECT 0.0000 16.4565 0.1170 17.5500 ;
      RECT 9.4590 16.4565 9.6120 17.3720 ;
      RECT 5.8950 16.4565 9.4410 17.5500 ;
      RECT 5.1480 16.4565 5.8770 17.3720 ;
      RECT 4.9860 16.6520 5.1120 17.5500 ;
      RECT 3.7350 16.5560 4.9590 17.3720 ;
      RECT 0.1710 16.4565 3.7170 17.5500 ;
      RECT 0.0000 16.4565 0.1530 17.3720 ;
      RECT 5.0940 16.4565 9.6120 17.2760 ;
      RECT 0.0000 16.5560 5.0760 17.2760 ;
      RECT 4.8690 16.4565 9.6120 16.6280 ;
      RECT 0.0000 16.4565 4.8510 17.2760 ;
      RECT 0.0000 16.4565 9.6120 16.5320 ;
      RECT 0.0000 24.8430 9.6120 26.1765 ;
      RECT 7.3530 17.5230 9.6120 26.1765 ;
      RECT 5.1530 21.3870 9.6120 26.1765 ;
      RECT 6.0570 18.7950 9.6120 26.1765 ;
      RECT 5.1010 17.5230 5.1350 26.1765 ;
      RECT 5.0490 17.5230 5.0830 26.1765 ;
      RECT 4.9970 17.5230 5.0310 26.1765 ;
      RECT 4.9450 17.5230 4.9790 26.1765 ;
      RECT 0.0000 24.4110 4.9270 26.1765 ;
      RECT 4.6850 21.6750 9.6120 24.6270 ;
      RECT 4.6330 17.5230 4.6670 26.1765 ;
      RECT 4.5810 17.5230 4.6150 26.1765 ;
      RECT 4.5290 17.5230 4.5630 26.1765 ;
      RECT 4.4770 17.5230 4.5110 26.1765 ;
      RECT 0.0000 19.0830 4.4590 26.1765 ;
      RECT 0.0000 21.2430 4.9270 24.1950 ;
      RECT 4.6850 18.5070 5.8230 21.4590 ;
      RECT 5.8410 18.9870 9.6120 26.1765 ;
      RECT 5.1930 17.6030 6.0390 21.3630 ;
      RECT 4.0050 18.0750 4.7790 21.0270 ;
      RECT 3.7890 18.2190 4.4590 26.1765 ;
      RECT 0.0000 18.7950 3.7710 26.1765 ;
      RECT 3.3570 17.5230 3.8070 19.0590 ;
      RECT 7.1370 17.5230 7.3350 26.1765 ;
      RECT 3.3570 18.6030 7.1190 18.9630 ;
      RECT 2.4930 18.2190 3.3390 26.1765 ;
      RECT 0.0000 18.5070 2.4750 26.1765 ;
      RECT 6.9210 17.5230 9.6120 18.7710 ;
      RECT 6.7050 18.2190 9.6120 18.7710 ;
      RECT 0.0000 18.5070 6.6870 18.7710 ;
      RECT 6.4890 17.5230 6.9030 18.5790 ;
      RECT 5.1530 18.2190 9.6120 18.5790 ;
      RECT 0.1710 18.2190 4.9270 18.7710 ;
      RECT 4.6850 18.1710 4.9270 26.1765 ;
      RECT 0.0000 18.0750 0.1530 26.1765 ;
      RECT 4.7970 17.5230 5.1750 18.2910 ;
      RECT 5.1930 18.1710 6.4710 18.9630 ;
      RECT 3.1410 18.1710 3.9870 18.7710 ;
      RECT 2.7090 18.1710 3.1230 26.1765 ;
      RECT 0.0000 18.0750 2.6910 18.2910 ;
      RECT 6.2730 17.5230 9.6120 18.1950 ;
      RECT 4.7970 17.6030 6.2550 18.1950 ;
      RECT 3.8250 18.0750 4.7790 18.1950 ;
      RECT 2.9250 17.5230 3.8070 18.1950 ;
      RECT 0.0000 18.0750 2.9070 18.1950 ;
      RECT 5.8410 17.5230 9.6120 18.1470 ;
      RECT 4.6850 17.6030 9.6120 18.1470 ;
      RECT 0.1350 17.5230 4.4590 18.1470 ;
      RECT 0.0000 17.5230 0.1170 26.1765 ;
      RECT 0.0000 17.5230 5.8230 17.8590 ;
      RECT 0.0000 17.5230 9.6120 17.5790 ;
        RECT 0.0000 26.6270 9.6120 26.7570 ;
        RECT 9.4950 25.6635 9.6120 26.7570 ;
        RECT 5.8410 26.5310 9.4770 26.7570 ;
        RECT 4.5090 26.5310 5.8230 26.7570 ;
        RECT 3.7890 25.6635 4.4190 26.7570 ;
        RECT 0.1350 26.5310 3.7710 26.7570 ;
        RECT 0.0000 25.6635 0.1170 26.7570 ;
        RECT 9.4590 25.6635 9.6120 26.5790 ;
        RECT 5.8950 25.6635 9.4410 26.7570 ;
        RECT 5.1480 25.6635 5.8770 26.5790 ;
        RECT 4.9860 25.8590 5.1120 26.7570 ;
        RECT 3.7350 25.7630 4.9590 26.5790 ;
        RECT 0.1710 25.6635 3.7170 26.7570 ;
        RECT 0.0000 25.6635 0.1530 26.5790 ;
        RECT 5.0940 25.6635 9.6120 26.4830 ;
        RECT 0.0000 25.7630 5.0760 26.4830 ;
        RECT 4.8690 25.6635 9.6120 25.8350 ;
        RECT 0.0000 25.6635 4.8510 26.4830 ;
        RECT 0.0000 25.6635 9.6120 25.7390 ;
        RECT 0.0000 27.7070 9.6120 27.8370 ;
        RECT 9.4950 26.7435 9.6120 27.8370 ;
        RECT 5.8410 27.6110 9.4770 27.8370 ;
        RECT 4.5090 27.6110 5.8230 27.8370 ;
        RECT 3.7890 26.7435 4.4190 27.8370 ;
        RECT 0.1350 27.6110 3.7710 27.8370 ;
        RECT 0.0000 26.7435 0.1170 27.8370 ;
        RECT 9.4590 26.7435 9.6120 27.6590 ;
        RECT 5.8950 26.7435 9.4410 27.8370 ;
        RECT 5.1480 26.7435 5.8770 27.6590 ;
        RECT 4.9860 26.9390 5.1120 27.8370 ;
        RECT 3.7350 26.8430 4.9590 27.6590 ;
        RECT 0.1710 26.7435 3.7170 27.8370 ;
        RECT 0.0000 26.7435 0.1530 27.6590 ;
        RECT 5.0940 26.7435 9.6120 27.5630 ;
        RECT 0.0000 26.8430 5.0760 27.5630 ;
        RECT 4.8690 26.7435 9.6120 26.9150 ;
        RECT 0.0000 26.7435 4.8510 27.5630 ;
        RECT 0.0000 26.7435 9.6120 26.8190 ;
        RECT 0.0000 28.7870 9.6120 28.9170 ;
        RECT 9.4950 27.8235 9.6120 28.9170 ;
        RECT 5.8410 28.6910 9.4770 28.9170 ;
        RECT 4.5090 28.6910 5.8230 28.9170 ;
        RECT 3.7890 27.8235 4.4190 28.9170 ;
        RECT 0.1350 28.6910 3.7710 28.9170 ;
        RECT 0.0000 27.8235 0.1170 28.9170 ;
        RECT 9.4590 27.8235 9.6120 28.7390 ;
        RECT 5.8950 27.8235 9.4410 28.9170 ;
        RECT 5.1480 27.8235 5.8770 28.7390 ;
        RECT 4.9860 28.0190 5.1120 28.9170 ;
        RECT 3.7350 27.9230 4.9590 28.7390 ;
        RECT 0.1710 27.8235 3.7170 28.9170 ;
        RECT 0.0000 27.8235 0.1530 28.7390 ;
        RECT 5.0940 27.8235 9.6120 28.6430 ;
        RECT 0.0000 27.9230 5.0760 28.6430 ;
        RECT 4.8690 27.8235 9.6120 27.9950 ;
        RECT 0.0000 27.8235 4.8510 28.6430 ;
        RECT 0.0000 27.8235 9.6120 27.8990 ;
        RECT 0.0000 29.8670 9.6120 29.9970 ;
        RECT 9.4950 28.9035 9.6120 29.9970 ;
        RECT 5.8410 29.7710 9.4770 29.9970 ;
        RECT 4.5090 29.7710 5.8230 29.9970 ;
        RECT 3.7890 28.9035 4.4190 29.9970 ;
        RECT 0.1350 29.7710 3.7710 29.9970 ;
        RECT 0.0000 28.9035 0.1170 29.9970 ;
        RECT 9.4590 28.9035 9.6120 29.8190 ;
        RECT 5.8950 28.9035 9.4410 29.9970 ;
        RECT 5.1480 28.9035 5.8770 29.8190 ;
        RECT 4.9860 29.0990 5.1120 29.9970 ;
        RECT 3.7350 29.0030 4.9590 29.8190 ;
        RECT 0.1710 28.9035 3.7170 29.9970 ;
        RECT 0.0000 28.9035 0.1530 29.8190 ;
        RECT 5.0940 28.9035 9.6120 29.7230 ;
        RECT 0.0000 29.0030 5.0760 29.7230 ;
        RECT 4.8690 28.9035 9.6120 29.0750 ;
        RECT 0.0000 28.9035 4.8510 29.7230 ;
        RECT 0.0000 28.9035 9.6120 28.9790 ;
        RECT 0.0000 30.9470 9.6120 31.0770 ;
        RECT 9.4950 29.9835 9.6120 31.0770 ;
        RECT 5.8410 30.8510 9.4770 31.0770 ;
        RECT 4.5090 30.8510 5.8230 31.0770 ;
        RECT 3.7890 29.9835 4.4190 31.0770 ;
        RECT 0.1350 30.8510 3.7710 31.0770 ;
        RECT 0.0000 29.9835 0.1170 31.0770 ;
        RECT 9.4590 29.9835 9.6120 30.8990 ;
        RECT 5.8950 29.9835 9.4410 31.0770 ;
        RECT 5.1480 29.9835 5.8770 30.8990 ;
        RECT 4.9860 30.1790 5.1120 31.0770 ;
        RECT 3.7350 30.0830 4.9590 30.8990 ;
        RECT 0.1710 29.9835 3.7170 31.0770 ;
        RECT 0.0000 29.9835 0.1530 30.8990 ;
        RECT 5.0940 29.9835 9.6120 30.8030 ;
        RECT 0.0000 30.0830 5.0760 30.8030 ;
        RECT 4.8690 29.9835 9.6120 30.1550 ;
        RECT 0.0000 29.9835 4.8510 30.8030 ;
        RECT 0.0000 29.9835 9.6120 30.0590 ;
        RECT 0.0000 32.0270 9.6120 32.1570 ;
        RECT 9.4950 31.0635 9.6120 32.1570 ;
        RECT 5.8410 31.9310 9.4770 32.1570 ;
        RECT 4.5090 31.9310 5.8230 32.1570 ;
        RECT 3.7890 31.0635 4.4190 32.1570 ;
        RECT 0.1350 31.9310 3.7710 32.1570 ;
        RECT 0.0000 31.0635 0.1170 32.1570 ;
        RECT 9.4590 31.0635 9.6120 31.9790 ;
        RECT 5.8950 31.0635 9.4410 32.1570 ;
        RECT 5.1480 31.0635 5.8770 31.9790 ;
        RECT 4.9860 31.2590 5.1120 32.1570 ;
        RECT 3.7350 31.1630 4.9590 31.9790 ;
        RECT 0.1710 31.0635 3.7170 32.1570 ;
        RECT 0.0000 31.0635 0.1530 31.9790 ;
        RECT 5.0940 31.0635 9.6120 31.8830 ;
        RECT 0.0000 31.1630 5.0760 31.8830 ;
        RECT 4.8690 31.0635 9.6120 31.2350 ;
        RECT 0.0000 31.0635 4.8510 31.8830 ;
        RECT 0.0000 31.0635 9.6120 31.1390 ;
        RECT 0.0000 33.1070 9.6120 33.2370 ;
        RECT 9.4950 32.1435 9.6120 33.2370 ;
        RECT 5.8410 33.0110 9.4770 33.2370 ;
        RECT 4.5090 33.0110 5.8230 33.2370 ;
        RECT 3.7890 32.1435 4.4190 33.2370 ;
        RECT 0.1350 33.0110 3.7710 33.2370 ;
        RECT 0.0000 32.1435 0.1170 33.2370 ;
        RECT 9.4590 32.1435 9.6120 33.0590 ;
        RECT 5.8950 32.1435 9.4410 33.2370 ;
        RECT 5.1480 32.1435 5.8770 33.0590 ;
        RECT 4.9860 32.3390 5.1120 33.2370 ;
        RECT 3.7350 32.2430 4.9590 33.0590 ;
        RECT 0.1710 32.1435 3.7170 33.2370 ;
        RECT 0.0000 32.1435 0.1530 33.0590 ;
        RECT 5.0940 32.1435 9.6120 32.9630 ;
        RECT 0.0000 32.2430 5.0760 32.9630 ;
        RECT 4.8690 32.1435 9.6120 32.3150 ;
        RECT 0.0000 32.1435 4.8510 32.9630 ;
        RECT 0.0000 32.1435 9.6120 32.2190 ;
        RECT 0.0000 34.1870 9.6120 34.3170 ;
        RECT 9.4950 33.2235 9.6120 34.3170 ;
        RECT 5.8410 34.0910 9.4770 34.3170 ;
        RECT 4.5090 34.0910 5.8230 34.3170 ;
        RECT 3.7890 33.2235 4.4190 34.3170 ;
        RECT 0.1350 34.0910 3.7710 34.3170 ;
        RECT 0.0000 33.2235 0.1170 34.3170 ;
        RECT 9.4590 33.2235 9.6120 34.1390 ;
        RECT 5.8950 33.2235 9.4410 34.3170 ;
        RECT 5.1480 33.2235 5.8770 34.1390 ;
        RECT 4.9860 33.4190 5.1120 34.3170 ;
        RECT 3.7350 33.3230 4.9590 34.1390 ;
        RECT 0.1710 33.2235 3.7170 34.3170 ;
        RECT 0.0000 33.2235 0.1530 34.1390 ;
        RECT 5.0940 33.2235 9.6120 34.0430 ;
        RECT 0.0000 33.3230 5.0760 34.0430 ;
        RECT 4.8690 33.2235 9.6120 33.3950 ;
        RECT 0.0000 33.2235 4.8510 34.0430 ;
        RECT 0.0000 33.2235 9.6120 33.2990 ;
        RECT 0.0000 35.2670 9.6120 35.3970 ;
        RECT 9.4950 34.3035 9.6120 35.3970 ;
        RECT 5.8410 35.1710 9.4770 35.3970 ;
        RECT 4.5090 35.1710 5.8230 35.3970 ;
        RECT 3.7890 34.3035 4.4190 35.3970 ;
        RECT 0.1350 35.1710 3.7710 35.3970 ;
        RECT 0.0000 34.3035 0.1170 35.3970 ;
        RECT 9.4590 34.3035 9.6120 35.2190 ;
        RECT 5.8950 34.3035 9.4410 35.3970 ;
        RECT 5.1480 34.3035 5.8770 35.2190 ;
        RECT 4.9860 34.4990 5.1120 35.3970 ;
        RECT 3.7350 34.4030 4.9590 35.2190 ;
        RECT 0.1710 34.3035 3.7170 35.3970 ;
        RECT 0.0000 34.3035 0.1530 35.2190 ;
        RECT 5.0940 34.3035 9.6120 35.1230 ;
        RECT 0.0000 34.4030 5.0760 35.1230 ;
        RECT 4.8690 34.3035 9.6120 34.4750 ;
        RECT 0.0000 34.3035 4.8510 35.1230 ;
        RECT 0.0000 34.3035 9.6120 34.3790 ;
        RECT 0.0000 36.3470 9.6120 36.4770 ;
        RECT 9.4950 35.3835 9.6120 36.4770 ;
        RECT 5.8410 36.2510 9.4770 36.4770 ;
        RECT 4.5090 36.2510 5.8230 36.4770 ;
        RECT 3.7890 35.3835 4.4190 36.4770 ;
        RECT 0.1350 36.2510 3.7710 36.4770 ;
        RECT 0.0000 35.3835 0.1170 36.4770 ;
        RECT 9.4590 35.3835 9.6120 36.2990 ;
        RECT 5.8950 35.3835 9.4410 36.4770 ;
        RECT 5.1480 35.3835 5.8770 36.2990 ;
        RECT 4.9860 35.5790 5.1120 36.4770 ;
        RECT 3.7350 35.4830 4.9590 36.2990 ;
        RECT 0.1710 35.3835 3.7170 36.4770 ;
        RECT 0.0000 35.3835 0.1530 36.2990 ;
        RECT 5.0940 35.3835 9.6120 36.2030 ;
        RECT 0.0000 35.4830 5.0760 36.2030 ;
        RECT 4.8690 35.3835 9.6120 35.5550 ;
        RECT 0.0000 35.3835 4.8510 36.2030 ;
        RECT 0.0000 35.3835 9.6120 35.4590 ;
        RECT 0.0000 37.4270 9.6120 37.5570 ;
        RECT 9.4950 36.4635 9.6120 37.5570 ;
        RECT 5.8410 37.3310 9.4770 37.5570 ;
        RECT 4.5090 37.3310 5.8230 37.5570 ;
        RECT 3.7890 36.4635 4.4190 37.5570 ;
        RECT 0.1350 37.3310 3.7710 37.5570 ;
        RECT 0.0000 36.4635 0.1170 37.5570 ;
        RECT 9.4590 36.4635 9.6120 37.3790 ;
        RECT 5.8950 36.4635 9.4410 37.5570 ;
        RECT 5.1480 36.4635 5.8770 37.3790 ;
        RECT 4.9860 36.6590 5.1120 37.5570 ;
        RECT 3.7350 36.5630 4.9590 37.3790 ;
        RECT 0.1710 36.4635 3.7170 37.5570 ;
        RECT 0.0000 36.4635 0.1530 37.3790 ;
        RECT 5.0940 36.4635 9.6120 37.2830 ;
        RECT 0.0000 36.5630 5.0760 37.2830 ;
        RECT 4.8690 36.4635 9.6120 36.6350 ;
        RECT 0.0000 36.4635 4.8510 37.2830 ;
        RECT 0.0000 36.4635 9.6120 36.5390 ;
        RECT 0.0000 38.5070 9.6120 38.6370 ;
        RECT 9.4950 37.5435 9.6120 38.6370 ;
        RECT 5.8410 38.4110 9.4770 38.6370 ;
        RECT 4.5090 38.4110 5.8230 38.6370 ;
        RECT 3.7890 37.5435 4.4190 38.6370 ;
        RECT 0.1350 38.4110 3.7710 38.6370 ;
        RECT 0.0000 37.5435 0.1170 38.6370 ;
        RECT 9.4590 37.5435 9.6120 38.4590 ;
        RECT 5.8950 37.5435 9.4410 38.6370 ;
        RECT 5.1480 37.5435 5.8770 38.4590 ;
        RECT 4.9860 37.7390 5.1120 38.6370 ;
        RECT 3.7350 37.6430 4.9590 38.4590 ;
        RECT 0.1710 37.5435 3.7170 38.6370 ;
        RECT 0.0000 37.5435 0.1530 38.4590 ;
        RECT 5.0940 37.5435 9.6120 38.3630 ;
        RECT 0.0000 37.6430 5.0760 38.3630 ;
        RECT 4.8690 37.5435 9.6120 37.7150 ;
        RECT 0.0000 37.5435 4.8510 38.3630 ;
        RECT 0.0000 37.5435 9.6120 37.6190 ;
        RECT 0.0000 39.5870 9.6120 39.7170 ;
        RECT 9.4950 38.6235 9.6120 39.7170 ;
        RECT 5.8410 39.4910 9.4770 39.7170 ;
        RECT 4.5090 39.4910 5.8230 39.7170 ;
        RECT 3.7890 38.6235 4.4190 39.7170 ;
        RECT 0.1350 39.4910 3.7710 39.7170 ;
        RECT 0.0000 38.6235 0.1170 39.7170 ;
        RECT 9.4590 38.6235 9.6120 39.5390 ;
        RECT 5.8950 38.6235 9.4410 39.7170 ;
        RECT 5.1480 38.6235 5.8770 39.5390 ;
        RECT 4.9860 38.8190 5.1120 39.7170 ;
        RECT 3.7350 38.7230 4.9590 39.5390 ;
        RECT 0.1710 38.6235 3.7170 39.7170 ;
        RECT 0.0000 38.6235 0.1530 39.5390 ;
        RECT 5.0940 38.6235 9.6120 39.4430 ;
        RECT 0.0000 38.7230 5.0760 39.4430 ;
        RECT 4.8690 38.6235 9.6120 38.7950 ;
        RECT 0.0000 38.6235 4.8510 39.4430 ;
        RECT 0.0000 38.6235 9.6120 38.6990 ;
        RECT 0.0000 40.6670 9.6120 40.7970 ;
        RECT 9.4950 39.7035 9.6120 40.7970 ;
        RECT 5.8410 40.5710 9.4770 40.7970 ;
        RECT 4.5090 40.5710 5.8230 40.7970 ;
        RECT 3.7890 39.7035 4.4190 40.7970 ;
        RECT 0.1350 40.5710 3.7710 40.7970 ;
        RECT 0.0000 39.7035 0.1170 40.7970 ;
        RECT 9.4590 39.7035 9.6120 40.6190 ;
        RECT 5.8950 39.7035 9.4410 40.7970 ;
        RECT 5.1480 39.7035 5.8770 40.6190 ;
        RECT 4.9860 39.8990 5.1120 40.7970 ;
        RECT 3.7350 39.8030 4.9590 40.6190 ;
        RECT 0.1710 39.7035 3.7170 40.7970 ;
        RECT 0.0000 39.7035 0.1530 40.6190 ;
        RECT 5.0940 39.7035 9.6120 40.5230 ;
        RECT 0.0000 39.8030 5.0760 40.5230 ;
        RECT 4.8690 39.7035 9.6120 39.8750 ;
        RECT 0.0000 39.7035 4.8510 40.5230 ;
        RECT 0.0000 39.7035 9.6120 39.7790 ;
        RECT 0.0000 41.7470 9.6120 41.8770 ;
        RECT 9.4950 40.7835 9.6120 41.8770 ;
        RECT 5.8410 41.6510 9.4770 41.8770 ;
        RECT 4.5090 41.6510 5.8230 41.8770 ;
        RECT 3.7890 40.7835 4.4190 41.8770 ;
        RECT 0.1350 41.6510 3.7710 41.8770 ;
        RECT 0.0000 40.7835 0.1170 41.8770 ;
        RECT 9.4590 40.7835 9.6120 41.6990 ;
        RECT 5.8950 40.7835 9.4410 41.8770 ;
        RECT 5.1480 40.7835 5.8770 41.6990 ;
        RECT 4.9860 40.9790 5.1120 41.8770 ;
        RECT 3.7350 40.8830 4.9590 41.6990 ;
        RECT 0.1710 40.7835 3.7170 41.8770 ;
        RECT 0.0000 40.7835 0.1530 41.6990 ;
        RECT 5.0940 40.7835 9.6120 41.6030 ;
        RECT 0.0000 40.8830 5.0760 41.6030 ;
        RECT 4.8690 40.7835 9.6120 40.9550 ;
        RECT 0.0000 40.7835 4.8510 41.6030 ;
        RECT 0.0000 40.7835 9.6120 40.8590 ;
        RECT 0.0000 42.8270 9.6120 42.9570 ;
        RECT 9.4950 41.8635 9.6120 42.9570 ;
        RECT 5.8410 42.7310 9.4770 42.9570 ;
        RECT 4.5090 42.7310 5.8230 42.9570 ;
        RECT 3.7890 41.8635 4.4190 42.9570 ;
        RECT 0.1350 42.7310 3.7710 42.9570 ;
        RECT 0.0000 41.8635 0.1170 42.9570 ;
        RECT 9.4590 41.8635 9.6120 42.7790 ;
        RECT 5.8950 41.8635 9.4410 42.9570 ;
        RECT 5.1480 41.8635 5.8770 42.7790 ;
        RECT 4.9860 42.0590 5.1120 42.9570 ;
        RECT 3.7350 41.9630 4.9590 42.7790 ;
        RECT 0.1710 41.8635 3.7170 42.9570 ;
        RECT 0.0000 41.8635 0.1530 42.7790 ;
        RECT 5.0940 41.8635 9.6120 42.6830 ;
        RECT 0.0000 41.9630 5.0760 42.6830 ;
        RECT 4.8690 41.8635 9.6120 42.0350 ;
        RECT 0.0000 41.8635 4.8510 42.6830 ;
        RECT 0.0000 41.8635 9.6120 41.9390 ;
  LAYER M4  ;
      RECT 1.6070 19.2360 8.0025 19.2600 ;
      RECT 1.6070 19.5240 8.0025 19.5480 ;
      RECT 1.6070 19.9080 8.0025 19.9320 ;
      RECT 1.6070 20.0040 8.0025 20.0280 ;
      RECT 1.6070 20.3400 8.0025 20.3640 ;
      RECT 7.4990 18.1950 7.5830 18.2190 ;
      RECT 7.3190 18.6270 7.4360 18.6510 ;
      RECT 7.3190 19.2840 7.4360 19.3080 ;
      RECT 7.3190 19.5720 7.4360 19.5960 ;
      RECT 6.6785 18.6270 7.2480 18.6510 ;
      RECT 6.7430 19.4040 6.8510 19.4280 ;
      RECT 5.4070 19.7790 6.5000 19.8030 ;
      RECT 6.0950 19.3470 6.1790 19.3710 ;
      RECT 5.3110 20.5470 6.1790 20.5710 ;
      RECT 6.0950 20.6430 6.1790 20.6670 ;
      RECT 5.9170 18.8670 6.0010 18.8910 ;
      RECT 5.8790 20.2110 5.9630 20.2350 ;
      RECT 5.7010 18.7710 5.7850 18.7950 ;
      RECT 5.4870 17.4830 5.7500 17.5070 ;
      RECT 5.4870 26.1230 5.7500 26.1470 ;
      RECT 5.5030 20.2590 5.7470 20.2830 ;
      RECT 5.6630 20.4030 5.7470 20.4270 ;
      RECT 4.2070 20.6430 5.7470 20.6670 ;
      RECT 5.6630 20.9310 5.7470 20.9550 ;
      RECT 5.4290 26.0270 5.6920 26.0510 ;
      RECT 5.4280 17.3870 5.6910 17.4110 ;
      RECT 5.3900 17.2910 5.6530 17.3150 ;
      RECT 5.3900 25.8350 5.6530 25.8590 ;
      RECT 5.5550 21.3630 5.6390 21.3870 ;
      RECT 4.7830 21.7470 5.6390 21.7710 ;
      RECT 5.1670 24.0030 5.6390 24.0270 ;
      RECT 5.5550 24.0990 5.6390 24.1230 ;
      RECT 5.3420 17.1950 5.6050 17.2190 ;
      RECT 5.3420 25.7390 5.6050 25.7630 ;
      RECT 5.1190 23.0910 5.5640 23.1150 ;
      RECT 5.2980 17.0990 5.5610 17.1230 ;
      RECT 5.2980 26.0750 5.5610 26.0990 ;
      RECT 5.2490 17.4350 5.5120 17.4590 ;
      RECT 5.2490 25.9790 5.5120 26.0030 ;
      RECT 5.3800 20.4030 5.5010 20.4270 ;
      RECT 5.3590 22.5150 5.4920 22.5390 ;
      RECT 5.2020 17.3390 5.4650 17.3630 ;
      RECT 5.2020 25.8830 5.4650 25.9070 ;
      RECT 5.1670 17.0510 5.4300 17.0750 ;
      RECT 5.1670 25.7870 5.4300 25.8110 ;
      RECT 4.3510 24.0990 5.4200 24.1230 ;
      RECT 5.3360 25.2510 5.4200 25.2750 ;
      RECT 5.1110 16.9070 5.3740 16.9310 ;
      RECT 5.1110 25.6910 5.3740 25.7150 ;
      RECT 5.2630 21.3630 5.3480 21.3870 ;
      RECT 4.1590 21.9390 5.2760 21.9630 ;
      RECT 4.8040 19.7790 5.2610 19.8030 ;
      RECT 4.6310 17.6270 4.8980 17.6510 ;
      RECT 4.6310 25.5470 4.8980 25.5710 ;
      RECT 4.7680 21.3150 4.8770 21.3390 ;
      RECT 4.6080 17.5310 4.8500 17.5550 ;
      RECT 4.6080 26.1710 4.8500 26.1950 ;
      RECT 4.5520 17.0510 4.7940 17.0750 ;
      RECT 4.5810 26.2670 4.7940 26.2910 ;
      RECT 4.6970 20.9310 4.7810 20.9550 ;
      RECT 4.4980 17.1470 4.7460 17.1710 ;
      RECT 4.4980 26.1230 4.7460 26.1470 ;
      RECT 4.2640 23.5230 4.6850 23.5470 ;
      RECT 4.2320 17.4830 4.4990 17.5070 ;
      RECT 4.2320 26.2670 4.4990 26.2910 ;
      RECT 4.3720 22.0830 4.4930 22.1070 ;
      RECT 4.3640 25.2510 4.4480 25.2750 ;
      RECT 4.1980 17.3870 4.4450 17.4110 ;
      RECT 4.1310 25.8350 4.4450 25.8590 ;
      RECT 4.1720 17.2910 4.4020 17.3150 ;
      RECT 4.1600 26.1710 4.4020 26.1950 ;
      RECT 4.1190 17.1950 4.3490 17.2190 ;
      RECT 4.2650 23.6670 4.3490 23.6910 ;
      RECT 4.0690 25.7390 4.3490 25.7630 ;
      RECT 4.0740 17.0990 4.3040 17.1230 ;
      RECT 4.0740 26.0750 4.3040 26.0990 ;
      RECT 3.1120 20.9310 4.3010 20.9550 ;
      RECT 4.0360 17.3390 4.2660 17.3630 ;
      RECT 4.0360 25.9790 4.2660 26.0030 ;
      RECT 4.0180 17.2430 4.2110 17.2670 ;
      RECT 4.0180 25.8830 4.2110 25.9070 ;
      RECT 3.9690 17.1470 4.1620 17.1710 ;
      RECT 3.9690 25.7870 4.1620 25.8110 ;
      RECT 3.9730 21.8430 4.1570 21.8670 ;
      RECT 3.9170 17.0510 4.1100 17.0750 ;
      RECT 3.9170 25.6910 4.1100 25.7150 ;
      RECT 3.4330 19.1550 4.1090 19.1790 ;
      RECT 3.9730 21.9390 4.0570 21.9630 ;
      RECT 3.7040 17.5790 3.9670 17.6030 ;
      RECT 3.7580 21.3630 3.8700 21.3870 ;
      RECT 3.3950 19.3470 3.4790 19.3710 ;
  LAYER V4  ;
      RECT 7.5480 18.1950 7.5720 18.2190 ;
      RECT 7.5480 19.2360 7.5720 19.2600 ;
      RECT 7.3800 18.6270 7.4040 18.6510 ;
      RECT 7.3800 19.2840 7.4040 19.3080 ;
      RECT 7.3800 19.5720 7.4040 19.5960 ;
      RECT 6.7560 18.6270 6.7800 18.6510 ;
      RECT 6.7560 19.4040 6.7800 19.4280 ;
      RECT 6.1440 19.3470 6.1680 19.3710 ;
      RECT 6.1440 19.5240 6.1680 19.5480 ;
      RECT 6.1440 20.5470 6.1680 20.5710 ;
      RECT 6.1440 20.6430 6.1680 20.6670 ;
      RECT 5.9280 18.8670 5.9520 18.8910 ;
      RECT 5.9280 19.9080 5.9520 19.9320 ;
      RECT 5.9280 20.2110 5.9520 20.2350 ;
      RECT 5.9280 20.3400 5.9520 20.3640 ;
      RECT 5.7120 18.7710 5.7360 18.7950 ;
      RECT 5.7120 20.0040 5.7360 20.0280 ;
      RECT 5.7120 20.2590 5.7360 20.2830 ;
      RECT 5.7120 20.4030 5.7360 20.4270 ;
      RECT 5.7120 20.6430 5.7360 20.6670 ;
      RECT 5.7120 20.9310 5.7360 20.9550 ;
      RECT 5.6040 21.3630 5.6280 21.3870 ;
      RECT 5.6040 21.7470 5.6280 21.7710 ;
      RECT 5.6040 24.0030 5.6280 24.0270 ;
      RECT 5.6040 24.0990 5.6280 24.1230 ;
      RECT 5.5140 17.4830 5.5380 17.5070 ;
      RECT 5.5140 20.2590 5.5380 20.2830 ;
      RECT 5.5140 26.1230 5.5380 26.1470 ;
      RECT 5.4660 17.3870 5.4900 17.4110 ;
      RECT 5.4660 20.4030 5.4900 20.4270 ;
      RECT 5.4660 26.0270 5.4900 26.0510 ;
      RECT 5.4180 17.2910 5.4420 17.3150 ;
      RECT 5.4180 19.7790 5.4420 19.8030 ;
      RECT 5.4180 25.8350 5.4420 25.8590 ;
      RECT 5.3700 17.1950 5.3940 17.2190 ;
      RECT 5.3700 22.5150 5.3940 22.5390 ;
      RECT 5.3700 25.2510 5.3940 25.2750 ;
      RECT 5.3700 25.7390 5.3940 25.7630 ;
      RECT 5.3220 17.0990 5.3460 17.1230 ;
      RECT 5.3220 20.5470 5.3460 20.5710 ;
      RECT 5.3220 26.0750 5.3460 26.0990 ;
      RECT 5.2740 17.4350 5.2980 17.4590 ;
      RECT 5.2740 21.3630 5.2980 21.3870 ;
      RECT 5.2740 25.9790 5.2980 26.0030 ;
      RECT 5.2260 17.3390 5.2500 17.3630 ;
      RECT 5.2260 19.7790 5.2500 19.8030 ;
      RECT 5.2260 25.8830 5.2500 25.9070 ;
      RECT 5.1780 17.0510 5.2020 17.0750 ;
      RECT 5.1780 24.0030 5.2020 24.0270 ;
      RECT 5.1780 25.7870 5.2020 25.8110 ;
      RECT 5.1300 16.9070 5.1540 16.9310 ;
      RECT 5.1300 23.0910 5.1540 23.1150 ;
      RECT 5.1300 25.6910 5.1540 25.7150 ;
      RECT 4.8420 17.6270 4.8660 17.6510 ;
      RECT 4.8420 21.3150 4.8660 21.3390 ;
      RECT 4.8420 25.5470 4.8660 25.5710 ;
      RECT 4.7940 17.5310 4.8180 17.5550 ;
      RECT 4.7940 21.7470 4.8180 21.7710 ;
      RECT 4.7940 26.1710 4.8180 26.1950 ;
      RECT 4.7460 17.0510 4.7700 17.0750 ;
      RECT 4.7460 20.9310 4.7700 20.9550 ;
      RECT 4.7460 26.2670 4.7700 26.2910 ;
      RECT 4.6500 17.1470 4.6740 17.1710 ;
      RECT 4.6500 23.5230 4.6740 23.5470 ;
      RECT 4.6500 26.1230 4.6740 26.1470 ;
      RECT 4.4580 17.4830 4.4820 17.5070 ;
      RECT 4.4580 22.0830 4.4820 22.1070 ;
      RECT 4.4580 26.2670 4.4820 26.2910 ;
      RECT 4.4100 17.3870 4.4340 17.4110 ;
      RECT 4.4100 25.2510 4.4340 25.2750 ;
      RECT 4.4100 25.8350 4.4340 25.8590 ;
      RECT 4.3620 17.2910 4.3860 17.3150 ;
      RECT 4.3620 24.0990 4.3860 24.1230 ;
      RECT 4.3620 26.1710 4.3860 26.1950 ;
      RECT 4.3140 17.1950 4.3380 17.2190 ;
      RECT 4.3140 23.6670 4.3380 23.6910 ;
      RECT 4.3140 25.7390 4.3380 25.7630 ;
      RECT 4.2660 17.0990 4.2900 17.1230 ;
      RECT 4.2660 20.9310 4.2900 20.9550 ;
      RECT 4.2660 26.0750 4.2900 26.0990 ;
      RECT 4.2180 17.3390 4.2420 17.3630 ;
      RECT 4.2180 20.6430 4.2420 20.6670 ;
      RECT 4.2180 25.9790 4.2420 26.0030 ;
      RECT 4.1700 17.2430 4.1940 17.2670 ;
      RECT 4.1700 21.9390 4.1940 21.9630 ;
      RECT 4.1700 25.8830 4.1940 25.9070 ;
      RECT 4.1220 17.1470 4.1460 17.1710 ;
      RECT 4.1220 21.8430 4.1460 21.8670 ;
      RECT 4.1220 25.7870 4.1460 25.8110 ;
      RECT 4.0740 17.0510 4.0980 17.0750 ;
      RECT 4.0740 19.1550 4.0980 19.1790 ;
      RECT 4.0740 25.6910 4.0980 25.7150 ;
      RECT 3.9840 21.8430 4.0080 21.8670 ;
      RECT 3.9840 21.9390 4.0080 21.9630 ;
      RECT 3.8170 17.5790 3.8410 17.6030 ;
      RECT 3.8170 21.3630 3.8410 21.3870 ;
      RECT 3.4440 19.1550 3.4680 19.1790 ;
      RECT 3.4440 19.3470 3.4680 19.3710 ;
  LAYER M5  ;
      RECT 7.5480 18.1840 7.5720 19.2710 ;
      RECT 7.3800 18.6135 7.4040 19.6460 ;
      RECT 6.7560 18.6075 6.7800 19.4400 ;
      RECT 6.1440 19.3360 6.1680 19.5590 ;
      RECT 6.1440 20.5360 6.1680 20.6780 ;
      RECT 5.9280 18.8560 5.9520 19.9430 ;
      RECT 5.9280 20.2000 5.9520 20.3750 ;
      RECT 5.7120 18.7600 5.7360 20.0390 ;
      RECT 5.7120 20.2480 5.7360 20.4380 ;
      RECT 5.7120 20.6320 5.7360 20.9660 ;
      RECT 5.6040 21.3520 5.6280 21.7820 ;
      RECT 5.6040 23.9920 5.6280 24.1340 ;
      RECT 5.5140 17.8200 5.5380 25.4030 ;
      RECT 5.4660 17.8200 5.4900 25.4030 ;
      RECT 5.4180 17.8200 5.4420 25.4030 ;
      RECT 5.3700 17.8200 5.3940 25.4030 ;
      RECT 5.3220 17.8200 5.3460 25.4030 ;
      RECT 5.2740 17.8200 5.2980 25.4030 ;
      RECT 5.2260 17.8200 5.2500 25.4030 ;
      RECT 5.1780 17.8200 5.2020 25.4030 ;
      RECT 5.1300 17.8200 5.1540 25.4030 ;
      RECT 4.8420 17.5580 4.8660 25.5910 ;
      RECT 4.7940 17.0370 4.8180 26.3660 ;
      RECT 4.7460 17.0060 4.7700 26.3650 ;
      RECT 4.6500 17.0520 4.6740 26.3660 ;
      RECT 4.4580 17.0510 4.4820 26.3190 ;
      RECT 4.4100 17.0510 4.4340 26.3190 ;
      RECT 4.3620 17.0510 4.3860 26.3190 ;
      RECT 4.3140 17.0510 4.3380 26.3190 ;
      RECT 4.2660 17.0510 4.2900 26.3190 ;
      RECT 4.2180 17.0220 4.2420 26.3190 ;
      RECT 4.1700 16.9780 4.1940 26.3200 ;
      RECT 4.1220 16.9410 4.1460 26.3210 ;
      RECT 4.0740 16.8810 4.0980 26.3210 ;
      RECT 3.9840 21.8320 4.0080 21.9740 ;
      RECT 3.8170 17.5610 3.8410 21.4050 ;
      RECT 3.4440 19.1440 3.4680 19.3820 ;
  LAYER M2  ;
    RECT 0.108 0.036 9.5040 43.1640 ;
  LAYER M1  ;
    RECT 0.108 0.036 9.5040 43.1640 ;
  END
END srambank_64x4x32_6t122 
