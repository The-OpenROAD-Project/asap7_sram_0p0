VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_256x4x48_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_256x4x48_6t122 0 0 ; 
  SIZE 121.392 BY 241.92 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.416 4.688 121.032 4.88 ; 
        RECT 0.416 9.008 121.032 9.2 ; 
        RECT 0.416 13.328 121.032 13.52 ; 
        RECT 0.416 17.648 121.032 17.84 ; 
        RECT 0.416 21.968 121.032 22.16 ; 
        RECT 0.416 26.288 121.032 26.48 ; 
        RECT 0.416 30.608 121.032 30.8 ; 
        RECT 0.416 34.928 121.032 35.12 ; 
        RECT 0.416 39.248 121.032 39.44 ; 
        RECT 0.416 43.568 121.032 43.76 ; 
        RECT 0.416 47.888 121.032 48.08 ; 
        RECT 0.416 52.208 121.032 52.4 ; 
        RECT 0.416 56.528 121.032 56.72 ; 
        RECT 0.416 60.848 121.032 61.04 ; 
        RECT 0.416 65.168 121.032 65.36 ; 
        RECT 0.416 69.488 121.032 69.68 ; 
        RECT 0.416 73.808 121.032 74 ; 
        RECT 0.416 78.128 121.032 78.32 ; 
        RECT 0.416 82.448 121.032 82.64 ; 
        RECT 0.416 86.768 121.032 86.96 ; 
        RECT 0.416 91.088 121.032 91.28 ; 
        RECT 0.416 95.408 121.032 95.6 ; 
        RECT 0.416 99.728 121.032 99.92 ; 
        RECT 0.416 104.048 121.032 104.24 ; 
        RECT 0.416 140.876 121.032 141.068 ; 
        RECT 0.416 145.196 121.032 145.388 ; 
        RECT 0.416 149.516 121.032 149.708 ; 
        RECT 0.416 153.836 121.032 154.028 ; 
        RECT 0.416 158.156 121.032 158.348 ; 
        RECT 0.416 162.476 121.032 162.668 ; 
        RECT 0.416 166.796 121.032 166.988 ; 
        RECT 0.416 171.116 121.032 171.308 ; 
        RECT 0.416 175.436 121.032 175.628 ; 
        RECT 0.416 179.756 121.032 179.948 ; 
        RECT 0.416 184.076 121.032 184.268 ; 
        RECT 0.416 188.396 121.032 188.588 ; 
        RECT 0.416 192.716 121.032 192.908 ; 
        RECT 0.416 197.036 121.032 197.228 ; 
        RECT 0.416 201.356 121.032 201.548 ; 
        RECT 0.416 205.676 121.032 205.868 ; 
        RECT 0.416 209.996 121.032 210.188 ; 
        RECT 0.416 214.316 121.032 214.508 ; 
        RECT 0.416 218.636 121.032 218.828 ; 
        RECT 0.416 222.956 121.032 223.148 ; 
        RECT 0.416 227.276 121.032 227.468 ; 
        RECT 0.416 231.596 121.032 231.788 ; 
        RECT 0.416 235.916 121.032 236.108 ; 
        RECT 0.416 240.236 121.032 240.428 ; 
      LAYER M3 ; 
        RECT 120.872 0.866 120.944 5.506 ; 
        RECT 64.784 0.868 64.856 5.504 ; 
        RECT 59.168 1.012 59.528 5.474 ; 
        RECT 56.576 0.868 56.648 5.504 ; 
        RECT 0.488 0.866 0.56 5.506 ; 
        RECT 120.872 5.186 120.944 9.826 ; 
        RECT 64.784 5.188 64.856 9.824 ; 
        RECT 59.168 5.332 59.528 9.794 ; 
        RECT 56.576 5.188 56.648 9.824 ; 
        RECT 0.488 5.186 0.56 9.826 ; 
        RECT 120.872 9.506 120.944 14.146 ; 
        RECT 64.784 9.508 64.856 14.144 ; 
        RECT 59.168 9.652 59.528 14.114 ; 
        RECT 56.576 9.508 56.648 14.144 ; 
        RECT 0.488 9.506 0.56 14.146 ; 
        RECT 120.872 13.826 120.944 18.466 ; 
        RECT 64.784 13.828 64.856 18.464 ; 
        RECT 59.168 13.972 59.528 18.434 ; 
        RECT 56.576 13.828 56.648 18.464 ; 
        RECT 0.488 13.826 0.56 18.466 ; 
        RECT 120.872 18.146 120.944 22.786 ; 
        RECT 64.784 18.148 64.856 22.784 ; 
        RECT 59.168 18.292 59.528 22.754 ; 
        RECT 56.576 18.148 56.648 22.784 ; 
        RECT 0.488 18.146 0.56 22.786 ; 
        RECT 120.872 22.466 120.944 27.106 ; 
        RECT 64.784 22.468 64.856 27.104 ; 
        RECT 59.168 22.612 59.528 27.074 ; 
        RECT 56.576 22.468 56.648 27.104 ; 
        RECT 0.488 22.466 0.56 27.106 ; 
        RECT 120.872 26.786 120.944 31.426 ; 
        RECT 64.784 26.788 64.856 31.424 ; 
        RECT 59.168 26.932 59.528 31.394 ; 
        RECT 56.576 26.788 56.648 31.424 ; 
        RECT 0.488 26.786 0.56 31.426 ; 
        RECT 120.872 31.106 120.944 35.746 ; 
        RECT 64.784 31.108 64.856 35.744 ; 
        RECT 59.168 31.252 59.528 35.714 ; 
        RECT 56.576 31.108 56.648 35.744 ; 
        RECT 0.488 31.106 0.56 35.746 ; 
        RECT 120.872 35.426 120.944 40.066 ; 
        RECT 64.784 35.428 64.856 40.064 ; 
        RECT 59.168 35.572 59.528 40.034 ; 
        RECT 56.576 35.428 56.648 40.064 ; 
        RECT 0.488 35.426 0.56 40.066 ; 
        RECT 120.872 39.746 120.944 44.386 ; 
        RECT 64.784 39.748 64.856 44.384 ; 
        RECT 59.168 39.892 59.528 44.354 ; 
        RECT 56.576 39.748 56.648 44.384 ; 
        RECT 0.488 39.746 0.56 44.386 ; 
        RECT 120.872 44.066 120.944 48.706 ; 
        RECT 64.784 44.068 64.856 48.704 ; 
        RECT 59.168 44.212 59.528 48.674 ; 
        RECT 56.576 44.068 56.648 48.704 ; 
        RECT 0.488 44.066 0.56 48.706 ; 
        RECT 120.872 48.386 120.944 53.026 ; 
        RECT 64.784 48.388 64.856 53.024 ; 
        RECT 59.168 48.532 59.528 52.994 ; 
        RECT 56.576 48.388 56.648 53.024 ; 
        RECT 0.488 48.386 0.56 53.026 ; 
        RECT 120.872 52.706 120.944 57.346 ; 
        RECT 64.784 52.708 64.856 57.344 ; 
        RECT 59.168 52.852 59.528 57.314 ; 
        RECT 56.576 52.708 56.648 57.344 ; 
        RECT 0.488 52.706 0.56 57.346 ; 
        RECT 120.872 57.026 120.944 61.666 ; 
        RECT 64.784 57.028 64.856 61.664 ; 
        RECT 59.168 57.172 59.528 61.634 ; 
        RECT 56.576 57.028 56.648 61.664 ; 
        RECT 0.488 57.026 0.56 61.666 ; 
        RECT 120.872 61.346 120.944 65.986 ; 
        RECT 64.784 61.348 64.856 65.984 ; 
        RECT 59.168 61.492 59.528 65.954 ; 
        RECT 56.576 61.348 56.648 65.984 ; 
        RECT 0.488 61.346 0.56 65.986 ; 
        RECT 120.872 65.666 120.944 70.306 ; 
        RECT 64.784 65.668 64.856 70.304 ; 
        RECT 59.168 65.812 59.528 70.274 ; 
        RECT 56.576 65.668 56.648 70.304 ; 
        RECT 0.488 65.666 0.56 70.306 ; 
        RECT 120.872 69.986 120.944 74.626 ; 
        RECT 64.784 69.988 64.856 74.624 ; 
        RECT 59.168 70.132 59.528 74.594 ; 
        RECT 56.576 69.988 56.648 74.624 ; 
        RECT 0.488 69.986 0.56 74.626 ; 
        RECT 120.872 74.306 120.944 78.946 ; 
        RECT 64.784 74.308 64.856 78.944 ; 
        RECT 59.168 74.452 59.528 78.914 ; 
        RECT 56.576 74.308 56.648 78.944 ; 
        RECT 0.488 74.306 0.56 78.946 ; 
        RECT 120.872 78.626 120.944 83.266 ; 
        RECT 64.784 78.628 64.856 83.264 ; 
        RECT 59.168 78.772 59.528 83.234 ; 
        RECT 56.576 78.628 56.648 83.264 ; 
        RECT 0.488 78.626 0.56 83.266 ; 
        RECT 120.872 82.946 120.944 87.586 ; 
        RECT 64.784 82.948 64.856 87.584 ; 
        RECT 59.168 83.092 59.528 87.554 ; 
        RECT 56.576 82.948 56.648 87.584 ; 
        RECT 0.488 82.946 0.56 87.586 ; 
        RECT 120.872 87.266 120.944 91.906 ; 
        RECT 64.784 87.268 64.856 91.904 ; 
        RECT 59.168 87.412 59.528 91.874 ; 
        RECT 56.576 87.268 56.648 91.904 ; 
        RECT 0.488 87.266 0.56 91.906 ; 
        RECT 120.872 91.586 120.944 96.226 ; 
        RECT 64.784 91.588 64.856 96.224 ; 
        RECT 59.168 91.732 59.528 96.194 ; 
        RECT 56.576 91.588 56.648 96.224 ; 
        RECT 0.488 91.586 0.56 96.226 ; 
        RECT 120.872 95.906 120.944 100.546 ; 
        RECT 64.784 95.908 64.856 100.544 ; 
        RECT 59.168 96.052 59.528 100.514 ; 
        RECT 56.576 95.908 56.648 100.544 ; 
        RECT 0.488 95.906 0.56 100.546 ; 
        RECT 120.872 100.226 120.944 104.866 ; 
        RECT 64.784 100.228 64.856 104.864 ; 
        RECT 59.168 100.372 59.528 104.834 ; 
        RECT 56.576 100.228 56.648 104.864 ; 
        RECT 0.488 100.226 0.56 104.866 ; 
        RECT 56.196 120.02 56.268 144.274 ; 
        RECT 120.872 137.054 120.944 141.694 ; 
        RECT 64.784 137.056 64.856 141.692 ; 
        RECT 59.168 137.2 59.528 141.662 ; 
        RECT 56.576 137.056 56.648 141.692 ; 
        RECT 0.488 137.054 0.56 141.694 ; 
        RECT 120.872 141.374 120.944 146.014 ; 
        RECT 64.784 141.376 64.856 146.012 ; 
        RECT 59.168 141.52 59.528 145.982 ; 
        RECT 56.576 141.376 56.648 146.012 ; 
        RECT 0.488 141.374 0.56 146.014 ; 
        RECT 120.872 145.694 120.944 150.334 ; 
        RECT 64.784 145.696 64.856 150.332 ; 
        RECT 59.168 145.84 59.528 150.302 ; 
        RECT 56.576 145.696 56.648 150.332 ; 
        RECT 0.488 145.694 0.56 150.334 ; 
        RECT 120.872 150.014 120.944 154.654 ; 
        RECT 64.784 150.016 64.856 154.652 ; 
        RECT 59.168 150.16 59.528 154.622 ; 
        RECT 56.576 150.016 56.648 154.652 ; 
        RECT 0.488 150.014 0.56 154.654 ; 
        RECT 120.872 154.334 120.944 158.974 ; 
        RECT 64.784 154.336 64.856 158.972 ; 
        RECT 59.168 154.48 59.528 158.942 ; 
        RECT 56.576 154.336 56.648 158.972 ; 
        RECT 0.488 154.334 0.56 158.974 ; 
        RECT 120.872 158.654 120.944 163.294 ; 
        RECT 64.784 158.656 64.856 163.292 ; 
        RECT 59.168 158.8 59.528 163.262 ; 
        RECT 56.576 158.656 56.648 163.292 ; 
        RECT 0.488 158.654 0.56 163.294 ; 
        RECT 120.872 162.974 120.944 167.614 ; 
        RECT 64.784 162.976 64.856 167.612 ; 
        RECT 59.168 163.12 59.528 167.582 ; 
        RECT 56.576 162.976 56.648 167.612 ; 
        RECT 0.488 162.974 0.56 167.614 ; 
        RECT 120.872 167.294 120.944 171.934 ; 
        RECT 64.784 167.296 64.856 171.932 ; 
        RECT 59.168 167.44 59.528 171.902 ; 
        RECT 56.576 167.296 56.648 171.932 ; 
        RECT 0.488 167.294 0.56 171.934 ; 
        RECT 120.872 171.614 120.944 176.254 ; 
        RECT 64.784 171.616 64.856 176.252 ; 
        RECT 59.168 171.76 59.528 176.222 ; 
        RECT 56.576 171.616 56.648 176.252 ; 
        RECT 0.488 171.614 0.56 176.254 ; 
        RECT 120.872 175.934 120.944 180.574 ; 
        RECT 64.784 175.936 64.856 180.572 ; 
        RECT 59.168 176.08 59.528 180.542 ; 
        RECT 56.576 175.936 56.648 180.572 ; 
        RECT 0.488 175.934 0.56 180.574 ; 
        RECT 120.872 180.254 120.944 184.894 ; 
        RECT 64.784 180.256 64.856 184.892 ; 
        RECT 59.168 180.4 59.528 184.862 ; 
        RECT 56.576 180.256 56.648 184.892 ; 
        RECT 0.488 180.254 0.56 184.894 ; 
        RECT 120.872 184.574 120.944 189.214 ; 
        RECT 64.784 184.576 64.856 189.212 ; 
        RECT 59.168 184.72 59.528 189.182 ; 
        RECT 56.576 184.576 56.648 189.212 ; 
        RECT 0.488 184.574 0.56 189.214 ; 
        RECT 120.872 188.894 120.944 193.534 ; 
        RECT 64.784 188.896 64.856 193.532 ; 
        RECT 59.168 189.04 59.528 193.502 ; 
        RECT 56.576 188.896 56.648 193.532 ; 
        RECT 0.488 188.894 0.56 193.534 ; 
        RECT 120.872 193.214 120.944 197.854 ; 
        RECT 64.784 193.216 64.856 197.852 ; 
        RECT 59.168 193.36 59.528 197.822 ; 
        RECT 56.576 193.216 56.648 197.852 ; 
        RECT 0.488 193.214 0.56 197.854 ; 
        RECT 120.872 197.534 120.944 202.174 ; 
        RECT 64.784 197.536 64.856 202.172 ; 
        RECT 59.168 197.68 59.528 202.142 ; 
        RECT 56.576 197.536 56.648 202.172 ; 
        RECT 0.488 197.534 0.56 202.174 ; 
        RECT 120.872 201.854 120.944 206.494 ; 
        RECT 64.784 201.856 64.856 206.492 ; 
        RECT 59.168 202 59.528 206.462 ; 
        RECT 56.576 201.856 56.648 206.492 ; 
        RECT 0.488 201.854 0.56 206.494 ; 
        RECT 120.872 206.174 120.944 210.814 ; 
        RECT 64.784 206.176 64.856 210.812 ; 
        RECT 59.168 206.32 59.528 210.782 ; 
        RECT 56.576 206.176 56.648 210.812 ; 
        RECT 0.488 206.174 0.56 210.814 ; 
        RECT 120.872 210.494 120.944 215.134 ; 
        RECT 64.784 210.496 64.856 215.132 ; 
        RECT 59.168 210.64 59.528 215.102 ; 
        RECT 56.576 210.496 56.648 215.132 ; 
        RECT 0.488 210.494 0.56 215.134 ; 
        RECT 120.872 214.814 120.944 219.454 ; 
        RECT 64.784 214.816 64.856 219.452 ; 
        RECT 59.168 214.96 59.528 219.422 ; 
        RECT 56.576 214.816 56.648 219.452 ; 
        RECT 0.488 214.814 0.56 219.454 ; 
        RECT 120.872 219.134 120.944 223.774 ; 
        RECT 64.784 219.136 64.856 223.772 ; 
        RECT 59.168 219.28 59.528 223.742 ; 
        RECT 56.576 219.136 56.648 223.772 ; 
        RECT 0.488 219.134 0.56 223.774 ; 
        RECT 120.872 223.454 120.944 228.094 ; 
        RECT 64.784 223.456 64.856 228.092 ; 
        RECT 59.168 223.6 59.528 228.062 ; 
        RECT 56.576 223.456 56.648 228.092 ; 
        RECT 0.488 223.454 0.56 228.094 ; 
        RECT 120.872 227.774 120.944 232.414 ; 
        RECT 64.784 227.776 64.856 232.412 ; 
        RECT 59.168 227.92 59.528 232.382 ; 
        RECT 56.576 227.776 56.648 232.412 ; 
        RECT 0.488 227.774 0.56 232.414 ; 
        RECT 120.872 232.094 120.944 236.734 ; 
        RECT 64.784 232.096 64.856 236.732 ; 
        RECT 59.168 232.24 59.528 236.702 ; 
        RECT 56.576 232.096 56.648 236.732 ; 
        RECT 0.488 232.094 0.56 236.734 ; 
        RECT 120.872 236.414 120.944 241.054 ; 
        RECT 64.784 236.416 64.856 241.052 ; 
        RECT 59.168 236.56 59.528 241.022 ; 
        RECT 56.576 236.416 56.648 241.052 ; 
        RECT 0.488 236.414 0.56 241.054 ; 
      LAYER V3 ; 
        RECT 0.488 4.688 0.56 4.88 ; 
        RECT 56.576 4.688 56.648 4.88 ; 
        RECT 59.168 4.688 59.528 4.88 ; 
        RECT 64.784 4.688 64.856 4.88 ; 
        RECT 120.872 4.688 120.944 4.88 ; 
        RECT 0.488 9.008 0.56 9.2 ; 
        RECT 56.576 9.008 56.648 9.2 ; 
        RECT 59.168 9.008 59.528 9.2 ; 
        RECT 64.784 9.008 64.856 9.2 ; 
        RECT 120.872 9.008 120.944 9.2 ; 
        RECT 0.488 13.328 0.56 13.52 ; 
        RECT 56.576 13.328 56.648 13.52 ; 
        RECT 59.168 13.328 59.528 13.52 ; 
        RECT 64.784 13.328 64.856 13.52 ; 
        RECT 120.872 13.328 120.944 13.52 ; 
        RECT 0.488 17.648 0.56 17.84 ; 
        RECT 56.576 17.648 56.648 17.84 ; 
        RECT 59.168 17.648 59.528 17.84 ; 
        RECT 64.784 17.648 64.856 17.84 ; 
        RECT 120.872 17.648 120.944 17.84 ; 
        RECT 0.488 21.968 0.56 22.16 ; 
        RECT 56.576 21.968 56.648 22.16 ; 
        RECT 59.168 21.968 59.528 22.16 ; 
        RECT 64.784 21.968 64.856 22.16 ; 
        RECT 120.872 21.968 120.944 22.16 ; 
        RECT 0.488 26.288 0.56 26.48 ; 
        RECT 56.576 26.288 56.648 26.48 ; 
        RECT 59.168 26.288 59.528 26.48 ; 
        RECT 64.784 26.288 64.856 26.48 ; 
        RECT 120.872 26.288 120.944 26.48 ; 
        RECT 0.488 30.608 0.56 30.8 ; 
        RECT 56.576 30.608 56.648 30.8 ; 
        RECT 59.168 30.608 59.528 30.8 ; 
        RECT 64.784 30.608 64.856 30.8 ; 
        RECT 120.872 30.608 120.944 30.8 ; 
        RECT 0.488 34.928 0.56 35.12 ; 
        RECT 56.576 34.928 56.648 35.12 ; 
        RECT 59.168 34.928 59.528 35.12 ; 
        RECT 64.784 34.928 64.856 35.12 ; 
        RECT 120.872 34.928 120.944 35.12 ; 
        RECT 0.488 39.248 0.56 39.44 ; 
        RECT 56.576 39.248 56.648 39.44 ; 
        RECT 59.168 39.248 59.528 39.44 ; 
        RECT 64.784 39.248 64.856 39.44 ; 
        RECT 120.872 39.248 120.944 39.44 ; 
        RECT 0.488 43.568 0.56 43.76 ; 
        RECT 56.576 43.568 56.648 43.76 ; 
        RECT 59.168 43.568 59.528 43.76 ; 
        RECT 64.784 43.568 64.856 43.76 ; 
        RECT 120.872 43.568 120.944 43.76 ; 
        RECT 0.488 47.888 0.56 48.08 ; 
        RECT 56.576 47.888 56.648 48.08 ; 
        RECT 59.168 47.888 59.528 48.08 ; 
        RECT 64.784 47.888 64.856 48.08 ; 
        RECT 120.872 47.888 120.944 48.08 ; 
        RECT 0.488 52.208 0.56 52.4 ; 
        RECT 56.576 52.208 56.648 52.4 ; 
        RECT 59.168 52.208 59.528 52.4 ; 
        RECT 64.784 52.208 64.856 52.4 ; 
        RECT 120.872 52.208 120.944 52.4 ; 
        RECT 0.488 56.528 0.56 56.72 ; 
        RECT 56.576 56.528 56.648 56.72 ; 
        RECT 59.168 56.528 59.528 56.72 ; 
        RECT 64.784 56.528 64.856 56.72 ; 
        RECT 120.872 56.528 120.944 56.72 ; 
        RECT 0.488 60.848 0.56 61.04 ; 
        RECT 56.576 60.848 56.648 61.04 ; 
        RECT 59.168 60.848 59.528 61.04 ; 
        RECT 64.784 60.848 64.856 61.04 ; 
        RECT 120.872 60.848 120.944 61.04 ; 
        RECT 0.488 65.168 0.56 65.36 ; 
        RECT 56.576 65.168 56.648 65.36 ; 
        RECT 59.168 65.168 59.528 65.36 ; 
        RECT 64.784 65.168 64.856 65.36 ; 
        RECT 120.872 65.168 120.944 65.36 ; 
        RECT 0.488 69.488 0.56 69.68 ; 
        RECT 56.576 69.488 56.648 69.68 ; 
        RECT 59.168 69.488 59.528 69.68 ; 
        RECT 64.784 69.488 64.856 69.68 ; 
        RECT 120.872 69.488 120.944 69.68 ; 
        RECT 0.488 73.808 0.56 74 ; 
        RECT 56.576 73.808 56.648 74 ; 
        RECT 59.168 73.808 59.528 74 ; 
        RECT 64.784 73.808 64.856 74 ; 
        RECT 120.872 73.808 120.944 74 ; 
        RECT 0.488 78.128 0.56 78.32 ; 
        RECT 56.576 78.128 56.648 78.32 ; 
        RECT 59.168 78.128 59.528 78.32 ; 
        RECT 64.784 78.128 64.856 78.32 ; 
        RECT 120.872 78.128 120.944 78.32 ; 
        RECT 0.488 82.448 0.56 82.64 ; 
        RECT 56.576 82.448 56.648 82.64 ; 
        RECT 59.168 82.448 59.528 82.64 ; 
        RECT 64.784 82.448 64.856 82.64 ; 
        RECT 120.872 82.448 120.944 82.64 ; 
        RECT 0.488 86.768 0.56 86.96 ; 
        RECT 56.576 86.768 56.648 86.96 ; 
        RECT 59.168 86.768 59.528 86.96 ; 
        RECT 64.784 86.768 64.856 86.96 ; 
        RECT 120.872 86.768 120.944 86.96 ; 
        RECT 0.488 91.088 0.56 91.28 ; 
        RECT 56.576 91.088 56.648 91.28 ; 
        RECT 59.168 91.088 59.528 91.28 ; 
        RECT 64.784 91.088 64.856 91.28 ; 
        RECT 120.872 91.088 120.944 91.28 ; 
        RECT 0.488 95.408 0.56 95.6 ; 
        RECT 56.576 95.408 56.648 95.6 ; 
        RECT 59.168 95.408 59.528 95.6 ; 
        RECT 64.784 95.408 64.856 95.6 ; 
        RECT 120.872 95.408 120.944 95.6 ; 
        RECT 0.488 99.728 0.56 99.92 ; 
        RECT 56.576 99.728 56.648 99.92 ; 
        RECT 59.168 99.728 59.528 99.92 ; 
        RECT 64.784 99.728 64.856 99.92 ; 
        RECT 120.872 99.728 120.944 99.92 ; 
        RECT 0.488 104.048 0.56 104.24 ; 
        RECT 56.576 104.048 56.648 104.24 ; 
        RECT 59.168 104.048 59.528 104.24 ; 
        RECT 64.784 104.048 64.856 104.24 ; 
        RECT 120.872 104.048 120.944 104.24 ; 
        RECT 0.488 140.876 0.56 141.068 ; 
        RECT 56.576 140.876 56.648 141.068 ; 
        RECT 59.168 140.876 59.528 141.068 ; 
        RECT 64.784 140.876 64.856 141.068 ; 
        RECT 120.872 140.876 120.944 141.068 ; 
        RECT 0.488 145.196 0.56 145.388 ; 
        RECT 56.576 145.196 56.648 145.388 ; 
        RECT 59.168 145.196 59.528 145.388 ; 
        RECT 64.784 145.196 64.856 145.388 ; 
        RECT 120.872 145.196 120.944 145.388 ; 
        RECT 0.488 149.516 0.56 149.708 ; 
        RECT 56.576 149.516 56.648 149.708 ; 
        RECT 59.168 149.516 59.528 149.708 ; 
        RECT 64.784 149.516 64.856 149.708 ; 
        RECT 120.872 149.516 120.944 149.708 ; 
        RECT 0.488 153.836 0.56 154.028 ; 
        RECT 56.576 153.836 56.648 154.028 ; 
        RECT 59.168 153.836 59.528 154.028 ; 
        RECT 64.784 153.836 64.856 154.028 ; 
        RECT 120.872 153.836 120.944 154.028 ; 
        RECT 0.488 158.156 0.56 158.348 ; 
        RECT 56.576 158.156 56.648 158.348 ; 
        RECT 59.168 158.156 59.528 158.348 ; 
        RECT 64.784 158.156 64.856 158.348 ; 
        RECT 120.872 158.156 120.944 158.348 ; 
        RECT 0.488 162.476 0.56 162.668 ; 
        RECT 56.576 162.476 56.648 162.668 ; 
        RECT 59.168 162.476 59.528 162.668 ; 
        RECT 64.784 162.476 64.856 162.668 ; 
        RECT 120.872 162.476 120.944 162.668 ; 
        RECT 0.488 166.796 0.56 166.988 ; 
        RECT 56.576 166.796 56.648 166.988 ; 
        RECT 59.168 166.796 59.528 166.988 ; 
        RECT 64.784 166.796 64.856 166.988 ; 
        RECT 120.872 166.796 120.944 166.988 ; 
        RECT 0.488 171.116 0.56 171.308 ; 
        RECT 56.576 171.116 56.648 171.308 ; 
        RECT 59.168 171.116 59.528 171.308 ; 
        RECT 64.784 171.116 64.856 171.308 ; 
        RECT 120.872 171.116 120.944 171.308 ; 
        RECT 0.488 175.436 0.56 175.628 ; 
        RECT 56.576 175.436 56.648 175.628 ; 
        RECT 59.168 175.436 59.528 175.628 ; 
        RECT 64.784 175.436 64.856 175.628 ; 
        RECT 120.872 175.436 120.944 175.628 ; 
        RECT 0.488 179.756 0.56 179.948 ; 
        RECT 56.576 179.756 56.648 179.948 ; 
        RECT 59.168 179.756 59.528 179.948 ; 
        RECT 64.784 179.756 64.856 179.948 ; 
        RECT 120.872 179.756 120.944 179.948 ; 
        RECT 0.488 184.076 0.56 184.268 ; 
        RECT 56.576 184.076 56.648 184.268 ; 
        RECT 59.168 184.076 59.528 184.268 ; 
        RECT 64.784 184.076 64.856 184.268 ; 
        RECT 120.872 184.076 120.944 184.268 ; 
        RECT 0.488 188.396 0.56 188.588 ; 
        RECT 56.576 188.396 56.648 188.588 ; 
        RECT 59.168 188.396 59.528 188.588 ; 
        RECT 64.784 188.396 64.856 188.588 ; 
        RECT 120.872 188.396 120.944 188.588 ; 
        RECT 0.488 192.716 0.56 192.908 ; 
        RECT 56.576 192.716 56.648 192.908 ; 
        RECT 59.168 192.716 59.528 192.908 ; 
        RECT 64.784 192.716 64.856 192.908 ; 
        RECT 120.872 192.716 120.944 192.908 ; 
        RECT 0.488 197.036 0.56 197.228 ; 
        RECT 56.576 197.036 56.648 197.228 ; 
        RECT 59.168 197.036 59.528 197.228 ; 
        RECT 64.784 197.036 64.856 197.228 ; 
        RECT 120.872 197.036 120.944 197.228 ; 
        RECT 0.488 201.356 0.56 201.548 ; 
        RECT 56.576 201.356 56.648 201.548 ; 
        RECT 59.168 201.356 59.528 201.548 ; 
        RECT 64.784 201.356 64.856 201.548 ; 
        RECT 120.872 201.356 120.944 201.548 ; 
        RECT 0.488 205.676 0.56 205.868 ; 
        RECT 56.576 205.676 56.648 205.868 ; 
        RECT 59.168 205.676 59.528 205.868 ; 
        RECT 64.784 205.676 64.856 205.868 ; 
        RECT 120.872 205.676 120.944 205.868 ; 
        RECT 0.488 209.996 0.56 210.188 ; 
        RECT 56.576 209.996 56.648 210.188 ; 
        RECT 59.168 209.996 59.528 210.188 ; 
        RECT 64.784 209.996 64.856 210.188 ; 
        RECT 120.872 209.996 120.944 210.188 ; 
        RECT 0.488 214.316 0.56 214.508 ; 
        RECT 56.576 214.316 56.648 214.508 ; 
        RECT 59.168 214.316 59.528 214.508 ; 
        RECT 64.784 214.316 64.856 214.508 ; 
        RECT 120.872 214.316 120.944 214.508 ; 
        RECT 0.488 218.636 0.56 218.828 ; 
        RECT 56.576 218.636 56.648 218.828 ; 
        RECT 59.168 218.636 59.528 218.828 ; 
        RECT 64.784 218.636 64.856 218.828 ; 
        RECT 120.872 218.636 120.944 218.828 ; 
        RECT 0.488 222.956 0.56 223.148 ; 
        RECT 56.576 222.956 56.648 223.148 ; 
        RECT 59.168 222.956 59.528 223.148 ; 
        RECT 64.784 222.956 64.856 223.148 ; 
        RECT 120.872 222.956 120.944 223.148 ; 
        RECT 0.488 227.276 0.56 227.468 ; 
        RECT 56.576 227.276 56.648 227.468 ; 
        RECT 59.168 227.276 59.528 227.468 ; 
        RECT 64.784 227.276 64.856 227.468 ; 
        RECT 120.872 227.276 120.944 227.468 ; 
        RECT 0.488 231.596 0.56 231.788 ; 
        RECT 56.576 231.596 56.648 231.788 ; 
        RECT 59.168 231.596 59.528 231.788 ; 
        RECT 64.784 231.596 64.856 231.788 ; 
        RECT 120.872 231.596 120.944 231.788 ; 
        RECT 0.488 235.916 0.56 236.108 ; 
        RECT 56.576 235.916 56.648 236.108 ; 
        RECT 59.168 235.916 59.528 236.108 ; 
        RECT 64.784 235.916 64.856 236.108 ; 
        RECT 120.872 235.916 120.944 236.108 ; 
        RECT 0.488 240.236 0.56 240.428 ; 
        RECT 56.576 240.236 56.648 240.428 ; 
        RECT 59.168 240.236 59.528 240.428 ; 
        RECT 64.784 240.236 64.856 240.428 ; 
        RECT 120.872 240.236 120.944 240.428 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.416 4.304 121.032 4.496 ; 
        RECT 0.416 8.624 121.032 8.816 ; 
        RECT 0.416 12.944 121.032 13.136 ; 
        RECT 0.416 17.264 121.032 17.456 ; 
        RECT 0.416 21.584 121.032 21.776 ; 
        RECT 0.416 25.904 121.032 26.096 ; 
        RECT 0.416 30.224 121.032 30.416 ; 
        RECT 0.416 34.544 121.032 34.736 ; 
        RECT 0.416 38.864 121.032 39.056 ; 
        RECT 0.416 43.184 121.032 43.376 ; 
        RECT 0.416 47.504 121.032 47.696 ; 
        RECT 0.416 51.824 121.032 52.016 ; 
        RECT 0.416 56.144 121.032 56.336 ; 
        RECT 0.416 60.464 121.032 60.656 ; 
        RECT 0.416 64.784 121.032 64.976 ; 
        RECT 0.416 69.104 121.032 69.296 ; 
        RECT 0.416 73.424 121.032 73.616 ; 
        RECT 0.416 77.744 121.032 77.936 ; 
        RECT 0.416 82.064 121.032 82.256 ; 
        RECT 0.416 86.384 121.032 86.576 ; 
        RECT 0.416 90.704 121.032 90.896 ; 
        RECT 0.416 95.024 121.032 95.216 ; 
        RECT 0.416 99.344 121.032 99.536 ; 
        RECT 0.416 103.664 121.032 103.856 ; 
        RECT 41.904 107.926 79.488 108.79 ; 
        RECT 57.24 120.598 64.152 121.462 ; 
        RECT 57.24 133.27 64.152 134.134 ; 
        RECT 0.416 140.492 121.032 140.684 ; 
        RECT 0.416 144.812 121.032 145.004 ; 
        RECT 0.416 149.132 121.032 149.324 ; 
        RECT 0.416 153.452 121.032 153.644 ; 
        RECT 0.416 157.772 121.032 157.964 ; 
        RECT 0.416 162.092 121.032 162.284 ; 
        RECT 0.416 166.412 121.032 166.604 ; 
        RECT 0.416 170.732 121.032 170.924 ; 
        RECT 0.416 175.052 121.032 175.244 ; 
        RECT 0.416 179.372 121.032 179.564 ; 
        RECT 0.416 183.692 121.032 183.884 ; 
        RECT 0.416 188.012 121.032 188.204 ; 
        RECT 0.416 192.332 121.032 192.524 ; 
        RECT 0.416 196.652 121.032 196.844 ; 
        RECT 0.416 200.972 121.032 201.164 ; 
        RECT 0.416 205.292 121.032 205.484 ; 
        RECT 0.416 209.612 121.032 209.804 ; 
        RECT 0.416 213.932 121.032 214.124 ; 
        RECT 0.416 218.252 121.032 218.444 ; 
        RECT 0.416 222.572 121.032 222.764 ; 
        RECT 0.416 226.892 121.032 227.084 ; 
        RECT 0.416 231.212 121.032 231.404 ; 
        RECT 0.416 235.532 121.032 235.724 ; 
        RECT 0.416 239.852 121.032 240.044 ; 
      LAYER M3 ; 
        RECT 120.728 0.866 120.8 5.506 ; 
        RECT 65 0.866 65.072 5.506 ; 
        RECT 61.94 1.012 62.084 5.47 ; 
        RECT 61.04 1.012 61.148 5.47 ; 
        RECT 56.36 0.866 56.432 5.506 ; 
        RECT 0.632 0.866 0.704 5.506 ; 
        RECT 120.728 5.186 120.8 9.826 ; 
        RECT 65 5.186 65.072 9.826 ; 
        RECT 61.94 5.332 62.084 9.79 ; 
        RECT 61.04 5.332 61.148 9.79 ; 
        RECT 56.36 5.186 56.432 9.826 ; 
        RECT 0.632 5.186 0.704 9.826 ; 
        RECT 120.728 9.506 120.8 14.146 ; 
        RECT 65 9.506 65.072 14.146 ; 
        RECT 61.94 9.652 62.084 14.11 ; 
        RECT 61.04 9.652 61.148 14.11 ; 
        RECT 56.36 9.506 56.432 14.146 ; 
        RECT 0.632 9.506 0.704 14.146 ; 
        RECT 120.728 13.826 120.8 18.466 ; 
        RECT 65 13.826 65.072 18.466 ; 
        RECT 61.94 13.972 62.084 18.43 ; 
        RECT 61.04 13.972 61.148 18.43 ; 
        RECT 56.36 13.826 56.432 18.466 ; 
        RECT 0.632 13.826 0.704 18.466 ; 
        RECT 120.728 18.146 120.8 22.786 ; 
        RECT 65 18.146 65.072 22.786 ; 
        RECT 61.94 18.292 62.084 22.75 ; 
        RECT 61.04 18.292 61.148 22.75 ; 
        RECT 56.36 18.146 56.432 22.786 ; 
        RECT 0.632 18.146 0.704 22.786 ; 
        RECT 120.728 22.466 120.8 27.106 ; 
        RECT 65 22.466 65.072 27.106 ; 
        RECT 61.94 22.612 62.084 27.07 ; 
        RECT 61.04 22.612 61.148 27.07 ; 
        RECT 56.36 22.466 56.432 27.106 ; 
        RECT 0.632 22.466 0.704 27.106 ; 
        RECT 120.728 26.786 120.8 31.426 ; 
        RECT 65 26.786 65.072 31.426 ; 
        RECT 61.94 26.932 62.084 31.39 ; 
        RECT 61.04 26.932 61.148 31.39 ; 
        RECT 56.36 26.786 56.432 31.426 ; 
        RECT 0.632 26.786 0.704 31.426 ; 
        RECT 120.728 31.106 120.8 35.746 ; 
        RECT 65 31.106 65.072 35.746 ; 
        RECT 61.94 31.252 62.084 35.71 ; 
        RECT 61.04 31.252 61.148 35.71 ; 
        RECT 56.36 31.106 56.432 35.746 ; 
        RECT 0.632 31.106 0.704 35.746 ; 
        RECT 120.728 35.426 120.8 40.066 ; 
        RECT 65 35.426 65.072 40.066 ; 
        RECT 61.94 35.572 62.084 40.03 ; 
        RECT 61.04 35.572 61.148 40.03 ; 
        RECT 56.36 35.426 56.432 40.066 ; 
        RECT 0.632 35.426 0.704 40.066 ; 
        RECT 120.728 39.746 120.8 44.386 ; 
        RECT 65 39.746 65.072 44.386 ; 
        RECT 61.94 39.892 62.084 44.35 ; 
        RECT 61.04 39.892 61.148 44.35 ; 
        RECT 56.36 39.746 56.432 44.386 ; 
        RECT 0.632 39.746 0.704 44.386 ; 
        RECT 120.728 44.066 120.8 48.706 ; 
        RECT 65 44.066 65.072 48.706 ; 
        RECT 61.94 44.212 62.084 48.67 ; 
        RECT 61.04 44.212 61.148 48.67 ; 
        RECT 56.36 44.066 56.432 48.706 ; 
        RECT 0.632 44.066 0.704 48.706 ; 
        RECT 120.728 48.386 120.8 53.026 ; 
        RECT 65 48.386 65.072 53.026 ; 
        RECT 61.94 48.532 62.084 52.99 ; 
        RECT 61.04 48.532 61.148 52.99 ; 
        RECT 56.36 48.386 56.432 53.026 ; 
        RECT 0.632 48.386 0.704 53.026 ; 
        RECT 120.728 52.706 120.8 57.346 ; 
        RECT 65 52.706 65.072 57.346 ; 
        RECT 61.94 52.852 62.084 57.31 ; 
        RECT 61.04 52.852 61.148 57.31 ; 
        RECT 56.36 52.706 56.432 57.346 ; 
        RECT 0.632 52.706 0.704 57.346 ; 
        RECT 120.728 57.026 120.8 61.666 ; 
        RECT 65 57.026 65.072 61.666 ; 
        RECT 61.94 57.172 62.084 61.63 ; 
        RECT 61.04 57.172 61.148 61.63 ; 
        RECT 56.36 57.026 56.432 61.666 ; 
        RECT 0.632 57.026 0.704 61.666 ; 
        RECT 120.728 61.346 120.8 65.986 ; 
        RECT 65 61.346 65.072 65.986 ; 
        RECT 61.94 61.492 62.084 65.95 ; 
        RECT 61.04 61.492 61.148 65.95 ; 
        RECT 56.36 61.346 56.432 65.986 ; 
        RECT 0.632 61.346 0.704 65.986 ; 
        RECT 120.728 65.666 120.8 70.306 ; 
        RECT 65 65.666 65.072 70.306 ; 
        RECT 61.94 65.812 62.084 70.27 ; 
        RECT 61.04 65.812 61.148 70.27 ; 
        RECT 56.36 65.666 56.432 70.306 ; 
        RECT 0.632 65.666 0.704 70.306 ; 
        RECT 120.728 69.986 120.8 74.626 ; 
        RECT 65 69.986 65.072 74.626 ; 
        RECT 61.94 70.132 62.084 74.59 ; 
        RECT 61.04 70.132 61.148 74.59 ; 
        RECT 56.36 69.986 56.432 74.626 ; 
        RECT 0.632 69.986 0.704 74.626 ; 
        RECT 120.728 74.306 120.8 78.946 ; 
        RECT 65 74.306 65.072 78.946 ; 
        RECT 61.94 74.452 62.084 78.91 ; 
        RECT 61.04 74.452 61.148 78.91 ; 
        RECT 56.36 74.306 56.432 78.946 ; 
        RECT 0.632 74.306 0.704 78.946 ; 
        RECT 120.728 78.626 120.8 83.266 ; 
        RECT 65 78.626 65.072 83.266 ; 
        RECT 61.94 78.772 62.084 83.23 ; 
        RECT 61.04 78.772 61.148 83.23 ; 
        RECT 56.36 78.626 56.432 83.266 ; 
        RECT 0.632 78.626 0.704 83.266 ; 
        RECT 120.728 82.946 120.8 87.586 ; 
        RECT 65 82.946 65.072 87.586 ; 
        RECT 61.94 83.092 62.084 87.55 ; 
        RECT 61.04 83.092 61.148 87.55 ; 
        RECT 56.36 82.946 56.432 87.586 ; 
        RECT 0.632 82.946 0.704 87.586 ; 
        RECT 120.728 87.266 120.8 91.906 ; 
        RECT 65 87.266 65.072 91.906 ; 
        RECT 61.94 87.412 62.084 91.87 ; 
        RECT 61.04 87.412 61.148 91.87 ; 
        RECT 56.36 87.266 56.432 91.906 ; 
        RECT 0.632 87.266 0.704 91.906 ; 
        RECT 120.728 91.586 120.8 96.226 ; 
        RECT 65 91.586 65.072 96.226 ; 
        RECT 61.94 91.732 62.084 96.19 ; 
        RECT 61.04 91.732 61.148 96.19 ; 
        RECT 56.36 91.586 56.432 96.226 ; 
        RECT 0.632 91.586 0.704 96.226 ; 
        RECT 120.728 95.906 120.8 100.546 ; 
        RECT 65 95.906 65.072 100.546 ; 
        RECT 61.94 96.052 62.084 100.51 ; 
        RECT 61.04 96.052 61.148 100.51 ; 
        RECT 56.36 95.906 56.432 100.546 ; 
        RECT 0.632 95.906 0.704 100.546 ; 
        RECT 120.728 100.226 120.8 104.866 ; 
        RECT 65 100.226 65.072 104.866 ; 
        RECT 61.94 100.372 62.084 104.83 ; 
        RECT 61.04 100.372 61.148 104.83 ; 
        RECT 56.36 100.226 56.432 104.866 ; 
        RECT 0.632 100.226 0.704 104.866 ; 
        RECT 64.98 104.748 65.052 137.576 ; 
        RECT 61.164 105.642 62.1 136.374 ; 
        RECT 56.34 104.748 56.412 144.274 ; 
        RECT 120.728 137.054 120.8 141.694 ; 
        RECT 65 137.054 65.072 141.694 ; 
        RECT 61.94 137.2 62.084 141.658 ; 
        RECT 61.04 137.2 61.148 141.658 ; 
        RECT 56.36 137.054 56.432 141.694 ; 
        RECT 0.632 137.054 0.704 141.694 ; 
        RECT 120.728 141.374 120.8 146.014 ; 
        RECT 65 141.374 65.072 146.014 ; 
        RECT 61.94 141.52 62.084 145.978 ; 
        RECT 61.04 141.52 61.148 145.978 ; 
        RECT 56.36 141.374 56.432 146.014 ; 
        RECT 0.632 141.374 0.704 146.014 ; 
        RECT 120.728 145.694 120.8 150.334 ; 
        RECT 65 145.694 65.072 150.334 ; 
        RECT 61.94 145.84 62.084 150.298 ; 
        RECT 61.04 145.84 61.148 150.298 ; 
        RECT 56.36 145.694 56.432 150.334 ; 
        RECT 0.632 145.694 0.704 150.334 ; 
        RECT 120.728 150.014 120.8 154.654 ; 
        RECT 65 150.014 65.072 154.654 ; 
        RECT 61.94 150.16 62.084 154.618 ; 
        RECT 61.04 150.16 61.148 154.618 ; 
        RECT 56.36 150.014 56.432 154.654 ; 
        RECT 0.632 150.014 0.704 154.654 ; 
        RECT 120.728 154.334 120.8 158.974 ; 
        RECT 65 154.334 65.072 158.974 ; 
        RECT 61.94 154.48 62.084 158.938 ; 
        RECT 61.04 154.48 61.148 158.938 ; 
        RECT 56.36 154.334 56.432 158.974 ; 
        RECT 0.632 154.334 0.704 158.974 ; 
        RECT 120.728 158.654 120.8 163.294 ; 
        RECT 65 158.654 65.072 163.294 ; 
        RECT 61.94 158.8 62.084 163.258 ; 
        RECT 61.04 158.8 61.148 163.258 ; 
        RECT 56.36 158.654 56.432 163.294 ; 
        RECT 0.632 158.654 0.704 163.294 ; 
        RECT 120.728 162.974 120.8 167.614 ; 
        RECT 65 162.974 65.072 167.614 ; 
        RECT 61.94 163.12 62.084 167.578 ; 
        RECT 61.04 163.12 61.148 167.578 ; 
        RECT 56.36 162.974 56.432 167.614 ; 
        RECT 0.632 162.974 0.704 167.614 ; 
        RECT 120.728 167.294 120.8 171.934 ; 
        RECT 65 167.294 65.072 171.934 ; 
        RECT 61.94 167.44 62.084 171.898 ; 
        RECT 61.04 167.44 61.148 171.898 ; 
        RECT 56.36 167.294 56.432 171.934 ; 
        RECT 0.632 167.294 0.704 171.934 ; 
        RECT 120.728 171.614 120.8 176.254 ; 
        RECT 65 171.614 65.072 176.254 ; 
        RECT 61.94 171.76 62.084 176.218 ; 
        RECT 61.04 171.76 61.148 176.218 ; 
        RECT 56.36 171.614 56.432 176.254 ; 
        RECT 0.632 171.614 0.704 176.254 ; 
        RECT 120.728 175.934 120.8 180.574 ; 
        RECT 65 175.934 65.072 180.574 ; 
        RECT 61.94 176.08 62.084 180.538 ; 
        RECT 61.04 176.08 61.148 180.538 ; 
        RECT 56.36 175.934 56.432 180.574 ; 
        RECT 0.632 175.934 0.704 180.574 ; 
        RECT 120.728 180.254 120.8 184.894 ; 
        RECT 65 180.254 65.072 184.894 ; 
        RECT 61.94 180.4 62.084 184.858 ; 
        RECT 61.04 180.4 61.148 184.858 ; 
        RECT 56.36 180.254 56.432 184.894 ; 
        RECT 0.632 180.254 0.704 184.894 ; 
        RECT 120.728 184.574 120.8 189.214 ; 
        RECT 65 184.574 65.072 189.214 ; 
        RECT 61.94 184.72 62.084 189.178 ; 
        RECT 61.04 184.72 61.148 189.178 ; 
        RECT 56.36 184.574 56.432 189.214 ; 
        RECT 0.632 184.574 0.704 189.214 ; 
        RECT 120.728 188.894 120.8 193.534 ; 
        RECT 65 188.894 65.072 193.534 ; 
        RECT 61.94 189.04 62.084 193.498 ; 
        RECT 61.04 189.04 61.148 193.498 ; 
        RECT 56.36 188.894 56.432 193.534 ; 
        RECT 0.632 188.894 0.704 193.534 ; 
        RECT 120.728 193.214 120.8 197.854 ; 
        RECT 65 193.214 65.072 197.854 ; 
        RECT 61.94 193.36 62.084 197.818 ; 
        RECT 61.04 193.36 61.148 197.818 ; 
        RECT 56.36 193.214 56.432 197.854 ; 
        RECT 0.632 193.214 0.704 197.854 ; 
        RECT 120.728 197.534 120.8 202.174 ; 
        RECT 65 197.534 65.072 202.174 ; 
        RECT 61.94 197.68 62.084 202.138 ; 
        RECT 61.04 197.68 61.148 202.138 ; 
        RECT 56.36 197.534 56.432 202.174 ; 
        RECT 0.632 197.534 0.704 202.174 ; 
        RECT 120.728 201.854 120.8 206.494 ; 
        RECT 65 201.854 65.072 206.494 ; 
        RECT 61.94 202 62.084 206.458 ; 
        RECT 61.04 202 61.148 206.458 ; 
        RECT 56.36 201.854 56.432 206.494 ; 
        RECT 0.632 201.854 0.704 206.494 ; 
        RECT 120.728 206.174 120.8 210.814 ; 
        RECT 65 206.174 65.072 210.814 ; 
        RECT 61.94 206.32 62.084 210.778 ; 
        RECT 61.04 206.32 61.148 210.778 ; 
        RECT 56.36 206.174 56.432 210.814 ; 
        RECT 0.632 206.174 0.704 210.814 ; 
        RECT 120.728 210.494 120.8 215.134 ; 
        RECT 65 210.494 65.072 215.134 ; 
        RECT 61.94 210.64 62.084 215.098 ; 
        RECT 61.04 210.64 61.148 215.098 ; 
        RECT 56.36 210.494 56.432 215.134 ; 
        RECT 0.632 210.494 0.704 215.134 ; 
        RECT 120.728 214.814 120.8 219.454 ; 
        RECT 65 214.814 65.072 219.454 ; 
        RECT 61.94 214.96 62.084 219.418 ; 
        RECT 61.04 214.96 61.148 219.418 ; 
        RECT 56.36 214.814 56.432 219.454 ; 
        RECT 0.632 214.814 0.704 219.454 ; 
        RECT 120.728 219.134 120.8 223.774 ; 
        RECT 65 219.134 65.072 223.774 ; 
        RECT 61.94 219.28 62.084 223.738 ; 
        RECT 61.04 219.28 61.148 223.738 ; 
        RECT 56.36 219.134 56.432 223.774 ; 
        RECT 0.632 219.134 0.704 223.774 ; 
        RECT 120.728 223.454 120.8 228.094 ; 
        RECT 65 223.454 65.072 228.094 ; 
        RECT 61.94 223.6 62.084 228.058 ; 
        RECT 61.04 223.6 61.148 228.058 ; 
        RECT 56.36 223.454 56.432 228.094 ; 
        RECT 0.632 223.454 0.704 228.094 ; 
        RECT 120.728 227.774 120.8 232.414 ; 
        RECT 65 227.774 65.072 232.414 ; 
        RECT 61.94 227.92 62.084 232.378 ; 
        RECT 61.04 227.92 61.148 232.378 ; 
        RECT 56.36 227.774 56.432 232.414 ; 
        RECT 0.632 227.774 0.704 232.414 ; 
        RECT 120.728 232.094 120.8 236.734 ; 
        RECT 65 232.094 65.072 236.734 ; 
        RECT 61.94 232.24 62.084 236.698 ; 
        RECT 61.04 232.24 61.148 236.698 ; 
        RECT 56.36 232.094 56.432 236.734 ; 
        RECT 0.632 232.094 0.704 236.734 ; 
        RECT 120.728 236.414 120.8 241.054 ; 
        RECT 65 236.414 65.072 241.054 ; 
        RECT 61.94 236.56 62.084 241.018 ; 
        RECT 61.04 236.56 61.148 241.018 ; 
        RECT 56.36 236.414 56.432 241.054 ; 
        RECT 0.632 236.414 0.704 241.054 ; 
      LAYER V3 ; 
        RECT 0.632 4.304 0.704 4.496 ; 
        RECT 56.36 4.304 56.432 4.496 ; 
        RECT 61.04 4.304 61.148 4.496 ; 
        RECT 61.94 4.304 62.084 4.496 ; 
        RECT 65 4.304 65.072 4.496 ; 
        RECT 120.728 4.304 120.8 4.496 ; 
        RECT 0.632 8.624 0.704 8.816 ; 
        RECT 56.36 8.624 56.432 8.816 ; 
        RECT 61.04 8.624 61.148 8.816 ; 
        RECT 61.94 8.624 62.084 8.816 ; 
        RECT 65 8.624 65.072 8.816 ; 
        RECT 120.728 8.624 120.8 8.816 ; 
        RECT 0.632 12.944 0.704 13.136 ; 
        RECT 56.36 12.944 56.432 13.136 ; 
        RECT 61.04 12.944 61.148 13.136 ; 
        RECT 61.94 12.944 62.084 13.136 ; 
        RECT 65 12.944 65.072 13.136 ; 
        RECT 120.728 12.944 120.8 13.136 ; 
        RECT 0.632 17.264 0.704 17.456 ; 
        RECT 56.36 17.264 56.432 17.456 ; 
        RECT 61.04 17.264 61.148 17.456 ; 
        RECT 61.94 17.264 62.084 17.456 ; 
        RECT 65 17.264 65.072 17.456 ; 
        RECT 120.728 17.264 120.8 17.456 ; 
        RECT 0.632 21.584 0.704 21.776 ; 
        RECT 56.36 21.584 56.432 21.776 ; 
        RECT 61.04 21.584 61.148 21.776 ; 
        RECT 61.94 21.584 62.084 21.776 ; 
        RECT 65 21.584 65.072 21.776 ; 
        RECT 120.728 21.584 120.8 21.776 ; 
        RECT 0.632 25.904 0.704 26.096 ; 
        RECT 56.36 25.904 56.432 26.096 ; 
        RECT 61.04 25.904 61.148 26.096 ; 
        RECT 61.94 25.904 62.084 26.096 ; 
        RECT 65 25.904 65.072 26.096 ; 
        RECT 120.728 25.904 120.8 26.096 ; 
        RECT 0.632 30.224 0.704 30.416 ; 
        RECT 56.36 30.224 56.432 30.416 ; 
        RECT 61.04 30.224 61.148 30.416 ; 
        RECT 61.94 30.224 62.084 30.416 ; 
        RECT 65 30.224 65.072 30.416 ; 
        RECT 120.728 30.224 120.8 30.416 ; 
        RECT 0.632 34.544 0.704 34.736 ; 
        RECT 56.36 34.544 56.432 34.736 ; 
        RECT 61.04 34.544 61.148 34.736 ; 
        RECT 61.94 34.544 62.084 34.736 ; 
        RECT 65 34.544 65.072 34.736 ; 
        RECT 120.728 34.544 120.8 34.736 ; 
        RECT 0.632 38.864 0.704 39.056 ; 
        RECT 56.36 38.864 56.432 39.056 ; 
        RECT 61.04 38.864 61.148 39.056 ; 
        RECT 61.94 38.864 62.084 39.056 ; 
        RECT 65 38.864 65.072 39.056 ; 
        RECT 120.728 38.864 120.8 39.056 ; 
        RECT 0.632 43.184 0.704 43.376 ; 
        RECT 56.36 43.184 56.432 43.376 ; 
        RECT 61.04 43.184 61.148 43.376 ; 
        RECT 61.94 43.184 62.084 43.376 ; 
        RECT 65 43.184 65.072 43.376 ; 
        RECT 120.728 43.184 120.8 43.376 ; 
        RECT 0.632 47.504 0.704 47.696 ; 
        RECT 56.36 47.504 56.432 47.696 ; 
        RECT 61.04 47.504 61.148 47.696 ; 
        RECT 61.94 47.504 62.084 47.696 ; 
        RECT 65 47.504 65.072 47.696 ; 
        RECT 120.728 47.504 120.8 47.696 ; 
        RECT 0.632 51.824 0.704 52.016 ; 
        RECT 56.36 51.824 56.432 52.016 ; 
        RECT 61.04 51.824 61.148 52.016 ; 
        RECT 61.94 51.824 62.084 52.016 ; 
        RECT 65 51.824 65.072 52.016 ; 
        RECT 120.728 51.824 120.8 52.016 ; 
        RECT 0.632 56.144 0.704 56.336 ; 
        RECT 56.36 56.144 56.432 56.336 ; 
        RECT 61.04 56.144 61.148 56.336 ; 
        RECT 61.94 56.144 62.084 56.336 ; 
        RECT 65 56.144 65.072 56.336 ; 
        RECT 120.728 56.144 120.8 56.336 ; 
        RECT 0.632 60.464 0.704 60.656 ; 
        RECT 56.36 60.464 56.432 60.656 ; 
        RECT 61.04 60.464 61.148 60.656 ; 
        RECT 61.94 60.464 62.084 60.656 ; 
        RECT 65 60.464 65.072 60.656 ; 
        RECT 120.728 60.464 120.8 60.656 ; 
        RECT 0.632 64.784 0.704 64.976 ; 
        RECT 56.36 64.784 56.432 64.976 ; 
        RECT 61.04 64.784 61.148 64.976 ; 
        RECT 61.94 64.784 62.084 64.976 ; 
        RECT 65 64.784 65.072 64.976 ; 
        RECT 120.728 64.784 120.8 64.976 ; 
        RECT 0.632 69.104 0.704 69.296 ; 
        RECT 56.36 69.104 56.432 69.296 ; 
        RECT 61.04 69.104 61.148 69.296 ; 
        RECT 61.94 69.104 62.084 69.296 ; 
        RECT 65 69.104 65.072 69.296 ; 
        RECT 120.728 69.104 120.8 69.296 ; 
        RECT 0.632 73.424 0.704 73.616 ; 
        RECT 56.36 73.424 56.432 73.616 ; 
        RECT 61.04 73.424 61.148 73.616 ; 
        RECT 61.94 73.424 62.084 73.616 ; 
        RECT 65 73.424 65.072 73.616 ; 
        RECT 120.728 73.424 120.8 73.616 ; 
        RECT 0.632 77.744 0.704 77.936 ; 
        RECT 56.36 77.744 56.432 77.936 ; 
        RECT 61.04 77.744 61.148 77.936 ; 
        RECT 61.94 77.744 62.084 77.936 ; 
        RECT 65 77.744 65.072 77.936 ; 
        RECT 120.728 77.744 120.8 77.936 ; 
        RECT 0.632 82.064 0.704 82.256 ; 
        RECT 56.36 82.064 56.432 82.256 ; 
        RECT 61.04 82.064 61.148 82.256 ; 
        RECT 61.94 82.064 62.084 82.256 ; 
        RECT 65 82.064 65.072 82.256 ; 
        RECT 120.728 82.064 120.8 82.256 ; 
        RECT 0.632 86.384 0.704 86.576 ; 
        RECT 56.36 86.384 56.432 86.576 ; 
        RECT 61.04 86.384 61.148 86.576 ; 
        RECT 61.94 86.384 62.084 86.576 ; 
        RECT 65 86.384 65.072 86.576 ; 
        RECT 120.728 86.384 120.8 86.576 ; 
        RECT 0.632 90.704 0.704 90.896 ; 
        RECT 56.36 90.704 56.432 90.896 ; 
        RECT 61.04 90.704 61.148 90.896 ; 
        RECT 61.94 90.704 62.084 90.896 ; 
        RECT 65 90.704 65.072 90.896 ; 
        RECT 120.728 90.704 120.8 90.896 ; 
        RECT 0.632 95.024 0.704 95.216 ; 
        RECT 56.36 95.024 56.432 95.216 ; 
        RECT 61.04 95.024 61.148 95.216 ; 
        RECT 61.94 95.024 62.084 95.216 ; 
        RECT 65 95.024 65.072 95.216 ; 
        RECT 120.728 95.024 120.8 95.216 ; 
        RECT 0.632 99.344 0.704 99.536 ; 
        RECT 56.36 99.344 56.432 99.536 ; 
        RECT 61.04 99.344 61.148 99.536 ; 
        RECT 61.94 99.344 62.084 99.536 ; 
        RECT 65 99.344 65.072 99.536 ; 
        RECT 120.728 99.344 120.8 99.536 ; 
        RECT 0.632 103.664 0.704 103.856 ; 
        RECT 56.36 103.664 56.432 103.856 ; 
        RECT 61.04 103.664 61.148 103.856 ; 
        RECT 61.94 103.664 62.084 103.856 ; 
        RECT 65 103.664 65.072 103.856 ; 
        RECT 120.728 103.664 120.8 103.856 ; 
        RECT 56.34 107.926 56.412 108.79 ; 
        RECT 61.18 133.27 61.252 134.134 ; 
        RECT 61.18 120.598 61.252 121.462 ; 
        RECT 61.18 107.926 61.252 108.79 ; 
        RECT 61.388 133.27 61.46 134.134 ; 
        RECT 61.388 120.598 61.46 121.462 ; 
        RECT 61.388 107.926 61.46 108.79 ; 
        RECT 61.596 133.27 61.668 134.134 ; 
        RECT 61.596 120.598 61.668 121.462 ; 
        RECT 61.596 107.926 61.668 108.79 ; 
        RECT 61.804 133.27 61.876 134.134 ; 
        RECT 61.804 120.598 61.876 121.462 ; 
        RECT 61.804 107.926 61.876 108.79 ; 
        RECT 62.012 133.27 62.084 134.134 ; 
        RECT 62.012 120.598 62.084 121.462 ; 
        RECT 62.012 107.926 62.084 108.79 ; 
        RECT 64.98 107.926 65.052 108.79 ; 
        RECT 0.632 140.492 0.704 140.684 ; 
        RECT 56.36 140.492 56.432 140.684 ; 
        RECT 61.04 140.492 61.148 140.684 ; 
        RECT 61.94 140.492 62.084 140.684 ; 
        RECT 65 140.492 65.072 140.684 ; 
        RECT 120.728 140.492 120.8 140.684 ; 
        RECT 0.632 144.812 0.704 145.004 ; 
        RECT 56.36 144.812 56.432 145.004 ; 
        RECT 61.04 144.812 61.148 145.004 ; 
        RECT 61.94 144.812 62.084 145.004 ; 
        RECT 65 144.812 65.072 145.004 ; 
        RECT 120.728 144.812 120.8 145.004 ; 
        RECT 0.632 149.132 0.704 149.324 ; 
        RECT 56.36 149.132 56.432 149.324 ; 
        RECT 61.04 149.132 61.148 149.324 ; 
        RECT 61.94 149.132 62.084 149.324 ; 
        RECT 65 149.132 65.072 149.324 ; 
        RECT 120.728 149.132 120.8 149.324 ; 
        RECT 0.632 153.452 0.704 153.644 ; 
        RECT 56.36 153.452 56.432 153.644 ; 
        RECT 61.04 153.452 61.148 153.644 ; 
        RECT 61.94 153.452 62.084 153.644 ; 
        RECT 65 153.452 65.072 153.644 ; 
        RECT 120.728 153.452 120.8 153.644 ; 
        RECT 0.632 157.772 0.704 157.964 ; 
        RECT 56.36 157.772 56.432 157.964 ; 
        RECT 61.04 157.772 61.148 157.964 ; 
        RECT 61.94 157.772 62.084 157.964 ; 
        RECT 65 157.772 65.072 157.964 ; 
        RECT 120.728 157.772 120.8 157.964 ; 
        RECT 0.632 162.092 0.704 162.284 ; 
        RECT 56.36 162.092 56.432 162.284 ; 
        RECT 61.04 162.092 61.148 162.284 ; 
        RECT 61.94 162.092 62.084 162.284 ; 
        RECT 65 162.092 65.072 162.284 ; 
        RECT 120.728 162.092 120.8 162.284 ; 
        RECT 0.632 166.412 0.704 166.604 ; 
        RECT 56.36 166.412 56.432 166.604 ; 
        RECT 61.04 166.412 61.148 166.604 ; 
        RECT 61.94 166.412 62.084 166.604 ; 
        RECT 65 166.412 65.072 166.604 ; 
        RECT 120.728 166.412 120.8 166.604 ; 
        RECT 0.632 170.732 0.704 170.924 ; 
        RECT 56.36 170.732 56.432 170.924 ; 
        RECT 61.04 170.732 61.148 170.924 ; 
        RECT 61.94 170.732 62.084 170.924 ; 
        RECT 65 170.732 65.072 170.924 ; 
        RECT 120.728 170.732 120.8 170.924 ; 
        RECT 0.632 175.052 0.704 175.244 ; 
        RECT 56.36 175.052 56.432 175.244 ; 
        RECT 61.04 175.052 61.148 175.244 ; 
        RECT 61.94 175.052 62.084 175.244 ; 
        RECT 65 175.052 65.072 175.244 ; 
        RECT 120.728 175.052 120.8 175.244 ; 
        RECT 0.632 179.372 0.704 179.564 ; 
        RECT 56.36 179.372 56.432 179.564 ; 
        RECT 61.04 179.372 61.148 179.564 ; 
        RECT 61.94 179.372 62.084 179.564 ; 
        RECT 65 179.372 65.072 179.564 ; 
        RECT 120.728 179.372 120.8 179.564 ; 
        RECT 0.632 183.692 0.704 183.884 ; 
        RECT 56.36 183.692 56.432 183.884 ; 
        RECT 61.04 183.692 61.148 183.884 ; 
        RECT 61.94 183.692 62.084 183.884 ; 
        RECT 65 183.692 65.072 183.884 ; 
        RECT 120.728 183.692 120.8 183.884 ; 
        RECT 0.632 188.012 0.704 188.204 ; 
        RECT 56.36 188.012 56.432 188.204 ; 
        RECT 61.04 188.012 61.148 188.204 ; 
        RECT 61.94 188.012 62.084 188.204 ; 
        RECT 65 188.012 65.072 188.204 ; 
        RECT 120.728 188.012 120.8 188.204 ; 
        RECT 0.632 192.332 0.704 192.524 ; 
        RECT 56.36 192.332 56.432 192.524 ; 
        RECT 61.04 192.332 61.148 192.524 ; 
        RECT 61.94 192.332 62.084 192.524 ; 
        RECT 65 192.332 65.072 192.524 ; 
        RECT 120.728 192.332 120.8 192.524 ; 
        RECT 0.632 196.652 0.704 196.844 ; 
        RECT 56.36 196.652 56.432 196.844 ; 
        RECT 61.04 196.652 61.148 196.844 ; 
        RECT 61.94 196.652 62.084 196.844 ; 
        RECT 65 196.652 65.072 196.844 ; 
        RECT 120.728 196.652 120.8 196.844 ; 
        RECT 0.632 200.972 0.704 201.164 ; 
        RECT 56.36 200.972 56.432 201.164 ; 
        RECT 61.04 200.972 61.148 201.164 ; 
        RECT 61.94 200.972 62.084 201.164 ; 
        RECT 65 200.972 65.072 201.164 ; 
        RECT 120.728 200.972 120.8 201.164 ; 
        RECT 0.632 205.292 0.704 205.484 ; 
        RECT 56.36 205.292 56.432 205.484 ; 
        RECT 61.04 205.292 61.148 205.484 ; 
        RECT 61.94 205.292 62.084 205.484 ; 
        RECT 65 205.292 65.072 205.484 ; 
        RECT 120.728 205.292 120.8 205.484 ; 
        RECT 0.632 209.612 0.704 209.804 ; 
        RECT 56.36 209.612 56.432 209.804 ; 
        RECT 61.04 209.612 61.148 209.804 ; 
        RECT 61.94 209.612 62.084 209.804 ; 
        RECT 65 209.612 65.072 209.804 ; 
        RECT 120.728 209.612 120.8 209.804 ; 
        RECT 0.632 213.932 0.704 214.124 ; 
        RECT 56.36 213.932 56.432 214.124 ; 
        RECT 61.04 213.932 61.148 214.124 ; 
        RECT 61.94 213.932 62.084 214.124 ; 
        RECT 65 213.932 65.072 214.124 ; 
        RECT 120.728 213.932 120.8 214.124 ; 
        RECT 0.632 218.252 0.704 218.444 ; 
        RECT 56.36 218.252 56.432 218.444 ; 
        RECT 61.04 218.252 61.148 218.444 ; 
        RECT 61.94 218.252 62.084 218.444 ; 
        RECT 65 218.252 65.072 218.444 ; 
        RECT 120.728 218.252 120.8 218.444 ; 
        RECT 0.632 222.572 0.704 222.764 ; 
        RECT 56.36 222.572 56.432 222.764 ; 
        RECT 61.04 222.572 61.148 222.764 ; 
        RECT 61.94 222.572 62.084 222.764 ; 
        RECT 65 222.572 65.072 222.764 ; 
        RECT 120.728 222.572 120.8 222.764 ; 
        RECT 0.632 226.892 0.704 227.084 ; 
        RECT 56.36 226.892 56.432 227.084 ; 
        RECT 61.04 226.892 61.148 227.084 ; 
        RECT 61.94 226.892 62.084 227.084 ; 
        RECT 65 226.892 65.072 227.084 ; 
        RECT 120.728 226.892 120.8 227.084 ; 
        RECT 0.632 231.212 0.704 231.404 ; 
        RECT 56.36 231.212 56.432 231.404 ; 
        RECT 61.04 231.212 61.148 231.404 ; 
        RECT 61.94 231.212 62.084 231.404 ; 
        RECT 65 231.212 65.072 231.404 ; 
        RECT 120.728 231.212 120.8 231.404 ; 
        RECT 0.632 235.532 0.704 235.724 ; 
        RECT 56.36 235.532 56.432 235.724 ; 
        RECT 61.04 235.532 61.148 235.724 ; 
        RECT 61.94 235.532 62.084 235.724 ; 
        RECT 65 235.532 65.072 235.724 ; 
        RECT 120.728 235.532 120.8 235.724 ; 
        RECT 0.632 239.852 0.704 240.044 ; 
        RECT 56.36 239.852 56.432 240.044 ; 
        RECT 61.04 239.852 61.148 240.044 ; 
        RECT 61.94 239.852 62.084 240.044 ; 
        RECT 65 239.852 65.072 240.044 ; 
        RECT 120.728 239.852 120.8 240.044 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 70.812 109.814 70.884 109.962 ; 
      LAYER M4 ; 
        RECT 70.604 109.846 70.94 109.942 ; 
      LAYER M5 ; 
        RECT 70.8 106.042 70.896 119.002 ; 
      LAYER V3 ; 
        RECT 70.812 109.846 70.884 109.942 ; 
      LAYER V4 ; 
        RECT 70.8 109.846 70.896 109.942 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 69.948 109.826 70.02 109.974 ; 
      LAYER M4 ; 
        RECT 69.74 109.846 70.076 109.942 ; 
      LAYER M5 ; 
        RECT 69.936 106.042 70.032 119.002 ; 
      LAYER V3 ; 
        RECT 69.948 109.846 70.02 109.942 ; 
      LAYER V4 ; 
        RECT 69.936 109.846 70.032 109.942 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 69.084 107.51 69.156 107.658 ; 
      LAYER M4 ; 
        RECT 68.876 107.542 69.212 107.638 ; 
      LAYER M5 ; 
        RECT 69.072 106.042 69.168 119.002 ; 
      LAYER V3 ; 
        RECT 69.084 107.542 69.156 107.638 ; 
      LAYER V4 ; 
        RECT 69.072 107.542 69.168 107.638 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 68.22 108.47 68.292 109.194 ; 
      LAYER M4 ; 
        RECT 68.012 109.078 68.348 109.174 ; 
      LAYER M5 ; 
        RECT 68.208 106.042 68.304 119.002 ; 
      LAYER V3 ; 
        RECT 68.22 109.078 68.292 109.174 ; 
      LAYER V4 ; 
        RECT 68.208 109.078 68.304 109.174 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 67.356 107.522 67.428 107.79 ; 
      LAYER M4 ; 
        RECT 67.148 107.542 67.484 107.638 ; 
      LAYER M5 ; 
        RECT 67.344 106.042 67.44 119.002 ; 
      LAYER V3 ; 
        RECT 67.356 107.542 67.428 107.638 ; 
      LAYER V4 ; 
        RECT 67.344 107.542 67.44 107.638 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 66.492 106.454 66.564 107.466 ; 
      LAYER M4 ; 
        RECT 66.284 107.35 66.62 107.446 ; 
      LAYER M5 ; 
        RECT 66.48 106.042 66.576 119.002 ; 
      LAYER V3 ; 
        RECT 66.492 107.35 66.564 107.446 ; 
      LAYER V4 ; 
        RECT 66.48 107.35 66.576 107.446 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 65.628 110.594 65.7 110.742 ; 
      LAYER M4 ; 
        RECT 65.42 110.614 65.756 110.71 ; 
      LAYER M5 ; 
        RECT 65.616 106.042 65.712 119.002 ; 
      LAYER V3 ; 
        RECT 65.628 110.614 65.7 110.71 ; 
      LAYER V4 ; 
        RECT 65.616 110.614 65.712 110.71 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 64.764 109.982 64.836 110.346 ; 
      LAYER M4 ; 
        RECT 64.556 110.23 64.892 110.326 ; 
      LAYER M5 ; 
        RECT 64.752 106.042 64.848 119.002 ; 
      LAYER V3 ; 
        RECT 64.764 110.23 64.836 110.326 ; 
      LAYER V4 ; 
        RECT 64.752 110.23 64.848 110.326 ; 
    END 
  END ADDRESS[7] 
  PIN ADDRESS[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 63.324 108.614 63.396 109.194 ; 
      LAYER M4 ; 
        RECT 63.28 109.078 64.028 109.174 ; 
      LAYER M5 ; 
        RECT 63.888 105.006 63.984 119.002 ; 
      LAYER V3 ; 
        RECT 63.324 109.078 63.396 109.174 ; 
      LAYER V4 ; 
        RECT 63.888 109.078 63.984 109.174 ; 
    END 
  END ADDRESS[8] 
  PIN ADDRESS[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 62.172 107.522 62.244 107.79 ; 
      LAYER M4 ; 
        RECT 61.036 107.542 62.288 107.638 ; 
      LAYER M5 ; 
        RECT 61.08 106.042 61.176 119.002 ; 
      LAYER V3 ; 
        RECT 62.172 107.542 62.244 107.638 ; 
      LAYER V4 ; 
        RECT 61.08 107.542 61.176 107.638 ; 
    END 
  END ADDRESS[9] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.588 106.454 60.66 107.466 ; 
      LAYER M4 ; 
        RECT 59.74 107.35 60.704 107.446 ; 
      LAYER M5 ; 
        RECT 59.784 106.042 59.88 119.002 ; 
      LAYER V3 ; 
        RECT 60.588 107.35 60.66 107.446 ; 
      LAYER V4 ; 
        RECT 59.784 107.35 59.88 107.446 ; 
    END 
  END banksel 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 56.556 110.978 56.628 111.174 ; 
      LAYER M4 ; 
        RECT 56.348 110.998 56.684 111.094 ; 
      LAYER M5 ; 
        RECT 56.544 106.042 56.64 119.002 ; 
      LAYER V3 ; 
        RECT 56.556 110.998 56.628 111.094 ; 
      LAYER V4 ; 
        RECT 56.544 110.998 56.64 111.094 ; 
    END 
  END clk 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 57.42 107.522 57.492 107.79 ; 
      LAYER M4 ; 
        RECT 57.212 107.542 57.548 107.638 ; 
      LAYER M5 ; 
        RECT 57.408 106.042 57.504 119.002 ; 
      LAYER V3 ; 
        RECT 57.42 107.542 57.492 107.638 ; 
      LAYER V4 ; 
        RECT 57.408 107.542 57.504 107.638 ; 
    END 
  END write 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 56.7 106.454 56.772 107.466 ; 
      LAYER M4 ; 
        RECT 55.636 107.35 56.816 107.446 ; 
      LAYER M5 ; 
        RECT 55.68 106.042 55.776 119.002 ; 
      LAYER V3 ; 
        RECT 56.7 107.35 56.772 107.446 ; 
      LAYER V4 ; 
        RECT 55.68 107.35 55.776 107.446 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 54.828 109.814 54.9 109.962 ; 
      LAYER M4 ; 
        RECT 54.62 109.846 54.956 109.942 ; 
      LAYER M5 ; 
        RECT 54.816 106.042 54.912 119.002 ; 
      LAYER V3 ; 
        RECT 54.828 109.846 54.9 109.942 ; 
      LAYER V4 ; 
        RECT 54.816 109.846 54.912 109.942 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 53.964 107.522 54.036 108.438 ; 
      LAYER M4 ; 
        RECT 53.756 107.542 54.092 107.638 ; 
      LAYER M5 ; 
        RECT 53.952 106.042 54.048 119.002 ; 
      LAYER V3 ; 
        RECT 53.964 107.542 54.036 107.638 ; 
      LAYER V4 ; 
        RECT 53.952 107.542 54.048 107.638 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 53.1 106.454 53.172 107.466 ; 
      LAYER M4 ; 
        RECT 52.892 107.35 53.228 107.446 ; 
      LAYER M5 ; 
        RECT 53.088 106.042 53.184 119.002 ; 
      LAYER V3 ; 
        RECT 53.1 107.35 53.172 107.446 ; 
      LAYER V4 ; 
        RECT 53.088 107.35 53.184 107.446 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 52.236 107.51 52.308 107.658 ; 
      LAYER M4 ; 
        RECT 52.028 107.542 52.364 107.638 ; 
      LAYER M5 ; 
        RECT 52.224 106.042 52.32 119.002 ; 
      LAYER V3 ; 
        RECT 52.236 107.542 52.308 107.638 ; 
      LAYER V4 ; 
        RECT 52.224 107.542 52.32 107.638 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 51.372 109.814 51.444 109.962 ; 
      LAYER M4 ; 
        RECT 51.164 109.846 51.5 109.942 ; 
      LAYER M5 ; 
        RECT 51.36 106.042 51.456 119.002 ; 
      LAYER V3 ; 
        RECT 51.372 109.846 51.444 109.942 ; 
      LAYER V4 ; 
        RECT 51.36 109.846 51.456 109.942 ; 
    END 
  END sdel[4] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 61.99 61.868 62.948 ; 
      LAYER M4 ; 
        RECT 59.444 62.192 62.036 62.288 ; 
      LAYER V3 ; 
        RECT 61.796 62.192 61.868 62.288 ; 
    END 
  END dataout[14] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 57.67 61.868 58.628 ; 
      LAYER M4 ; 
        RECT 59.444 57.872 62.036 57.968 ; 
      LAYER V3 ; 
        RECT 61.796 57.872 61.868 57.968 ; 
    END 
  END dataout[13] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 53.35 61.868 54.308 ; 
      LAYER M4 ; 
        RECT 59.444 53.552 62.036 53.648 ; 
      LAYER V3 ; 
        RECT 61.796 53.552 61.868 53.648 ; 
    END 
  END dataout[12] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 49.03 61.868 49.988 ; 
      LAYER M4 ; 
        RECT 59.444 49.232 62.036 49.328 ; 
      LAYER V3 ; 
        RECT 61.796 49.232 61.868 49.328 ; 
    END 
  END dataout[11] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 44.71 61.868 45.668 ; 
      LAYER M4 ; 
        RECT 59.444 44.912 62.036 45.008 ; 
      LAYER V3 ; 
        RECT 61.796 44.912 61.868 45.008 ; 
    END 
  END dataout[10] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 1.51 61.868 2.468 ; 
      LAYER M4 ; 
        RECT 59.444 1.712 62.036 1.808 ; 
      LAYER V3 ; 
        RECT 61.796 1.712 61.868 1.808 ; 
    END 
  END dataout[0] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 66.31 61.868 67.268 ; 
      LAYER M4 ; 
        RECT 59.444 66.512 62.036 66.608 ; 
      LAYER V3 ; 
        RECT 61.796 66.512 61.868 66.608 ; 
    END 
  END dataout[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 70.63 61.868 71.588 ; 
      LAYER M4 ; 
        RECT 59.444 70.832 62.036 70.928 ; 
      LAYER V3 ; 
        RECT 61.796 70.832 61.868 70.928 ; 
    END 
  END dataout[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 74.95 61.868 75.908 ; 
      LAYER M4 ; 
        RECT 59.444 75.152 62.036 75.248 ; 
      LAYER V3 ; 
        RECT 61.796 75.152 61.868 75.248 ; 
    END 
  END dataout[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 79.27 61.868 80.228 ; 
      LAYER M4 ; 
        RECT 59.444 79.472 62.036 79.568 ; 
      LAYER V3 ; 
        RECT 61.796 79.472 61.868 79.568 ; 
    END 
  END dataout[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 83.59 61.868 84.548 ; 
      LAYER M4 ; 
        RECT 59.444 83.792 62.036 83.888 ; 
      LAYER V3 ; 
        RECT 61.796 83.792 61.868 83.888 ; 
    END 
  END dataout[19] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 5.83 61.868 6.788 ; 
      LAYER M4 ; 
        RECT 59.444 6.032 62.036 6.128 ; 
      LAYER V3 ; 
        RECT 61.796 6.032 61.868 6.128 ; 
    END 
  END dataout[1] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 87.91 61.868 88.868 ; 
      LAYER M4 ; 
        RECT 59.444 88.112 62.036 88.208 ; 
      LAYER V3 ; 
        RECT 61.796 88.112 61.868 88.208 ; 
    END 
  END dataout[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 92.23 61.868 93.188 ; 
      LAYER M4 ; 
        RECT 59.444 92.432 62.036 92.528 ; 
      LAYER V3 ; 
        RECT 61.796 92.432 61.868 92.528 ; 
    END 
  END dataout[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 96.55 61.868 97.508 ; 
      LAYER M4 ; 
        RECT 59.444 96.752 62.036 96.848 ; 
      LAYER V3 ; 
        RECT 61.796 96.752 61.868 96.848 ; 
    END 
  END dataout[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 100.87 61.868 101.828 ; 
      LAYER M4 ; 
        RECT 59.444 101.072 62.036 101.168 ; 
      LAYER V3 ; 
        RECT 61.796 101.072 61.868 101.168 ; 
    END 
  END dataout[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 137.698 61.868 138.656 ; 
      LAYER M4 ; 
        RECT 59.444 137.9 62.036 137.996 ; 
      LAYER V3 ; 
        RECT 61.796 137.9 61.868 137.996 ; 
    END 
  END dataout[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 142.018 61.868 142.976 ; 
      LAYER M4 ; 
        RECT 59.444 142.22 62.036 142.316 ; 
      LAYER V3 ; 
        RECT 61.796 142.22 61.868 142.316 ; 
    END 
  END dataout[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 146.338 61.868 147.296 ; 
      LAYER M4 ; 
        RECT 59.444 146.54 62.036 146.636 ; 
      LAYER V3 ; 
        RECT 61.796 146.54 61.868 146.636 ; 
    END 
  END dataout[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 150.658 61.868 151.616 ; 
      LAYER M4 ; 
        RECT 59.444 150.86 62.036 150.956 ; 
      LAYER V3 ; 
        RECT 61.796 150.86 61.868 150.956 ; 
    END 
  END dataout[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 154.978 61.868 155.936 ; 
      LAYER M4 ; 
        RECT 59.444 155.18 62.036 155.276 ; 
      LAYER V3 ; 
        RECT 61.796 155.18 61.868 155.276 ; 
    END 
  END dataout[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 159.298 61.868 160.256 ; 
      LAYER M4 ; 
        RECT 59.444 159.5 62.036 159.596 ; 
      LAYER V3 ; 
        RECT 61.796 159.5 61.868 159.596 ; 
    END 
  END dataout[29] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 10.15 61.868 11.108 ; 
      LAYER M4 ; 
        RECT 59.444 10.352 62.036 10.448 ; 
      LAYER V3 ; 
        RECT 61.796 10.352 61.868 10.448 ; 
    END 
  END dataout[2] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 163.618 61.868 164.576 ; 
      LAYER M4 ; 
        RECT 59.444 163.82 62.036 163.916 ; 
      LAYER V3 ; 
        RECT 61.796 163.82 61.868 163.916 ; 
    END 
  END dataout[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 167.938 61.868 168.896 ; 
      LAYER M4 ; 
        RECT 59.444 168.14 62.036 168.236 ; 
      LAYER V3 ; 
        RECT 61.796 168.14 61.868 168.236 ; 
    END 
  END dataout[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 172.258 61.868 173.216 ; 
      LAYER M4 ; 
        RECT 59.444 172.46 62.036 172.556 ; 
      LAYER V3 ; 
        RECT 61.796 172.46 61.868 172.556 ; 
    END 
  END dataout[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 176.578 61.868 177.536 ; 
      LAYER M4 ; 
        RECT 59.444 176.78 62.036 176.876 ; 
      LAYER V3 ; 
        RECT 61.796 176.78 61.868 176.876 ; 
    END 
  END dataout[33] 
  PIN dataout[34] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 180.898 61.868 181.856 ; 
      LAYER M4 ; 
        RECT 59.444 181.1 62.036 181.196 ; 
      LAYER V3 ; 
        RECT 61.796 181.1 61.868 181.196 ; 
    END 
  END dataout[34] 
  PIN dataout[35] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 185.218 61.868 186.176 ; 
      LAYER M4 ; 
        RECT 59.444 185.42 62.036 185.516 ; 
      LAYER V3 ; 
        RECT 61.796 185.42 61.868 185.516 ; 
    END 
  END dataout[35] 
  PIN dataout[36] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 189.538 61.868 190.496 ; 
      LAYER M4 ; 
        RECT 59.444 189.74 62.036 189.836 ; 
      LAYER V3 ; 
        RECT 61.796 189.74 61.868 189.836 ; 
    END 
  END dataout[36] 
  PIN dataout[37] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 193.858 61.868 194.816 ; 
      LAYER M4 ; 
        RECT 59.444 194.06 62.036 194.156 ; 
      LAYER V3 ; 
        RECT 61.796 194.06 61.868 194.156 ; 
    END 
  END dataout[37] 
  PIN dataout[38] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 198.178 61.868 199.136 ; 
      LAYER M4 ; 
        RECT 59.444 198.38 62.036 198.476 ; 
      LAYER V3 ; 
        RECT 61.796 198.38 61.868 198.476 ; 
    END 
  END dataout[38] 
  PIN dataout[39] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 202.498 61.868 203.456 ; 
      LAYER M4 ; 
        RECT 59.444 202.7 62.036 202.796 ; 
      LAYER V3 ; 
        RECT 61.796 202.7 61.868 202.796 ; 
    END 
  END dataout[39] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 14.47 61.868 15.428 ; 
      LAYER M4 ; 
        RECT 59.444 14.672 62.036 14.768 ; 
      LAYER V3 ; 
        RECT 61.796 14.672 61.868 14.768 ; 
    END 
  END dataout[3] 
  PIN dataout[40] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 206.818 61.868 207.776 ; 
      LAYER M4 ; 
        RECT 59.444 207.02 62.036 207.116 ; 
      LAYER V3 ; 
        RECT 61.796 207.02 61.868 207.116 ; 
    END 
  END dataout[40] 
  PIN dataout[41] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 211.138 61.868 212.096 ; 
      LAYER M4 ; 
        RECT 59.444 211.34 62.036 211.436 ; 
      LAYER V3 ; 
        RECT 61.796 211.34 61.868 211.436 ; 
    END 
  END dataout[41] 
  PIN dataout[42] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 215.458 61.868 216.416 ; 
      LAYER M4 ; 
        RECT 59.444 215.66 62.036 215.756 ; 
      LAYER V3 ; 
        RECT 61.796 215.66 61.868 215.756 ; 
    END 
  END dataout[42] 
  PIN dataout[43] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 219.778 61.868 220.736 ; 
      LAYER M4 ; 
        RECT 59.444 219.98 62.036 220.076 ; 
      LAYER V3 ; 
        RECT 61.796 219.98 61.868 220.076 ; 
    END 
  END dataout[43] 
  PIN dataout[44] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 224.098 61.868 225.056 ; 
      LAYER M4 ; 
        RECT 59.444 224.3 62.036 224.396 ; 
      LAYER V3 ; 
        RECT 61.796 224.3 61.868 224.396 ; 
    END 
  END dataout[44] 
  PIN dataout[45] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 228.418 61.868 229.376 ; 
      LAYER M4 ; 
        RECT 59.444 228.62 62.036 228.716 ; 
      LAYER V3 ; 
        RECT 61.796 228.62 61.868 228.716 ; 
    END 
  END dataout[45] 
  PIN dataout[46] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 232.738 61.868 233.696 ; 
      LAYER M4 ; 
        RECT 59.444 232.94 62.036 233.036 ; 
      LAYER V3 ; 
        RECT 61.796 232.94 61.868 233.036 ; 
    END 
  END dataout[46] 
  PIN dataout[47] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 237.058 61.868 238.016 ; 
      LAYER M4 ; 
        RECT 59.444 237.26 62.036 237.356 ; 
      LAYER V3 ; 
        RECT 61.796 237.26 61.868 237.356 ; 
    END 
  END dataout[47] 
  PIN dataout[48] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[48] 
  PIN dataout[49] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[49] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 18.79 61.868 19.748 ; 
      LAYER M4 ; 
        RECT 59.444 18.992 62.036 19.088 ; 
      LAYER V3 ; 
        RECT 61.796 18.992 61.868 19.088 ; 
    END 
  END dataout[4] 
  PIN dataout[50] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[50] 
  PIN dataout[51] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[51] 
  PIN dataout[52] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[52] 
  PIN dataout[53] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[53] 
  PIN dataout[54] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[54] 
  PIN dataout[55] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[55] 
  PIN dataout[56] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[56] 
  PIN dataout[57] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[57] 
  PIN dataout[58] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[58] 
  PIN dataout[59] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[59] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 23.11 61.868 24.068 ; 
      LAYER M4 ; 
        RECT 59.444 23.312 62.036 23.408 ; 
      LAYER V3 ; 
        RECT 61.796 23.312 61.868 23.408 ; 
    END 
  END dataout[5] 
  PIN dataout[60] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[60] 
  PIN dataout[61] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[61] 
  PIN dataout[62] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[62] 
  PIN dataout[63] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[63] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 27.43 61.868 28.388 ; 
      LAYER M4 ; 
        RECT 59.444 27.632 62.036 27.728 ; 
      LAYER V3 ; 
        RECT 61.796 27.632 61.868 27.728 ; 
    END 
  END dataout[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 31.75 61.868 32.708 ; 
      LAYER M4 ; 
        RECT 59.444 31.952 62.036 32.048 ; 
      LAYER V3 ; 
        RECT 61.796 31.952 61.868 32.048 ; 
    END 
  END dataout[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 36.07 61.868 37.028 ; 
      LAYER M4 ; 
        RECT 59.444 36.272 62.036 36.368 ; 
      LAYER V3 ; 
        RECT 61.796 36.272 61.868 36.368 ; 
    END 
  END dataout[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 40.39 61.868 41.348 ; 
      LAYER M4 ; 
        RECT 59.444 40.592 62.036 40.688 ; 
      LAYER V3 ; 
        RECT 61.796 40.592 61.868 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 1.08 60.968 2.7 ; 
      LAYER M4 ; 
        RECT 59.444 1.328 61.988 1.424 ; 
      LAYER V3 ; 
        RECT 60.896 1.328 60.968 1.424 ; 
    END 
  END wd[0] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 44.28 60.968 45.9 ; 
      LAYER M4 ; 
        RECT 59.444 44.528 61.988 44.624 ; 
      LAYER V3 ; 
        RECT 60.896 44.528 60.968 44.624 ; 
    END 
  END wd[10] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 48.6 60.968 50.22 ; 
      LAYER M4 ; 
        RECT 59.444 48.848 61.988 48.944 ; 
      LAYER V3 ; 
        RECT 60.896 48.848 60.968 48.944 ; 
    END 
  END wd[11] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 52.92 60.968 54.54 ; 
      LAYER M4 ; 
        RECT 59.444 53.168 61.988 53.264 ; 
      LAYER V3 ; 
        RECT 60.896 53.168 60.968 53.264 ; 
    END 
  END wd[12] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 57.24 60.968 58.86 ; 
      LAYER M4 ; 
        RECT 59.444 57.488 61.988 57.584 ; 
      LAYER V3 ; 
        RECT 60.896 57.488 60.968 57.584 ; 
    END 
  END wd[13] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 61.56 60.968 63.18 ; 
      LAYER M4 ; 
        RECT 59.444 61.808 61.988 61.904 ; 
      LAYER V3 ; 
        RECT 60.896 61.808 60.968 61.904 ; 
    END 
  END wd[14] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 65.88 60.968 67.5 ; 
      LAYER M4 ; 
        RECT 59.444 66.128 61.988 66.224 ; 
      LAYER V3 ; 
        RECT 60.896 66.128 60.968 66.224 ; 
    END 
  END wd[15] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 70.2 60.968 71.82 ; 
      LAYER M4 ; 
        RECT 59.444 70.448 61.988 70.544 ; 
      LAYER V3 ; 
        RECT 60.896 70.448 60.968 70.544 ; 
    END 
  END wd[16] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 74.52 60.968 76.14 ; 
      LAYER M4 ; 
        RECT 59.444 74.768 61.988 74.864 ; 
      LAYER V3 ; 
        RECT 60.896 74.768 60.968 74.864 ; 
    END 
  END wd[17] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 78.84 60.968 80.46 ; 
      LAYER M4 ; 
        RECT 59.444 79.088 61.988 79.184 ; 
      LAYER V3 ; 
        RECT 60.896 79.088 60.968 79.184 ; 
    END 
  END wd[18] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 83.16 60.968 84.78 ; 
      LAYER M4 ; 
        RECT 59.444 83.408 61.988 83.504 ; 
      LAYER V3 ; 
        RECT 60.896 83.408 60.968 83.504 ; 
    END 
  END wd[19] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 5.4 60.968 7.02 ; 
      LAYER M4 ; 
        RECT 59.444 5.648 61.988 5.744 ; 
      LAYER V3 ; 
        RECT 60.896 5.648 60.968 5.744 ; 
    END 
  END wd[1] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 87.48 60.968 89.1 ; 
      LAYER M4 ; 
        RECT 59.444 87.728 61.988 87.824 ; 
      LAYER V3 ; 
        RECT 60.896 87.728 60.968 87.824 ; 
    END 
  END wd[20] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 91.8 60.968 93.42 ; 
      LAYER M4 ; 
        RECT 59.444 92.048 61.988 92.144 ; 
      LAYER V3 ; 
        RECT 60.896 92.048 60.968 92.144 ; 
    END 
  END wd[21] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 96.12 60.968 97.74 ; 
      LAYER M4 ; 
        RECT 59.444 96.368 61.988 96.464 ; 
      LAYER V3 ; 
        RECT 60.896 96.368 60.968 96.464 ; 
    END 
  END wd[22] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 100.44 60.968 102.06 ; 
      LAYER M4 ; 
        RECT 59.444 100.688 61.988 100.784 ; 
      LAYER V3 ; 
        RECT 60.896 100.688 60.968 100.784 ; 
    END 
  END wd[23] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 137.268 60.968 138.888 ; 
      LAYER M4 ; 
        RECT 59.444 137.516 61.988 137.612 ; 
      LAYER V3 ; 
        RECT 60.896 137.516 60.968 137.612 ; 
    END 
  END wd[24] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 141.588 60.968 143.208 ; 
      LAYER M4 ; 
        RECT 59.444 141.836 61.988 141.932 ; 
      LAYER V3 ; 
        RECT 60.896 141.836 60.968 141.932 ; 
    END 
  END wd[25] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 145.908 60.968 147.528 ; 
      LAYER M4 ; 
        RECT 59.444 146.156 61.988 146.252 ; 
      LAYER V3 ; 
        RECT 60.896 146.156 60.968 146.252 ; 
    END 
  END wd[26] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 150.228 60.968 151.848 ; 
      LAYER M4 ; 
        RECT 59.444 150.476 61.988 150.572 ; 
      LAYER V3 ; 
        RECT 60.896 150.476 60.968 150.572 ; 
    END 
  END wd[27] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 154.548 60.968 156.168 ; 
      LAYER M4 ; 
        RECT 59.444 154.796 61.988 154.892 ; 
      LAYER V3 ; 
        RECT 60.896 154.796 60.968 154.892 ; 
    END 
  END wd[28] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 158.868 60.968 160.488 ; 
      LAYER M4 ; 
        RECT 59.444 159.116 61.988 159.212 ; 
      LAYER V3 ; 
        RECT 60.896 159.116 60.968 159.212 ; 
    END 
  END wd[29] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 9.72 60.968 11.34 ; 
      LAYER M4 ; 
        RECT 59.444 9.968 61.988 10.064 ; 
      LAYER V3 ; 
        RECT 60.896 9.968 60.968 10.064 ; 
    END 
  END wd[2] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 163.188 60.968 164.808 ; 
      LAYER M4 ; 
        RECT 59.444 163.436 61.988 163.532 ; 
      LAYER V3 ; 
        RECT 60.896 163.436 60.968 163.532 ; 
    END 
  END wd[30] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 167.508 60.968 169.128 ; 
      LAYER M4 ; 
        RECT 59.444 167.756 61.988 167.852 ; 
      LAYER V3 ; 
        RECT 60.896 167.756 60.968 167.852 ; 
    END 
  END wd[31] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 171.828 60.968 173.448 ; 
      LAYER M4 ; 
        RECT 59.444 172.076 61.988 172.172 ; 
      LAYER V3 ; 
        RECT 60.896 172.076 60.968 172.172 ; 
    END 
  END wd[32] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 176.148 60.968 177.768 ; 
      LAYER M4 ; 
        RECT 59.444 176.396 61.988 176.492 ; 
      LAYER V3 ; 
        RECT 60.896 176.396 60.968 176.492 ; 
    END 
  END wd[33] 
  PIN wd[34] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 180.468 60.968 182.088 ; 
      LAYER M4 ; 
        RECT 59.444 180.716 61.988 180.812 ; 
      LAYER V3 ; 
        RECT 60.896 180.716 60.968 180.812 ; 
    END 
  END wd[34] 
  PIN wd[35] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 184.788 60.968 186.408 ; 
      LAYER M4 ; 
        RECT 59.444 185.036 61.988 185.132 ; 
      LAYER V3 ; 
        RECT 60.896 185.036 60.968 185.132 ; 
    END 
  END wd[35] 
  PIN wd[36] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 189.108 60.968 190.728 ; 
      LAYER M4 ; 
        RECT 59.444 189.356 61.988 189.452 ; 
      LAYER V3 ; 
        RECT 60.896 189.356 60.968 189.452 ; 
    END 
  END wd[36] 
  PIN wd[37] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 193.428 60.968 195.048 ; 
      LAYER M4 ; 
        RECT 59.444 193.676 61.988 193.772 ; 
      LAYER V3 ; 
        RECT 60.896 193.676 60.968 193.772 ; 
    END 
  END wd[37] 
  PIN wd[38] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 197.748 60.968 199.368 ; 
      LAYER M4 ; 
        RECT 59.444 197.996 61.988 198.092 ; 
      LAYER V3 ; 
        RECT 60.896 197.996 60.968 198.092 ; 
    END 
  END wd[38] 
  PIN wd[39] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 202.068 60.968 203.688 ; 
      LAYER M4 ; 
        RECT 59.444 202.316 61.988 202.412 ; 
      LAYER V3 ; 
        RECT 60.896 202.316 60.968 202.412 ; 
    END 
  END wd[39] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 14.04 60.968 15.66 ; 
      LAYER M4 ; 
        RECT 59.444 14.288 61.988 14.384 ; 
      LAYER V3 ; 
        RECT 60.896 14.288 60.968 14.384 ; 
    END 
  END wd[3] 
  PIN wd[40] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 206.388 60.968 208.008 ; 
      LAYER M4 ; 
        RECT 59.444 206.636 61.988 206.732 ; 
      LAYER V3 ; 
        RECT 60.896 206.636 60.968 206.732 ; 
    END 
  END wd[40] 
  PIN wd[41] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 210.708 60.968 212.328 ; 
      LAYER M4 ; 
        RECT 59.444 210.956 61.988 211.052 ; 
      LAYER V3 ; 
        RECT 60.896 210.956 60.968 211.052 ; 
    END 
  END wd[41] 
  PIN wd[42] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 215.028 60.968 216.648 ; 
      LAYER M4 ; 
        RECT 59.444 215.276 61.988 215.372 ; 
      LAYER V3 ; 
        RECT 60.896 215.276 60.968 215.372 ; 
    END 
  END wd[42] 
  PIN wd[43] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 219.348 60.968 220.968 ; 
      LAYER M4 ; 
        RECT 59.444 219.596 61.988 219.692 ; 
      LAYER V3 ; 
        RECT 60.896 219.596 60.968 219.692 ; 
    END 
  END wd[43] 
  PIN wd[44] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 223.668 60.968 225.288 ; 
      LAYER M4 ; 
        RECT 59.444 223.916 61.988 224.012 ; 
      LAYER V3 ; 
        RECT 60.896 223.916 60.968 224.012 ; 
    END 
  END wd[44] 
  PIN wd[45] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 227.988 60.968 229.608 ; 
      LAYER M4 ; 
        RECT 59.444 228.236 61.988 228.332 ; 
      LAYER V3 ; 
        RECT 60.896 228.236 60.968 228.332 ; 
    END 
  END wd[45] 
  PIN wd[46] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 232.308 60.968 233.928 ; 
      LAYER M4 ; 
        RECT 59.444 232.556 61.988 232.652 ; 
      LAYER V3 ; 
        RECT 60.896 232.556 60.968 232.652 ; 
    END 
  END wd[46] 
  PIN wd[47] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 236.628 60.968 238.248 ; 
      LAYER M4 ; 
        RECT 59.444 236.876 61.988 236.972 ; 
      LAYER V3 ; 
        RECT 60.896 236.876 60.968 236.972 ; 
    END 
  END wd[47] 
  PIN wd[48] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[48] 
  PIN wd[49] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[49] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 18.36 60.968 19.98 ; 
      LAYER M4 ; 
        RECT 59.444 18.608 61.988 18.704 ; 
      LAYER V3 ; 
        RECT 60.896 18.608 60.968 18.704 ; 
    END 
  END wd[4] 
  PIN wd[50] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[50] 
  PIN wd[51] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[51] 
  PIN wd[52] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[52] 
  PIN wd[53] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[53] 
  PIN wd[54] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[54] 
  PIN wd[55] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[55] 
  PIN wd[56] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[56] 
  PIN wd[57] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[57] 
  PIN wd[58] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[58] 
  PIN wd[59] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[59] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 22.68 60.968 24.3 ; 
      LAYER M4 ; 
        RECT 59.444 22.928 61.988 23.024 ; 
      LAYER V3 ; 
        RECT 60.896 22.928 60.968 23.024 ; 
    END 
  END wd[5] 
  PIN wd[60] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[60] 
  PIN wd[61] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[61] 
  PIN wd[62] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[62] 
  PIN wd[63] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[63] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 27 60.968 28.62 ; 
      LAYER M4 ; 
        RECT 59.444 27.248 61.988 27.344 ; 
      LAYER V3 ; 
        RECT 60.896 27.248 60.968 27.344 ; 
    END 
  END wd[6] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 31.32 60.968 32.94 ; 
      LAYER M4 ; 
        RECT 59.444 31.568 61.988 31.664 ; 
      LAYER V3 ; 
        RECT 60.896 31.568 60.968 31.664 ; 
    END 
  END wd[7] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 35.64 60.968 37.26 ; 
      LAYER M4 ; 
        RECT 59.444 35.888 61.988 35.984 ; 
      LAYER V3 ; 
        RECT 60.896 35.888 60.968 35.984 ; 
    END 
  END wd[8] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 39.96 60.968 41.58 ; 
      LAYER M4 ; 
        RECT 59.444 40.208 61.988 40.304 ; 
      LAYER V3 ; 
        RECT 60.896 40.208 60.968 40.304 ; 
    END 
  END wd[9] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0.02 39.906 121.412 44.28 ; 
      RECT 0.02 44.226 121.412 48.6 ; 
      RECT 0.02 48.546 121.412 52.92 ; 
      RECT 0.02 52.866 121.412 57.24 ; 
      RECT 0.02 57.186 121.412 61.56 ; 
      RECT 0.02 61.506 121.412 65.88 ; 
      RECT 0.02 65.826 121.412 70.2 ; 
      RECT 0.02 70.146 121.412 74.52 ; 
      RECT 0.02 74.466 121.412 78.84 ; 
      RECT 0.02 78.786 121.412 83.16 ; 
      RECT 0.02 83.106 121.412 87.48 ; 
      RECT 0.02 87.426 121.412 91.8 ; 
      RECT 0.02 91.746 121.412 96.12 ; 
      RECT 0.02 96.066 121.412 100.44 ; 
      RECT 0.02 100.386 121.412 104.76 ; 
      RECT 0 104.854 121.392 139.468 ; 
        RECT 0.02 137.214 121.412 141.588 ; 
        RECT 0.02 141.534 121.412 145.908 ; 
        RECT 0.02 145.854 121.412 150.228 ; 
        RECT 0.02 150.174 121.412 154.548 ; 
        RECT 0.02 154.494 121.412 158.868 ; 
        RECT 0.02 158.814 121.412 163.188 ; 
        RECT 0.02 163.134 121.412 167.508 ; 
        RECT 0.02 167.454 121.412 171.828 ; 
        RECT 0.02 171.774 121.412 176.148 ; 
        RECT 0.02 176.094 121.412 180.468 ; 
        RECT 0.02 180.414 121.412 184.788 ; 
        RECT 0.02 184.734 121.412 189.108 ; 
        RECT 0.02 189.054 121.412 193.428 ; 
        RECT 0.02 193.374 121.412 197.748 ; 
        RECT 0.02 197.694 121.412 202.068 ; 
        RECT 0.02 202.014 121.412 206.388 ; 
        RECT 0.02 206.334 121.412 210.708 ; 
        RECT 0.02 210.654 121.412 215.028 ; 
        RECT 0.02 214.974 121.412 219.348 ; 
        RECT 0.02 219.294 121.412 223.668 ; 
        RECT 0.02 223.614 121.412 227.988 ; 
        RECT 0.02 227.934 121.412 232.308 ; 
        RECT 0.02 232.254 121.412 236.628 ; 
        RECT 0.02 236.574 121.412 240.948 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0.02 39.906 121.412 44.28 ; 
      RECT 0.02 44.226 121.412 48.6 ; 
      RECT 0.02 48.546 121.412 52.92 ; 
      RECT 0.02 52.866 121.412 57.24 ; 
      RECT 0.02 57.186 121.412 61.56 ; 
      RECT 0.02 61.506 121.412 65.88 ; 
      RECT 0.02 65.826 121.412 70.2 ; 
      RECT 0.02 70.146 121.412 74.52 ; 
      RECT 0.02 74.466 121.412 78.84 ; 
      RECT 0.02 78.786 121.412 83.16 ; 
      RECT 0.02 83.106 121.412 87.48 ; 
      RECT 0.02 87.426 121.412 91.8 ; 
      RECT 0.02 91.746 121.412 96.12 ; 
      RECT 0.02 96.066 121.412 100.44 ; 
      RECT 0.02 100.386 121.412 104.76 ; 
      RECT 0 104.854 121.392 139.468 ; 
        RECT 0.02 137.214 121.412 141.588 ; 
        RECT 0.02 141.534 121.412 145.908 ; 
        RECT 0.02 145.854 121.412 150.228 ; 
        RECT 0.02 150.174 121.412 154.548 ; 
        RECT 0.02 154.494 121.412 158.868 ; 
        RECT 0.02 158.814 121.412 163.188 ; 
        RECT 0.02 163.134 121.412 167.508 ; 
        RECT 0.02 167.454 121.412 171.828 ; 
        RECT 0.02 171.774 121.412 176.148 ; 
        RECT 0.02 176.094 121.412 180.468 ; 
        RECT 0.02 180.414 121.412 184.788 ; 
        RECT 0.02 184.734 121.412 189.108 ; 
        RECT 0.02 189.054 121.412 193.428 ; 
        RECT 0.02 193.374 121.412 197.748 ; 
        RECT 0.02 197.694 121.412 202.068 ; 
        RECT 0.02 202.014 121.412 206.388 ; 
        RECT 0.02 206.334 121.412 210.708 ; 
        RECT 0.02 210.654 121.412 215.028 ; 
        RECT 0.02 214.974 121.412 219.348 ; 
        RECT 0.02 219.294 121.412 223.668 ; 
        RECT 0.02 223.614 121.412 227.988 ; 
        RECT 0.02 227.934 121.412 232.308 ; 
        RECT 0.02 232.254 121.412 236.628 ; 
        RECT 0.02 236.574 121.412 240.948 ; 
  LAYER V1 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0.02 39.906 121.412 44.28 ; 
      RECT 0.02 44.226 121.412 48.6 ; 
      RECT 0.02 48.546 121.412 52.92 ; 
      RECT 0.02 52.866 121.412 57.24 ; 
      RECT 0.02 57.186 121.412 61.56 ; 
      RECT 0.02 61.506 121.412 65.88 ; 
      RECT 0.02 65.826 121.412 70.2 ; 
      RECT 0.02 70.146 121.412 74.52 ; 
      RECT 0.02 74.466 121.412 78.84 ; 
      RECT 0.02 78.786 121.412 83.16 ; 
      RECT 0.02 83.106 121.412 87.48 ; 
      RECT 0.02 87.426 121.412 91.8 ; 
      RECT 0.02 91.746 121.412 96.12 ; 
      RECT 0.02 96.066 121.412 100.44 ; 
      RECT 0.02 100.386 121.412 104.76 ; 
      RECT 0 104.854 121.392 139.468 ; 
        RECT 0.02 137.214 121.412 141.588 ; 
        RECT 0.02 141.534 121.412 145.908 ; 
        RECT 0.02 145.854 121.412 150.228 ; 
        RECT 0.02 150.174 121.412 154.548 ; 
        RECT 0.02 154.494 121.412 158.868 ; 
        RECT 0.02 158.814 121.412 163.188 ; 
        RECT 0.02 163.134 121.412 167.508 ; 
        RECT 0.02 167.454 121.412 171.828 ; 
        RECT 0.02 171.774 121.412 176.148 ; 
        RECT 0.02 176.094 121.412 180.468 ; 
        RECT 0.02 180.414 121.412 184.788 ; 
        RECT 0.02 184.734 121.412 189.108 ; 
        RECT 0.02 189.054 121.412 193.428 ; 
        RECT 0.02 193.374 121.412 197.748 ; 
        RECT 0.02 197.694 121.412 202.068 ; 
        RECT 0.02 202.014 121.412 206.388 ; 
        RECT 0.02 206.334 121.412 210.708 ; 
        RECT 0.02 210.654 121.412 215.028 ; 
        RECT 0.02 214.974 121.412 219.348 ; 
        RECT 0.02 219.294 121.412 223.668 ; 
        RECT 0.02 223.614 121.412 227.988 ; 
        RECT 0.02 227.934 121.412 232.308 ; 
        RECT 0.02 232.254 121.412 236.628 ; 
        RECT 0.02 236.574 121.412 240.948 ; 
  LAYER V2 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0.02 39.906 121.412 44.28 ; 
      RECT 0.02 44.226 121.412 48.6 ; 
      RECT 0.02 48.546 121.412 52.92 ; 
      RECT 0.02 52.866 121.412 57.24 ; 
      RECT 0.02 57.186 121.412 61.56 ; 
      RECT 0.02 61.506 121.412 65.88 ; 
      RECT 0.02 65.826 121.412 70.2 ; 
      RECT 0.02 70.146 121.412 74.52 ; 
      RECT 0.02 74.466 121.412 78.84 ; 
      RECT 0.02 78.786 121.412 83.16 ; 
      RECT 0.02 83.106 121.412 87.48 ; 
      RECT 0.02 87.426 121.412 91.8 ; 
      RECT 0.02 91.746 121.412 96.12 ; 
      RECT 0.02 96.066 121.412 100.44 ; 
      RECT 0.02 100.386 121.412 104.76 ; 
      RECT 0 104.854 121.392 139.468 ; 
        RECT 0.02 137.214 121.412 141.588 ; 
        RECT 0.02 141.534 121.412 145.908 ; 
        RECT 0.02 145.854 121.412 150.228 ; 
        RECT 0.02 150.174 121.412 154.548 ; 
        RECT 0.02 154.494 121.412 158.868 ; 
        RECT 0.02 158.814 121.412 163.188 ; 
        RECT 0.02 163.134 121.412 167.508 ; 
        RECT 0.02 167.454 121.412 171.828 ; 
        RECT 0.02 171.774 121.412 176.148 ; 
        RECT 0.02 176.094 121.412 180.468 ; 
        RECT 0.02 180.414 121.412 184.788 ; 
        RECT 0.02 184.734 121.412 189.108 ; 
        RECT 0.02 189.054 121.412 193.428 ; 
        RECT 0.02 193.374 121.412 197.748 ; 
        RECT 0.02 197.694 121.412 202.068 ; 
        RECT 0.02 202.014 121.412 206.388 ; 
        RECT 0.02 206.334 121.412 210.708 ; 
        RECT 0.02 210.654 121.412 215.028 ; 
        RECT 0.02 214.974 121.412 219.348 ; 
        RECT 0.02 219.294 121.412 223.668 ; 
        RECT 0.02 223.614 121.412 227.988 ; 
        RECT 0.02 227.934 121.412 232.308 ; 
        RECT 0.02 232.254 121.412 236.628 ; 
        RECT 0.02 236.574 121.412 240.948 ; 
  LAYER M3 ; 
      RECT 62.444 1.38 62.516 5.122 ; 
      RECT 62.3 1.38 62.372 5.122 ; 
      RECT 62.156 3.688 62.228 4.978 ; 
      RECT 61.688 4.476 61.76 4.914 ; 
      RECT 61.652 1.51 61.724 2.468 ; 
      RECT 61.508 3.834 61.58 4.448 ; 
      RECT 61.184 3.936 61.256 4.968 ; 
      RECT 59.024 1.38 59.096 5.122 ; 
      RECT 58.88 1.38 58.952 5.122 ; 
      RECT 58.736 2.104 58.808 4.376 ; 
      RECT 62.444 5.7 62.516 9.442 ; 
      RECT 62.3 5.7 62.372 9.442 ; 
      RECT 62.156 8.008 62.228 9.298 ; 
      RECT 61.688 8.796 61.76 9.234 ; 
      RECT 61.652 5.83 61.724 6.788 ; 
      RECT 61.508 8.154 61.58 8.768 ; 
      RECT 61.184 8.256 61.256 9.288 ; 
      RECT 59.024 5.7 59.096 9.442 ; 
      RECT 58.88 5.7 58.952 9.442 ; 
      RECT 58.736 6.424 58.808 8.696 ; 
      RECT 62.444 10.02 62.516 13.762 ; 
      RECT 62.3 10.02 62.372 13.762 ; 
      RECT 62.156 12.328 62.228 13.618 ; 
      RECT 61.688 13.116 61.76 13.554 ; 
      RECT 61.652 10.15 61.724 11.108 ; 
      RECT 61.508 12.474 61.58 13.088 ; 
      RECT 61.184 12.576 61.256 13.608 ; 
      RECT 59.024 10.02 59.096 13.762 ; 
      RECT 58.88 10.02 58.952 13.762 ; 
      RECT 58.736 10.744 58.808 13.016 ; 
      RECT 62.444 14.34 62.516 18.082 ; 
      RECT 62.3 14.34 62.372 18.082 ; 
      RECT 62.156 16.648 62.228 17.938 ; 
      RECT 61.688 17.436 61.76 17.874 ; 
      RECT 61.652 14.47 61.724 15.428 ; 
      RECT 61.508 16.794 61.58 17.408 ; 
      RECT 61.184 16.896 61.256 17.928 ; 
      RECT 59.024 14.34 59.096 18.082 ; 
      RECT 58.88 14.34 58.952 18.082 ; 
      RECT 58.736 15.064 58.808 17.336 ; 
      RECT 62.444 18.66 62.516 22.402 ; 
      RECT 62.3 18.66 62.372 22.402 ; 
      RECT 62.156 20.968 62.228 22.258 ; 
      RECT 61.688 21.756 61.76 22.194 ; 
      RECT 61.652 18.79 61.724 19.748 ; 
      RECT 61.508 21.114 61.58 21.728 ; 
      RECT 61.184 21.216 61.256 22.248 ; 
      RECT 59.024 18.66 59.096 22.402 ; 
      RECT 58.88 18.66 58.952 22.402 ; 
      RECT 58.736 19.384 58.808 21.656 ; 
      RECT 62.444 22.98 62.516 26.722 ; 
      RECT 62.3 22.98 62.372 26.722 ; 
      RECT 62.156 25.288 62.228 26.578 ; 
      RECT 61.688 26.076 61.76 26.514 ; 
      RECT 61.652 23.11 61.724 24.068 ; 
      RECT 61.508 25.434 61.58 26.048 ; 
      RECT 61.184 25.536 61.256 26.568 ; 
      RECT 59.024 22.98 59.096 26.722 ; 
      RECT 58.88 22.98 58.952 26.722 ; 
      RECT 58.736 23.704 58.808 25.976 ; 
      RECT 62.444 27.3 62.516 31.042 ; 
      RECT 62.3 27.3 62.372 31.042 ; 
      RECT 62.156 29.608 62.228 30.898 ; 
      RECT 61.688 30.396 61.76 30.834 ; 
      RECT 61.652 27.43 61.724 28.388 ; 
      RECT 61.508 29.754 61.58 30.368 ; 
      RECT 61.184 29.856 61.256 30.888 ; 
      RECT 59.024 27.3 59.096 31.042 ; 
      RECT 58.88 27.3 58.952 31.042 ; 
      RECT 58.736 28.024 58.808 30.296 ; 
      RECT 62.444 31.62 62.516 35.362 ; 
      RECT 62.3 31.62 62.372 35.362 ; 
      RECT 62.156 33.928 62.228 35.218 ; 
      RECT 61.688 34.716 61.76 35.154 ; 
      RECT 61.652 31.75 61.724 32.708 ; 
      RECT 61.508 34.074 61.58 34.688 ; 
      RECT 61.184 34.176 61.256 35.208 ; 
      RECT 59.024 31.62 59.096 35.362 ; 
      RECT 58.88 31.62 58.952 35.362 ; 
      RECT 58.736 32.344 58.808 34.616 ; 
      RECT 62.444 35.94 62.516 39.682 ; 
      RECT 62.3 35.94 62.372 39.682 ; 
      RECT 62.156 38.248 62.228 39.538 ; 
      RECT 61.688 39.036 61.76 39.474 ; 
      RECT 61.652 36.07 61.724 37.028 ; 
      RECT 61.508 38.394 61.58 39.008 ; 
      RECT 61.184 38.496 61.256 39.528 ; 
      RECT 59.024 35.94 59.096 39.682 ; 
      RECT 58.88 35.94 58.952 39.682 ; 
      RECT 58.736 36.664 58.808 38.936 ; 
      RECT 62.444 40.26 62.516 44.002 ; 
      RECT 62.3 40.26 62.372 44.002 ; 
      RECT 62.156 42.568 62.228 43.858 ; 
      RECT 61.688 43.356 61.76 43.794 ; 
      RECT 61.652 40.39 61.724 41.348 ; 
      RECT 61.508 42.714 61.58 43.328 ; 
      RECT 61.184 42.816 61.256 43.848 ; 
      RECT 59.024 40.26 59.096 44.002 ; 
      RECT 58.88 40.26 58.952 44.002 ; 
      RECT 58.736 40.984 58.808 43.256 ; 
      RECT 62.444 44.58 62.516 48.322 ; 
      RECT 62.3 44.58 62.372 48.322 ; 
      RECT 62.156 46.888 62.228 48.178 ; 
      RECT 61.688 47.676 61.76 48.114 ; 
      RECT 61.652 44.71 61.724 45.668 ; 
      RECT 61.508 47.034 61.58 47.648 ; 
      RECT 61.184 47.136 61.256 48.168 ; 
      RECT 59.024 44.58 59.096 48.322 ; 
      RECT 58.88 44.58 58.952 48.322 ; 
      RECT 58.736 45.304 58.808 47.576 ; 
      RECT 62.444 48.9 62.516 52.642 ; 
      RECT 62.3 48.9 62.372 52.642 ; 
      RECT 62.156 51.208 62.228 52.498 ; 
      RECT 61.688 51.996 61.76 52.434 ; 
      RECT 61.652 49.03 61.724 49.988 ; 
      RECT 61.508 51.354 61.58 51.968 ; 
      RECT 61.184 51.456 61.256 52.488 ; 
      RECT 59.024 48.9 59.096 52.642 ; 
      RECT 58.88 48.9 58.952 52.642 ; 
      RECT 58.736 49.624 58.808 51.896 ; 
      RECT 62.444 53.22 62.516 56.962 ; 
      RECT 62.3 53.22 62.372 56.962 ; 
      RECT 62.156 55.528 62.228 56.818 ; 
      RECT 61.688 56.316 61.76 56.754 ; 
      RECT 61.652 53.35 61.724 54.308 ; 
      RECT 61.508 55.674 61.58 56.288 ; 
      RECT 61.184 55.776 61.256 56.808 ; 
      RECT 59.024 53.22 59.096 56.962 ; 
      RECT 58.88 53.22 58.952 56.962 ; 
      RECT 58.736 53.944 58.808 56.216 ; 
      RECT 62.444 57.54 62.516 61.282 ; 
      RECT 62.3 57.54 62.372 61.282 ; 
      RECT 62.156 59.848 62.228 61.138 ; 
      RECT 61.688 60.636 61.76 61.074 ; 
      RECT 61.652 57.67 61.724 58.628 ; 
      RECT 61.508 59.994 61.58 60.608 ; 
      RECT 61.184 60.096 61.256 61.128 ; 
      RECT 59.024 57.54 59.096 61.282 ; 
      RECT 58.88 57.54 58.952 61.282 ; 
      RECT 58.736 58.264 58.808 60.536 ; 
      RECT 62.444 61.86 62.516 65.602 ; 
      RECT 62.3 61.86 62.372 65.602 ; 
      RECT 62.156 64.168 62.228 65.458 ; 
      RECT 61.688 64.956 61.76 65.394 ; 
      RECT 61.652 61.99 61.724 62.948 ; 
      RECT 61.508 64.314 61.58 64.928 ; 
      RECT 61.184 64.416 61.256 65.448 ; 
      RECT 59.024 61.86 59.096 65.602 ; 
      RECT 58.88 61.86 58.952 65.602 ; 
      RECT 58.736 62.584 58.808 64.856 ; 
      RECT 62.444 66.18 62.516 69.922 ; 
      RECT 62.3 66.18 62.372 69.922 ; 
      RECT 62.156 68.488 62.228 69.778 ; 
      RECT 61.688 69.276 61.76 69.714 ; 
      RECT 61.652 66.31 61.724 67.268 ; 
      RECT 61.508 68.634 61.58 69.248 ; 
      RECT 61.184 68.736 61.256 69.768 ; 
      RECT 59.024 66.18 59.096 69.922 ; 
      RECT 58.88 66.18 58.952 69.922 ; 
      RECT 58.736 66.904 58.808 69.176 ; 
      RECT 62.444 70.5 62.516 74.242 ; 
      RECT 62.3 70.5 62.372 74.242 ; 
      RECT 62.156 72.808 62.228 74.098 ; 
      RECT 61.688 73.596 61.76 74.034 ; 
      RECT 61.652 70.63 61.724 71.588 ; 
      RECT 61.508 72.954 61.58 73.568 ; 
      RECT 61.184 73.056 61.256 74.088 ; 
      RECT 59.024 70.5 59.096 74.242 ; 
      RECT 58.88 70.5 58.952 74.242 ; 
      RECT 58.736 71.224 58.808 73.496 ; 
      RECT 62.444 74.82 62.516 78.562 ; 
      RECT 62.3 74.82 62.372 78.562 ; 
      RECT 62.156 77.128 62.228 78.418 ; 
      RECT 61.688 77.916 61.76 78.354 ; 
      RECT 61.652 74.95 61.724 75.908 ; 
      RECT 61.508 77.274 61.58 77.888 ; 
      RECT 61.184 77.376 61.256 78.408 ; 
      RECT 59.024 74.82 59.096 78.562 ; 
      RECT 58.88 74.82 58.952 78.562 ; 
      RECT 58.736 75.544 58.808 77.816 ; 
      RECT 62.444 79.14 62.516 82.882 ; 
      RECT 62.3 79.14 62.372 82.882 ; 
      RECT 62.156 81.448 62.228 82.738 ; 
      RECT 61.688 82.236 61.76 82.674 ; 
      RECT 61.652 79.27 61.724 80.228 ; 
      RECT 61.508 81.594 61.58 82.208 ; 
      RECT 61.184 81.696 61.256 82.728 ; 
      RECT 59.024 79.14 59.096 82.882 ; 
      RECT 58.88 79.14 58.952 82.882 ; 
      RECT 58.736 79.864 58.808 82.136 ; 
      RECT 62.444 83.46 62.516 87.202 ; 
      RECT 62.3 83.46 62.372 87.202 ; 
      RECT 62.156 85.768 62.228 87.058 ; 
      RECT 61.688 86.556 61.76 86.994 ; 
      RECT 61.652 83.59 61.724 84.548 ; 
      RECT 61.508 85.914 61.58 86.528 ; 
      RECT 61.184 86.016 61.256 87.048 ; 
      RECT 59.024 83.46 59.096 87.202 ; 
      RECT 58.88 83.46 58.952 87.202 ; 
      RECT 58.736 84.184 58.808 86.456 ; 
      RECT 62.444 87.78 62.516 91.522 ; 
      RECT 62.3 87.78 62.372 91.522 ; 
      RECT 62.156 90.088 62.228 91.378 ; 
      RECT 61.688 90.876 61.76 91.314 ; 
      RECT 61.652 87.91 61.724 88.868 ; 
      RECT 61.508 90.234 61.58 90.848 ; 
      RECT 61.184 90.336 61.256 91.368 ; 
      RECT 59.024 87.78 59.096 91.522 ; 
      RECT 58.88 87.78 58.952 91.522 ; 
      RECT 58.736 88.504 58.808 90.776 ; 
      RECT 62.444 92.1 62.516 95.842 ; 
      RECT 62.3 92.1 62.372 95.842 ; 
      RECT 62.156 94.408 62.228 95.698 ; 
      RECT 61.688 95.196 61.76 95.634 ; 
      RECT 61.652 92.23 61.724 93.188 ; 
      RECT 61.508 94.554 61.58 95.168 ; 
      RECT 61.184 94.656 61.256 95.688 ; 
      RECT 59.024 92.1 59.096 95.842 ; 
      RECT 58.88 92.1 58.952 95.842 ; 
      RECT 58.736 92.824 58.808 95.096 ; 
      RECT 62.444 96.42 62.516 100.162 ; 
      RECT 62.3 96.42 62.372 100.162 ; 
      RECT 62.156 98.728 62.228 100.018 ; 
      RECT 61.688 99.516 61.76 99.954 ; 
      RECT 61.652 96.55 61.724 97.508 ; 
      RECT 61.508 98.874 61.58 99.488 ; 
      RECT 61.184 98.976 61.256 100.008 ; 
      RECT 59.024 96.42 59.096 100.162 ; 
      RECT 58.88 96.42 58.952 100.162 ; 
      RECT 58.736 97.144 58.808 99.416 ; 
      RECT 62.444 100.74 62.516 104.482 ; 
      RECT 62.3 100.74 62.372 104.482 ; 
      RECT 62.156 103.048 62.228 104.338 ; 
      RECT 61.688 103.836 61.76 104.274 ; 
      RECT 61.652 100.87 61.724 101.828 ; 
      RECT 61.508 103.194 61.58 103.808 ; 
      RECT 61.184 103.296 61.256 104.328 ; 
      RECT 59.024 100.74 59.096 104.482 ; 
      RECT 58.88 100.74 58.952 104.482 ; 
      RECT 58.736 101.464 58.808 103.736 ; 
      RECT 120.852 104.094 120.924 137.576 ; 
      RECT 120.708 104.094 120.78 137.576 ; 
      RECT 120.276 104.094 120.348 119.058 ; 
      RECT 119.844 104.094 119.916 119.058 ; 
      RECT 119.412 104.094 119.484 119.058 ; 
      RECT 118.98 104.094 119.052 119.058 ; 
      RECT 118.548 104.094 118.62 119.058 ; 
      RECT 118.116 104.094 118.188 119.058 ; 
      RECT 117.684 104.094 117.756 119.058 ; 
      RECT 117.252 104.094 117.324 119.058 ; 
      RECT 116.82 104.094 116.892 119.058 ; 
      RECT 116.388 104.094 116.46 119.058 ; 
      RECT 115.956 104.094 116.028 119.058 ; 
      RECT 115.524 104.094 115.596 119.058 ; 
      RECT 115.092 104.094 115.164 119.058 ; 
      RECT 114.66 104.094 114.732 119.058 ; 
      RECT 114.228 104.094 114.3 119.058 ; 
      RECT 113.796 104.094 113.868 119.058 ; 
      RECT 113.364 104.094 113.436 119.058 ; 
      RECT 112.932 104.094 113.004 119.058 ; 
      RECT 112.5 104.094 112.572 119.058 ; 
      RECT 112.068 104.094 112.14 119.058 ; 
      RECT 111.636 104.094 111.708 119.058 ; 
      RECT 111.204 104.094 111.276 119.058 ; 
      RECT 110.772 104.094 110.844 119.058 ; 
      RECT 110.34 104.094 110.412 119.058 ; 
      RECT 109.908 104.094 109.98 119.058 ; 
      RECT 109.476 104.094 109.548 119.058 ; 
      RECT 109.044 104.094 109.116 119.058 ; 
      RECT 108.612 104.094 108.684 119.058 ; 
      RECT 108.18 104.094 108.252 119.058 ; 
      RECT 107.748 104.094 107.82 119.058 ; 
      RECT 107.316 104.094 107.388 119.058 ; 
      RECT 106.884 104.094 106.956 119.058 ; 
      RECT 106.452 104.094 106.524 119.058 ; 
      RECT 106.02 104.094 106.092 119.058 ; 
      RECT 105.588 104.094 105.66 119.058 ; 
      RECT 105.156 104.094 105.228 119.058 ; 
      RECT 104.724 104.094 104.796 119.058 ; 
      RECT 104.292 104.094 104.364 119.058 ; 
      RECT 103.86 104.094 103.932 119.058 ; 
      RECT 103.428 104.094 103.5 119.058 ; 
      RECT 102.996 104.094 103.068 119.058 ; 
      RECT 102.564 104.094 102.636 119.058 ; 
      RECT 102.132 104.094 102.204 119.058 ; 
      RECT 101.7 104.094 101.772 119.058 ; 
      RECT 101.268 104.094 101.34 119.058 ; 
      RECT 100.836 104.094 100.908 119.058 ; 
      RECT 100.404 104.094 100.476 119.058 ; 
      RECT 99.972 104.094 100.044 119.058 ; 
      RECT 99.54 104.094 99.612 119.058 ; 
      RECT 99.108 104.094 99.18 119.058 ; 
      RECT 98.676 104.094 98.748 119.058 ; 
      RECT 98.244 104.094 98.316 119.058 ; 
      RECT 97.812 104.094 97.884 119.058 ; 
      RECT 97.38 104.094 97.452 119.058 ; 
      RECT 96.948 104.094 97.02 119.058 ; 
      RECT 96.516 104.094 96.588 119.058 ; 
      RECT 96.084 104.094 96.156 119.058 ; 
      RECT 95.652 104.094 95.724 119.058 ; 
      RECT 95.22 104.094 95.292 119.058 ; 
      RECT 94.788 104.094 94.86 119.058 ; 
      RECT 94.356 104.094 94.428 119.058 ; 
      RECT 93.924 104.094 93.996 119.058 ; 
      RECT 93.492 104.094 93.564 119.058 ; 
      RECT 93.06 104.094 93.132 119.058 ; 
      RECT 92.628 104.094 92.7 119.058 ; 
      RECT 92.196 104.094 92.268 119.058 ; 
      RECT 91.764 104.094 91.836 119.058 ; 
      RECT 91.332 104.094 91.404 119.058 ; 
      RECT 90.9 104.094 90.972 119.058 ; 
      RECT 90.468 104.094 90.54 119.058 ; 
      RECT 90.036 104.094 90.108 119.058 ; 
      RECT 89.604 104.094 89.676 119.058 ; 
      RECT 89.172 104.094 89.244 119.058 ; 
      RECT 88.74 104.094 88.812 119.058 ; 
      RECT 88.308 104.094 88.38 119.058 ; 
      RECT 87.876 104.094 87.948 119.058 ; 
      RECT 87.444 104.094 87.516 119.058 ; 
      RECT 87.012 104.094 87.084 119.058 ; 
      RECT 86.58 104.094 86.652 119.058 ; 
      RECT 86.148 104.094 86.22 119.058 ; 
      RECT 85.716 104.094 85.788 119.058 ; 
      RECT 85.284 104.094 85.356 119.058 ; 
      RECT 84.852 104.094 84.924 119.058 ; 
      RECT 84.42 104.094 84.492 119.058 ; 
      RECT 83.988 104.094 84.06 119.058 ; 
      RECT 83.556 104.094 83.628 119.058 ; 
      RECT 83.124 104.094 83.196 119.058 ; 
      RECT 82.692 104.094 82.764 119.058 ; 
      RECT 82.26 104.094 82.332 119.058 ; 
      RECT 81.828 104.094 81.9 119.058 ; 
      RECT 81.396 104.094 81.468 119.058 ; 
      RECT 80.964 104.094 81.036 119.058 ; 
      RECT 80.532 104.094 80.604 119.058 ; 
      RECT 80.1 104.094 80.172 119.058 ; 
      RECT 79.668 104.094 79.74 119.058 ; 
      RECT 79.236 104.748 79.308 106.148 ; 
      RECT 78.804 104.094 78.876 119.058 ; 
      RECT 78.372 104.094 78.444 119.058 ; 
      RECT 77.94 104.094 78.012 119.058 ; 
      RECT 77.508 104.094 77.58 119.058 ; 
      RECT 77.076 104.094 77.148 119.058 ; 
      RECT 76.644 104.094 76.716 119.058 ; 
      RECT 76.212 104.094 76.284 119.058 ; 
      RECT 75.78 104.094 75.852 119.058 ; 
      RECT 75.348 104.094 75.42 119.058 ; 
      RECT 74.916 104.094 74.988 119.058 ; 
      RECT 74.484 104.094 74.556 119.058 ; 
      RECT 74.052 104.094 74.124 119.058 ; 
      RECT 73.62 104.094 73.692 119.058 ; 
      RECT 73.188 104.094 73.26 119.058 ; 
      RECT 72.756 104.094 72.828 119.058 ; 
      RECT 72.324 104.094 72.396 119.058 ; 
      RECT 71.892 104.094 71.964 119.058 ; 
      RECT 71.46 104.094 71.532 119.058 ; 
      RECT 71.028 104.094 71.1 119.058 ; 
      RECT 70.596 104.094 70.668 119.058 ; 
      RECT 70.164 104.094 70.236 119.058 ; 
      RECT 69.732 104.094 69.804 119.058 ; 
      RECT 69.3 104.094 69.372 119.058 ; 
      RECT 68.868 104.094 68.94 119.058 ; 
      RECT 68.436 104.094 68.508 119.058 ; 
      RECT 68.004 104.094 68.076 119.058 ; 
      RECT 67.572 104.094 67.644 119.058 ; 
      RECT 67.14 104.094 67.212 119.058 ; 
      RECT 66.708 104.094 66.78 119.058 ; 
      RECT 66.276 104.094 66.348 119.058 ; 
      RECT 65.844 104.094 65.916 119.058 ; 
      RECT 65.7 119.902 65.772 122.7208 ; 
      RECT 65.7 125.674 65.772 130.318 ; 
      RECT 65.628 107.39 65.7 110.094 ; 
      RECT 65.628 113.078 65.7 114.27 ; 
      RECT 65.628 117.542 65.7 118.59 ; 
      RECT 65.556 120.156 65.628 122.916 ; 
      RECT 65.556 123.12 65.628 127.062 ; 
      RECT 65.556 127.226 65.628 129.694 ; 
      RECT 65.412 104.094 65.484 137.576 ; 
      RECT 65.268 121.246 65.34 121.578 ; 
      RECT 65.196 107.822 65.268 110.346 ; 
      RECT 65.196 111.998 65.268 112.758 ; 
      RECT 65.196 115.526 65.268 115.722 ; 
      RECT 65.196 118.454 65.268 118.602 ; 
      RECT 65.124 120.026 65.196 134.398 ; 
      RECT 64.764 104.88 64.836 105.432 ; 
      RECT 64.764 106.31 64.836 109.518 ; 
      RECT 64.764 111.71 64.836 113.982 ; 
      RECT 64.764 120.026 64.836 134.398 ; 
      RECT 64.62 111.998 64.692 113.478 ; 
      RECT 64.476 109.406 64.548 109.95 ; 
      RECT 64.476 113.366 64.548 114.27 ; 
      RECT 64.476 118.334 64.548 118.59 ; 
      RECT 64.332 109.814 64.404 109.962 ; 
      RECT 64.332 116.318 64.404 116.49 ; 
      RECT 64.332 118.454 64.404 118.602 ; 
      RECT 64.188 111.062 64.26 113.046 ; 
      RECT 64.188 113.222 64.26 113.982 ; 
      RECT 64.188 117.062 64.26 118.302 ; 
      RECT 64.044 110.63 64.116 115.618 ; 
      RECT 60.156 104.854 60.228 105.47 ; 
      RECT 60.012 104.854 60.084 105.054 ; 
      RECT 59.724 104.854 59.796 105.14 ; 
      RECT 57.132 109.406 57.204 111.03 ; 
      RECT 56.988 113.846 57.06 113.994 ; 
      RECT 56.844 109.55 56.916 111.966 ; 
      RECT 56.7 108.902 56.772 109.158 ; 
      RECT 56.556 105.066 56.628 105.27 ; 
      RECT 56.556 117.542 56.628 118.302 ; 
      RECT 56.556 120.026 56.628 134.398 ; 
      RECT 56.124 106.742 56.196 107.502 ; 
      RECT 56.124 109.838 56.196 118.878 ; 
      RECT 56.052 121.246 56.124 121.578 ; 
      RECT 55.908 104.748 55.98 137.576 ; 
      RECT 55.764 120.156 55.836 122.916 ; 
      RECT 55.764 123.12 55.836 127.062 ; 
      RECT 55.764 127.226 55.836 129.694 ; 
      RECT 55.692 106.742 55.764 108.726 ; 
      RECT 55.692 111.854 55.764 114.126 ; 
      RECT 55.692 115.382 55.764 118.302 ; 
      RECT 55.62 119.902 55.692 122.7208 ; 
      RECT 55.62 125.674 55.692 130.318 ; 
      RECT 55.476 104.748 55.548 106.148 ; 
      RECT 55.476 118.924 55.548 137.576 ; 
      RECT 55.044 104.748 55.116 106.148 ; 
      RECT 54.612 104.748 54.684 106.148 ; 
      RECT 54.18 104.748 54.252 106.148 ; 
      RECT 53.748 104.748 53.82 106.148 ; 
      RECT 53.316 104.748 53.388 106.148 ; 
      RECT 52.884 104.748 52.956 106.148 ; 
      RECT 52.452 104.748 52.524 106.148 ; 
      RECT 52.02 104.748 52.092 106.148 ; 
      RECT 51.588 104.748 51.66 106.148 ; 
      RECT 51.156 104.748 51.228 106.148 ; 
      RECT 50.724 104.748 50.796 106.148 ; 
      RECT 50.292 104.748 50.364 106.148 ; 
      RECT 49.86 104.748 49.932 106.148 ; 
      RECT 49.428 104.748 49.5 106.148 ; 
      RECT 48.996 104.748 49.068 106.148 ; 
      RECT 48.564 104.748 48.636 106.148 ; 
      RECT 48.132 104.748 48.204 106.148 ; 
      RECT 47.7 104.748 47.772 106.148 ; 
      RECT 47.268 104.748 47.34 106.148 ; 
      RECT 46.836 104.748 46.908 106.148 ; 
      RECT 46.404 104.748 46.476 106.148 ; 
      RECT 45.972 104.748 46.044 106.148 ; 
      RECT 45.54 104.748 45.612 106.148 ; 
      RECT 45.108 104.748 45.18 106.148 ; 
      RECT 44.676 104.748 44.748 106.148 ; 
      RECT 44.244 104.748 44.316 106.148 ; 
      RECT 43.812 104.748 43.884 106.148 ; 
      RECT 43.38 104.748 43.452 106.148 ; 
      RECT 42.948 104.748 43.02 106.148 ; 
      RECT 42.516 104.748 42.588 106.148 ; 
      RECT 42.084 104.748 42.156 106.148 ; 
      RECT 41.652 104.748 41.724 106.148 ; 
      RECT 41.22 104.748 41.292 106.148 ; 
      RECT 40.788 104.748 40.86 106.148 ; 
      RECT 40.356 104.748 40.428 106.148 ; 
      RECT 39.924 104.748 39.996 106.148 ; 
      RECT 39.492 104.748 39.564 106.148 ; 
      RECT 39.06 104.748 39.132 106.148 ; 
      RECT 38.628 104.748 38.7 106.148 ; 
      RECT 38.196 104.748 38.268 106.148 ; 
      RECT 37.764 104.748 37.836 106.148 ; 
      RECT 37.332 104.748 37.404 106.148 ; 
      RECT 36.9 104.748 36.972 106.148 ; 
      RECT 36.468 104.748 36.54 106.148 ; 
      RECT 36.036 104.748 36.108 106.148 ; 
      RECT 35.604 104.748 35.676 106.148 ; 
      RECT 35.172 104.748 35.244 106.148 ; 
      RECT 34.74 104.748 34.812 106.148 ; 
      RECT 34.308 104.748 34.38 106.148 ; 
      RECT 33.876 104.748 33.948 106.148 ; 
      RECT 33.444 104.748 33.516 106.148 ; 
      RECT 33.012 104.748 33.084 106.148 ; 
      RECT 32.58 104.748 32.652 106.148 ; 
      RECT 32.148 104.748 32.22 106.148 ; 
      RECT 31.716 104.748 31.788 106.148 ; 
      RECT 31.284 104.748 31.356 106.148 ; 
      RECT 30.852 104.748 30.924 106.148 ; 
      RECT 30.42 104.748 30.492 106.148 ; 
      RECT 29.988 104.748 30.06 106.148 ; 
      RECT 29.556 104.748 29.628 106.148 ; 
      RECT 29.124 104.748 29.196 106.148 ; 
      RECT 28.692 104.748 28.764 106.148 ; 
      RECT 28.26 104.748 28.332 106.148 ; 
      RECT 27.828 104.748 27.9 106.148 ; 
      RECT 27.396 104.748 27.468 106.148 ; 
      RECT 26.964 104.748 27.036 106.148 ; 
      RECT 26.532 104.748 26.604 106.148 ; 
      RECT 26.1 104.748 26.172 106.148 ; 
      RECT 25.668 104.748 25.74 106.148 ; 
      RECT 25.236 104.748 25.308 106.148 ; 
      RECT 24.804 104.748 24.876 106.148 ; 
      RECT 24.372 104.748 24.444 106.148 ; 
      RECT 23.94 104.748 24.012 106.148 ; 
      RECT 23.508 104.748 23.58 106.148 ; 
      RECT 23.076 104.748 23.148 106.148 ; 
      RECT 22.644 104.748 22.716 106.148 ; 
      RECT 22.212 104.748 22.284 106.148 ; 
      RECT 21.78 104.748 21.852 106.148 ; 
      RECT 21.348 104.748 21.42 106.148 ; 
      RECT 20.916 104.748 20.988 106.148 ; 
      RECT 20.484 104.748 20.556 106.148 ; 
      RECT 20.052 104.748 20.124 106.148 ; 
      RECT 19.62 104.748 19.692 106.148 ; 
      RECT 19.188 104.748 19.26 106.148 ; 
      RECT 18.756 104.748 18.828 106.148 ; 
      RECT 18.324 104.748 18.396 106.148 ; 
      RECT 17.892 104.748 17.964 106.148 ; 
      RECT 17.46 104.748 17.532 106.148 ; 
      RECT 17.028 104.748 17.1 106.148 ; 
      RECT 16.596 104.748 16.668 106.148 ; 
      RECT 16.164 104.748 16.236 106.148 ; 
      RECT 15.732 104.748 15.804 106.148 ; 
      RECT 15.3 104.748 15.372 106.148 ; 
      RECT 14.868 104.748 14.94 106.148 ; 
      RECT 14.436 104.748 14.508 106.148 ; 
      RECT 14.004 104.748 14.076 106.148 ; 
      RECT 13.572 104.748 13.644 106.148 ; 
      RECT 13.14 104.748 13.212 106.148 ; 
      RECT 12.708 104.748 12.78 106.148 ; 
      RECT 12.276 104.748 12.348 106.148 ; 
      RECT 11.844 104.748 11.916 106.148 ; 
      RECT 11.412 104.748 11.484 106.148 ; 
      RECT 10.98 104.748 11.052 106.148 ; 
      RECT 10.548 104.748 10.62 106.148 ; 
      RECT 10.116 104.748 10.188 106.148 ; 
      RECT 9.684 104.748 9.756 106.148 ; 
      RECT 9.252 104.748 9.324 106.148 ; 
      RECT 8.82 104.748 8.892 106.148 ; 
      RECT 8.388 104.748 8.46 106.148 ; 
      RECT 7.956 104.748 8.028 106.148 ; 
      RECT 7.524 104.748 7.596 106.148 ; 
      RECT 7.092 104.748 7.164 106.148 ; 
      RECT 6.66 104.748 6.732 106.148 ; 
      RECT 6.228 104.748 6.3 106.148 ; 
      RECT 5.796 104.748 5.868 106.148 ; 
      RECT 5.364 104.748 5.436 106.148 ; 
      RECT 4.932 104.748 5.004 106.148 ; 
      RECT 4.5 104.748 4.572 106.148 ; 
      RECT 4.068 104.748 4.14 106.148 ; 
      RECT 3.636 104.748 3.708 106.148 ; 
      RECT 3.204 104.748 3.276 106.148 ; 
      RECT 2.772 104.748 2.844 106.148 ; 
      RECT 2.34 104.748 2.412 106.148 ; 
      RECT 1.908 104.748 1.98 106.148 ; 
      RECT 1.476 104.748 1.548 106.148 ; 
      RECT 1.044 104.748 1.116 106.148 ; 
      RECT 0.612 104.748 0.684 137.576 ; 
      RECT 0.468 104.748 0.54 137.576 ; 
        RECT 62.444 137.568 62.516 141.31 ; 
        RECT 62.3 137.568 62.372 141.31 ; 
        RECT 62.156 139.876 62.228 141.166 ; 
        RECT 61.688 140.664 61.76 141.102 ; 
        RECT 61.652 137.698 61.724 138.656 ; 
        RECT 61.508 140.022 61.58 140.636 ; 
        RECT 61.184 140.124 61.256 141.156 ; 
        RECT 59.024 137.568 59.096 141.31 ; 
        RECT 58.88 137.568 58.952 141.31 ; 
        RECT 58.736 138.292 58.808 140.564 ; 
        RECT 62.444 141.888 62.516 145.63 ; 
        RECT 62.3 141.888 62.372 145.63 ; 
        RECT 62.156 144.196 62.228 145.486 ; 
        RECT 61.688 144.984 61.76 145.422 ; 
        RECT 61.652 142.018 61.724 142.976 ; 
        RECT 61.508 144.342 61.58 144.956 ; 
        RECT 61.184 144.444 61.256 145.476 ; 
        RECT 59.024 141.888 59.096 145.63 ; 
        RECT 58.88 141.888 58.952 145.63 ; 
        RECT 58.736 142.612 58.808 144.884 ; 
        RECT 62.444 146.208 62.516 149.95 ; 
        RECT 62.3 146.208 62.372 149.95 ; 
        RECT 62.156 148.516 62.228 149.806 ; 
        RECT 61.688 149.304 61.76 149.742 ; 
        RECT 61.652 146.338 61.724 147.296 ; 
        RECT 61.508 148.662 61.58 149.276 ; 
        RECT 61.184 148.764 61.256 149.796 ; 
        RECT 59.024 146.208 59.096 149.95 ; 
        RECT 58.88 146.208 58.952 149.95 ; 
        RECT 58.736 146.932 58.808 149.204 ; 
        RECT 62.444 150.528 62.516 154.27 ; 
        RECT 62.3 150.528 62.372 154.27 ; 
        RECT 62.156 152.836 62.228 154.126 ; 
        RECT 61.688 153.624 61.76 154.062 ; 
        RECT 61.652 150.658 61.724 151.616 ; 
        RECT 61.508 152.982 61.58 153.596 ; 
        RECT 61.184 153.084 61.256 154.116 ; 
        RECT 59.024 150.528 59.096 154.27 ; 
        RECT 58.88 150.528 58.952 154.27 ; 
        RECT 58.736 151.252 58.808 153.524 ; 
        RECT 62.444 154.848 62.516 158.59 ; 
        RECT 62.3 154.848 62.372 158.59 ; 
        RECT 62.156 157.156 62.228 158.446 ; 
        RECT 61.688 157.944 61.76 158.382 ; 
        RECT 61.652 154.978 61.724 155.936 ; 
        RECT 61.508 157.302 61.58 157.916 ; 
        RECT 61.184 157.404 61.256 158.436 ; 
        RECT 59.024 154.848 59.096 158.59 ; 
        RECT 58.88 154.848 58.952 158.59 ; 
        RECT 58.736 155.572 58.808 157.844 ; 
        RECT 62.444 159.168 62.516 162.91 ; 
        RECT 62.3 159.168 62.372 162.91 ; 
        RECT 62.156 161.476 62.228 162.766 ; 
        RECT 61.688 162.264 61.76 162.702 ; 
        RECT 61.652 159.298 61.724 160.256 ; 
        RECT 61.508 161.622 61.58 162.236 ; 
        RECT 61.184 161.724 61.256 162.756 ; 
        RECT 59.024 159.168 59.096 162.91 ; 
        RECT 58.88 159.168 58.952 162.91 ; 
        RECT 58.736 159.892 58.808 162.164 ; 
        RECT 62.444 163.488 62.516 167.23 ; 
        RECT 62.3 163.488 62.372 167.23 ; 
        RECT 62.156 165.796 62.228 167.086 ; 
        RECT 61.688 166.584 61.76 167.022 ; 
        RECT 61.652 163.618 61.724 164.576 ; 
        RECT 61.508 165.942 61.58 166.556 ; 
        RECT 61.184 166.044 61.256 167.076 ; 
        RECT 59.024 163.488 59.096 167.23 ; 
        RECT 58.88 163.488 58.952 167.23 ; 
        RECT 58.736 164.212 58.808 166.484 ; 
        RECT 62.444 167.808 62.516 171.55 ; 
        RECT 62.3 167.808 62.372 171.55 ; 
        RECT 62.156 170.116 62.228 171.406 ; 
        RECT 61.688 170.904 61.76 171.342 ; 
        RECT 61.652 167.938 61.724 168.896 ; 
        RECT 61.508 170.262 61.58 170.876 ; 
        RECT 61.184 170.364 61.256 171.396 ; 
        RECT 59.024 167.808 59.096 171.55 ; 
        RECT 58.88 167.808 58.952 171.55 ; 
        RECT 58.736 168.532 58.808 170.804 ; 
        RECT 62.444 172.128 62.516 175.87 ; 
        RECT 62.3 172.128 62.372 175.87 ; 
        RECT 62.156 174.436 62.228 175.726 ; 
        RECT 61.688 175.224 61.76 175.662 ; 
        RECT 61.652 172.258 61.724 173.216 ; 
        RECT 61.508 174.582 61.58 175.196 ; 
        RECT 61.184 174.684 61.256 175.716 ; 
        RECT 59.024 172.128 59.096 175.87 ; 
        RECT 58.88 172.128 58.952 175.87 ; 
        RECT 58.736 172.852 58.808 175.124 ; 
        RECT 62.444 176.448 62.516 180.19 ; 
        RECT 62.3 176.448 62.372 180.19 ; 
        RECT 62.156 178.756 62.228 180.046 ; 
        RECT 61.688 179.544 61.76 179.982 ; 
        RECT 61.652 176.578 61.724 177.536 ; 
        RECT 61.508 178.902 61.58 179.516 ; 
        RECT 61.184 179.004 61.256 180.036 ; 
        RECT 59.024 176.448 59.096 180.19 ; 
        RECT 58.88 176.448 58.952 180.19 ; 
        RECT 58.736 177.172 58.808 179.444 ; 
        RECT 62.444 180.768 62.516 184.51 ; 
        RECT 62.3 180.768 62.372 184.51 ; 
        RECT 62.156 183.076 62.228 184.366 ; 
        RECT 61.688 183.864 61.76 184.302 ; 
        RECT 61.652 180.898 61.724 181.856 ; 
        RECT 61.508 183.222 61.58 183.836 ; 
        RECT 61.184 183.324 61.256 184.356 ; 
        RECT 59.024 180.768 59.096 184.51 ; 
        RECT 58.88 180.768 58.952 184.51 ; 
        RECT 58.736 181.492 58.808 183.764 ; 
        RECT 62.444 185.088 62.516 188.83 ; 
        RECT 62.3 185.088 62.372 188.83 ; 
        RECT 62.156 187.396 62.228 188.686 ; 
        RECT 61.688 188.184 61.76 188.622 ; 
        RECT 61.652 185.218 61.724 186.176 ; 
        RECT 61.508 187.542 61.58 188.156 ; 
        RECT 61.184 187.644 61.256 188.676 ; 
        RECT 59.024 185.088 59.096 188.83 ; 
        RECT 58.88 185.088 58.952 188.83 ; 
        RECT 58.736 185.812 58.808 188.084 ; 
        RECT 62.444 189.408 62.516 193.15 ; 
        RECT 62.3 189.408 62.372 193.15 ; 
        RECT 62.156 191.716 62.228 193.006 ; 
        RECT 61.688 192.504 61.76 192.942 ; 
        RECT 61.652 189.538 61.724 190.496 ; 
        RECT 61.508 191.862 61.58 192.476 ; 
        RECT 61.184 191.964 61.256 192.996 ; 
        RECT 59.024 189.408 59.096 193.15 ; 
        RECT 58.88 189.408 58.952 193.15 ; 
        RECT 58.736 190.132 58.808 192.404 ; 
        RECT 62.444 193.728 62.516 197.47 ; 
        RECT 62.3 193.728 62.372 197.47 ; 
        RECT 62.156 196.036 62.228 197.326 ; 
        RECT 61.688 196.824 61.76 197.262 ; 
        RECT 61.652 193.858 61.724 194.816 ; 
        RECT 61.508 196.182 61.58 196.796 ; 
        RECT 61.184 196.284 61.256 197.316 ; 
        RECT 59.024 193.728 59.096 197.47 ; 
        RECT 58.88 193.728 58.952 197.47 ; 
        RECT 58.736 194.452 58.808 196.724 ; 
        RECT 62.444 198.048 62.516 201.79 ; 
        RECT 62.3 198.048 62.372 201.79 ; 
        RECT 62.156 200.356 62.228 201.646 ; 
        RECT 61.688 201.144 61.76 201.582 ; 
        RECT 61.652 198.178 61.724 199.136 ; 
        RECT 61.508 200.502 61.58 201.116 ; 
        RECT 61.184 200.604 61.256 201.636 ; 
        RECT 59.024 198.048 59.096 201.79 ; 
        RECT 58.88 198.048 58.952 201.79 ; 
        RECT 58.736 198.772 58.808 201.044 ; 
        RECT 62.444 202.368 62.516 206.11 ; 
        RECT 62.3 202.368 62.372 206.11 ; 
        RECT 62.156 204.676 62.228 205.966 ; 
        RECT 61.688 205.464 61.76 205.902 ; 
        RECT 61.652 202.498 61.724 203.456 ; 
        RECT 61.508 204.822 61.58 205.436 ; 
        RECT 61.184 204.924 61.256 205.956 ; 
        RECT 59.024 202.368 59.096 206.11 ; 
        RECT 58.88 202.368 58.952 206.11 ; 
        RECT 58.736 203.092 58.808 205.364 ; 
        RECT 62.444 206.688 62.516 210.43 ; 
        RECT 62.3 206.688 62.372 210.43 ; 
        RECT 62.156 208.996 62.228 210.286 ; 
        RECT 61.688 209.784 61.76 210.222 ; 
        RECT 61.652 206.818 61.724 207.776 ; 
        RECT 61.508 209.142 61.58 209.756 ; 
        RECT 61.184 209.244 61.256 210.276 ; 
        RECT 59.024 206.688 59.096 210.43 ; 
        RECT 58.88 206.688 58.952 210.43 ; 
        RECT 58.736 207.412 58.808 209.684 ; 
        RECT 62.444 211.008 62.516 214.75 ; 
        RECT 62.3 211.008 62.372 214.75 ; 
        RECT 62.156 213.316 62.228 214.606 ; 
        RECT 61.688 214.104 61.76 214.542 ; 
        RECT 61.652 211.138 61.724 212.096 ; 
        RECT 61.508 213.462 61.58 214.076 ; 
        RECT 61.184 213.564 61.256 214.596 ; 
        RECT 59.024 211.008 59.096 214.75 ; 
        RECT 58.88 211.008 58.952 214.75 ; 
        RECT 58.736 211.732 58.808 214.004 ; 
        RECT 62.444 215.328 62.516 219.07 ; 
        RECT 62.3 215.328 62.372 219.07 ; 
        RECT 62.156 217.636 62.228 218.926 ; 
        RECT 61.688 218.424 61.76 218.862 ; 
        RECT 61.652 215.458 61.724 216.416 ; 
        RECT 61.508 217.782 61.58 218.396 ; 
        RECT 61.184 217.884 61.256 218.916 ; 
        RECT 59.024 215.328 59.096 219.07 ; 
        RECT 58.88 215.328 58.952 219.07 ; 
        RECT 58.736 216.052 58.808 218.324 ; 
        RECT 62.444 219.648 62.516 223.39 ; 
        RECT 62.3 219.648 62.372 223.39 ; 
        RECT 62.156 221.956 62.228 223.246 ; 
        RECT 61.688 222.744 61.76 223.182 ; 
        RECT 61.652 219.778 61.724 220.736 ; 
        RECT 61.508 222.102 61.58 222.716 ; 
        RECT 61.184 222.204 61.256 223.236 ; 
        RECT 59.024 219.648 59.096 223.39 ; 
        RECT 58.88 219.648 58.952 223.39 ; 
        RECT 58.736 220.372 58.808 222.644 ; 
        RECT 62.444 223.968 62.516 227.71 ; 
        RECT 62.3 223.968 62.372 227.71 ; 
        RECT 62.156 226.276 62.228 227.566 ; 
        RECT 61.688 227.064 61.76 227.502 ; 
        RECT 61.652 224.098 61.724 225.056 ; 
        RECT 61.508 226.422 61.58 227.036 ; 
        RECT 61.184 226.524 61.256 227.556 ; 
        RECT 59.024 223.968 59.096 227.71 ; 
        RECT 58.88 223.968 58.952 227.71 ; 
        RECT 58.736 224.692 58.808 226.964 ; 
        RECT 62.444 228.288 62.516 232.03 ; 
        RECT 62.3 228.288 62.372 232.03 ; 
        RECT 62.156 230.596 62.228 231.886 ; 
        RECT 61.688 231.384 61.76 231.822 ; 
        RECT 61.652 228.418 61.724 229.376 ; 
        RECT 61.508 230.742 61.58 231.356 ; 
        RECT 61.184 230.844 61.256 231.876 ; 
        RECT 59.024 228.288 59.096 232.03 ; 
        RECT 58.88 228.288 58.952 232.03 ; 
        RECT 58.736 229.012 58.808 231.284 ; 
        RECT 62.444 232.608 62.516 236.35 ; 
        RECT 62.3 232.608 62.372 236.35 ; 
        RECT 62.156 234.916 62.228 236.206 ; 
        RECT 61.688 235.704 61.76 236.142 ; 
        RECT 61.652 232.738 61.724 233.696 ; 
        RECT 61.508 235.062 61.58 235.676 ; 
        RECT 61.184 235.164 61.256 236.196 ; 
        RECT 59.024 232.608 59.096 236.35 ; 
        RECT 58.88 232.608 58.952 236.35 ; 
        RECT 58.736 233.332 58.808 235.604 ; 
        RECT 62.444 236.928 62.516 240.67 ; 
        RECT 62.3 236.928 62.372 240.67 ; 
        RECT 62.156 239.236 62.228 240.526 ; 
        RECT 61.688 240.024 61.76 240.462 ; 
        RECT 61.652 237.058 61.724 238.016 ; 
        RECT 61.508 239.382 61.58 239.996 ; 
        RECT 61.184 239.484 61.256 240.516 ; 
        RECT 59.024 236.928 59.096 240.67 ; 
        RECT 58.88 236.928 58.952 240.67 ; 
        RECT 58.736 237.652 58.808 239.924 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 62.212 1.026 62.724 5.4 ; 
      RECT 62.156 3.688 62.724 4.978 ; 
      RECT 61.276 2.596 61.812 5.4 ; 
      RECT 61.184 3.936 61.812 4.968 ; 
      RECT 61.276 1.026 61.668 5.4 ; 
      RECT 61.276 1.51 61.724 2.468 ; 
      RECT 61.276 1.026 61.812 1.382 ; 
      RECT 60.376 2.828 60.912 5.4 ; 
      RECT 60.376 1.026 60.768 5.4 ; 
      RECT 58.708 1.026 59.04 5.4 ; 
      RECT 58.708 1.38 59.096 5.122 ; 
      RECT 121.072 1.026 121.412 5.4 ; 
      RECT 120.496 1.026 120.6 5.4 ; 
      RECT 120.064 1.026 120.168 5.4 ; 
      RECT 119.632 1.026 119.736 5.4 ; 
      RECT 119.2 1.026 119.304 5.4 ; 
      RECT 118.768 1.026 118.872 5.4 ; 
      RECT 118.336 1.026 118.44 5.4 ; 
      RECT 117.904 1.026 118.008 5.4 ; 
      RECT 117.472 1.026 117.576 5.4 ; 
      RECT 117.04 1.026 117.144 5.4 ; 
      RECT 116.608 1.026 116.712 5.4 ; 
      RECT 116.176 1.026 116.28 5.4 ; 
      RECT 115.744 1.026 115.848 5.4 ; 
      RECT 115.312 1.026 115.416 5.4 ; 
      RECT 114.88 1.026 114.984 5.4 ; 
      RECT 114.448 1.026 114.552 5.4 ; 
      RECT 114.016 1.026 114.12 5.4 ; 
      RECT 113.584 1.026 113.688 5.4 ; 
      RECT 113.152 1.026 113.256 5.4 ; 
      RECT 112.72 1.026 112.824 5.4 ; 
      RECT 112.288 1.026 112.392 5.4 ; 
      RECT 111.856 1.026 111.96 5.4 ; 
      RECT 111.424 1.026 111.528 5.4 ; 
      RECT 110.992 1.026 111.096 5.4 ; 
      RECT 110.56 1.026 110.664 5.4 ; 
      RECT 110.128 1.026 110.232 5.4 ; 
      RECT 109.696 1.026 109.8 5.4 ; 
      RECT 109.264 1.026 109.368 5.4 ; 
      RECT 108.832 1.026 108.936 5.4 ; 
      RECT 108.4 1.026 108.504 5.4 ; 
      RECT 107.968 1.026 108.072 5.4 ; 
      RECT 107.536 1.026 107.64 5.4 ; 
      RECT 107.104 1.026 107.208 5.4 ; 
      RECT 106.672 1.026 106.776 5.4 ; 
      RECT 106.24 1.026 106.344 5.4 ; 
      RECT 105.808 1.026 105.912 5.4 ; 
      RECT 105.376 1.026 105.48 5.4 ; 
      RECT 104.944 1.026 105.048 5.4 ; 
      RECT 104.512 1.026 104.616 5.4 ; 
      RECT 104.08 1.026 104.184 5.4 ; 
      RECT 103.648 1.026 103.752 5.4 ; 
      RECT 103.216 1.026 103.32 5.4 ; 
      RECT 102.784 1.026 102.888 5.4 ; 
      RECT 102.352 1.026 102.456 5.4 ; 
      RECT 101.92 1.026 102.024 5.4 ; 
      RECT 101.488 1.026 101.592 5.4 ; 
      RECT 101.056 1.026 101.16 5.4 ; 
      RECT 100.624 1.026 100.728 5.4 ; 
      RECT 100.192 1.026 100.296 5.4 ; 
      RECT 99.76 1.026 99.864 5.4 ; 
      RECT 99.328 1.026 99.432 5.4 ; 
      RECT 98.896 1.026 99 5.4 ; 
      RECT 98.464 1.026 98.568 5.4 ; 
      RECT 98.032 1.026 98.136 5.4 ; 
      RECT 97.6 1.026 97.704 5.4 ; 
      RECT 97.168 1.026 97.272 5.4 ; 
      RECT 96.736 1.026 96.84 5.4 ; 
      RECT 96.304 1.026 96.408 5.4 ; 
      RECT 95.872 1.026 95.976 5.4 ; 
      RECT 95.44 1.026 95.544 5.4 ; 
      RECT 95.008 1.026 95.112 5.4 ; 
      RECT 94.576 1.026 94.68 5.4 ; 
      RECT 94.144 1.026 94.248 5.4 ; 
      RECT 93.712 1.026 93.816 5.4 ; 
      RECT 93.28 1.026 93.384 5.4 ; 
      RECT 92.848 1.026 92.952 5.4 ; 
      RECT 92.416 1.026 92.52 5.4 ; 
      RECT 91.984 1.026 92.088 5.4 ; 
      RECT 91.552 1.026 91.656 5.4 ; 
      RECT 91.12 1.026 91.224 5.4 ; 
      RECT 90.688 1.026 90.792 5.4 ; 
      RECT 90.256 1.026 90.36 5.4 ; 
      RECT 89.824 1.026 89.928 5.4 ; 
      RECT 89.392 1.026 89.496 5.4 ; 
      RECT 88.96 1.026 89.064 5.4 ; 
      RECT 88.528 1.026 88.632 5.4 ; 
      RECT 88.096 1.026 88.2 5.4 ; 
      RECT 87.664 1.026 87.768 5.4 ; 
      RECT 87.232 1.026 87.336 5.4 ; 
      RECT 86.8 1.026 86.904 5.4 ; 
      RECT 86.368 1.026 86.472 5.4 ; 
      RECT 85.936 1.026 86.04 5.4 ; 
      RECT 85.504 1.026 85.608 5.4 ; 
      RECT 85.072 1.026 85.176 5.4 ; 
      RECT 84.64 1.026 84.744 5.4 ; 
      RECT 84.208 1.026 84.312 5.4 ; 
      RECT 83.776 1.026 83.88 5.4 ; 
      RECT 83.344 1.026 83.448 5.4 ; 
      RECT 82.912 1.026 83.016 5.4 ; 
      RECT 82.48 1.026 82.584 5.4 ; 
      RECT 82.048 1.026 82.152 5.4 ; 
      RECT 81.616 1.026 81.72 5.4 ; 
      RECT 81.184 1.026 81.288 5.4 ; 
      RECT 80.752 1.026 80.856 5.4 ; 
      RECT 80.32 1.026 80.424 5.4 ; 
      RECT 79.888 1.026 79.992 5.4 ; 
      RECT 79.456 1.026 79.56 5.4 ; 
      RECT 79.024 1.026 79.128 5.4 ; 
      RECT 78.592 1.026 78.696 5.4 ; 
      RECT 78.16 1.026 78.264 5.4 ; 
      RECT 77.728 1.026 77.832 5.4 ; 
      RECT 77.296 1.026 77.4 5.4 ; 
      RECT 76.864 1.026 76.968 5.4 ; 
      RECT 76.432 1.026 76.536 5.4 ; 
      RECT 76 1.026 76.104 5.4 ; 
      RECT 75.568 1.026 75.672 5.4 ; 
      RECT 75.136 1.026 75.24 5.4 ; 
      RECT 74.704 1.026 74.808 5.4 ; 
      RECT 74.272 1.026 74.376 5.4 ; 
      RECT 73.84 1.026 73.944 5.4 ; 
      RECT 73.408 1.026 73.512 5.4 ; 
      RECT 72.976 1.026 73.08 5.4 ; 
      RECT 72.544 1.026 72.648 5.4 ; 
      RECT 72.112 1.026 72.216 5.4 ; 
      RECT 71.68 1.026 71.784 5.4 ; 
      RECT 71.248 1.026 71.352 5.4 ; 
      RECT 70.816 1.026 70.92 5.4 ; 
      RECT 70.384 1.026 70.488 5.4 ; 
      RECT 69.952 1.026 70.056 5.4 ; 
      RECT 69.52 1.026 69.624 5.4 ; 
      RECT 69.088 1.026 69.192 5.4 ; 
      RECT 68.656 1.026 68.76 5.4 ; 
      RECT 68.224 1.026 68.328 5.4 ; 
      RECT 67.792 1.026 67.896 5.4 ; 
      RECT 67.36 1.026 67.464 5.4 ; 
      RECT 66.928 1.026 67.032 5.4 ; 
      RECT 66.496 1.026 66.6 5.4 ; 
      RECT 66.064 1.026 66.168 5.4 ; 
      RECT 65.632 1.026 65.736 5.4 ; 
      RECT 65.2 1.026 65.304 5.4 ; 
      RECT 64.348 1.026 64.656 5.4 ; 
      RECT 56.776 1.026 57.084 5.4 ; 
      RECT 56.128 1.026 56.232 5.4 ; 
      RECT 55.696 1.026 55.8 5.4 ; 
      RECT 55.264 1.026 55.368 5.4 ; 
      RECT 54.832 1.026 54.936 5.4 ; 
      RECT 54.4 1.026 54.504 5.4 ; 
      RECT 53.968 1.026 54.072 5.4 ; 
      RECT 53.536 1.026 53.64 5.4 ; 
      RECT 53.104 1.026 53.208 5.4 ; 
      RECT 52.672 1.026 52.776 5.4 ; 
      RECT 52.24 1.026 52.344 5.4 ; 
      RECT 51.808 1.026 51.912 5.4 ; 
      RECT 51.376 1.026 51.48 5.4 ; 
      RECT 50.944 1.026 51.048 5.4 ; 
      RECT 50.512 1.026 50.616 5.4 ; 
      RECT 50.08 1.026 50.184 5.4 ; 
      RECT 49.648 1.026 49.752 5.4 ; 
      RECT 49.216 1.026 49.32 5.4 ; 
      RECT 48.784 1.026 48.888 5.4 ; 
      RECT 48.352 1.026 48.456 5.4 ; 
      RECT 47.92 1.026 48.024 5.4 ; 
      RECT 47.488 1.026 47.592 5.4 ; 
      RECT 47.056 1.026 47.16 5.4 ; 
      RECT 46.624 1.026 46.728 5.4 ; 
      RECT 46.192 1.026 46.296 5.4 ; 
      RECT 45.76 1.026 45.864 5.4 ; 
      RECT 45.328 1.026 45.432 5.4 ; 
      RECT 44.896 1.026 45 5.4 ; 
      RECT 44.464 1.026 44.568 5.4 ; 
      RECT 44.032 1.026 44.136 5.4 ; 
      RECT 43.6 1.026 43.704 5.4 ; 
      RECT 43.168 1.026 43.272 5.4 ; 
      RECT 42.736 1.026 42.84 5.4 ; 
      RECT 42.304 1.026 42.408 5.4 ; 
      RECT 41.872 1.026 41.976 5.4 ; 
      RECT 41.44 1.026 41.544 5.4 ; 
      RECT 41.008 1.026 41.112 5.4 ; 
      RECT 40.576 1.026 40.68 5.4 ; 
      RECT 40.144 1.026 40.248 5.4 ; 
      RECT 39.712 1.026 39.816 5.4 ; 
      RECT 39.28 1.026 39.384 5.4 ; 
      RECT 38.848 1.026 38.952 5.4 ; 
      RECT 38.416 1.026 38.52 5.4 ; 
      RECT 37.984 1.026 38.088 5.4 ; 
      RECT 37.552 1.026 37.656 5.4 ; 
      RECT 37.12 1.026 37.224 5.4 ; 
      RECT 36.688 1.026 36.792 5.4 ; 
      RECT 36.256 1.026 36.36 5.4 ; 
      RECT 35.824 1.026 35.928 5.4 ; 
      RECT 35.392 1.026 35.496 5.4 ; 
      RECT 34.96 1.026 35.064 5.4 ; 
      RECT 34.528 1.026 34.632 5.4 ; 
      RECT 34.096 1.026 34.2 5.4 ; 
      RECT 33.664 1.026 33.768 5.4 ; 
      RECT 33.232 1.026 33.336 5.4 ; 
      RECT 32.8 1.026 32.904 5.4 ; 
      RECT 32.368 1.026 32.472 5.4 ; 
      RECT 31.936 1.026 32.04 5.4 ; 
      RECT 31.504 1.026 31.608 5.4 ; 
      RECT 31.072 1.026 31.176 5.4 ; 
      RECT 30.64 1.026 30.744 5.4 ; 
      RECT 30.208 1.026 30.312 5.4 ; 
      RECT 29.776 1.026 29.88 5.4 ; 
      RECT 29.344 1.026 29.448 5.4 ; 
      RECT 28.912 1.026 29.016 5.4 ; 
      RECT 28.48 1.026 28.584 5.4 ; 
      RECT 28.048 1.026 28.152 5.4 ; 
      RECT 27.616 1.026 27.72 5.4 ; 
      RECT 27.184 1.026 27.288 5.4 ; 
      RECT 26.752 1.026 26.856 5.4 ; 
      RECT 26.32 1.026 26.424 5.4 ; 
      RECT 25.888 1.026 25.992 5.4 ; 
      RECT 25.456 1.026 25.56 5.4 ; 
      RECT 25.024 1.026 25.128 5.4 ; 
      RECT 24.592 1.026 24.696 5.4 ; 
      RECT 24.16 1.026 24.264 5.4 ; 
      RECT 23.728 1.026 23.832 5.4 ; 
      RECT 23.296 1.026 23.4 5.4 ; 
      RECT 22.864 1.026 22.968 5.4 ; 
      RECT 22.432 1.026 22.536 5.4 ; 
      RECT 22 1.026 22.104 5.4 ; 
      RECT 21.568 1.026 21.672 5.4 ; 
      RECT 21.136 1.026 21.24 5.4 ; 
      RECT 20.704 1.026 20.808 5.4 ; 
      RECT 20.272 1.026 20.376 5.4 ; 
      RECT 19.84 1.026 19.944 5.4 ; 
      RECT 19.408 1.026 19.512 5.4 ; 
      RECT 18.976 1.026 19.08 5.4 ; 
      RECT 18.544 1.026 18.648 5.4 ; 
      RECT 18.112 1.026 18.216 5.4 ; 
      RECT 17.68 1.026 17.784 5.4 ; 
      RECT 17.248 1.026 17.352 5.4 ; 
      RECT 16.816 1.026 16.92 5.4 ; 
      RECT 16.384 1.026 16.488 5.4 ; 
      RECT 15.952 1.026 16.056 5.4 ; 
      RECT 15.52 1.026 15.624 5.4 ; 
      RECT 15.088 1.026 15.192 5.4 ; 
      RECT 14.656 1.026 14.76 5.4 ; 
      RECT 14.224 1.026 14.328 5.4 ; 
      RECT 13.792 1.026 13.896 5.4 ; 
      RECT 13.36 1.026 13.464 5.4 ; 
      RECT 12.928 1.026 13.032 5.4 ; 
      RECT 12.496 1.026 12.6 5.4 ; 
      RECT 12.064 1.026 12.168 5.4 ; 
      RECT 11.632 1.026 11.736 5.4 ; 
      RECT 11.2 1.026 11.304 5.4 ; 
      RECT 10.768 1.026 10.872 5.4 ; 
      RECT 10.336 1.026 10.44 5.4 ; 
      RECT 9.904 1.026 10.008 5.4 ; 
      RECT 9.472 1.026 9.576 5.4 ; 
      RECT 9.04 1.026 9.144 5.4 ; 
      RECT 8.608 1.026 8.712 5.4 ; 
      RECT 8.176 1.026 8.28 5.4 ; 
      RECT 7.744 1.026 7.848 5.4 ; 
      RECT 7.312 1.026 7.416 5.4 ; 
      RECT 6.88 1.026 6.984 5.4 ; 
      RECT 6.448 1.026 6.552 5.4 ; 
      RECT 6.016 1.026 6.12 5.4 ; 
      RECT 5.584 1.026 5.688 5.4 ; 
      RECT 5.152 1.026 5.256 5.4 ; 
      RECT 4.72 1.026 4.824 5.4 ; 
      RECT 4.288 1.026 4.392 5.4 ; 
      RECT 3.856 1.026 3.96 5.4 ; 
      RECT 3.424 1.026 3.528 5.4 ; 
      RECT 2.992 1.026 3.096 5.4 ; 
      RECT 2.56 1.026 2.664 5.4 ; 
      RECT 2.128 1.026 2.232 5.4 ; 
      RECT 1.696 1.026 1.8 5.4 ; 
      RECT 1.264 1.026 1.368 5.4 ; 
      RECT 0.832 1.026 0.936 5.4 ; 
      RECT 0.02 1.026 0.36 5.4 ; 
      RECT 62.212 5.346 62.724 9.72 ; 
      RECT 62.156 8.008 62.724 9.298 ; 
      RECT 61.276 6.916 61.812 9.72 ; 
      RECT 61.184 8.256 61.812 9.288 ; 
      RECT 61.276 5.346 61.668 9.72 ; 
      RECT 61.276 5.83 61.724 6.788 ; 
      RECT 61.276 5.346 61.812 5.702 ; 
      RECT 60.376 7.148 60.912 9.72 ; 
      RECT 60.376 5.346 60.768 9.72 ; 
      RECT 58.708 5.346 59.04 9.72 ; 
      RECT 58.708 5.7 59.096 9.442 ; 
      RECT 121.072 5.346 121.412 9.72 ; 
      RECT 120.496 5.346 120.6 9.72 ; 
      RECT 120.064 5.346 120.168 9.72 ; 
      RECT 119.632 5.346 119.736 9.72 ; 
      RECT 119.2 5.346 119.304 9.72 ; 
      RECT 118.768 5.346 118.872 9.72 ; 
      RECT 118.336 5.346 118.44 9.72 ; 
      RECT 117.904 5.346 118.008 9.72 ; 
      RECT 117.472 5.346 117.576 9.72 ; 
      RECT 117.04 5.346 117.144 9.72 ; 
      RECT 116.608 5.346 116.712 9.72 ; 
      RECT 116.176 5.346 116.28 9.72 ; 
      RECT 115.744 5.346 115.848 9.72 ; 
      RECT 115.312 5.346 115.416 9.72 ; 
      RECT 114.88 5.346 114.984 9.72 ; 
      RECT 114.448 5.346 114.552 9.72 ; 
      RECT 114.016 5.346 114.12 9.72 ; 
      RECT 113.584 5.346 113.688 9.72 ; 
      RECT 113.152 5.346 113.256 9.72 ; 
      RECT 112.72 5.346 112.824 9.72 ; 
      RECT 112.288 5.346 112.392 9.72 ; 
      RECT 111.856 5.346 111.96 9.72 ; 
      RECT 111.424 5.346 111.528 9.72 ; 
      RECT 110.992 5.346 111.096 9.72 ; 
      RECT 110.56 5.346 110.664 9.72 ; 
      RECT 110.128 5.346 110.232 9.72 ; 
      RECT 109.696 5.346 109.8 9.72 ; 
      RECT 109.264 5.346 109.368 9.72 ; 
      RECT 108.832 5.346 108.936 9.72 ; 
      RECT 108.4 5.346 108.504 9.72 ; 
      RECT 107.968 5.346 108.072 9.72 ; 
      RECT 107.536 5.346 107.64 9.72 ; 
      RECT 107.104 5.346 107.208 9.72 ; 
      RECT 106.672 5.346 106.776 9.72 ; 
      RECT 106.24 5.346 106.344 9.72 ; 
      RECT 105.808 5.346 105.912 9.72 ; 
      RECT 105.376 5.346 105.48 9.72 ; 
      RECT 104.944 5.346 105.048 9.72 ; 
      RECT 104.512 5.346 104.616 9.72 ; 
      RECT 104.08 5.346 104.184 9.72 ; 
      RECT 103.648 5.346 103.752 9.72 ; 
      RECT 103.216 5.346 103.32 9.72 ; 
      RECT 102.784 5.346 102.888 9.72 ; 
      RECT 102.352 5.346 102.456 9.72 ; 
      RECT 101.92 5.346 102.024 9.72 ; 
      RECT 101.488 5.346 101.592 9.72 ; 
      RECT 101.056 5.346 101.16 9.72 ; 
      RECT 100.624 5.346 100.728 9.72 ; 
      RECT 100.192 5.346 100.296 9.72 ; 
      RECT 99.76 5.346 99.864 9.72 ; 
      RECT 99.328 5.346 99.432 9.72 ; 
      RECT 98.896 5.346 99 9.72 ; 
      RECT 98.464 5.346 98.568 9.72 ; 
      RECT 98.032 5.346 98.136 9.72 ; 
      RECT 97.6 5.346 97.704 9.72 ; 
      RECT 97.168 5.346 97.272 9.72 ; 
      RECT 96.736 5.346 96.84 9.72 ; 
      RECT 96.304 5.346 96.408 9.72 ; 
      RECT 95.872 5.346 95.976 9.72 ; 
      RECT 95.44 5.346 95.544 9.72 ; 
      RECT 95.008 5.346 95.112 9.72 ; 
      RECT 94.576 5.346 94.68 9.72 ; 
      RECT 94.144 5.346 94.248 9.72 ; 
      RECT 93.712 5.346 93.816 9.72 ; 
      RECT 93.28 5.346 93.384 9.72 ; 
      RECT 92.848 5.346 92.952 9.72 ; 
      RECT 92.416 5.346 92.52 9.72 ; 
      RECT 91.984 5.346 92.088 9.72 ; 
      RECT 91.552 5.346 91.656 9.72 ; 
      RECT 91.12 5.346 91.224 9.72 ; 
      RECT 90.688 5.346 90.792 9.72 ; 
      RECT 90.256 5.346 90.36 9.72 ; 
      RECT 89.824 5.346 89.928 9.72 ; 
      RECT 89.392 5.346 89.496 9.72 ; 
      RECT 88.96 5.346 89.064 9.72 ; 
      RECT 88.528 5.346 88.632 9.72 ; 
      RECT 88.096 5.346 88.2 9.72 ; 
      RECT 87.664 5.346 87.768 9.72 ; 
      RECT 87.232 5.346 87.336 9.72 ; 
      RECT 86.8 5.346 86.904 9.72 ; 
      RECT 86.368 5.346 86.472 9.72 ; 
      RECT 85.936 5.346 86.04 9.72 ; 
      RECT 85.504 5.346 85.608 9.72 ; 
      RECT 85.072 5.346 85.176 9.72 ; 
      RECT 84.64 5.346 84.744 9.72 ; 
      RECT 84.208 5.346 84.312 9.72 ; 
      RECT 83.776 5.346 83.88 9.72 ; 
      RECT 83.344 5.346 83.448 9.72 ; 
      RECT 82.912 5.346 83.016 9.72 ; 
      RECT 82.48 5.346 82.584 9.72 ; 
      RECT 82.048 5.346 82.152 9.72 ; 
      RECT 81.616 5.346 81.72 9.72 ; 
      RECT 81.184 5.346 81.288 9.72 ; 
      RECT 80.752 5.346 80.856 9.72 ; 
      RECT 80.32 5.346 80.424 9.72 ; 
      RECT 79.888 5.346 79.992 9.72 ; 
      RECT 79.456 5.346 79.56 9.72 ; 
      RECT 79.024 5.346 79.128 9.72 ; 
      RECT 78.592 5.346 78.696 9.72 ; 
      RECT 78.16 5.346 78.264 9.72 ; 
      RECT 77.728 5.346 77.832 9.72 ; 
      RECT 77.296 5.346 77.4 9.72 ; 
      RECT 76.864 5.346 76.968 9.72 ; 
      RECT 76.432 5.346 76.536 9.72 ; 
      RECT 76 5.346 76.104 9.72 ; 
      RECT 75.568 5.346 75.672 9.72 ; 
      RECT 75.136 5.346 75.24 9.72 ; 
      RECT 74.704 5.346 74.808 9.72 ; 
      RECT 74.272 5.346 74.376 9.72 ; 
      RECT 73.84 5.346 73.944 9.72 ; 
      RECT 73.408 5.346 73.512 9.72 ; 
      RECT 72.976 5.346 73.08 9.72 ; 
      RECT 72.544 5.346 72.648 9.72 ; 
      RECT 72.112 5.346 72.216 9.72 ; 
      RECT 71.68 5.346 71.784 9.72 ; 
      RECT 71.248 5.346 71.352 9.72 ; 
      RECT 70.816 5.346 70.92 9.72 ; 
      RECT 70.384 5.346 70.488 9.72 ; 
      RECT 69.952 5.346 70.056 9.72 ; 
      RECT 69.52 5.346 69.624 9.72 ; 
      RECT 69.088 5.346 69.192 9.72 ; 
      RECT 68.656 5.346 68.76 9.72 ; 
      RECT 68.224 5.346 68.328 9.72 ; 
      RECT 67.792 5.346 67.896 9.72 ; 
      RECT 67.36 5.346 67.464 9.72 ; 
      RECT 66.928 5.346 67.032 9.72 ; 
      RECT 66.496 5.346 66.6 9.72 ; 
      RECT 66.064 5.346 66.168 9.72 ; 
      RECT 65.632 5.346 65.736 9.72 ; 
      RECT 65.2 5.346 65.304 9.72 ; 
      RECT 64.348 5.346 64.656 9.72 ; 
      RECT 56.776 5.346 57.084 9.72 ; 
      RECT 56.128 5.346 56.232 9.72 ; 
      RECT 55.696 5.346 55.8 9.72 ; 
      RECT 55.264 5.346 55.368 9.72 ; 
      RECT 54.832 5.346 54.936 9.72 ; 
      RECT 54.4 5.346 54.504 9.72 ; 
      RECT 53.968 5.346 54.072 9.72 ; 
      RECT 53.536 5.346 53.64 9.72 ; 
      RECT 53.104 5.346 53.208 9.72 ; 
      RECT 52.672 5.346 52.776 9.72 ; 
      RECT 52.24 5.346 52.344 9.72 ; 
      RECT 51.808 5.346 51.912 9.72 ; 
      RECT 51.376 5.346 51.48 9.72 ; 
      RECT 50.944 5.346 51.048 9.72 ; 
      RECT 50.512 5.346 50.616 9.72 ; 
      RECT 50.08 5.346 50.184 9.72 ; 
      RECT 49.648 5.346 49.752 9.72 ; 
      RECT 49.216 5.346 49.32 9.72 ; 
      RECT 48.784 5.346 48.888 9.72 ; 
      RECT 48.352 5.346 48.456 9.72 ; 
      RECT 47.92 5.346 48.024 9.72 ; 
      RECT 47.488 5.346 47.592 9.72 ; 
      RECT 47.056 5.346 47.16 9.72 ; 
      RECT 46.624 5.346 46.728 9.72 ; 
      RECT 46.192 5.346 46.296 9.72 ; 
      RECT 45.76 5.346 45.864 9.72 ; 
      RECT 45.328 5.346 45.432 9.72 ; 
      RECT 44.896 5.346 45 9.72 ; 
      RECT 44.464 5.346 44.568 9.72 ; 
      RECT 44.032 5.346 44.136 9.72 ; 
      RECT 43.6 5.346 43.704 9.72 ; 
      RECT 43.168 5.346 43.272 9.72 ; 
      RECT 42.736 5.346 42.84 9.72 ; 
      RECT 42.304 5.346 42.408 9.72 ; 
      RECT 41.872 5.346 41.976 9.72 ; 
      RECT 41.44 5.346 41.544 9.72 ; 
      RECT 41.008 5.346 41.112 9.72 ; 
      RECT 40.576 5.346 40.68 9.72 ; 
      RECT 40.144 5.346 40.248 9.72 ; 
      RECT 39.712 5.346 39.816 9.72 ; 
      RECT 39.28 5.346 39.384 9.72 ; 
      RECT 38.848 5.346 38.952 9.72 ; 
      RECT 38.416 5.346 38.52 9.72 ; 
      RECT 37.984 5.346 38.088 9.72 ; 
      RECT 37.552 5.346 37.656 9.72 ; 
      RECT 37.12 5.346 37.224 9.72 ; 
      RECT 36.688 5.346 36.792 9.72 ; 
      RECT 36.256 5.346 36.36 9.72 ; 
      RECT 35.824 5.346 35.928 9.72 ; 
      RECT 35.392 5.346 35.496 9.72 ; 
      RECT 34.96 5.346 35.064 9.72 ; 
      RECT 34.528 5.346 34.632 9.72 ; 
      RECT 34.096 5.346 34.2 9.72 ; 
      RECT 33.664 5.346 33.768 9.72 ; 
      RECT 33.232 5.346 33.336 9.72 ; 
      RECT 32.8 5.346 32.904 9.72 ; 
      RECT 32.368 5.346 32.472 9.72 ; 
      RECT 31.936 5.346 32.04 9.72 ; 
      RECT 31.504 5.346 31.608 9.72 ; 
      RECT 31.072 5.346 31.176 9.72 ; 
      RECT 30.64 5.346 30.744 9.72 ; 
      RECT 30.208 5.346 30.312 9.72 ; 
      RECT 29.776 5.346 29.88 9.72 ; 
      RECT 29.344 5.346 29.448 9.72 ; 
      RECT 28.912 5.346 29.016 9.72 ; 
      RECT 28.48 5.346 28.584 9.72 ; 
      RECT 28.048 5.346 28.152 9.72 ; 
      RECT 27.616 5.346 27.72 9.72 ; 
      RECT 27.184 5.346 27.288 9.72 ; 
      RECT 26.752 5.346 26.856 9.72 ; 
      RECT 26.32 5.346 26.424 9.72 ; 
      RECT 25.888 5.346 25.992 9.72 ; 
      RECT 25.456 5.346 25.56 9.72 ; 
      RECT 25.024 5.346 25.128 9.72 ; 
      RECT 24.592 5.346 24.696 9.72 ; 
      RECT 24.16 5.346 24.264 9.72 ; 
      RECT 23.728 5.346 23.832 9.72 ; 
      RECT 23.296 5.346 23.4 9.72 ; 
      RECT 22.864 5.346 22.968 9.72 ; 
      RECT 22.432 5.346 22.536 9.72 ; 
      RECT 22 5.346 22.104 9.72 ; 
      RECT 21.568 5.346 21.672 9.72 ; 
      RECT 21.136 5.346 21.24 9.72 ; 
      RECT 20.704 5.346 20.808 9.72 ; 
      RECT 20.272 5.346 20.376 9.72 ; 
      RECT 19.84 5.346 19.944 9.72 ; 
      RECT 19.408 5.346 19.512 9.72 ; 
      RECT 18.976 5.346 19.08 9.72 ; 
      RECT 18.544 5.346 18.648 9.72 ; 
      RECT 18.112 5.346 18.216 9.72 ; 
      RECT 17.68 5.346 17.784 9.72 ; 
      RECT 17.248 5.346 17.352 9.72 ; 
      RECT 16.816 5.346 16.92 9.72 ; 
      RECT 16.384 5.346 16.488 9.72 ; 
      RECT 15.952 5.346 16.056 9.72 ; 
      RECT 15.52 5.346 15.624 9.72 ; 
      RECT 15.088 5.346 15.192 9.72 ; 
      RECT 14.656 5.346 14.76 9.72 ; 
      RECT 14.224 5.346 14.328 9.72 ; 
      RECT 13.792 5.346 13.896 9.72 ; 
      RECT 13.36 5.346 13.464 9.72 ; 
      RECT 12.928 5.346 13.032 9.72 ; 
      RECT 12.496 5.346 12.6 9.72 ; 
      RECT 12.064 5.346 12.168 9.72 ; 
      RECT 11.632 5.346 11.736 9.72 ; 
      RECT 11.2 5.346 11.304 9.72 ; 
      RECT 10.768 5.346 10.872 9.72 ; 
      RECT 10.336 5.346 10.44 9.72 ; 
      RECT 9.904 5.346 10.008 9.72 ; 
      RECT 9.472 5.346 9.576 9.72 ; 
      RECT 9.04 5.346 9.144 9.72 ; 
      RECT 8.608 5.346 8.712 9.72 ; 
      RECT 8.176 5.346 8.28 9.72 ; 
      RECT 7.744 5.346 7.848 9.72 ; 
      RECT 7.312 5.346 7.416 9.72 ; 
      RECT 6.88 5.346 6.984 9.72 ; 
      RECT 6.448 5.346 6.552 9.72 ; 
      RECT 6.016 5.346 6.12 9.72 ; 
      RECT 5.584 5.346 5.688 9.72 ; 
      RECT 5.152 5.346 5.256 9.72 ; 
      RECT 4.72 5.346 4.824 9.72 ; 
      RECT 4.288 5.346 4.392 9.72 ; 
      RECT 3.856 5.346 3.96 9.72 ; 
      RECT 3.424 5.346 3.528 9.72 ; 
      RECT 2.992 5.346 3.096 9.72 ; 
      RECT 2.56 5.346 2.664 9.72 ; 
      RECT 2.128 5.346 2.232 9.72 ; 
      RECT 1.696 5.346 1.8 9.72 ; 
      RECT 1.264 5.346 1.368 9.72 ; 
      RECT 0.832 5.346 0.936 9.72 ; 
      RECT 0.02 5.346 0.36 9.72 ; 
      RECT 62.212 9.666 62.724 14.04 ; 
      RECT 62.156 12.328 62.724 13.618 ; 
      RECT 61.276 11.236 61.812 14.04 ; 
      RECT 61.184 12.576 61.812 13.608 ; 
      RECT 61.276 9.666 61.668 14.04 ; 
      RECT 61.276 10.15 61.724 11.108 ; 
      RECT 61.276 9.666 61.812 10.022 ; 
      RECT 60.376 11.468 60.912 14.04 ; 
      RECT 60.376 9.666 60.768 14.04 ; 
      RECT 58.708 9.666 59.04 14.04 ; 
      RECT 58.708 10.02 59.096 13.762 ; 
      RECT 121.072 9.666 121.412 14.04 ; 
      RECT 120.496 9.666 120.6 14.04 ; 
      RECT 120.064 9.666 120.168 14.04 ; 
      RECT 119.632 9.666 119.736 14.04 ; 
      RECT 119.2 9.666 119.304 14.04 ; 
      RECT 118.768 9.666 118.872 14.04 ; 
      RECT 118.336 9.666 118.44 14.04 ; 
      RECT 117.904 9.666 118.008 14.04 ; 
      RECT 117.472 9.666 117.576 14.04 ; 
      RECT 117.04 9.666 117.144 14.04 ; 
      RECT 116.608 9.666 116.712 14.04 ; 
      RECT 116.176 9.666 116.28 14.04 ; 
      RECT 115.744 9.666 115.848 14.04 ; 
      RECT 115.312 9.666 115.416 14.04 ; 
      RECT 114.88 9.666 114.984 14.04 ; 
      RECT 114.448 9.666 114.552 14.04 ; 
      RECT 114.016 9.666 114.12 14.04 ; 
      RECT 113.584 9.666 113.688 14.04 ; 
      RECT 113.152 9.666 113.256 14.04 ; 
      RECT 112.72 9.666 112.824 14.04 ; 
      RECT 112.288 9.666 112.392 14.04 ; 
      RECT 111.856 9.666 111.96 14.04 ; 
      RECT 111.424 9.666 111.528 14.04 ; 
      RECT 110.992 9.666 111.096 14.04 ; 
      RECT 110.56 9.666 110.664 14.04 ; 
      RECT 110.128 9.666 110.232 14.04 ; 
      RECT 109.696 9.666 109.8 14.04 ; 
      RECT 109.264 9.666 109.368 14.04 ; 
      RECT 108.832 9.666 108.936 14.04 ; 
      RECT 108.4 9.666 108.504 14.04 ; 
      RECT 107.968 9.666 108.072 14.04 ; 
      RECT 107.536 9.666 107.64 14.04 ; 
      RECT 107.104 9.666 107.208 14.04 ; 
      RECT 106.672 9.666 106.776 14.04 ; 
      RECT 106.24 9.666 106.344 14.04 ; 
      RECT 105.808 9.666 105.912 14.04 ; 
      RECT 105.376 9.666 105.48 14.04 ; 
      RECT 104.944 9.666 105.048 14.04 ; 
      RECT 104.512 9.666 104.616 14.04 ; 
      RECT 104.08 9.666 104.184 14.04 ; 
      RECT 103.648 9.666 103.752 14.04 ; 
      RECT 103.216 9.666 103.32 14.04 ; 
      RECT 102.784 9.666 102.888 14.04 ; 
      RECT 102.352 9.666 102.456 14.04 ; 
      RECT 101.92 9.666 102.024 14.04 ; 
      RECT 101.488 9.666 101.592 14.04 ; 
      RECT 101.056 9.666 101.16 14.04 ; 
      RECT 100.624 9.666 100.728 14.04 ; 
      RECT 100.192 9.666 100.296 14.04 ; 
      RECT 99.76 9.666 99.864 14.04 ; 
      RECT 99.328 9.666 99.432 14.04 ; 
      RECT 98.896 9.666 99 14.04 ; 
      RECT 98.464 9.666 98.568 14.04 ; 
      RECT 98.032 9.666 98.136 14.04 ; 
      RECT 97.6 9.666 97.704 14.04 ; 
      RECT 97.168 9.666 97.272 14.04 ; 
      RECT 96.736 9.666 96.84 14.04 ; 
      RECT 96.304 9.666 96.408 14.04 ; 
      RECT 95.872 9.666 95.976 14.04 ; 
      RECT 95.44 9.666 95.544 14.04 ; 
      RECT 95.008 9.666 95.112 14.04 ; 
      RECT 94.576 9.666 94.68 14.04 ; 
      RECT 94.144 9.666 94.248 14.04 ; 
      RECT 93.712 9.666 93.816 14.04 ; 
      RECT 93.28 9.666 93.384 14.04 ; 
      RECT 92.848 9.666 92.952 14.04 ; 
      RECT 92.416 9.666 92.52 14.04 ; 
      RECT 91.984 9.666 92.088 14.04 ; 
      RECT 91.552 9.666 91.656 14.04 ; 
      RECT 91.12 9.666 91.224 14.04 ; 
      RECT 90.688 9.666 90.792 14.04 ; 
      RECT 90.256 9.666 90.36 14.04 ; 
      RECT 89.824 9.666 89.928 14.04 ; 
      RECT 89.392 9.666 89.496 14.04 ; 
      RECT 88.96 9.666 89.064 14.04 ; 
      RECT 88.528 9.666 88.632 14.04 ; 
      RECT 88.096 9.666 88.2 14.04 ; 
      RECT 87.664 9.666 87.768 14.04 ; 
      RECT 87.232 9.666 87.336 14.04 ; 
      RECT 86.8 9.666 86.904 14.04 ; 
      RECT 86.368 9.666 86.472 14.04 ; 
      RECT 85.936 9.666 86.04 14.04 ; 
      RECT 85.504 9.666 85.608 14.04 ; 
      RECT 85.072 9.666 85.176 14.04 ; 
      RECT 84.64 9.666 84.744 14.04 ; 
      RECT 84.208 9.666 84.312 14.04 ; 
      RECT 83.776 9.666 83.88 14.04 ; 
      RECT 83.344 9.666 83.448 14.04 ; 
      RECT 82.912 9.666 83.016 14.04 ; 
      RECT 82.48 9.666 82.584 14.04 ; 
      RECT 82.048 9.666 82.152 14.04 ; 
      RECT 81.616 9.666 81.72 14.04 ; 
      RECT 81.184 9.666 81.288 14.04 ; 
      RECT 80.752 9.666 80.856 14.04 ; 
      RECT 80.32 9.666 80.424 14.04 ; 
      RECT 79.888 9.666 79.992 14.04 ; 
      RECT 79.456 9.666 79.56 14.04 ; 
      RECT 79.024 9.666 79.128 14.04 ; 
      RECT 78.592 9.666 78.696 14.04 ; 
      RECT 78.16 9.666 78.264 14.04 ; 
      RECT 77.728 9.666 77.832 14.04 ; 
      RECT 77.296 9.666 77.4 14.04 ; 
      RECT 76.864 9.666 76.968 14.04 ; 
      RECT 76.432 9.666 76.536 14.04 ; 
      RECT 76 9.666 76.104 14.04 ; 
      RECT 75.568 9.666 75.672 14.04 ; 
      RECT 75.136 9.666 75.24 14.04 ; 
      RECT 74.704 9.666 74.808 14.04 ; 
      RECT 74.272 9.666 74.376 14.04 ; 
      RECT 73.84 9.666 73.944 14.04 ; 
      RECT 73.408 9.666 73.512 14.04 ; 
      RECT 72.976 9.666 73.08 14.04 ; 
      RECT 72.544 9.666 72.648 14.04 ; 
      RECT 72.112 9.666 72.216 14.04 ; 
      RECT 71.68 9.666 71.784 14.04 ; 
      RECT 71.248 9.666 71.352 14.04 ; 
      RECT 70.816 9.666 70.92 14.04 ; 
      RECT 70.384 9.666 70.488 14.04 ; 
      RECT 69.952 9.666 70.056 14.04 ; 
      RECT 69.52 9.666 69.624 14.04 ; 
      RECT 69.088 9.666 69.192 14.04 ; 
      RECT 68.656 9.666 68.76 14.04 ; 
      RECT 68.224 9.666 68.328 14.04 ; 
      RECT 67.792 9.666 67.896 14.04 ; 
      RECT 67.36 9.666 67.464 14.04 ; 
      RECT 66.928 9.666 67.032 14.04 ; 
      RECT 66.496 9.666 66.6 14.04 ; 
      RECT 66.064 9.666 66.168 14.04 ; 
      RECT 65.632 9.666 65.736 14.04 ; 
      RECT 65.2 9.666 65.304 14.04 ; 
      RECT 64.348 9.666 64.656 14.04 ; 
      RECT 56.776 9.666 57.084 14.04 ; 
      RECT 56.128 9.666 56.232 14.04 ; 
      RECT 55.696 9.666 55.8 14.04 ; 
      RECT 55.264 9.666 55.368 14.04 ; 
      RECT 54.832 9.666 54.936 14.04 ; 
      RECT 54.4 9.666 54.504 14.04 ; 
      RECT 53.968 9.666 54.072 14.04 ; 
      RECT 53.536 9.666 53.64 14.04 ; 
      RECT 53.104 9.666 53.208 14.04 ; 
      RECT 52.672 9.666 52.776 14.04 ; 
      RECT 52.24 9.666 52.344 14.04 ; 
      RECT 51.808 9.666 51.912 14.04 ; 
      RECT 51.376 9.666 51.48 14.04 ; 
      RECT 50.944 9.666 51.048 14.04 ; 
      RECT 50.512 9.666 50.616 14.04 ; 
      RECT 50.08 9.666 50.184 14.04 ; 
      RECT 49.648 9.666 49.752 14.04 ; 
      RECT 49.216 9.666 49.32 14.04 ; 
      RECT 48.784 9.666 48.888 14.04 ; 
      RECT 48.352 9.666 48.456 14.04 ; 
      RECT 47.92 9.666 48.024 14.04 ; 
      RECT 47.488 9.666 47.592 14.04 ; 
      RECT 47.056 9.666 47.16 14.04 ; 
      RECT 46.624 9.666 46.728 14.04 ; 
      RECT 46.192 9.666 46.296 14.04 ; 
      RECT 45.76 9.666 45.864 14.04 ; 
      RECT 45.328 9.666 45.432 14.04 ; 
      RECT 44.896 9.666 45 14.04 ; 
      RECT 44.464 9.666 44.568 14.04 ; 
      RECT 44.032 9.666 44.136 14.04 ; 
      RECT 43.6 9.666 43.704 14.04 ; 
      RECT 43.168 9.666 43.272 14.04 ; 
      RECT 42.736 9.666 42.84 14.04 ; 
      RECT 42.304 9.666 42.408 14.04 ; 
      RECT 41.872 9.666 41.976 14.04 ; 
      RECT 41.44 9.666 41.544 14.04 ; 
      RECT 41.008 9.666 41.112 14.04 ; 
      RECT 40.576 9.666 40.68 14.04 ; 
      RECT 40.144 9.666 40.248 14.04 ; 
      RECT 39.712 9.666 39.816 14.04 ; 
      RECT 39.28 9.666 39.384 14.04 ; 
      RECT 38.848 9.666 38.952 14.04 ; 
      RECT 38.416 9.666 38.52 14.04 ; 
      RECT 37.984 9.666 38.088 14.04 ; 
      RECT 37.552 9.666 37.656 14.04 ; 
      RECT 37.12 9.666 37.224 14.04 ; 
      RECT 36.688 9.666 36.792 14.04 ; 
      RECT 36.256 9.666 36.36 14.04 ; 
      RECT 35.824 9.666 35.928 14.04 ; 
      RECT 35.392 9.666 35.496 14.04 ; 
      RECT 34.96 9.666 35.064 14.04 ; 
      RECT 34.528 9.666 34.632 14.04 ; 
      RECT 34.096 9.666 34.2 14.04 ; 
      RECT 33.664 9.666 33.768 14.04 ; 
      RECT 33.232 9.666 33.336 14.04 ; 
      RECT 32.8 9.666 32.904 14.04 ; 
      RECT 32.368 9.666 32.472 14.04 ; 
      RECT 31.936 9.666 32.04 14.04 ; 
      RECT 31.504 9.666 31.608 14.04 ; 
      RECT 31.072 9.666 31.176 14.04 ; 
      RECT 30.64 9.666 30.744 14.04 ; 
      RECT 30.208 9.666 30.312 14.04 ; 
      RECT 29.776 9.666 29.88 14.04 ; 
      RECT 29.344 9.666 29.448 14.04 ; 
      RECT 28.912 9.666 29.016 14.04 ; 
      RECT 28.48 9.666 28.584 14.04 ; 
      RECT 28.048 9.666 28.152 14.04 ; 
      RECT 27.616 9.666 27.72 14.04 ; 
      RECT 27.184 9.666 27.288 14.04 ; 
      RECT 26.752 9.666 26.856 14.04 ; 
      RECT 26.32 9.666 26.424 14.04 ; 
      RECT 25.888 9.666 25.992 14.04 ; 
      RECT 25.456 9.666 25.56 14.04 ; 
      RECT 25.024 9.666 25.128 14.04 ; 
      RECT 24.592 9.666 24.696 14.04 ; 
      RECT 24.16 9.666 24.264 14.04 ; 
      RECT 23.728 9.666 23.832 14.04 ; 
      RECT 23.296 9.666 23.4 14.04 ; 
      RECT 22.864 9.666 22.968 14.04 ; 
      RECT 22.432 9.666 22.536 14.04 ; 
      RECT 22 9.666 22.104 14.04 ; 
      RECT 21.568 9.666 21.672 14.04 ; 
      RECT 21.136 9.666 21.24 14.04 ; 
      RECT 20.704 9.666 20.808 14.04 ; 
      RECT 20.272 9.666 20.376 14.04 ; 
      RECT 19.84 9.666 19.944 14.04 ; 
      RECT 19.408 9.666 19.512 14.04 ; 
      RECT 18.976 9.666 19.08 14.04 ; 
      RECT 18.544 9.666 18.648 14.04 ; 
      RECT 18.112 9.666 18.216 14.04 ; 
      RECT 17.68 9.666 17.784 14.04 ; 
      RECT 17.248 9.666 17.352 14.04 ; 
      RECT 16.816 9.666 16.92 14.04 ; 
      RECT 16.384 9.666 16.488 14.04 ; 
      RECT 15.952 9.666 16.056 14.04 ; 
      RECT 15.52 9.666 15.624 14.04 ; 
      RECT 15.088 9.666 15.192 14.04 ; 
      RECT 14.656 9.666 14.76 14.04 ; 
      RECT 14.224 9.666 14.328 14.04 ; 
      RECT 13.792 9.666 13.896 14.04 ; 
      RECT 13.36 9.666 13.464 14.04 ; 
      RECT 12.928 9.666 13.032 14.04 ; 
      RECT 12.496 9.666 12.6 14.04 ; 
      RECT 12.064 9.666 12.168 14.04 ; 
      RECT 11.632 9.666 11.736 14.04 ; 
      RECT 11.2 9.666 11.304 14.04 ; 
      RECT 10.768 9.666 10.872 14.04 ; 
      RECT 10.336 9.666 10.44 14.04 ; 
      RECT 9.904 9.666 10.008 14.04 ; 
      RECT 9.472 9.666 9.576 14.04 ; 
      RECT 9.04 9.666 9.144 14.04 ; 
      RECT 8.608 9.666 8.712 14.04 ; 
      RECT 8.176 9.666 8.28 14.04 ; 
      RECT 7.744 9.666 7.848 14.04 ; 
      RECT 7.312 9.666 7.416 14.04 ; 
      RECT 6.88 9.666 6.984 14.04 ; 
      RECT 6.448 9.666 6.552 14.04 ; 
      RECT 6.016 9.666 6.12 14.04 ; 
      RECT 5.584 9.666 5.688 14.04 ; 
      RECT 5.152 9.666 5.256 14.04 ; 
      RECT 4.72 9.666 4.824 14.04 ; 
      RECT 4.288 9.666 4.392 14.04 ; 
      RECT 3.856 9.666 3.96 14.04 ; 
      RECT 3.424 9.666 3.528 14.04 ; 
      RECT 2.992 9.666 3.096 14.04 ; 
      RECT 2.56 9.666 2.664 14.04 ; 
      RECT 2.128 9.666 2.232 14.04 ; 
      RECT 1.696 9.666 1.8 14.04 ; 
      RECT 1.264 9.666 1.368 14.04 ; 
      RECT 0.832 9.666 0.936 14.04 ; 
      RECT 0.02 9.666 0.36 14.04 ; 
      RECT 62.212 13.986 62.724 18.36 ; 
      RECT 62.156 16.648 62.724 17.938 ; 
      RECT 61.276 15.556 61.812 18.36 ; 
      RECT 61.184 16.896 61.812 17.928 ; 
      RECT 61.276 13.986 61.668 18.36 ; 
      RECT 61.276 14.47 61.724 15.428 ; 
      RECT 61.276 13.986 61.812 14.342 ; 
      RECT 60.376 15.788 60.912 18.36 ; 
      RECT 60.376 13.986 60.768 18.36 ; 
      RECT 58.708 13.986 59.04 18.36 ; 
      RECT 58.708 14.34 59.096 18.082 ; 
      RECT 121.072 13.986 121.412 18.36 ; 
      RECT 120.496 13.986 120.6 18.36 ; 
      RECT 120.064 13.986 120.168 18.36 ; 
      RECT 119.632 13.986 119.736 18.36 ; 
      RECT 119.2 13.986 119.304 18.36 ; 
      RECT 118.768 13.986 118.872 18.36 ; 
      RECT 118.336 13.986 118.44 18.36 ; 
      RECT 117.904 13.986 118.008 18.36 ; 
      RECT 117.472 13.986 117.576 18.36 ; 
      RECT 117.04 13.986 117.144 18.36 ; 
      RECT 116.608 13.986 116.712 18.36 ; 
      RECT 116.176 13.986 116.28 18.36 ; 
      RECT 115.744 13.986 115.848 18.36 ; 
      RECT 115.312 13.986 115.416 18.36 ; 
      RECT 114.88 13.986 114.984 18.36 ; 
      RECT 114.448 13.986 114.552 18.36 ; 
      RECT 114.016 13.986 114.12 18.36 ; 
      RECT 113.584 13.986 113.688 18.36 ; 
      RECT 113.152 13.986 113.256 18.36 ; 
      RECT 112.72 13.986 112.824 18.36 ; 
      RECT 112.288 13.986 112.392 18.36 ; 
      RECT 111.856 13.986 111.96 18.36 ; 
      RECT 111.424 13.986 111.528 18.36 ; 
      RECT 110.992 13.986 111.096 18.36 ; 
      RECT 110.56 13.986 110.664 18.36 ; 
      RECT 110.128 13.986 110.232 18.36 ; 
      RECT 109.696 13.986 109.8 18.36 ; 
      RECT 109.264 13.986 109.368 18.36 ; 
      RECT 108.832 13.986 108.936 18.36 ; 
      RECT 108.4 13.986 108.504 18.36 ; 
      RECT 107.968 13.986 108.072 18.36 ; 
      RECT 107.536 13.986 107.64 18.36 ; 
      RECT 107.104 13.986 107.208 18.36 ; 
      RECT 106.672 13.986 106.776 18.36 ; 
      RECT 106.24 13.986 106.344 18.36 ; 
      RECT 105.808 13.986 105.912 18.36 ; 
      RECT 105.376 13.986 105.48 18.36 ; 
      RECT 104.944 13.986 105.048 18.36 ; 
      RECT 104.512 13.986 104.616 18.36 ; 
      RECT 104.08 13.986 104.184 18.36 ; 
      RECT 103.648 13.986 103.752 18.36 ; 
      RECT 103.216 13.986 103.32 18.36 ; 
      RECT 102.784 13.986 102.888 18.36 ; 
      RECT 102.352 13.986 102.456 18.36 ; 
      RECT 101.92 13.986 102.024 18.36 ; 
      RECT 101.488 13.986 101.592 18.36 ; 
      RECT 101.056 13.986 101.16 18.36 ; 
      RECT 100.624 13.986 100.728 18.36 ; 
      RECT 100.192 13.986 100.296 18.36 ; 
      RECT 99.76 13.986 99.864 18.36 ; 
      RECT 99.328 13.986 99.432 18.36 ; 
      RECT 98.896 13.986 99 18.36 ; 
      RECT 98.464 13.986 98.568 18.36 ; 
      RECT 98.032 13.986 98.136 18.36 ; 
      RECT 97.6 13.986 97.704 18.36 ; 
      RECT 97.168 13.986 97.272 18.36 ; 
      RECT 96.736 13.986 96.84 18.36 ; 
      RECT 96.304 13.986 96.408 18.36 ; 
      RECT 95.872 13.986 95.976 18.36 ; 
      RECT 95.44 13.986 95.544 18.36 ; 
      RECT 95.008 13.986 95.112 18.36 ; 
      RECT 94.576 13.986 94.68 18.36 ; 
      RECT 94.144 13.986 94.248 18.36 ; 
      RECT 93.712 13.986 93.816 18.36 ; 
      RECT 93.28 13.986 93.384 18.36 ; 
      RECT 92.848 13.986 92.952 18.36 ; 
      RECT 92.416 13.986 92.52 18.36 ; 
      RECT 91.984 13.986 92.088 18.36 ; 
      RECT 91.552 13.986 91.656 18.36 ; 
      RECT 91.12 13.986 91.224 18.36 ; 
      RECT 90.688 13.986 90.792 18.36 ; 
      RECT 90.256 13.986 90.36 18.36 ; 
      RECT 89.824 13.986 89.928 18.36 ; 
      RECT 89.392 13.986 89.496 18.36 ; 
      RECT 88.96 13.986 89.064 18.36 ; 
      RECT 88.528 13.986 88.632 18.36 ; 
      RECT 88.096 13.986 88.2 18.36 ; 
      RECT 87.664 13.986 87.768 18.36 ; 
      RECT 87.232 13.986 87.336 18.36 ; 
      RECT 86.8 13.986 86.904 18.36 ; 
      RECT 86.368 13.986 86.472 18.36 ; 
      RECT 85.936 13.986 86.04 18.36 ; 
      RECT 85.504 13.986 85.608 18.36 ; 
      RECT 85.072 13.986 85.176 18.36 ; 
      RECT 84.64 13.986 84.744 18.36 ; 
      RECT 84.208 13.986 84.312 18.36 ; 
      RECT 83.776 13.986 83.88 18.36 ; 
      RECT 83.344 13.986 83.448 18.36 ; 
      RECT 82.912 13.986 83.016 18.36 ; 
      RECT 82.48 13.986 82.584 18.36 ; 
      RECT 82.048 13.986 82.152 18.36 ; 
      RECT 81.616 13.986 81.72 18.36 ; 
      RECT 81.184 13.986 81.288 18.36 ; 
      RECT 80.752 13.986 80.856 18.36 ; 
      RECT 80.32 13.986 80.424 18.36 ; 
      RECT 79.888 13.986 79.992 18.36 ; 
      RECT 79.456 13.986 79.56 18.36 ; 
      RECT 79.024 13.986 79.128 18.36 ; 
      RECT 78.592 13.986 78.696 18.36 ; 
      RECT 78.16 13.986 78.264 18.36 ; 
      RECT 77.728 13.986 77.832 18.36 ; 
      RECT 77.296 13.986 77.4 18.36 ; 
      RECT 76.864 13.986 76.968 18.36 ; 
      RECT 76.432 13.986 76.536 18.36 ; 
      RECT 76 13.986 76.104 18.36 ; 
      RECT 75.568 13.986 75.672 18.36 ; 
      RECT 75.136 13.986 75.24 18.36 ; 
      RECT 74.704 13.986 74.808 18.36 ; 
      RECT 74.272 13.986 74.376 18.36 ; 
      RECT 73.84 13.986 73.944 18.36 ; 
      RECT 73.408 13.986 73.512 18.36 ; 
      RECT 72.976 13.986 73.08 18.36 ; 
      RECT 72.544 13.986 72.648 18.36 ; 
      RECT 72.112 13.986 72.216 18.36 ; 
      RECT 71.68 13.986 71.784 18.36 ; 
      RECT 71.248 13.986 71.352 18.36 ; 
      RECT 70.816 13.986 70.92 18.36 ; 
      RECT 70.384 13.986 70.488 18.36 ; 
      RECT 69.952 13.986 70.056 18.36 ; 
      RECT 69.52 13.986 69.624 18.36 ; 
      RECT 69.088 13.986 69.192 18.36 ; 
      RECT 68.656 13.986 68.76 18.36 ; 
      RECT 68.224 13.986 68.328 18.36 ; 
      RECT 67.792 13.986 67.896 18.36 ; 
      RECT 67.36 13.986 67.464 18.36 ; 
      RECT 66.928 13.986 67.032 18.36 ; 
      RECT 66.496 13.986 66.6 18.36 ; 
      RECT 66.064 13.986 66.168 18.36 ; 
      RECT 65.632 13.986 65.736 18.36 ; 
      RECT 65.2 13.986 65.304 18.36 ; 
      RECT 64.348 13.986 64.656 18.36 ; 
      RECT 56.776 13.986 57.084 18.36 ; 
      RECT 56.128 13.986 56.232 18.36 ; 
      RECT 55.696 13.986 55.8 18.36 ; 
      RECT 55.264 13.986 55.368 18.36 ; 
      RECT 54.832 13.986 54.936 18.36 ; 
      RECT 54.4 13.986 54.504 18.36 ; 
      RECT 53.968 13.986 54.072 18.36 ; 
      RECT 53.536 13.986 53.64 18.36 ; 
      RECT 53.104 13.986 53.208 18.36 ; 
      RECT 52.672 13.986 52.776 18.36 ; 
      RECT 52.24 13.986 52.344 18.36 ; 
      RECT 51.808 13.986 51.912 18.36 ; 
      RECT 51.376 13.986 51.48 18.36 ; 
      RECT 50.944 13.986 51.048 18.36 ; 
      RECT 50.512 13.986 50.616 18.36 ; 
      RECT 50.08 13.986 50.184 18.36 ; 
      RECT 49.648 13.986 49.752 18.36 ; 
      RECT 49.216 13.986 49.32 18.36 ; 
      RECT 48.784 13.986 48.888 18.36 ; 
      RECT 48.352 13.986 48.456 18.36 ; 
      RECT 47.92 13.986 48.024 18.36 ; 
      RECT 47.488 13.986 47.592 18.36 ; 
      RECT 47.056 13.986 47.16 18.36 ; 
      RECT 46.624 13.986 46.728 18.36 ; 
      RECT 46.192 13.986 46.296 18.36 ; 
      RECT 45.76 13.986 45.864 18.36 ; 
      RECT 45.328 13.986 45.432 18.36 ; 
      RECT 44.896 13.986 45 18.36 ; 
      RECT 44.464 13.986 44.568 18.36 ; 
      RECT 44.032 13.986 44.136 18.36 ; 
      RECT 43.6 13.986 43.704 18.36 ; 
      RECT 43.168 13.986 43.272 18.36 ; 
      RECT 42.736 13.986 42.84 18.36 ; 
      RECT 42.304 13.986 42.408 18.36 ; 
      RECT 41.872 13.986 41.976 18.36 ; 
      RECT 41.44 13.986 41.544 18.36 ; 
      RECT 41.008 13.986 41.112 18.36 ; 
      RECT 40.576 13.986 40.68 18.36 ; 
      RECT 40.144 13.986 40.248 18.36 ; 
      RECT 39.712 13.986 39.816 18.36 ; 
      RECT 39.28 13.986 39.384 18.36 ; 
      RECT 38.848 13.986 38.952 18.36 ; 
      RECT 38.416 13.986 38.52 18.36 ; 
      RECT 37.984 13.986 38.088 18.36 ; 
      RECT 37.552 13.986 37.656 18.36 ; 
      RECT 37.12 13.986 37.224 18.36 ; 
      RECT 36.688 13.986 36.792 18.36 ; 
      RECT 36.256 13.986 36.36 18.36 ; 
      RECT 35.824 13.986 35.928 18.36 ; 
      RECT 35.392 13.986 35.496 18.36 ; 
      RECT 34.96 13.986 35.064 18.36 ; 
      RECT 34.528 13.986 34.632 18.36 ; 
      RECT 34.096 13.986 34.2 18.36 ; 
      RECT 33.664 13.986 33.768 18.36 ; 
      RECT 33.232 13.986 33.336 18.36 ; 
      RECT 32.8 13.986 32.904 18.36 ; 
      RECT 32.368 13.986 32.472 18.36 ; 
      RECT 31.936 13.986 32.04 18.36 ; 
      RECT 31.504 13.986 31.608 18.36 ; 
      RECT 31.072 13.986 31.176 18.36 ; 
      RECT 30.64 13.986 30.744 18.36 ; 
      RECT 30.208 13.986 30.312 18.36 ; 
      RECT 29.776 13.986 29.88 18.36 ; 
      RECT 29.344 13.986 29.448 18.36 ; 
      RECT 28.912 13.986 29.016 18.36 ; 
      RECT 28.48 13.986 28.584 18.36 ; 
      RECT 28.048 13.986 28.152 18.36 ; 
      RECT 27.616 13.986 27.72 18.36 ; 
      RECT 27.184 13.986 27.288 18.36 ; 
      RECT 26.752 13.986 26.856 18.36 ; 
      RECT 26.32 13.986 26.424 18.36 ; 
      RECT 25.888 13.986 25.992 18.36 ; 
      RECT 25.456 13.986 25.56 18.36 ; 
      RECT 25.024 13.986 25.128 18.36 ; 
      RECT 24.592 13.986 24.696 18.36 ; 
      RECT 24.16 13.986 24.264 18.36 ; 
      RECT 23.728 13.986 23.832 18.36 ; 
      RECT 23.296 13.986 23.4 18.36 ; 
      RECT 22.864 13.986 22.968 18.36 ; 
      RECT 22.432 13.986 22.536 18.36 ; 
      RECT 22 13.986 22.104 18.36 ; 
      RECT 21.568 13.986 21.672 18.36 ; 
      RECT 21.136 13.986 21.24 18.36 ; 
      RECT 20.704 13.986 20.808 18.36 ; 
      RECT 20.272 13.986 20.376 18.36 ; 
      RECT 19.84 13.986 19.944 18.36 ; 
      RECT 19.408 13.986 19.512 18.36 ; 
      RECT 18.976 13.986 19.08 18.36 ; 
      RECT 18.544 13.986 18.648 18.36 ; 
      RECT 18.112 13.986 18.216 18.36 ; 
      RECT 17.68 13.986 17.784 18.36 ; 
      RECT 17.248 13.986 17.352 18.36 ; 
      RECT 16.816 13.986 16.92 18.36 ; 
      RECT 16.384 13.986 16.488 18.36 ; 
      RECT 15.952 13.986 16.056 18.36 ; 
      RECT 15.52 13.986 15.624 18.36 ; 
      RECT 15.088 13.986 15.192 18.36 ; 
      RECT 14.656 13.986 14.76 18.36 ; 
      RECT 14.224 13.986 14.328 18.36 ; 
      RECT 13.792 13.986 13.896 18.36 ; 
      RECT 13.36 13.986 13.464 18.36 ; 
      RECT 12.928 13.986 13.032 18.36 ; 
      RECT 12.496 13.986 12.6 18.36 ; 
      RECT 12.064 13.986 12.168 18.36 ; 
      RECT 11.632 13.986 11.736 18.36 ; 
      RECT 11.2 13.986 11.304 18.36 ; 
      RECT 10.768 13.986 10.872 18.36 ; 
      RECT 10.336 13.986 10.44 18.36 ; 
      RECT 9.904 13.986 10.008 18.36 ; 
      RECT 9.472 13.986 9.576 18.36 ; 
      RECT 9.04 13.986 9.144 18.36 ; 
      RECT 8.608 13.986 8.712 18.36 ; 
      RECT 8.176 13.986 8.28 18.36 ; 
      RECT 7.744 13.986 7.848 18.36 ; 
      RECT 7.312 13.986 7.416 18.36 ; 
      RECT 6.88 13.986 6.984 18.36 ; 
      RECT 6.448 13.986 6.552 18.36 ; 
      RECT 6.016 13.986 6.12 18.36 ; 
      RECT 5.584 13.986 5.688 18.36 ; 
      RECT 5.152 13.986 5.256 18.36 ; 
      RECT 4.72 13.986 4.824 18.36 ; 
      RECT 4.288 13.986 4.392 18.36 ; 
      RECT 3.856 13.986 3.96 18.36 ; 
      RECT 3.424 13.986 3.528 18.36 ; 
      RECT 2.992 13.986 3.096 18.36 ; 
      RECT 2.56 13.986 2.664 18.36 ; 
      RECT 2.128 13.986 2.232 18.36 ; 
      RECT 1.696 13.986 1.8 18.36 ; 
      RECT 1.264 13.986 1.368 18.36 ; 
      RECT 0.832 13.986 0.936 18.36 ; 
      RECT 0.02 13.986 0.36 18.36 ; 
      RECT 62.212 18.306 62.724 22.68 ; 
      RECT 62.156 20.968 62.724 22.258 ; 
      RECT 61.276 19.876 61.812 22.68 ; 
      RECT 61.184 21.216 61.812 22.248 ; 
      RECT 61.276 18.306 61.668 22.68 ; 
      RECT 61.276 18.79 61.724 19.748 ; 
      RECT 61.276 18.306 61.812 18.662 ; 
      RECT 60.376 20.108 60.912 22.68 ; 
      RECT 60.376 18.306 60.768 22.68 ; 
      RECT 58.708 18.306 59.04 22.68 ; 
      RECT 58.708 18.66 59.096 22.402 ; 
      RECT 121.072 18.306 121.412 22.68 ; 
      RECT 120.496 18.306 120.6 22.68 ; 
      RECT 120.064 18.306 120.168 22.68 ; 
      RECT 119.632 18.306 119.736 22.68 ; 
      RECT 119.2 18.306 119.304 22.68 ; 
      RECT 118.768 18.306 118.872 22.68 ; 
      RECT 118.336 18.306 118.44 22.68 ; 
      RECT 117.904 18.306 118.008 22.68 ; 
      RECT 117.472 18.306 117.576 22.68 ; 
      RECT 117.04 18.306 117.144 22.68 ; 
      RECT 116.608 18.306 116.712 22.68 ; 
      RECT 116.176 18.306 116.28 22.68 ; 
      RECT 115.744 18.306 115.848 22.68 ; 
      RECT 115.312 18.306 115.416 22.68 ; 
      RECT 114.88 18.306 114.984 22.68 ; 
      RECT 114.448 18.306 114.552 22.68 ; 
      RECT 114.016 18.306 114.12 22.68 ; 
      RECT 113.584 18.306 113.688 22.68 ; 
      RECT 113.152 18.306 113.256 22.68 ; 
      RECT 112.72 18.306 112.824 22.68 ; 
      RECT 112.288 18.306 112.392 22.68 ; 
      RECT 111.856 18.306 111.96 22.68 ; 
      RECT 111.424 18.306 111.528 22.68 ; 
      RECT 110.992 18.306 111.096 22.68 ; 
      RECT 110.56 18.306 110.664 22.68 ; 
      RECT 110.128 18.306 110.232 22.68 ; 
      RECT 109.696 18.306 109.8 22.68 ; 
      RECT 109.264 18.306 109.368 22.68 ; 
      RECT 108.832 18.306 108.936 22.68 ; 
      RECT 108.4 18.306 108.504 22.68 ; 
      RECT 107.968 18.306 108.072 22.68 ; 
      RECT 107.536 18.306 107.64 22.68 ; 
      RECT 107.104 18.306 107.208 22.68 ; 
      RECT 106.672 18.306 106.776 22.68 ; 
      RECT 106.24 18.306 106.344 22.68 ; 
      RECT 105.808 18.306 105.912 22.68 ; 
      RECT 105.376 18.306 105.48 22.68 ; 
      RECT 104.944 18.306 105.048 22.68 ; 
      RECT 104.512 18.306 104.616 22.68 ; 
      RECT 104.08 18.306 104.184 22.68 ; 
      RECT 103.648 18.306 103.752 22.68 ; 
      RECT 103.216 18.306 103.32 22.68 ; 
      RECT 102.784 18.306 102.888 22.68 ; 
      RECT 102.352 18.306 102.456 22.68 ; 
      RECT 101.92 18.306 102.024 22.68 ; 
      RECT 101.488 18.306 101.592 22.68 ; 
      RECT 101.056 18.306 101.16 22.68 ; 
      RECT 100.624 18.306 100.728 22.68 ; 
      RECT 100.192 18.306 100.296 22.68 ; 
      RECT 99.76 18.306 99.864 22.68 ; 
      RECT 99.328 18.306 99.432 22.68 ; 
      RECT 98.896 18.306 99 22.68 ; 
      RECT 98.464 18.306 98.568 22.68 ; 
      RECT 98.032 18.306 98.136 22.68 ; 
      RECT 97.6 18.306 97.704 22.68 ; 
      RECT 97.168 18.306 97.272 22.68 ; 
      RECT 96.736 18.306 96.84 22.68 ; 
      RECT 96.304 18.306 96.408 22.68 ; 
      RECT 95.872 18.306 95.976 22.68 ; 
      RECT 95.44 18.306 95.544 22.68 ; 
      RECT 95.008 18.306 95.112 22.68 ; 
      RECT 94.576 18.306 94.68 22.68 ; 
      RECT 94.144 18.306 94.248 22.68 ; 
      RECT 93.712 18.306 93.816 22.68 ; 
      RECT 93.28 18.306 93.384 22.68 ; 
      RECT 92.848 18.306 92.952 22.68 ; 
      RECT 92.416 18.306 92.52 22.68 ; 
      RECT 91.984 18.306 92.088 22.68 ; 
      RECT 91.552 18.306 91.656 22.68 ; 
      RECT 91.12 18.306 91.224 22.68 ; 
      RECT 90.688 18.306 90.792 22.68 ; 
      RECT 90.256 18.306 90.36 22.68 ; 
      RECT 89.824 18.306 89.928 22.68 ; 
      RECT 89.392 18.306 89.496 22.68 ; 
      RECT 88.96 18.306 89.064 22.68 ; 
      RECT 88.528 18.306 88.632 22.68 ; 
      RECT 88.096 18.306 88.2 22.68 ; 
      RECT 87.664 18.306 87.768 22.68 ; 
      RECT 87.232 18.306 87.336 22.68 ; 
      RECT 86.8 18.306 86.904 22.68 ; 
      RECT 86.368 18.306 86.472 22.68 ; 
      RECT 85.936 18.306 86.04 22.68 ; 
      RECT 85.504 18.306 85.608 22.68 ; 
      RECT 85.072 18.306 85.176 22.68 ; 
      RECT 84.64 18.306 84.744 22.68 ; 
      RECT 84.208 18.306 84.312 22.68 ; 
      RECT 83.776 18.306 83.88 22.68 ; 
      RECT 83.344 18.306 83.448 22.68 ; 
      RECT 82.912 18.306 83.016 22.68 ; 
      RECT 82.48 18.306 82.584 22.68 ; 
      RECT 82.048 18.306 82.152 22.68 ; 
      RECT 81.616 18.306 81.72 22.68 ; 
      RECT 81.184 18.306 81.288 22.68 ; 
      RECT 80.752 18.306 80.856 22.68 ; 
      RECT 80.32 18.306 80.424 22.68 ; 
      RECT 79.888 18.306 79.992 22.68 ; 
      RECT 79.456 18.306 79.56 22.68 ; 
      RECT 79.024 18.306 79.128 22.68 ; 
      RECT 78.592 18.306 78.696 22.68 ; 
      RECT 78.16 18.306 78.264 22.68 ; 
      RECT 77.728 18.306 77.832 22.68 ; 
      RECT 77.296 18.306 77.4 22.68 ; 
      RECT 76.864 18.306 76.968 22.68 ; 
      RECT 76.432 18.306 76.536 22.68 ; 
      RECT 76 18.306 76.104 22.68 ; 
      RECT 75.568 18.306 75.672 22.68 ; 
      RECT 75.136 18.306 75.24 22.68 ; 
      RECT 74.704 18.306 74.808 22.68 ; 
      RECT 74.272 18.306 74.376 22.68 ; 
      RECT 73.84 18.306 73.944 22.68 ; 
      RECT 73.408 18.306 73.512 22.68 ; 
      RECT 72.976 18.306 73.08 22.68 ; 
      RECT 72.544 18.306 72.648 22.68 ; 
      RECT 72.112 18.306 72.216 22.68 ; 
      RECT 71.68 18.306 71.784 22.68 ; 
      RECT 71.248 18.306 71.352 22.68 ; 
      RECT 70.816 18.306 70.92 22.68 ; 
      RECT 70.384 18.306 70.488 22.68 ; 
      RECT 69.952 18.306 70.056 22.68 ; 
      RECT 69.52 18.306 69.624 22.68 ; 
      RECT 69.088 18.306 69.192 22.68 ; 
      RECT 68.656 18.306 68.76 22.68 ; 
      RECT 68.224 18.306 68.328 22.68 ; 
      RECT 67.792 18.306 67.896 22.68 ; 
      RECT 67.36 18.306 67.464 22.68 ; 
      RECT 66.928 18.306 67.032 22.68 ; 
      RECT 66.496 18.306 66.6 22.68 ; 
      RECT 66.064 18.306 66.168 22.68 ; 
      RECT 65.632 18.306 65.736 22.68 ; 
      RECT 65.2 18.306 65.304 22.68 ; 
      RECT 64.348 18.306 64.656 22.68 ; 
      RECT 56.776 18.306 57.084 22.68 ; 
      RECT 56.128 18.306 56.232 22.68 ; 
      RECT 55.696 18.306 55.8 22.68 ; 
      RECT 55.264 18.306 55.368 22.68 ; 
      RECT 54.832 18.306 54.936 22.68 ; 
      RECT 54.4 18.306 54.504 22.68 ; 
      RECT 53.968 18.306 54.072 22.68 ; 
      RECT 53.536 18.306 53.64 22.68 ; 
      RECT 53.104 18.306 53.208 22.68 ; 
      RECT 52.672 18.306 52.776 22.68 ; 
      RECT 52.24 18.306 52.344 22.68 ; 
      RECT 51.808 18.306 51.912 22.68 ; 
      RECT 51.376 18.306 51.48 22.68 ; 
      RECT 50.944 18.306 51.048 22.68 ; 
      RECT 50.512 18.306 50.616 22.68 ; 
      RECT 50.08 18.306 50.184 22.68 ; 
      RECT 49.648 18.306 49.752 22.68 ; 
      RECT 49.216 18.306 49.32 22.68 ; 
      RECT 48.784 18.306 48.888 22.68 ; 
      RECT 48.352 18.306 48.456 22.68 ; 
      RECT 47.92 18.306 48.024 22.68 ; 
      RECT 47.488 18.306 47.592 22.68 ; 
      RECT 47.056 18.306 47.16 22.68 ; 
      RECT 46.624 18.306 46.728 22.68 ; 
      RECT 46.192 18.306 46.296 22.68 ; 
      RECT 45.76 18.306 45.864 22.68 ; 
      RECT 45.328 18.306 45.432 22.68 ; 
      RECT 44.896 18.306 45 22.68 ; 
      RECT 44.464 18.306 44.568 22.68 ; 
      RECT 44.032 18.306 44.136 22.68 ; 
      RECT 43.6 18.306 43.704 22.68 ; 
      RECT 43.168 18.306 43.272 22.68 ; 
      RECT 42.736 18.306 42.84 22.68 ; 
      RECT 42.304 18.306 42.408 22.68 ; 
      RECT 41.872 18.306 41.976 22.68 ; 
      RECT 41.44 18.306 41.544 22.68 ; 
      RECT 41.008 18.306 41.112 22.68 ; 
      RECT 40.576 18.306 40.68 22.68 ; 
      RECT 40.144 18.306 40.248 22.68 ; 
      RECT 39.712 18.306 39.816 22.68 ; 
      RECT 39.28 18.306 39.384 22.68 ; 
      RECT 38.848 18.306 38.952 22.68 ; 
      RECT 38.416 18.306 38.52 22.68 ; 
      RECT 37.984 18.306 38.088 22.68 ; 
      RECT 37.552 18.306 37.656 22.68 ; 
      RECT 37.12 18.306 37.224 22.68 ; 
      RECT 36.688 18.306 36.792 22.68 ; 
      RECT 36.256 18.306 36.36 22.68 ; 
      RECT 35.824 18.306 35.928 22.68 ; 
      RECT 35.392 18.306 35.496 22.68 ; 
      RECT 34.96 18.306 35.064 22.68 ; 
      RECT 34.528 18.306 34.632 22.68 ; 
      RECT 34.096 18.306 34.2 22.68 ; 
      RECT 33.664 18.306 33.768 22.68 ; 
      RECT 33.232 18.306 33.336 22.68 ; 
      RECT 32.8 18.306 32.904 22.68 ; 
      RECT 32.368 18.306 32.472 22.68 ; 
      RECT 31.936 18.306 32.04 22.68 ; 
      RECT 31.504 18.306 31.608 22.68 ; 
      RECT 31.072 18.306 31.176 22.68 ; 
      RECT 30.64 18.306 30.744 22.68 ; 
      RECT 30.208 18.306 30.312 22.68 ; 
      RECT 29.776 18.306 29.88 22.68 ; 
      RECT 29.344 18.306 29.448 22.68 ; 
      RECT 28.912 18.306 29.016 22.68 ; 
      RECT 28.48 18.306 28.584 22.68 ; 
      RECT 28.048 18.306 28.152 22.68 ; 
      RECT 27.616 18.306 27.72 22.68 ; 
      RECT 27.184 18.306 27.288 22.68 ; 
      RECT 26.752 18.306 26.856 22.68 ; 
      RECT 26.32 18.306 26.424 22.68 ; 
      RECT 25.888 18.306 25.992 22.68 ; 
      RECT 25.456 18.306 25.56 22.68 ; 
      RECT 25.024 18.306 25.128 22.68 ; 
      RECT 24.592 18.306 24.696 22.68 ; 
      RECT 24.16 18.306 24.264 22.68 ; 
      RECT 23.728 18.306 23.832 22.68 ; 
      RECT 23.296 18.306 23.4 22.68 ; 
      RECT 22.864 18.306 22.968 22.68 ; 
      RECT 22.432 18.306 22.536 22.68 ; 
      RECT 22 18.306 22.104 22.68 ; 
      RECT 21.568 18.306 21.672 22.68 ; 
      RECT 21.136 18.306 21.24 22.68 ; 
      RECT 20.704 18.306 20.808 22.68 ; 
      RECT 20.272 18.306 20.376 22.68 ; 
      RECT 19.84 18.306 19.944 22.68 ; 
      RECT 19.408 18.306 19.512 22.68 ; 
      RECT 18.976 18.306 19.08 22.68 ; 
      RECT 18.544 18.306 18.648 22.68 ; 
      RECT 18.112 18.306 18.216 22.68 ; 
      RECT 17.68 18.306 17.784 22.68 ; 
      RECT 17.248 18.306 17.352 22.68 ; 
      RECT 16.816 18.306 16.92 22.68 ; 
      RECT 16.384 18.306 16.488 22.68 ; 
      RECT 15.952 18.306 16.056 22.68 ; 
      RECT 15.52 18.306 15.624 22.68 ; 
      RECT 15.088 18.306 15.192 22.68 ; 
      RECT 14.656 18.306 14.76 22.68 ; 
      RECT 14.224 18.306 14.328 22.68 ; 
      RECT 13.792 18.306 13.896 22.68 ; 
      RECT 13.36 18.306 13.464 22.68 ; 
      RECT 12.928 18.306 13.032 22.68 ; 
      RECT 12.496 18.306 12.6 22.68 ; 
      RECT 12.064 18.306 12.168 22.68 ; 
      RECT 11.632 18.306 11.736 22.68 ; 
      RECT 11.2 18.306 11.304 22.68 ; 
      RECT 10.768 18.306 10.872 22.68 ; 
      RECT 10.336 18.306 10.44 22.68 ; 
      RECT 9.904 18.306 10.008 22.68 ; 
      RECT 9.472 18.306 9.576 22.68 ; 
      RECT 9.04 18.306 9.144 22.68 ; 
      RECT 8.608 18.306 8.712 22.68 ; 
      RECT 8.176 18.306 8.28 22.68 ; 
      RECT 7.744 18.306 7.848 22.68 ; 
      RECT 7.312 18.306 7.416 22.68 ; 
      RECT 6.88 18.306 6.984 22.68 ; 
      RECT 6.448 18.306 6.552 22.68 ; 
      RECT 6.016 18.306 6.12 22.68 ; 
      RECT 5.584 18.306 5.688 22.68 ; 
      RECT 5.152 18.306 5.256 22.68 ; 
      RECT 4.72 18.306 4.824 22.68 ; 
      RECT 4.288 18.306 4.392 22.68 ; 
      RECT 3.856 18.306 3.96 22.68 ; 
      RECT 3.424 18.306 3.528 22.68 ; 
      RECT 2.992 18.306 3.096 22.68 ; 
      RECT 2.56 18.306 2.664 22.68 ; 
      RECT 2.128 18.306 2.232 22.68 ; 
      RECT 1.696 18.306 1.8 22.68 ; 
      RECT 1.264 18.306 1.368 22.68 ; 
      RECT 0.832 18.306 0.936 22.68 ; 
      RECT 0.02 18.306 0.36 22.68 ; 
      RECT 62.212 22.626 62.724 27 ; 
      RECT 62.156 25.288 62.724 26.578 ; 
      RECT 61.276 24.196 61.812 27 ; 
      RECT 61.184 25.536 61.812 26.568 ; 
      RECT 61.276 22.626 61.668 27 ; 
      RECT 61.276 23.11 61.724 24.068 ; 
      RECT 61.276 22.626 61.812 22.982 ; 
      RECT 60.376 24.428 60.912 27 ; 
      RECT 60.376 22.626 60.768 27 ; 
      RECT 58.708 22.626 59.04 27 ; 
      RECT 58.708 22.98 59.096 26.722 ; 
      RECT 121.072 22.626 121.412 27 ; 
      RECT 120.496 22.626 120.6 27 ; 
      RECT 120.064 22.626 120.168 27 ; 
      RECT 119.632 22.626 119.736 27 ; 
      RECT 119.2 22.626 119.304 27 ; 
      RECT 118.768 22.626 118.872 27 ; 
      RECT 118.336 22.626 118.44 27 ; 
      RECT 117.904 22.626 118.008 27 ; 
      RECT 117.472 22.626 117.576 27 ; 
      RECT 117.04 22.626 117.144 27 ; 
      RECT 116.608 22.626 116.712 27 ; 
      RECT 116.176 22.626 116.28 27 ; 
      RECT 115.744 22.626 115.848 27 ; 
      RECT 115.312 22.626 115.416 27 ; 
      RECT 114.88 22.626 114.984 27 ; 
      RECT 114.448 22.626 114.552 27 ; 
      RECT 114.016 22.626 114.12 27 ; 
      RECT 113.584 22.626 113.688 27 ; 
      RECT 113.152 22.626 113.256 27 ; 
      RECT 112.72 22.626 112.824 27 ; 
      RECT 112.288 22.626 112.392 27 ; 
      RECT 111.856 22.626 111.96 27 ; 
      RECT 111.424 22.626 111.528 27 ; 
      RECT 110.992 22.626 111.096 27 ; 
      RECT 110.56 22.626 110.664 27 ; 
      RECT 110.128 22.626 110.232 27 ; 
      RECT 109.696 22.626 109.8 27 ; 
      RECT 109.264 22.626 109.368 27 ; 
      RECT 108.832 22.626 108.936 27 ; 
      RECT 108.4 22.626 108.504 27 ; 
      RECT 107.968 22.626 108.072 27 ; 
      RECT 107.536 22.626 107.64 27 ; 
      RECT 107.104 22.626 107.208 27 ; 
      RECT 106.672 22.626 106.776 27 ; 
      RECT 106.24 22.626 106.344 27 ; 
      RECT 105.808 22.626 105.912 27 ; 
      RECT 105.376 22.626 105.48 27 ; 
      RECT 104.944 22.626 105.048 27 ; 
      RECT 104.512 22.626 104.616 27 ; 
      RECT 104.08 22.626 104.184 27 ; 
      RECT 103.648 22.626 103.752 27 ; 
      RECT 103.216 22.626 103.32 27 ; 
      RECT 102.784 22.626 102.888 27 ; 
      RECT 102.352 22.626 102.456 27 ; 
      RECT 101.92 22.626 102.024 27 ; 
      RECT 101.488 22.626 101.592 27 ; 
      RECT 101.056 22.626 101.16 27 ; 
      RECT 100.624 22.626 100.728 27 ; 
      RECT 100.192 22.626 100.296 27 ; 
      RECT 99.76 22.626 99.864 27 ; 
      RECT 99.328 22.626 99.432 27 ; 
      RECT 98.896 22.626 99 27 ; 
      RECT 98.464 22.626 98.568 27 ; 
      RECT 98.032 22.626 98.136 27 ; 
      RECT 97.6 22.626 97.704 27 ; 
      RECT 97.168 22.626 97.272 27 ; 
      RECT 96.736 22.626 96.84 27 ; 
      RECT 96.304 22.626 96.408 27 ; 
      RECT 95.872 22.626 95.976 27 ; 
      RECT 95.44 22.626 95.544 27 ; 
      RECT 95.008 22.626 95.112 27 ; 
      RECT 94.576 22.626 94.68 27 ; 
      RECT 94.144 22.626 94.248 27 ; 
      RECT 93.712 22.626 93.816 27 ; 
      RECT 93.28 22.626 93.384 27 ; 
      RECT 92.848 22.626 92.952 27 ; 
      RECT 92.416 22.626 92.52 27 ; 
      RECT 91.984 22.626 92.088 27 ; 
      RECT 91.552 22.626 91.656 27 ; 
      RECT 91.12 22.626 91.224 27 ; 
      RECT 90.688 22.626 90.792 27 ; 
      RECT 90.256 22.626 90.36 27 ; 
      RECT 89.824 22.626 89.928 27 ; 
      RECT 89.392 22.626 89.496 27 ; 
      RECT 88.96 22.626 89.064 27 ; 
      RECT 88.528 22.626 88.632 27 ; 
      RECT 88.096 22.626 88.2 27 ; 
      RECT 87.664 22.626 87.768 27 ; 
      RECT 87.232 22.626 87.336 27 ; 
      RECT 86.8 22.626 86.904 27 ; 
      RECT 86.368 22.626 86.472 27 ; 
      RECT 85.936 22.626 86.04 27 ; 
      RECT 85.504 22.626 85.608 27 ; 
      RECT 85.072 22.626 85.176 27 ; 
      RECT 84.64 22.626 84.744 27 ; 
      RECT 84.208 22.626 84.312 27 ; 
      RECT 83.776 22.626 83.88 27 ; 
      RECT 83.344 22.626 83.448 27 ; 
      RECT 82.912 22.626 83.016 27 ; 
      RECT 82.48 22.626 82.584 27 ; 
      RECT 82.048 22.626 82.152 27 ; 
      RECT 81.616 22.626 81.72 27 ; 
      RECT 81.184 22.626 81.288 27 ; 
      RECT 80.752 22.626 80.856 27 ; 
      RECT 80.32 22.626 80.424 27 ; 
      RECT 79.888 22.626 79.992 27 ; 
      RECT 79.456 22.626 79.56 27 ; 
      RECT 79.024 22.626 79.128 27 ; 
      RECT 78.592 22.626 78.696 27 ; 
      RECT 78.16 22.626 78.264 27 ; 
      RECT 77.728 22.626 77.832 27 ; 
      RECT 77.296 22.626 77.4 27 ; 
      RECT 76.864 22.626 76.968 27 ; 
      RECT 76.432 22.626 76.536 27 ; 
      RECT 76 22.626 76.104 27 ; 
      RECT 75.568 22.626 75.672 27 ; 
      RECT 75.136 22.626 75.24 27 ; 
      RECT 74.704 22.626 74.808 27 ; 
      RECT 74.272 22.626 74.376 27 ; 
      RECT 73.84 22.626 73.944 27 ; 
      RECT 73.408 22.626 73.512 27 ; 
      RECT 72.976 22.626 73.08 27 ; 
      RECT 72.544 22.626 72.648 27 ; 
      RECT 72.112 22.626 72.216 27 ; 
      RECT 71.68 22.626 71.784 27 ; 
      RECT 71.248 22.626 71.352 27 ; 
      RECT 70.816 22.626 70.92 27 ; 
      RECT 70.384 22.626 70.488 27 ; 
      RECT 69.952 22.626 70.056 27 ; 
      RECT 69.52 22.626 69.624 27 ; 
      RECT 69.088 22.626 69.192 27 ; 
      RECT 68.656 22.626 68.76 27 ; 
      RECT 68.224 22.626 68.328 27 ; 
      RECT 67.792 22.626 67.896 27 ; 
      RECT 67.36 22.626 67.464 27 ; 
      RECT 66.928 22.626 67.032 27 ; 
      RECT 66.496 22.626 66.6 27 ; 
      RECT 66.064 22.626 66.168 27 ; 
      RECT 65.632 22.626 65.736 27 ; 
      RECT 65.2 22.626 65.304 27 ; 
      RECT 64.348 22.626 64.656 27 ; 
      RECT 56.776 22.626 57.084 27 ; 
      RECT 56.128 22.626 56.232 27 ; 
      RECT 55.696 22.626 55.8 27 ; 
      RECT 55.264 22.626 55.368 27 ; 
      RECT 54.832 22.626 54.936 27 ; 
      RECT 54.4 22.626 54.504 27 ; 
      RECT 53.968 22.626 54.072 27 ; 
      RECT 53.536 22.626 53.64 27 ; 
      RECT 53.104 22.626 53.208 27 ; 
      RECT 52.672 22.626 52.776 27 ; 
      RECT 52.24 22.626 52.344 27 ; 
      RECT 51.808 22.626 51.912 27 ; 
      RECT 51.376 22.626 51.48 27 ; 
      RECT 50.944 22.626 51.048 27 ; 
      RECT 50.512 22.626 50.616 27 ; 
      RECT 50.08 22.626 50.184 27 ; 
      RECT 49.648 22.626 49.752 27 ; 
      RECT 49.216 22.626 49.32 27 ; 
      RECT 48.784 22.626 48.888 27 ; 
      RECT 48.352 22.626 48.456 27 ; 
      RECT 47.92 22.626 48.024 27 ; 
      RECT 47.488 22.626 47.592 27 ; 
      RECT 47.056 22.626 47.16 27 ; 
      RECT 46.624 22.626 46.728 27 ; 
      RECT 46.192 22.626 46.296 27 ; 
      RECT 45.76 22.626 45.864 27 ; 
      RECT 45.328 22.626 45.432 27 ; 
      RECT 44.896 22.626 45 27 ; 
      RECT 44.464 22.626 44.568 27 ; 
      RECT 44.032 22.626 44.136 27 ; 
      RECT 43.6 22.626 43.704 27 ; 
      RECT 43.168 22.626 43.272 27 ; 
      RECT 42.736 22.626 42.84 27 ; 
      RECT 42.304 22.626 42.408 27 ; 
      RECT 41.872 22.626 41.976 27 ; 
      RECT 41.44 22.626 41.544 27 ; 
      RECT 41.008 22.626 41.112 27 ; 
      RECT 40.576 22.626 40.68 27 ; 
      RECT 40.144 22.626 40.248 27 ; 
      RECT 39.712 22.626 39.816 27 ; 
      RECT 39.28 22.626 39.384 27 ; 
      RECT 38.848 22.626 38.952 27 ; 
      RECT 38.416 22.626 38.52 27 ; 
      RECT 37.984 22.626 38.088 27 ; 
      RECT 37.552 22.626 37.656 27 ; 
      RECT 37.12 22.626 37.224 27 ; 
      RECT 36.688 22.626 36.792 27 ; 
      RECT 36.256 22.626 36.36 27 ; 
      RECT 35.824 22.626 35.928 27 ; 
      RECT 35.392 22.626 35.496 27 ; 
      RECT 34.96 22.626 35.064 27 ; 
      RECT 34.528 22.626 34.632 27 ; 
      RECT 34.096 22.626 34.2 27 ; 
      RECT 33.664 22.626 33.768 27 ; 
      RECT 33.232 22.626 33.336 27 ; 
      RECT 32.8 22.626 32.904 27 ; 
      RECT 32.368 22.626 32.472 27 ; 
      RECT 31.936 22.626 32.04 27 ; 
      RECT 31.504 22.626 31.608 27 ; 
      RECT 31.072 22.626 31.176 27 ; 
      RECT 30.64 22.626 30.744 27 ; 
      RECT 30.208 22.626 30.312 27 ; 
      RECT 29.776 22.626 29.88 27 ; 
      RECT 29.344 22.626 29.448 27 ; 
      RECT 28.912 22.626 29.016 27 ; 
      RECT 28.48 22.626 28.584 27 ; 
      RECT 28.048 22.626 28.152 27 ; 
      RECT 27.616 22.626 27.72 27 ; 
      RECT 27.184 22.626 27.288 27 ; 
      RECT 26.752 22.626 26.856 27 ; 
      RECT 26.32 22.626 26.424 27 ; 
      RECT 25.888 22.626 25.992 27 ; 
      RECT 25.456 22.626 25.56 27 ; 
      RECT 25.024 22.626 25.128 27 ; 
      RECT 24.592 22.626 24.696 27 ; 
      RECT 24.16 22.626 24.264 27 ; 
      RECT 23.728 22.626 23.832 27 ; 
      RECT 23.296 22.626 23.4 27 ; 
      RECT 22.864 22.626 22.968 27 ; 
      RECT 22.432 22.626 22.536 27 ; 
      RECT 22 22.626 22.104 27 ; 
      RECT 21.568 22.626 21.672 27 ; 
      RECT 21.136 22.626 21.24 27 ; 
      RECT 20.704 22.626 20.808 27 ; 
      RECT 20.272 22.626 20.376 27 ; 
      RECT 19.84 22.626 19.944 27 ; 
      RECT 19.408 22.626 19.512 27 ; 
      RECT 18.976 22.626 19.08 27 ; 
      RECT 18.544 22.626 18.648 27 ; 
      RECT 18.112 22.626 18.216 27 ; 
      RECT 17.68 22.626 17.784 27 ; 
      RECT 17.248 22.626 17.352 27 ; 
      RECT 16.816 22.626 16.92 27 ; 
      RECT 16.384 22.626 16.488 27 ; 
      RECT 15.952 22.626 16.056 27 ; 
      RECT 15.52 22.626 15.624 27 ; 
      RECT 15.088 22.626 15.192 27 ; 
      RECT 14.656 22.626 14.76 27 ; 
      RECT 14.224 22.626 14.328 27 ; 
      RECT 13.792 22.626 13.896 27 ; 
      RECT 13.36 22.626 13.464 27 ; 
      RECT 12.928 22.626 13.032 27 ; 
      RECT 12.496 22.626 12.6 27 ; 
      RECT 12.064 22.626 12.168 27 ; 
      RECT 11.632 22.626 11.736 27 ; 
      RECT 11.2 22.626 11.304 27 ; 
      RECT 10.768 22.626 10.872 27 ; 
      RECT 10.336 22.626 10.44 27 ; 
      RECT 9.904 22.626 10.008 27 ; 
      RECT 9.472 22.626 9.576 27 ; 
      RECT 9.04 22.626 9.144 27 ; 
      RECT 8.608 22.626 8.712 27 ; 
      RECT 8.176 22.626 8.28 27 ; 
      RECT 7.744 22.626 7.848 27 ; 
      RECT 7.312 22.626 7.416 27 ; 
      RECT 6.88 22.626 6.984 27 ; 
      RECT 6.448 22.626 6.552 27 ; 
      RECT 6.016 22.626 6.12 27 ; 
      RECT 5.584 22.626 5.688 27 ; 
      RECT 5.152 22.626 5.256 27 ; 
      RECT 4.72 22.626 4.824 27 ; 
      RECT 4.288 22.626 4.392 27 ; 
      RECT 3.856 22.626 3.96 27 ; 
      RECT 3.424 22.626 3.528 27 ; 
      RECT 2.992 22.626 3.096 27 ; 
      RECT 2.56 22.626 2.664 27 ; 
      RECT 2.128 22.626 2.232 27 ; 
      RECT 1.696 22.626 1.8 27 ; 
      RECT 1.264 22.626 1.368 27 ; 
      RECT 0.832 22.626 0.936 27 ; 
      RECT 0.02 22.626 0.36 27 ; 
      RECT 62.212 26.946 62.724 31.32 ; 
      RECT 62.156 29.608 62.724 30.898 ; 
      RECT 61.276 28.516 61.812 31.32 ; 
      RECT 61.184 29.856 61.812 30.888 ; 
      RECT 61.276 26.946 61.668 31.32 ; 
      RECT 61.276 27.43 61.724 28.388 ; 
      RECT 61.276 26.946 61.812 27.302 ; 
      RECT 60.376 28.748 60.912 31.32 ; 
      RECT 60.376 26.946 60.768 31.32 ; 
      RECT 58.708 26.946 59.04 31.32 ; 
      RECT 58.708 27.3 59.096 31.042 ; 
      RECT 121.072 26.946 121.412 31.32 ; 
      RECT 120.496 26.946 120.6 31.32 ; 
      RECT 120.064 26.946 120.168 31.32 ; 
      RECT 119.632 26.946 119.736 31.32 ; 
      RECT 119.2 26.946 119.304 31.32 ; 
      RECT 118.768 26.946 118.872 31.32 ; 
      RECT 118.336 26.946 118.44 31.32 ; 
      RECT 117.904 26.946 118.008 31.32 ; 
      RECT 117.472 26.946 117.576 31.32 ; 
      RECT 117.04 26.946 117.144 31.32 ; 
      RECT 116.608 26.946 116.712 31.32 ; 
      RECT 116.176 26.946 116.28 31.32 ; 
      RECT 115.744 26.946 115.848 31.32 ; 
      RECT 115.312 26.946 115.416 31.32 ; 
      RECT 114.88 26.946 114.984 31.32 ; 
      RECT 114.448 26.946 114.552 31.32 ; 
      RECT 114.016 26.946 114.12 31.32 ; 
      RECT 113.584 26.946 113.688 31.32 ; 
      RECT 113.152 26.946 113.256 31.32 ; 
      RECT 112.72 26.946 112.824 31.32 ; 
      RECT 112.288 26.946 112.392 31.32 ; 
      RECT 111.856 26.946 111.96 31.32 ; 
      RECT 111.424 26.946 111.528 31.32 ; 
      RECT 110.992 26.946 111.096 31.32 ; 
      RECT 110.56 26.946 110.664 31.32 ; 
      RECT 110.128 26.946 110.232 31.32 ; 
      RECT 109.696 26.946 109.8 31.32 ; 
      RECT 109.264 26.946 109.368 31.32 ; 
      RECT 108.832 26.946 108.936 31.32 ; 
      RECT 108.4 26.946 108.504 31.32 ; 
      RECT 107.968 26.946 108.072 31.32 ; 
      RECT 107.536 26.946 107.64 31.32 ; 
      RECT 107.104 26.946 107.208 31.32 ; 
      RECT 106.672 26.946 106.776 31.32 ; 
      RECT 106.24 26.946 106.344 31.32 ; 
      RECT 105.808 26.946 105.912 31.32 ; 
      RECT 105.376 26.946 105.48 31.32 ; 
      RECT 104.944 26.946 105.048 31.32 ; 
      RECT 104.512 26.946 104.616 31.32 ; 
      RECT 104.08 26.946 104.184 31.32 ; 
      RECT 103.648 26.946 103.752 31.32 ; 
      RECT 103.216 26.946 103.32 31.32 ; 
      RECT 102.784 26.946 102.888 31.32 ; 
      RECT 102.352 26.946 102.456 31.32 ; 
      RECT 101.92 26.946 102.024 31.32 ; 
      RECT 101.488 26.946 101.592 31.32 ; 
      RECT 101.056 26.946 101.16 31.32 ; 
      RECT 100.624 26.946 100.728 31.32 ; 
      RECT 100.192 26.946 100.296 31.32 ; 
      RECT 99.76 26.946 99.864 31.32 ; 
      RECT 99.328 26.946 99.432 31.32 ; 
      RECT 98.896 26.946 99 31.32 ; 
      RECT 98.464 26.946 98.568 31.32 ; 
      RECT 98.032 26.946 98.136 31.32 ; 
      RECT 97.6 26.946 97.704 31.32 ; 
      RECT 97.168 26.946 97.272 31.32 ; 
      RECT 96.736 26.946 96.84 31.32 ; 
      RECT 96.304 26.946 96.408 31.32 ; 
      RECT 95.872 26.946 95.976 31.32 ; 
      RECT 95.44 26.946 95.544 31.32 ; 
      RECT 95.008 26.946 95.112 31.32 ; 
      RECT 94.576 26.946 94.68 31.32 ; 
      RECT 94.144 26.946 94.248 31.32 ; 
      RECT 93.712 26.946 93.816 31.32 ; 
      RECT 93.28 26.946 93.384 31.32 ; 
      RECT 92.848 26.946 92.952 31.32 ; 
      RECT 92.416 26.946 92.52 31.32 ; 
      RECT 91.984 26.946 92.088 31.32 ; 
      RECT 91.552 26.946 91.656 31.32 ; 
      RECT 91.12 26.946 91.224 31.32 ; 
      RECT 90.688 26.946 90.792 31.32 ; 
      RECT 90.256 26.946 90.36 31.32 ; 
      RECT 89.824 26.946 89.928 31.32 ; 
      RECT 89.392 26.946 89.496 31.32 ; 
      RECT 88.96 26.946 89.064 31.32 ; 
      RECT 88.528 26.946 88.632 31.32 ; 
      RECT 88.096 26.946 88.2 31.32 ; 
      RECT 87.664 26.946 87.768 31.32 ; 
      RECT 87.232 26.946 87.336 31.32 ; 
      RECT 86.8 26.946 86.904 31.32 ; 
      RECT 86.368 26.946 86.472 31.32 ; 
      RECT 85.936 26.946 86.04 31.32 ; 
      RECT 85.504 26.946 85.608 31.32 ; 
      RECT 85.072 26.946 85.176 31.32 ; 
      RECT 84.64 26.946 84.744 31.32 ; 
      RECT 84.208 26.946 84.312 31.32 ; 
      RECT 83.776 26.946 83.88 31.32 ; 
      RECT 83.344 26.946 83.448 31.32 ; 
      RECT 82.912 26.946 83.016 31.32 ; 
      RECT 82.48 26.946 82.584 31.32 ; 
      RECT 82.048 26.946 82.152 31.32 ; 
      RECT 81.616 26.946 81.72 31.32 ; 
      RECT 81.184 26.946 81.288 31.32 ; 
      RECT 80.752 26.946 80.856 31.32 ; 
      RECT 80.32 26.946 80.424 31.32 ; 
      RECT 79.888 26.946 79.992 31.32 ; 
      RECT 79.456 26.946 79.56 31.32 ; 
      RECT 79.024 26.946 79.128 31.32 ; 
      RECT 78.592 26.946 78.696 31.32 ; 
      RECT 78.16 26.946 78.264 31.32 ; 
      RECT 77.728 26.946 77.832 31.32 ; 
      RECT 77.296 26.946 77.4 31.32 ; 
      RECT 76.864 26.946 76.968 31.32 ; 
      RECT 76.432 26.946 76.536 31.32 ; 
      RECT 76 26.946 76.104 31.32 ; 
      RECT 75.568 26.946 75.672 31.32 ; 
      RECT 75.136 26.946 75.24 31.32 ; 
      RECT 74.704 26.946 74.808 31.32 ; 
      RECT 74.272 26.946 74.376 31.32 ; 
      RECT 73.84 26.946 73.944 31.32 ; 
      RECT 73.408 26.946 73.512 31.32 ; 
      RECT 72.976 26.946 73.08 31.32 ; 
      RECT 72.544 26.946 72.648 31.32 ; 
      RECT 72.112 26.946 72.216 31.32 ; 
      RECT 71.68 26.946 71.784 31.32 ; 
      RECT 71.248 26.946 71.352 31.32 ; 
      RECT 70.816 26.946 70.92 31.32 ; 
      RECT 70.384 26.946 70.488 31.32 ; 
      RECT 69.952 26.946 70.056 31.32 ; 
      RECT 69.52 26.946 69.624 31.32 ; 
      RECT 69.088 26.946 69.192 31.32 ; 
      RECT 68.656 26.946 68.76 31.32 ; 
      RECT 68.224 26.946 68.328 31.32 ; 
      RECT 67.792 26.946 67.896 31.32 ; 
      RECT 67.36 26.946 67.464 31.32 ; 
      RECT 66.928 26.946 67.032 31.32 ; 
      RECT 66.496 26.946 66.6 31.32 ; 
      RECT 66.064 26.946 66.168 31.32 ; 
      RECT 65.632 26.946 65.736 31.32 ; 
      RECT 65.2 26.946 65.304 31.32 ; 
      RECT 64.348 26.946 64.656 31.32 ; 
      RECT 56.776 26.946 57.084 31.32 ; 
      RECT 56.128 26.946 56.232 31.32 ; 
      RECT 55.696 26.946 55.8 31.32 ; 
      RECT 55.264 26.946 55.368 31.32 ; 
      RECT 54.832 26.946 54.936 31.32 ; 
      RECT 54.4 26.946 54.504 31.32 ; 
      RECT 53.968 26.946 54.072 31.32 ; 
      RECT 53.536 26.946 53.64 31.32 ; 
      RECT 53.104 26.946 53.208 31.32 ; 
      RECT 52.672 26.946 52.776 31.32 ; 
      RECT 52.24 26.946 52.344 31.32 ; 
      RECT 51.808 26.946 51.912 31.32 ; 
      RECT 51.376 26.946 51.48 31.32 ; 
      RECT 50.944 26.946 51.048 31.32 ; 
      RECT 50.512 26.946 50.616 31.32 ; 
      RECT 50.08 26.946 50.184 31.32 ; 
      RECT 49.648 26.946 49.752 31.32 ; 
      RECT 49.216 26.946 49.32 31.32 ; 
      RECT 48.784 26.946 48.888 31.32 ; 
      RECT 48.352 26.946 48.456 31.32 ; 
      RECT 47.92 26.946 48.024 31.32 ; 
      RECT 47.488 26.946 47.592 31.32 ; 
      RECT 47.056 26.946 47.16 31.32 ; 
      RECT 46.624 26.946 46.728 31.32 ; 
      RECT 46.192 26.946 46.296 31.32 ; 
      RECT 45.76 26.946 45.864 31.32 ; 
      RECT 45.328 26.946 45.432 31.32 ; 
      RECT 44.896 26.946 45 31.32 ; 
      RECT 44.464 26.946 44.568 31.32 ; 
      RECT 44.032 26.946 44.136 31.32 ; 
      RECT 43.6 26.946 43.704 31.32 ; 
      RECT 43.168 26.946 43.272 31.32 ; 
      RECT 42.736 26.946 42.84 31.32 ; 
      RECT 42.304 26.946 42.408 31.32 ; 
      RECT 41.872 26.946 41.976 31.32 ; 
      RECT 41.44 26.946 41.544 31.32 ; 
      RECT 41.008 26.946 41.112 31.32 ; 
      RECT 40.576 26.946 40.68 31.32 ; 
      RECT 40.144 26.946 40.248 31.32 ; 
      RECT 39.712 26.946 39.816 31.32 ; 
      RECT 39.28 26.946 39.384 31.32 ; 
      RECT 38.848 26.946 38.952 31.32 ; 
      RECT 38.416 26.946 38.52 31.32 ; 
      RECT 37.984 26.946 38.088 31.32 ; 
      RECT 37.552 26.946 37.656 31.32 ; 
      RECT 37.12 26.946 37.224 31.32 ; 
      RECT 36.688 26.946 36.792 31.32 ; 
      RECT 36.256 26.946 36.36 31.32 ; 
      RECT 35.824 26.946 35.928 31.32 ; 
      RECT 35.392 26.946 35.496 31.32 ; 
      RECT 34.96 26.946 35.064 31.32 ; 
      RECT 34.528 26.946 34.632 31.32 ; 
      RECT 34.096 26.946 34.2 31.32 ; 
      RECT 33.664 26.946 33.768 31.32 ; 
      RECT 33.232 26.946 33.336 31.32 ; 
      RECT 32.8 26.946 32.904 31.32 ; 
      RECT 32.368 26.946 32.472 31.32 ; 
      RECT 31.936 26.946 32.04 31.32 ; 
      RECT 31.504 26.946 31.608 31.32 ; 
      RECT 31.072 26.946 31.176 31.32 ; 
      RECT 30.64 26.946 30.744 31.32 ; 
      RECT 30.208 26.946 30.312 31.32 ; 
      RECT 29.776 26.946 29.88 31.32 ; 
      RECT 29.344 26.946 29.448 31.32 ; 
      RECT 28.912 26.946 29.016 31.32 ; 
      RECT 28.48 26.946 28.584 31.32 ; 
      RECT 28.048 26.946 28.152 31.32 ; 
      RECT 27.616 26.946 27.72 31.32 ; 
      RECT 27.184 26.946 27.288 31.32 ; 
      RECT 26.752 26.946 26.856 31.32 ; 
      RECT 26.32 26.946 26.424 31.32 ; 
      RECT 25.888 26.946 25.992 31.32 ; 
      RECT 25.456 26.946 25.56 31.32 ; 
      RECT 25.024 26.946 25.128 31.32 ; 
      RECT 24.592 26.946 24.696 31.32 ; 
      RECT 24.16 26.946 24.264 31.32 ; 
      RECT 23.728 26.946 23.832 31.32 ; 
      RECT 23.296 26.946 23.4 31.32 ; 
      RECT 22.864 26.946 22.968 31.32 ; 
      RECT 22.432 26.946 22.536 31.32 ; 
      RECT 22 26.946 22.104 31.32 ; 
      RECT 21.568 26.946 21.672 31.32 ; 
      RECT 21.136 26.946 21.24 31.32 ; 
      RECT 20.704 26.946 20.808 31.32 ; 
      RECT 20.272 26.946 20.376 31.32 ; 
      RECT 19.84 26.946 19.944 31.32 ; 
      RECT 19.408 26.946 19.512 31.32 ; 
      RECT 18.976 26.946 19.08 31.32 ; 
      RECT 18.544 26.946 18.648 31.32 ; 
      RECT 18.112 26.946 18.216 31.32 ; 
      RECT 17.68 26.946 17.784 31.32 ; 
      RECT 17.248 26.946 17.352 31.32 ; 
      RECT 16.816 26.946 16.92 31.32 ; 
      RECT 16.384 26.946 16.488 31.32 ; 
      RECT 15.952 26.946 16.056 31.32 ; 
      RECT 15.52 26.946 15.624 31.32 ; 
      RECT 15.088 26.946 15.192 31.32 ; 
      RECT 14.656 26.946 14.76 31.32 ; 
      RECT 14.224 26.946 14.328 31.32 ; 
      RECT 13.792 26.946 13.896 31.32 ; 
      RECT 13.36 26.946 13.464 31.32 ; 
      RECT 12.928 26.946 13.032 31.32 ; 
      RECT 12.496 26.946 12.6 31.32 ; 
      RECT 12.064 26.946 12.168 31.32 ; 
      RECT 11.632 26.946 11.736 31.32 ; 
      RECT 11.2 26.946 11.304 31.32 ; 
      RECT 10.768 26.946 10.872 31.32 ; 
      RECT 10.336 26.946 10.44 31.32 ; 
      RECT 9.904 26.946 10.008 31.32 ; 
      RECT 9.472 26.946 9.576 31.32 ; 
      RECT 9.04 26.946 9.144 31.32 ; 
      RECT 8.608 26.946 8.712 31.32 ; 
      RECT 8.176 26.946 8.28 31.32 ; 
      RECT 7.744 26.946 7.848 31.32 ; 
      RECT 7.312 26.946 7.416 31.32 ; 
      RECT 6.88 26.946 6.984 31.32 ; 
      RECT 6.448 26.946 6.552 31.32 ; 
      RECT 6.016 26.946 6.12 31.32 ; 
      RECT 5.584 26.946 5.688 31.32 ; 
      RECT 5.152 26.946 5.256 31.32 ; 
      RECT 4.72 26.946 4.824 31.32 ; 
      RECT 4.288 26.946 4.392 31.32 ; 
      RECT 3.856 26.946 3.96 31.32 ; 
      RECT 3.424 26.946 3.528 31.32 ; 
      RECT 2.992 26.946 3.096 31.32 ; 
      RECT 2.56 26.946 2.664 31.32 ; 
      RECT 2.128 26.946 2.232 31.32 ; 
      RECT 1.696 26.946 1.8 31.32 ; 
      RECT 1.264 26.946 1.368 31.32 ; 
      RECT 0.832 26.946 0.936 31.32 ; 
      RECT 0.02 26.946 0.36 31.32 ; 
      RECT 62.212 31.266 62.724 35.64 ; 
      RECT 62.156 33.928 62.724 35.218 ; 
      RECT 61.276 32.836 61.812 35.64 ; 
      RECT 61.184 34.176 61.812 35.208 ; 
      RECT 61.276 31.266 61.668 35.64 ; 
      RECT 61.276 31.75 61.724 32.708 ; 
      RECT 61.276 31.266 61.812 31.622 ; 
      RECT 60.376 33.068 60.912 35.64 ; 
      RECT 60.376 31.266 60.768 35.64 ; 
      RECT 58.708 31.266 59.04 35.64 ; 
      RECT 58.708 31.62 59.096 35.362 ; 
      RECT 121.072 31.266 121.412 35.64 ; 
      RECT 120.496 31.266 120.6 35.64 ; 
      RECT 120.064 31.266 120.168 35.64 ; 
      RECT 119.632 31.266 119.736 35.64 ; 
      RECT 119.2 31.266 119.304 35.64 ; 
      RECT 118.768 31.266 118.872 35.64 ; 
      RECT 118.336 31.266 118.44 35.64 ; 
      RECT 117.904 31.266 118.008 35.64 ; 
      RECT 117.472 31.266 117.576 35.64 ; 
      RECT 117.04 31.266 117.144 35.64 ; 
      RECT 116.608 31.266 116.712 35.64 ; 
      RECT 116.176 31.266 116.28 35.64 ; 
      RECT 115.744 31.266 115.848 35.64 ; 
      RECT 115.312 31.266 115.416 35.64 ; 
      RECT 114.88 31.266 114.984 35.64 ; 
      RECT 114.448 31.266 114.552 35.64 ; 
      RECT 114.016 31.266 114.12 35.64 ; 
      RECT 113.584 31.266 113.688 35.64 ; 
      RECT 113.152 31.266 113.256 35.64 ; 
      RECT 112.72 31.266 112.824 35.64 ; 
      RECT 112.288 31.266 112.392 35.64 ; 
      RECT 111.856 31.266 111.96 35.64 ; 
      RECT 111.424 31.266 111.528 35.64 ; 
      RECT 110.992 31.266 111.096 35.64 ; 
      RECT 110.56 31.266 110.664 35.64 ; 
      RECT 110.128 31.266 110.232 35.64 ; 
      RECT 109.696 31.266 109.8 35.64 ; 
      RECT 109.264 31.266 109.368 35.64 ; 
      RECT 108.832 31.266 108.936 35.64 ; 
      RECT 108.4 31.266 108.504 35.64 ; 
      RECT 107.968 31.266 108.072 35.64 ; 
      RECT 107.536 31.266 107.64 35.64 ; 
      RECT 107.104 31.266 107.208 35.64 ; 
      RECT 106.672 31.266 106.776 35.64 ; 
      RECT 106.24 31.266 106.344 35.64 ; 
      RECT 105.808 31.266 105.912 35.64 ; 
      RECT 105.376 31.266 105.48 35.64 ; 
      RECT 104.944 31.266 105.048 35.64 ; 
      RECT 104.512 31.266 104.616 35.64 ; 
      RECT 104.08 31.266 104.184 35.64 ; 
      RECT 103.648 31.266 103.752 35.64 ; 
      RECT 103.216 31.266 103.32 35.64 ; 
      RECT 102.784 31.266 102.888 35.64 ; 
      RECT 102.352 31.266 102.456 35.64 ; 
      RECT 101.92 31.266 102.024 35.64 ; 
      RECT 101.488 31.266 101.592 35.64 ; 
      RECT 101.056 31.266 101.16 35.64 ; 
      RECT 100.624 31.266 100.728 35.64 ; 
      RECT 100.192 31.266 100.296 35.64 ; 
      RECT 99.76 31.266 99.864 35.64 ; 
      RECT 99.328 31.266 99.432 35.64 ; 
      RECT 98.896 31.266 99 35.64 ; 
      RECT 98.464 31.266 98.568 35.64 ; 
      RECT 98.032 31.266 98.136 35.64 ; 
      RECT 97.6 31.266 97.704 35.64 ; 
      RECT 97.168 31.266 97.272 35.64 ; 
      RECT 96.736 31.266 96.84 35.64 ; 
      RECT 96.304 31.266 96.408 35.64 ; 
      RECT 95.872 31.266 95.976 35.64 ; 
      RECT 95.44 31.266 95.544 35.64 ; 
      RECT 95.008 31.266 95.112 35.64 ; 
      RECT 94.576 31.266 94.68 35.64 ; 
      RECT 94.144 31.266 94.248 35.64 ; 
      RECT 93.712 31.266 93.816 35.64 ; 
      RECT 93.28 31.266 93.384 35.64 ; 
      RECT 92.848 31.266 92.952 35.64 ; 
      RECT 92.416 31.266 92.52 35.64 ; 
      RECT 91.984 31.266 92.088 35.64 ; 
      RECT 91.552 31.266 91.656 35.64 ; 
      RECT 91.12 31.266 91.224 35.64 ; 
      RECT 90.688 31.266 90.792 35.64 ; 
      RECT 90.256 31.266 90.36 35.64 ; 
      RECT 89.824 31.266 89.928 35.64 ; 
      RECT 89.392 31.266 89.496 35.64 ; 
      RECT 88.96 31.266 89.064 35.64 ; 
      RECT 88.528 31.266 88.632 35.64 ; 
      RECT 88.096 31.266 88.2 35.64 ; 
      RECT 87.664 31.266 87.768 35.64 ; 
      RECT 87.232 31.266 87.336 35.64 ; 
      RECT 86.8 31.266 86.904 35.64 ; 
      RECT 86.368 31.266 86.472 35.64 ; 
      RECT 85.936 31.266 86.04 35.64 ; 
      RECT 85.504 31.266 85.608 35.64 ; 
      RECT 85.072 31.266 85.176 35.64 ; 
      RECT 84.64 31.266 84.744 35.64 ; 
      RECT 84.208 31.266 84.312 35.64 ; 
      RECT 83.776 31.266 83.88 35.64 ; 
      RECT 83.344 31.266 83.448 35.64 ; 
      RECT 82.912 31.266 83.016 35.64 ; 
      RECT 82.48 31.266 82.584 35.64 ; 
      RECT 82.048 31.266 82.152 35.64 ; 
      RECT 81.616 31.266 81.72 35.64 ; 
      RECT 81.184 31.266 81.288 35.64 ; 
      RECT 80.752 31.266 80.856 35.64 ; 
      RECT 80.32 31.266 80.424 35.64 ; 
      RECT 79.888 31.266 79.992 35.64 ; 
      RECT 79.456 31.266 79.56 35.64 ; 
      RECT 79.024 31.266 79.128 35.64 ; 
      RECT 78.592 31.266 78.696 35.64 ; 
      RECT 78.16 31.266 78.264 35.64 ; 
      RECT 77.728 31.266 77.832 35.64 ; 
      RECT 77.296 31.266 77.4 35.64 ; 
      RECT 76.864 31.266 76.968 35.64 ; 
      RECT 76.432 31.266 76.536 35.64 ; 
      RECT 76 31.266 76.104 35.64 ; 
      RECT 75.568 31.266 75.672 35.64 ; 
      RECT 75.136 31.266 75.24 35.64 ; 
      RECT 74.704 31.266 74.808 35.64 ; 
      RECT 74.272 31.266 74.376 35.64 ; 
      RECT 73.84 31.266 73.944 35.64 ; 
      RECT 73.408 31.266 73.512 35.64 ; 
      RECT 72.976 31.266 73.08 35.64 ; 
      RECT 72.544 31.266 72.648 35.64 ; 
      RECT 72.112 31.266 72.216 35.64 ; 
      RECT 71.68 31.266 71.784 35.64 ; 
      RECT 71.248 31.266 71.352 35.64 ; 
      RECT 70.816 31.266 70.92 35.64 ; 
      RECT 70.384 31.266 70.488 35.64 ; 
      RECT 69.952 31.266 70.056 35.64 ; 
      RECT 69.52 31.266 69.624 35.64 ; 
      RECT 69.088 31.266 69.192 35.64 ; 
      RECT 68.656 31.266 68.76 35.64 ; 
      RECT 68.224 31.266 68.328 35.64 ; 
      RECT 67.792 31.266 67.896 35.64 ; 
      RECT 67.36 31.266 67.464 35.64 ; 
      RECT 66.928 31.266 67.032 35.64 ; 
      RECT 66.496 31.266 66.6 35.64 ; 
      RECT 66.064 31.266 66.168 35.64 ; 
      RECT 65.632 31.266 65.736 35.64 ; 
      RECT 65.2 31.266 65.304 35.64 ; 
      RECT 64.348 31.266 64.656 35.64 ; 
      RECT 56.776 31.266 57.084 35.64 ; 
      RECT 56.128 31.266 56.232 35.64 ; 
      RECT 55.696 31.266 55.8 35.64 ; 
      RECT 55.264 31.266 55.368 35.64 ; 
      RECT 54.832 31.266 54.936 35.64 ; 
      RECT 54.4 31.266 54.504 35.64 ; 
      RECT 53.968 31.266 54.072 35.64 ; 
      RECT 53.536 31.266 53.64 35.64 ; 
      RECT 53.104 31.266 53.208 35.64 ; 
      RECT 52.672 31.266 52.776 35.64 ; 
      RECT 52.24 31.266 52.344 35.64 ; 
      RECT 51.808 31.266 51.912 35.64 ; 
      RECT 51.376 31.266 51.48 35.64 ; 
      RECT 50.944 31.266 51.048 35.64 ; 
      RECT 50.512 31.266 50.616 35.64 ; 
      RECT 50.08 31.266 50.184 35.64 ; 
      RECT 49.648 31.266 49.752 35.64 ; 
      RECT 49.216 31.266 49.32 35.64 ; 
      RECT 48.784 31.266 48.888 35.64 ; 
      RECT 48.352 31.266 48.456 35.64 ; 
      RECT 47.92 31.266 48.024 35.64 ; 
      RECT 47.488 31.266 47.592 35.64 ; 
      RECT 47.056 31.266 47.16 35.64 ; 
      RECT 46.624 31.266 46.728 35.64 ; 
      RECT 46.192 31.266 46.296 35.64 ; 
      RECT 45.76 31.266 45.864 35.64 ; 
      RECT 45.328 31.266 45.432 35.64 ; 
      RECT 44.896 31.266 45 35.64 ; 
      RECT 44.464 31.266 44.568 35.64 ; 
      RECT 44.032 31.266 44.136 35.64 ; 
      RECT 43.6 31.266 43.704 35.64 ; 
      RECT 43.168 31.266 43.272 35.64 ; 
      RECT 42.736 31.266 42.84 35.64 ; 
      RECT 42.304 31.266 42.408 35.64 ; 
      RECT 41.872 31.266 41.976 35.64 ; 
      RECT 41.44 31.266 41.544 35.64 ; 
      RECT 41.008 31.266 41.112 35.64 ; 
      RECT 40.576 31.266 40.68 35.64 ; 
      RECT 40.144 31.266 40.248 35.64 ; 
      RECT 39.712 31.266 39.816 35.64 ; 
      RECT 39.28 31.266 39.384 35.64 ; 
      RECT 38.848 31.266 38.952 35.64 ; 
      RECT 38.416 31.266 38.52 35.64 ; 
      RECT 37.984 31.266 38.088 35.64 ; 
      RECT 37.552 31.266 37.656 35.64 ; 
      RECT 37.12 31.266 37.224 35.64 ; 
      RECT 36.688 31.266 36.792 35.64 ; 
      RECT 36.256 31.266 36.36 35.64 ; 
      RECT 35.824 31.266 35.928 35.64 ; 
      RECT 35.392 31.266 35.496 35.64 ; 
      RECT 34.96 31.266 35.064 35.64 ; 
      RECT 34.528 31.266 34.632 35.64 ; 
      RECT 34.096 31.266 34.2 35.64 ; 
      RECT 33.664 31.266 33.768 35.64 ; 
      RECT 33.232 31.266 33.336 35.64 ; 
      RECT 32.8 31.266 32.904 35.64 ; 
      RECT 32.368 31.266 32.472 35.64 ; 
      RECT 31.936 31.266 32.04 35.64 ; 
      RECT 31.504 31.266 31.608 35.64 ; 
      RECT 31.072 31.266 31.176 35.64 ; 
      RECT 30.64 31.266 30.744 35.64 ; 
      RECT 30.208 31.266 30.312 35.64 ; 
      RECT 29.776 31.266 29.88 35.64 ; 
      RECT 29.344 31.266 29.448 35.64 ; 
      RECT 28.912 31.266 29.016 35.64 ; 
      RECT 28.48 31.266 28.584 35.64 ; 
      RECT 28.048 31.266 28.152 35.64 ; 
      RECT 27.616 31.266 27.72 35.64 ; 
      RECT 27.184 31.266 27.288 35.64 ; 
      RECT 26.752 31.266 26.856 35.64 ; 
      RECT 26.32 31.266 26.424 35.64 ; 
      RECT 25.888 31.266 25.992 35.64 ; 
      RECT 25.456 31.266 25.56 35.64 ; 
      RECT 25.024 31.266 25.128 35.64 ; 
      RECT 24.592 31.266 24.696 35.64 ; 
      RECT 24.16 31.266 24.264 35.64 ; 
      RECT 23.728 31.266 23.832 35.64 ; 
      RECT 23.296 31.266 23.4 35.64 ; 
      RECT 22.864 31.266 22.968 35.64 ; 
      RECT 22.432 31.266 22.536 35.64 ; 
      RECT 22 31.266 22.104 35.64 ; 
      RECT 21.568 31.266 21.672 35.64 ; 
      RECT 21.136 31.266 21.24 35.64 ; 
      RECT 20.704 31.266 20.808 35.64 ; 
      RECT 20.272 31.266 20.376 35.64 ; 
      RECT 19.84 31.266 19.944 35.64 ; 
      RECT 19.408 31.266 19.512 35.64 ; 
      RECT 18.976 31.266 19.08 35.64 ; 
      RECT 18.544 31.266 18.648 35.64 ; 
      RECT 18.112 31.266 18.216 35.64 ; 
      RECT 17.68 31.266 17.784 35.64 ; 
      RECT 17.248 31.266 17.352 35.64 ; 
      RECT 16.816 31.266 16.92 35.64 ; 
      RECT 16.384 31.266 16.488 35.64 ; 
      RECT 15.952 31.266 16.056 35.64 ; 
      RECT 15.52 31.266 15.624 35.64 ; 
      RECT 15.088 31.266 15.192 35.64 ; 
      RECT 14.656 31.266 14.76 35.64 ; 
      RECT 14.224 31.266 14.328 35.64 ; 
      RECT 13.792 31.266 13.896 35.64 ; 
      RECT 13.36 31.266 13.464 35.64 ; 
      RECT 12.928 31.266 13.032 35.64 ; 
      RECT 12.496 31.266 12.6 35.64 ; 
      RECT 12.064 31.266 12.168 35.64 ; 
      RECT 11.632 31.266 11.736 35.64 ; 
      RECT 11.2 31.266 11.304 35.64 ; 
      RECT 10.768 31.266 10.872 35.64 ; 
      RECT 10.336 31.266 10.44 35.64 ; 
      RECT 9.904 31.266 10.008 35.64 ; 
      RECT 9.472 31.266 9.576 35.64 ; 
      RECT 9.04 31.266 9.144 35.64 ; 
      RECT 8.608 31.266 8.712 35.64 ; 
      RECT 8.176 31.266 8.28 35.64 ; 
      RECT 7.744 31.266 7.848 35.64 ; 
      RECT 7.312 31.266 7.416 35.64 ; 
      RECT 6.88 31.266 6.984 35.64 ; 
      RECT 6.448 31.266 6.552 35.64 ; 
      RECT 6.016 31.266 6.12 35.64 ; 
      RECT 5.584 31.266 5.688 35.64 ; 
      RECT 5.152 31.266 5.256 35.64 ; 
      RECT 4.72 31.266 4.824 35.64 ; 
      RECT 4.288 31.266 4.392 35.64 ; 
      RECT 3.856 31.266 3.96 35.64 ; 
      RECT 3.424 31.266 3.528 35.64 ; 
      RECT 2.992 31.266 3.096 35.64 ; 
      RECT 2.56 31.266 2.664 35.64 ; 
      RECT 2.128 31.266 2.232 35.64 ; 
      RECT 1.696 31.266 1.8 35.64 ; 
      RECT 1.264 31.266 1.368 35.64 ; 
      RECT 0.832 31.266 0.936 35.64 ; 
      RECT 0.02 31.266 0.36 35.64 ; 
      RECT 62.212 35.586 62.724 39.96 ; 
      RECT 62.156 38.248 62.724 39.538 ; 
      RECT 61.276 37.156 61.812 39.96 ; 
      RECT 61.184 38.496 61.812 39.528 ; 
      RECT 61.276 35.586 61.668 39.96 ; 
      RECT 61.276 36.07 61.724 37.028 ; 
      RECT 61.276 35.586 61.812 35.942 ; 
      RECT 60.376 37.388 60.912 39.96 ; 
      RECT 60.376 35.586 60.768 39.96 ; 
      RECT 58.708 35.586 59.04 39.96 ; 
      RECT 58.708 35.94 59.096 39.682 ; 
      RECT 121.072 35.586 121.412 39.96 ; 
      RECT 120.496 35.586 120.6 39.96 ; 
      RECT 120.064 35.586 120.168 39.96 ; 
      RECT 119.632 35.586 119.736 39.96 ; 
      RECT 119.2 35.586 119.304 39.96 ; 
      RECT 118.768 35.586 118.872 39.96 ; 
      RECT 118.336 35.586 118.44 39.96 ; 
      RECT 117.904 35.586 118.008 39.96 ; 
      RECT 117.472 35.586 117.576 39.96 ; 
      RECT 117.04 35.586 117.144 39.96 ; 
      RECT 116.608 35.586 116.712 39.96 ; 
      RECT 116.176 35.586 116.28 39.96 ; 
      RECT 115.744 35.586 115.848 39.96 ; 
      RECT 115.312 35.586 115.416 39.96 ; 
      RECT 114.88 35.586 114.984 39.96 ; 
      RECT 114.448 35.586 114.552 39.96 ; 
      RECT 114.016 35.586 114.12 39.96 ; 
      RECT 113.584 35.586 113.688 39.96 ; 
      RECT 113.152 35.586 113.256 39.96 ; 
      RECT 112.72 35.586 112.824 39.96 ; 
      RECT 112.288 35.586 112.392 39.96 ; 
      RECT 111.856 35.586 111.96 39.96 ; 
      RECT 111.424 35.586 111.528 39.96 ; 
      RECT 110.992 35.586 111.096 39.96 ; 
      RECT 110.56 35.586 110.664 39.96 ; 
      RECT 110.128 35.586 110.232 39.96 ; 
      RECT 109.696 35.586 109.8 39.96 ; 
      RECT 109.264 35.586 109.368 39.96 ; 
      RECT 108.832 35.586 108.936 39.96 ; 
      RECT 108.4 35.586 108.504 39.96 ; 
      RECT 107.968 35.586 108.072 39.96 ; 
      RECT 107.536 35.586 107.64 39.96 ; 
      RECT 107.104 35.586 107.208 39.96 ; 
      RECT 106.672 35.586 106.776 39.96 ; 
      RECT 106.24 35.586 106.344 39.96 ; 
      RECT 105.808 35.586 105.912 39.96 ; 
      RECT 105.376 35.586 105.48 39.96 ; 
      RECT 104.944 35.586 105.048 39.96 ; 
      RECT 104.512 35.586 104.616 39.96 ; 
      RECT 104.08 35.586 104.184 39.96 ; 
      RECT 103.648 35.586 103.752 39.96 ; 
      RECT 103.216 35.586 103.32 39.96 ; 
      RECT 102.784 35.586 102.888 39.96 ; 
      RECT 102.352 35.586 102.456 39.96 ; 
      RECT 101.92 35.586 102.024 39.96 ; 
      RECT 101.488 35.586 101.592 39.96 ; 
      RECT 101.056 35.586 101.16 39.96 ; 
      RECT 100.624 35.586 100.728 39.96 ; 
      RECT 100.192 35.586 100.296 39.96 ; 
      RECT 99.76 35.586 99.864 39.96 ; 
      RECT 99.328 35.586 99.432 39.96 ; 
      RECT 98.896 35.586 99 39.96 ; 
      RECT 98.464 35.586 98.568 39.96 ; 
      RECT 98.032 35.586 98.136 39.96 ; 
      RECT 97.6 35.586 97.704 39.96 ; 
      RECT 97.168 35.586 97.272 39.96 ; 
      RECT 96.736 35.586 96.84 39.96 ; 
      RECT 96.304 35.586 96.408 39.96 ; 
      RECT 95.872 35.586 95.976 39.96 ; 
      RECT 95.44 35.586 95.544 39.96 ; 
      RECT 95.008 35.586 95.112 39.96 ; 
      RECT 94.576 35.586 94.68 39.96 ; 
      RECT 94.144 35.586 94.248 39.96 ; 
      RECT 93.712 35.586 93.816 39.96 ; 
      RECT 93.28 35.586 93.384 39.96 ; 
      RECT 92.848 35.586 92.952 39.96 ; 
      RECT 92.416 35.586 92.52 39.96 ; 
      RECT 91.984 35.586 92.088 39.96 ; 
      RECT 91.552 35.586 91.656 39.96 ; 
      RECT 91.12 35.586 91.224 39.96 ; 
      RECT 90.688 35.586 90.792 39.96 ; 
      RECT 90.256 35.586 90.36 39.96 ; 
      RECT 89.824 35.586 89.928 39.96 ; 
      RECT 89.392 35.586 89.496 39.96 ; 
      RECT 88.96 35.586 89.064 39.96 ; 
      RECT 88.528 35.586 88.632 39.96 ; 
      RECT 88.096 35.586 88.2 39.96 ; 
      RECT 87.664 35.586 87.768 39.96 ; 
      RECT 87.232 35.586 87.336 39.96 ; 
      RECT 86.8 35.586 86.904 39.96 ; 
      RECT 86.368 35.586 86.472 39.96 ; 
      RECT 85.936 35.586 86.04 39.96 ; 
      RECT 85.504 35.586 85.608 39.96 ; 
      RECT 85.072 35.586 85.176 39.96 ; 
      RECT 84.64 35.586 84.744 39.96 ; 
      RECT 84.208 35.586 84.312 39.96 ; 
      RECT 83.776 35.586 83.88 39.96 ; 
      RECT 83.344 35.586 83.448 39.96 ; 
      RECT 82.912 35.586 83.016 39.96 ; 
      RECT 82.48 35.586 82.584 39.96 ; 
      RECT 82.048 35.586 82.152 39.96 ; 
      RECT 81.616 35.586 81.72 39.96 ; 
      RECT 81.184 35.586 81.288 39.96 ; 
      RECT 80.752 35.586 80.856 39.96 ; 
      RECT 80.32 35.586 80.424 39.96 ; 
      RECT 79.888 35.586 79.992 39.96 ; 
      RECT 79.456 35.586 79.56 39.96 ; 
      RECT 79.024 35.586 79.128 39.96 ; 
      RECT 78.592 35.586 78.696 39.96 ; 
      RECT 78.16 35.586 78.264 39.96 ; 
      RECT 77.728 35.586 77.832 39.96 ; 
      RECT 77.296 35.586 77.4 39.96 ; 
      RECT 76.864 35.586 76.968 39.96 ; 
      RECT 76.432 35.586 76.536 39.96 ; 
      RECT 76 35.586 76.104 39.96 ; 
      RECT 75.568 35.586 75.672 39.96 ; 
      RECT 75.136 35.586 75.24 39.96 ; 
      RECT 74.704 35.586 74.808 39.96 ; 
      RECT 74.272 35.586 74.376 39.96 ; 
      RECT 73.84 35.586 73.944 39.96 ; 
      RECT 73.408 35.586 73.512 39.96 ; 
      RECT 72.976 35.586 73.08 39.96 ; 
      RECT 72.544 35.586 72.648 39.96 ; 
      RECT 72.112 35.586 72.216 39.96 ; 
      RECT 71.68 35.586 71.784 39.96 ; 
      RECT 71.248 35.586 71.352 39.96 ; 
      RECT 70.816 35.586 70.92 39.96 ; 
      RECT 70.384 35.586 70.488 39.96 ; 
      RECT 69.952 35.586 70.056 39.96 ; 
      RECT 69.52 35.586 69.624 39.96 ; 
      RECT 69.088 35.586 69.192 39.96 ; 
      RECT 68.656 35.586 68.76 39.96 ; 
      RECT 68.224 35.586 68.328 39.96 ; 
      RECT 67.792 35.586 67.896 39.96 ; 
      RECT 67.36 35.586 67.464 39.96 ; 
      RECT 66.928 35.586 67.032 39.96 ; 
      RECT 66.496 35.586 66.6 39.96 ; 
      RECT 66.064 35.586 66.168 39.96 ; 
      RECT 65.632 35.586 65.736 39.96 ; 
      RECT 65.2 35.586 65.304 39.96 ; 
      RECT 64.348 35.586 64.656 39.96 ; 
      RECT 56.776 35.586 57.084 39.96 ; 
      RECT 56.128 35.586 56.232 39.96 ; 
      RECT 55.696 35.586 55.8 39.96 ; 
      RECT 55.264 35.586 55.368 39.96 ; 
      RECT 54.832 35.586 54.936 39.96 ; 
      RECT 54.4 35.586 54.504 39.96 ; 
      RECT 53.968 35.586 54.072 39.96 ; 
      RECT 53.536 35.586 53.64 39.96 ; 
      RECT 53.104 35.586 53.208 39.96 ; 
      RECT 52.672 35.586 52.776 39.96 ; 
      RECT 52.24 35.586 52.344 39.96 ; 
      RECT 51.808 35.586 51.912 39.96 ; 
      RECT 51.376 35.586 51.48 39.96 ; 
      RECT 50.944 35.586 51.048 39.96 ; 
      RECT 50.512 35.586 50.616 39.96 ; 
      RECT 50.08 35.586 50.184 39.96 ; 
      RECT 49.648 35.586 49.752 39.96 ; 
      RECT 49.216 35.586 49.32 39.96 ; 
      RECT 48.784 35.586 48.888 39.96 ; 
      RECT 48.352 35.586 48.456 39.96 ; 
      RECT 47.92 35.586 48.024 39.96 ; 
      RECT 47.488 35.586 47.592 39.96 ; 
      RECT 47.056 35.586 47.16 39.96 ; 
      RECT 46.624 35.586 46.728 39.96 ; 
      RECT 46.192 35.586 46.296 39.96 ; 
      RECT 45.76 35.586 45.864 39.96 ; 
      RECT 45.328 35.586 45.432 39.96 ; 
      RECT 44.896 35.586 45 39.96 ; 
      RECT 44.464 35.586 44.568 39.96 ; 
      RECT 44.032 35.586 44.136 39.96 ; 
      RECT 43.6 35.586 43.704 39.96 ; 
      RECT 43.168 35.586 43.272 39.96 ; 
      RECT 42.736 35.586 42.84 39.96 ; 
      RECT 42.304 35.586 42.408 39.96 ; 
      RECT 41.872 35.586 41.976 39.96 ; 
      RECT 41.44 35.586 41.544 39.96 ; 
      RECT 41.008 35.586 41.112 39.96 ; 
      RECT 40.576 35.586 40.68 39.96 ; 
      RECT 40.144 35.586 40.248 39.96 ; 
      RECT 39.712 35.586 39.816 39.96 ; 
      RECT 39.28 35.586 39.384 39.96 ; 
      RECT 38.848 35.586 38.952 39.96 ; 
      RECT 38.416 35.586 38.52 39.96 ; 
      RECT 37.984 35.586 38.088 39.96 ; 
      RECT 37.552 35.586 37.656 39.96 ; 
      RECT 37.12 35.586 37.224 39.96 ; 
      RECT 36.688 35.586 36.792 39.96 ; 
      RECT 36.256 35.586 36.36 39.96 ; 
      RECT 35.824 35.586 35.928 39.96 ; 
      RECT 35.392 35.586 35.496 39.96 ; 
      RECT 34.96 35.586 35.064 39.96 ; 
      RECT 34.528 35.586 34.632 39.96 ; 
      RECT 34.096 35.586 34.2 39.96 ; 
      RECT 33.664 35.586 33.768 39.96 ; 
      RECT 33.232 35.586 33.336 39.96 ; 
      RECT 32.8 35.586 32.904 39.96 ; 
      RECT 32.368 35.586 32.472 39.96 ; 
      RECT 31.936 35.586 32.04 39.96 ; 
      RECT 31.504 35.586 31.608 39.96 ; 
      RECT 31.072 35.586 31.176 39.96 ; 
      RECT 30.64 35.586 30.744 39.96 ; 
      RECT 30.208 35.586 30.312 39.96 ; 
      RECT 29.776 35.586 29.88 39.96 ; 
      RECT 29.344 35.586 29.448 39.96 ; 
      RECT 28.912 35.586 29.016 39.96 ; 
      RECT 28.48 35.586 28.584 39.96 ; 
      RECT 28.048 35.586 28.152 39.96 ; 
      RECT 27.616 35.586 27.72 39.96 ; 
      RECT 27.184 35.586 27.288 39.96 ; 
      RECT 26.752 35.586 26.856 39.96 ; 
      RECT 26.32 35.586 26.424 39.96 ; 
      RECT 25.888 35.586 25.992 39.96 ; 
      RECT 25.456 35.586 25.56 39.96 ; 
      RECT 25.024 35.586 25.128 39.96 ; 
      RECT 24.592 35.586 24.696 39.96 ; 
      RECT 24.16 35.586 24.264 39.96 ; 
      RECT 23.728 35.586 23.832 39.96 ; 
      RECT 23.296 35.586 23.4 39.96 ; 
      RECT 22.864 35.586 22.968 39.96 ; 
      RECT 22.432 35.586 22.536 39.96 ; 
      RECT 22 35.586 22.104 39.96 ; 
      RECT 21.568 35.586 21.672 39.96 ; 
      RECT 21.136 35.586 21.24 39.96 ; 
      RECT 20.704 35.586 20.808 39.96 ; 
      RECT 20.272 35.586 20.376 39.96 ; 
      RECT 19.84 35.586 19.944 39.96 ; 
      RECT 19.408 35.586 19.512 39.96 ; 
      RECT 18.976 35.586 19.08 39.96 ; 
      RECT 18.544 35.586 18.648 39.96 ; 
      RECT 18.112 35.586 18.216 39.96 ; 
      RECT 17.68 35.586 17.784 39.96 ; 
      RECT 17.248 35.586 17.352 39.96 ; 
      RECT 16.816 35.586 16.92 39.96 ; 
      RECT 16.384 35.586 16.488 39.96 ; 
      RECT 15.952 35.586 16.056 39.96 ; 
      RECT 15.52 35.586 15.624 39.96 ; 
      RECT 15.088 35.586 15.192 39.96 ; 
      RECT 14.656 35.586 14.76 39.96 ; 
      RECT 14.224 35.586 14.328 39.96 ; 
      RECT 13.792 35.586 13.896 39.96 ; 
      RECT 13.36 35.586 13.464 39.96 ; 
      RECT 12.928 35.586 13.032 39.96 ; 
      RECT 12.496 35.586 12.6 39.96 ; 
      RECT 12.064 35.586 12.168 39.96 ; 
      RECT 11.632 35.586 11.736 39.96 ; 
      RECT 11.2 35.586 11.304 39.96 ; 
      RECT 10.768 35.586 10.872 39.96 ; 
      RECT 10.336 35.586 10.44 39.96 ; 
      RECT 9.904 35.586 10.008 39.96 ; 
      RECT 9.472 35.586 9.576 39.96 ; 
      RECT 9.04 35.586 9.144 39.96 ; 
      RECT 8.608 35.586 8.712 39.96 ; 
      RECT 8.176 35.586 8.28 39.96 ; 
      RECT 7.744 35.586 7.848 39.96 ; 
      RECT 7.312 35.586 7.416 39.96 ; 
      RECT 6.88 35.586 6.984 39.96 ; 
      RECT 6.448 35.586 6.552 39.96 ; 
      RECT 6.016 35.586 6.12 39.96 ; 
      RECT 5.584 35.586 5.688 39.96 ; 
      RECT 5.152 35.586 5.256 39.96 ; 
      RECT 4.72 35.586 4.824 39.96 ; 
      RECT 4.288 35.586 4.392 39.96 ; 
      RECT 3.856 35.586 3.96 39.96 ; 
      RECT 3.424 35.586 3.528 39.96 ; 
      RECT 2.992 35.586 3.096 39.96 ; 
      RECT 2.56 35.586 2.664 39.96 ; 
      RECT 2.128 35.586 2.232 39.96 ; 
      RECT 1.696 35.586 1.8 39.96 ; 
      RECT 1.264 35.586 1.368 39.96 ; 
      RECT 0.832 35.586 0.936 39.96 ; 
      RECT 0.02 35.586 0.36 39.96 ; 
      RECT 62.212 39.906 62.724 44.28 ; 
      RECT 62.156 42.568 62.724 43.858 ; 
      RECT 61.276 41.476 61.812 44.28 ; 
      RECT 61.184 42.816 61.812 43.848 ; 
      RECT 61.276 39.906 61.668 44.28 ; 
      RECT 61.276 40.39 61.724 41.348 ; 
      RECT 61.276 39.906 61.812 40.262 ; 
      RECT 60.376 41.708 60.912 44.28 ; 
      RECT 60.376 39.906 60.768 44.28 ; 
      RECT 58.708 39.906 59.04 44.28 ; 
      RECT 58.708 40.26 59.096 44.002 ; 
      RECT 121.072 39.906 121.412 44.28 ; 
      RECT 120.496 39.906 120.6 44.28 ; 
      RECT 120.064 39.906 120.168 44.28 ; 
      RECT 119.632 39.906 119.736 44.28 ; 
      RECT 119.2 39.906 119.304 44.28 ; 
      RECT 118.768 39.906 118.872 44.28 ; 
      RECT 118.336 39.906 118.44 44.28 ; 
      RECT 117.904 39.906 118.008 44.28 ; 
      RECT 117.472 39.906 117.576 44.28 ; 
      RECT 117.04 39.906 117.144 44.28 ; 
      RECT 116.608 39.906 116.712 44.28 ; 
      RECT 116.176 39.906 116.28 44.28 ; 
      RECT 115.744 39.906 115.848 44.28 ; 
      RECT 115.312 39.906 115.416 44.28 ; 
      RECT 114.88 39.906 114.984 44.28 ; 
      RECT 114.448 39.906 114.552 44.28 ; 
      RECT 114.016 39.906 114.12 44.28 ; 
      RECT 113.584 39.906 113.688 44.28 ; 
      RECT 113.152 39.906 113.256 44.28 ; 
      RECT 112.72 39.906 112.824 44.28 ; 
      RECT 112.288 39.906 112.392 44.28 ; 
      RECT 111.856 39.906 111.96 44.28 ; 
      RECT 111.424 39.906 111.528 44.28 ; 
      RECT 110.992 39.906 111.096 44.28 ; 
      RECT 110.56 39.906 110.664 44.28 ; 
      RECT 110.128 39.906 110.232 44.28 ; 
      RECT 109.696 39.906 109.8 44.28 ; 
      RECT 109.264 39.906 109.368 44.28 ; 
      RECT 108.832 39.906 108.936 44.28 ; 
      RECT 108.4 39.906 108.504 44.28 ; 
      RECT 107.968 39.906 108.072 44.28 ; 
      RECT 107.536 39.906 107.64 44.28 ; 
      RECT 107.104 39.906 107.208 44.28 ; 
      RECT 106.672 39.906 106.776 44.28 ; 
      RECT 106.24 39.906 106.344 44.28 ; 
      RECT 105.808 39.906 105.912 44.28 ; 
      RECT 105.376 39.906 105.48 44.28 ; 
      RECT 104.944 39.906 105.048 44.28 ; 
      RECT 104.512 39.906 104.616 44.28 ; 
      RECT 104.08 39.906 104.184 44.28 ; 
      RECT 103.648 39.906 103.752 44.28 ; 
      RECT 103.216 39.906 103.32 44.28 ; 
      RECT 102.784 39.906 102.888 44.28 ; 
      RECT 102.352 39.906 102.456 44.28 ; 
      RECT 101.92 39.906 102.024 44.28 ; 
      RECT 101.488 39.906 101.592 44.28 ; 
      RECT 101.056 39.906 101.16 44.28 ; 
      RECT 100.624 39.906 100.728 44.28 ; 
      RECT 100.192 39.906 100.296 44.28 ; 
      RECT 99.76 39.906 99.864 44.28 ; 
      RECT 99.328 39.906 99.432 44.28 ; 
      RECT 98.896 39.906 99 44.28 ; 
      RECT 98.464 39.906 98.568 44.28 ; 
      RECT 98.032 39.906 98.136 44.28 ; 
      RECT 97.6 39.906 97.704 44.28 ; 
      RECT 97.168 39.906 97.272 44.28 ; 
      RECT 96.736 39.906 96.84 44.28 ; 
      RECT 96.304 39.906 96.408 44.28 ; 
      RECT 95.872 39.906 95.976 44.28 ; 
      RECT 95.44 39.906 95.544 44.28 ; 
      RECT 95.008 39.906 95.112 44.28 ; 
      RECT 94.576 39.906 94.68 44.28 ; 
      RECT 94.144 39.906 94.248 44.28 ; 
      RECT 93.712 39.906 93.816 44.28 ; 
      RECT 93.28 39.906 93.384 44.28 ; 
      RECT 92.848 39.906 92.952 44.28 ; 
      RECT 92.416 39.906 92.52 44.28 ; 
      RECT 91.984 39.906 92.088 44.28 ; 
      RECT 91.552 39.906 91.656 44.28 ; 
      RECT 91.12 39.906 91.224 44.28 ; 
      RECT 90.688 39.906 90.792 44.28 ; 
      RECT 90.256 39.906 90.36 44.28 ; 
      RECT 89.824 39.906 89.928 44.28 ; 
      RECT 89.392 39.906 89.496 44.28 ; 
      RECT 88.96 39.906 89.064 44.28 ; 
      RECT 88.528 39.906 88.632 44.28 ; 
      RECT 88.096 39.906 88.2 44.28 ; 
      RECT 87.664 39.906 87.768 44.28 ; 
      RECT 87.232 39.906 87.336 44.28 ; 
      RECT 86.8 39.906 86.904 44.28 ; 
      RECT 86.368 39.906 86.472 44.28 ; 
      RECT 85.936 39.906 86.04 44.28 ; 
      RECT 85.504 39.906 85.608 44.28 ; 
      RECT 85.072 39.906 85.176 44.28 ; 
      RECT 84.64 39.906 84.744 44.28 ; 
      RECT 84.208 39.906 84.312 44.28 ; 
      RECT 83.776 39.906 83.88 44.28 ; 
      RECT 83.344 39.906 83.448 44.28 ; 
      RECT 82.912 39.906 83.016 44.28 ; 
      RECT 82.48 39.906 82.584 44.28 ; 
      RECT 82.048 39.906 82.152 44.28 ; 
      RECT 81.616 39.906 81.72 44.28 ; 
      RECT 81.184 39.906 81.288 44.28 ; 
      RECT 80.752 39.906 80.856 44.28 ; 
      RECT 80.32 39.906 80.424 44.28 ; 
      RECT 79.888 39.906 79.992 44.28 ; 
      RECT 79.456 39.906 79.56 44.28 ; 
      RECT 79.024 39.906 79.128 44.28 ; 
      RECT 78.592 39.906 78.696 44.28 ; 
      RECT 78.16 39.906 78.264 44.28 ; 
      RECT 77.728 39.906 77.832 44.28 ; 
      RECT 77.296 39.906 77.4 44.28 ; 
      RECT 76.864 39.906 76.968 44.28 ; 
      RECT 76.432 39.906 76.536 44.28 ; 
      RECT 76 39.906 76.104 44.28 ; 
      RECT 75.568 39.906 75.672 44.28 ; 
      RECT 75.136 39.906 75.24 44.28 ; 
      RECT 74.704 39.906 74.808 44.28 ; 
      RECT 74.272 39.906 74.376 44.28 ; 
      RECT 73.84 39.906 73.944 44.28 ; 
      RECT 73.408 39.906 73.512 44.28 ; 
      RECT 72.976 39.906 73.08 44.28 ; 
      RECT 72.544 39.906 72.648 44.28 ; 
      RECT 72.112 39.906 72.216 44.28 ; 
      RECT 71.68 39.906 71.784 44.28 ; 
      RECT 71.248 39.906 71.352 44.28 ; 
      RECT 70.816 39.906 70.92 44.28 ; 
      RECT 70.384 39.906 70.488 44.28 ; 
      RECT 69.952 39.906 70.056 44.28 ; 
      RECT 69.52 39.906 69.624 44.28 ; 
      RECT 69.088 39.906 69.192 44.28 ; 
      RECT 68.656 39.906 68.76 44.28 ; 
      RECT 68.224 39.906 68.328 44.28 ; 
      RECT 67.792 39.906 67.896 44.28 ; 
      RECT 67.36 39.906 67.464 44.28 ; 
      RECT 66.928 39.906 67.032 44.28 ; 
      RECT 66.496 39.906 66.6 44.28 ; 
      RECT 66.064 39.906 66.168 44.28 ; 
      RECT 65.632 39.906 65.736 44.28 ; 
      RECT 65.2 39.906 65.304 44.28 ; 
      RECT 64.348 39.906 64.656 44.28 ; 
      RECT 56.776 39.906 57.084 44.28 ; 
      RECT 56.128 39.906 56.232 44.28 ; 
      RECT 55.696 39.906 55.8 44.28 ; 
      RECT 55.264 39.906 55.368 44.28 ; 
      RECT 54.832 39.906 54.936 44.28 ; 
      RECT 54.4 39.906 54.504 44.28 ; 
      RECT 53.968 39.906 54.072 44.28 ; 
      RECT 53.536 39.906 53.64 44.28 ; 
      RECT 53.104 39.906 53.208 44.28 ; 
      RECT 52.672 39.906 52.776 44.28 ; 
      RECT 52.24 39.906 52.344 44.28 ; 
      RECT 51.808 39.906 51.912 44.28 ; 
      RECT 51.376 39.906 51.48 44.28 ; 
      RECT 50.944 39.906 51.048 44.28 ; 
      RECT 50.512 39.906 50.616 44.28 ; 
      RECT 50.08 39.906 50.184 44.28 ; 
      RECT 49.648 39.906 49.752 44.28 ; 
      RECT 49.216 39.906 49.32 44.28 ; 
      RECT 48.784 39.906 48.888 44.28 ; 
      RECT 48.352 39.906 48.456 44.28 ; 
      RECT 47.92 39.906 48.024 44.28 ; 
      RECT 47.488 39.906 47.592 44.28 ; 
      RECT 47.056 39.906 47.16 44.28 ; 
      RECT 46.624 39.906 46.728 44.28 ; 
      RECT 46.192 39.906 46.296 44.28 ; 
      RECT 45.76 39.906 45.864 44.28 ; 
      RECT 45.328 39.906 45.432 44.28 ; 
      RECT 44.896 39.906 45 44.28 ; 
      RECT 44.464 39.906 44.568 44.28 ; 
      RECT 44.032 39.906 44.136 44.28 ; 
      RECT 43.6 39.906 43.704 44.28 ; 
      RECT 43.168 39.906 43.272 44.28 ; 
      RECT 42.736 39.906 42.84 44.28 ; 
      RECT 42.304 39.906 42.408 44.28 ; 
      RECT 41.872 39.906 41.976 44.28 ; 
      RECT 41.44 39.906 41.544 44.28 ; 
      RECT 41.008 39.906 41.112 44.28 ; 
      RECT 40.576 39.906 40.68 44.28 ; 
      RECT 40.144 39.906 40.248 44.28 ; 
      RECT 39.712 39.906 39.816 44.28 ; 
      RECT 39.28 39.906 39.384 44.28 ; 
      RECT 38.848 39.906 38.952 44.28 ; 
      RECT 38.416 39.906 38.52 44.28 ; 
      RECT 37.984 39.906 38.088 44.28 ; 
      RECT 37.552 39.906 37.656 44.28 ; 
      RECT 37.12 39.906 37.224 44.28 ; 
      RECT 36.688 39.906 36.792 44.28 ; 
      RECT 36.256 39.906 36.36 44.28 ; 
      RECT 35.824 39.906 35.928 44.28 ; 
      RECT 35.392 39.906 35.496 44.28 ; 
      RECT 34.96 39.906 35.064 44.28 ; 
      RECT 34.528 39.906 34.632 44.28 ; 
      RECT 34.096 39.906 34.2 44.28 ; 
      RECT 33.664 39.906 33.768 44.28 ; 
      RECT 33.232 39.906 33.336 44.28 ; 
      RECT 32.8 39.906 32.904 44.28 ; 
      RECT 32.368 39.906 32.472 44.28 ; 
      RECT 31.936 39.906 32.04 44.28 ; 
      RECT 31.504 39.906 31.608 44.28 ; 
      RECT 31.072 39.906 31.176 44.28 ; 
      RECT 30.64 39.906 30.744 44.28 ; 
      RECT 30.208 39.906 30.312 44.28 ; 
      RECT 29.776 39.906 29.88 44.28 ; 
      RECT 29.344 39.906 29.448 44.28 ; 
      RECT 28.912 39.906 29.016 44.28 ; 
      RECT 28.48 39.906 28.584 44.28 ; 
      RECT 28.048 39.906 28.152 44.28 ; 
      RECT 27.616 39.906 27.72 44.28 ; 
      RECT 27.184 39.906 27.288 44.28 ; 
      RECT 26.752 39.906 26.856 44.28 ; 
      RECT 26.32 39.906 26.424 44.28 ; 
      RECT 25.888 39.906 25.992 44.28 ; 
      RECT 25.456 39.906 25.56 44.28 ; 
      RECT 25.024 39.906 25.128 44.28 ; 
      RECT 24.592 39.906 24.696 44.28 ; 
      RECT 24.16 39.906 24.264 44.28 ; 
      RECT 23.728 39.906 23.832 44.28 ; 
      RECT 23.296 39.906 23.4 44.28 ; 
      RECT 22.864 39.906 22.968 44.28 ; 
      RECT 22.432 39.906 22.536 44.28 ; 
      RECT 22 39.906 22.104 44.28 ; 
      RECT 21.568 39.906 21.672 44.28 ; 
      RECT 21.136 39.906 21.24 44.28 ; 
      RECT 20.704 39.906 20.808 44.28 ; 
      RECT 20.272 39.906 20.376 44.28 ; 
      RECT 19.84 39.906 19.944 44.28 ; 
      RECT 19.408 39.906 19.512 44.28 ; 
      RECT 18.976 39.906 19.08 44.28 ; 
      RECT 18.544 39.906 18.648 44.28 ; 
      RECT 18.112 39.906 18.216 44.28 ; 
      RECT 17.68 39.906 17.784 44.28 ; 
      RECT 17.248 39.906 17.352 44.28 ; 
      RECT 16.816 39.906 16.92 44.28 ; 
      RECT 16.384 39.906 16.488 44.28 ; 
      RECT 15.952 39.906 16.056 44.28 ; 
      RECT 15.52 39.906 15.624 44.28 ; 
      RECT 15.088 39.906 15.192 44.28 ; 
      RECT 14.656 39.906 14.76 44.28 ; 
      RECT 14.224 39.906 14.328 44.28 ; 
      RECT 13.792 39.906 13.896 44.28 ; 
      RECT 13.36 39.906 13.464 44.28 ; 
      RECT 12.928 39.906 13.032 44.28 ; 
      RECT 12.496 39.906 12.6 44.28 ; 
      RECT 12.064 39.906 12.168 44.28 ; 
      RECT 11.632 39.906 11.736 44.28 ; 
      RECT 11.2 39.906 11.304 44.28 ; 
      RECT 10.768 39.906 10.872 44.28 ; 
      RECT 10.336 39.906 10.44 44.28 ; 
      RECT 9.904 39.906 10.008 44.28 ; 
      RECT 9.472 39.906 9.576 44.28 ; 
      RECT 9.04 39.906 9.144 44.28 ; 
      RECT 8.608 39.906 8.712 44.28 ; 
      RECT 8.176 39.906 8.28 44.28 ; 
      RECT 7.744 39.906 7.848 44.28 ; 
      RECT 7.312 39.906 7.416 44.28 ; 
      RECT 6.88 39.906 6.984 44.28 ; 
      RECT 6.448 39.906 6.552 44.28 ; 
      RECT 6.016 39.906 6.12 44.28 ; 
      RECT 5.584 39.906 5.688 44.28 ; 
      RECT 5.152 39.906 5.256 44.28 ; 
      RECT 4.72 39.906 4.824 44.28 ; 
      RECT 4.288 39.906 4.392 44.28 ; 
      RECT 3.856 39.906 3.96 44.28 ; 
      RECT 3.424 39.906 3.528 44.28 ; 
      RECT 2.992 39.906 3.096 44.28 ; 
      RECT 2.56 39.906 2.664 44.28 ; 
      RECT 2.128 39.906 2.232 44.28 ; 
      RECT 1.696 39.906 1.8 44.28 ; 
      RECT 1.264 39.906 1.368 44.28 ; 
      RECT 0.832 39.906 0.936 44.28 ; 
      RECT 0.02 39.906 0.36 44.28 ; 
      RECT 62.212 44.226 62.724 48.6 ; 
      RECT 62.156 46.888 62.724 48.178 ; 
      RECT 61.276 45.796 61.812 48.6 ; 
      RECT 61.184 47.136 61.812 48.168 ; 
      RECT 61.276 44.226 61.668 48.6 ; 
      RECT 61.276 44.71 61.724 45.668 ; 
      RECT 61.276 44.226 61.812 44.582 ; 
      RECT 60.376 46.028 60.912 48.6 ; 
      RECT 60.376 44.226 60.768 48.6 ; 
      RECT 58.708 44.226 59.04 48.6 ; 
      RECT 58.708 44.58 59.096 48.322 ; 
      RECT 121.072 44.226 121.412 48.6 ; 
      RECT 120.496 44.226 120.6 48.6 ; 
      RECT 120.064 44.226 120.168 48.6 ; 
      RECT 119.632 44.226 119.736 48.6 ; 
      RECT 119.2 44.226 119.304 48.6 ; 
      RECT 118.768 44.226 118.872 48.6 ; 
      RECT 118.336 44.226 118.44 48.6 ; 
      RECT 117.904 44.226 118.008 48.6 ; 
      RECT 117.472 44.226 117.576 48.6 ; 
      RECT 117.04 44.226 117.144 48.6 ; 
      RECT 116.608 44.226 116.712 48.6 ; 
      RECT 116.176 44.226 116.28 48.6 ; 
      RECT 115.744 44.226 115.848 48.6 ; 
      RECT 115.312 44.226 115.416 48.6 ; 
      RECT 114.88 44.226 114.984 48.6 ; 
      RECT 114.448 44.226 114.552 48.6 ; 
      RECT 114.016 44.226 114.12 48.6 ; 
      RECT 113.584 44.226 113.688 48.6 ; 
      RECT 113.152 44.226 113.256 48.6 ; 
      RECT 112.72 44.226 112.824 48.6 ; 
      RECT 112.288 44.226 112.392 48.6 ; 
      RECT 111.856 44.226 111.96 48.6 ; 
      RECT 111.424 44.226 111.528 48.6 ; 
      RECT 110.992 44.226 111.096 48.6 ; 
      RECT 110.56 44.226 110.664 48.6 ; 
      RECT 110.128 44.226 110.232 48.6 ; 
      RECT 109.696 44.226 109.8 48.6 ; 
      RECT 109.264 44.226 109.368 48.6 ; 
      RECT 108.832 44.226 108.936 48.6 ; 
      RECT 108.4 44.226 108.504 48.6 ; 
      RECT 107.968 44.226 108.072 48.6 ; 
      RECT 107.536 44.226 107.64 48.6 ; 
      RECT 107.104 44.226 107.208 48.6 ; 
      RECT 106.672 44.226 106.776 48.6 ; 
      RECT 106.24 44.226 106.344 48.6 ; 
      RECT 105.808 44.226 105.912 48.6 ; 
      RECT 105.376 44.226 105.48 48.6 ; 
      RECT 104.944 44.226 105.048 48.6 ; 
      RECT 104.512 44.226 104.616 48.6 ; 
      RECT 104.08 44.226 104.184 48.6 ; 
      RECT 103.648 44.226 103.752 48.6 ; 
      RECT 103.216 44.226 103.32 48.6 ; 
      RECT 102.784 44.226 102.888 48.6 ; 
      RECT 102.352 44.226 102.456 48.6 ; 
      RECT 101.92 44.226 102.024 48.6 ; 
      RECT 101.488 44.226 101.592 48.6 ; 
      RECT 101.056 44.226 101.16 48.6 ; 
      RECT 100.624 44.226 100.728 48.6 ; 
      RECT 100.192 44.226 100.296 48.6 ; 
      RECT 99.76 44.226 99.864 48.6 ; 
      RECT 99.328 44.226 99.432 48.6 ; 
      RECT 98.896 44.226 99 48.6 ; 
      RECT 98.464 44.226 98.568 48.6 ; 
      RECT 98.032 44.226 98.136 48.6 ; 
      RECT 97.6 44.226 97.704 48.6 ; 
      RECT 97.168 44.226 97.272 48.6 ; 
      RECT 96.736 44.226 96.84 48.6 ; 
      RECT 96.304 44.226 96.408 48.6 ; 
      RECT 95.872 44.226 95.976 48.6 ; 
      RECT 95.44 44.226 95.544 48.6 ; 
      RECT 95.008 44.226 95.112 48.6 ; 
      RECT 94.576 44.226 94.68 48.6 ; 
      RECT 94.144 44.226 94.248 48.6 ; 
      RECT 93.712 44.226 93.816 48.6 ; 
      RECT 93.28 44.226 93.384 48.6 ; 
      RECT 92.848 44.226 92.952 48.6 ; 
      RECT 92.416 44.226 92.52 48.6 ; 
      RECT 91.984 44.226 92.088 48.6 ; 
      RECT 91.552 44.226 91.656 48.6 ; 
      RECT 91.12 44.226 91.224 48.6 ; 
      RECT 90.688 44.226 90.792 48.6 ; 
      RECT 90.256 44.226 90.36 48.6 ; 
      RECT 89.824 44.226 89.928 48.6 ; 
      RECT 89.392 44.226 89.496 48.6 ; 
      RECT 88.96 44.226 89.064 48.6 ; 
      RECT 88.528 44.226 88.632 48.6 ; 
      RECT 88.096 44.226 88.2 48.6 ; 
      RECT 87.664 44.226 87.768 48.6 ; 
      RECT 87.232 44.226 87.336 48.6 ; 
      RECT 86.8 44.226 86.904 48.6 ; 
      RECT 86.368 44.226 86.472 48.6 ; 
      RECT 85.936 44.226 86.04 48.6 ; 
      RECT 85.504 44.226 85.608 48.6 ; 
      RECT 85.072 44.226 85.176 48.6 ; 
      RECT 84.64 44.226 84.744 48.6 ; 
      RECT 84.208 44.226 84.312 48.6 ; 
      RECT 83.776 44.226 83.88 48.6 ; 
      RECT 83.344 44.226 83.448 48.6 ; 
      RECT 82.912 44.226 83.016 48.6 ; 
      RECT 82.48 44.226 82.584 48.6 ; 
      RECT 82.048 44.226 82.152 48.6 ; 
      RECT 81.616 44.226 81.72 48.6 ; 
      RECT 81.184 44.226 81.288 48.6 ; 
      RECT 80.752 44.226 80.856 48.6 ; 
      RECT 80.32 44.226 80.424 48.6 ; 
      RECT 79.888 44.226 79.992 48.6 ; 
      RECT 79.456 44.226 79.56 48.6 ; 
      RECT 79.024 44.226 79.128 48.6 ; 
      RECT 78.592 44.226 78.696 48.6 ; 
      RECT 78.16 44.226 78.264 48.6 ; 
      RECT 77.728 44.226 77.832 48.6 ; 
      RECT 77.296 44.226 77.4 48.6 ; 
      RECT 76.864 44.226 76.968 48.6 ; 
      RECT 76.432 44.226 76.536 48.6 ; 
      RECT 76 44.226 76.104 48.6 ; 
      RECT 75.568 44.226 75.672 48.6 ; 
      RECT 75.136 44.226 75.24 48.6 ; 
      RECT 74.704 44.226 74.808 48.6 ; 
      RECT 74.272 44.226 74.376 48.6 ; 
      RECT 73.84 44.226 73.944 48.6 ; 
      RECT 73.408 44.226 73.512 48.6 ; 
      RECT 72.976 44.226 73.08 48.6 ; 
      RECT 72.544 44.226 72.648 48.6 ; 
      RECT 72.112 44.226 72.216 48.6 ; 
      RECT 71.68 44.226 71.784 48.6 ; 
      RECT 71.248 44.226 71.352 48.6 ; 
      RECT 70.816 44.226 70.92 48.6 ; 
      RECT 70.384 44.226 70.488 48.6 ; 
      RECT 69.952 44.226 70.056 48.6 ; 
      RECT 69.52 44.226 69.624 48.6 ; 
      RECT 69.088 44.226 69.192 48.6 ; 
      RECT 68.656 44.226 68.76 48.6 ; 
      RECT 68.224 44.226 68.328 48.6 ; 
      RECT 67.792 44.226 67.896 48.6 ; 
      RECT 67.36 44.226 67.464 48.6 ; 
      RECT 66.928 44.226 67.032 48.6 ; 
      RECT 66.496 44.226 66.6 48.6 ; 
      RECT 66.064 44.226 66.168 48.6 ; 
      RECT 65.632 44.226 65.736 48.6 ; 
      RECT 65.2 44.226 65.304 48.6 ; 
      RECT 64.348 44.226 64.656 48.6 ; 
      RECT 56.776 44.226 57.084 48.6 ; 
      RECT 56.128 44.226 56.232 48.6 ; 
      RECT 55.696 44.226 55.8 48.6 ; 
      RECT 55.264 44.226 55.368 48.6 ; 
      RECT 54.832 44.226 54.936 48.6 ; 
      RECT 54.4 44.226 54.504 48.6 ; 
      RECT 53.968 44.226 54.072 48.6 ; 
      RECT 53.536 44.226 53.64 48.6 ; 
      RECT 53.104 44.226 53.208 48.6 ; 
      RECT 52.672 44.226 52.776 48.6 ; 
      RECT 52.24 44.226 52.344 48.6 ; 
      RECT 51.808 44.226 51.912 48.6 ; 
      RECT 51.376 44.226 51.48 48.6 ; 
      RECT 50.944 44.226 51.048 48.6 ; 
      RECT 50.512 44.226 50.616 48.6 ; 
      RECT 50.08 44.226 50.184 48.6 ; 
      RECT 49.648 44.226 49.752 48.6 ; 
      RECT 49.216 44.226 49.32 48.6 ; 
      RECT 48.784 44.226 48.888 48.6 ; 
      RECT 48.352 44.226 48.456 48.6 ; 
      RECT 47.92 44.226 48.024 48.6 ; 
      RECT 47.488 44.226 47.592 48.6 ; 
      RECT 47.056 44.226 47.16 48.6 ; 
      RECT 46.624 44.226 46.728 48.6 ; 
      RECT 46.192 44.226 46.296 48.6 ; 
      RECT 45.76 44.226 45.864 48.6 ; 
      RECT 45.328 44.226 45.432 48.6 ; 
      RECT 44.896 44.226 45 48.6 ; 
      RECT 44.464 44.226 44.568 48.6 ; 
      RECT 44.032 44.226 44.136 48.6 ; 
      RECT 43.6 44.226 43.704 48.6 ; 
      RECT 43.168 44.226 43.272 48.6 ; 
      RECT 42.736 44.226 42.84 48.6 ; 
      RECT 42.304 44.226 42.408 48.6 ; 
      RECT 41.872 44.226 41.976 48.6 ; 
      RECT 41.44 44.226 41.544 48.6 ; 
      RECT 41.008 44.226 41.112 48.6 ; 
      RECT 40.576 44.226 40.68 48.6 ; 
      RECT 40.144 44.226 40.248 48.6 ; 
      RECT 39.712 44.226 39.816 48.6 ; 
      RECT 39.28 44.226 39.384 48.6 ; 
      RECT 38.848 44.226 38.952 48.6 ; 
      RECT 38.416 44.226 38.52 48.6 ; 
      RECT 37.984 44.226 38.088 48.6 ; 
      RECT 37.552 44.226 37.656 48.6 ; 
      RECT 37.12 44.226 37.224 48.6 ; 
      RECT 36.688 44.226 36.792 48.6 ; 
      RECT 36.256 44.226 36.36 48.6 ; 
      RECT 35.824 44.226 35.928 48.6 ; 
      RECT 35.392 44.226 35.496 48.6 ; 
      RECT 34.96 44.226 35.064 48.6 ; 
      RECT 34.528 44.226 34.632 48.6 ; 
      RECT 34.096 44.226 34.2 48.6 ; 
      RECT 33.664 44.226 33.768 48.6 ; 
      RECT 33.232 44.226 33.336 48.6 ; 
      RECT 32.8 44.226 32.904 48.6 ; 
      RECT 32.368 44.226 32.472 48.6 ; 
      RECT 31.936 44.226 32.04 48.6 ; 
      RECT 31.504 44.226 31.608 48.6 ; 
      RECT 31.072 44.226 31.176 48.6 ; 
      RECT 30.64 44.226 30.744 48.6 ; 
      RECT 30.208 44.226 30.312 48.6 ; 
      RECT 29.776 44.226 29.88 48.6 ; 
      RECT 29.344 44.226 29.448 48.6 ; 
      RECT 28.912 44.226 29.016 48.6 ; 
      RECT 28.48 44.226 28.584 48.6 ; 
      RECT 28.048 44.226 28.152 48.6 ; 
      RECT 27.616 44.226 27.72 48.6 ; 
      RECT 27.184 44.226 27.288 48.6 ; 
      RECT 26.752 44.226 26.856 48.6 ; 
      RECT 26.32 44.226 26.424 48.6 ; 
      RECT 25.888 44.226 25.992 48.6 ; 
      RECT 25.456 44.226 25.56 48.6 ; 
      RECT 25.024 44.226 25.128 48.6 ; 
      RECT 24.592 44.226 24.696 48.6 ; 
      RECT 24.16 44.226 24.264 48.6 ; 
      RECT 23.728 44.226 23.832 48.6 ; 
      RECT 23.296 44.226 23.4 48.6 ; 
      RECT 22.864 44.226 22.968 48.6 ; 
      RECT 22.432 44.226 22.536 48.6 ; 
      RECT 22 44.226 22.104 48.6 ; 
      RECT 21.568 44.226 21.672 48.6 ; 
      RECT 21.136 44.226 21.24 48.6 ; 
      RECT 20.704 44.226 20.808 48.6 ; 
      RECT 20.272 44.226 20.376 48.6 ; 
      RECT 19.84 44.226 19.944 48.6 ; 
      RECT 19.408 44.226 19.512 48.6 ; 
      RECT 18.976 44.226 19.08 48.6 ; 
      RECT 18.544 44.226 18.648 48.6 ; 
      RECT 18.112 44.226 18.216 48.6 ; 
      RECT 17.68 44.226 17.784 48.6 ; 
      RECT 17.248 44.226 17.352 48.6 ; 
      RECT 16.816 44.226 16.92 48.6 ; 
      RECT 16.384 44.226 16.488 48.6 ; 
      RECT 15.952 44.226 16.056 48.6 ; 
      RECT 15.52 44.226 15.624 48.6 ; 
      RECT 15.088 44.226 15.192 48.6 ; 
      RECT 14.656 44.226 14.76 48.6 ; 
      RECT 14.224 44.226 14.328 48.6 ; 
      RECT 13.792 44.226 13.896 48.6 ; 
      RECT 13.36 44.226 13.464 48.6 ; 
      RECT 12.928 44.226 13.032 48.6 ; 
      RECT 12.496 44.226 12.6 48.6 ; 
      RECT 12.064 44.226 12.168 48.6 ; 
      RECT 11.632 44.226 11.736 48.6 ; 
      RECT 11.2 44.226 11.304 48.6 ; 
      RECT 10.768 44.226 10.872 48.6 ; 
      RECT 10.336 44.226 10.44 48.6 ; 
      RECT 9.904 44.226 10.008 48.6 ; 
      RECT 9.472 44.226 9.576 48.6 ; 
      RECT 9.04 44.226 9.144 48.6 ; 
      RECT 8.608 44.226 8.712 48.6 ; 
      RECT 8.176 44.226 8.28 48.6 ; 
      RECT 7.744 44.226 7.848 48.6 ; 
      RECT 7.312 44.226 7.416 48.6 ; 
      RECT 6.88 44.226 6.984 48.6 ; 
      RECT 6.448 44.226 6.552 48.6 ; 
      RECT 6.016 44.226 6.12 48.6 ; 
      RECT 5.584 44.226 5.688 48.6 ; 
      RECT 5.152 44.226 5.256 48.6 ; 
      RECT 4.72 44.226 4.824 48.6 ; 
      RECT 4.288 44.226 4.392 48.6 ; 
      RECT 3.856 44.226 3.96 48.6 ; 
      RECT 3.424 44.226 3.528 48.6 ; 
      RECT 2.992 44.226 3.096 48.6 ; 
      RECT 2.56 44.226 2.664 48.6 ; 
      RECT 2.128 44.226 2.232 48.6 ; 
      RECT 1.696 44.226 1.8 48.6 ; 
      RECT 1.264 44.226 1.368 48.6 ; 
      RECT 0.832 44.226 0.936 48.6 ; 
      RECT 0.02 44.226 0.36 48.6 ; 
      RECT 62.212 48.546 62.724 52.92 ; 
      RECT 62.156 51.208 62.724 52.498 ; 
      RECT 61.276 50.116 61.812 52.92 ; 
      RECT 61.184 51.456 61.812 52.488 ; 
      RECT 61.276 48.546 61.668 52.92 ; 
      RECT 61.276 49.03 61.724 49.988 ; 
      RECT 61.276 48.546 61.812 48.902 ; 
      RECT 60.376 50.348 60.912 52.92 ; 
      RECT 60.376 48.546 60.768 52.92 ; 
      RECT 58.708 48.546 59.04 52.92 ; 
      RECT 58.708 48.9 59.096 52.642 ; 
      RECT 121.072 48.546 121.412 52.92 ; 
      RECT 120.496 48.546 120.6 52.92 ; 
      RECT 120.064 48.546 120.168 52.92 ; 
      RECT 119.632 48.546 119.736 52.92 ; 
      RECT 119.2 48.546 119.304 52.92 ; 
      RECT 118.768 48.546 118.872 52.92 ; 
      RECT 118.336 48.546 118.44 52.92 ; 
      RECT 117.904 48.546 118.008 52.92 ; 
      RECT 117.472 48.546 117.576 52.92 ; 
      RECT 117.04 48.546 117.144 52.92 ; 
      RECT 116.608 48.546 116.712 52.92 ; 
      RECT 116.176 48.546 116.28 52.92 ; 
      RECT 115.744 48.546 115.848 52.92 ; 
      RECT 115.312 48.546 115.416 52.92 ; 
      RECT 114.88 48.546 114.984 52.92 ; 
      RECT 114.448 48.546 114.552 52.92 ; 
      RECT 114.016 48.546 114.12 52.92 ; 
      RECT 113.584 48.546 113.688 52.92 ; 
      RECT 113.152 48.546 113.256 52.92 ; 
      RECT 112.72 48.546 112.824 52.92 ; 
      RECT 112.288 48.546 112.392 52.92 ; 
      RECT 111.856 48.546 111.96 52.92 ; 
      RECT 111.424 48.546 111.528 52.92 ; 
      RECT 110.992 48.546 111.096 52.92 ; 
      RECT 110.56 48.546 110.664 52.92 ; 
      RECT 110.128 48.546 110.232 52.92 ; 
      RECT 109.696 48.546 109.8 52.92 ; 
      RECT 109.264 48.546 109.368 52.92 ; 
      RECT 108.832 48.546 108.936 52.92 ; 
      RECT 108.4 48.546 108.504 52.92 ; 
      RECT 107.968 48.546 108.072 52.92 ; 
      RECT 107.536 48.546 107.64 52.92 ; 
      RECT 107.104 48.546 107.208 52.92 ; 
      RECT 106.672 48.546 106.776 52.92 ; 
      RECT 106.24 48.546 106.344 52.92 ; 
      RECT 105.808 48.546 105.912 52.92 ; 
      RECT 105.376 48.546 105.48 52.92 ; 
      RECT 104.944 48.546 105.048 52.92 ; 
      RECT 104.512 48.546 104.616 52.92 ; 
      RECT 104.08 48.546 104.184 52.92 ; 
      RECT 103.648 48.546 103.752 52.92 ; 
      RECT 103.216 48.546 103.32 52.92 ; 
      RECT 102.784 48.546 102.888 52.92 ; 
      RECT 102.352 48.546 102.456 52.92 ; 
      RECT 101.92 48.546 102.024 52.92 ; 
      RECT 101.488 48.546 101.592 52.92 ; 
      RECT 101.056 48.546 101.16 52.92 ; 
      RECT 100.624 48.546 100.728 52.92 ; 
      RECT 100.192 48.546 100.296 52.92 ; 
      RECT 99.76 48.546 99.864 52.92 ; 
      RECT 99.328 48.546 99.432 52.92 ; 
      RECT 98.896 48.546 99 52.92 ; 
      RECT 98.464 48.546 98.568 52.92 ; 
      RECT 98.032 48.546 98.136 52.92 ; 
      RECT 97.6 48.546 97.704 52.92 ; 
      RECT 97.168 48.546 97.272 52.92 ; 
      RECT 96.736 48.546 96.84 52.92 ; 
      RECT 96.304 48.546 96.408 52.92 ; 
      RECT 95.872 48.546 95.976 52.92 ; 
      RECT 95.44 48.546 95.544 52.92 ; 
      RECT 95.008 48.546 95.112 52.92 ; 
      RECT 94.576 48.546 94.68 52.92 ; 
      RECT 94.144 48.546 94.248 52.92 ; 
      RECT 93.712 48.546 93.816 52.92 ; 
      RECT 93.28 48.546 93.384 52.92 ; 
      RECT 92.848 48.546 92.952 52.92 ; 
      RECT 92.416 48.546 92.52 52.92 ; 
      RECT 91.984 48.546 92.088 52.92 ; 
      RECT 91.552 48.546 91.656 52.92 ; 
      RECT 91.12 48.546 91.224 52.92 ; 
      RECT 90.688 48.546 90.792 52.92 ; 
      RECT 90.256 48.546 90.36 52.92 ; 
      RECT 89.824 48.546 89.928 52.92 ; 
      RECT 89.392 48.546 89.496 52.92 ; 
      RECT 88.96 48.546 89.064 52.92 ; 
      RECT 88.528 48.546 88.632 52.92 ; 
      RECT 88.096 48.546 88.2 52.92 ; 
      RECT 87.664 48.546 87.768 52.92 ; 
      RECT 87.232 48.546 87.336 52.92 ; 
      RECT 86.8 48.546 86.904 52.92 ; 
      RECT 86.368 48.546 86.472 52.92 ; 
      RECT 85.936 48.546 86.04 52.92 ; 
      RECT 85.504 48.546 85.608 52.92 ; 
      RECT 85.072 48.546 85.176 52.92 ; 
      RECT 84.64 48.546 84.744 52.92 ; 
      RECT 84.208 48.546 84.312 52.92 ; 
      RECT 83.776 48.546 83.88 52.92 ; 
      RECT 83.344 48.546 83.448 52.92 ; 
      RECT 82.912 48.546 83.016 52.92 ; 
      RECT 82.48 48.546 82.584 52.92 ; 
      RECT 82.048 48.546 82.152 52.92 ; 
      RECT 81.616 48.546 81.72 52.92 ; 
      RECT 81.184 48.546 81.288 52.92 ; 
      RECT 80.752 48.546 80.856 52.92 ; 
      RECT 80.32 48.546 80.424 52.92 ; 
      RECT 79.888 48.546 79.992 52.92 ; 
      RECT 79.456 48.546 79.56 52.92 ; 
      RECT 79.024 48.546 79.128 52.92 ; 
      RECT 78.592 48.546 78.696 52.92 ; 
      RECT 78.16 48.546 78.264 52.92 ; 
      RECT 77.728 48.546 77.832 52.92 ; 
      RECT 77.296 48.546 77.4 52.92 ; 
      RECT 76.864 48.546 76.968 52.92 ; 
      RECT 76.432 48.546 76.536 52.92 ; 
      RECT 76 48.546 76.104 52.92 ; 
      RECT 75.568 48.546 75.672 52.92 ; 
      RECT 75.136 48.546 75.24 52.92 ; 
      RECT 74.704 48.546 74.808 52.92 ; 
      RECT 74.272 48.546 74.376 52.92 ; 
      RECT 73.84 48.546 73.944 52.92 ; 
      RECT 73.408 48.546 73.512 52.92 ; 
      RECT 72.976 48.546 73.08 52.92 ; 
      RECT 72.544 48.546 72.648 52.92 ; 
      RECT 72.112 48.546 72.216 52.92 ; 
      RECT 71.68 48.546 71.784 52.92 ; 
      RECT 71.248 48.546 71.352 52.92 ; 
      RECT 70.816 48.546 70.92 52.92 ; 
      RECT 70.384 48.546 70.488 52.92 ; 
      RECT 69.952 48.546 70.056 52.92 ; 
      RECT 69.52 48.546 69.624 52.92 ; 
      RECT 69.088 48.546 69.192 52.92 ; 
      RECT 68.656 48.546 68.76 52.92 ; 
      RECT 68.224 48.546 68.328 52.92 ; 
      RECT 67.792 48.546 67.896 52.92 ; 
      RECT 67.36 48.546 67.464 52.92 ; 
      RECT 66.928 48.546 67.032 52.92 ; 
      RECT 66.496 48.546 66.6 52.92 ; 
      RECT 66.064 48.546 66.168 52.92 ; 
      RECT 65.632 48.546 65.736 52.92 ; 
      RECT 65.2 48.546 65.304 52.92 ; 
      RECT 64.348 48.546 64.656 52.92 ; 
      RECT 56.776 48.546 57.084 52.92 ; 
      RECT 56.128 48.546 56.232 52.92 ; 
      RECT 55.696 48.546 55.8 52.92 ; 
      RECT 55.264 48.546 55.368 52.92 ; 
      RECT 54.832 48.546 54.936 52.92 ; 
      RECT 54.4 48.546 54.504 52.92 ; 
      RECT 53.968 48.546 54.072 52.92 ; 
      RECT 53.536 48.546 53.64 52.92 ; 
      RECT 53.104 48.546 53.208 52.92 ; 
      RECT 52.672 48.546 52.776 52.92 ; 
      RECT 52.24 48.546 52.344 52.92 ; 
      RECT 51.808 48.546 51.912 52.92 ; 
      RECT 51.376 48.546 51.48 52.92 ; 
      RECT 50.944 48.546 51.048 52.92 ; 
      RECT 50.512 48.546 50.616 52.92 ; 
      RECT 50.08 48.546 50.184 52.92 ; 
      RECT 49.648 48.546 49.752 52.92 ; 
      RECT 49.216 48.546 49.32 52.92 ; 
      RECT 48.784 48.546 48.888 52.92 ; 
      RECT 48.352 48.546 48.456 52.92 ; 
      RECT 47.92 48.546 48.024 52.92 ; 
      RECT 47.488 48.546 47.592 52.92 ; 
      RECT 47.056 48.546 47.16 52.92 ; 
      RECT 46.624 48.546 46.728 52.92 ; 
      RECT 46.192 48.546 46.296 52.92 ; 
      RECT 45.76 48.546 45.864 52.92 ; 
      RECT 45.328 48.546 45.432 52.92 ; 
      RECT 44.896 48.546 45 52.92 ; 
      RECT 44.464 48.546 44.568 52.92 ; 
      RECT 44.032 48.546 44.136 52.92 ; 
      RECT 43.6 48.546 43.704 52.92 ; 
      RECT 43.168 48.546 43.272 52.92 ; 
      RECT 42.736 48.546 42.84 52.92 ; 
      RECT 42.304 48.546 42.408 52.92 ; 
      RECT 41.872 48.546 41.976 52.92 ; 
      RECT 41.44 48.546 41.544 52.92 ; 
      RECT 41.008 48.546 41.112 52.92 ; 
      RECT 40.576 48.546 40.68 52.92 ; 
      RECT 40.144 48.546 40.248 52.92 ; 
      RECT 39.712 48.546 39.816 52.92 ; 
      RECT 39.28 48.546 39.384 52.92 ; 
      RECT 38.848 48.546 38.952 52.92 ; 
      RECT 38.416 48.546 38.52 52.92 ; 
      RECT 37.984 48.546 38.088 52.92 ; 
      RECT 37.552 48.546 37.656 52.92 ; 
      RECT 37.12 48.546 37.224 52.92 ; 
      RECT 36.688 48.546 36.792 52.92 ; 
      RECT 36.256 48.546 36.36 52.92 ; 
      RECT 35.824 48.546 35.928 52.92 ; 
      RECT 35.392 48.546 35.496 52.92 ; 
      RECT 34.96 48.546 35.064 52.92 ; 
      RECT 34.528 48.546 34.632 52.92 ; 
      RECT 34.096 48.546 34.2 52.92 ; 
      RECT 33.664 48.546 33.768 52.92 ; 
      RECT 33.232 48.546 33.336 52.92 ; 
      RECT 32.8 48.546 32.904 52.92 ; 
      RECT 32.368 48.546 32.472 52.92 ; 
      RECT 31.936 48.546 32.04 52.92 ; 
      RECT 31.504 48.546 31.608 52.92 ; 
      RECT 31.072 48.546 31.176 52.92 ; 
      RECT 30.64 48.546 30.744 52.92 ; 
      RECT 30.208 48.546 30.312 52.92 ; 
      RECT 29.776 48.546 29.88 52.92 ; 
      RECT 29.344 48.546 29.448 52.92 ; 
      RECT 28.912 48.546 29.016 52.92 ; 
      RECT 28.48 48.546 28.584 52.92 ; 
      RECT 28.048 48.546 28.152 52.92 ; 
      RECT 27.616 48.546 27.72 52.92 ; 
      RECT 27.184 48.546 27.288 52.92 ; 
      RECT 26.752 48.546 26.856 52.92 ; 
      RECT 26.32 48.546 26.424 52.92 ; 
      RECT 25.888 48.546 25.992 52.92 ; 
      RECT 25.456 48.546 25.56 52.92 ; 
      RECT 25.024 48.546 25.128 52.92 ; 
      RECT 24.592 48.546 24.696 52.92 ; 
      RECT 24.16 48.546 24.264 52.92 ; 
      RECT 23.728 48.546 23.832 52.92 ; 
      RECT 23.296 48.546 23.4 52.92 ; 
      RECT 22.864 48.546 22.968 52.92 ; 
      RECT 22.432 48.546 22.536 52.92 ; 
      RECT 22 48.546 22.104 52.92 ; 
      RECT 21.568 48.546 21.672 52.92 ; 
      RECT 21.136 48.546 21.24 52.92 ; 
      RECT 20.704 48.546 20.808 52.92 ; 
      RECT 20.272 48.546 20.376 52.92 ; 
      RECT 19.84 48.546 19.944 52.92 ; 
      RECT 19.408 48.546 19.512 52.92 ; 
      RECT 18.976 48.546 19.08 52.92 ; 
      RECT 18.544 48.546 18.648 52.92 ; 
      RECT 18.112 48.546 18.216 52.92 ; 
      RECT 17.68 48.546 17.784 52.92 ; 
      RECT 17.248 48.546 17.352 52.92 ; 
      RECT 16.816 48.546 16.92 52.92 ; 
      RECT 16.384 48.546 16.488 52.92 ; 
      RECT 15.952 48.546 16.056 52.92 ; 
      RECT 15.52 48.546 15.624 52.92 ; 
      RECT 15.088 48.546 15.192 52.92 ; 
      RECT 14.656 48.546 14.76 52.92 ; 
      RECT 14.224 48.546 14.328 52.92 ; 
      RECT 13.792 48.546 13.896 52.92 ; 
      RECT 13.36 48.546 13.464 52.92 ; 
      RECT 12.928 48.546 13.032 52.92 ; 
      RECT 12.496 48.546 12.6 52.92 ; 
      RECT 12.064 48.546 12.168 52.92 ; 
      RECT 11.632 48.546 11.736 52.92 ; 
      RECT 11.2 48.546 11.304 52.92 ; 
      RECT 10.768 48.546 10.872 52.92 ; 
      RECT 10.336 48.546 10.44 52.92 ; 
      RECT 9.904 48.546 10.008 52.92 ; 
      RECT 9.472 48.546 9.576 52.92 ; 
      RECT 9.04 48.546 9.144 52.92 ; 
      RECT 8.608 48.546 8.712 52.92 ; 
      RECT 8.176 48.546 8.28 52.92 ; 
      RECT 7.744 48.546 7.848 52.92 ; 
      RECT 7.312 48.546 7.416 52.92 ; 
      RECT 6.88 48.546 6.984 52.92 ; 
      RECT 6.448 48.546 6.552 52.92 ; 
      RECT 6.016 48.546 6.12 52.92 ; 
      RECT 5.584 48.546 5.688 52.92 ; 
      RECT 5.152 48.546 5.256 52.92 ; 
      RECT 4.72 48.546 4.824 52.92 ; 
      RECT 4.288 48.546 4.392 52.92 ; 
      RECT 3.856 48.546 3.96 52.92 ; 
      RECT 3.424 48.546 3.528 52.92 ; 
      RECT 2.992 48.546 3.096 52.92 ; 
      RECT 2.56 48.546 2.664 52.92 ; 
      RECT 2.128 48.546 2.232 52.92 ; 
      RECT 1.696 48.546 1.8 52.92 ; 
      RECT 1.264 48.546 1.368 52.92 ; 
      RECT 0.832 48.546 0.936 52.92 ; 
      RECT 0.02 48.546 0.36 52.92 ; 
      RECT 62.212 52.866 62.724 57.24 ; 
      RECT 62.156 55.528 62.724 56.818 ; 
      RECT 61.276 54.436 61.812 57.24 ; 
      RECT 61.184 55.776 61.812 56.808 ; 
      RECT 61.276 52.866 61.668 57.24 ; 
      RECT 61.276 53.35 61.724 54.308 ; 
      RECT 61.276 52.866 61.812 53.222 ; 
      RECT 60.376 54.668 60.912 57.24 ; 
      RECT 60.376 52.866 60.768 57.24 ; 
      RECT 58.708 52.866 59.04 57.24 ; 
      RECT 58.708 53.22 59.096 56.962 ; 
      RECT 121.072 52.866 121.412 57.24 ; 
      RECT 120.496 52.866 120.6 57.24 ; 
      RECT 120.064 52.866 120.168 57.24 ; 
      RECT 119.632 52.866 119.736 57.24 ; 
      RECT 119.2 52.866 119.304 57.24 ; 
      RECT 118.768 52.866 118.872 57.24 ; 
      RECT 118.336 52.866 118.44 57.24 ; 
      RECT 117.904 52.866 118.008 57.24 ; 
      RECT 117.472 52.866 117.576 57.24 ; 
      RECT 117.04 52.866 117.144 57.24 ; 
      RECT 116.608 52.866 116.712 57.24 ; 
      RECT 116.176 52.866 116.28 57.24 ; 
      RECT 115.744 52.866 115.848 57.24 ; 
      RECT 115.312 52.866 115.416 57.24 ; 
      RECT 114.88 52.866 114.984 57.24 ; 
      RECT 114.448 52.866 114.552 57.24 ; 
      RECT 114.016 52.866 114.12 57.24 ; 
      RECT 113.584 52.866 113.688 57.24 ; 
      RECT 113.152 52.866 113.256 57.24 ; 
      RECT 112.72 52.866 112.824 57.24 ; 
      RECT 112.288 52.866 112.392 57.24 ; 
      RECT 111.856 52.866 111.96 57.24 ; 
      RECT 111.424 52.866 111.528 57.24 ; 
      RECT 110.992 52.866 111.096 57.24 ; 
      RECT 110.56 52.866 110.664 57.24 ; 
      RECT 110.128 52.866 110.232 57.24 ; 
      RECT 109.696 52.866 109.8 57.24 ; 
      RECT 109.264 52.866 109.368 57.24 ; 
      RECT 108.832 52.866 108.936 57.24 ; 
      RECT 108.4 52.866 108.504 57.24 ; 
      RECT 107.968 52.866 108.072 57.24 ; 
      RECT 107.536 52.866 107.64 57.24 ; 
      RECT 107.104 52.866 107.208 57.24 ; 
      RECT 106.672 52.866 106.776 57.24 ; 
      RECT 106.24 52.866 106.344 57.24 ; 
      RECT 105.808 52.866 105.912 57.24 ; 
      RECT 105.376 52.866 105.48 57.24 ; 
      RECT 104.944 52.866 105.048 57.24 ; 
      RECT 104.512 52.866 104.616 57.24 ; 
      RECT 104.08 52.866 104.184 57.24 ; 
      RECT 103.648 52.866 103.752 57.24 ; 
      RECT 103.216 52.866 103.32 57.24 ; 
      RECT 102.784 52.866 102.888 57.24 ; 
      RECT 102.352 52.866 102.456 57.24 ; 
      RECT 101.92 52.866 102.024 57.24 ; 
      RECT 101.488 52.866 101.592 57.24 ; 
      RECT 101.056 52.866 101.16 57.24 ; 
      RECT 100.624 52.866 100.728 57.24 ; 
      RECT 100.192 52.866 100.296 57.24 ; 
      RECT 99.76 52.866 99.864 57.24 ; 
      RECT 99.328 52.866 99.432 57.24 ; 
      RECT 98.896 52.866 99 57.24 ; 
      RECT 98.464 52.866 98.568 57.24 ; 
      RECT 98.032 52.866 98.136 57.24 ; 
      RECT 97.6 52.866 97.704 57.24 ; 
      RECT 97.168 52.866 97.272 57.24 ; 
      RECT 96.736 52.866 96.84 57.24 ; 
      RECT 96.304 52.866 96.408 57.24 ; 
      RECT 95.872 52.866 95.976 57.24 ; 
      RECT 95.44 52.866 95.544 57.24 ; 
      RECT 95.008 52.866 95.112 57.24 ; 
      RECT 94.576 52.866 94.68 57.24 ; 
      RECT 94.144 52.866 94.248 57.24 ; 
      RECT 93.712 52.866 93.816 57.24 ; 
      RECT 93.28 52.866 93.384 57.24 ; 
      RECT 92.848 52.866 92.952 57.24 ; 
      RECT 92.416 52.866 92.52 57.24 ; 
      RECT 91.984 52.866 92.088 57.24 ; 
      RECT 91.552 52.866 91.656 57.24 ; 
      RECT 91.12 52.866 91.224 57.24 ; 
      RECT 90.688 52.866 90.792 57.24 ; 
      RECT 90.256 52.866 90.36 57.24 ; 
      RECT 89.824 52.866 89.928 57.24 ; 
      RECT 89.392 52.866 89.496 57.24 ; 
      RECT 88.96 52.866 89.064 57.24 ; 
      RECT 88.528 52.866 88.632 57.24 ; 
      RECT 88.096 52.866 88.2 57.24 ; 
      RECT 87.664 52.866 87.768 57.24 ; 
      RECT 87.232 52.866 87.336 57.24 ; 
      RECT 86.8 52.866 86.904 57.24 ; 
      RECT 86.368 52.866 86.472 57.24 ; 
      RECT 85.936 52.866 86.04 57.24 ; 
      RECT 85.504 52.866 85.608 57.24 ; 
      RECT 85.072 52.866 85.176 57.24 ; 
      RECT 84.64 52.866 84.744 57.24 ; 
      RECT 84.208 52.866 84.312 57.24 ; 
      RECT 83.776 52.866 83.88 57.24 ; 
      RECT 83.344 52.866 83.448 57.24 ; 
      RECT 82.912 52.866 83.016 57.24 ; 
      RECT 82.48 52.866 82.584 57.24 ; 
      RECT 82.048 52.866 82.152 57.24 ; 
      RECT 81.616 52.866 81.72 57.24 ; 
      RECT 81.184 52.866 81.288 57.24 ; 
      RECT 80.752 52.866 80.856 57.24 ; 
      RECT 80.32 52.866 80.424 57.24 ; 
      RECT 79.888 52.866 79.992 57.24 ; 
      RECT 79.456 52.866 79.56 57.24 ; 
      RECT 79.024 52.866 79.128 57.24 ; 
      RECT 78.592 52.866 78.696 57.24 ; 
      RECT 78.16 52.866 78.264 57.24 ; 
      RECT 77.728 52.866 77.832 57.24 ; 
      RECT 77.296 52.866 77.4 57.24 ; 
      RECT 76.864 52.866 76.968 57.24 ; 
      RECT 76.432 52.866 76.536 57.24 ; 
      RECT 76 52.866 76.104 57.24 ; 
      RECT 75.568 52.866 75.672 57.24 ; 
      RECT 75.136 52.866 75.24 57.24 ; 
      RECT 74.704 52.866 74.808 57.24 ; 
      RECT 74.272 52.866 74.376 57.24 ; 
      RECT 73.84 52.866 73.944 57.24 ; 
      RECT 73.408 52.866 73.512 57.24 ; 
      RECT 72.976 52.866 73.08 57.24 ; 
      RECT 72.544 52.866 72.648 57.24 ; 
      RECT 72.112 52.866 72.216 57.24 ; 
      RECT 71.68 52.866 71.784 57.24 ; 
      RECT 71.248 52.866 71.352 57.24 ; 
      RECT 70.816 52.866 70.92 57.24 ; 
      RECT 70.384 52.866 70.488 57.24 ; 
      RECT 69.952 52.866 70.056 57.24 ; 
      RECT 69.52 52.866 69.624 57.24 ; 
      RECT 69.088 52.866 69.192 57.24 ; 
      RECT 68.656 52.866 68.76 57.24 ; 
      RECT 68.224 52.866 68.328 57.24 ; 
      RECT 67.792 52.866 67.896 57.24 ; 
      RECT 67.36 52.866 67.464 57.24 ; 
      RECT 66.928 52.866 67.032 57.24 ; 
      RECT 66.496 52.866 66.6 57.24 ; 
      RECT 66.064 52.866 66.168 57.24 ; 
      RECT 65.632 52.866 65.736 57.24 ; 
      RECT 65.2 52.866 65.304 57.24 ; 
      RECT 64.348 52.866 64.656 57.24 ; 
      RECT 56.776 52.866 57.084 57.24 ; 
      RECT 56.128 52.866 56.232 57.24 ; 
      RECT 55.696 52.866 55.8 57.24 ; 
      RECT 55.264 52.866 55.368 57.24 ; 
      RECT 54.832 52.866 54.936 57.24 ; 
      RECT 54.4 52.866 54.504 57.24 ; 
      RECT 53.968 52.866 54.072 57.24 ; 
      RECT 53.536 52.866 53.64 57.24 ; 
      RECT 53.104 52.866 53.208 57.24 ; 
      RECT 52.672 52.866 52.776 57.24 ; 
      RECT 52.24 52.866 52.344 57.24 ; 
      RECT 51.808 52.866 51.912 57.24 ; 
      RECT 51.376 52.866 51.48 57.24 ; 
      RECT 50.944 52.866 51.048 57.24 ; 
      RECT 50.512 52.866 50.616 57.24 ; 
      RECT 50.08 52.866 50.184 57.24 ; 
      RECT 49.648 52.866 49.752 57.24 ; 
      RECT 49.216 52.866 49.32 57.24 ; 
      RECT 48.784 52.866 48.888 57.24 ; 
      RECT 48.352 52.866 48.456 57.24 ; 
      RECT 47.92 52.866 48.024 57.24 ; 
      RECT 47.488 52.866 47.592 57.24 ; 
      RECT 47.056 52.866 47.16 57.24 ; 
      RECT 46.624 52.866 46.728 57.24 ; 
      RECT 46.192 52.866 46.296 57.24 ; 
      RECT 45.76 52.866 45.864 57.24 ; 
      RECT 45.328 52.866 45.432 57.24 ; 
      RECT 44.896 52.866 45 57.24 ; 
      RECT 44.464 52.866 44.568 57.24 ; 
      RECT 44.032 52.866 44.136 57.24 ; 
      RECT 43.6 52.866 43.704 57.24 ; 
      RECT 43.168 52.866 43.272 57.24 ; 
      RECT 42.736 52.866 42.84 57.24 ; 
      RECT 42.304 52.866 42.408 57.24 ; 
      RECT 41.872 52.866 41.976 57.24 ; 
      RECT 41.44 52.866 41.544 57.24 ; 
      RECT 41.008 52.866 41.112 57.24 ; 
      RECT 40.576 52.866 40.68 57.24 ; 
      RECT 40.144 52.866 40.248 57.24 ; 
      RECT 39.712 52.866 39.816 57.24 ; 
      RECT 39.28 52.866 39.384 57.24 ; 
      RECT 38.848 52.866 38.952 57.24 ; 
      RECT 38.416 52.866 38.52 57.24 ; 
      RECT 37.984 52.866 38.088 57.24 ; 
      RECT 37.552 52.866 37.656 57.24 ; 
      RECT 37.12 52.866 37.224 57.24 ; 
      RECT 36.688 52.866 36.792 57.24 ; 
      RECT 36.256 52.866 36.36 57.24 ; 
      RECT 35.824 52.866 35.928 57.24 ; 
      RECT 35.392 52.866 35.496 57.24 ; 
      RECT 34.96 52.866 35.064 57.24 ; 
      RECT 34.528 52.866 34.632 57.24 ; 
      RECT 34.096 52.866 34.2 57.24 ; 
      RECT 33.664 52.866 33.768 57.24 ; 
      RECT 33.232 52.866 33.336 57.24 ; 
      RECT 32.8 52.866 32.904 57.24 ; 
      RECT 32.368 52.866 32.472 57.24 ; 
      RECT 31.936 52.866 32.04 57.24 ; 
      RECT 31.504 52.866 31.608 57.24 ; 
      RECT 31.072 52.866 31.176 57.24 ; 
      RECT 30.64 52.866 30.744 57.24 ; 
      RECT 30.208 52.866 30.312 57.24 ; 
      RECT 29.776 52.866 29.88 57.24 ; 
      RECT 29.344 52.866 29.448 57.24 ; 
      RECT 28.912 52.866 29.016 57.24 ; 
      RECT 28.48 52.866 28.584 57.24 ; 
      RECT 28.048 52.866 28.152 57.24 ; 
      RECT 27.616 52.866 27.72 57.24 ; 
      RECT 27.184 52.866 27.288 57.24 ; 
      RECT 26.752 52.866 26.856 57.24 ; 
      RECT 26.32 52.866 26.424 57.24 ; 
      RECT 25.888 52.866 25.992 57.24 ; 
      RECT 25.456 52.866 25.56 57.24 ; 
      RECT 25.024 52.866 25.128 57.24 ; 
      RECT 24.592 52.866 24.696 57.24 ; 
      RECT 24.16 52.866 24.264 57.24 ; 
      RECT 23.728 52.866 23.832 57.24 ; 
      RECT 23.296 52.866 23.4 57.24 ; 
      RECT 22.864 52.866 22.968 57.24 ; 
      RECT 22.432 52.866 22.536 57.24 ; 
      RECT 22 52.866 22.104 57.24 ; 
      RECT 21.568 52.866 21.672 57.24 ; 
      RECT 21.136 52.866 21.24 57.24 ; 
      RECT 20.704 52.866 20.808 57.24 ; 
      RECT 20.272 52.866 20.376 57.24 ; 
      RECT 19.84 52.866 19.944 57.24 ; 
      RECT 19.408 52.866 19.512 57.24 ; 
      RECT 18.976 52.866 19.08 57.24 ; 
      RECT 18.544 52.866 18.648 57.24 ; 
      RECT 18.112 52.866 18.216 57.24 ; 
      RECT 17.68 52.866 17.784 57.24 ; 
      RECT 17.248 52.866 17.352 57.24 ; 
      RECT 16.816 52.866 16.92 57.24 ; 
      RECT 16.384 52.866 16.488 57.24 ; 
      RECT 15.952 52.866 16.056 57.24 ; 
      RECT 15.52 52.866 15.624 57.24 ; 
      RECT 15.088 52.866 15.192 57.24 ; 
      RECT 14.656 52.866 14.76 57.24 ; 
      RECT 14.224 52.866 14.328 57.24 ; 
      RECT 13.792 52.866 13.896 57.24 ; 
      RECT 13.36 52.866 13.464 57.24 ; 
      RECT 12.928 52.866 13.032 57.24 ; 
      RECT 12.496 52.866 12.6 57.24 ; 
      RECT 12.064 52.866 12.168 57.24 ; 
      RECT 11.632 52.866 11.736 57.24 ; 
      RECT 11.2 52.866 11.304 57.24 ; 
      RECT 10.768 52.866 10.872 57.24 ; 
      RECT 10.336 52.866 10.44 57.24 ; 
      RECT 9.904 52.866 10.008 57.24 ; 
      RECT 9.472 52.866 9.576 57.24 ; 
      RECT 9.04 52.866 9.144 57.24 ; 
      RECT 8.608 52.866 8.712 57.24 ; 
      RECT 8.176 52.866 8.28 57.24 ; 
      RECT 7.744 52.866 7.848 57.24 ; 
      RECT 7.312 52.866 7.416 57.24 ; 
      RECT 6.88 52.866 6.984 57.24 ; 
      RECT 6.448 52.866 6.552 57.24 ; 
      RECT 6.016 52.866 6.12 57.24 ; 
      RECT 5.584 52.866 5.688 57.24 ; 
      RECT 5.152 52.866 5.256 57.24 ; 
      RECT 4.72 52.866 4.824 57.24 ; 
      RECT 4.288 52.866 4.392 57.24 ; 
      RECT 3.856 52.866 3.96 57.24 ; 
      RECT 3.424 52.866 3.528 57.24 ; 
      RECT 2.992 52.866 3.096 57.24 ; 
      RECT 2.56 52.866 2.664 57.24 ; 
      RECT 2.128 52.866 2.232 57.24 ; 
      RECT 1.696 52.866 1.8 57.24 ; 
      RECT 1.264 52.866 1.368 57.24 ; 
      RECT 0.832 52.866 0.936 57.24 ; 
      RECT 0.02 52.866 0.36 57.24 ; 
      RECT 62.212 57.186 62.724 61.56 ; 
      RECT 62.156 59.848 62.724 61.138 ; 
      RECT 61.276 58.756 61.812 61.56 ; 
      RECT 61.184 60.096 61.812 61.128 ; 
      RECT 61.276 57.186 61.668 61.56 ; 
      RECT 61.276 57.67 61.724 58.628 ; 
      RECT 61.276 57.186 61.812 57.542 ; 
      RECT 60.376 58.988 60.912 61.56 ; 
      RECT 60.376 57.186 60.768 61.56 ; 
      RECT 58.708 57.186 59.04 61.56 ; 
      RECT 58.708 57.54 59.096 61.282 ; 
      RECT 121.072 57.186 121.412 61.56 ; 
      RECT 120.496 57.186 120.6 61.56 ; 
      RECT 120.064 57.186 120.168 61.56 ; 
      RECT 119.632 57.186 119.736 61.56 ; 
      RECT 119.2 57.186 119.304 61.56 ; 
      RECT 118.768 57.186 118.872 61.56 ; 
      RECT 118.336 57.186 118.44 61.56 ; 
      RECT 117.904 57.186 118.008 61.56 ; 
      RECT 117.472 57.186 117.576 61.56 ; 
      RECT 117.04 57.186 117.144 61.56 ; 
      RECT 116.608 57.186 116.712 61.56 ; 
      RECT 116.176 57.186 116.28 61.56 ; 
      RECT 115.744 57.186 115.848 61.56 ; 
      RECT 115.312 57.186 115.416 61.56 ; 
      RECT 114.88 57.186 114.984 61.56 ; 
      RECT 114.448 57.186 114.552 61.56 ; 
      RECT 114.016 57.186 114.12 61.56 ; 
      RECT 113.584 57.186 113.688 61.56 ; 
      RECT 113.152 57.186 113.256 61.56 ; 
      RECT 112.72 57.186 112.824 61.56 ; 
      RECT 112.288 57.186 112.392 61.56 ; 
      RECT 111.856 57.186 111.96 61.56 ; 
      RECT 111.424 57.186 111.528 61.56 ; 
      RECT 110.992 57.186 111.096 61.56 ; 
      RECT 110.56 57.186 110.664 61.56 ; 
      RECT 110.128 57.186 110.232 61.56 ; 
      RECT 109.696 57.186 109.8 61.56 ; 
      RECT 109.264 57.186 109.368 61.56 ; 
      RECT 108.832 57.186 108.936 61.56 ; 
      RECT 108.4 57.186 108.504 61.56 ; 
      RECT 107.968 57.186 108.072 61.56 ; 
      RECT 107.536 57.186 107.64 61.56 ; 
      RECT 107.104 57.186 107.208 61.56 ; 
      RECT 106.672 57.186 106.776 61.56 ; 
      RECT 106.24 57.186 106.344 61.56 ; 
      RECT 105.808 57.186 105.912 61.56 ; 
      RECT 105.376 57.186 105.48 61.56 ; 
      RECT 104.944 57.186 105.048 61.56 ; 
      RECT 104.512 57.186 104.616 61.56 ; 
      RECT 104.08 57.186 104.184 61.56 ; 
      RECT 103.648 57.186 103.752 61.56 ; 
      RECT 103.216 57.186 103.32 61.56 ; 
      RECT 102.784 57.186 102.888 61.56 ; 
      RECT 102.352 57.186 102.456 61.56 ; 
      RECT 101.92 57.186 102.024 61.56 ; 
      RECT 101.488 57.186 101.592 61.56 ; 
      RECT 101.056 57.186 101.16 61.56 ; 
      RECT 100.624 57.186 100.728 61.56 ; 
      RECT 100.192 57.186 100.296 61.56 ; 
      RECT 99.76 57.186 99.864 61.56 ; 
      RECT 99.328 57.186 99.432 61.56 ; 
      RECT 98.896 57.186 99 61.56 ; 
      RECT 98.464 57.186 98.568 61.56 ; 
      RECT 98.032 57.186 98.136 61.56 ; 
      RECT 97.6 57.186 97.704 61.56 ; 
      RECT 97.168 57.186 97.272 61.56 ; 
      RECT 96.736 57.186 96.84 61.56 ; 
      RECT 96.304 57.186 96.408 61.56 ; 
      RECT 95.872 57.186 95.976 61.56 ; 
      RECT 95.44 57.186 95.544 61.56 ; 
      RECT 95.008 57.186 95.112 61.56 ; 
      RECT 94.576 57.186 94.68 61.56 ; 
      RECT 94.144 57.186 94.248 61.56 ; 
      RECT 93.712 57.186 93.816 61.56 ; 
      RECT 93.28 57.186 93.384 61.56 ; 
      RECT 92.848 57.186 92.952 61.56 ; 
      RECT 92.416 57.186 92.52 61.56 ; 
      RECT 91.984 57.186 92.088 61.56 ; 
      RECT 91.552 57.186 91.656 61.56 ; 
      RECT 91.12 57.186 91.224 61.56 ; 
      RECT 90.688 57.186 90.792 61.56 ; 
      RECT 90.256 57.186 90.36 61.56 ; 
      RECT 89.824 57.186 89.928 61.56 ; 
      RECT 89.392 57.186 89.496 61.56 ; 
      RECT 88.96 57.186 89.064 61.56 ; 
      RECT 88.528 57.186 88.632 61.56 ; 
      RECT 88.096 57.186 88.2 61.56 ; 
      RECT 87.664 57.186 87.768 61.56 ; 
      RECT 87.232 57.186 87.336 61.56 ; 
      RECT 86.8 57.186 86.904 61.56 ; 
      RECT 86.368 57.186 86.472 61.56 ; 
      RECT 85.936 57.186 86.04 61.56 ; 
      RECT 85.504 57.186 85.608 61.56 ; 
      RECT 85.072 57.186 85.176 61.56 ; 
      RECT 84.64 57.186 84.744 61.56 ; 
      RECT 84.208 57.186 84.312 61.56 ; 
      RECT 83.776 57.186 83.88 61.56 ; 
      RECT 83.344 57.186 83.448 61.56 ; 
      RECT 82.912 57.186 83.016 61.56 ; 
      RECT 82.48 57.186 82.584 61.56 ; 
      RECT 82.048 57.186 82.152 61.56 ; 
      RECT 81.616 57.186 81.72 61.56 ; 
      RECT 81.184 57.186 81.288 61.56 ; 
      RECT 80.752 57.186 80.856 61.56 ; 
      RECT 80.32 57.186 80.424 61.56 ; 
      RECT 79.888 57.186 79.992 61.56 ; 
      RECT 79.456 57.186 79.56 61.56 ; 
      RECT 79.024 57.186 79.128 61.56 ; 
      RECT 78.592 57.186 78.696 61.56 ; 
      RECT 78.16 57.186 78.264 61.56 ; 
      RECT 77.728 57.186 77.832 61.56 ; 
      RECT 77.296 57.186 77.4 61.56 ; 
      RECT 76.864 57.186 76.968 61.56 ; 
      RECT 76.432 57.186 76.536 61.56 ; 
      RECT 76 57.186 76.104 61.56 ; 
      RECT 75.568 57.186 75.672 61.56 ; 
      RECT 75.136 57.186 75.24 61.56 ; 
      RECT 74.704 57.186 74.808 61.56 ; 
      RECT 74.272 57.186 74.376 61.56 ; 
      RECT 73.84 57.186 73.944 61.56 ; 
      RECT 73.408 57.186 73.512 61.56 ; 
      RECT 72.976 57.186 73.08 61.56 ; 
      RECT 72.544 57.186 72.648 61.56 ; 
      RECT 72.112 57.186 72.216 61.56 ; 
      RECT 71.68 57.186 71.784 61.56 ; 
      RECT 71.248 57.186 71.352 61.56 ; 
      RECT 70.816 57.186 70.92 61.56 ; 
      RECT 70.384 57.186 70.488 61.56 ; 
      RECT 69.952 57.186 70.056 61.56 ; 
      RECT 69.52 57.186 69.624 61.56 ; 
      RECT 69.088 57.186 69.192 61.56 ; 
      RECT 68.656 57.186 68.76 61.56 ; 
      RECT 68.224 57.186 68.328 61.56 ; 
      RECT 67.792 57.186 67.896 61.56 ; 
      RECT 67.36 57.186 67.464 61.56 ; 
      RECT 66.928 57.186 67.032 61.56 ; 
      RECT 66.496 57.186 66.6 61.56 ; 
      RECT 66.064 57.186 66.168 61.56 ; 
      RECT 65.632 57.186 65.736 61.56 ; 
      RECT 65.2 57.186 65.304 61.56 ; 
      RECT 64.348 57.186 64.656 61.56 ; 
      RECT 56.776 57.186 57.084 61.56 ; 
      RECT 56.128 57.186 56.232 61.56 ; 
      RECT 55.696 57.186 55.8 61.56 ; 
      RECT 55.264 57.186 55.368 61.56 ; 
      RECT 54.832 57.186 54.936 61.56 ; 
      RECT 54.4 57.186 54.504 61.56 ; 
      RECT 53.968 57.186 54.072 61.56 ; 
      RECT 53.536 57.186 53.64 61.56 ; 
      RECT 53.104 57.186 53.208 61.56 ; 
      RECT 52.672 57.186 52.776 61.56 ; 
      RECT 52.24 57.186 52.344 61.56 ; 
      RECT 51.808 57.186 51.912 61.56 ; 
      RECT 51.376 57.186 51.48 61.56 ; 
      RECT 50.944 57.186 51.048 61.56 ; 
      RECT 50.512 57.186 50.616 61.56 ; 
      RECT 50.08 57.186 50.184 61.56 ; 
      RECT 49.648 57.186 49.752 61.56 ; 
      RECT 49.216 57.186 49.32 61.56 ; 
      RECT 48.784 57.186 48.888 61.56 ; 
      RECT 48.352 57.186 48.456 61.56 ; 
      RECT 47.92 57.186 48.024 61.56 ; 
      RECT 47.488 57.186 47.592 61.56 ; 
      RECT 47.056 57.186 47.16 61.56 ; 
      RECT 46.624 57.186 46.728 61.56 ; 
      RECT 46.192 57.186 46.296 61.56 ; 
      RECT 45.76 57.186 45.864 61.56 ; 
      RECT 45.328 57.186 45.432 61.56 ; 
      RECT 44.896 57.186 45 61.56 ; 
      RECT 44.464 57.186 44.568 61.56 ; 
      RECT 44.032 57.186 44.136 61.56 ; 
      RECT 43.6 57.186 43.704 61.56 ; 
      RECT 43.168 57.186 43.272 61.56 ; 
      RECT 42.736 57.186 42.84 61.56 ; 
      RECT 42.304 57.186 42.408 61.56 ; 
      RECT 41.872 57.186 41.976 61.56 ; 
      RECT 41.44 57.186 41.544 61.56 ; 
      RECT 41.008 57.186 41.112 61.56 ; 
      RECT 40.576 57.186 40.68 61.56 ; 
      RECT 40.144 57.186 40.248 61.56 ; 
      RECT 39.712 57.186 39.816 61.56 ; 
      RECT 39.28 57.186 39.384 61.56 ; 
      RECT 38.848 57.186 38.952 61.56 ; 
      RECT 38.416 57.186 38.52 61.56 ; 
      RECT 37.984 57.186 38.088 61.56 ; 
      RECT 37.552 57.186 37.656 61.56 ; 
      RECT 37.12 57.186 37.224 61.56 ; 
      RECT 36.688 57.186 36.792 61.56 ; 
      RECT 36.256 57.186 36.36 61.56 ; 
      RECT 35.824 57.186 35.928 61.56 ; 
      RECT 35.392 57.186 35.496 61.56 ; 
      RECT 34.96 57.186 35.064 61.56 ; 
      RECT 34.528 57.186 34.632 61.56 ; 
      RECT 34.096 57.186 34.2 61.56 ; 
      RECT 33.664 57.186 33.768 61.56 ; 
      RECT 33.232 57.186 33.336 61.56 ; 
      RECT 32.8 57.186 32.904 61.56 ; 
      RECT 32.368 57.186 32.472 61.56 ; 
      RECT 31.936 57.186 32.04 61.56 ; 
      RECT 31.504 57.186 31.608 61.56 ; 
      RECT 31.072 57.186 31.176 61.56 ; 
      RECT 30.64 57.186 30.744 61.56 ; 
      RECT 30.208 57.186 30.312 61.56 ; 
      RECT 29.776 57.186 29.88 61.56 ; 
      RECT 29.344 57.186 29.448 61.56 ; 
      RECT 28.912 57.186 29.016 61.56 ; 
      RECT 28.48 57.186 28.584 61.56 ; 
      RECT 28.048 57.186 28.152 61.56 ; 
      RECT 27.616 57.186 27.72 61.56 ; 
      RECT 27.184 57.186 27.288 61.56 ; 
      RECT 26.752 57.186 26.856 61.56 ; 
      RECT 26.32 57.186 26.424 61.56 ; 
      RECT 25.888 57.186 25.992 61.56 ; 
      RECT 25.456 57.186 25.56 61.56 ; 
      RECT 25.024 57.186 25.128 61.56 ; 
      RECT 24.592 57.186 24.696 61.56 ; 
      RECT 24.16 57.186 24.264 61.56 ; 
      RECT 23.728 57.186 23.832 61.56 ; 
      RECT 23.296 57.186 23.4 61.56 ; 
      RECT 22.864 57.186 22.968 61.56 ; 
      RECT 22.432 57.186 22.536 61.56 ; 
      RECT 22 57.186 22.104 61.56 ; 
      RECT 21.568 57.186 21.672 61.56 ; 
      RECT 21.136 57.186 21.24 61.56 ; 
      RECT 20.704 57.186 20.808 61.56 ; 
      RECT 20.272 57.186 20.376 61.56 ; 
      RECT 19.84 57.186 19.944 61.56 ; 
      RECT 19.408 57.186 19.512 61.56 ; 
      RECT 18.976 57.186 19.08 61.56 ; 
      RECT 18.544 57.186 18.648 61.56 ; 
      RECT 18.112 57.186 18.216 61.56 ; 
      RECT 17.68 57.186 17.784 61.56 ; 
      RECT 17.248 57.186 17.352 61.56 ; 
      RECT 16.816 57.186 16.92 61.56 ; 
      RECT 16.384 57.186 16.488 61.56 ; 
      RECT 15.952 57.186 16.056 61.56 ; 
      RECT 15.52 57.186 15.624 61.56 ; 
      RECT 15.088 57.186 15.192 61.56 ; 
      RECT 14.656 57.186 14.76 61.56 ; 
      RECT 14.224 57.186 14.328 61.56 ; 
      RECT 13.792 57.186 13.896 61.56 ; 
      RECT 13.36 57.186 13.464 61.56 ; 
      RECT 12.928 57.186 13.032 61.56 ; 
      RECT 12.496 57.186 12.6 61.56 ; 
      RECT 12.064 57.186 12.168 61.56 ; 
      RECT 11.632 57.186 11.736 61.56 ; 
      RECT 11.2 57.186 11.304 61.56 ; 
      RECT 10.768 57.186 10.872 61.56 ; 
      RECT 10.336 57.186 10.44 61.56 ; 
      RECT 9.904 57.186 10.008 61.56 ; 
      RECT 9.472 57.186 9.576 61.56 ; 
      RECT 9.04 57.186 9.144 61.56 ; 
      RECT 8.608 57.186 8.712 61.56 ; 
      RECT 8.176 57.186 8.28 61.56 ; 
      RECT 7.744 57.186 7.848 61.56 ; 
      RECT 7.312 57.186 7.416 61.56 ; 
      RECT 6.88 57.186 6.984 61.56 ; 
      RECT 6.448 57.186 6.552 61.56 ; 
      RECT 6.016 57.186 6.12 61.56 ; 
      RECT 5.584 57.186 5.688 61.56 ; 
      RECT 5.152 57.186 5.256 61.56 ; 
      RECT 4.72 57.186 4.824 61.56 ; 
      RECT 4.288 57.186 4.392 61.56 ; 
      RECT 3.856 57.186 3.96 61.56 ; 
      RECT 3.424 57.186 3.528 61.56 ; 
      RECT 2.992 57.186 3.096 61.56 ; 
      RECT 2.56 57.186 2.664 61.56 ; 
      RECT 2.128 57.186 2.232 61.56 ; 
      RECT 1.696 57.186 1.8 61.56 ; 
      RECT 1.264 57.186 1.368 61.56 ; 
      RECT 0.832 57.186 0.936 61.56 ; 
      RECT 0.02 57.186 0.36 61.56 ; 
      RECT 62.212 61.506 62.724 65.88 ; 
      RECT 62.156 64.168 62.724 65.458 ; 
      RECT 61.276 63.076 61.812 65.88 ; 
      RECT 61.184 64.416 61.812 65.448 ; 
      RECT 61.276 61.506 61.668 65.88 ; 
      RECT 61.276 61.99 61.724 62.948 ; 
      RECT 61.276 61.506 61.812 61.862 ; 
      RECT 60.376 63.308 60.912 65.88 ; 
      RECT 60.376 61.506 60.768 65.88 ; 
      RECT 58.708 61.506 59.04 65.88 ; 
      RECT 58.708 61.86 59.096 65.602 ; 
      RECT 121.072 61.506 121.412 65.88 ; 
      RECT 120.496 61.506 120.6 65.88 ; 
      RECT 120.064 61.506 120.168 65.88 ; 
      RECT 119.632 61.506 119.736 65.88 ; 
      RECT 119.2 61.506 119.304 65.88 ; 
      RECT 118.768 61.506 118.872 65.88 ; 
      RECT 118.336 61.506 118.44 65.88 ; 
      RECT 117.904 61.506 118.008 65.88 ; 
      RECT 117.472 61.506 117.576 65.88 ; 
      RECT 117.04 61.506 117.144 65.88 ; 
      RECT 116.608 61.506 116.712 65.88 ; 
      RECT 116.176 61.506 116.28 65.88 ; 
      RECT 115.744 61.506 115.848 65.88 ; 
      RECT 115.312 61.506 115.416 65.88 ; 
      RECT 114.88 61.506 114.984 65.88 ; 
      RECT 114.448 61.506 114.552 65.88 ; 
      RECT 114.016 61.506 114.12 65.88 ; 
      RECT 113.584 61.506 113.688 65.88 ; 
      RECT 113.152 61.506 113.256 65.88 ; 
      RECT 112.72 61.506 112.824 65.88 ; 
      RECT 112.288 61.506 112.392 65.88 ; 
      RECT 111.856 61.506 111.96 65.88 ; 
      RECT 111.424 61.506 111.528 65.88 ; 
      RECT 110.992 61.506 111.096 65.88 ; 
      RECT 110.56 61.506 110.664 65.88 ; 
      RECT 110.128 61.506 110.232 65.88 ; 
      RECT 109.696 61.506 109.8 65.88 ; 
      RECT 109.264 61.506 109.368 65.88 ; 
      RECT 108.832 61.506 108.936 65.88 ; 
      RECT 108.4 61.506 108.504 65.88 ; 
      RECT 107.968 61.506 108.072 65.88 ; 
      RECT 107.536 61.506 107.64 65.88 ; 
      RECT 107.104 61.506 107.208 65.88 ; 
      RECT 106.672 61.506 106.776 65.88 ; 
      RECT 106.24 61.506 106.344 65.88 ; 
      RECT 105.808 61.506 105.912 65.88 ; 
      RECT 105.376 61.506 105.48 65.88 ; 
      RECT 104.944 61.506 105.048 65.88 ; 
      RECT 104.512 61.506 104.616 65.88 ; 
      RECT 104.08 61.506 104.184 65.88 ; 
      RECT 103.648 61.506 103.752 65.88 ; 
      RECT 103.216 61.506 103.32 65.88 ; 
      RECT 102.784 61.506 102.888 65.88 ; 
      RECT 102.352 61.506 102.456 65.88 ; 
      RECT 101.92 61.506 102.024 65.88 ; 
      RECT 101.488 61.506 101.592 65.88 ; 
      RECT 101.056 61.506 101.16 65.88 ; 
      RECT 100.624 61.506 100.728 65.88 ; 
      RECT 100.192 61.506 100.296 65.88 ; 
      RECT 99.76 61.506 99.864 65.88 ; 
      RECT 99.328 61.506 99.432 65.88 ; 
      RECT 98.896 61.506 99 65.88 ; 
      RECT 98.464 61.506 98.568 65.88 ; 
      RECT 98.032 61.506 98.136 65.88 ; 
      RECT 97.6 61.506 97.704 65.88 ; 
      RECT 97.168 61.506 97.272 65.88 ; 
      RECT 96.736 61.506 96.84 65.88 ; 
      RECT 96.304 61.506 96.408 65.88 ; 
      RECT 95.872 61.506 95.976 65.88 ; 
      RECT 95.44 61.506 95.544 65.88 ; 
      RECT 95.008 61.506 95.112 65.88 ; 
      RECT 94.576 61.506 94.68 65.88 ; 
      RECT 94.144 61.506 94.248 65.88 ; 
      RECT 93.712 61.506 93.816 65.88 ; 
      RECT 93.28 61.506 93.384 65.88 ; 
      RECT 92.848 61.506 92.952 65.88 ; 
      RECT 92.416 61.506 92.52 65.88 ; 
      RECT 91.984 61.506 92.088 65.88 ; 
      RECT 91.552 61.506 91.656 65.88 ; 
      RECT 91.12 61.506 91.224 65.88 ; 
      RECT 90.688 61.506 90.792 65.88 ; 
      RECT 90.256 61.506 90.36 65.88 ; 
      RECT 89.824 61.506 89.928 65.88 ; 
      RECT 89.392 61.506 89.496 65.88 ; 
      RECT 88.96 61.506 89.064 65.88 ; 
      RECT 88.528 61.506 88.632 65.88 ; 
      RECT 88.096 61.506 88.2 65.88 ; 
      RECT 87.664 61.506 87.768 65.88 ; 
      RECT 87.232 61.506 87.336 65.88 ; 
      RECT 86.8 61.506 86.904 65.88 ; 
      RECT 86.368 61.506 86.472 65.88 ; 
      RECT 85.936 61.506 86.04 65.88 ; 
      RECT 85.504 61.506 85.608 65.88 ; 
      RECT 85.072 61.506 85.176 65.88 ; 
      RECT 84.64 61.506 84.744 65.88 ; 
      RECT 84.208 61.506 84.312 65.88 ; 
      RECT 83.776 61.506 83.88 65.88 ; 
      RECT 83.344 61.506 83.448 65.88 ; 
      RECT 82.912 61.506 83.016 65.88 ; 
      RECT 82.48 61.506 82.584 65.88 ; 
      RECT 82.048 61.506 82.152 65.88 ; 
      RECT 81.616 61.506 81.72 65.88 ; 
      RECT 81.184 61.506 81.288 65.88 ; 
      RECT 80.752 61.506 80.856 65.88 ; 
      RECT 80.32 61.506 80.424 65.88 ; 
      RECT 79.888 61.506 79.992 65.88 ; 
      RECT 79.456 61.506 79.56 65.88 ; 
      RECT 79.024 61.506 79.128 65.88 ; 
      RECT 78.592 61.506 78.696 65.88 ; 
      RECT 78.16 61.506 78.264 65.88 ; 
      RECT 77.728 61.506 77.832 65.88 ; 
      RECT 77.296 61.506 77.4 65.88 ; 
      RECT 76.864 61.506 76.968 65.88 ; 
      RECT 76.432 61.506 76.536 65.88 ; 
      RECT 76 61.506 76.104 65.88 ; 
      RECT 75.568 61.506 75.672 65.88 ; 
      RECT 75.136 61.506 75.24 65.88 ; 
      RECT 74.704 61.506 74.808 65.88 ; 
      RECT 74.272 61.506 74.376 65.88 ; 
      RECT 73.84 61.506 73.944 65.88 ; 
      RECT 73.408 61.506 73.512 65.88 ; 
      RECT 72.976 61.506 73.08 65.88 ; 
      RECT 72.544 61.506 72.648 65.88 ; 
      RECT 72.112 61.506 72.216 65.88 ; 
      RECT 71.68 61.506 71.784 65.88 ; 
      RECT 71.248 61.506 71.352 65.88 ; 
      RECT 70.816 61.506 70.92 65.88 ; 
      RECT 70.384 61.506 70.488 65.88 ; 
      RECT 69.952 61.506 70.056 65.88 ; 
      RECT 69.52 61.506 69.624 65.88 ; 
      RECT 69.088 61.506 69.192 65.88 ; 
      RECT 68.656 61.506 68.76 65.88 ; 
      RECT 68.224 61.506 68.328 65.88 ; 
      RECT 67.792 61.506 67.896 65.88 ; 
      RECT 67.36 61.506 67.464 65.88 ; 
      RECT 66.928 61.506 67.032 65.88 ; 
      RECT 66.496 61.506 66.6 65.88 ; 
      RECT 66.064 61.506 66.168 65.88 ; 
      RECT 65.632 61.506 65.736 65.88 ; 
      RECT 65.2 61.506 65.304 65.88 ; 
      RECT 64.348 61.506 64.656 65.88 ; 
      RECT 56.776 61.506 57.084 65.88 ; 
      RECT 56.128 61.506 56.232 65.88 ; 
      RECT 55.696 61.506 55.8 65.88 ; 
      RECT 55.264 61.506 55.368 65.88 ; 
      RECT 54.832 61.506 54.936 65.88 ; 
      RECT 54.4 61.506 54.504 65.88 ; 
      RECT 53.968 61.506 54.072 65.88 ; 
      RECT 53.536 61.506 53.64 65.88 ; 
      RECT 53.104 61.506 53.208 65.88 ; 
      RECT 52.672 61.506 52.776 65.88 ; 
      RECT 52.24 61.506 52.344 65.88 ; 
      RECT 51.808 61.506 51.912 65.88 ; 
      RECT 51.376 61.506 51.48 65.88 ; 
      RECT 50.944 61.506 51.048 65.88 ; 
      RECT 50.512 61.506 50.616 65.88 ; 
      RECT 50.08 61.506 50.184 65.88 ; 
      RECT 49.648 61.506 49.752 65.88 ; 
      RECT 49.216 61.506 49.32 65.88 ; 
      RECT 48.784 61.506 48.888 65.88 ; 
      RECT 48.352 61.506 48.456 65.88 ; 
      RECT 47.92 61.506 48.024 65.88 ; 
      RECT 47.488 61.506 47.592 65.88 ; 
      RECT 47.056 61.506 47.16 65.88 ; 
      RECT 46.624 61.506 46.728 65.88 ; 
      RECT 46.192 61.506 46.296 65.88 ; 
      RECT 45.76 61.506 45.864 65.88 ; 
      RECT 45.328 61.506 45.432 65.88 ; 
      RECT 44.896 61.506 45 65.88 ; 
      RECT 44.464 61.506 44.568 65.88 ; 
      RECT 44.032 61.506 44.136 65.88 ; 
      RECT 43.6 61.506 43.704 65.88 ; 
      RECT 43.168 61.506 43.272 65.88 ; 
      RECT 42.736 61.506 42.84 65.88 ; 
      RECT 42.304 61.506 42.408 65.88 ; 
      RECT 41.872 61.506 41.976 65.88 ; 
      RECT 41.44 61.506 41.544 65.88 ; 
      RECT 41.008 61.506 41.112 65.88 ; 
      RECT 40.576 61.506 40.68 65.88 ; 
      RECT 40.144 61.506 40.248 65.88 ; 
      RECT 39.712 61.506 39.816 65.88 ; 
      RECT 39.28 61.506 39.384 65.88 ; 
      RECT 38.848 61.506 38.952 65.88 ; 
      RECT 38.416 61.506 38.52 65.88 ; 
      RECT 37.984 61.506 38.088 65.88 ; 
      RECT 37.552 61.506 37.656 65.88 ; 
      RECT 37.12 61.506 37.224 65.88 ; 
      RECT 36.688 61.506 36.792 65.88 ; 
      RECT 36.256 61.506 36.36 65.88 ; 
      RECT 35.824 61.506 35.928 65.88 ; 
      RECT 35.392 61.506 35.496 65.88 ; 
      RECT 34.96 61.506 35.064 65.88 ; 
      RECT 34.528 61.506 34.632 65.88 ; 
      RECT 34.096 61.506 34.2 65.88 ; 
      RECT 33.664 61.506 33.768 65.88 ; 
      RECT 33.232 61.506 33.336 65.88 ; 
      RECT 32.8 61.506 32.904 65.88 ; 
      RECT 32.368 61.506 32.472 65.88 ; 
      RECT 31.936 61.506 32.04 65.88 ; 
      RECT 31.504 61.506 31.608 65.88 ; 
      RECT 31.072 61.506 31.176 65.88 ; 
      RECT 30.64 61.506 30.744 65.88 ; 
      RECT 30.208 61.506 30.312 65.88 ; 
      RECT 29.776 61.506 29.88 65.88 ; 
      RECT 29.344 61.506 29.448 65.88 ; 
      RECT 28.912 61.506 29.016 65.88 ; 
      RECT 28.48 61.506 28.584 65.88 ; 
      RECT 28.048 61.506 28.152 65.88 ; 
      RECT 27.616 61.506 27.72 65.88 ; 
      RECT 27.184 61.506 27.288 65.88 ; 
      RECT 26.752 61.506 26.856 65.88 ; 
      RECT 26.32 61.506 26.424 65.88 ; 
      RECT 25.888 61.506 25.992 65.88 ; 
      RECT 25.456 61.506 25.56 65.88 ; 
      RECT 25.024 61.506 25.128 65.88 ; 
      RECT 24.592 61.506 24.696 65.88 ; 
      RECT 24.16 61.506 24.264 65.88 ; 
      RECT 23.728 61.506 23.832 65.88 ; 
      RECT 23.296 61.506 23.4 65.88 ; 
      RECT 22.864 61.506 22.968 65.88 ; 
      RECT 22.432 61.506 22.536 65.88 ; 
      RECT 22 61.506 22.104 65.88 ; 
      RECT 21.568 61.506 21.672 65.88 ; 
      RECT 21.136 61.506 21.24 65.88 ; 
      RECT 20.704 61.506 20.808 65.88 ; 
      RECT 20.272 61.506 20.376 65.88 ; 
      RECT 19.84 61.506 19.944 65.88 ; 
      RECT 19.408 61.506 19.512 65.88 ; 
      RECT 18.976 61.506 19.08 65.88 ; 
      RECT 18.544 61.506 18.648 65.88 ; 
      RECT 18.112 61.506 18.216 65.88 ; 
      RECT 17.68 61.506 17.784 65.88 ; 
      RECT 17.248 61.506 17.352 65.88 ; 
      RECT 16.816 61.506 16.92 65.88 ; 
      RECT 16.384 61.506 16.488 65.88 ; 
      RECT 15.952 61.506 16.056 65.88 ; 
      RECT 15.52 61.506 15.624 65.88 ; 
      RECT 15.088 61.506 15.192 65.88 ; 
      RECT 14.656 61.506 14.76 65.88 ; 
      RECT 14.224 61.506 14.328 65.88 ; 
      RECT 13.792 61.506 13.896 65.88 ; 
      RECT 13.36 61.506 13.464 65.88 ; 
      RECT 12.928 61.506 13.032 65.88 ; 
      RECT 12.496 61.506 12.6 65.88 ; 
      RECT 12.064 61.506 12.168 65.88 ; 
      RECT 11.632 61.506 11.736 65.88 ; 
      RECT 11.2 61.506 11.304 65.88 ; 
      RECT 10.768 61.506 10.872 65.88 ; 
      RECT 10.336 61.506 10.44 65.88 ; 
      RECT 9.904 61.506 10.008 65.88 ; 
      RECT 9.472 61.506 9.576 65.88 ; 
      RECT 9.04 61.506 9.144 65.88 ; 
      RECT 8.608 61.506 8.712 65.88 ; 
      RECT 8.176 61.506 8.28 65.88 ; 
      RECT 7.744 61.506 7.848 65.88 ; 
      RECT 7.312 61.506 7.416 65.88 ; 
      RECT 6.88 61.506 6.984 65.88 ; 
      RECT 6.448 61.506 6.552 65.88 ; 
      RECT 6.016 61.506 6.12 65.88 ; 
      RECT 5.584 61.506 5.688 65.88 ; 
      RECT 5.152 61.506 5.256 65.88 ; 
      RECT 4.72 61.506 4.824 65.88 ; 
      RECT 4.288 61.506 4.392 65.88 ; 
      RECT 3.856 61.506 3.96 65.88 ; 
      RECT 3.424 61.506 3.528 65.88 ; 
      RECT 2.992 61.506 3.096 65.88 ; 
      RECT 2.56 61.506 2.664 65.88 ; 
      RECT 2.128 61.506 2.232 65.88 ; 
      RECT 1.696 61.506 1.8 65.88 ; 
      RECT 1.264 61.506 1.368 65.88 ; 
      RECT 0.832 61.506 0.936 65.88 ; 
      RECT 0.02 61.506 0.36 65.88 ; 
      RECT 62.212 65.826 62.724 70.2 ; 
      RECT 62.156 68.488 62.724 69.778 ; 
      RECT 61.276 67.396 61.812 70.2 ; 
      RECT 61.184 68.736 61.812 69.768 ; 
      RECT 61.276 65.826 61.668 70.2 ; 
      RECT 61.276 66.31 61.724 67.268 ; 
      RECT 61.276 65.826 61.812 66.182 ; 
      RECT 60.376 67.628 60.912 70.2 ; 
      RECT 60.376 65.826 60.768 70.2 ; 
      RECT 58.708 65.826 59.04 70.2 ; 
      RECT 58.708 66.18 59.096 69.922 ; 
      RECT 121.072 65.826 121.412 70.2 ; 
      RECT 120.496 65.826 120.6 70.2 ; 
      RECT 120.064 65.826 120.168 70.2 ; 
      RECT 119.632 65.826 119.736 70.2 ; 
      RECT 119.2 65.826 119.304 70.2 ; 
      RECT 118.768 65.826 118.872 70.2 ; 
      RECT 118.336 65.826 118.44 70.2 ; 
      RECT 117.904 65.826 118.008 70.2 ; 
      RECT 117.472 65.826 117.576 70.2 ; 
      RECT 117.04 65.826 117.144 70.2 ; 
      RECT 116.608 65.826 116.712 70.2 ; 
      RECT 116.176 65.826 116.28 70.2 ; 
      RECT 115.744 65.826 115.848 70.2 ; 
      RECT 115.312 65.826 115.416 70.2 ; 
      RECT 114.88 65.826 114.984 70.2 ; 
      RECT 114.448 65.826 114.552 70.2 ; 
      RECT 114.016 65.826 114.12 70.2 ; 
      RECT 113.584 65.826 113.688 70.2 ; 
      RECT 113.152 65.826 113.256 70.2 ; 
      RECT 112.72 65.826 112.824 70.2 ; 
      RECT 112.288 65.826 112.392 70.2 ; 
      RECT 111.856 65.826 111.96 70.2 ; 
      RECT 111.424 65.826 111.528 70.2 ; 
      RECT 110.992 65.826 111.096 70.2 ; 
      RECT 110.56 65.826 110.664 70.2 ; 
      RECT 110.128 65.826 110.232 70.2 ; 
      RECT 109.696 65.826 109.8 70.2 ; 
      RECT 109.264 65.826 109.368 70.2 ; 
      RECT 108.832 65.826 108.936 70.2 ; 
      RECT 108.4 65.826 108.504 70.2 ; 
      RECT 107.968 65.826 108.072 70.2 ; 
      RECT 107.536 65.826 107.64 70.2 ; 
      RECT 107.104 65.826 107.208 70.2 ; 
      RECT 106.672 65.826 106.776 70.2 ; 
      RECT 106.24 65.826 106.344 70.2 ; 
      RECT 105.808 65.826 105.912 70.2 ; 
      RECT 105.376 65.826 105.48 70.2 ; 
      RECT 104.944 65.826 105.048 70.2 ; 
      RECT 104.512 65.826 104.616 70.2 ; 
      RECT 104.08 65.826 104.184 70.2 ; 
      RECT 103.648 65.826 103.752 70.2 ; 
      RECT 103.216 65.826 103.32 70.2 ; 
      RECT 102.784 65.826 102.888 70.2 ; 
      RECT 102.352 65.826 102.456 70.2 ; 
      RECT 101.92 65.826 102.024 70.2 ; 
      RECT 101.488 65.826 101.592 70.2 ; 
      RECT 101.056 65.826 101.16 70.2 ; 
      RECT 100.624 65.826 100.728 70.2 ; 
      RECT 100.192 65.826 100.296 70.2 ; 
      RECT 99.76 65.826 99.864 70.2 ; 
      RECT 99.328 65.826 99.432 70.2 ; 
      RECT 98.896 65.826 99 70.2 ; 
      RECT 98.464 65.826 98.568 70.2 ; 
      RECT 98.032 65.826 98.136 70.2 ; 
      RECT 97.6 65.826 97.704 70.2 ; 
      RECT 97.168 65.826 97.272 70.2 ; 
      RECT 96.736 65.826 96.84 70.2 ; 
      RECT 96.304 65.826 96.408 70.2 ; 
      RECT 95.872 65.826 95.976 70.2 ; 
      RECT 95.44 65.826 95.544 70.2 ; 
      RECT 95.008 65.826 95.112 70.2 ; 
      RECT 94.576 65.826 94.68 70.2 ; 
      RECT 94.144 65.826 94.248 70.2 ; 
      RECT 93.712 65.826 93.816 70.2 ; 
      RECT 93.28 65.826 93.384 70.2 ; 
      RECT 92.848 65.826 92.952 70.2 ; 
      RECT 92.416 65.826 92.52 70.2 ; 
      RECT 91.984 65.826 92.088 70.2 ; 
      RECT 91.552 65.826 91.656 70.2 ; 
      RECT 91.12 65.826 91.224 70.2 ; 
      RECT 90.688 65.826 90.792 70.2 ; 
      RECT 90.256 65.826 90.36 70.2 ; 
      RECT 89.824 65.826 89.928 70.2 ; 
      RECT 89.392 65.826 89.496 70.2 ; 
      RECT 88.96 65.826 89.064 70.2 ; 
      RECT 88.528 65.826 88.632 70.2 ; 
      RECT 88.096 65.826 88.2 70.2 ; 
      RECT 87.664 65.826 87.768 70.2 ; 
      RECT 87.232 65.826 87.336 70.2 ; 
      RECT 86.8 65.826 86.904 70.2 ; 
      RECT 86.368 65.826 86.472 70.2 ; 
      RECT 85.936 65.826 86.04 70.2 ; 
      RECT 85.504 65.826 85.608 70.2 ; 
      RECT 85.072 65.826 85.176 70.2 ; 
      RECT 84.64 65.826 84.744 70.2 ; 
      RECT 84.208 65.826 84.312 70.2 ; 
      RECT 83.776 65.826 83.88 70.2 ; 
      RECT 83.344 65.826 83.448 70.2 ; 
      RECT 82.912 65.826 83.016 70.2 ; 
      RECT 82.48 65.826 82.584 70.2 ; 
      RECT 82.048 65.826 82.152 70.2 ; 
      RECT 81.616 65.826 81.72 70.2 ; 
      RECT 81.184 65.826 81.288 70.2 ; 
      RECT 80.752 65.826 80.856 70.2 ; 
      RECT 80.32 65.826 80.424 70.2 ; 
      RECT 79.888 65.826 79.992 70.2 ; 
      RECT 79.456 65.826 79.56 70.2 ; 
      RECT 79.024 65.826 79.128 70.2 ; 
      RECT 78.592 65.826 78.696 70.2 ; 
      RECT 78.16 65.826 78.264 70.2 ; 
      RECT 77.728 65.826 77.832 70.2 ; 
      RECT 77.296 65.826 77.4 70.2 ; 
      RECT 76.864 65.826 76.968 70.2 ; 
      RECT 76.432 65.826 76.536 70.2 ; 
      RECT 76 65.826 76.104 70.2 ; 
      RECT 75.568 65.826 75.672 70.2 ; 
      RECT 75.136 65.826 75.24 70.2 ; 
      RECT 74.704 65.826 74.808 70.2 ; 
      RECT 74.272 65.826 74.376 70.2 ; 
      RECT 73.84 65.826 73.944 70.2 ; 
      RECT 73.408 65.826 73.512 70.2 ; 
      RECT 72.976 65.826 73.08 70.2 ; 
      RECT 72.544 65.826 72.648 70.2 ; 
      RECT 72.112 65.826 72.216 70.2 ; 
      RECT 71.68 65.826 71.784 70.2 ; 
      RECT 71.248 65.826 71.352 70.2 ; 
      RECT 70.816 65.826 70.92 70.2 ; 
      RECT 70.384 65.826 70.488 70.2 ; 
      RECT 69.952 65.826 70.056 70.2 ; 
      RECT 69.52 65.826 69.624 70.2 ; 
      RECT 69.088 65.826 69.192 70.2 ; 
      RECT 68.656 65.826 68.76 70.2 ; 
      RECT 68.224 65.826 68.328 70.2 ; 
      RECT 67.792 65.826 67.896 70.2 ; 
      RECT 67.36 65.826 67.464 70.2 ; 
      RECT 66.928 65.826 67.032 70.2 ; 
      RECT 66.496 65.826 66.6 70.2 ; 
      RECT 66.064 65.826 66.168 70.2 ; 
      RECT 65.632 65.826 65.736 70.2 ; 
      RECT 65.2 65.826 65.304 70.2 ; 
      RECT 64.348 65.826 64.656 70.2 ; 
      RECT 56.776 65.826 57.084 70.2 ; 
      RECT 56.128 65.826 56.232 70.2 ; 
      RECT 55.696 65.826 55.8 70.2 ; 
      RECT 55.264 65.826 55.368 70.2 ; 
      RECT 54.832 65.826 54.936 70.2 ; 
      RECT 54.4 65.826 54.504 70.2 ; 
      RECT 53.968 65.826 54.072 70.2 ; 
      RECT 53.536 65.826 53.64 70.2 ; 
      RECT 53.104 65.826 53.208 70.2 ; 
      RECT 52.672 65.826 52.776 70.2 ; 
      RECT 52.24 65.826 52.344 70.2 ; 
      RECT 51.808 65.826 51.912 70.2 ; 
      RECT 51.376 65.826 51.48 70.2 ; 
      RECT 50.944 65.826 51.048 70.2 ; 
      RECT 50.512 65.826 50.616 70.2 ; 
      RECT 50.08 65.826 50.184 70.2 ; 
      RECT 49.648 65.826 49.752 70.2 ; 
      RECT 49.216 65.826 49.32 70.2 ; 
      RECT 48.784 65.826 48.888 70.2 ; 
      RECT 48.352 65.826 48.456 70.2 ; 
      RECT 47.92 65.826 48.024 70.2 ; 
      RECT 47.488 65.826 47.592 70.2 ; 
      RECT 47.056 65.826 47.16 70.2 ; 
      RECT 46.624 65.826 46.728 70.2 ; 
      RECT 46.192 65.826 46.296 70.2 ; 
      RECT 45.76 65.826 45.864 70.2 ; 
      RECT 45.328 65.826 45.432 70.2 ; 
      RECT 44.896 65.826 45 70.2 ; 
      RECT 44.464 65.826 44.568 70.2 ; 
      RECT 44.032 65.826 44.136 70.2 ; 
      RECT 43.6 65.826 43.704 70.2 ; 
      RECT 43.168 65.826 43.272 70.2 ; 
      RECT 42.736 65.826 42.84 70.2 ; 
      RECT 42.304 65.826 42.408 70.2 ; 
      RECT 41.872 65.826 41.976 70.2 ; 
      RECT 41.44 65.826 41.544 70.2 ; 
      RECT 41.008 65.826 41.112 70.2 ; 
      RECT 40.576 65.826 40.68 70.2 ; 
      RECT 40.144 65.826 40.248 70.2 ; 
      RECT 39.712 65.826 39.816 70.2 ; 
      RECT 39.28 65.826 39.384 70.2 ; 
      RECT 38.848 65.826 38.952 70.2 ; 
      RECT 38.416 65.826 38.52 70.2 ; 
      RECT 37.984 65.826 38.088 70.2 ; 
      RECT 37.552 65.826 37.656 70.2 ; 
      RECT 37.12 65.826 37.224 70.2 ; 
      RECT 36.688 65.826 36.792 70.2 ; 
      RECT 36.256 65.826 36.36 70.2 ; 
      RECT 35.824 65.826 35.928 70.2 ; 
      RECT 35.392 65.826 35.496 70.2 ; 
      RECT 34.96 65.826 35.064 70.2 ; 
      RECT 34.528 65.826 34.632 70.2 ; 
      RECT 34.096 65.826 34.2 70.2 ; 
      RECT 33.664 65.826 33.768 70.2 ; 
      RECT 33.232 65.826 33.336 70.2 ; 
      RECT 32.8 65.826 32.904 70.2 ; 
      RECT 32.368 65.826 32.472 70.2 ; 
      RECT 31.936 65.826 32.04 70.2 ; 
      RECT 31.504 65.826 31.608 70.2 ; 
      RECT 31.072 65.826 31.176 70.2 ; 
      RECT 30.64 65.826 30.744 70.2 ; 
      RECT 30.208 65.826 30.312 70.2 ; 
      RECT 29.776 65.826 29.88 70.2 ; 
      RECT 29.344 65.826 29.448 70.2 ; 
      RECT 28.912 65.826 29.016 70.2 ; 
      RECT 28.48 65.826 28.584 70.2 ; 
      RECT 28.048 65.826 28.152 70.2 ; 
      RECT 27.616 65.826 27.72 70.2 ; 
      RECT 27.184 65.826 27.288 70.2 ; 
      RECT 26.752 65.826 26.856 70.2 ; 
      RECT 26.32 65.826 26.424 70.2 ; 
      RECT 25.888 65.826 25.992 70.2 ; 
      RECT 25.456 65.826 25.56 70.2 ; 
      RECT 25.024 65.826 25.128 70.2 ; 
      RECT 24.592 65.826 24.696 70.2 ; 
      RECT 24.16 65.826 24.264 70.2 ; 
      RECT 23.728 65.826 23.832 70.2 ; 
      RECT 23.296 65.826 23.4 70.2 ; 
      RECT 22.864 65.826 22.968 70.2 ; 
      RECT 22.432 65.826 22.536 70.2 ; 
      RECT 22 65.826 22.104 70.2 ; 
      RECT 21.568 65.826 21.672 70.2 ; 
      RECT 21.136 65.826 21.24 70.2 ; 
      RECT 20.704 65.826 20.808 70.2 ; 
      RECT 20.272 65.826 20.376 70.2 ; 
      RECT 19.84 65.826 19.944 70.2 ; 
      RECT 19.408 65.826 19.512 70.2 ; 
      RECT 18.976 65.826 19.08 70.2 ; 
      RECT 18.544 65.826 18.648 70.2 ; 
      RECT 18.112 65.826 18.216 70.2 ; 
      RECT 17.68 65.826 17.784 70.2 ; 
      RECT 17.248 65.826 17.352 70.2 ; 
      RECT 16.816 65.826 16.92 70.2 ; 
      RECT 16.384 65.826 16.488 70.2 ; 
      RECT 15.952 65.826 16.056 70.2 ; 
      RECT 15.52 65.826 15.624 70.2 ; 
      RECT 15.088 65.826 15.192 70.2 ; 
      RECT 14.656 65.826 14.76 70.2 ; 
      RECT 14.224 65.826 14.328 70.2 ; 
      RECT 13.792 65.826 13.896 70.2 ; 
      RECT 13.36 65.826 13.464 70.2 ; 
      RECT 12.928 65.826 13.032 70.2 ; 
      RECT 12.496 65.826 12.6 70.2 ; 
      RECT 12.064 65.826 12.168 70.2 ; 
      RECT 11.632 65.826 11.736 70.2 ; 
      RECT 11.2 65.826 11.304 70.2 ; 
      RECT 10.768 65.826 10.872 70.2 ; 
      RECT 10.336 65.826 10.44 70.2 ; 
      RECT 9.904 65.826 10.008 70.2 ; 
      RECT 9.472 65.826 9.576 70.2 ; 
      RECT 9.04 65.826 9.144 70.2 ; 
      RECT 8.608 65.826 8.712 70.2 ; 
      RECT 8.176 65.826 8.28 70.2 ; 
      RECT 7.744 65.826 7.848 70.2 ; 
      RECT 7.312 65.826 7.416 70.2 ; 
      RECT 6.88 65.826 6.984 70.2 ; 
      RECT 6.448 65.826 6.552 70.2 ; 
      RECT 6.016 65.826 6.12 70.2 ; 
      RECT 5.584 65.826 5.688 70.2 ; 
      RECT 5.152 65.826 5.256 70.2 ; 
      RECT 4.72 65.826 4.824 70.2 ; 
      RECT 4.288 65.826 4.392 70.2 ; 
      RECT 3.856 65.826 3.96 70.2 ; 
      RECT 3.424 65.826 3.528 70.2 ; 
      RECT 2.992 65.826 3.096 70.2 ; 
      RECT 2.56 65.826 2.664 70.2 ; 
      RECT 2.128 65.826 2.232 70.2 ; 
      RECT 1.696 65.826 1.8 70.2 ; 
      RECT 1.264 65.826 1.368 70.2 ; 
      RECT 0.832 65.826 0.936 70.2 ; 
      RECT 0.02 65.826 0.36 70.2 ; 
      RECT 62.212 70.146 62.724 74.52 ; 
      RECT 62.156 72.808 62.724 74.098 ; 
      RECT 61.276 71.716 61.812 74.52 ; 
      RECT 61.184 73.056 61.812 74.088 ; 
      RECT 61.276 70.146 61.668 74.52 ; 
      RECT 61.276 70.63 61.724 71.588 ; 
      RECT 61.276 70.146 61.812 70.502 ; 
      RECT 60.376 71.948 60.912 74.52 ; 
      RECT 60.376 70.146 60.768 74.52 ; 
      RECT 58.708 70.146 59.04 74.52 ; 
      RECT 58.708 70.5 59.096 74.242 ; 
      RECT 121.072 70.146 121.412 74.52 ; 
      RECT 120.496 70.146 120.6 74.52 ; 
      RECT 120.064 70.146 120.168 74.52 ; 
      RECT 119.632 70.146 119.736 74.52 ; 
      RECT 119.2 70.146 119.304 74.52 ; 
      RECT 118.768 70.146 118.872 74.52 ; 
      RECT 118.336 70.146 118.44 74.52 ; 
      RECT 117.904 70.146 118.008 74.52 ; 
      RECT 117.472 70.146 117.576 74.52 ; 
      RECT 117.04 70.146 117.144 74.52 ; 
      RECT 116.608 70.146 116.712 74.52 ; 
      RECT 116.176 70.146 116.28 74.52 ; 
      RECT 115.744 70.146 115.848 74.52 ; 
      RECT 115.312 70.146 115.416 74.52 ; 
      RECT 114.88 70.146 114.984 74.52 ; 
      RECT 114.448 70.146 114.552 74.52 ; 
      RECT 114.016 70.146 114.12 74.52 ; 
      RECT 113.584 70.146 113.688 74.52 ; 
      RECT 113.152 70.146 113.256 74.52 ; 
      RECT 112.72 70.146 112.824 74.52 ; 
      RECT 112.288 70.146 112.392 74.52 ; 
      RECT 111.856 70.146 111.96 74.52 ; 
      RECT 111.424 70.146 111.528 74.52 ; 
      RECT 110.992 70.146 111.096 74.52 ; 
      RECT 110.56 70.146 110.664 74.52 ; 
      RECT 110.128 70.146 110.232 74.52 ; 
      RECT 109.696 70.146 109.8 74.52 ; 
      RECT 109.264 70.146 109.368 74.52 ; 
      RECT 108.832 70.146 108.936 74.52 ; 
      RECT 108.4 70.146 108.504 74.52 ; 
      RECT 107.968 70.146 108.072 74.52 ; 
      RECT 107.536 70.146 107.64 74.52 ; 
      RECT 107.104 70.146 107.208 74.52 ; 
      RECT 106.672 70.146 106.776 74.52 ; 
      RECT 106.24 70.146 106.344 74.52 ; 
      RECT 105.808 70.146 105.912 74.52 ; 
      RECT 105.376 70.146 105.48 74.52 ; 
      RECT 104.944 70.146 105.048 74.52 ; 
      RECT 104.512 70.146 104.616 74.52 ; 
      RECT 104.08 70.146 104.184 74.52 ; 
      RECT 103.648 70.146 103.752 74.52 ; 
      RECT 103.216 70.146 103.32 74.52 ; 
      RECT 102.784 70.146 102.888 74.52 ; 
      RECT 102.352 70.146 102.456 74.52 ; 
      RECT 101.92 70.146 102.024 74.52 ; 
      RECT 101.488 70.146 101.592 74.52 ; 
      RECT 101.056 70.146 101.16 74.52 ; 
      RECT 100.624 70.146 100.728 74.52 ; 
      RECT 100.192 70.146 100.296 74.52 ; 
      RECT 99.76 70.146 99.864 74.52 ; 
      RECT 99.328 70.146 99.432 74.52 ; 
      RECT 98.896 70.146 99 74.52 ; 
      RECT 98.464 70.146 98.568 74.52 ; 
      RECT 98.032 70.146 98.136 74.52 ; 
      RECT 97.6 70.146 97.704 74.52 ; 
      RECT 97.168 70.146 97.272 74.52 ; 
      RECT 96.736 70.146 96.84 74.52 ; 
      RECT 96.304 70.146 96.408 74.52 ; 
      RECT 95.872 70.146 95.976 74.52 ; 
      RECT 95.44 70.146 95.544 74.52 ; 
      RECT 95.008 70.146 95.112 74.52 ; 
      RECT 94.576 70.146 94.68 74.52 ; 
      RECT 94.144 70.146 94.248 74.52 ; 
      RECT 93.712 70.146 93.816 74.52 ; 
      RECT 93.28 70.146 93.384 74.52 ; 
      RECT 92.848 70.146 92.952 74.52 ; 
      RECT 92.416 70.146 92.52 74.52 ; 
      RECT 91.984 70.146 92.088 74.52 ; 
      RECT 91.552 70.146 91.656 74.52 ; 
      RECT 91.12 70.146 91.224 74.52 ; 
      RECT 90.688 70.146 90.792 74.52 ; 
      RECT 90.256 70.146 90.36 74.52 ; 
      RECT 89.824 70.146 89.928 74.52 ; 
      RECT 89.392 70.146 89.496 74.52 ; 
      RECT 88.96 70.146 89.064 74.52 ; 
      RECT 88.528 70.146 88.632 74.52 ; 
      RECT 88.096 70.146 88.2 74.52 ; 
      RECT 87.664 70.146 87.768 74.52 ; 
      RECT 87.232 70.146 87.336 74.52 ; 
      RECT 86.8 70.146 86.904 74.52 ; 
      RECT 86.368 70.146 86.472 74.52 ; 
      RECT 85.936 70.146 86.04 74.52 ; 
      RECT 85.504 70.146 85.608 74.52 ; 
      RECT 85.072 70.146 85.176 74.52 ; 
      RECT 84.64 70.146 84.744 74.52 ; 
      RECT 84.208 70.146 84.312 74.52 ; 
      RECT 83.776 70.146 83.88 74.52 ; 
      RECT 83.344 70.146 83.448 74.52 ; 
      RECT 82.912 70.146 83.016 74.52 ; 
      RECT 82.48 70.146 82.584 74.52 ; 
      RECT 82.048 70.146 82.152 74.52 ; 
      RECT 81.616 70.146 81.72 74.52 ; 
      RECT 81.184 70.146 81.288 74.52 ; 
      RECT 80.752 70.146 80.856 74.52 ; 
      RECT 80.32 70.146 80.424 74.52 ; 
      RECT 79.888 70.146 79.992 74.52 ; 
      RECT 79.456 70.146 79.56 74.52 ; 
      RECT 79.024 70.146 79.128 74.52 ; 
      RECT 78.592 70.146 78.696 74.52 ; 
      RECT 78.16 70.146 78.264 74.52 ; 
      RECT 77.728 70.146 77.832 74.52 ; 
      RECT 77.296 70.146 77.4 74.52 ; 
      RECT 76.864 70.146 76.968 74.52 ; 
      RECT 76.432 70.146 76.536 74.52 ; 
      RECT 76 70.146 76.104 74.52 ; 
      RECT 75.568 70.146 75.672 74.52 ; 
      RECT 75.136 70.146 75.24 74.52 ; 
      RECT 74.704 70.146 74.808 74.52 ; 
      RECT 74.272 70.146 74.376 74.52 ; 
      RECT 73.84 70.146 73.944 74.52 ; 
      RECT 73.408 70.146 73.512 74.52 ; 
      RECT 72.976 70.146 73.08 74.52 ; 
      RECT 72.544 70.146 72.648 74.52 ; 
      RECT 72.112 70.146 72.216 74.52 ; 
      RECT 71.68 70.146 71.784 74.52 ; 
      RECT 71.248 70.146 71.352 74.52 ; 
      RECT 70.816 70.146 70.92 74.52 ; 
      RECT 70.384 70.146 70.488 74.52 ; 
      RECT 69.952 70.146 70.056 74.52 ; 
      RECT 69.52 70.146 69.624 74.52 ; 
      RECT 69.088 70.146 69.192 74.52 ; 
      RECT 68.656 70.146 68.76 74.52 ; 
      RECT 68.224 70.146 68.328 74.52 ; 
      RECT 67.792 70.146 67.896 74.52 ; 
      RECT 67.36 70.146 67.464 74.52 ; 
      RECT 66.928 70.146 67.032 74.52 ; 
      RECT 66.496 70.146 66.6 74.52 ; 
      RECT 66.064 70.146 66.168 74.52 ; 
      RECT 65.632 70.146 65.736 74.52 ; 
      RECT 65.2 70.146 65.304 74.52 ; 
      RECT 64.348 70.146 64.656 74.52 ; 
      RECT 56.776 70.146 57.084 74.52 ; 
      RECT 56.128 70.146 56.232 74.52 ; 
      RECT 55.696 70.146 55.8 74.52 ; 
      RECT 55.264 70.146 55.368 74.52 ; 
      RECT 54.832 70.146 54.936 74.52 ; 
      RECT 54.4 70.146 54.504 74.52 ; 
      RECT 53.968 70.146 54.072 74.52 ; 
      RECT 53.536 70.146 53.64 74.52 ; 
      RECT 53.104 70.146 53.208 74.52 ; 
      RECT 52.672 70.146 52.776 74.52 ; 
      RECT 52.24 70.146 52.344 74.52 ; 
      RECT 51.808 70.146 51.912 74.52 ; 
      RECT 51.376 70.146 51.48 74.52 ; 
      RECT 50.944 70.146 51.048 74.52 ; 
      RECT 50.512 70.146 50.616 74.52 ; 
      RECT 50.08 70.146 50.184 74.52 ; 
      RECT 49.648 70.146 49.752 74.52 ; 
      RECT 49.216 70.146 49.32 74.52 ; 
      RECT 48.784 70.146 48.888 74.52 ; 
      RECT 48.352 70.146 48.456 74.52 ; 
      RECT 47.92 70.146 48.024 74.52 ; 
      RECT 47.488 70.146 47.592 74.52 ; 
      RECT 47.056 70.146 47.16 74.52 ; 
      RECT 46.624 70.146 46.728 74.52 ; 
      RECT 46.192 70.146 46.296 74.52 ; 
      RECT 45.76 70.146 45.864 74.52 ; 
      RECT 45.328 70.146 45.432 74.52 ; 
      RECT 44.896 70.146 45 74.52 ; 
      RECT 44.464 70.146 44.568 74.52 ; 
      RECT 44.032 70.146 44.136 74.52 ; 
      RECT 43.6 70.146 43.704 74.52 ; 
      RECT 43.168 70.146 43.272 74.52 ; 
      RECT 42.736 70.146 42.84 74.52 ; 
      RECT 42.304 70.146 42.408 74.52 ; 
      RECT 41.872 70.146 41.976 74.52 ; 
      RECT 41.44 70.146 41.544 74.52 ; 
      RECT 41.008 70.146 41.112 74.52 ; 
      RECT 40.576 70.146 40.68 74.52 ; 
      RECT 40.144 70.146 40.248 74.52 ; 
      RECT 39.712 70.146 39.816 74.52 ; 
      RECT 39.28 70.146 39.384 74.52 ; 
      RECT 38.848 70.146 38.952 74.52 ; 
      RECT 38.416 70.146 38.52 74.52 ; 
      RECT 37.984 70.146 38.088 74.52 ; 
      RECT 37.552 70.146 37.656 74.52 ; 
      RECT 37.12 70.146 37.224 74.52 ; 
      RECT 36.688 70.146 36.792 74.52 ; 
      RECT 36.256 70.146 36.36 74.52 ; 
      RECT 35.824 70.146 35.928 74.52 ; 
      RECT 35.392 70.146 35.496 74.52 ; 
      RECT 34.96 70.146 35.064 74.52 ; 
      RECT 34.528 70.146 34.632 74.52 ; 
      RECT 34.096 70.146 34.2 74.52 ; 
      RECT 33.664 70.146 33.768 74.52 ; 
      RECT 33.232 70.146 33.336 74.52 ; 
      RECT 32.8 70.146 32.904 74.52 ; 
      RECT 32.368 70.146 32.472 74.52 ; 
      RECT 31.936 70.146 32.04 74.52 ; 
      RECT 31.504 70.146 31.608 74.52 ; 
      RECT 31.072 70.146 31.176 74.52 ; 
      RECT 30.64 70.146 30.744 74.52 ; 
      RECT 30.208 70.146 30.312 74.52 ; 
      RECT 29.776 70.146 29.88 74.52 ; 
      RECT 29.344 70.146 29.448 74.52 ; 
      RECT 28.912 70.146 29.016 74.52 ; 
      RECT 28.48 70.146 28.584 74.52 ; 
      RECT 28.048 70.146 28.152 74.52 ; 
      RECT 27.616 70.146 27.72 74.52 ; 
      RECT 27.184 70.146 27.288 74.52 ; 
      RECT 26.752 70.146 26.856 74.52 ; 
      RECT 26.32 70.146 26.424 74.52 ; 
      RECT 25.888 70.146 25.992 74.52 ; 
      RECT 25.456 70.146 25.56 74.52 ; 
      RECT 25.024 70.146 25.128 74.52 ; 
      RECT 24.592 70.146 24.696 74.52 ; 
      RECT 24.16 70.146 24.264 74.52 ; 
      RECT 23.728 70.146 23.832 74.52 ; 
      RECT 23.296 70.146 23.4 74.52 ; 
      RECT 22.864 70.146 22.968 74.52 ; 
      RECT 22.432 70.146 22.536 74.52 ; 
      RECT 22 70.146 22.104 74.52 ; 
      RECT 21.568 70.146 21.672 74.52 ; 
      RECT 21.136 70.146 21.24 74.52 ; 
      RECT 20.704 70.146 20.808 74.52 ; 
      RECT 20.272 70.146 20.376 74.52 ; 
      RECT 19.84 70.146 19.944 74.52 ; 
      RECT 19.408 70.146 19.512 74.52 ; 
      RECT 18.976 70.146 19.08 74.52 ; 
      RECT 18.544 70.146 18.648 74.52 ; 
      RECT 18.112 70.146 18.216 74.52 ; 
      RECT 17.68 70.146 17.784 74.52 ; 
      RECT 17.248 70.146 17.352 74.52 ; 
      RECT 16.816 70.146 16.92 74.52 ; 
      RECT 16.384 70.146 16.488 74.52 ; 
      RECT 15.952 70.146 16.056 74.52 ; 
      RECT 15.52 70.146 15.624 74.52 ; 
      RECT 15.088 70.146 15.192 74.52 ; 
      RECT 14.656 70.146 14.76 74.52 ; 
      RECT 14.224 70.146 14.328 74.52 ; 
      RECT 13.792 70.146 13.896 74.52 ; 
      RECT 13.36 70.146 13.464 74.52 ; 
      RECT 12.928 70.146 13.032 74.52 ; 
      RECT 12.496 70.146 12.6 74.52 ; 
      RECT 12.064 70.146 12.168 74.52 ; 
      RECT 11.632 70.146 11.736 74.52 ; 
      RECT 11.2 70.146 11.304 74.52 ; 
      RECT 10.768 70.146 10.872 74.52 ; 
      RECT 10.336 70.146 10.44 74.52 ; 
      RECT 9.904 70.146 10.008 74.52 ; 
      RECT 9.472 70.146 9.576 74.52 ; 
      RECT 9.04 70.146 9.144 74.52 ; 
      RECT 8.608 70.146 8.712 74.52 ; 
      RECT 8.176 70.146 8.28 74.52 ; 
      RECT 7.744 70.146 7.848 74.52 ; 
      RECT 7.312 70.146 7.416 74.52 ; 
      RECT 6.88 70.146 6.984 74.52 ; 
      RECT 6.448 70.146 6.552 74.52 ; 
      RECT 6.016 70.146 6.12 74.52 ; 
      RECT 5.584 70.146 5.688 74.52 ; 
      RECT 5.152 70.146 5.256 74.52 ; 
      RECT 4.72 70.146 4.824 74.52 ; 
      RECT 4.288 70.146 4.392 74.52 ; 
      RECT 3.856 70.146 3.96 74.52 ; 
      RECT 3.424 70.146 3.528 74.52 ; 
      RECT 2.992 70.146 3.096 74.52 ; 
      RECT 2.56 70.146 2.664 74.52 ; 
      RECT 2.128 70.146 2.232 74.52 ; 
      RECT 1.696 70.146 1.8 74.52 ; 
      RECT 1.264 70.146 1.368 74.52 ; 
      RECT 0.832 70.146 0.936 74.52 ; 
      RECT 0.02 70.146 0.36 74.52 ; 
      RECT 62.212 74.466 62.724 78.84 ; 
      RECT 62.156 77.128 62.724 78.418 ; 
      RECT 61.276 76.036 61.812 78.84 ; 
      RECT 61.184 77.376 61.812 78.408 ; 
      RECT 61.276 74.466 61.668 78.84 ; 
      RECT 61.276 74.95 61.724 75.908 ; 
      RECT 61.276 74.466 61.812 74.822 ; 
      RECT 60.376 76.268 60.912 78.84 ; 
      RECT 60.376 74.466 60.768 78.84 ; 
      RECT 58.708 74.466 59.04 78.84 ; 
      RECT 58.708 74.82 59.096 78.562 ; 
      RECT 121.072 74.466 121.412 78.84 ; 
      RECT 120.496 74.466 120.6 78.84 ; 
      RECT 120.064 74.466 120.168 78.84 ; 
      RECT 119.632 74.466 119.736 78.84 ; 
      RECT 119.2 74.466 119.304 78.84 ; 
      RECT 118.768 74.466 118.872 78.84 ; 
      RECT 118.336 74.466 118.44 78.84 ; 
      RECT 117.904 74.466 118.008 78.84 ; 
      RECT 117.472 74.466 117.576 78.84 ; 
      RECT 117.04 74.466 117.144 78.84 ; 
      RECT 116.608 74.466 116.712 78.84 ; 
      RECT 116.176 74.466 116.28 78.84 ; 
      RECT 115.744 74.466 115.848 78.84 ; 
      RECT 115.312 74.466 115.416 78.84 ; 
      RECT 114.88 74.466 114.984 78.84 ; 
      RECT 114.448 74.466 114.552 78.84 ; 
      RECT 114.016 74.466 114.12 78.84 ; 
      RECT 113.584 74.466 113.688 78.84 ; 
      RECT 113.152 74.466 113.256 78.84 ; 
      RECT 112.72 74.466 112.824 78.84 ; 
      RECT 112.288 74.466 112.392 78.84 ; 
      RECT 111.856 74.466 111.96 78.84 ; 
      RECT 111.424 74.466 111.528 78.84 ; 
      RECT 110.992 74.466 111.096 78.84 ; 
      RECT 110.56 74.466 110.664 78.84 ; 
      RECT 110.128 74.466 110.232 78.84 ; 
      RECT 109.696 74.466 109.8 78.84 ; 
      RECT 109.264 74.466 109.368 78.84 ; 
      RECT 108.832 74.466 108.936 78.84 ; 
      RECT 108.4 74.466 108.504 78.84 ; 
      RECT 107.968 74.466 108.072 78.84 ; 
      RECT 107.536 74.466 107.64 78.84 ; 
      RECT 107.104 74.466 107.208 78.84 ; 
      RECT 106.672 74.466 106.776 78.84 ; 
      RECT 106.24 74.466 106.344 78.84 ; 
      RECT 105.808 74.466 105.912 78.84 ; 
      RECT 105.376 74.466 105.48 78.84 ; 
      RECT 104.944 74.466 105.048 78.84 ; 
      RECT 104.512 74.466 104.616 78.84 ; 
      RECT 104.08 74.466 104.184 78.84 ; 
      RECT 103.648 74.466 103.752 78.84 ; 
      RECT 103.216 74.466 103.32 78.84 ; 
      RECT 102.784 74.466 102.888 78.84 ; 
      RECT 102.352 74.466 102.456 78.84 ; 
      RECT 101.92 74.466 102.024 78.84 ; 
      RECT 101.488 74.466 101.592 78.84 ; 
      RECT 101.056 74.466 101.16 78.84 ; 
      RECT 100.624 74.466 100.728 78.84 ; 
      RECT 100.192 74.466 100.296 78.84 ; 
      RECT 99.76 74.466 99.864 78.84 ; 
      RECT 99.328 74.466 99.432 78.84 ; 
      RECT 98.896 74.466 99 78.84 ; 
      RECT 98.464 74.466 98.568 78.84 ; 
      RECT 98.032 74.466 98.136 78.84 ; 
      RECT 97.6 74.466 97.704 78.84 ; 
      RECT 97.168 74.466 97.272 78.84 ; 
      RECT 96.736 74.466 96.84 78.84 ; 
      RECT 96.304 74.466 96.408 78.84 ; 
      RECT 95.872 74.466 95.976 78.84 ; 
      RECT 95.44 74.466 95.544 78.84 ; 
      RECT 95.008 74.466 95.112 78.84 ; 
      RECT 94.576 74.466 94.68 78.84 ; 
      RECT 94.144 74.466 94.248 78.84 ; 
      RECT 93.712 74.466 93.816 78.84 ; 
      RECT 93.28 74.466 93.384 78.84 ; 
      RECT 92.848 74.466 92.952 78.84 ; 
      RECT 92.416 74.466 92.52 78.84 ; 
      RECT 91.984 74.466 92.088 78.84 ; 
      RECT 91.552 74.466 91.656 78.84 ; 
      RECT 91.12 74.466 91.224 78.84 ; 
      RECT 90.688 74.466 90.792 78.84 ; 
      RECT 90.256 74.466 90.36 78.84 ; 
      RECT 89.824 74.466 89.928 78.84 ; 
      RECT 89.392 74.466 89.496 78.84 ; 
      RECT 88.96 74.466 89.064 78.84 ; 
      RECT 88.528 74.466 88.632 78.84 ; 
      RECT 88.096 74.466 88.2 78.84 ; 
      RECT 87.664 74.466 87.768 78.84 ; 
      RECT 87.232 74.466 87.336 78.84 ; 
      RECT 86.8 74.466 86.904 78.84 ; 
      RECT 86.368 74.466 86.472 78.84 ; 
      RECT 85.936 74.466 86.04 78.84 ; 
      RECT 85.504 74.466 85.608 78.84 ; 
      RECT 85.072 74.466 85.176 78.84 ; 
      RECT 84.64 74.466 84.744 78.84 ; 
      RECT 84.208 74.466 84.312 78.84 ; 
      RECT 83.776 74.466 83.88 78.84 ; 
      RECT 83.344 74.466 83.448 78.84 ; 
      RECT 82.912 74.466 83.016 78.84 ; 
      RECT 82.48 74.466 82.584 78.84 ; 
      RECT 82.048 74.466 82.152 78.84 ; 
      RECT 81.616 74.466 81.72 78.84 ; 
      RECT 81.184 74.466 81.288 78.84 ; 
      RECT 80.752 74.466 80.856 78.84 ; 
      RECT 80.32 74.466 80.424 78.84 ; 
      RECT 79.888 74.466 79.992 78.84 ; 
      RECT 79.456 74.466 79.56 78.84 ; 
      RECT 79.024 74.466 79.128 78.84 ; 
      RECT 78.592 74.466 78.696 78.84 ; 
      RECT 78.16 74.466 78.264 78.84 ; 
      RECT 77.728 74.466 77.832 78.84 ; 
      RECT 77.296 74.466 77.4 78.84 ; 
      RECT 76.864 74.466 76.968 78.84 ; 
      RECT 76.432 74.466 76.536 78.84 ; 
      RECT 76 74.466 76.104 78.84 ; 
      RECT 75.568 74.466 75.672 78.84 ; 
      RECT 75.136 74.466 75.24 78.84 ; 
      RECT 74.704 74.466 74.808 78.84 ; 
      RECT 74.272 74.466 74.376 78.84 ; 
      RECT 73.84 74.466 73.944 78.84 ; 
      RECT 73.408 74.466 73.512 78.84 ; 
      RECT 72.976 74.466 73.08 78.84 ; 
      RECT 72.544 74.466 72.648 78.84 ; 
      RECT 72.112 74.466 72.216 78.84 ; 
      RECT 71.68 74.466 71.784 78.84 ; 
      RECT 71.248 74.466 71.352 78.84 ; 
      RECT 70.816 74.466 70.92 78.84 ; 
      RECT 70.384 74.466 70.488 78.84 ; 
      RECT 69.952 74.466 70.056 78.84 ; 
      RECT 69.52 74.466 69.624 78.84 ; 
      RECT 69.088 74.466 69.192 78.84 ; 
      RECT 68.656 74.466 68.76 78.84 ; 
      RECT 68.224 74.466 68.328 78.84 ; 
      RECT 67.792 74.466 67.896 78.84 ; 
      RECT 67.36 74.466 67.464 78.84 ; 
      RECT 66.928 74.466 67.032 78.84 ; 
      RECT 66.496 74.466 66.6 78.84 ; 
      RECT 66.064 74.466 66.168 78.84 ; 
      RECT 65.632 74.466 65.736 78.84 ; 
      RECT 65.2 74.466 65.304 78.84 ; 
      RECT 64.348 74.466 64.656 78.84 ; 
      RECT 56.776 74.466 57.084 78.84 ; 
      RECT 56.128 74.466 56.232 78.84 ; 
      RECT 55.696 74.466 55.8 78.84 ; 
      RECT 55.264 74.466 55.368 78.84 ; 
      RECT 54.832 74.466 54.936 78.84 ; 
      RECT 54.4 74.466 54.504 78.84 ; 
      RECT 53.968 74.466 54.072 78.84 ; 
      RECT 53.536 74.466 53.64 78.84 ; 
      RECT 53.104 74.466 53.208 78.84 ; 
      RECT 52.672 74.466 52.776 78.84 ; 
      RECT 52.24 74.466 52.344 78.84 ; 
      RECT 51.808 74.466 51.912 78.84 ; 
      RECT 51.376 74.466 51.48 78.84 ; 
      RECT 50.944 74.466 51.048 78.84 ; 
      RECT 50.512 74.466 50.616 78.84 ; 
      RECT 50.08 74.466 50.184 78.84 ; 
      RECT 49.648 74.466 49.752 78.84 ; 
      RECT 49.216 74.466 49.32 78.84 ; 
      RECT 48.784 74.466 48.888 78.84 ; 
      RECT 48.352 74.466 48.456 78.84 ; 
      RECT 47.92 74.466 48.024 78.84 ; 
      RECT 47.488 74.466 47.592 78.84 ; 
      RECT 47.056 74.466 47.16 78.84 ; 
      RECT 46.624 74.466 46.728 78.84 ; 
      RECT 46.192 74.466 46.296 78.84 ; 
      RECT 45.76 74.466 45.864 78.84 ; 
      RECT 45.328 74.466 45.432 78.84 ; 
      RECT 44.896 74.466 45 78.84 ; 
      RECT 44.464 74.466 44.568 78.84 ; 
      RECT 44.032 74.466 44.136 78.84 ; 
      RECT 43.6 74.466 43.704 78.84 ; 
      RECT 43.168 74.466 43.272 78.84 ; 
      RECT 42.736 74.466 42.84 78.84 ; 
      RECT 42.304 74.466 42.408 78.84 ; 
      RECT 41.872 74.466 41.976 78.84 ; 
      RECT 41.44 74.466 41.544 78.84 ; 
      RECT 41.008 74.466 41.112 78.84 ; 
      RECT 40.576 74.466 40.68 78.84 ; 
      RECT 40.144 74.466 40.248 78.84 ; 
      RECT 39.712 74.466 39.816 78.84 ; 
      RECT 39.28 74.466 39.384 78.84 ; 
      RECT 38.848 74.466 38.952 78.84 ; 
      RECT 38.416 74.466 38.52 78.84 ; 
      RECT 37.984 74.466 38.088 78.84 ; 
      RECT 37.552 74.466 37.656 78.84 ; 
      RECT 37.12 74.466 37.224 78.84 ; 
      RECT 36.688 74.466 36.792 78.84 ; 
      RECT 36.256 74.466 36.36 78.84 ; 
      RECT 35.824 74.466 35.928 78.84 ; 
      RECT 35.392 74.466 35.496 78.84 ; 
      RECT 34.96 74.466 35.064 78.84 ; 
      RECT 34.528 74.466 34.632 78.84 ; 
      RECT 34.096 74.466 34.2 78.84 ; 
      RECT 33.664 74.466 33.768 78.84 ; 
      RECT 33.232 74.466 33.336 78.84 ; 
      RECT 32.8 74.466 32.904 78.84 ; 
      RECT 32.368 74.466 32.472 78.84 ; 
      RECT 31.936 74.466 32.04 78.84 ; 
      RECT 31.504 74.466 31.608 78.84 ; 
      RECT 31.072 74.466 31.176 78.84 ; 
      RECT 30.64 74.466 30.744 78.84 ; 
      RECT 30.208 74.466 30.312 78.84 ; 
      RECT 29.776 74.466 29.88 78.84 ; 
      RECT 29.344 74.466 29.448 78.84 ; 
      RECT 28.912 74.466 29.016 78.84 ; 
      RECT 28.48 74.466 28.584 78.84 ; 
      RECT 28.048 74.466 28.152 78.84 ; 
      RECT 27.616 74.466 27.72 78.84 ; 
      RECT 27.184 74.466 27.288 78.84 ; 
      RECT 26.752 74.466 26.856 78.84 ; 
      RECT 26.32 74.466 26.424 78.84 ; 
      RECT 25.888 74.466 25.992 78.84 ; 
      RECT 25.456 74.466 25.56 78.84 ; 
      RECT 25.024 74.466 25.128 78.84 ; 
      RECT 24.592 74.466 24.696 78.84 ; 
      RECT 24.16 74.466 24.264 78.84 ; 
      RECT 23.728 74.466 23.832 78.84 ; 
      RECT 23.296 74.466 23.4 78.84 ; 
      RECT 22.864 74.466 22.968 78.84 ; 
      RECT 22.432 74.466 22.536 78.84 ; 
      RECT 22 74.466 22.104 78.84 ; 
      RECT 21.568 74.466 21.672 78.84 ; 
      RECT 21.136 74.466 21.24 78.84 ; 
      RECT 20.704 74.466 20.808 78.84 ; 
      RECT 20.272 74.466 20.376 78.84 ; 
      RECT 19.84 74.466 19.944 78.84 ; 
      RECT 19.408 74.466 19.512 78.84 ; 
      RECT 18.976 74.466 19.08 78.84 ; 
      RECT 18.544 74.466 18.648 78.84 ; 
      RECT 18.112 74.466 18.216 78.84 ; 
      RECT 17.68 74.466 17.784 78.84 ; 
      RECT 17.248 74.466 17.352 78.84 ; 
      RECT 16.816 74.466 16.92 78.84 ; 
      RECT 16.384 74.466 16.488 78.84 ; 
      RECT 15.952 74.466 16.056 78.84 ; 
      RECT 15.52 74.466 15.624 78.84 ; 
      RECT 15.088 74.466 15.192 78.84 ; 
      RECT 14.656 74.466 14.76 78.84 ; 
      RECT 14.224 74.466 14.328 78.84 ; 
      RECT 13.792 74.466 13.896 78.84 ; 
      RECT 13.36 74.466 13.464 78.84 ; 
      RECT 12.928 74.466 13.032 78.84 ; 
      RECT 12.496 74.466 12.6 78.84 ; 
      RECT 12.064 74.466 12.168 78.84 ; 
      RECT 11.632 74.466 11.736 78.84 ; 
      RECT 11.2 74.466 11.304 78.84 ; 
      RECT 10.768 74.466 10.872 78.84 ; 
      RECT 10.336 74.466 10.44 78.84 ; 
      RECT 9.904 74.466 10.008 78.84 ; 
      RECT 9.472 74.466 9.576 78.84 ; 
      RECT 9.04 74.466 9.144 78.84 ; 
      RECT 8.608 74.466 8.712 78.84 ; 
      RECT 8.176 74.466 8.28 78.84 ; 
      RECT 7.744 74.466 7.848 78.84 ; 
      RECT 7.312 74.466 7.416 78.84 ; 
      RECT 6.88 74.466 6.984 78.84 ; 
      RECT 6.448 74.466 6.552 78.84 ; 
      RECT 6.016 74.466 6.12 78.84 ; 
      RECT 5.584 74.466 5.688 78.84 ; 
      RECT 5.152 74.466 5.256 78.84 ; 
      RECT 4.72 74.466 4.824 78.84 ; 
      RECT 4.288 74.466 4.392 78.84 ; 
      RECT 3.856 74.466 3.96 78.84 ; 
      RECT 3.424 74.466 3.528 78.84 ; 
      RECT 2.992 74.466 3.096 78.84 ; 
      RECT 2.56 74.466 2.664 78.84 ; 
      RECT 2.128 74.466 2.232 78.84 ; 
      RECT 1.696 74.466 1.8 78.84 ; 
      RECT 1.264 74.466 1.368 78.84 ; 
      RECT 0.832 74.466 0.936 78.84 ; 
      RECT 0.02 74.466 0.36 78.84 ; 
      RECT 62.212 78.786 62.724 83.16 ; 
      RECT 62.156 81.448 62.724 82.738 ; 
      RECT 61.276 80.356 61.812 83.16 ; 
      RECT 61.184 81.696 61.812 82.728 ; 
      RECT 61.276 78.786 61.668 83.16 ; 
      RECT 61.276 79.27 61.724 80.228 ; 
      RECT 61.276 78.786 61.812 79.142 ; 
      RECT 60.376 80.588 60.912 83.16 ; 
      RECT 60.376 78.786 60.768 83.16 ; 
      RECT 58.708 78.786 59.04 83.16 ; 
      RECT 58.708 79.14 59.096 82.882 ; 
      RECT 121.072 78.786 121.412 83.16 ; 
      RECT 120.496 78.786 120.6 83.16 ; 
      RECT 120.064 78.786 120.168 83.16 ; 
      RECT 119.632 78.786 119.736 83.16 ; 
      RECT 119.2 78.786 119.304 83.16 ; 
      RECT 118.768 78.786 118.872 83.16 ; 
      RECT 118.336 78.786 118.44 83.16 ; 
      RECT 117.904 78.786 118.008 83.16 ; 
      RECT 117.472 78.786 117.576 83.16 ; 
      RECT 117.04 78.786 117.144 83.16 ; 
      RECT 116.608 78.786 116.712 83.16 ; 
      RECT 116.176 78.786 116.28 83.16 ; 
      RECT 115.744 78.786 115.848 83.16 ; 
      RECT 115.312 78.786 115.416 83.16 ; 
      RECT 114.88 78.786 114.984 83.16 ; 
      RECT 114.448 78.786 114.552 83.16 ; 
      RECT 114.016 78.786 114.12 83.16 ; 
      RECT 113.584 78.786 113.688 83.16 ; 
      RECT 113.152 78.786 113.256 83.16 ; 
      RECT 112.72 78.786 112.824 83.16 ; 
      RECT 112.288 78.786 112.392 83.16 ; 
      RECT 111.856 78.786 111.96 83.16 ; 
      RECT 111.424 78.786 111.528 83.16 ; 
      RECT 110.992 78.786 111.096 83.16 ; 
      RECT 110.56 78.786 110.664 83.16 ; 
      RECT 110.128 78.786 110.232 83.16 ; 
      RECT 109.696 78.786 109.8 83.16 ; 
      RECT 109.264 78.786 109.368 83.16 ; 
      RECT 108.832 78.786 108.936 83.16 ; 
      RECT 108.4 78.786 108.504 83.16 ; 
      RECT 107.968 78.786 108.072 83.16 ; 
      RECT 107.536 78.786 107.64 83.16 ; 
      RECT 107.104 78.786 107.208 83.16 ; 
      RECT 106.672 78.786 106.776 83.16 ; 
      RECT 106.24 78.786 106.344 83.16 ; 
      RECT 105.808 78.786 105.912 83.16 ; 
      RECT 105.376 78.786 105.48 83.16 ; 
      RECT 104.944 78.786 105.048 83.16 ; 
      RECT 104.512 78.786 104.616 83.16 ; 
      RECT 104.08 78.786 104.184 83.16 ; 
      RECT 103.648 78.786 103.752 83.16 ; 
      RECT 103.216 78.786 103.32 83.16 ; 
      RECT 102.784 78.786 102.888 83.16 ; 
      RECT 102.352 78.786 102.456 83.16 ; 
      RECT 101.92 78.786 102.024 83.16 ; 
      RECT 101.488 78.786 101.592 83.16 ; 
      RECT 101.056 78.786 101.16 83.16 ; 
      RECT 100.624 78.786 100.728 83.16 ; 
      RECT 100.192 78.786 100.296 83.16 ; 
      RECT 99.76 78.786 99.864 83.16 ; 
      RECT 99.328 78.786 99.432 83.16 ; 
      RECT 98.896 78.786 99 83.16 ; 
      RECT 98.464 78.786 98.568 83.16 ; 
      RECT 98.032 78.786 98.136 83.16 ; 
      RECT 97.6 78.786 97.704 83.16 ; 
      RECT 97.168 78.786 97.272 83.16 ; 
      RECT 96.736 78.786 96.84 83.16 ; 
      RECT 96.304 78.786 96.408 83.16 ; 
      RECT 95.872 78.786 95.976 83.16 ; 
      RECT 95.44 78.786 95.544 83.16 ; 
      RECT 95.008 78.786 95.112 83.16 ; 
      RECT 94.576 78.786 94.68 83.16 ; 
      RECT 94.144 78.786 94.248 83.16 ; 
      RECT 93.712 78.786 93.816 83.16 ; 
      RECT 93.28 78.786 93.384 83.16 ; 
      RECT 92.848 78.786 92.952 83.16 ; 
      RECT 92.416 78.786 92.52 83.16 ; 
      RECT 91.984 78.786 92.088 83.16 ; 
      RECT 91.552 78.786 91.656 83.16 ; 
      RECT 91.12 78.786 91.224 83.16 ; 
      RECT 90.688 78.786 90.792 83.16 ; 
      RECT 90.256 78.786 90.36 83.16 ; 
      RECT 89.824 78.786 89.928 83.16 ; 
      RECT 89.392 78.786 89.496 83.16 ; 
      RECT 88.96 78.786 89.064 83.16 ; 
      RECT 88.528 78.786 88.632 83.16 ; 
      RECT 88.096 78.786 88.2 83.16 ; 
      RECT 87.664 78.786 87.768 83.16 ; 
      RECT 87.232 78.786 87.336 83.16 ; 
      RECT 86.8 78.786 86.904 83.16 ; 
      RECT 86.368 78.786 86.472 83.16 ; 
      RECT 85.936 78.786 86.04 83.16 ; 
      RECT 85.504 78.786 85.608 83.16 ; 
      RECT 85.072 78.786 85.176 83.16 ; 
      RECT 84.64 78.786 84.744 83.16 ; 
      RECT 84.208 78.786 84.312 83.16 ; 
      RECT 83.776 78.786 83.88 83.16 ; 
      RECT 83.344 78.786 83.448 83.16 ; 
      RECT 82.912 78.786 83.016 83.16 ; 
      RECT 82.48 78.786 82.584 83.16 ; 
      RECT 82.048 78.786 82.152 83.16 ; 
      RECT 81.616 78.786 81.72 83.16 ; 
      RECT 81.184 78.786 81.288 83.16 ; 
      RECT 80.752 78.786 80.856 83.16 ; 
      RECT 80.32 78.786 80.424 83.16 ; 
      RECT 79.888 78.786 79.992 83.16 ; 
      RECT 79.456 78.786 79.56 83.16 ; 
      RECT 79.024 78.786 79.128 83.16 ; 
      RECT 78.592 78.786 78.696 83.16 ; 
      RECT 78.16 78.786 78.264 83.16 ; 
      RECT 77.728 78.786 77.832 83.16 ; 
      RECT 77.296 78.786 77.4 83.16 ; 
      RECT 76.864 78.786 76.968 83.16 ; 
      RECT 76.432 78.786 76.536 83.16 ; 
      RECT 76 78.786 76.104 83.16 ; 
      RECT 75.568 78.786 75.672 83.16 ; 
      RECT 75.136 78.786 75.24 83.16 ; 
      RECT 74.704 78.786 74.808 83.16 ; 
      RECT 74.272 78.786 74.376 83.16 ; 
      RECT 73.84 78.786 73.944 83.16 ; 
      RECT 73.408 78.786 73.512 83.16 ; 
      RECT 72.976 78.786 73.08 83.16 ; 
      RECT 72.544 78.786 72.648 83.16 ; 
      RECT 72.112 78.786 72.216 83.16 ; 
      RECT 71.68 78.786 71.784 83.16 ; 
      RECT 71.248 78.786 71.352 83.16 ; 
      RECT 70.816 78.786 70.92 83.16 ; 
      RECT 70.384 78.786 70.488 83.16 ; 
      RECT 69.952 78.786 70.056 83.16 ; 
      RECT 69.52 78.786 69.624 83.16 ; 
      RECT 69.088 78.786 69.192 83.16 ; 
      RECT 68.656 78.786 68.76 83.16 ; 
      RECT 68.224 78.786 68.328 83.16 ; 
      RECT 67.792 78.786 67.896 83.16 ; 
      RECT 67.36 78.786 67.464 83.16 ; 
      RECT 66.928 78.786 67.032 83.16 ; 
      RECT 66.496 78.786 66.6 83.16 ; 
      RECT 66.064 78.786 66.168 83.16 ; 
      RECT 65.632 78.786 65.736 83.16 ; 
      RECT 65.2 78.786 65.304 83.16 ; 
      RECT 64.348 78.786 64.656 83.16 ; 
      RECT 56.776 78.786 57.084 83.16 ; 
      RECT 56.128 78.786 56.232 83.16 ; 
      RECT 55.696 78.786 55.8 83.16 ; 
      RECT 55.264 78.786 55.368 83.16 ; 
      RECT 54.832 78.786 54.936 83.16 ; 
      RECT 54.4 78.786 54.504 83.16 ; 
      RECT 53.968 78.786 54.072 83.16 ; 
      RECT 53.536 78.786 53.64 83.16 ; 
      RECT 53.104 78.786 53.208 83.16 ; 
      RECT 52.672 78.786 52.776 83.16 ; 
      RECT 52.24 78.786 52.344 83.16 ; 
      RECT 51.808 78.786 51.912 83.16 ; 
      RECT 51.376 78.786 51.48 83.16 ; 
      RECT 50.944 78.786 51.048 83.16 ; 
      RECT 50.512 78.786 50.616 83.16 ; 
      RECT 50.08 78.786 50.184 83.16 ; 
      RECT 49.648 78.786 49.752 83.16 ; 
      RECT 49.216 78.786 49.32 83.16 ; 
      RECT 48.784 78.786 48.888 83.16 ; 
      RECT 48.352 78.786 48.456 83.16 ; 
      RECT 47.92 78.786 48.024 83.16 ; 
      RECT 47.488 78.786 47.592 83.16 ; 
      RECT 47.056 78.786 47.16 83.16 ; 
      RECT 46.624 78.786 46.728 83.16 ; 
      RECT 46.192 78.786 46.296 83.16 ; 
      RECT 45.76 78.786 45.864 83.16 ; 
      RECT 45.328 78.786 45.432 83.16 ; 
      RECT 44.896 78.786 45 83.16 ; 
      RECT 44.464 78.786 44.568 83.16 ; 
      RECT 44.032 78.786 44.136 83.16 ; 
      RECT 43.6 78.786 43.704 83.16 ; 
      RECT 43.168 78.786 43.272 83.16 ; 
      RECT 42.736 78.786 42.84 83.16 ; 
      RECT 42.304 78.786 42.408 83.16 ; 
      RECT 41.872 78.786 41.976 83.16 ; 
      RECT 41.44 78.786 41.544 83.16 ; 
      RECT 41.008 78.786 41.112 83.16 ; 
      RECT 40.576 78.786 40.68 83.16 ; 
      RECT 40.144 78.786 40.248 83.16 ; 
      RECT 39.712 78.786 39.816 83.16 ; 
      RECT 39.28 78.786 39.384 83.16 ; 
      RECT 38.848 78.786 38.952 83.16 ; 
      RECT 38.416 78.786 38.52 83.16 ; 
      RECT 37.984 78.786 38.088 83.16 ; 
      RECT 37.552 78.786 37.656 83.16 ; 
      RECT 37.12 78.786 37.224 83.16 ; 
      RECT 36.688 78.786 36.792 83.16 ; 
      RECT 36.256 78.786 36.36 83.16 ; 
      RECT 35.824 78.786 35.928 83.16 ; 
      RECT 35.392 78.786 35.496 83.16 ; 
      RECT 34.96 78.786 35.064 83.16 ; 
      RECT 34.528 78.786 34.632 83.16 ; 
      RECT 34.096 78.786 34.2 83.16 ; 
      RECT 33.664 78.786 33.768 83.16 ; 
      RECT 33.232 78.786 33.336 83.16 ; 
      RECT 32.8 78.786 32.904 83.16 ; 
      RECT 32.368 78.786 32.472 83.16 ; 
      RECT 31.936 78.786 32.04 83.16 ; 
      RECT 31.504 78.786 31.608 83.16 ; 
      RECT 31.072 78.786 31.176 83.16 ; 
      RECT 30.64 78.786 30.744 83.16 ; 
      RECT 30.208 78.786 30.312 83.16 ; 
      RECT 29.776 78.786 29.88 83.16 ; 
      RECT 29.344 78.786 29.448 83.16 ; 
      RECT 28.912 78.786 29.016 83.16 ; 
      RECT 28.48 78.786 28.584 83.16 ; 
      RECT 28.048 78.786 28.152 83.16 ; 
      RECT 27.616 78.786 27.72 83.16 ; 
      RECT 27.184 78.786 27.288 83.16 ; 
      RECT 26.752 78.786 26.856 83.16 ; 
      RECT 26.32 78.786 26.424 83.16 ; 
      RECT 25.888 78.786 25.992 83.16 ; 
      RECT 25.456 78.786 25.56 83.16 ; 
      RECT 25.024 78.786 25.128 83.16 ; 
      RECT 24.592 78.786 24.696 83.16 ; 
      RECT 24.16 78.786 24.264 83.16 ; 
      RECT 23.728 78.786 23.832 83.16 ; 
      RECT 23.296 78.786 23.4 83.16 ; 
      RECT 22.864 78.786 22.968 83.16 ; 
      RECT 22.432 78.786 22.536 83.16 ; 
      RECT 22 78.786 22.104 83.16 ; 
      RECT 21.568 78.786 21.672 83.16 ; 
      RECT 21.136 78.786 21.24 83.16 ; 
      RECT 20.704 78.786 20.808 83.16 ; 
      RECT 20.272 78.786 20.376 83.16 ; 
      RECT 19.84 78.786 19.944 83.16 ; 
      RECT 19.408 78.786 19.512 83.16 ; 
      RECT 18.976 78.786 19.08 83.16 ; 
      RECT 18.544 78.786 18.648 83.16 ; 
      RECT 18.112 78.786 18.216 83.16 ; 
      RECT 17.68 78.786 17.784 83.16 ; 
      RECT 17.248 78.786 17.352 83.16 ; 
      RECT 16.816 78.786 16.92 83.16 ; 
      RECT 16.384 78.786 16.488 83.16 ; 
      RECT 15.952 78.786 16.056 83.16 ; 
      RECT 15.52 78.786 15.624 83.16 ; 
      RECT 15.088 78.786 15.192 83.16 ; 
      RECT 14.656 78.786 14.76 83.16 ; 
      RECT 14.224 78.786 14.328 83.16 ; 
      RECT 13.792 78.786 13.896 83.16 ; 
      RECT 13.36 78.786 13.464 83.16 ; 
      RECT 12.928 78.786 13.032 83.16 ; 
      RECT 12.496 78.786 12.6 83.16 ; 
      RECT 12.064 78.786 12.168 83.16 ; 
      RECT 11.632 78.786 11.736 83.16 ; 
      RECT 11.2 78.786 11.304 83.16 ; 
      RECT 10.768 78.786 10.872 83.16 ; 
      RECT 10.336 78.786 10.44 83.16 ; 
      RECT 9.904 78.786 10.008 83.16 ; 
      RECT 9.472 78.786 9.576 83.16 ; 
      RECT 9.04 78.786 9.144 83.16 ; 
      RECT 8.608 78.786 8.712 83.16 ; 
      RECT 8.176 78.786 8.28 83.16 ; 
      RECT 7.744 78.786 7.848 83.16 ; 
      RECT 7.312 78.786 7.416 83.16 ; 
      RECT 6.88 78.786 6.984 83.16 ; 
      RECT 6.448 78.786 6.552 83.16 ; 
      RECT 6.016 78.786 6.12 83.16 ; 
      RECT 5.584 78.786 5.688 83.16 ; 
      RECT 5.152 78.786 5.256 83.16 ; 
      RECT 4.72 78.786 4.824 83.16 ; 
      RECT 4.288 78.786 4.392 83.16 ; 
      RECT 3.856 78.786 3.96 83.16 ; 
      RECT 3.424 78.786 3.528 83.16 ; 
      RECT 2.992 78.786 3.096 83.16 ; 
      RECT 2.56 78.786 2.664 83.16 ; 
      RECT 2.128 78.786 2.232 83.16 ; 
      RECT 1.696 78.786 1.8 83.16 ; 
      RECT 1.264 78.786 1.368 83.16 ; 
      RECT 0.832 78.786 0.936 83.16 ; 
      RECT 0.02 78.786 0.36 83.16 ; 
      RECT 62.212 83.106 62.724 87.48 ; 
      RECT 62.156 85.768 62.724 87.058 ; 
      RECT 61.276 84.676 61.812 87.48 ; 
      RECT 61.184 86.016 61.812 87.048 ; 
      RECT 61.276 83.106 61.668 87.48 ; 
      RECT 61.276 83.59 61.724 84.548 ; 
      RECT 61.276 83.106 61.812 83.462 ; 
      RECT 60.376 84.908 60.912 87.48 ; 
      RECT 60.376 83.106 60.768 87.48 ; 
      RECT 58.708 83.106 59.04 87.48 ; 
      RECT 58.708 83.46 59.096 87.202 ; 
      RECT 121.072 83.106 121.412 87.48 ; 
      RECT 120.496 83.106 120.6 87.48 ; 
      RECT 120.064 83.106 120.168 87.48 ; 
      RECT 119.632 83.106 119.736 87.48 ; 
      RECT 119.2 83.106 119.304 87.48 ; 
      RECT 118.768 83.106 118.872 87.48 ; 
      RECT 118.336 83.106 118.44 87.48 ; 
      RECT 117.904 83.106 118.008 87.48 ; 
      RECT 117.472 83.106 117.576 87.48 ; 
      RECT 117.04 83.106 117.144 87.48 ; 
      RECT 116.608 83.106 116.712 87.48 ; 
      RECT 116.176 83.106 116.28 87.48 ; 
      RECT 115.744 83.106 115.848 87.48 ; 
      RECT 115.312 83.106 115.416 87.48 ; 
      RECT 114.88 83.106 114.984 87.48 ; 
      RECT 114.448 83.106 114.552 87.48 ; 
      RECT 114.016 83.106 114.12 87.48 ; 
      RECT 113.584 83.106 113.688 87.48 ; 
      RECT 113.152 83.106 113.256 87.48 ; 
      RECT 112.72 83.106 112.824 87.48 ; 
      RECT 112.288 83.106 112.392 87.48 ; 
      RECT 111.856 83.106 111.96 87.48 ; 
      RECT 111.424 83.106 111.528 87.48 ; 
      RECT 110.992 83.106 111.096 87.48 ; 
      RECT 110.56 83.106 110.664 87.48 ; 
      RECT 110.128 83.106 110.232 87.48 ; 
      RECT 109.696 83.106 109.8 87.48 ; 
      RECT 109.264 83.106 109.368 87.48 ; 
      RECT 108.832 83.106 108.936 87.48 ; 
      RECT 108.4 83.106 108.504 87.48 ; 
      RECT 107.968 83.106 108.072 87.48 ; 
      RECT 107.536 83.106 107.64 87.48 ; 
      RECT 107.104 83.106 107.208 87.48 ; 
      RECT 106.672 83.106 106.776 87.48 ; 
      RECT 106.24 83.106 106.344 87.48 ; 
      RECT 105.808 83.106 105.912 87.48 ; 
      RECT 105.376 83.106 105.48 87.48 ; 
      RECT 104.944 83.106 105.048 87.48 ; 
      RECT 104.512 83.106 104.616 87.48 ; 
      RECT 104.08 83.106 104.184 87.48 ; 
      RECT 103.648 83.106 103.752 87.48 ; 
      RECT 103.216 83.106 103.32 87.48 ; 
      RECT 102.784 83.106 102.888 87.48 ; 
      RECT 102.352 83.106 102.456 87.48 ; 
      RECT 101.92 83.106 102.024 87.48 ; 
      RECT 101.488 83.106 101.592 87.48 ; 
      RECT 101.056 83.106 101.16 87.48 ; 
      RECT 100.624 83.106 100.728 87.48 ; 
      RECT 100.192 83.106 100.296 87.48 ; 
      RECT 99.76 83.106 99.864 87.48 ; 
      RECT 99.328 83.106 99.432 87.48 ; 
      RECT 98.896 83.106 99 87.48 ; 
      RECT 98.464 83.106 98.568 87.48 ; 
      RECT 98.032 83.106 98.136 87.48 ; 
      RECT 97.6 83.106 97.704 87.48 ; 
      RECT 97.168 83.106 97.272 87.48 ; 
      RECT 96.736 83.106 96.84 87.48 ; 
      RECT 96.304 83.106 96.408 87.48 ; 
      RECT 95.872 83.106 95.976 87.48 ; 
      RECT 95.44 83.106 95.544 87.48 ; 
      RECT 95.008 83.106 95.112 87.48 ; 
      RECT 94.576 83.106 94.68 87.48 ; 
      RECT 94.144 83.106 94.248 87.48 ; 
      RECT 93.712 83.106 93.816 87.48 ; 
      RECT 93.28 83.106 93.384 87.48 ; 
      RECT 92.848 83.106 92.952 87.48 ; 
      RECT 92.416 83.106 92.52 87.48 ; 
      RECT 91.984 83.106 92.088 87.48 ; 
      RECT 91.552 83.106 91.656 87.48 ; 
      RECT 91.12 83.106 91.224 87.48 ; 
      RECT 90.688 83.106 90.792 87.48 ; 
      RECT 90.256 83.106 90.36 87.48 ; 
      RECT 89.824 83.106 89.928 87.48 ; 
      RECT 89.392 83.106 89.496 87.48 ; 
      RECT 88.96 83.106 89.064 87.48 ; 
      RECT 88.528 83.106 88.632 87.48 ; 
      RECT 88.096 83.106 88.2 87.48 ; 
      RECT 87.664 83.106 87.768 87.48 ; 
      RECT 87.232 83.106 87.336 87.48 ; 
      RECT 86.8 83.106 86.904 87.48 ; 
      RECT 86.368 83.106 86.472 87.48 ; 
      RECT 85.936 83.106 86.04 87.48 ; 
      RECT 85.504 83.106 85.608 87.48 ; 
      RECT 85.072 83.106 85.176 87.48 ; 
      RECT 84.64 83.106 84.744 87.48 ; 
      RECT 84.208 83.106 84.312 87.48 ; 
      RECT 83.776 83.106 83.88 87.48 ; 
      RECT 83.344 83.106 83.448 87.48 ; 
      RECT 82.912 83.106 83.016 87.48 ; 
      RECT 82.48 83.106 82.584 87.48 ; 
      RECT 82.048 83.106 82.152 87.48 ; 
      RECT 81.616 83.106 81.72 87.48 ; 
      RECT 81.184 83.106 81.288 87.48 ; 
      RECT 80.752 83.106 80.856 87.48 ; 
      RECT 80.32 83.106 80.424 87.48 ; 
      RECT 79.888 83.106 79.992 87.48 ; 
      RECT 79.456 83.106 79.56 87.48 ; 
      RECT 79.024 83.106 79.128 87.48 ; 
      RECT 78.592 83.106 78.696 87.48 ; 
      RECT 78.16 83.106 78.264 87.48 ; 
      RECT 77.728 83.106 77.832 87.48 ; 
      RECT 77.296 83.106 77.4 87.48 ; 
      RECT 76.864 83.106 76.968 87.48 ; 
      RECT 76.432 83.106 76.536 87.48 ; 
      RECT 76 83.106 76.104 87.48 ; 
      RECT 75.568 83.106 75.672 87.48 ; 
      RECT 75.136 83.106 75.24 87.48 ; 
      RECT 74.704 83.106 74.808 87.48 ; 
      RECT 74.272 83.106 74.376 87.48 ; 
      RECT 73.84 83.106 73.944 87.48 ; 
      RECT 73.408 83.106 73.512 87.48 ; 
      RECT 72.976 83.106 73.08 87.48 ; 
      RECT 72.544 83.106 72.648 87.48 ; 
      RECT 72.112 83.106 72.216 87.48 ; 
      RECT 71.68 83.106 71.784 87.48 ; 
      RECT 71.248 83.106 71.352 87.48 ; 
      RECT 70.816 83.106 70.92 87.48 ; 
      RECT 70.384 83.106 70.488 87.48 ; 
      RECT 69.952 83.106 70.056 87.48 ; 
      RECT 69.52 83.106 69.624 87.48 ; 
      RECT 69.088 83.106 69.192 87.48 ; 
      RECT 68.656 83.106 68.76 87.48 ; 
      RECT 68.224 83.106 68.328 87.48 ; 
      RECT 67.792 83.106 67.896 87.48 ; 
      RECT 67.36 83.106 67.464 87.48 ; 
      RECT 66.928 83.106 67.032 87.48 ; 
      RECT 66.496 83.106 66.6 87.48 ; 
      RECT 66.064 83.106 66.168 87.48 ; 
      RECT 65.632 83.106 65.736 87.48 ; 
      RECT 65.2 83.106 65.304 87.48 ; 
      RECT 64.348 83.106 64.656 87.48 ; 
      RECT 56.776 83.106 57.084 87.48 ; 
      RECT 56.128 83.106 56.232 87.48 ; 
      RECT 55.696 83.106 55.8 87.48 ; 
      RECT 55.264 83.106 55.368 87.48 ; 
      RECT 54.832 83.106 54.936 87.48 ; 
      RECT 54.4 83.106 54.504 87.48 ; 
      RECT 53.968 83.106 54.072 87.48 ; 
      RECT 53.536 83.106 53.64 87.48 ; 
      RECT 53.104 83.106 53.208 87.48 ; 
      RECT 52.672 83.106 52.776 87.48 ; 
      RECT 52.24 83.106 52.344 87.48 ; 
      RECT 51.808 83.106 51.912 87.48 ; 
      RECT 51.376 83.106 51.48 87.48 ; 
      RECT 50.944 83.106 51.048 87.48 ; 
      RECT 50.512 83.106 50.616 87.48 ; 
      RECT 50.08 83.106 50.184 87.48 ; 
      RECT 49.648 83.106 49.752 87.48 ; 
      RECT 49.216 83.106 49.32 87.48 ; 
      RECT 48.784 83.106 48.888 87.48 ; 
      RECT 48.352 83.106 48.456 87.48 ; 
      RECT 47.92 83.106 48.024 87.48 ; 
      RECT 47.488 83.106 47.592 87.48 ; 
      RECT 47.056 83.106 47.16 87.48 ; 
      RECT 46.624 83.106 46.728 87.48 ; 
      RECT 46.192 83.106 46.296 87.48 ; 
      RECT 45.76 83.106 45.864 87.48 ; 
      RECT 45.328 83.106 45.432 87.48 ; 
      RECT 44.896 83.106 45 87.48 ; 
      RECT 44.464 83.106 44.568 87.48 ; 
      RECT 44.032 83.106 44.136 87.48 ; 
      RECT 43.6 83.106 43.704 87.48 ; 
      RECT 43.168 83.106 43.272 87.48 ; 
      RECT 42.736 83.106 42.84 87.48 ; 
      RECT 42.304 83.106 42.408 87.48 ; 
      RECT 41.872 83.106 41.976 87.48 ; 
      RECT 41.44 83.106 41.544 87.48 ; 
      RECT 41.008 83.106 41.112 87.48 ; 
      RECT 40.576 83.106 40.68 87.48 ; 
      RECT 40.144 83.106 40.248 87.48 ; 
      RECT 39.712 83.106 39.816 87.48 ; 
      RECT 39.28 83.106 39.384 87.48 ; 
      RECT 38.848 83.106 38.952 87.48 ; 
      RECT 38.416 83.106 38.52 87.48 ; 
      RECT 37.984 83.106 38.088 87.48 ; 
      RECT 37.552 83.106 37.656 87.48 ; 
      RECT 37.12 83.106 37.224 87.48 ; 
      RECT 36.688 83.106 36.792 87.48 ; 
      RECT 36.256 83.106 36.36 87.48 ; 
      RECT 35.824 83.106 35.928 87.48 ; 
      RECT 35.392 83.106 35.496 87.48 ; 
      RECT 34.96 83.106 35.064 87.48 ; 
      RECT 34.528 83.106 34.632 87.48 ; 
      RECT 34.096 83.106 34.2 87.48 ; 
      RECT 33.664 83.106 33.768 87.48 ; 
      RECT 33.232 83.106 33.336 87.48 ; 
      RECT 32.8 83.106 32.904 87.48 ; 
      RECT 32.368 83.106 32.472 87.48 ; 
      RECT 31.936 83.106 32.04 87.48 ; 
      RECT 31.504 83.106 31.608 87.48 ; 
      RECT 31.072 83.106 31.176 87.48 ; 
      RECT 30.64 83.106 30.744 87.48 ; 
      RECT 30.208 83.106 30.312 87.48 ; 
      RECT 29.776 83.106 29.88 87.48 ; 
      RECT 29.344 83.106 29.448 87.48 ; 
      RECT 28.912 83.106 29.016 87.48 ; 
      RECT 28.48 83.106 28.584 87.48 ; 
      RECT 28.048 83.106 28.152 87.48 ; 
      RECT 27.616 83.106 27.72 87.48 ; 
      RECT 27.184 83.106 27.288 87.48 ; 
      RECT 26.752 83.106 26.856 87.48 ; 
      RECT 26.32 83.106 26.424 87.48 ; 
      RECT 25.888 83.106 25.992 87.48 ; 
      RECT 25.456 83.106 25.56 87.48 ; 
      RECT 25.024 83.106 25.128 87.48 ; 
      RECT 24.592 83.106 24.696 87.48 ; 
      RECT 24.16 83.106 24.264 87.48 ; 
      RECT 23.728 83.106 23.832 87.48 ; 
      RECT 23.296 83.106 23.4 87.48 ; 
      RECT 22.864 83.106 22.968 87.48 ; 
      RECT 22.432 83.106 22.536 87.48 ; 
      RECT 22 83.106 22.104 87.48 ; 
      RECT 21.568 83.106 21.672 87.48 ; 
      RECT 21.136 83.106 21.24 87.48 ; 
      RECT 20.704 83.106 20.808 87.48 ; 
      RECT 20.272 83.106 20.376 87.48 ; 
      RECT 19.84 83.106 19.944 87.48 ; 
      RECT 19.408 83.106 19.512 87.48 ; 
      RECT 18.976 83.106 19.08 87.48 ; 
      RECT 18.544 83.106 18.648 87.48 ; 
      RECT 18.112 83.106 18.216 87.48 ; 
      RECT 17.68 83.106 17.784 87.48 ; 
      RECT 17.248 83.106 17.352 87.48 ; 
      RECT 16.816 83.106 16.92 87.48 ; 
      RECT 16.384 83.106 16.488 87.48 ; 
      RECT 15.952 83.106 16.056 87.48 ; 
      RECT 15.52 83.106 15.624 87.48 ; 
      RECT 15.088 83.106 15.192 87.48 ; 
      RECT 14.656 83.106 14.76 87.48 ; 
      RECT 14.224 83.106 14.328 87.48 ; 
      RECT 13.792 83.106 13.896 87.48 ; 
      RECT 13.36 83.106 13.464 87.48 ; 
      RECT 12.928 83.106 13.032 87.48 ; 
      RECT 12.496 83.106 12.6 87.48 ; 
      RECT 12.064 83.106 12.168 87.48 ; 
      RECT 11.632 83.106 11.736 87.48 ; 
      RECT 11.2 83.106 11.304 87.48 ; 
      RECT 10.768 83.106 10.872 87.48 ; 
      RECT 10.336 83.106 10.44 87.48 ; 
      RECT 9.904 83.106 10.008 87.48 ; 
      RECT 9.472 83.106 9.576 87.48 ; 
      RECT 9.04 83.106 9.144 87.48 ; 
      RECT 8.608 83.106 8.712 87.48 ; 
      RECT 8.176 83.106 8.28 87.48 ; 
      RECT 7.744 83.106 7.848 87.48 ; 
      RECT 7.312 83.106 7.416 87.48 ; 
      RECT 6.88 83.106 6.984 87.48 ; 
      RECT 6.448 83.106 6.552 87.48 ; 
      RECT 6.016 83.106 6.12 87.48 ; 
      RECT 5.584 83.106 5.688 87.48 ; 
      RECT 5.152 83.106 5.256 87.48 ; 
      RECT 4.72 83.106 4.824 87.48 ; 
      RECT 4.288 83.106 4.392 87.48 ; 
      RECT 3.856 83.106 3.96 87.48 ; 
      RECT 3.424 83.106 3.528 87.48 ; 
      RECT 2.992 83.106 3.096 87.48 ; 
      RECT 2.56 83.106 2.664 87.48 ; 
      RECT 2.128 83.106 2.232 87.48 ; 
      RECT 1.696 83.106 1.8 87.48 ; 
      RECT 1.264 83.106 1.368 87.48 ; 
      RECT 0.832 83.106 0.936 87.48 ; 
      RECT 0.02 83.106 0.36 87.48 ; 
      RECT 62.212 87.426 62.724 91.8 ; 
      RECT 62.156 90.088 62.724 91.378 ; 
      RECT 61.276 88.996 61.812 91.8 ; 
      RECT 61.184 90.336 61.812 91.368 ; 
      RECT 61.276 87.426 61.668 91.8 ; 
      RECT 61.276 87.91 61.724 88.868 ; 
      RECT 61.276 87.426 61.812 87.782 ; 
      RECT 60.376 89.228 60.912 91.8 ; 
      RECT 60.376 87.426 60.768 91.8 ; 
      RECT 58.708 87.426 59.04 91.8 ; 
      RECT 58.708 87.78 59.096 91.522 ; 
      RECT 121.072 87.426 121.412 91.8 ; 
      RECT 120.496 87.426 120.6 91.8 ; 
      RECT 120.064 87.426 120.168 91.8 ; 
      RECT 119.632 87.426 119.736 91.8 ; 
      RECT 119.2 87.426 119.304 91.8 ; 
      RECT 118.768 87.426 118.872 91.8 ; 
      RECT 118.336 87.426 118.44 91.8 ; 
      RECT 117.904 87.426 118.008 91.8 ; 
      RECT 117.472 87.426 117.576 91.8 ; 
      RECT 117.04 87.426 117.144 91.8 ; 
      RECT 116.608 87.426 116.712 91.8 ; 
      RECT 116.176 87.426 116.28 91.8 ; 
      RECT 115.744 87.426 115.848 91.8 ; 
      RECT 115.312 87.426 115.416 91.8 ; 
      RECT 114.88 87.426 114.984 91.8 ; 
      RECT 114.448 87.426 114.552 91.8 ; 
      RECT 114.016 87.426 114.12 91.8 ; 
      RECT 113.584 87.426 113.688 91.8 ; 
      RECT 113.152 87.426 113.256 91.8 ; 
      RECT 112.72 87.426 112.824 91.8 ; 
      RECT 112.288 87.426 112.392 91.8 ; 
      RECT 111.856 87.426 111.96 91.8 ; 
      RECT 111.424 87.426 111.528 91.8 ; 
      RECT 110.992 87.426 111.096 91.8 ; 
      RECT 110.56 87.426 110.664 91.8 ; 
      RECT 110.128 87.426 110.232 91.8 ; 
      RECT 109.696 87.426 109.8 91.8 ; 
      RECT 109.264 87.426 109.368 91.8 ; 
      RECT 108.832 87.426 108.936 91.8 ; 
      RECT 108.4 87.426 108.504 91.8 ; 
      RECT 107.968 87.426 108.072 91.8 ; 
      RECT 107.536 87.426 107.64 91.8 ; 
      RECT 107.104 87.426 107.208 91.8 ; 
      RECT 106.672 87.426 106.776 91.8 ; 
      RECT 106.24 87.426 106.344 91.8 ; 
      RECT 105.808 87.426 105.912 91.8 ; 
      RECT 105.376 87.426 105.48 91.8 ; 
      RECT 104.944 87.426 105.048 91.8 ; 
      RECT 104.512 87.426 104.616 91.8 ; 
      RECT 104.08 87.426 104.184 91.8 ; 
      RECT 103.648 87.426 103.752 91.8 ; 
      RECT 103.216 87.426 103.32 91.8 ; 
      RECT 102.784 87.426 102.888 91.8 ; 
      RECT 102.352 87.426 102.456 91.8 ; 
      RECT 101.92 87.426 102.024 91.8 ; 
      RECT 101.488 87.426 101.592 91.8 ; 
      RECT 101.056 87.426 101.16 91.8 ; 
      RECT 100.624 87.426 100.728 91.8 ; 
      RECT 100.192 87.426 100.296 91.8 ; 
      RECT 99.76 87.426 99.864 91.8 ; 
      RECT 99.328 87.426 99.432 91.8 ; 
      RECT 98.896 87.426 99 91.8 ; 
      RECT 98.464 87.426 98.568 91.8 ; 
      RECT 98.032 87.426 98.136 91.8 ; 
      RECT 97.6 87.426 97.704 91.8 ; 
      RECT 97.168 87.426 97.272 91.8 ; 
      RECT 96.736 87.426 96.84 91.8 ; 
      RECT 96.304 87.426 96.408 91.8 ; 
      RECT 95.872 87.426 95.976 91.8 ; 
      RECT 95.44 87.426 95.544 91.8 ; 
      RECT 95.008 87.426 95.112 91.8 ; 
      RECT 94.576 87.426 94.68 91.8 ; 
      RECT 94.144 87.426 94.248 91.8 ; 
      RECT 93.712 87.426 93.816 91.8 ; 
      RECT 93.28 87.426 93.384 91.8 ; 
      RECT 92.848 87.426 92.952 91.8 ; 
      RECT 92.416 87.426 92.52 91.8 ; 
      RECT 91.984 87.426 92.088 91.8 ; 
      RECT 91.552 87.426 91.656 91.8 ; 
      RECT 91.12 87.426 91.224 91.8 ; 
      RECT 90.688 87.426 90.792 91.8 ; 
      RECT 90.256 87.426 90.36 91.8 ; 
      RECT 89.824 87.426 89.928 91.8 ; 
      RECT 89.392 87.426 89.496 91.8 ; 
      RECT 88.96 87.426 89.064 91.8 ; 
      RECT 88.528 87.426 88.632 91.8 ; 
      RECT 88.096 87.426 88.2 91.8 ; 
      RECT 87.664 87.426 87.768 91.8 ; 
      RECT 87.232 87.426 87.336 91.8 ; 
      RECT 86.8 87.426 86.904 91.8 ; 
      RECT 86.368 87.426 86.472 91.8 ; 
      RECT 85.936 87.426 86.04 91.8 ; 
      RECT 85.504 87.426 85.608 91.8 ; 
      RECT 85.072 87.426 85.176 91.8 ; 
      RECT 84.64 87.426 84.744 91.8 ; 
      RECT 84.208 87.426 84.312 91.8 ; 
      RECT 83.776 87.426 83.88 91.8 ; 
      RECT 83.344 87.426 83.448 91.8 ; 
      RECT 82.912 87.426 83.016 91.8 ; 
      RECT 82.48 87.426 82.584 91.8 ; 
      RECT 82.048 87.426 82.152 91.8 ; 
      RECT 81.616 87.426 81.72 91.8 ; 
      RECT 81.184 87.426 81.288 91.8 ; 
      RECT 80.752 87.426 80.856 91.8 ; 
      RECT 80.32 87.426 80.424 91.8 ; 
      RECT 79.888 87.426 79.992 91.8 ; 
      RECT 79.456 87.426 79.56 91.8 ; 
      RECT 79.024 87.426 79.128 91.8 ; 
      RECT 78.592 87.426 78.696 91.8 ; 
      RECT 78.16 87.426 78.264 91.8 ; 
      RECT 77.728 87.426 77.832 91.8 ; 
      RECT 77.296 87.426 77.4 91.8 ; 
      RECT 76.864 87.426 76.968 91.8 ; 
      RECT 76.432 87.426 76.536 91.8 ; 
      RECT 76 87.426 76.104 91.8 ; 
      RECT 75.568 87.426 75.672 91.8 ; 
      RECT 75.136 87.426 75.24 91.8 ; 
      RECT 74.704 87.426 74.808 91.8 ; 
      RECT 74.272 87.426 74.376 91.8 ; 
      RECT 73.84 87.426 73.944 91.8 ; 
      RECT 73.408 87.426 73.512 91.8 ; 
      RECT 72.976 87.426 73.08 91.8 ; 
      RECT 72.544 87.426 72.648 91.8 ; 
      RECT 72.112 87.426 72.216 91.8 ; 
      RECT 71.68 87.426 71.784 91.8 ; 
      RECT 71.248 87.426 71.352 91.8 ; 
      RECT 70.816 87.426 70.92 91.8 ; 
      RECT 70.384 87.426 70.488 91.8 ; 
      RECT 69.952 87.426 70.056 91.8 ; 
      RECT 69.52 87.426 69.624 91.8 ; 
      RECT 69.088 87.426 69.192 91.8 ; 
      RECT 68.656 87.426 68.76 91.8 ; 
      RECT 68.224 87.426 68.328 91.8 ; 
      RECT 67.792 87.426 67.896 91.8 ; 
      RECT 67.36 87.426 67.464 91.8 ; 
      RECT 66.928 87.426 67.032 91.8 ; 
      RECT 66.496 87.426 66.6 91.8 ; 
      RECT 66.064 87.426 66.168 91.8 ; 
      RECT 65.632 87.426 65.736 91.8 ; 
      RECT 65.2 87.426 65.304 91.8 ; 
      RECT 64.348 87.426 64.656 91.8 ; 
      RECT 56.776 87.426 57.084 91.8 ; 
      RECT 56.128 87.426 56.232 91.8 ; 
      RECT 55.696 87.426 55.8 91.8 ; 
      RECT 55.264 87.426 55.368 91.8 ; 
      RECT 54.832 87.426 54.936 91.8 ; 
      RECT 54.4 87.426 54.504 91.8 ; 
      RECT 53.968 87.426 54.072 91.8 ; 
      RECT 53.536 87.426 53.64 91.8 ; 
      RECT 53.104 87.426 53.208 91.8 ; 
      RECT 52.672 87.426 52.776 91.8 ; 
      RECT 52.24 87.426 52.344 91.8 ; 
      RECT 51.808 87.426 51.912 91.8 ; 
      RECT 51.376 87.426 51.48 91.8 ; 
      RECT 50.944 87.426 51.048 91.8 ; 
      RECT 50.512 87.426 50.616 91.8 ; 
      RECT 50.08 87.426 50.184 91.8 ; 
      RECT 49.648 87.426 49.752 91.8 ; 
      RECT 49.216 87.426 49.32 91.8 ; 
      RECT 48.784 87.426 48.888 91.8 ; 
      RECT 48.352 87.426 48.456 91.8 ; 
      RECT 47.92 87.426 48.024 91.8 ; 
      RECT 47.488 87.426 47.592 91.8 ; 
      RECT 47.056 87.426 47.16 91.8 ; 
      RECT 46.624 87.426 46.728 91.8 ; 
      RECT 46.192 87.426 46.296 91.8 ; 
      RECT 45.76 87.426 45.864 91.8 ; 
      RECT 45.328 87.426 45.432 91.8 ; 
      RECT 44.896 87.426 45 91.8 ; 
      RECT 44.464 87.426 44.568 91.8 ; 
      RECT 44.032 87.426 44.136 91.8 ; 
      RECT 43.6 87.426 43.704 91.8 ; 
      RECT 43.168 87.426 43.272 91.8 ; 
      RECT 42.736 87.426 42.84 91.8 ; 
      RECT 42.304 87.426 42.408 91.8 ; 
      RECT 41.872 87.426 41.976 91.8 ; 
      RECT 41.44 87.426 41.544 91.8 ; 
      RECT 41.008 87.426 41.112 91.8 ; 
      RECT 40.576 87.426 40.68 91.8 ; 
      RECT 40.144 87.426 40.248 91.8 ; 
      RECT 39.712 87.426 39.816 91.8 ; 
      RECT 39.28 87.426 39.384 91.8 ; 
      RECT 38.848 87.426 38.952 91.8 ; 
      RECT 38.416 87.426 38.52 91.8 ; 
      RECT 37.984 87.426 38.088 91.8 ; 
      RECT 37.552 87.426 37.656 91.8 ; 
      RECT 37.12 87.426 37.224 91.8 ; 
      RECT 36.688 87.426 36.792 91.8 ; 
      RECT 36.256 87.426 36.36 91.8 ; 
      RECT 35.824 87.426 35.928 91.8 ; 
      RECT 35.392 87.426 35.496 91.8 ; 
      RECT 34.96 87.426 35.064 91.8 ; 
      RECT 34.528 87.426 34.632 91.8 ; 
      RECT 34.096 87.426 34.2 91.8 ; 
      RECT 33.664 87.426 33.768 91.8 ; 
      RECT 33.232 87.426 33.336 91.8 ; 
      RECT 32.8 87.426 32.904 91.8 ; 
      RECT 32.368 87.426 32.472 91.8 ; 
      RECT 31.936 87.426 32.04 91.8 ; 
      RECT 31.504 87.426 31.608 91.8 ; 
      RECT 31.072 87.426 31.176 91.8 ; 
      RECT 30.64 87.426 30.744 91.8 ; 
      RECT 30.208 87.426 30.312 91.8 ; 
      RECT 29.776 87.426 29.88 91.8 ; 
      RECT 29.344 87.426 29.448 91.8 ; 
      RECT 28.912 87.426 29.016 91.8 ; 
      RECT 28.48 87.426 28.584 91.8 ; 
      RECT 28.048 87.426 28.152 91.8 ; 
      RECT 27.616 87.426 27.72 91.8 ; 
      RECT 27.184 87.426 27.288 91.8 ; 
      RECT 26.752 87.426 26.856 91.8 ; 
      RECT 26.32 87.426 26.424 91.8 ; 
      RECT 25.888 87.426 25.992 91.8 ; 
      RECT 25.456 87.426 25.56 91.8 ; 
      RECT 25.024 87.426 25.128 91.8 ; 
      RECT 24.592 87.426 24.696 91.8 ; 
      RECT 24.16 87.426 24.264 91.8 ; 
      RECT 23.728 87.426 23.832 91.8 ; 
      RECT 23.296 87.426 23.4 91.8 ; 
      RECT 22.864 87.426 22.968 91.8 ; 
      RECT 22.432 87.426 22.536 91.8 ; 
      RECT 22 87.426 22.104 91.8 ; 
      RECT 21.568 87.426 21.672 91.8 ; 
      RECT 21.136 87.426 21.24 91.8 ; 
      RECT 20.704 87.426 20.808 91.8 ; 
      RECT 20.272 87.426 20.376 91.8 ; 
      RECT 19.84 87.426 19.944 91.8 ; 
      RECT 19.408 87.426 19.512 91.8 ; 
      RECT 18.976 87.426 19.08 91.8 ; 
      RECT 18.544 87.426 18.648 91.8 ; 
      RECT 18.112 87.426 18.216 91.8 ; 
      RECT 17.68 87.426 17.784 91.8 ; 
      RECT 17.248 87.426 17.352 91.8 ; 
      RECT 16.816 87.426 16.92 91.8 ; 
      RECT 16.384 87.426 16.488 91.8 ; 
      RECT 15.952 87.426 16.056 91.8 ; 
      RECT 15.52 87.426 15.624 91.8 ; 
      RECT 15.088 87.426 15.192 91.8 ; 
      RECT 14.656 87.426 14.76 91.8 ; 
      RECT 14.224 87.426 14.328 91.8 ; 
      RECT 13.792 87.426 13.896 91.8 ; 
      RECT 13.36 87.426 13.464 91.8 ; 
      RECT 12.928 87.426 13.032 91.8 ; 
      RECT 12.496 87.426 12.6 91.8 ; 
      RECT 12.064 87.426 12.168 91.8 ; 
      RECT 11.632 87.426 11.736 91.8 ; 
      RECT 11.2 87.426 11.304 91.8 ; 
      RECT 10.768 87.426 10.872 91.8 ; 
      RECT 10.336 87.426 10.44 91.8 ; 
      RECT 9.904 87.426 10.008 91.8 ; 
      RECT 9.472 87.426 9.576 91.8 ; 
      RECT 9.04 87.426 9.144 91.8 ; 
      RECT 8.608 87.426 8.712 91.8 ; 
      RECT 8.176 87.426 8.28 91.8 ; 
      RECT 7.744 87.426 7.848 91.8 ; 
      RECT 7.312 87.426 7.416 91.8 ; 
      RECT 6.88 87.426 6.984 91.8 ; 
      RECT 6.448 87.426 6.552 91.8 ; 
      RECT 6.016 87.426 6.12 91.8 ; 
      RECT 5.584 87.426 5.688 91.8 ; 
      RECT 5.152 87.426 5.256 91.8 ; 
      RECT 4.72 87.426 4.824 91.8 ; 
      RECT 4.288 87.426 4.392 91.8 ; 
      RECT 3.856 87.426 3.96 91.8 ; 
      RECT 3.424 87.426 3.528 91.8 ; 
      RECT 2.992 87.426 3.096 91.8 ; 
      RECT 2.56 87.426 2.664 91.8 ; 
      RECT 2.128 87.426 2.232 91.8 ; 
      RECT 1.696 87.426 1.8 91.8 ; 
      RECT 1.264 87.426 1.368 91.8 ; 
      RECT 0.832 87.426 0.936 91.8 ; 
      RECT 0.02 87.426 0.36 91.8 ; 
      RECT 62.212 91.746 62.724 96.12 ; 
      RECT 62.156 94.408 62.724 95.698 ; 
      RECT 61.276 93.316 61.812 96.12 ; 
      RECT 61.184 94.656 61.812 95.688 ; 
      RECT 61.276 91.746 61.668 96.12 ; 
      RECT 61.276 92.23 61.724 93.188 ; 
      RECT 61.276 91.746 61.812 92.102 ; 
      RECT 60.376 93.548 60.912 96.12 ; 
      RECT 60.376 91.746 60.768 96.12 ; 
      RECT 58.708 91.746 59.04 96.12 ; 
      RECT 58.708 92.1 59.096 95.842 ; 
      RECT 121.072 91.746 121.412 96.12 ; 
      RECT 120.496 91.746 120.6 96.12 ; 
      RECT 120.064 91.746 120.168 96.12 ; 
      RECT 119.632 91.746 119.736 96.12 ; 
      RECT 119.2 91.746 119.304 96.12 ; 
      RECT 118.768 91.746 118.872 96.12 ; 
      RECT 118.336 91.746 118.44 96.12 ; 
      RECT 117.904 91.746 118.008 96.12 ; 
      RECT 117.472 91.746 117.576 96.12 ; 
      RECT 117.04 91.746 117.144 96.12 ; 
      RECT 116.608 91.746 116.712 96.12 ; 
      RECT 116.176 91.746 116.28 96.12 ; 
      RECT 115.744 91.746 115.848 96.12 ; 
      RECT 115.312 91.746 115.416 96.12 ; 
      RECT 114.88 91.746 114.984 96.12 ; 
      RECT 114.448 91.746 114.552 96.12 ; 
      RECT 114.016 91.746 114.12 96.12 ; 
      RECT 113.584 91.746 113.688 96.12 ; 
      RECT 113.152 91.746 113.256 96.12 ; 
      RECT 112.72 91.746 112.824 96.12 ; 
      RECT 112.288 91.746 112.392 96.12 ; 
      RECT 111.856 91.746 111.96 96.12 ; 
      RECT 111.424 91.746 111.528 96.12 ; 
      RECT 110.992 91.746 111.096 96.12 ; 
      RECT 110.56 91.746 110.664 96.12 ; 
      RECT 110.128 91.746 110.232 96.12 ; 
      RECT 109.696 91.746 109.8 96.12 ; 
      RECT 109.264 91.746 109.368 96.12 ; 
      RECT 108.832 91.746 108.936 96.12 ; 
      RECT 108.4 91.746 108.504 96.12 ; 
      RECT 107.968 91.746 108.072 96.12 ; 
      RECT 107.536 91.746 107.64 96.12 ; 
      RECT 107.104 91.746 107.208 96.12 ; 
      RECT 106.672 91.746 106.776 96.12 ; 
      RECT 106.24 91.746 106.344 96.12 ; 
      RECT 105.808 91.746 105.912 96.12 ; 
      RECT 105.376 91.746 105.48 96.12 ; 
      RECT 104.944 91.746 105.048 96.12 ; 
      RECT 104.512 91.746 104.616 96.12 ; 
      RECT 104.08 91.746 104.184 96.12 ; 
      RECT 103.648 91.746 103.752 96.12 ; 
      RECT 103.216 91.746 103.32 96.12 ; 
      RECT 102.784 91.746 102.888 96.12 ; 
      RECT 102.352 91.746 102.456 96.12 ; 
      RECT 101.92 91.746 102.024 96.12 ; 
      RECT 101.488 91.746 101.592 96.12 ; 
      RECT 101.056 91.746 101.16 96.12 ; 
      RECT 100.624 91.746 100.728 96.12 ; 
      RECT 100.192 91.746 100.296 96.12 ; 
      RECT 99.76 91.746 99.864 96.12 ; 
      RECT 99.328 91.746 99.432 96.12 ; 
      RECT 98.896 91.746 99 96.12 ; 
      RECT 98.464 91.746 98.568 96.12 ; 
      RECT 98.032 91.746 98.136 96.12 ; 
      RECT 97.6 91.746 97.704 96.12 ; 
      RECT 97.168 91.746 97.272 96.12 ; 
      RECT 96.736 91.746 96.84 96.12 ; 
      RECT 96.304 91.746 96.408 96.12 ; 
      RECT 95.872 91.746 95.976 96.12 ; 
      RECT 95.44 91.746 95.544 96.12 ; 
      RECT 95.008 91.746 95.112 96.12 ; 
      RECT 94.576 91.746 94.68 96.12 ; 
      RECT 94.144 91.746 94.248 96.12 ; 
      RECT 93.712 91.746 93.816 96.12 ; 
      RECT 93.28 91.746 93.384 96.12 ; 
      RECT 92.848 91.746 92.952 96.12 ; 
      RECT 92.416 91.746 92.52 96.12 ; 
      RECT 91.984 91.746 92.088 96.12 ; 
      RECT 91.552 91.746 91.656 96.12 ; 
      RECT 91.12 91.746 91.224 96.12 ; 
      RECT 90.688 91.746 90.792 96.12 ; 
      RECT 90.256 91.746 90.36 96.12 ; 
      RECT 89.824 91.746 89.928 96.12 ; 
      RECT 89.392 91.746 89.496 96.12 ; 
      RECT 88.96 91.746 89.064 96.12 ; 
      RECT 88.528 91.746 88.632 96.12 ; 
      RECT 88.096 91.746 88.2 96.12 ; 
      RECT 87.664 91.746 87.768 96.12 ; 
      RECT 87.232 91.746 87.336 96.12 ; 
      RECT 86.8 91.746 86.904 96.12 ; 
      RECT 86.368 91.746 86.472 96.12 ; 
      RECT 85.936 91.746 86.04 96.12 ; 
      RECT 85.504 91.746 85.608 96.12 ; 
      RECT 85.072 91.746 85.176 96.12 ; 
      RECT 84.64 91.746 84.744 96.12 ; 
      RECT 84.208 91.746 84.312 96.12 ; 
      RECT 83.776 91.746 83.88 96.12 ; 
      RECT 83.344 91.746 83.448 96.12 ; 
      RECT 82.912 91.746 83.016 96.12 ; 
      RECT 82.48 91.746 82.584 96.12 ; 
      RECT 82.048 91.746 82.152 96.12 ; 
      RECT 81.616 91.746 81.72 96.12 ; 
      RECT 81.184 91.746 81.288 96.12 ; 
      RECT 80.752 91.746 80.856 96.12 ; 
      RECT 80.32 91.746 80.424 96.12 ; 
      RECT 79.888 91.746 79.992 96.12 ; 
      RECT 79.456 91.746 79.56 96.12 ; 
      RECT 79.024 91.746 79.128 96.12 ; 
      RECT 78.592 91.746 78.696 96.12 ; 
      RECT 78.16 91.746 78.264 96.12 ; 
      RECT 77.728 91.746 77.832 96.12 ; 
      RECT 77.296 91.746 77.4 96.12 ; 
      RECT 76.864 91.746 76.968 96.12 ; 
      RECT 76.432 91.746 76.536 96.12 ; 
      RECT 76 91.746 76.104 96.12 ; 
      RECT 75.568 91.746 75.672 96.12 ; 
      RECT 75.136 91.746 75.24 96.12 ; 
      RECT 74.704 91.746 74.808 96.12 ; 
      RECT 74.272 91.746 74.376 96.12 ; 
      RECT 73.84 91.746 73.944 96.12 ; 
      RECT 73.408 91.746 73.512 96.12 ; 
      RECT 72.976 91.746 73.08 96.12 ; 
      RECT 72.544 91.746 72.648 96.12 ; 
      RECT 72.112 91.746 72.216 96.12 ; 
      RECT 71.68 91.746 71.784 96.12 ; 
      RECT 71.248 91.746 71.352 96.12 ; 
      RECT 70.816 91.746 70.92 96.12 ; 
      RECT 70.384 91.746 70.488 96.12 ; 
      RECT 69.952 91.746 70.056 96.12 ; 
      RECT 69.52 91.746 69.624 96.12 ; 
      RECT 69.088 91.746 69.192 96.12 ; 
      RECT 68.656 91.746 68.76 96.12 ; 
      RECT 68.224 91.746 68.328 96.12 ; 
      RECT 67.792 91.746 67.896 96.12 ; 
      RECT 67.36 91.746 67.464 96.12 ; 
      RECT 66.928 91.746 67.032 96.12 ; 
      RECT 66.496 91.746 66.6 96.12 ; 
      RECT 66.064 91.746 66.168 96.12 ; 
      RECT 65.632 91.746 65.736 96.12 ; 
      RECT 65.2 91.746 65.304 96.12 ; 
      RECT 64.348 91.746 64.656 96.12 ; 
      RECT 56.776 91.746 57.084 96.12 ; 
      RECT 56.128 91.746 56.232 96.12 ; 
      RECT 55.696 91.746 55.8 96.12 ; 
      RECT 55.264 91.746 55.368 96.12 ; 
      RECT 54.832 91.746 54.936 96.12 ; 
      RECT 54.4 91.746 54.504 96.12 ; 
      RECT 53.968 91.746 54.072 96.12 ; 
      RECT 53.536 91.746 53.64 96.12 ; 
      RECT 53.104 91.746 53.208 96.12 ; 
      RECT 52.672 91.746 52.776 96.12 ; 
      RECT 52.24 91.746 52.344 96.12 ; 
      RECT 51.808 91.746 51.912 96.12 ; 
      RECT 51.376 91.746 51.48 96.12 ; 
      RECT 50.944 91.746 51.048 96.12 ; 
      RECT 50.512 91.746 50.616 96.12 ; 
      RECT 50.08 91.746 50.184 96.12 ; 
      RECT 49.648 91.746 49.752 96.12 ; 
      RECT 49.216 91.746 49.32 96.12 ; 
      RECT 48.784 91.746 48.888 96.12 ; 
      RECT 48.352 91.746 48.456 96.12 ; 
      RECT 47.92 91.746 48.024 96.12 ; 
      RECT 47.488 91.746 47.592 96.12 ; 
      RECT 47.056 91.746 47.16 96.12 ; 
      RECT 46.624 91.746 46.728 96.12 ; 
      RECT 46.192 91.746 46.296 96.12 ; 
      RECT 45.76 91.746 45.864 96.12 ; 
      RECT 45.328 91.746 45.432 96.12 ; 
      RECT 44.896 91.746 45 96.12 ; 
      RECT 44.464 91.746 44.568 96.12 ; 
      RECT 44.032 91.746 44.136 96.12 ; 
      RECT 43.6 91.746 43.704 96.12 ; 
      RECT 43.168 91.746 43.272 96.12 ; 
      RECT 42.736 91.746 42.84 96.12 ; 
      RECT 42.304 91.746 42.408 96.12 ; 
      RECT 41.872 91.746 41.976 96.12 ; 
      RECT 41.44 91.746 41.544 96.12 ; 
      RECT 41.008 91.746 41.112 96.12 ; 
      RECT 40.576 91.746 40.68 96.12 ; 
      RECT 40.144 91.746 40.248 96.12 ; 
      RECT 39.712 91.746 39.816 96.12 ; 
      RECT 39.28 91.746 39.384 96.12 ; 
      RECT 38.848 91.746 38.952 96.12 ; 
      RECT 38.416 91.746 38.52 96.12 ; 
      RECT 37.984 91.746 38.088 96.12 ; 
      RECT 37.552 91.746 37.656 96.12 ; 
      RECT 37.12 91.746 37.224 96.12 ; 
      RECT 36.688 91.746 36.792 96.12 ; 
      RECT 36.256 91.746 36.36 96.12 ; 
      RECT 35.824 91.746 35.928 96.12 ; 
      RECT 35.392 91.746 35.496 96.12 ; 
      RECT 34.96 91.746 35.064 96.12 ; 
      RECT 34.528 91.746 34.632 96.12 ; 
      RECT 34.096 91.746 34.2 96.12 ; 
      RECT 33.664 91.746 33.768 96.12 ; 
      RECT 33.232 91.746 33.336 96.12 ; 
      RECT 32.8 91.746 32.904 96.12 ; 
      RECT 32.368 91.746 32.472 96.12 ; 
      RECT 31.936 91.746 32.04 96.12 ; 
      RECT 31.504 91.746 31.608 96.12 ; 
      RECT 31.072 91.746 31.176 96.12 ; 
      RECT 30.64 91.746 30.744 96.12 ; 
      RECT 30.208 91.746 30.312 96.12 ; 
      RECT 29.776 91.746 29.88 96.12 ; 
      RECT 29.344 91.746 29.448 96.12 ; 
      RECT 28.912 91.746 29.016 96.12 ; 
      RECT 28.48 91.746 28.584 96.12 ; 
      RECT 28.048 91.746 28.152 96.12 ; 
      RECT 27.616 91.746 27.72 96.12 ; 
      RECT 27.184 91.746 27.288 96.12 ; 
      RECT 26.752 91.746 26.856 96.12 ; 
      RECT 26.32 91.746 26.424 96.12 ; 
      RECT 25.888 91.746 25.992 96.12 ; 
      RECT 25.456 91.746 25.56 96.12 ; 
      RECT 25.024 91.746 25.128 96.12 ; 
      RECT 24.592 91.746 24.696 96.12 ; 
      RECT 24.16 91.746 24.264 96.12 ; 
      RECT 23.728 91.746 23.832 96.12 ; 
      RECT 23.296 91.746 23.4 96.12 ; 
      RECT 22.864 91.746 22.968 96.12 ; 
      RECT 22.432 91.746 22.536 96.12 ; 
      RECT 22 91.746 22.104 96.12 ; 
      RECT 21.568 91.746 21.672 96.12 ; 
      RECT 21.136 91.746 21.24 96.12 ; 
      RECT 20.704 91.746 20.808 96.12 ; 
      RECT 20.272 91.746 20.376 96.12 ; 
      RECT 19.84 91.746 19.944 96.12 ; 
      RECT 19.408 91.746 19.512 96.12 ; 
      RECT 18.976 91.746 19.08 96.12 ; 
      RECT 18.544 91.746 18.648 96.12 ; 
      RECT 18.112 91.746 18.216 96.12 ; 
      RECT 17.68 91.746 17.784 96.12 ; 
      RECT 17.248 91.746 17.352 96.12 ; 
      RECT 16.816 91.746 16.92 96.12 ; 
      RECT 16.384 91.746 16.488 96.12 ; 
      RECT 15.952 91.746 16.056 96.12 ; 
      RECT 15.52 91.746 15.624 96.12 ; 
      RECT 15.088 91.746 15.192 96.12 ; 
      RECT 14.656 91.746 14.76 96.12 ; 
      RECT 14.224 91.746 14.328 96.12 ; 
      RECT 13.792 91.746 13.896 96.12 ; 
      RECT 13.36 91.746 13.464 96.12 ; 
      RECT 12.928 91.746 13.032 96.12 ; 
      RECT 12.496 91.746 12.6 96.12 ; 
      RECT 12.064 91.746 12.168 96.12 ; 
      RECT 11.632 91.746 11.736 96.12 ; 
      RECT 11.2 91.746 11.304 96.12 ; 
      RECT 10.768 91.746 10.872 96.12 ; 
      RECT 10.336 91.746 10.44 96.12 ; 
      RECT 9.904 91.746 10.008 96.12 ; 
      RECT 9.472 91.746 9.576 96.12 ; 
      RECT 9.04 91.746 9.144 96.12 ; 
      RECT 8.608 91.746 8.712 96.12 ; 
      RECT 8.176 91.746 8.28 96.12 ; 
      RECT 7.744 91.746 7.848 96.12 ; 
      RECT 7.312 91.746 7.416 96.12 ; 
      RECT 6.88 91.746 6.984 96.12 ; 
      RECT 6.448 91.746 6.552 96.12 ; 
      RECT 6.016 91.746 6.12 96.12 ; 
      RECT 5.584 91.746 5.688 96.12 ; 
      RECT 5.152 91.746 5.256 96.12 ; 
      RECT 4.72 91.746 4.824 96.12 ; 
      RECT 4.288 91.746 4.392 96.12 ; 
      RECT 3.856 91.746 3.96 96.12 ; 
      RECT 3.424 91.746 3.528 96.12 ; 
      RECT 2.992 91.746 3.096 96.12 ; 
      RECT 2.56 91.746 2.664 96.12 ; 
      RECT 2.128 91.746 2.232 96.12 ; 
      RECT 1.696 91.746 1.8 96.12 ; 
      RECT 1.264 91.746 1.368 96.12 ; 
      RECT 0.832 91.746 0.936 96.12 ; 
      RECT 0.02 91.746 0.36 96.12 ; 
      RECT 62.212 96.066 62.724 100.44 ; 
      RECT 62.156 98.728 62.724 100.018 ; 
      RECT 61.276 97.636 61.812 100.44 ; 
      RECT 61.184 98.976 61.812 100.008 ; 
      RECT 61.276 96.066 61.668 100.44 ; 
      RECT 61.276 96.55 61.724 97.508 ; 
      RECT 61.276 96.066 61.812 96.422 ; 
      RECT 60.376 97.868 60.912 100.44 ; 
      RECT 60.376 96.066 60.768 100.44 ; 
      RECT 58.708 96.066 59.04 100.44 ; 
      RECT 58.708 96.42 59.096 100.162 ; 
      RECT 121.072 96.066 121.412 100.44 ; 
      RECT 120.496 96.066 120.6 100.44 ; 
      RECT 120.064 96.066 120.168 100.44 ; 
      RECT 119.632 96.066 119.736 100.44 ; 
      RECT 119.2 96.066 119.304 100.44 ; 
      RECT 118.768 96.066 118.872 100.44 ; 
      RECT 118.336 96.066 118.44 100.44 ; 
      RECT 117.904 96.066 118.008 100.44 ; 
      RECT 117.472 96.066 117.576 100.44 ; 
      RECT 117.04 96.066 117.144 100.44 ; 
      RECT 116.608 96.066 116.712 100.44 ; 
      RECT 116.176 96.066 116.28 100.44 ; 
      RECT 115.744 96.066 115.848 100.44 ; 
      RECT 115.312 96.066 115.416 100.44 ; 
      RECT 114.88 96.066 114.984 100.44 ; 
      RECT 114.448 96.066 114.552 100.44 ; 
      RECT 114.016 96.066 114.12 100.44 ; 
      RECT 113.584 96.066 113.688 100.44 ; 
      RECT 113.152 96.066 113.256 100.44 ; 
      RECT 112.72 96.066 112.824 100.44 ; 
      RECT 112.288 96.066 112.392 100.44 ; 
      RECT 111.856 96.066 111.96 100.44 ; 
      RECT 111.424 96.066 111.528 100.44 ; 
      RECT 110.992 96.066 111.096 100.44 ; 
      RECT 110.56 96.066 110.664 100.44 ; 
      RECT 110.128 96.066 110.232 100.44 ; 
      RECT 109.696 96.066 109.8 100.44 ; 
      RECT 109.264 96.066 109.368 100.44 ; 
      RECT 108.832 96.066 108.936 100.44 ; 
      RECT 108.4 96.066 108.504 100.44 ; 
      RECT 107.968 96.066 108.072 100.44 ; 
      RECT 107.536 96.066 107.64 100.44 ; 
      RECT 107.104 96.066 107.208 100.44 ; 
      RECT 106.672 96.066 106.776 100.44 ; 
      RECT 106.24 96.066 106.344 100.44 ; 
      RECT 105.808 96.066 105.912 100.44 ; 
      RECT 105.376 96.066 105.48 100.44 ; 
      RECT 104.944 96.066 105.048 100.44 ; 
      RECT 104.512 96.066 104.616 100.44 ; 
      RECT 104.08 96.066 104.184 100.44 ; 
      RECT 103.648 96.066 103.752 100.44 ; 
      RECT 103.216 96.066 103.32 100.44 ; 
      RECT 102.784 96.066 102.888 100.44 ; 
      RECT 102.352 96.066 102.456 100.44 ; 
      RECT 101.92 96.066 102.024 100.44 ; 
      RECT 101.488 96.066 101.592 100.44 ; 
      RECT 101.056 96.066 101.16 100.44 ; 
      RECT 100.624 96.066 100.728 100.44 ; 
      RECT 100.192 96.066 100.296 100.44 ; 
      RECT 99.76 96.066 99.864 100.44 ; 
      RECT 99.328 96.066 99.432 100.44 ; 
      RECT 98.896 96.066 99 100.44 ; 
      RECT 98.464 96.066 98.568 100.44 ; 
      RECT 98.032 96.066 98.136 100.44 ; 
      RECT 97.6 96.066 97.704 100.44 ; 
      RECT 97.168 96.066 97.272 100.44 ; 
      RECT 96.736 96.066 96.84 100.44 ; 
      RECT 96.304 96.066 96.408 100.44 ; 
      RECT 95.872 96.066 95.976 100.44 ; 
      RECT 95.44 96.066 95.544 100.44 ; 
      RECT 95.008 96.066 95.112 100.44 ; 
      RECT 94.576 96.066 94.68 100.44 ; 
      RECT 94.144 96.066 94.248 100.44 ; 
      RECT 93.712 96.066 93.816 100.44 ; 
      RECT 93.28 96.066 93.384 100.44 ; 
      RECT 92.848 96.066 92.952 100.44 ; 
      RECT 92.416 96.066 92.52 100.44 ; 
      RECT 91.984 96.066 92.088 100.44 ; 
      RECT 91.552 96.066 91.656 100.44 ; 
      RECT 91.12 96.066 91.224 100.44 ; 
      RECT 90.688 96.066 90.792 100.44 ; 
      RECT 90.256 96.066 90.36 100.44 ; 
      RECT 89.824 96.066 89.928 100.44 ; 
      RECT 89.392 96.066 89.496 100.44 ; 
      RECT 88.96 96.066 89.064 100.44 ; 
      RECT 88.528 96.066 88.632 100.44 ; 
      RECT 88.096 96.066 88.2 100.44 ; 
      RECT 87.664 96.066 87.768 100.44 ; 
      RECT 87.232 96.066 87.336 100.44 ; 
      RECT 86.8 96.066 86.904 100.44 ; 
      RECT 86.368 96.066 86.472 100.44 ; 
      RECT 85.936 96.066 86.04 100.44 ; 
      RECT 85.504 96.066 85.608 100.44 ; 
      RECT 85.072 96.066 85.176 100.44 ; 
      RECT 84.64 96.066 84.744 100.44 ; 
      RECT 84.208 96.066 84.312 100.44 ; 
      RECT 83.776 96.066 83.88 100.44 ; 
      RECT 83.344 96.066 83.448 100.44 ; 
      RECT 82.912 96.066 83.016 100.44 ; 
      RECT 82.48 96.066 82.584 100.44 ; 
      RECT 82.048 96.066 82.152 100.44 ; 
      RECT 81.616 96.066 81.72 100.44 ; 
      RECT 81.184 96.066 81.288 100.44 ; 
      RECT 80.752 96.066 80.856 100.44 ; 
      RECT 80.32 96.066 80.424 100.44 ; 
      RECT 79.888 96.066 79.992 100.44 ; 
      RECT 79.456 96.066 79.56 100.44 ; 
      RECT 79.024 96.066 79.128 100.44 ; 
      RECT 78.592 96.066 78.696 100.44 ; 
      RECT 78.16 96.066 78.264 100.44 ; 
      RECT 77.728 96.066 77.832 100.44 ; 
      RECT 77.296 96.066 77.4 100.44 ; 
      RECT 76.864 96.066 76.968 100.44 ; 
      RECT 76.432 96.066 76.536 100.44 ; 
      RECT 76 96.066 76.104 100.44 ; 
      RECT 75.568 96.066 75.672 100.44 ; 
      RECT 75.136 96.066 75.24 100.44 ; 
      RECT 74.704 96.066 74.808 100.44 ; 
      RECT 74.272 96.066 74.376 100.44 ; 
      RECT 73.84 96.066 73.944 100.44 ; 
      RECT 73.408 96.066 73.512 100.44 ; 
      RECT 72.976 96.066 73.08 100.44 ; 
      RECT 72.544 96.066 72.648 100.44 ; 
      RECT 72.112 96.066 72.216 100.44 ; 
      RECT 71.68 96.066 71.784 100.44 ; 
      RECT 71.248 96.066 71.352 100.44 ; 
      RECT 70.816 96.066 70.92 100.44 ; 
      RECT 70.384 96.066 70.488 100.44 ; 
      RECT 69.952 96.066 70.056 100.44 ; 
      RECT 69.52 96.066 69.624 100.44 ; 
      RECT 69.088 96.066 69.192 100.44 ; 
      RECT 68.656 96.066 68.76 100.44 ; 
      RECT 68.224 96.066 68.328 100.44 ; 
      RECT 67.792 96.066 67.896 100.44 ; 
      RECT 67.36 96.066 67.464 100.44 ; 
      RECT 66.928 96.066 67.032 100.44 ; 
      RECT 66.496 96.066 66.6 100.44 ; 
      RECT 66.064 96.066 66.168 100.44 ; 
      RECT 65.632 96.066 65.736 100.44 ; 
      RECT 65.2 96.066 65.304 100.44 ; 
      RECT 64.348 96.066 64.656 100.44 ; 
      RECT 56.776 96.066 57.084 100.44 ; 
      RECT 56.128 96.066 56.232 100.44 ; 
      RECT 55.696 96.066 55.8 100.44 ; 
      RECT 55.264 96.066 55.368 100.44 ; 
      RECT 54.832 96.066 54.936 100.44 ; 
      RECT 54.4 96.066 54.504 100.44 ; 
      RECT 53.968 96.066 54.072 100.44 ; 
      RECT 53.536 96.066 53.64 100.44 ; 
      RECT 53.104 96.066 53.208 100.44 ; 
      RECT 52.672 96.066 52.776 100.44 ; 
      RECT 52.24 96.066 52.344 100.44 ; 
      RECT 51.808 96.066 51.912 100.44 ; 
      RECT 51.376 96.066 51.48 100.44 ; 
      RECT 50.944 96.066 51.048 100.44 ; 
      RECT 50.512 96.066 50.616 100.44 ; 
      RECT 50.08 96.066 50.184 100.44 ; 
      RECT 49.648 96.066 49.752 100.44 ; 
      RECT 49.216 96.066 49.32 100.44 ; 
      RECT 48.784 96.066 48.888 100.44 ; 
      RECT 48.352 96.066 48.456 100.44 ; 
      RECT 47.92 96.066 48.024 100.44 ; 
      RECT 47.488 96.066 47.592 100.44 ; 
      RECT 47.056 96.066 47.16 100.44 ; 
      RECT 46.624 96.066 46.728 100.44 ; 
      RECT 46.192 96.066 46.296 100.44 ; 
      RECT 45.76 96.066 45.864 100.44 ; 
      RECT 45.328 96.066 45.432 100.44 ; 
      RECT 44.896 96.066 45 100.44 ; 
      RECT 44.464 96.066 44.568 100.44 ; 
      RECT 44.032 96.066 44.136 100.44 ; 
      RECT 43.6 96.066 43.704 100.44 ; 
      RECT 43.168 96.066 43.272 100.44 ; 
      RECT 42.736 96.066 42.84 100.44 ; 
      RECT 42.304 96.066 42.408 100.44 ; 
      RECT 41.872 96.066 41.976 100.44 ; 
      RECT 41.44 96.066 41.544 100.44 ; 
      RECT 41.008 96.066 41.112 100.44 ; 
      RECT 40.576 96.066 40.68 100.44 ; 
      RECT 40.144 96.066 40.248 100.44 ; 
      RECT 39.712 96.066 39.816 100.44 ; 
      RECT 39.28 96.066 39.384 100.44 ; 
      RECT 38.848 96.066 38.952 100.44 ; 
      RECT 38.416 96.066 38.52 100.44 ; 
      RECT 37.984 96.066 38.088 100.44 ; 
      RECT 37.552 96.066 37.656 100.44 ; 
      RECT 37.12 96.066 37.224 100.44 ; 
      RECT 36.688 96.066 36.792 100.44 ; 
      RECT 36.256 96.066 36.36 100.44 ; 
      RECT 35.824 96.066 35.928 100.44 ; 
      RECT 35.392 96.066 35.496 100.44 ; 
      RECT 34.96 96.066 35.064 100.44 ; 
      RECT 34.528 96.066 34.632 100.44 ; 
      RECT 34.096 96.066 34.2 100.44 ; 
      RECT 33.664 96.066 33.768 100.44 ; 
      RECT 33.232 96.066 33.336 100.44 ; 
      RECT 32.8 96.066 32.904 100.44 ; 
      RECT 32.368 96.066 32.472 100.44 ; 
      RECT 31.936 96.066 32.04 100.44 ; 
      RECT 31.504 96.066 31.608 100.44 ; 
      RECT 31.072 96.066 31.176 100.44 ; 
      RECT 30.64 96.066 30.744 100.44 ; 
      RECT 30.208 96.066 30.312 100.44 ; 
      RECT 29.776 96.066 29.88 100.44 ; 
      RECT 29.344 96.066 29.448 100.44 ; 
      RECT 28.912 96.066 29.016 100.44 ; 
      RECT 28.48 96.066 28.584 100.44 ; 
      RECT 28.048 96.066 28.152 100.44 ; 
      RECT 27.616 96.066 27.72 100.44 ; 
      RECT 27.184 96.066 27.288 100.44 ; 
      RECT 26.752 96.066 26.856 100.44 ; 
      RECT 26.32 96.066 26.424 100.44 ; 
      RECT 25.888 96.066 25.992 100.44 ; 
      RECT 25.456 96.066 25.56 100.44 ; 
      RECT 25.024 96.066 25.128 100.44 ; 
      RECT 24.592 96.066 24.696 100.44 ; 
      RECT 24.16 96.066 24.264 100.44 ; 
      RECT 23.728 96.066 23.832 100.44 ; 
      RECT 23.296 96.066 23.4 100.44 ; 
      RECT 22.864 96.066 22.968 100.44 ; 
      RECT 22.432 96.066 22.536 100.44 ; 
      RECT 22 96.066 22.104 100.44 ; 
      RECT 21.568 96.066 21.672 100.44 ; 
      RECT 21.136 96.066 21.24 100.44 ; 
      RECT 20.704 96.066 20.808 100.44 ; 
      RECT 20.272 96.066 20.376 100.44 ; 
      RECT 19.84 96.066 19.944 100.44 ; 
      RECT 19.408 96.066 19.512 100.44 ; 
      RECT 18.976 96.066 19.08 100.44 ; 
      RECT 18.544 96.066 18.648 100.44 ; 
      RECT 18.112 96.066 18.216 100.44 ; 
      RECT 17.68 96.066 17.784 100.44 ; 
      RECT 17.248 96.066 17.352 100.44 ; 
      RECT 16.816 96.066 16.92 100.44 ; 
      RECT 16.384 96.066 16.488 100.44 ; 
      RECT 15.952 96.066 16.056 100.44 ; 
      RECT 15.52 96.066 15.624 100.44 ; 
      RECT 15.088 96.066 15.192 100.44 ; 
      RECT 14.656 96.066 14.76 100.44 ; 
      RECT 14.224 96.066 14.328 100.44 ; 
      RECT 13.792 96.066 13.896 100.44 ; 
      RECT 13.36 96.066 13.464 100.44 ; 
      RECT 12.928 96.066 13.032 100.44 ; 
      RECT 12.496 96.066 12.6 100.44 ; 
      RECT 12.064 96.066 12.168 100.44 ; 
      RECT 11.632 96.066 11.736 100.44 ; 
      RECT 11.2 96.066 11.304 100.44 ; 
      RECT 10.768 96.066 10.872 100.44 ; 
      RECT 10.336 96.066 10.44 100.44 ; 
      RECT 9.904 96.066 10.008 100.44 ; 
      RECT 9.472 96.066 9.576 100.44 ; 
      RECT 9.04 96.066 9.144 100.44 ; 
      RECT 8.608 96.066 8.712 100.44 ; 
      RECT 8.176 96.066 8.28 100.44 ; 
      RECT 7.744 96.066 7.848 100.44 ; 
      RECT 7.312 96.066 7.416 100.44 ; 
      RECT 6.88 96.066 6.984 100.44 ; 
      RECT 6.448 96.066 6.552 100.44 ; 
      RECT 6.016 96.066 6.12 100.44 ; 
      RECT 5.584 96.066 5.688 100.44 ; 
      RECT 5.152 96.066 5.256 100.44 ; 
      RECT 4.72 96.066 4.824 100.44 ; 
      RECT 4.288 96.066 4.392 100.44 ; 
      RECT 3.856 96.066 3.96 100.44 ; 
      RECT 3.424 96.066 3.528 100.44 ; 
      RECT 2.992 96.066 3.096 100.44 ; 
      RECT 2.56 96.066 2.664 100.44 ; 
      RECT 2.128 96.066 2.232 100.44 ; 
      RECT 1.696 96.066 1.8 100.44 ; 
      RECT 1.264 96.066 1.368 100.44 ; 
      RECT 0.832 96.066 0.936 100.44 ; 
      RECT 0.02 96.066 0.36 100.44 ; 
      RECT 62.212 100.386 62.724 104.76 ; 
      RECT 62.156 103.048 62.724 104.338 ; 
      RECT 61.276 101.956 61.812 104.76 ; 
      RECT 61.184 103.296 61.812 104.328 ; 
      RECT 61.276 100.386 61.668 104.76 ; 
      RECT 61.276 100.87 61.724 101.828 ; 
      RECT 61.276 100.386 61.812 100.742 ; 
      RECT 60.376 102.188 60.912 104.76 ; 
      RECT 60.376 100.386 60.768 104.76 ; 
      RECT 58.708 100.386 59.04 104.76 ; 
      RECT 58.708 100.74 59.096 104.482 ; 
      RECT 121.072 100.386 121.412 104.76 ; 
      RECT 120.496 100.386 120.6 104.76 ; 
      RECT 120.064 100.386 120.168 104.76 ; 
      RECT 119.632 100.386 119.736 104.76 ; 
      RECT 119.2 100.386 119.304 104.76 ; 
      RECT 118.768 100.386 118.872 104.76 ; 
      RECT 118.336 100.386 118.44 104.76 ; 
      RECT 117.904 100.386 118.008 104.76 ; 
      RECT 117.472 100.386 117.576 104.76 ; 
      RECT 117.04 100.386 117.144 104.76 ; 
      RECT 116.608 100.386 116.712 104.76 ; 
      RECT 116.176 100.386 116.28 104.76 ; 
      RECT 115.744 100.386 115.848 104.76 ; 
      RECT 115.312 100.386 115.416 104.76 ; 
      RECT 114.88 100.386 114.984 104.76 ; 
      RECT 114.448 100.386 114.552 104.76 ; 
      RECT 114.016 100.386 114.12 104.76 ; 
      RECT 113.584 100.386 113.688 104.76 ; 
      RECT 113.152 100.386 113.256 104.76 ; 
      RECT 112.72 100.386 112.824 104.76 ; 
      RECT 112.288 100.386 112.392 104.76 ; 
      RECT 111.856 100.386 111.96 104.76 ; 
      RECT 111.424 100.386 111.528 104.76 ; 
      RECT 110.992 100.386 111.096 104.76 ; 
      RECT 110.56 100.386 110.664 104.76 ; 
      RECT 110.128 100.386 110.232 104.76 ; 
      RECT 109.696 100.386 109.8 104.76 ; 
      RECT 109.264 100.386 109.368 104.76 ; 
      RECT 108.832 100.386 108.936 104.76 ; 
      RECT 108.4 100.386 108.504 104.76 ; 
      RECT 107.968 100.386 108.072 104.76 ; 
      RECT 107.536 100.386 107.64 104.76 ; 
      RECT 107.104 100.386 107.208 104.76 ; 
      RECT 106.672 100.386 106.776 104.76 ; 
      RECT 106.24 100.386 106.344 104.76 ; 
      RECT 105.808 100.386 105.912 104.76 ; 
      RECT 105.376 100.386 105.48 104.76 ; 
      RECT 104.944 100.386 105.048 104.76 ; 
      RECT 104.512 100.386 104.616 104.76 ; 
      RECT 104.08 100.386 104.184 104.76 ; 
      RECT 103.648 100.386 103.752 104.76 ; 
      RECT 103.216 100.386 103.32 104.76 ; 
      RECT 102.784 100.386 102.888 104.76 ; 
      RECT 102.352 100.386 102.456 104.76 ; 
      RECT 101.92 100.386 102.024 104.76 ; 
      RECT 101.488 100.386 101.592 104.76 ; 
      RECT 101.056 100.386 101.16 104.76 ; 
      RECT 100.624 100.386 100.728 104.76 ; 
      RECT 100.192 100.386 100.296 104.76 ; 
      RECT 99.76 100.386 99.864 104.76 ; 
      RECT 99.328 100.386 99.432 104.76 ; 
      RECT 98.896 100.386 99 104.76 ; 
      RECT 98.464 100.386 98.568 104.76 ; 
      RECT 98.032 100.386 98.136 104.76 ; 
      RECT 97.6 100.386 97.704 104.76 ; 
      RECT 97.168 100.386 97.272 104.76 ; 
      RECT 96.736 100.386 96.84 104.76 ; 
      RECT 96.304 100.386 96.408 104.76 ; 
      RECT 95.872 100.386 95.976 104.76 ; 
      RECT 95.44 100.386 95.544 104.76 ; 
      RECT 95.008 100.386 95.112 104.76 ; 
      RECT 94.576 100.386 94.68 104.76 ; 
      RECT 94.144 100.386 94.248 104.76 ; 
      RECT 93.712 100.386 93.816 104.76 ; 
      RECT 93.28 100.386 93.384 104.76 ; 
      RECT 92.848 100.386 92.952 104.76 ; 
      RECT 92.416 100.386 92.52 104.76 ; 
      RECT 91.984 100.386 92.088 104.76 ; 
      RECT 91.552 100.386 91.656 104.76 ; 
      RECT 91.12 100.386 91.224 104.76 ; 
      RECT 90.688 100.386 90.792 104.76 ; 
      RECT 90.256 100.386 90.36 104.76 ; 
      RECT 89.824 100.386 89.928 104.76 ; 
      RECT 89.392 100.386 89.496 104.76 ; 
      RECT 88.96 100.386 89.064 104.76 ; 
      RECT 88.528 100.386 88.632 104.76 ; 
      RECT 88.096 100.386 88.2 104.76 ; 
      RECT 87.664 100.386 87.768 104.76 ; 
      RECT 87.232 100.386 87.336 104.76 ; 
      RECT 86.8 100.386 86.904 104.76 ; 
      RECT 86.368 100.386 86.472 104.76 ; 
      RECT 85.936 100.386 86.04 104.76 ; 
      RECT 85.504 100.386 85.608 104.76 ; 
      RECT 85.072 100.386 85.176 104.76 ; 
      RECT 84.64 100.386 84.744 104.76 ; 
      RECT 84.208 100.386 84.312 104.76 ; 
      RECT 83.776 100.386 83.88 104.76 ; 
      RECT 83.344 100.386 83.448 104.76 ; 
      RECT 82.912 100.386 83.016 104.76 ; 
      RECT 82.48 100.386 82.584 104.76 ; 
      RECT 82.048 100.386 82.152 104.76 ; 
      RECT 81.616 100.386 81.72 104.76 ; 
      RECT 81.184 100.386 81.288 104.76 ; 
      RECT 80.752 100.386 80.856 104.76 ; 
      RECT 80.32 100.386 80.424 104.76 ; 
      RECT 79.888 100.386 79.992 104.76 ; 
      RECT 79.456 100.386 79.56 104.76 ; 
      RECT 79.024 100.386 79.128 104.76 ; 
      RECT 78.592 100.386 78.696 104.76 ; 
      RECT 78.16 100.386 78.264 104.76 ; 
      RECT 77.728 100.386 77.832 104.76 ; 
      RECT 77.296 100.386 77.4 104.76 ; 
      RECT 76.864 100.386 76.968 104.76 ; 
      RECT 76.432 100.386 76.536 104.76 ; 
      RECT 76 100.386 76.104 104.76 ; 
      RECT 75.568 100.386 75.672 104.76 ; 
      RECT 75.136 100.386 75.24 104.76 ; 
      RECT 74.704 100.386 74.808 104.76 ; 
      RECT 74.272 100.386 74.376 104.76 ; 
      RECT 73.84 100.386 73.944 104.76 ; 
      RECT 73.408 100.386 73.512 104.76 ; 
      RECT 72.976 100.386 73.08 104.76 ; 
      RECT 72.544 100.386 72.648 104.76 ; 
      RECT 72.112 100.386 72.216 104.76 ; 
      RECT 71.68 100.386 71.784 104.76 ; 
      RECT 71.248 100.386 71.352 104.76 ; 
      RECT 70.816 100.386 70.92 104.76 ; 
      RECT 70.384 100.386 70.488 104.76 ; 
      RECT 69.952 100.386 70.056 104.76 ; 
      RECT 69.52 100.386 69.624 104.76 ; 
      RECT 69.088 100.386 69.192 104.76 ; 
      RECT 68.656 100.386 68.76 104.76 ; 
      RECT 68.224 100.386 68.328 104.76 ; 
      RECT 67.792 100.386 67.896 104.76 ; 
      RECT 67.36 100.386 67.464 104.76 ; 
      RECT 66.928 100.386 67.032 104.76 ; 
      RECT 66.496 100.386 66.6 104.76 ; 
      RECT 66.064 100.386 66.168 104.76 ; 
      RECT 65.632 100.386 65.736 104.76 ; 
      RECT 65.2 100.386 65.304 104.76 ; 
      RECT 64.348 100.386 64.656 104.76 ; 
      RECT 56.776 100.386 57.084 104.76 ; 
      RECT 56.128 100.386 56.232 104.76 ; 
      RECT 55.696 100.386 55.8 104.76 ; 
      RECT 55.264 100.386 55.368 104.76 ; 
      RECT 54.832 100.386 54.936 104.76 ; 
      RECT 54.4 100.386 54.504 104.76 ; 
      RECT 53.968 100.386 54.072 104.76 ; 
      RECT 53.536 100.386 53.64 104.76 ; 
      RECT 53.104 100.386 53.208 104.76 ; 
      RECT 52.672 100.386 52.776 104.76 ; 
      RECT 52.24 100.386 52.344 104.76 ; 
      RECT 51.808 100.386 51.912 104.76 ; 
      RECT 51.376 100.386 51.48 104.76 ; 
      RECT 50.944 100.386 51.048 104.76 ; 
      RECT 50.512 100.386 50.616 104.76 ; 
      RECT 50.08 100.386 50.184 104.76 ; 
      RECT 49.648 100.386 49.752 104.76 ; 
      RECT 49.216 100.386 49.32 104.76 ; 
      RECT 48.784 100.386 48.888 104.76 ; 
      RECT 48.352 100.386 48.456 104.76 ; 
      RECT 47.92 100.386 48.024 104.76 ; 
      RECT 47.488 100.386 47.592 104.76 ; 
      RECT 47.056 100.386 47.16 104.76 ; 
      RECT 46.624 100.386 46.728 104.76 ; 
      RECT 46.192 100.386 46.296 104.76 ; 
      RECT 45.76 100.386 45.864 104.76 ; 
      RECT 45.328 100.386 45.432 104.76 ; 
      RECT 44.896 100.386 45 104.76 ; 
      RECT 44.464 100.386 44.568 104.76 ; 
      RECT 44.032 100.386 44.136 104.76 ; 
      RECT 43.6 100.386 43.704 104.76 ; 
      RECT 43.168 100.386 43.272 104.76 ; 
      RECT 42.736 100.386 42.84 104.76 ; 
      RECT 42.304 100.386 42.408 104.76 ; 
      RECT 41.872 100.386 41.976 104.76 ; 
      RECT 41.44 100.386 41.544 104.76 ; 
      RECT 41.008 100.386 41.112 104.76 ; 
      RECT 40.576 100.386 40.68 104.76 ; 
      RECT 40.144 100.386 40.248 104.76 ; 
      RECT 39.712 100.386 39.816 104.76 ; 
      RECT 39.28 100.386 39.384 104.76 ; 
      RECT 38.848 100.386 38.952 104.76 ; 
      RECT 38.416 100.386 38.52 104.76 ; 
      RECT 37.984 100.386 38.088 104.76 ; 
      RECT 37.552 100.386 37.656 104.76 ; 
      RECT 37.12 100.386 37.224 104.76 ; 
      RECT 36.688 100.386 36.792 104.76 ; 
      RECT 36.256 100.386 36.36 104.76 ; 
      RECT 35.824 100.386 35.928 104.76 ; 
      RECT 35.392 100.386 35.496 104.76 ; 
      RECT 34.96 100.386 35.064 104.76 ; 
      RECT 34.528 100.386 34.632 104.76 ; 
      RECT 34.096 100.386 34.2 104.76 ; 
      RECT 33.664 100.386 33.768 104.76 ; 
      RECT 33.232 100.386 33.336 104.76 ; 
      RECT 32.8 100.386 32.904 104.76 ; 
      RECT 32.368 100.386 32.472 104.76 ; 
      RECT 31.936 100.386 32.04 104.76 ; 
      RECT 31.504 100.386 31.608 104.76 ; 
      RECT 31.072 100.386 31.176 104.76 ; 
      RECT 30.64 100.386 30.744 104.76 ; 
      RECT 30.208 100.386 30.312 104.76 ; 
      RECT 29.776 100.386 29.88 104.76 ; 
      RECT 29.344 100.386 29.448 104.76 ; 
      RECT 28.912 100.386 29.016 104.76 ; 
      RECT 28.48 100.386 28.584 104.76 ; 
      RECT 28.048 100.386 28.152 104.76 ; 
      RECT 27.616 100.386 27.72 104.76 ; 
      RECT 27.184 100.386 27.288 104.76 ; 
      RECT 26.752 100.386 26.856 104.76 ; 
      RECT 26.32 100.386 26.424 104.76 ; 
      RECT 25.888 100.386 25.992 104.76 ; 
      RECT 25.456 100.386 25.56 104.76 ; 
      RECT 25.024 100.386 25.128 104.76 ; 
      RECT 24.592 100.386 24.696 104.76 ; 
      RECT 24.16 100.386 24.264 104.76 ; 
      RECT 23.728 100.386 23.832 104.76 ; 
      RECT 23.296 100.386 23.4 104.76 ; 
      RECT 22.864 100.386 22.968 104.76 ; 
      RECT 22.432 100.386 22.536 104.76 ; 
      RECT 22 100.386 22.104 104.76 ; 
      RECT 21.568 100.386 21.672 104.76 ; 
      RECT 21.136 100.386 21.24 104.76 ; 
      RECT 20.704 100.386 20.808 104.76 ; 
      RECT 20.272 100.386 20.376 104.76 ; 
      RECT 19.84 100.386 19.944 104.76 ; 
      RECT 19.408 100.386 19.512 104.76 ; 
      RECT 18.976 100.386 19.08 104.76 ; 
      RECT 18.544 100.386 18.648 104.76 ; 
      RECT 18.112 100.386 18.216 104.76 ; 
      RECT 17.68 100.386 17.784 104.76 ; 
      RECT 17.248 100.386 17.352 104.76 ; 
      RECT 16.816 100.386 16.92 104.76 ; 
      RECT 16.384 100.386 16.488 104.76 ; 
      RECT 15.952 100.386 16.056 104.76 ; 
      RECT 15.52 100.386 15.624 104.76 ; 
      RECT 15.088 100.386 15.192 104.76 ; 
      RECT 14.656 100.386 14.76 104.76 ; 
      RECT 14.224 100.386 14.328 104.76 ; 
      RECT 13.792 100.386 13.896 104.76 ; 
      RECT 13.36 100.386 13.464 104.76 ; 
      RECT 12.928 100.386 13.032 104.76 ; 
      RECT 12.496 100.386 12.6 104.76 ; 
      RECT 12.064 100.386 12.168 104.76 ; 
      RECT 11.632 100.386 11.736 104.76 ; 
      RECT 11.2 100.386 11.304 104.76 ; 
      RECT 10.768 100.386 10.872 104.76 ; 
      RECT 10.336 100.386 10.44 104.76 ; 
      RECT 9.904 100.386 10.008 104.76 ; 
      RECT 9.472 100.386 9.576 104.76 ; 
      RECT 9.04 100.386 9.144 104.76 ; 
      RECT 8.608 100.386 8.712 104.76 ; 
      RECT 8.176 100.386 8.28 104.76 ; 
      RECT 7.744 100.386 7.848 104.76 ; 
      RECT 7.312 100.386 7.416 104.76 ; 
      RECT 6.88 100.386 6.984 104.76 ; 
      RECT 6.448 100.386 6.552 104.76 ; 
      RECT 6.016 100.386 6.12 104.76 ; 
      RECT 5.584 100.386 5.688 104.76 ; 
      RECT 5.152 100.386 5.256 104.76 ; 
      RECT 4.72 100.386 4.824 104.76 ; 
      RECT 4.288 100.386 4.392 104.76 ; 
      RECT 3.856 100.386 3.96 104.76 ; 
      RECT 3.424 100.386 3.528 104.76 ; 
      RECT 2.992 100.386 3.096 104.76 ; 
      RECT 2.56 100.386 2.664 104.76 ; 
      RECT 2.128 100.386 2.232 104.76 ; 
      RECT 1.696 100.386 1.8 104.76 ; 
      RECT 1.264 100.386 1.368 104.76 ; 
      RECT 0.832 100.386 0.936 104.76 ; 
      RECT 0.02 100.386 0.36 104.76 ; 
      RECT 56.54 137.704 121.392 139.468 ; 
      RECT 71.012 104.854 121.392 139.468 ; 
      RECT 65.18 110.87 121.392 139.468 ; 
      RECT 70.148 110.09 121.392 139.468 ; 
      RECT 56.54 136.502 64.852 139.468 ; 
      RECT 62.228 110.474 64.852 139.468 ; 
      RECT 56.54 111.302 61.036 139.468 ; 
      RECT 60.788 104.854 61.036 139.468 ; 
      RECT 62.172 131.438 64.852 135.87 ; 
      RECT 65.124 120.026 121.392 134.398 ; 
      RECT 56.54 132.374 61.092 133.422 ; 
      RECT 62.172 121.286 64.852 130.614 ; 
      RECT 56.54 122.798 61.092 128.022 ; 
      RECT 56.54 112.142 61.092 122.622 ; 
      RECT 62.172 109.982 64.636 117.126 ; 
      RECT 56.756 111.062 61.092 111.822 ; 
      RECT 56.756 107.918 61.036 139.468 ; 
      RECT 57.62 107.594 61.036 139.468 ; 
      RECT 56.756 109.982 61.092 110.886 ; 
      RECT 65.828 110.102 121.392 139.468 ; 
      RECT 65.18 104.854 65.5 139.468 ; 
      RECT 56.54 107.594 57.292 110.85 ; 
      RECT 65.18 104.854 66.364 110.466 ; 
      RECT 65.18 109.322 69.82 110.466 ; 
      RECT 70.148 104.854 70.684 139.468 ; 
      RECT 62.228 109.322 64.636 139.468 ; 
      RECT 63.524 104.854 64.852 109.854 ; 
      RECT 65.18 109.322 70.684 109.698 ; 
      RECT 69.284 104.854 121.392 109.686 ; 
      RECT 56.54 109.406 61.092 109.662 ; 
      RECT 68.42 107.786 121.392 109.686 ; 
      RECT 65.18 107.918 68.092 110.466 ; 
      RECT 62.228 107.918 63.196 139.468 ; 
      RECT 57.62 107.822 61.092 108.87 ; 
      RECT 62.372 104.854 64.852 108.486 ; 
      RECT 67.556 104.854 68.956 108.342 ; 
      RECT 65.18 107.594 67.228 110.466 ; 
      RECT 66.692 104.854 67.228 139.468 ; 
      RECT 57.62 104.854 60.46 139.468 ; 
      RECT 56.9 104.854 57.292 139.468 ; 
      RECT 66.692 104.854 68.956 107.394 ; 
      RECT 62.228 104.854 64.852 107.394 ; 
      RECT 56.9 104.854 60.46 107.394 ; 
      RECT 66.692 104.854 121.392 107.382 ; 
      RECT 62.172 106.742 64.852 107.358 ; 
      RECT 65.18 104.854 121.392 106.326 ; 
      RECT 56.54 104.854 61.036 106.326 ; 
      RECT 56.54 104.854 64.852 105.514 ; 
      RECT 71.028 104.094 71.1 139.468 ; 
      RECT 70.596 104.094 70.668 139.468 ; 
      RECT 70.164 104.094 70.236 139.468 ; 
      RECT 69.732 104.094 69.804 139.468 ; 
      RECT 69.3 104.094 69.372 139.468 ; 
      RECT 68.868 104.094 68.94 139.468 ; 
      RECT 68.436 104.094 68.508 139.468 ; 
      RECT 68.004 104.094 68.076 139.468 ; 
      RECT 67.572 104.094 67.644 139.468 ; 
      RECT 67.14 104.094 67.212 139.468 ; 
      RECT 66.708 104.094 66.78 139.468 ; 
      RECT 66.276 104.094 66.348 139.468 ; 
      RECT 65.844 104.094 65.916 139.468 ; 
      RECT 65.412 104.094 65.484 139.468 ; 
      RECT 0 110.09 56.068 139.468 ; 
      RECT 0 121.246 56.124 121.578 ; 
      RECT 55.028 104.854 56.212 119.892 ; 
      RECT 51.572 108.566 54.7 139.468 ; 
      RECT 0 104.854 51.244 139.468 ; 
      RECT 54.164 104.854 56.212 109.686 ; 
      RECT 0 107.786 53.836 109.686 ; 
      RECT 53.3 104.854 53.836 139.468 ; 
      RECT 52.436 107.594 53.836 139.468 ; 
      RECT 0 104.854 52.108 109.686 ; 
      RECT 52.436 104.854 52.972 139.468 ; 
      RECT 53.3 104.854 56.212 107.394 ; 
      RECT 0 104.854 52.972 107.382 ; 
      RECT 0 104.854 56.212 106.326 ; 
      RECT 53.316 104.748 53.388 139.468 ; 
      RECT 52.884 104.748 52.956 139.468 ; 
        RECT 62.212 137.214 62.724 141.588 ; 
        RECT 62.156 139.876 62.724 141.166 ; 
        RECT 61.276 138.784 61.812 141.588 ; 
        RECT 61.184 140.124 61.812 141.156 ; 
        RECT 61.276 137.214 61.668 141.588 ; 
        RECT 61.276 137.698 61.724 138.656 ; 
        RECT 61.276 137.214 61.812 137.57 ; 
        RECT 60.376 139.016 60.912 141.588 ; 
        RECT 60.376 137.214 60.768 141.588 ; 
        RECT 58.708 137.214 59.04 141.588 ; 
        RECT 58.708 137.568 59.096 141.31 ; 
        RECT 121.072 137.214 121.412 141.588 ; 
        RECT 120.496 137.214 120.6 141.588 ; 
        RECT 120.064 137.214 120.168 141.588 ; 
        RECT 119.632 137.214 119.736 141.588 ; 
        RECT 119.2 137.214 119.304 141.588 ; 
        RECT 118.768 137.214 118.872 141.588 ; 
        RECT 118.336 137.214 118.44 141.588 ; 
        RECT 117.904 137.214 118.008 141.588 ; 
        RECT 117.472 137.214 117.576 141.588 ; 
        RECT 117.04 137.214 117.144 141.588 ; 
        RECT 116.608 137.214 116.712 141.588 ; 
        RECT 116.176 137.214 116.28 141.588 ; 
        RECT 115.744 137.214 115.848 141.588 ; 
        RECT 115.312 137.214 115.416 141.588 ; 
        RECT 114.88 137.214 114.984 141.588 ; 
        RECT 114.448 137.214 114.552 141.588 ; 
        RECT 114.016 137.214 114.12 141.588 ; 
        RECT 113.584 137.214 113.688 141.588 ; 
        RECT 113.152 137.214 113.256 141.588 ; 
        RECT 112.72 137.214 112.824 141.588 ; 
        RECT 112.288 137.214 112.392 141.588 ; 
        RECT 111.856 137.214 111.96 141.588 ; 
        RECT 111.424 137.214 111.528 141.588 ; 
        RECT 110.992 137.214 111.096 141.588 ; 
        RECT 110.56 137.214 110.664 141.588 ; 
        RECT 110.128 137.214 110.232 141.588 ; 
        RECT 109.696 137.214 109.8 141.588 ; 
        RECT 109.264 137.214 109.368 141.588 ; 
        RECT 108.832 137.214 108.936 141.588 ; 
        RECT 108.4 137.214 108.504 141.588 ; 
        RECT 107.968 137.214 108.072 141.588 ; 
        RECT 107.536 137.214 107.64 141.588 ; 
        RECT 107.104 137.214 107.208 141.588 ; 
        RECT 106.672 137.214 106.776 141.588 ; 
        RECT 106.24 137.214 106.344 141.588 ; 
        RECT 105.808 137.214 105.912 141.588 ; 
        RECT 105.376 137.214 105.48 141.588 ; 
        RECT 104.944 137.214 105.048 141.588 ; 
        RECT 104.512 137.214 104.616 141.588 ; 
        RECT 104.08 137.214 104.184 141.588 ; 
        RECT 103.648 137.214 103.752 141.588 ; 
        RECT 103.216 137.214 103.32 141.588 ; 
        RECT 102.784 137.214 102.888 141.588 ; 
        RECT 102.352 137.214 102.456 141.588 ; 
        RECT 101.92 137.214 102.024 141.588 ; 
        RECT 101.488 137.214 101.592 141.588 ; 
        RECT 101.056 137.214 101.16 141.588 ; 
        RECT 100.624 137.214 100.728 141.588 ; 
        RECT 100.192 137.214 100.296 141.588 ; 
        RECT 99.76 137.214 99.864 141.588 ; 
        RECT 99.328 137.214 99.432 141.588 ; 
        RECT 98.896 137.214 99 141.588 ; 
        RECT 98.464 137.214 98.568 141.588 ; 
        RECT 98.032 137.214 98.136 141.588 ; 
        RECT 97.6 137.214 97.704 141.588 ; 
        RECT 97.168 137.214 97.272 141.588 ; 
        RECT 96.736 137.214 96.84 141.588 ; 
        RECT 96.304 137.214 96.408 141.588 ; 
        RECT 95.872 137.214 95.976 141.588 ; 
        RECT 95.44 137.214 95.544 141.588 ; 
        RECT 95.008 137.214 95.112 141.588 ; 
        RECT 94.576 137.214 94.68 141.588 ; 
        RECT 94.144 137.214 94.248 141.588 ; 
        RECT 93.712 137.214 93.816 141.588 ; 
        RECT 93.28 137.214 93.384 141.588 ; 
        RECT 92.848 137.214 92.952 141.588 ; 
        RECT 92.416 137.214 92.52 141.588 ; 
        RECT 91.984 137.214 92.088 141.588 ; 
        RECT 91.552 137.214 91.656 141.588 ; 
        RECT 91.12 137.214 91.224 141.588 ; 
        RECT 90.688 137.214 90.792 141.588 ; 
        RECT 90.256 137.214 90.36 141.588 ; 
        RECT 89.824 137.214 89.928 141.588 ; 
        RECT 89.392 137.214 89.496 141.588 ; 
        RECT 88.96 137.214 89.064 141.588 ; 
        RECT 88.528 137.214 88.632 141.588 ; 
        RECT 88.096 137.214 88.2 141.588 ; 
        RECT 87.664 137.214 87.768 141.588 ; 
        RECT 87.232 137.214 87.336 141.588 ; 
        RECT 86.8 137.214 86.904 141.588 ; 
        RECT 86.368 137.214 86.472 141.588 ; 
        RECT 85.936 137.214 86.04 141.588 ; 
        RECT 85.504 137.214 85.608 141.588 ; 
        RECT 85.072 137.214 85.176 141.588 ; 
        RECT 84.64 137.214 84.744 141.588 ; 
        RECT 84.208 137.214 84.312 141.588 ; 
        RECT 83.776 137.214 83.88 141.588 ; 
        RECT 83.344 137.214 83.448 141.588 ; 
        RECT 82.912 137.214 83.016 141.588 ; 
        RECT 82.48 137.214 82.584 141.588 ; 
        RECT 82.048 137.214 82.152 141.588 ; 
        RECT 81.616 137.214 81.72 141.588 ; 
        RECT 81.184 137.214 81.288 141.588 ; 
        RECT 80.752 137.214 80.856 141.588 ; 
        RECT 80.32 137.214 80.424 141.588 ; 
        RECT 79.888 137.214 79.992 141.588 ; 
        RECT 79.456 137.214 79.56 141.588 ; 
        RECT 79.024 137.214 79.128 141.588 ; 
        RECT 78.592 137.214 78.696 141.588 ; 
        RECT 78.16 137.214 78.264 141.588 ; 
        RECT 77.728 137.214 77.832 141.588 ; 
        RECT 77.296 137.214 77.4 141.588 ; 
        RECT 76.864 137.214 76.968 141.588 ; 
        RECT 76.432 137.214 76.536 141.588 ; 
        RECT 76 137.214 76.104 141.588 ; 
        RECT 75.568 137.214 75.672 141.588 ; 
        RECT 75.136 137.214 75.24 141.588 ; 
        RECT 74.704 137.214 74.808 141.588 ; 
        RECT 74.272 137.214 74.376 141.588 ; 
        RECT 73.84 137.214 73.944 141.588 ; 
        RECT 73.408 137.214 73.512 141.588 ; 
        RECT 72.976 137.214 73.08 141.588 ; 
        RECT 72.544 137.214 72.648 141.588 ; 
        RECT 72.112 137.214 72.216 141.588 ; 
        RECT 71.68 137.214 71.784 141.588 ; 
        RECT 71.248 137.214 71.352 141.588 ; 
        RECT 70.816 137.214 70.92 141.588 ; 
        RECT 70.384 137.214 70.488 141.588 ; 
        RECT 69.952 137.214 70.056 141.588 ; 
        RECT 69.52 137.214 69.624 141.588 ; 
        RECT 69.088 137.214 69.192 141.588 ; 
        RECT 68.656 137.214 68.76 141.588 ; 
        RECT 68.224 137.214 68.328 141.588 ; 
        RECT 67.792 137.214 67.896 141.588 ; 
        RECT 67.36 137.214 67.464 141.588 ; 
        RECT 66.928 137.214 67.032 141.588 ; 
        RECT 66.496 137.214 66.6 141.588 ; 
        RECT 66.064 137.214 66.168 141.588 ; 
        RECT 65.632 137.214 65.736 141.588 ; 
        RECT 65.2 137.214 65.304 141.588 ; 
        RECT 64.348 137.214 64.656 141.588 ; 
        RECT 56.776 137.214 57.084 141.588 ; 
        RECT 56.128 137.214 56.232 141.588 ; 
        RECT 55.696 137.214 55.8 141.588 ; 
        RECT 55.264 137.214 55.368 141.588 ; 
        RECT 54.832 137.214 54.936 141.588 ; 
        RECT 54.4 137.214 54.504 141.588 ; 
        RECT 53.968 137.214 54.072 141.588 ; 
        RECT 53.536 137.214 53.64 141.588 ; 
        RECT 53.104 137.214 53.208 141.588 ; 
        RECT 52.672 137.214 52.776 141.588 ; 
        RECT 52.24 137.214 52.344 141.588 ; 
        RECT 51.808 137.214 51.912 141.588 ; 
        RECT 51.376 137.214 51.48 141.588 ; 
        RECT 50.944 137.214 51.048 141.588 ; 
        RECT 50.512 137.214 50.616 141.588 ; 
        RECT 50.08 137.214 50.184 141.588 ; 
        RECT 49.648 137.214 49.752 141.588 ; 
        RECT 49.216 137.214 49.32 141.588 ; 
        RECT 48.784 137.214 48.888 141.588 ; 
        RECT 48.352 137.214 48.456 141.588 ; 
        RECT 47.92 137.214 48.024 141.588 ; 
        RECT 47.488 137.214 47.592 141.588 ; 
        RECT 47.056 137.214 47.16 141.588 ; 
        RECT 46.624 137.214 46.728 141.588 ; 
        RECT 46.192 137.214 46.296 141.588 ; 
        RECT 45.76 137.214 45.864 141.588 ; 
        RECT 45.328 137.214 45.432 141.588 ; 
        RECT 44.896 137.214 45 141.588 ; 
        RECT 44.464 137.214 44.568 141.588 ; 
        RECT 44.032 137.214 44.136 141.588 ; 
        RECT 43.6 137.214 43.704 141.588 ; 
        RECT 43.168 137.214 43.272 141.588 ; 
        RECT 42.736 137.214 42.84 141.588 ; 
        RECT 42.304 137.214 42.408 141.588 ; 
        RECT 41.872 137.214 41.976 141.588 ; 
        RECT 41.44 137.214 41.544 141.588 ; 
        RECT 41.008 137.214 41.112 141.588 ; 
        RECT 40.576 137.214 40.68 141.588 ; 
        RECT 40.144 137.214 40.248 141.588 ; 
        RECT 39.712 137.214 39.816 141.588 ; 
        RECT 39.28 137.214 39.384 141.588 ; 
        RECT 38.848 137.214 38.952 141.588 ; 
        RECT 38.416 137.214 38.52 141.588 ; 
        RECT 37.984 137.214 38.088 141.588 ; 
        RECT 37.552 137.214 37.656 141.588 ; 
        RECT 37.12 137.214 37.224 141.588 ; 
        RECT 36.688 137.214 36.792 141.588 ; 
        RECT 36.256 137.214 36.36 141.588 ; 
        RECT 35.824 137.214 35.928 141.588 ; 
        RECT 35.392 137.214 35.496 141.588 ; 
        RECT 34.96 137.214 35.064 141.588 ; 
        RECT 34.528 137.214 34.632 141.588 ; 
        RECT 34.096 137.214 34.2 141.588 ; 
        RECT 33.664 137.214 33.768 141.588 ; 
        RECT 33.232 137.214 33.336 141.588 ; 
        RECT 32.8 137.214 32.904 141.588 ; 
        RECT 32.368 137.214 32.472 141.588 ; 
        RECT 31.936 137.214 32.04 141.588 ; 
        RECT 31.504 137.214 31.608 141.588 ; 
        RECT 31.072 137.214 31.176 141.588 ; 
        RECT 30.64 137.214 30.744 141.588 ; 
        RECT 30.208 137.214 30.312 141.588 ; 
        RECT 29.776 137.214 29.88 141.588 ; 
        RECT 29.344 137.214 29.448 141.588 ; 
        RECT 28.912 137.214 29.016 141.588 ; 
        RECT 28.48 137.214 28.584 141.588 ; 
        RECT 28.048 137.214 28.152 141.588 ; 
        RECT 27.616 137.214 27.72 141.588 ; 
        RECT 27.184 137.214 27.288 141.588 ; 
        RECT 26.752 137.214 26.856 141.588 ; 
        RECT 26.32 137.214 26.424 141.588 ; 
        RECT 25.888 137.214 25.992 141.588 ; 
        RECT 25.456 137.214 25.56 141.588 ; 
        RECT 25.024 137.214 25.128 141.588 ; 
        RECT 24.592 137.214 24.696 141.588 ; 
        RECT 24.16 137.214 24.264 141.588 ; 
        RECT 23.728 137.214 23.832 141.588 ; 
        RECT 23.296 137.214 23.4 141.588 ; 
        RECT 22.864 137.214 22.968 141.588 ; 
        RECT 22.432 137.214 22.536 141.588 ; 
        RECT 22 137.214 22.104 141.588 ; 
        RECT 21.568 137.214 21.672 141.588 ; 
        RECT 21.136 137.214 21.24 141.588 ; 
        RECT 20.704 137.214 20.808 141.588 ; 
        RECT 20.272 137.214 20.376 141.588 ; 
        RECT 19.84 137.214 19.944 141.588 ; 
        RECT 19.408 137.214 19.512 141.588 ; 
        RECT 18.976 137.214 19.08 141.588 ; 
        RECT 18.544 137.214 18.648 141.588 ; 
        RECT 18.112 137.214 18.216 141.588 ; 
        RECT 17.68 137.214 17.784 141.588 ; 
        RECT 17.248 137.214 17.352 141.588 ; 
        RECT 16.816 137.214 16.92 141.588 ; 
        RECT 16.384 137.214 16.488 141.588 ; 
        RECT 15.952 137.214 16.056 141.588 ; 
        RECT 15.52 137.214 15.624 141.588 ; 
        RECT 15.088 137.214 15.192 141.588 ; 
        RECT 14.656 137.214 14.76 141.588 ; 
        RECT 14.224 137.214 14.328 141.588 ; 
        RECT 13.792 137.214 13.896 141.588 ; 
        RECT 13.36 137.214 13.464 141.588 ; 
        RECT 12.928 137.214 13.032 141.588 ; 
        RECT 12.496 137.214 12.6 141.588 ; 
        RECT 12.064 137.214 12.168 141.588 ; 
        RECT 11.632 137.214 11.736 141.588 ; 
        RECT 11.2 137.214 11.304 141.588 ; 
        RECT 10.768 137.214 10.872 141.588 ; 
        RECT 10.336 137.214 10.44 141.588 ; 
        RECT 9.904 137.214 10.008 141.588 ; 
        RECT 9.472 137.214 9.576 141.588 ; 
        RECT 9.04 137.214 9.144 141.588 ; 
        RECT 8.608 137.214 8.712 141.588 ; 
        RECT 8.176 137.214 8.28 141.588 ; 
        RECT 7.744 137.214 7.848 141.588 ; 
        RECT 7.312 137.214 7.416 141.588 ; 
        RECT 6.88 137.214 6.984 141.588 ; 
        RECT 6.448 137.214 6.552 141.588 ; 
        RECT 6.016 137.214 6.12 141.588 ; 
        RECT 5.584 137.214 5.688 141.588 ; 
        RECT 5.152 137.214 5.256 141.588 ; 
        RECT 4.72 137.214 4.824 141.588 ; 
        RECT 4.288 137.214 4.392 141.588 ; 
        RECT 3.856 137.214 3.96 141.588 ; 
        RECT 3.424 137.214 3.528 141.588 ; 
        RECT 2.992 137.214 3.096 141.588 ; 
        RECT 2.56 137.214 2.664 141.588 ; 
        RECT 2.128 137.214 2.232 141.588 ; 
        RECT 1.696 137.214 1.8 141.588 ; 
        RECT 1.264 137.214 1.368 141.588 ; 
        RECT 0.832 137.214 0.936 141.588 ; 
        RECT 0.02 137.214 0.36 141.588 ; 
        RECT 62.212 141.534 62.724 145.908 ; 
        RECT 62.156 144.196 62.724 145.486 ; 
        RECT 61.276 143.104 61.812 145.908 ; 
        RECT 61.184 144.444 61.812 145.476 ; 
        RECT 61.276 141.534 61.668 145.908 ; 
        RECT 61.276 142.018 61.724 142.976 ; 
        RECT 61.276 141.534 61.812 141.89 ; 
        RECT 60.376 143.336 60.912 145.908 ; 
        RECT 60.376 141.534 60.768 145.908 ; 
        RECT 58.708 141.534 59.04 145.908 ; 
        RECT 58.708 141.888 59.096 145.63 ; 
        RECT 121.072 141.534 121.412 145.908 ; 
        RECT 120.496 141.534 120.6 145.908 ; 
        RECT 120.064 141.534 120.168 145.908 ; 
        RECT 119.632 141.534 119.736 145.908 ; 
        RECT 119.2 141.534 119.304 145.908 ; 
        RECT 118.768 141.534 118.872 145.908 ; 
        RECT 118.336 141.534 118.44 145.908 ; 
        RECT 117.904 141.534 118.008 145.908 ; 
        RECT 117.472 141.534 117.576 145.908 ; 
        RECT 117.04 141.534 117.144 145.908 ; 
        RECT 116.608 141.534 116.712 145.908 ; 
        RECT 116.176 141.534 116.28 145.908 ; 
        RECT 115.744 141.534 115.848 145.908 ; 
        RECT 115.312 141.534 115.416 145.908 ; 
        RECT 114.88 141.534 114.984 145.908 ; 
        RECT 114.448 141.534 114.552 145.908 ; 
        RECT 114.016 141.534 114.12 145.908 ; 
        RECT 113.584 141.534 113.688 145.908 ; 
        RECT 113.152 141.534 113.256 145.908 ; 
        RECT 112.72 141.534 112.824 145.908 ; 
        RECT 112.288 141.534 112.392 145.908 ; 
        RECT 111.856 141.534 111.96 145.908 ; 
        RECT 111.424 141.534 111.528 145.908 ; 
        RECT 110.992 141.534 111.096 145.908 ; 
        RECT 110.56 141.534 110.664 145.908 ; 
        RECT 110.128 141.534 110.232 145.908 ; 
        RECT 109.696 141.534 109.8 145.908 ; 
        RECT 109.264 141.534 109.368 145.908 ; 
        RECT 108.832 141.534 108.936 145.908 ; 
        RECT 108.4 141.534 108.504 145.908 ; 
        RECT 107.968 141.534 108.072 145.908 ; 
        RECT 107.536 141.534 107.64 145.908 ; 
        RECT 107.104 141.534 107.208 145.908 ; 
        RECT 106.672 141.534 106.776 145.908 ; 
        RECT 106.24 141.534 106.344 145.908 ; 
        RECT 105.808 141.534 105.912 145.908 ; 
        RECT 105.376 141.534 105.48 145.908 ; 
        RECT 104.944 141.534 105.048 145.908 ; 
        RECT 104.512 141.534 104.616 145.908 ; 
        RECT 104.08 141.534 104.184 145.908 ; 
        RECT 103.648 141.534 103.752 145.908 ; 
        RECT 103.216 141.534 103.32 145.908 ; 
        RECT 102.784 141.534 102.888 145.908 ; 
        RECT 102.352 141.534 102.456 145.908 ; 
        RECT 101.92 141.534 102.024 145.908 ; 
        RECT 101.488 141.534 101.592 145.908 ; 
        RECT 101.056 141.534 101.16 145.908 ; 
        RECT 100.624 141.534 100.728 145.908 ; 
        RECT 100.192 141.534 100.296 145.908 ; 
        RECT 99.76 141.534 99.864 145.908 ; 
        RECT 99.328 141.534 99.432 145.908 ; 
        RECT 98.896 141.534 99 145.908 ; 
        RECT 98.464 141.534 98.568 145.908 ; 
        RECT 98.032 141.534 98.136 145.908 ; 
        RECT 97.6 141.534 97.704 145.908 ; 
        RECT 97.168 141.534 97.272 145.908 ; 
        RECT 96.736 141.534 96.84 145.908 ; 
        RECT 96.304 141.534 96.408 145.908 ; 
        RECT 95.872 141.534 95.976 145.908 ; 
        RECT 95.44 141.534 95.544 145.908 ; 
        RECT 95.008 141.534 95.112 145.908 ; 
        RECT 94.576 141.534 94.68 145.908 ; 
        RECT 94.144 141.534 94.248 145.908 ; 
        RECT 93.712 141.534 93.816 145.908 ; 
        RECT 93.28 141.534 93.384 145.908 ; 
        RECT 92.848 141.534 92.952 145.908 ; 
        RECT 92.416 141.534 92.52 145.908 ; 
        RECT 91.984 141.534 92.088 145.908 ; 
        RECT 91.552 141.534 91.656 145.908 ; 
        RECT 91.12 141.534 91.224 145.908 ; 
        RECT 90.688 141.534 90.792 145.908 ; 
        RECT 90.256 141.534 90.36 145.908 ; 
        RECT 89.824 141.534 89.928 145.908 ; 
        RECT 89.392 141.534 89.496 145.908 ; 
        RECT 88.96 141.534 89.064 145.908 ; 
        RECT 88.528 141.534 88.632 145.908 ; 
        RECT 88.096 141.534 88.2 145.908 ; 
        RECT 87.664 141.534 87.768 145.908 ; 
        RECT 87.232 141.534 87.336 145.908 ; 
        RECT 86.8 141.534 86.904 145.908 ; 
        RECT 86.368 141.534 86.472 145.908 ; 
        RECT 85.936 141.534 86.04 145.908 ; 
        RECT 85.504 141.534 85.608 145.908 ; 
        RECT 85.072 141.534 85.176 145.908 ; 
        RECT 84.64 141.534 84.744 145.908 ; 
        RECT 84.208 141.534 84.312 145.908 ; 
        RECT 83.776 141.534 83.88 145.908 ; 
        RECT 83.344 141.534 83.448 145.908 ; 
        RECT 82.912 141.534 83.016 145.908 ; 
        RECT 82.48 141.534 82.584 145.908 ; 
        RECT 82.048 141.534 82.152 145.908 ; 
        RECT 81.616 141.534 81.72 145.908 ; 
        RECT 81.184 141.534 81.288 145.908 ; 
        RECT 80.752 141.534 80.856 145.908 ; 
        RECT 80.32 141.534 80.424 145.908 ; 
        RECT 79.888 141.534 79.992 145.908 ; 
        RECT 79.456 141.534 79.56 145.908 ; 
        RECT 79.024 141.534 79.128 145.908 ; 
        RECT 78.592 141.534 78.696 145.908 ; 
        RECT 78.16 141.534 78.264 145.908 ; 
        RECT 77.728 141.534 77.832 145.908 ; 
        RECT 77.296 141.534 77.4 145.908 ; 
        RECT 76.864 141.534 76.968 145.908 ; 
        RECT 76.432 141.534 76.536 145.908 ; 
        RECT 76 141.534 76.104 145.908 ; 
        RECT 75.568 141.534 75.672 145.908 ; 
        RECT 75.136 141.534 75.24 145.908 ; 
        RECT 74.704 141.534 74.808 145.908 ; 
        RECT 74.272 141.534 74.376 145.908 ; 
        RECT 73.84 141.534 73.944 145.908 ; 
        RECT 73.408 141.534 73.512 145.908 ; 
        RECT 72.976 141.534 73.08 145.908 ; 
        RECT 72.544 141.534 72.648 145.908 ; 
        RECT 72.112 141.534 72.216 145.908 ; 
        RECT 71.68 141.534 71.784 145.908 ; 
        RECT 71.248 141.534 71.352 145.908 ; 
        RECT 70.816 141.534 70.92 145.908 ; 
        RECT 70.384 141.534 70.488 145.908 ; 
        RECT 69.952 141.534 70.056 145.908 ; 
        RECT 69.52 141.534 69.624 145.908 ; 
        RECT 69.088 141.534 69.192 145.908 ; 
        RECT 68.656 141.534 68.76 145.908 ; 
        RECT 68.224 141.534 68.328 145.908 ; 
        RECT 67.792 141.534 67.896 145.908 ; 
        RECT 67.36 141.534 67.464 145.908 ; 
        RECT 66.928 141.534 67.032 145.908 ; 
        RECT 66.496 141.534 66.6 145.908 ; 
        RECT 66.064 141.534 66.168 145.908 ; 
        RECT 65.632 141.534 65.736 145.908 ; 
        RECT 65.2 141.534 65.304 145.908 ; 
        RECT 64.348 141.534 64.656 145.908 ; 
        RECT 56.776 141.534 57.084 145.908 ; 
        RECT 56.128 141.534 56.232 145.908 ; 
        RECT 55.696 141.534 55.8 145.908 ; 
        RECT 55.264 141.534 55.368 145.908 ; 
        RECT 54.832 141.534 54.936 145.908 ; 
        RECT 54.4 141.534 54.504 145.908 ; 
        RECT 53.968 141.534 54.072 145.908 ; 
        RECT 53.536 141.534 53.64 145.908 ; 
        RECT 53.104 141.534 53.208 145.908 ; 
        RECT 52.672 141.534 52.776 145.908 ; 
        RECT 52.24 141.534 52.344 145.908 ; 
        RECT 51.808 141.534 51.912 145.908 ; 
        RECT 51.376 141.534 51.48 145.908 ; 
        RECT 50.944 141.534 51.048 145.908 ; 
        RECT 50.512 141.534 50.616 145.908 ; 
        RECT 50.08 141.534 50.184 145.908 ; 
        RECT 49.648 141.534 49.752 145.908 ; 
        RECT 49.216 141.534 49.32 145.908 ; 
        RECT 48.784 141.534 48.888 145.908 ; 
        RECT 48.352 141.534 48.456 145.908 ; 
        RECT 47.92 141.534 48.024 145.908 ; 
        RECT 47.488 141.534 47.592 145.908 ; 
        RECT 47.056 141.534 47.16 145.908 ; 
        RECT 46.624 141.534 46.728 145.908 ; 
        RECT 46.192 141.534 46.296 145.908 ; 
        RECT 45.76 141.534 45.864 145.908 ; 
        RECT 45.328 141.534 45.432 145.908 ; 
        RECT 44.896 141.534 45 145.908 ; 
        RECT 44.464 141.534 44.568 145.908 ; 
        RECT 44.032 141.534 44.136 145.908 ; 
        RECT 43.6 141.534 43.704 145.908 ; 
        RECT 43.168 141.534 43.272 145.908 ; 
        RECT 42.736 141.534 42.84 145.908 ; 
        RECT 42.304 141.534 42.408 145.908 ; 
        RECT 41.872 141.534 41.976 145.908 ; 
        RECT 41.44 141.534 41.544 145.908 ; 
        RECT 41.008 141.534 41.112 145.908 ; 
        RECT 40.576 141.534 40.68 145.908 ; 
        RECT 40.144 141.534 40.248 145.908 ; 
        RECT 39.712 141.534 39.816 145.908 ; 
        RECT 39.28 141.534 39.384 145.908 ; 
        RECT 38.848 141.534 38.952 145.908 ; 
        RECT 38.416 141.534 38.52 145.908 ; 
        RECT 37.984 141.534 38.088 145.908 ; 
        RECT 37.552 141.534 37.656 145.908 ; 
        RECT 37.12 141.534 37.224 145.908 ; 
        RECT 36.688 141.534 36.792 145.908 ; 
        RECT 36.256 141.534 36.36 145.908 ; 
        RECT 35.824 141.534 35.928 145.908 ; 
        RECT 35.392 141.534 35.496 145.908 ; 
        RECT 34.96 141.534 35.064 145.908 ; 
        RECT 34.528 141.534 34.632 145.908 ; 
        RECT 34.096 141.534 34.2 145.908 ; 
        RECT 33.664 141.534 33.768 145.908 ; 
        RECT 33.232 141.534 33.336 145.908 ; 
        RECT 32.8 141.534 32.904 145.908 ; 
        RECT 32.368 141.534 32.472 145.908 ; 
        RECT 31.936 141.534 32.04 145.908 ; 
        RECT 31.504 141.534 31.608 145.908 ; 
        RECT 31.072 141.534 31.176 145.908 ; 
        RECT 30.64 141.534 30.744 145.908 ; 
        RECT 30.208 141.534 30.312 145.908 ; 
        RECT 29.776 141.534 29.88 145.908 ; 
        RECT 29.344 141.534 29.448 145.908 ; 
        RECT 28.912 141.534 29.016 145.908 ; 
        RECT 28.48 141.534 28.584 145.908 ; 
        RECT 28.048 141.534 28.152 145.908 ; 
        RECT 27.616 141.534 27.72 145.908 ; 
        RECT 27.184 141.534 27.288 145.908 ; 
        RECT 26.752 141.534 26.856 145.908 ; 
        RECT 26.32 141.534 26.424 145.908 ; 
        RECT 25.888 141.534 25.992 145.908 ; 
        RECT 25.456 141.534 25.56 145.908 ; 
        RECT 25.024 141.534 25.128 145.908 ; 
        RECT 24.592 141.534 24.696 145.908 ; 
        RECT 24.16 141.534 24.264 145.908 ; 
        RECT 23.728 141.534 23.832 145.908 ; 
        RECT 23.296 141.534 23.4 145.908 ; 
        RECT 22.864 141.534 22.968 145.908 ; 
        RECT 22.432 141.534 22.536 145.908 ; 
        RECT 22 141.534 22.104 145.908 ; 
        RECT 21.568 141.534 21.672 145.908 ; 
        RECT 21.136 141.534 21.24 145.908 ; 
        RECT 20.704 141.534 20.808 145.908 ; 
        RECT 20.272 141.534 20.376 145.908 ; 
        RECT 19.84 141.534 19.944 145.908 ; 
        RECT 19.408 141.534 19.512 145.908 ; 
        RECT 18.976 141.534 19.08 145.908 ; 
        RECT 18.544 141.534 18.648 145.908 ; 
        RECT 18.112 141.534 18.216 145.908 ; 
        RECT 17.68 141.534 17.784 145.908 ; 
        RECT 17.248 141.534 17.352 145.908 ; 
        RECT 16.816 141.534 16.92 145.908 ; 
        RECT 16.384 141.534 16.488 145.908 ; 
        RECT 15.952 141.534 16.056 145.908 ; 
        RECT 15.52 141.534 15.624 145.908 ; 
        RECT 15.088 141.534 15.192 145.908 ; 
        RECT 14.656 141.534 14.76 145.908 ; 
        RECT 14.224 141.534 14.328 145.908 ; 
        RECT 13.792 141.534 13.896 145.908 ; 
        RECT 13.36 141.534 13.464 145.908 ; 
        RECT 12.928 141.534 13.032 145.908 ; 
        RECT 12.496 141.534 12.6 145.908 ; 
        RECT 12.064 141.534 12.168 145.908 ; 
        RECT 11.632 141.534 11.736 145.908 ; 
        RECT 11.2 141.534 11.304 145.908 ; 
        RECT 10.768 141.534 10.872 145.908 ; 
        RECT 10.336 141.534 10.44 145.908 ; 
        RECT 9.904 141.534 10.008 145.908 ; 
        RECT 9.472 141.534 9.576 145.908 ; 
        RECT 9.04 141.534 9.144 145.908 ; 
        RECT 8.608 141.534 8.712 145.908 ; 
        RECT 8.176 141.534 8.28 145.908 ; 
        RECT 7.744 141.534 7.848 145.908 ; 
        RECT 7.312 141.534 7.416 145.908 ; 
        RECT 6.88 141.534 6.984 145.908 ; 
        RECT 6.448 141.534 6.552 145.908 ; 
        RECT 6.016 141.534 6.12 145.908 ; 
        RECT 5.584 141.534 5.688 145.908 ; 
        RECT 5.152 141.534 5.256 145.908 ; 
        RECT 4.72 141.534 4.824 145.908 ; 
        RECT 4.288 141.534 4.392 145.908 ; 
        RECT 3.856 141.534 3.96 145.908 ; 
        RECT 3.424 141.534 3.528 145.908 ; 
        RECT 2.992 141.534 3.096 145.908 ; 
        RECT 2.56 141.534 2.664 145.908 ; 
        RECT 2.128 141.534 2.232 145.908 ; 
        RECT 1.696 141.534 1.8 145.908 ; 
        RECT 1.264 141.534 1.368 145.908 ; 
        RECT 0.832 141.534 0.936 145.908 ; 
        RECT 0.02 141.534 0.36 145.908 ; 
        RECT 62.212 145.854 62.724 150.228 ; 
        RECT 62.156 148.516 62.724 149.806 ; 
        RECT 61.276 147.424 61.812 150.228 ; 
        RECT 61.184 148.764 61.812 149.796 ; 
        RECT 61.276 145.854 61.668 150.228 ; 
        RECT 61.276 146.338 61.724 147.296 ; 
        RECT 61.276 145.854 61.812 146.21 ; 
        RECT 60.376 147.656 60.912 150.228 ; 
        RECT 60.376 145.854 60.768 150.228 ; 
        RECT 58.708 145.854 59.04 150.228 ; 
        RECT 58.708 146.208 59.096 149.95 ; 
        RECT 121.072 145.854 121.412 150.228 ; 
        RECT 120.496 145.854 120.6 150.228 ; 
        RECT 120.064 145.854 120.168 150.228 ; 
        RECT 119.632 145.854 119.736 150.228 ; 
        RECT 119.2 145.854 119.304 150.228 ; 
        RECT 118.768 145.854 118.872 150.228 ; 
        RECT 118.336 145.854 118.44 150.228 ; 
        RECT 117.904 145.854 118.008 150.228 ; 
        RECT 117.472 145.854 117.576 150.228 ; 
        RECT 117.04 145.854 117.144 150.228 ; 
        RECT 116.608 145.854 116.712 150.228 ; 
        RECT 116.176 145.854 116.28 150.228 ; 
        RECT 115.744 145.854 115.848 150.228 ; 
        RECT 115.312 145.854 115.416 150.228 ; 
        RECT 114.88 145.854 114.984 150.228 ; 
        RECT 114.448 145.854 114.552 150.228 ; 
        RECT 114.016 145.854 114.12 150.228 ; 
        RECT 113.584 145.854 113.688 150.228 ; 
        RECT 113.152 145.854 113.256 150.228 ; 
        RECT 112.72 145.854 112.824 150.228 ; 
        RECT 112.288 145.854 112.392 150.228 ; 
        RECT 111.856 145.854 111.96 150.228 ; 
        RECT 111.424 145.854 111.528 150.228 ; 
        RECT 110.992 145.854 111.096 150.228 ; 
        RECT 110.56 145.854 110.664 150.228 ; 
        RECT 110.128 145.854 110.232 150.228 ; 
        RECT 109.696 145.854 109.8 150.228 ; 
        RECT 109.264 145.854 109.368 150.228 ; 
        RECT 108.832 145.854 108.936 150.228 ; 
        RECT 108.4 145.854 108.504 150.228 ; 
        RECT 107.968 145.854 108.072 150.228 ; 
        RECT 107.536 145.854 107.64 150.228 ; 
        RECT 107.104 145.854 107.208 150.228 ; 
        RECT 106.672 145.854 106.776 150.228 ; 
        RECT 106.24 145.854 106.344 150.228 ; 
        RECT 105.808 145.854 105.912 150.228 ; 
        RECT 105.376 145.854 105.48 150.228 ; 
        RECT 104.944 145.854 105.048 150.228 ; 
        RECT 104.512 145.854 104.616 150.228 ; 
        RECT 104.08 145.854 104.184 150.228 ; 
        RECT 103.648 145.854 103.752 150.228 ; 
        RECT 103.216 145.854 103.32 150.228 ; 
        RECT 102.784 145.854 102.888 150.228 ; 
        RECT 102.352 145.854 102.456 150.228 ; 
        RECT 101.92 145.854 102.024 150.228 ; 
        RECT 101.488 145.854 101.592 150.228 ; 
        RECT 101.056 145.854 101.16 150.228 ; 
        RECT 100.624 145.854 100.728 150.228 ; 
        RECT 100.192 145.854 100.296 150.228 ; 
        RECT 99.76 145.854 99.864 150.228 ; 
        RECT 99.328 145.854 99.432 150.228 ; 
        RECT 98.896 145.854 99 150.228 ; 
        RECT 98.464 145.854 98.568 150.228 ; 
        RECT 98.032 145.854 98.136 150.228 ; 
        RECT 97.6 145.854 97.704 150.228 ; 
        RECT 97.168 145.854 97.272 150.228 ; 
        RECT 96.736 145.854 96.84 150.228 ; 
        RECT 96.304 145.854 96.408 150.228 ; 
        RECT 95.872 145.854 95.976 150.228 ; 
        RECT 95.44 145.854 95.544 150.228 ; 
        RECT 95.008 145.854 95.112 150.228 ; 
        RECT 94.576 145.854 94.68 150.228 ; 
        RECT 94.144 145.854 94.248 150.228 ; 
        RECT 93.712 145.854 93.816 150.228 ; 
        RECT 93.28 145.854 93.384 150.228 ; 
        RECT 92.848 145.854 92.952 150.228 ; 
        RECT 92.416 145.854 92.52 150.228 ; 
        RECT 91.984 145.854 92.088 150.228 ; 
        RECT 91.552 145.854 91.656 150.228 ; 
        RECT 91.12 145.854 91.224 150.228 ; 
        RECT 90.688 145.854 90.792 150.228 ; 
        RECT 90.256 145.854 90.36 150.228 ; 
        RECT 89.824 145.854 89.928 150.228 ; 
        RECT 89.392 145.854 89.496 150.228 ; 
        RECT 88.96 145.854 89.064 150.228 ; 
        RECT 88.528 145.854 88.632 150.228 ; 
        RECT 88.096 145.854 88.2 150.228 ; 
        RECT 87.664 145.854 87.768 150.228 ; 
        RECT 87.232 145.854 87.336 150.228 ; 
        RECT 86.8 145.854 86.904 150.228 ; 
        RECT 86.368 145.854 86.472 150.228 ; 
        RECT 85.936 145.854 86.04 150.228 ; 
        RECT 85.504 145.854 85.608 150.228 ; 
        RECT 85.072 145.854 85.176 150.228 ; 
        RECT 84.64 145.854 84.744 150.228 ; 
        RECT 84.208 145.854 84.312 150.228 ; 
        RECT 83.776 145.854 83.88 150.228 ; 
        RECT 83.344 145.854 83.448 150.228 ; 
        RECT 82.912 145.854 83.016 150.228 ; 
        RECT 82.48 145.854 82.584 150.228 ; 
        RECT 82.048 145.854 82.152 150.228 ; 
        RECT 81.616 145.854 81.72 150.228 ; 
        RECT 81.184 145.854 81.288 150.228 ; 
        RECT 80.752 145.854 80.856 150.228 ; 
        RECT 80.32 145.854 80.424 150.228 ; 
        RECT 79.888 145.854 79.992 150.228 ; 
        RECT 79.456 145.854 79.56 150.228 ; 
        RECT 79.024 145.854 79.128 150.228 ; 
        RECT 78.592 145.854 78.696 150.228 ; 
        RECT 78.16 145.854 78.264 150.228 ; 
        RECT 77.728 145.854 77.832 150.228 ; 
        RECT 77.296 145.854 77.4 150.228 ; 
        RECT 76.864 145.854 76.968 150.228 ; 
        RECT 76.432 145.854 76.536 150.228 ; 
        RECT 76 145.854 76.104 150.228 ; 
        RECT 75.568 145.854 75.672 150.228 ; 
        RECT 75.136 145.854 75.24 150.228 ; 
        RECT 74.704 145.854 74.808 150.228 ; 
        RECT 74.272 145.854 74.376 150.228 ; 
        RECT 73.84 145.854 73.944 150.228 ; 
        RECT 73.408 145.854 73.512 150.228 ; 
        RECT 72.976 145.854 73.08 150.228 ; 
        RECT 72.544 145.854 72.648 150.228 ; 
        RECT 72.112 145.854 72.216 150.228 ; 
        RECT 71.68 145.854 71.784 150.228 ; 
        RECT 71.248 145.854 71.352 150.228 ; 
        RECT 70.816 145.854 70.92 150.228 ; 
        RECT 70.384 145.854 70.488 150.228 ; 
        RECT 69.952 145.854 70.056 150.228 ; 
        RECT 69.52 145.854 69.624 150.228 ; 
        RECT 69.088 145.854 69.192 150.228 ; 
        RECT 68.656 145.854 68.76 150.228 ; 
        RECT 68.224 145.854 68.328 150.228 ; 
        RECT 67.792 145.854 67.896 150.228 ; 
        RECT 67.36 145.854 67.464 150.228 ; 
        RECT 66.928 145.854 67.032 150.228 ; 
        RECT 66.496 145.854 66.6 150.228 ; 
        RECT 66.064 145.854 66.168 150.228 ; 
        RECT 65.632 145.854 65.736 150.228 ; 
        RECT 65.2 145.854 65.304 150.228 ; 
        RECT 64.348 145.854 64.656 150.228 ; 
        RECT 56.776 145.854 57.084 150.228 ; 
        RECT 56.128 145.854 56.232 150.228 ; 
        RECT 55.696 145.854 55.8 150.228 ; 
        RECT 55.264 145.854 55.368 150.228 ; 
        RECT 54.832 145.854 54.936 150.228 ; 
        RECT 54.4 145.854 54.504 150.228 ; 
        RECT 53.968 145.854 54.072 150.228 ; 
        RECT 53.536 145.854 53.64 150.228 ; 
        RECT 53.104 145.854 53.208 150.228 ; 
        RECT 52.672 145.854 52.776 150.228 ; 
        RECT 52.24 145.854 52.344 150.228 ; 
        RECT 51.808 145.854 51.912 150.228 ; 
        RECT 51.376 145.854 51.48 150.228 ; 
        RECT 50.944 145.854 51.048 150.228 ; 
        RECT 50.512 145.854 50.616 150.228 ; 
        RECT 50.08 145.854 50.184 150.228 ; 
        RECT 49.648 145.854 49.752 150.228 ; 
        RECT 49.216 145.854 49.32 150.228 ; 
        RECT 48.784 145.854 48.888 150.228 ; 
        RECT 48.352 145.854 48.456 150.228 ; 
        RECT 47.92 145.854 48.024 150.228 ; 
        RECT 47.488 145.854 47.592 150.228 ; 
        RECT 47.056 145.854 47.16 150.228 ; 
        RECT 46.624 145.854 46.728 150.228 ; 
        RECT 46.192 145.854 46.296 150.228 ; 
        RECT 45.76 145.854 45.864 150.228 ; 
        RECT 45.328 145.854 45.432 150.228 ; 
        RECT 44.896 145.854 45 150.228 ; 
        RECT 44.464 145.854 44.568 150.228 ; 
        RECT 44.032 145.854 44.136 150.228 ; 
        RECT 43.6 145.854 43.704 150.228 ; 
        RECT 43.168 145.854 43.272 150.228 ; 
        RECT 42.736 145.854 42.84 150.228 ; 
        RECT 42.304 145.854 42.408 150.228 ; 
        RECT 41.872 145.854 41.976 150.228 ; 
        RECT 41.44 145.854 41.544 150.228 ; 
        RECT 41.008 145.854 41.112 150.228 ; 
        RECT 40.576 145.854 40.68 150.228 ; 
        RECT 40.144 145.854 40.248 150.228 ; 
        RECT 39.712 145.854 39.816 150.228 ; 
        RECT 39.28 145.854 39.384 150.228 ; 
        RECT 38.848 145.854 38.952 150.228 ; 
        RECT 38.416 145.854 38.52 150.228 ; 
        RECT 37.984 145.854 38.088 150.228 ; 
        RECT 37.552 145.854 37.656 150.228 ; 
        RECT 37.12 145.854 37.224 150.228 ; 
        RECT 36.688 145.854 36.792 150.228 ; 
        RECT 36.256 145.854 36.36 150.228 ; 
        RECT 35.824 145.854 35.928 150.228 ; 
        RECT 35.392 145.854 35.496 150.228 ; 
        RECT 34.96 145.854 35.064 150.228 ; 
        RECT 34.528 145.854 34.632 150.228 ; 
        RECT 34.096 145.854 34.2 150.228 ; 
        RECT 33.664 145.854 33.768 150.228 ; 
        RECT 33.232 145.854 33.336 150.228 ; 
        RECT 32.8 145.854 32.904 150.228 ; 
        RECT 32.368 145.854 32.472 150.228 ; 
        RECT 31.936 145.854 32.04 150.228 ; 
        RECT 31.504 145.854 31.608 150.228 ; 
        RECT 31.072 145.854 31.176 150.228 ; 
        RECT 30.64 145.854 30.744 150.228 ; 
        RECT 30.208 145.854 30.312 150.228 ; 
        RECT 29.776 145.854 29.88 150.228 ; 
        RECT 29.344 145.854 29.448 150.228 ; 
        RECT 28.912 145.854 29.016 150.228 ; 
        RECT 28.48 145.854 28.584 150.228 ; 
        RECT 28.048 145.854 28.152 150.228 ; 
        RECT 27.616 145.854 27.72 150.228 ; 
        RECT 27.184 145.854 27.288 150.228 ; 
        RECT 26.752 145.854 26.856 150.228 ; 
        RECT 26.32 145.854 26.424 150.228 ; 
        RECT 25.888 145.854 25.992 150.228 ; 
        RECT 25.456 145.854 25.56 150.228 ; 
        RECT 25.024 145.854 25.128 150.228 ; 
        RECT 24.592 145.854 24.696 150.228 ; 
        RECT 24.16 145.854 24.264 150.228 ; 
        RECT 23.728 145.854 23.832 150.228 ; 
        RECT 23.296 145.854 23.4 150.228 ; 
        RECT 22.864 145.854 22.968 150.228 ; 
        RECT 22.432 145.854 22.536 150.228 ; 
        RECT 22 145.854 22.104 150.228 ; 
        RECT 21.568 145.854 21.672 150.228 ; 
        RECT 21.136 145.854 21.24 150.228 ; 
        RECT 20.704 145.854 20.808 150.228 ; 
        RECT 20.272 145.854 20.376 150.228 ; 
        RECT 19.84 145.854 19.944 150.228 ; 
        RECT 19.408 145.854 19.512 150.228 ; 
        RECT 18.976 145.854 19.08 150.228 ; 
        RECT 18.544 145.854 18.648 150.228 ; 
        RECT 18.112 145.854 18.216 150.228 ; 
        RECT 17.68 145.854 17.784 150.228 ; 
        RECT 17.248 145.854 17.352 150.228 ; 
        RECT 16.816 145.854 16.92 150.228 ; 
        RECT 16.384 145.854 16.488 150.228 ; 
        RECT 15.952 145.854 16.056 150.228 ; 
        RECT 15.52 145.854 15.624 150.228 ; 
        RECT 15.088 145.854 15.192 150.228 ; 
        RECT 14.656 145.854 14.76 150.228 ; 
        RECT 14.224 145.854 14.328 150.228 ; 
        RECT 13.792 145.854 13.896 150.228 ; 
        RECT 13.36 145.854 13.464 150.228 ; 
        RECT 12.928 145.854 13.032 150.228 ; 
        RECT 12.496 145.854 12.6 150.228 ; 
        RECT 12.064 145.854 12.168 150.228 ; 
        RECT 11.632 145.854 11.736 150.228 ; 
        RECT 11.2 145.854 11.304 150.228 ; 
        RECT 10.768 145.854 10.872 150.228 ; 
        RECT 10.336 145.854 10.44 150.228 ; 
        RECT 9.904 145.854 10.008 150.228 ; 
        RECT 9.472 145.854 9.576 150.228 ; 
        RECT 9.04 145.854 9.144 150.228 ; 
        RECT 8.608 145.854 8.712 150.228 ; 
        RECT 8.176 145.854 8.28 150.228 ; 
        RECT 7.744 145.854 7.848 150.228 ; 
        RECT 7.312 145.854 7.416 150.228 ; 
        RECT 6.88 145.854 6.984 150.228 ; 
        RECT 6.448 145.854 6.552 150.228 ; 
        RECT 6.016 145.854 6.12 150.228 ; 
        RECT 5.584 145.854 5.688 150.228 ; 
        RECT 5.152 145.854 5.256 150.228 ; 
        RECT 4.72 145.854 4.824 150.228 ; 
        RECT 4.288 145.854 4.392 150.228 ; 
        RECT 3.856 145.854 3.96 150.228 ; 
        RECT 3.424 145.854 3.528 150.228 ; 
        RECT 2.992 145.854 3.096 150.228 ; 
        RECT 2.56 145.854 2.664 150.228 ; 
        RECT 2.128 145.854 2.232 150.228 ; 
        RECT 1.696 145.854 1.8 150.228 ; 
        RECT 1.264 145.854 1.368 150.228 ; 
        RECT 0.832 145.854 0.936 150.228 ; 
        RECT 0.02 145.854 0.36 150.228 ; 
        RECT 62.212 150.174 62.724 154.548 ; 
        RECT 62.156 152.836 62.724 154.126 ; 
        RECT 61.276 151.744 61.812 154.548 ; 
        RECT 61.184 153.084 61.812 154.116 ; 
        RECT 61.276 150.174 61.668 154.548 ; 
        RECT 61.276 150.658 61.724 151.616 ; 
        RECT 61.276 150.174 61.812 150.53 ; 
        RECT 60.376 151.976 60.912 154.548 ; 
        RECT 60.376 150.174 60.768 154.548 ; 
        RECT 58.708 150.174 59.04 154.548 ; 
        RECT 58.708 150.528 59.096 154.27 ; 
        RECT 121.072 150.174 121.412 154.548 ; 
        RECT 120.496 150.174 120.6 154.548 ; 
        RECT 120.064 150.174 120.168 154.548 ; 
        RECT 119.632 150.174 119.736 154.548 ; 
        RECT 119.2 150.174 119.304 154.548 ; 
        RECT 118.768 150.174 118.872 154.548 ; 
        RECT 118.336 150.174 118.44 154.548 ; 
        RECT 117.904 150.174 118.008 154.548 ; 
        RECT 117.472 150.174 117.576 154.548 ; 
        RECT 117.04 150.174 117.144 154.548 ; 
        RECT 116.608 150.174 116.712 154.548 ; 
        RECT 116.176 150.174 116.28 154.548 ; 
        RECT 115.744 150.174 115.848 154.548 ; 
        RECT 115.312 150.174 115.416 154.548 ; 
        RECT 114.88 150.174 114.984 154.548 ; 
        RECT 114.448 150.174 114.552 154.548 ; 
        RECT 114.016 150.174 114.12 154.548 ; 
        RECT 113.584 150.174 113.688 154.548 ; 
        RECT 113.152 150.174 113.256 154.548 ; 
        RECT 112.72 150.174 112.824 154.548 ; 
        RECT 112.288 150.174 112.392 154.548 ; 
        RECT 111.856 150.174 111.96 154.548 ; 
        RECT 111.424 150.174 111.528 154.548 ; 
        RECT 110.992 150.174 111.096 154.548 ; 
        RECT 110.56 150.174 110.664 154.548 ; 
        RECT 110.128 150.174 110.232 154.548 ; 
        RECT 109.696 150.174 109.8 154.548 ; 
        RECT 109.264 150.174 109.368 154.548 ; 
        RECT 108.832 150.174 108.936 154.548 ; 
        RECT 108.4 150.174 108.504 154.548 ; 
        RECT 107.968 150.174 108.072 154.548 ; 
        RECT 107.536 150.174 107.64 154.548 ; 
        RECT 107.104 150.174 107.208 154.548 ; 
        RECT 106.672 150.174 106.776 154.548 ; 
        RECT 106.24 150.174 106.344 154.548 ; 
        RECT 105.808 150.174 105.912 154.548 ; 
        RECT 105.376 150.174 105.48 154.548 ; 
        RECT 104.944 150.174 105.048 154.548 ; 
        RECT 104.512 150.174 104.616 154.548 ; 
        RECT 104.08 150.174 104.184 154.548 ; 
        RECT 103.648 150.174 103.752 154.548 ; 
        RECT 103.216 150.174 103.32 154.548 ; 
        RECT 102.784 150.174 102.888 154.548 ; 
        RECT 102.352 150.174 102.456 154.548 ; 
        RECT 101.92 150.174 102.024 154.548 ; 
        RECT 101.488 150.174 101.592 154.548 ; 
        RECT 101.056 150.174 101.16 154.548 ; 
        RECT 100.624 150.174 100.728 154.548 ; 
        RECT 100.192 150.174 100.296 154.548 ; 
        RECT 99.76 150.174 99.864 154.548 ; 
        RECT 99.328 150.174 99.432 154.548 ; 
        RECT 98.896 150.174 99 154.548 ; 
        RECT 98.464 150.174 98.568 154.548 ; 
        RECT 98.032 150.174 98.136 154.548 ; 
        RECT 97.6 150.174 97.704 154.548 ; 
        RECT 97.168 150.174 97.272 154.548 ; 
        RECT 96.736 150.174 96.84 154.548 ; 
        RECT 96.304 150.174 96.408 154.548 ; 
        RECT 95.872 150.174 95.976 154.548 ; 
        RECT 95.44 150.174 95.544 154.548 ; 
        RECT 95.008 150.174 95.112 154.548 ; 
        RECT 94.576 150.174 94.68 154.548 ; 
        RECT 94.144 150.174 94.248 154.548 ; 
        RECT 93.712 150.174 93.816 154.548 ; 
        RECT 93.28 150.174 93.384 154.548 ; 
        RECT 92.848 150.174 92.952 154.548 ; 
        RECT 92.416 150.174 92.52 154.548 ; 
        RECT 91.984 150.174 92.088 154.548 ; 
        RECT 91.552 150.174 91.656 154.548 ; 
        RECT 91.12 150.174 91.224 154.548 ; 
        RECT 90.688 150.174 90.792 154.548 ; 
        RECT 90.256 150.174 90.36 154.548 ; 
        RECT 89.824 150.174 89.928 154.548 ; 
        RECT 89.392 150.174 89.496 154.548 ; 
        RECT 88.96 150.174 89.064 154.548 ; 
        RECT 88.528 150.174 88.632 154.548 ; 
        RECT 88.096 150.174 88.2 154.548 ; 
        RECT 87.664 150.174 87.768 154.548 ; 
        RECT 87.232 150.174 87.336 154.548 ; 
        RECT 86.8 150.174 86.904 154.548 ; 
        RECT 86.368 150.174 86.472 154.548 ; 
        RECT 85.936 150.174 86.04 154.548 ; 
        RECT 85.504 150.174 85.608 154.548 ; 
        RECT 85.072 150.174 85.176 154.548 ; 
        RECT 84.64 150.174 84.744 154.548 ; 
        RECT 84.208 150.174 84.312 154.548 ; 
        RECT 83.776 150.174 83.88 154.548 ; 
        RECT 83.344 150.174 83.448 154.548 ; 
        RECT 82.912 150.174 83.016 154.548 ; 
        RECT 82.48 150.174 82.584 154.548 ; 
        RECT 82.048 150.174 82.152 154.548 ; 
        RECT 81.616 150.174 81.72 154.548 ; 
        RECT 81.184 150.174 81.288 154.548 ; 
        RECT 80.752 150.174 80.856 154.548 ; 
        RECT 80.32 150.174 80.424 154.548 ; 
        RECT 79.888 150.174 79.992 154.548 ; 
        RECT 79.456 150.174 79.56 154.548 ; 
        RECT 79.024 150.174 79.128 154.548 ; 
        RECT 78.592 150.174 78.696 154.548 ; 
        RECT 78.16 150.174 78.264 154.548 ; 
        RECT 77.728 150.174 77.832 154.548 ; 
        RECT 77.296 150.174 77.4 154.548 ; 
        RECT 76.864 150.174 76.968 154.548 ; 
        RECT 76.432 150.174 76.536 154.548 ; 
        RECT 76 150.174 76.104 154.548 ; 
        RECT 75.568 150.174 75.672 154.548 ; 
        RECT 75.136 150.174 75.24 154.548 ; 
        RECT 74.704 150.174 74.808 154.548 ; 
        RECT 74.272 150.174 74.376 154.548 ; 
        RECT 73.84 150.174 73.944 154.548 ; 
        RECT 73.408 150.174 73.512 154.548 ; 
        RECT 72.976 150.174 73.08 154.548 ; 
        RECT 72.544 150.174 72.648 154.548 ; 
        RECT 72.112 150.174 72.216 154.548 ; 
        RECT 71.68 150.174 71.784 154.548 ; 
        RECT 71.248 150.174 71.352 154.548 ; 
        RECT 70.816 150.174 70.92 154.548 ; 
        RECT 70.384 150.174 70.488 154.548 ; 
        RECT 69.952 150.174 70.056 154.548 ; 
        RECT 69.52 150.174 69.624 154.548 ; 
        RECT 69.088 150.174 69.192 154.548 ; 
        RECT 68.656 150.174 68.76 154.548 ; 
        RECT 68.224 150.174 68.328 154.548 ; 
        RECT 67.792 150.174 67.896 154.548 ; 
        RECT 67.36 150.174 67.464 154.548 ; 
        RECT 66.928 150.174 67.032 154.548 ; 
        RECT 66.496 150.174 66.6 154.548 ; 
        RECT 66.064 150.174 66.168 154.548 ; 
        RECT 65.632 150.174 65.736 154.548 ; 
        RECT 65.2 150.174 65.304 154.548 ; 
        RECT 64.348 150.174 64.656 154.548 ; 
        RECT 56.776 150.174 57.084 154.548 ; 
        RECT 56.128 150.174 56.232 154.548 ; 
        RECT 55.696 150.174 55.8 154.548 ; 
        RECT 55.264 150.174 55.368 154.548 ; 
        RECT 54.832 150.174 54.936 154.548 ; 
        RECT 54.4 150.174 54.504 154.548 ; 
        RECT 53.968 150.174 54.072 154.548 ; 
        RECT 53.536 150.174 53.64 154.548 ; 
        RECT 53.104 150.174 53.208 154.548 ; 
        RECT 52.672 150.174 52.776 154.548 ; 
        RECT 52.24 150.174 52.344 154.548 ; 
        RECT 51.808 150.174 51.912 154.548 ; 
        RECT 51.376 150.174 51.48 154.548 ; 
        RECT 50.944 150.174 51.048 154.548 ; 
        RECT 50.512 150.174 50.616 154.548 ; 
        RECT 50.08 150.174 50.184 154.548 ; 
        RECT 49.648 150.174 49.752 154.548 ; 
        RECT 49.216 150.174 49.32 154.548 ; 
        RECT 48.784 150.174 48.888 154.548 ; 
        RECT 48.352 150.174 48.456 154.548 ; 
        RECT 47.92 150.174 48.024 154.548 ; 
        RECT 47.488 150.174 47.592 154.548 ; 
        RECT 47.056 150.174 47.16 154.548 ; 
        RECT 46.624 150.174 46.728 154.548 ; 
        RECT 46.192 150.174 46.296 154.548 ; 
        RECT 45.76 150.174 45.864 154.548 ; 
        RECT 45.328 150.174 45.432 154.548 ; 
        RECT 44.896 150.174 45 154.548 ; 
        RECT 44.464 150.174 44.568 154.548 ; 
        RECT 44.032 150.174 44.136 154.548 ; 
        RECT 43.6 150.174 43.704 154.548 ; 
        RECT 43.168 150.174 43.272 154.548 ; 
        RECT 42.736 150.174 42.84 154.548 ; 
        RECT 42.304 150.174 42.408 154.548 ; 
        RECT 41.872 150.174 41.976 154.548 ; 
        RECT 41.44 150.174 41.544 154.548 ; 
        RECT 41.008 150.174 41.112 154.548 ; 
        RECT 40.576 150.174 40.68 154.548 ; 
        RECT 40.144 150.174 40.248 154.548 ; 
        RECT 39.712 150.174 39.816 154.548 ; 
        RECT 39.28 150.174 39.384 154.548 ; 
        RECT 38.848 150.174 38.952 154.548 ; 
        RECT 38.416 150.174 38.52 154.548 ; 
        RECT 37.984 150.174 38.088 154.548 ; 
        RECT 37.552 150.174 37.656 154.548 ; 
        RECT 37.12 150.174 37.224 154.548 ; 
        RECT 36.688 150.174 36.792 154.548 ; 
        RECT 36.256 150.174 36.36 154.548 ; 
        RECT 35.824 150.174 35.928 154.548 ; 
        RECT 35.392 150.174 35.496 154.548 ; 
        RECT 34.96 150.174 35.064 154.548 ; 
        RECT 34.528 150.174 34.632 154.548 ; 
        RECT 34.096 150.174 34.2 154.548 ; 
        RECT 33.664 150.174 33.768 154.548 ; 
        RECT 33.232 150.174 33.336 154.548 ; 
        RECT 32.8 150.174 32.904 154.548 ; 
        RECT 32.368 150.174 32.472 154.548 ; 
        RECT 31.936 150.174 32.04 154.548 ; 
        RECT 31.504 150.174 31.608 154.548 ; 
        RECT 31.072 150.174 31.176 154.548 ; 
        RECT 30.64 150.174 30.744 154.548 ; 
        RECT 30.208 150.174 30.312 154.548 ; 
        RECT 29.776 150.174 29.88 154.548 ; 
        RECT 29.344 150.174 29.448 154.548 ; 
        RECT 28.912 150.174 29.016 154.548 ; 
        RECT 28.48 150.174 28.584 154.548 ; 
        RECT 28.048 150.174 28.152 154.548 ; 
        RECT 27.616 150.174 27.72 154.548 ; 
        RECT 27.184 150.174 27.288 154.548 ; 
        RECT 26.752 150.174 26.856 154.548 ; 
        RECT 26.32 150.174 26.424 154.548 ; 
        RECT 25.888 150.174 25.992 154.548 ; 
        RECT 25.456 150.174 25.56 154.548 ; 
        RECT 25.024 150.174 25.128 154.548 ; 
        RECT 24.592 150.174 24.696 154.548 ; 
        RECT 24.16 150.174 24.264 154.548 ; 
        RECT 23.728 150.174 23.832 154.548 ; 
        RECT 23.296 150.174 23.4 154.548 ; 
        RECT 22.864 150.174 22.968 154.548 ; 
        RECT 22.432 150.174 22.536 154.548 ; 
        RECT 22 150.174 22.104 154.548 ; 
        RECT 21.568 150.174 21.672 154.548 ; 
        RECT 21.136 150.174 21.24 154.548 ; 
        RECT 20.704 150.174 20.808 154.548 ; 
        RECT 20.272 150.174 20.376 154.548 ; 
        RECT 19.84 150.174 19.944 154.548 ; 
        RECT 19.408 150.174 19.512 154.548 ; 
        RECT 18.976 150.174 19.08 154.548 ; 
        RECT 18.544 150.174 18.648 154.548 ; 
        RECT 18.112 150.174 18.216 154.548 ; 
        RECT 17.68 150.174 17.784 154.548 ; 
        RECT 17.248 150.174 17.352 154.548 ; 
        RECT 16.816 150.174 16.92 154.548 ; 
        RECT 16.384 150.174 16.488 154.548 ; 
        RECT 15.952 150.174 16.056 154.548 ; 
        RECT 15.52 150.174 15.624 154.548 ; 
        RECT 15.088 150.174 15.192 154.548 ; 
        RECT 14.656 150.174 14.76 154.548 ; 
        RECT 14.224 150.174 14.328 154.548 ; 
        RECT 13.792 150.174 13.896 154.548 ; 
        RECT 13.36 150.174 13.464 154.548 ; 
        RECT 12.928 150.174 13.032 154.548 ; 
        RECT 12.496 150.174 12.6 154.548 ; 
        RECT 12.064 150.174 12.168 154.548 ; 
        RECT 11.632 150.174 11.736 154.548 ; 
        RECT 11.2 150.174 11.304 154.548 ; 
        RECT 10.768 150.174 10.872 154.548 ; 
        RECT 10.336 150.174 10.44 154.548 ; 
        RECT 9.904 150.174 10.008 154.548 ; 
        RECT 9.472 150.174 9.576 154.548 ; 
        RECT 9.04 150.174 9.144 154.548 ; 
        RECT 8.608 150.174 8.712 154.548 ; 
        RECT 8.176 150.174 8.28 154.548 ; 
        RECT 7.744 150.174 7.848 154.548 ; 
        RECT 7.312 150.174 7.416 154.548 ; 
        RECT 6.88 150.174 6.984 154.548 ; 
        RECT 6.448 150.174 6.552 154.548 ; 
        RECT 6.016 150.174 6.12 154.548 ; 
        RECT 5.584 150.174 5.688 154.548 ; 
        RECT 5.152 150.174 5.256 154.548 ; 
        RECT 4.72 150.174 4.824 154.548 ; 
        RECT 4.288 150.174 4.392 154.548 ; 
        RECT 3.856 150.174 3.96 154.548 ; 
        RECT 3.424 150.174 3.528 154.548 ; 
        RECT 2.992 150.174 3.096 154.548 ; 
        RECT 2.56 150.174 2.664 154.548 ; 
        RECT 2.128 150.174 2.232 154.548 ; 
        RECT 1.696 150.174 1.8 154.548 ; 
        RECT 1.264 150.174 1.368 154.548 ; 
        RECT 0.832 150.174 0.936 154.548 ; 
        RECT 0.02 150.174 0.36 154.548 ; 
        RECT 62.212 154.494 62.724 158.868 ; 
        RECT 62.156 157.156 62.724 158.446 ; 
        RECT 61.276 156.064 61.812 158.868 ; 
        RECT 61.184 157.404 61.812 158.436 ; 
        RECT 61.276 154.494 61.668 158.868 ; 
        RECT 61.276 154.978 61.724 155.936 ; 
        RECT 61.276 154.494 61.812 154.85 ; 
        RECT 60.376 156.296 60.912 158.868 ; 
        RECT 60.376 154.494 60.768 158.868 ; 
        RECT 58.708 154.494 59.04 158.868 ; 
        RECT 58.708 154.848 59.096 158.59 ; 
        RECT 121.072 154.494 121.412 158.868 ; 
        RECT 120.496 154.494 120.6 158.868 ; 
        RECT 120.064 154.494 120.168 158.868 ; 
        RECT 119.632 154.494 119.736 158.868 ; 
        RECT 119.2 154.494 119.304 158.868 ; 
        RECT 118.768 154.494 118.872 158.868 ; 
        RECT 118.336 154.494 118.44 158.868 ; 
        RECT 117.904 154.494 118.008 158.868 ; 
        RECT 117.472 154.494 117.576 158.868 ; 
        RECT 117.04 154.494 117.144 158.868 ; 
        RECT 116.608 154.494 116.712 158.868 ; 
        RECT 116.176 154.494 116.28 158.868 ; 
        RECT 115.744 154.494 115.848 158.868 ; 
        RECT 115.312 154.494 115.416 158.868 ; 
        RECT 114.88 154.494 114.984 158.868 ; 
        RECT 114.448 154.494 114.552 158.868 ; 
        RECT 114.016 154.494 114.12 158.868 ; 
        RECT 113.584 154.494 113.688 158.868 ; 
        RECT 113.152 154.494 113.256 158.868 ; 
        RECT 112.72 154.494 112.824 158.868 ; 
        RECT 112.288 154.494 112.392 158.868 ; 
        RECT 111.856 154.494 111.96 158.868 ; 
        RECT 111.424 154.494 111.528 158.868 ; 
        RECT 110.992 154.494 111.096 158.868 ; 
        RECT 110.56 154.494 110.664 158.868 ; 
        RECT 110.128 154.494 110.232 158.868 ; 
        RECT 109.696 154.494 109.8 158.868 ; 
        RECT 109.264 154.494 109.368 158.868 ; 
        RECT 108.832 154.494 108.936 158.868 ; 
        RECT 108.4 154.494 108.504 158.868 ; 
        RECT 107.968 154.494 108.072 158.868 ; 
        RECT 107.536 154.494 107.64 158.868 ; 
        RECT 107.104 154.494 107.208 158.868 ; 
        RECT 106.672 154.494 106.776 158.868 ; 
        RECT 106.24 154.494 106.344 158.868 ; 
        RECT 105.808 154.494 105.912 158.868 ; 
        RECT 105.376 154.494 105.48 158.868 ; 
        RECT 104.944 154.494 105.048 158.868 ; 
        RECT 104.512 154.494 104.616 158.868 ; 
        RECT 104.08 154.494 104.184 158.868 ; 
        RECT 103.648 154.494 103.752 158.868 ; 
        RECT 103.216 154.494 103.32 158.868 ; 
        RECT 102.784 154.494 102.888 158.868 ; 
        RECT 102.352 154.494 102.456 158.868 ; 
        RECT 101.92 154.494 102.024 158.868 ; 
        RECT 101.488 154.494 101.592 158.868 ; 
        RECT 101.056 154.494 101.16 158.868 ; 
        RECT 100.624 154.494 100.728 158.868 ; 
        RECT 100.192 154.494 100.296 158.868 ; 
        RECT 99.76 154.494 99.864 158.868 ; 
        RECT 99.328 154.494 99.432 158.868 ; 
        RECT 98.896 154.494 99 158.868 ; 
        RECT 98.464 154.494 98.568 158.868 ; 
        RECT 98.032 154.494 98.136 158.868 ; 
        RECT 97.6 154.494 97.704 158.868 ; 
        RECT 97.168 154.494 97.272 158.868 ; 
        RECT 96.736 154.494 96.84 158.868 ; 
        RECT 96.304 154.494 96.408 158.868 ; 
        RECT 95.872 154.494 95.976 158.868 ; 
        RECT 95.44 154.494 95.544 158.868 ; 
        RECT 95.008 154.494 95.112 158.868 ; 
        RECT 94.576 154.494 94.68 158.868 ; 
        RECT 94.144 154.494 94.248 158.868 ; 
        RECT 93.712 154.494 93.816 158.868 ; 
        RECT 93.28 154.494 93.384 158.868 ; 
        RECT 92.848 154.494 92.952 158.868 ; 
        RECT 92.416 154.494 92.52 158.868 ; 
        RECT 91.984 154.494 92.088 158.868 ; 
        RECT 91.552 154.494 91.656 158.868 ; 
        RECT 91.12 154.494 91.224 158.868 ; 
        RECT 90.688 154.494 90.792 158.868 ; 
        RECT 90.256 154.494 90.36 158.868 ; 
        RECT 89.824 154.494 89.928 158.868 ; 
        RECT 89.392 154.494 89.496 158.868 ; 
        RECT 88.96 154.494 89.064 158.868 ; 
        RECT 88.528 154.494 88.632 158.868 ; 
        RECT 88.096 154.494 88.2 158.868 ; 
        RECT 87.664 154.494 87.768 158.868 ; 
        RECT 87.232 154.494 87.336 158.868 ; 
        RECT 86.8 154.494 86.904 158.868 ; 
        RECT 86.368 154.494 86.472 158.868 ; 
        RECT 85.936 154.494 86.04 158.868 ; 
        RECT 85.504 154.494 85.608 158.868 ; 
        RECT 85.072 154.494 85.176 158.868 ; 
        RECT 84.64 154.494 84.744 158.868 ; 
        RECT 84.208 154.494 84.312 158.868 ; 
        RECT 83.776 154.494 83.88 158.868 ; 
        RECT 83.344 154.494 83.448 158.868 ; 
        RECT 82.912 154.494 83.016 158.868 ; 
        RECT 82.48 154.494 82.584 158.868 ; 
        RECT 82.048 154.494 82.152 158.868 ; 
        RECT 81.616 154.494 81.72 158.868 ; 
        RECT 81.184 154.494 81.288 158.868 ; 
        RECT 80.752 154.494 80.856 158.868 ; 
        RECT 80.32 154.494 80.424 158.868 ; 
        RECT 79.888 154.494 79.992 158.868 ; 
        RECT 79.456 154.494 79.56 158.868 ; 
        RECT 79.024 154.494 79.128 158.868 ; 
        RECT 78.592 154.494 78.696 158.868 ; 
        RECT 78.16 154.494 78.264 158.868 ; 
        RECT 77.728 154.494 77.832 158.868 ; 
        RECT 77.296 154.494 77.4 158.868 ; 
        RECT 76.864 154.494 76.968 158.868 ; 
        RECT 76.432 154.494 76.536 158.868 ; 
        RECT 76 154.494 76.104 158.868 ; 
        RECT 75.568 154.494 75.672 158.868 ; 
        RECT 75.136 154.494 75.24 158.868 ; 
        RECT 74.704 154.494 74.808 158.868 ; 
        RECT 74.272 154.494 74.376 158.868 ; 
        RECT 73.84 154.494 73.944 158.868 ; 
        RECT 73.408 154.494 73.512 158.868 ; 
        RECT 72.976 154.494 73.08 158.868 ; 
        RECT 72.544 154.494 72.648 158.868 ; 
        RECT 72.112 154.494 72.216 158.868 ; 
        RECT 71.68 154.494 71.784 158.868 ; 
        RECT 71.248 154.494 71.352 158.868 ; 
        RECT 70.816 154.494 70.92 158.868 ; 
        RECT 70.384 154.494 70.488 158.868 ; 
        RECT 69.952 154.494 70.056 158.868 ; 
        RECT 69.52 154.494 69.624 158.868 ; 
        RECT 69.088 154.494 69.192 158.868 ; 
        RECT 68.656 154.494 68.76 158.868 ; 
        RECT 68.224 154.494 68.328 158.868 ; 
        RECT 67.792 154.494 67.896 158.868 ; 
        RECT 67.36 154.494 67.464 158.868 ; 
        RECT 66.928 154.494 67.032 158.868 ; 
        RECT 66.496 154.494 66.6 158.868 ; 
        RECT 66.064 154.494 66.168 158.868 ; 
        RECT 65.632 154.494 65.736 158.868 ; 
        RECT 65.2 154.494 65.304 158.868 ; 
        RECT 64.348 154.494 64.656 158.868 ; 
        RECT 56.776 154.494 57.084 158.868 ; 
        RECT 56.128 154.494 56.232 158.868 ; 
        RECT 55.696 154.494 55.8 158.868 ; 
        RECT 55.264 154.494 55.368 158.868 ; 
        RECT 54.832 154.494 54.936 158.868 ; 
        RECT 54.4 154.494 54.504 158.868 ; 
        RECT 53.968 154.494 54.072 158.868 ; 
        RECT 53.536 154.494 53.64 158.868 ; 
        RECT 53.104 154.494 53.208 158.868 ; 
        RECT 52.672 154.494 52.776 158.868 ; 
        RECT 52.24 154.494 52.344 158.868 ; 
        RECT 51.808 154.494 51.912 158.868 ; 
        RECT 51.376 154.494 51.48 158.868 ; 
        RECT 50.944 154.494 51.048 158.868 ; 
        RECT 50.512 154.494 50.616 158.868 ; 
        RECT 50.08 154.494 50.184 158.868 ; 
        RECT 49.648 154.494 49.752 158.868 ; 
        RECT 49.216 154.494 49.32 158.868 ; 
        RECT 48.784 154.494 48.888 158.868 ; 
        RECT 48.352 154.494 48.456 158.868 ; 
        RECT 47.92 154.494 48.024 158.868 ; 
        RECT 47.488 154.494 47.592 158.868 ; 
        RECT 47.056 154.494 47.16 158.868 ; 
        RECT 46.624 154.494 46.728 158.868 ; 
        RECT 46.192 154.494 46.296 158.868 ; 
        RECT 45.76 154.494 45.864 158.868 ; 
        RECT 45.328 154.494 45.432 158.868 ; 
        RECT 44.896 154.494 45 158.868 ; 
        RECT 44.464 154.494 44.568 158.868 ; 
        RECT 44.032 154.494 44.136 158.868 ; 
        RECT 43.6 154.494 43.704 158.868 ; 
        RECT 43.168 154.494 43.272 158.868 ; 
        RECT 42.736 154.494 42.84 158.868 ; 
        RECT 42.304 154.494 42.408 158.868 ; 
        RECT 41.872 154.494 41.976 158.868 ; 
        RECT 41.44 154.494 41.544 158.868 ; 
        RECT 41.008 154.494 41.112 158.868 ; 
        RECT 40.576 154.494 40.68 158.868 ; 
        RECT 40.144 154.494 40.248 158.868 ; 
        RECT 39.712 154.494 39.816 158.868 ; 
        RECT 39.28 154.494 39.384 158.868 ; 
        RECT 38.848 154.494 38.952 158.868 ; 
        RECT 38.416 154.494 38.52 158.868 ; 
        RECT 37.984 154.494 38.088 158.868 ; 
        RECT 37.552 154.494 37.656 158.868 ; 
        RECT 37.12 154.494 37.224 158.868 ; 
        RECT 36.688 154.494 36.792 158.868 ; 
        RECT 36.256 154.494 36.36 158.868 ; 
        RECT 35.824 154.494 35.928 158.868 ; 
        RECT 35.392 154.494 35.496 158.868 ; 
        RECT 34.96 154.494 35.064 158.868 ; 
        RECT 34.528 154.494 34.632 158.868 ; 
        RECT 34.096 154.494 34.2 158.868 ; 
        RECT 33.664 154.494 33.768 158.868 ; 
        RECT 33.232 154.494 33.336 158.868 ; 
        RECT 32.8 154.494 32.904 158.868 ; 
        RECT 32.368 154.494 32.472 158.868 ; 
        RECT 31.936 154.494 32.04 158.868 ; 
        RECT 31.504 154.494 31.608 158.868 ; 
        RECT 31.072 154.494 31.176 158.868 ; 
        RECT 30.64 154.494 30.744 158.868 ; 
        RECT 30.208 154.494 30.312 158.868 ; 
        RECT 29.776 154.494 29.88 158.868 ; 
        RECT 29.344 154.494 29.448 158.868 ; 
        RECT 28.912 154.494 29.016 158.868 ; 
        RECT 28.48 154.494 28.584 158.868 ; 
        RECT 28.048 154.494 28.152 158.868 ; 
        RECT 27.616 154.494 27.72 158.868 ; 
        RECT 27.184 154.494 27.288 158.868 ; 
        RECT 26.752 154.494 26.856 158.868 ; 
        RECT 26.32 154.494 26.424 158.868 ; 
        RECT 25.888 154.494 25.992 158.868 ; 
        RECT 25.456 154.494 25.56 158.868 ; 
        RECT 25.024 154.494 25.128 158.868 ; 
        RECT 24.592 154.494 24.696 158.868 ; 
        RECT 24.16 154.494 24.264 158.868 ; 
        RECT 23.728 154.494 23.832 158.868 ; 
        RECT 23.296 154.494 23.4 158.868 ; 
        RECT 22.864 154.494 22.968 158.868 ; 
        RECT 22.432 154.494 22.536 158.868 ; 
        RECT 22 154.494 22.104 158.868 ; 
        RECT 21.568 154.494 21.672 158.868 ; 
        RECT 21.136 154.494 21.24 158.868 ; 
        RECT 20.704 154.494 20.808 158.868 ; 
        RECT 20.272 154.494 20.376 158.868 ; 
        RECT 19.84 154.494 19.944 158.868 ; 
        RECT 19.408 154.494 19.512 158.868 ; 
        RECT 18.976 154.494 19.08 158.868 ; 
        RECT 18.544 154.494 18.648 158.868 ; 
        RECT 18.112 154.494 18.216 158.868 ; 
        RECT 17.68 154.494 17.784 158.868 ; 
        RECT 17.248 154.494 17.352 158.868 ; 
        RECT 16.816 154.494 16.92 158.868 ; 
        RECT 16.384 154.494 16.488 158.868 ; 
        RECT 15.952 154.494 16.056 158.868 ; 
        RECT 15.52 154.494 15.624 158.868 ; 
        RECT 15.088 154.494 15.192 158.868 ; 
        RECT 14.656 154.494 14.76 158.868 ; 
        RECT 14.224 154.494 14.328 158.868 ; 
        RECT 13.792 154.494 13.896 158.868 ; 
        RECT 13.36 154.494 13.464 158.868 ; 
        RECT 12.928 154.494 13.032 158.868 ; 
        RECT 12.496 154.494 12.6 158.868 ; 
        RECT 12.064 154.494 12.168 158.868 ; 
        RECT 11.632 154.494 11.736 158.868 ; 
        RECT 11.2 154.494 11.304 158.868 ; 
        RECT 10.768 154.494 10.872 158.868 ; 
        RECT 10.336 154.494 10.44 158.868 ; 
        RECT 9.904 154.494 10.008 158.868 ; 
        RECT 9.472 154.494 9.576 158.868 ; 
        RECT 9.04 154.494 9.144 158.868 ; 
        RECT 8.608 154.494 8.712 158.868 ; 
        RECT 8.176 154.494 8.28 158.868 ; 
        RECT 7.744 154.494 7.848 158.868 ; 
        RECT 7.312 154.494 7.416 158.868 ; 
        RECT 6.88 154.494 6.984 158.868 ; 
        RECT 6.448 154.494 6.552 158.868 ; 
        RECT 6.016 154.494 6.12 158.868 ; 
        RECT 5.584 154.494 5.688 158.868 ; 
        RECT 5.152 154.494 5.256 158.868 ; 
        RECT 4.72 154.494 4.824 158.868 ; 
        RECT 4.288 154.494 4.392 158.868 ; 
        RECT 3.856 154.494 3.96 158.868 ; 
        RECT 3.424 154.494 3.528 158.868 ; 
        RECT 2.992 154.494 3.096 158.868 ; 
        RECT 2.56 154.494 2.664 158.868 ; 
        RECT 2.128 154.494 2.232 158.868 ; 
        RECT 1.696 154.494 1.8 158.868 ; 
        RECT 1.264 154.494 1.368 158.868 ; 
        RECT 0.832 154.494 0.936 158.868 ; 
        RECT 0.02 154.494 0.36 158.868 ; 
        RECT 62.212 158.814 62.724 163.188 ; 
        RECT 62.156 161.476 62.724 162.766 ; 
        RECT 61.276 160.384 61.812 163.188 ; 
        RECT 61.184 161.724 61.812 162.756 ; 
        RECT 61.276 158.814 61.668 163.188 ; 
        RECT 61.276 159.298 61.724 160.256 ; 
        RECT 61.276 158.814 61.812 159.17 ; 
        RECT 60.376 160.616 60.912 163.188 ; 
        RECT 60.376 158.814 60.768 163.188 ; 
        RECT 58.708 158.814 59.04 163.188 ; 
        RECT 58.708 159.168 59.096 162.91 ; 
        RECT 121.072 158.814 121.412 163.188 ; 
        RECT 120.496 158.814 120.6 163.188 ; 
        RECT 120.064 158.814 120.168 163.188 ; 
        RECT 119.632 158.814 119.736 163.188 ; 
        RECT 119.2 158.814 119.304 163.188 ; 
        RECT 118.768 158.814 118.872 163.188 ; 
        RECT 118.336 158.814 118.44 163.188 ; 
        RECT 117.904 158.814 118.008 163.188 ; 
        RECT 117.472 158.814 117.576 163.188 ; 
        RECT 117.04 158.814 117.144 163.188 ; 
        RECT 116.608 158.814 116.712 163.188 ; 
        RECT 116.176 158.814 116.28 163.188 ; 
        RECT 115.744 158.814 115.848 163.188 ; 
        RECT 115.312 158.814 115.416 163.188 ; 
        RECT 114.88 158.814 114.984 163.188 ; 
        RECT 114.448 158.814 114.552 163.188 ; 
        RECT 114.016 158.814 114.12 163.188 ; 
        RECT 113.584 158.814 113.688 163.188 ; 
        RECT 113.152 158.814 113.256 163.188 ; 
        RECT 112.72 158.814 112.824 163.188 ; 
        RECT 112.288 158.814 112.392 163.188 ; 
        RECT 111.856 158.814 111.96 163.188 ; 
        RECT 111.424 158.814 111.528 163.188 ; 
        RECT 110.992 158.814 111.096 163.188 ; 
        RECT 110.56 158.814 110.664 163.188 ; 
        RECT 110.128 158.814 110.232 163.188 ; 
        RECT 109.696 158.814 109.8 163.188 ; 
        RECT 109.264 158.814 109.368 163.188 ; 
        RECT 108.832 158.814 108.936 163.188 ; 
        RECT 108.4 158.814 108.504 163.188 ; 
        RECT 107.968 158.814 108.072 163.188 ; 
        RECT 107.536 158.814 107.64 163.188 ; 
        RECT 107.104 158.814 107.208 163.188 ; 
        RECT 106.672 158.814 106.776 163.188 ; 
        RECT 106.24 158.814 106.344 163.188 ; 
        RECT 105.808 158.814 105.912 163.188 ; 
        RECT 105.376 158.814 105.48 163.188 ; 
        RECT 104.944 158.814 105.048 163.188 ; 
        RECT 104.512 158.814 104.616 163.188 ; 
        RECT 104.08 158.814 104.184 163.188 ; 
        RECT 103.648 158.814 103.752 163.188 ; 
        RECT 103.216 158.814 103.32 163.188 ; 
        RECT 102.784 158.814 102.888 163.188 ; 
        RECT 102.352 158.814 102.456 163.188 ; 
        RECT 101.92 158.814 102.024 163.188 ; 
        RECT 101.488 158.814 101.592 163.188 ; 
        RECT 101.056 158.814 101.16 163.188 ; 
        RECT 100.624 158.814 100.728 163.188 ; 
        RECT 100.192 158.814 100.296 163.188 ; 
        RECT 99.76 158.814 99.864 163.188 ; 
        RECT 99.328 158.814 99.432 163.188 ; 
        RECT 98.896 158.814 99 163.188 ; 
        RECT 98.464 158.814 98.568 163.188 ; 
        RECT 98.032 158.814 98.136 163.188 ; 
        RECT 97.6 158.814 97.704 163.188 ; 
        RECT 97.168 158.814 97.272 163.188 ; 
        RECT 96.736 158.814 96.84 163.188 ; 
        RECT 96.304 158.814 96.408 163.188 ; 
        RECT 95.872 158.814 95.976 163.188 ; 
        RECT 95.44 158.814 95.544 163.188 ; 
        RECT 95.008 158.814 95.112 163.188 ; 
        RECT 94.576 158.814 94.68 163.188 ; 
        RECT 94.144 158.814 94.248 163.188 ; 
        RECT 93.712 158.814 93.816 163.188 ; 
        RECT 93.28 158.814 93.384 163.188 ; 
        RECT 92.848 158.814 92.952 163.188 ; 
        RECT 92.416 158.814 92.52 163.188 ; 
        RECT 91.984 158.814 92.088 163.188 ; 
        RECT 91.552 158.814 91.656 163.188 ; 
        RECT 91.12 158.814 91.224 163.188 ; 
        RECT 90.688 158.814 90.792 163.188 ; 
        RECT 90.256 158.814 90.36 163.188 ; 
        RECT 89.824 158.814 89.928 163.188 ; 
        RECT 89.392 158.814 89.496 163.188 ; 
        RECT 88.96 158.814 89.064 163.188 ; 
        RECT 88.528 158.814 88.632 163.188 ; 
        RECT 88.096 158.814 88.2 163.188 ; 
        RECT 87.664 158.814 87.768 163.188 ; 
        RECT 87.232 158.814 87.336 163.188 ; 
        RECT 86.8 158.814 86.904 163.188 ; 
        RECT 86.368 158.814 86.472 163.188 ; 
        RECT 85.936 158.814 86.04 163.188 ; 
        RECT 85.504 158.814 85.608 163.188 ; 
        RECT 85.072 158.814 85.176 163.188 ; 
        RECT 84.64 158.814 84.744 163.188 ; 
        RECT 84.208 158.814 84.312 163.188 ; 
        RECT 83.776 158.814 83.88 163.188 ; 
        RECT 83.344 158.814 83.448 163.188 ; 
        RECT 82.912 158.814 83.016 163.188 ; 
        RECT 82.48 158.814 82.584 163.188 ; 
        RECT 82.048 158.814 82.152 163.188 ; 
        RECT 81.616 158.814 81.72 163.188 ; 
        RECT 81.184 158.814 81.288 163.188 ; 
        RECT 80.752 158.814 80.856 163.188 ; 
        RECT 80.32 158.814 80.424 163.188 ; 
        RECT 79.888 158.814 79.992 163.188 ; 
        RECT 79.456 158.814 79.56 163.188 ; 
        RECT 79.024 158.814 79.128 163.188 ; 
        RECT 78.592 158.814 78.696 163.188 ; 
        RECT 78.16 158.814 78.264 163.188 ; 
        RECT 77.728 158.814 77.832 163.188 ; 
        RECT 77.296 158.814 77.4 163.188 ; 
        RECT 76.864 158.814 76.968 163.188 ; 
        RECT 76.432 158.814 76.536 163.188 ; 
        RECT 76 158.814 76.104 163.188 ; 
        RECT 75.568 158.814 75.672 163.188 ; 
        RECT 75.136 158.814 75.24 163.188 ; 
        RECT 74.704 158.814 74.808 163.188 ; 
        RECT 74.272 158.814 74.376 163.188 ; 
        RECT 73.84 158.814 73.944 163.188 ; 
        RECT 73.408 158.814 73.512 163.188 ; 
        RECT 72.976 158.814 73.08 163.188 ; 
        RECT 72.544 158.814 72.648 163.188 ; 
        RECT 72.112 158.814 72.216 163.188 ; 
        RECT 71.68 158.814 71.784 163.188 ; 
        RECT 71.248 158.814 71.352 163.188 ; 
        RECT 70.816 158.814 70.92 163.188 ; 
        RECT 70.384 158.814 70.488 163.188 ; 
        RECT 69.952 158.814 70.056 163.188 ; 
        RECT 69.52 158.814 69.624 163.188 ; 
        RECT 69.088 158.814 69.192 163.188 ; 
        RECT 68.656 158.814 68.76 163.188 ; 
        RECT 68.224 158.814 68.328 163.188 ; 
        RECT 67.792 158.814 67.896 163.188 ; 
        RECT 67.36 158.814 67.464 163.188 ; 
        RECT 66.928 158.814 67.032 163.188 ; 
        RECT 66.496 158.814 66.6 163.188 ; 
        RECT 66.064 158.814 66.168 163.188 ; 
        RECT 65.632 158.814 65.736 163.188 ; 
        RECT 65.2 158.814 65.304 163.188 ; 
        RECT 64.348 158.814 64.656 163.188 ; 
        RECT 56.776 158.814 57.084 163.188 ; 
        RECT 56.128 158.814 56.232 163.188 ; 
        RECT 55.696 158.814 55.8 163.188 ; 
        RECT 55.264 158.814 55.368 163.188 ; 
        RECT 54.832 158.814 54.936 163.188 ; 
        RECT 54.4 158.814 54.504 163.188 ; 
        RECT 53.968 158.814 54.072 163.188 ; 
        RECT 53.536 158.814 53.64 163.188 ; 
        RECT 53.104 158.814 53.208 163.188 ; 
        RECT 52.672 158.814 52.776 163.188 ; 
        RECT 52.24 158.814 52.344 163.188 ; 
        RECT 51.808 158.814 51.912 163.188 ; 
        RECT 51.376 158.814 51.48 163.188 ; 
        RECT 50.944 158.814 51.048 163.188 ; 
        RECT 50.512 158.814 50.616 163.188 ; 
        RECT 50.08 158.814 50.184 163.188 ; 
        RECT 49.648 158.814 49.752 163.188 ; 
        RECT 49.216 158.814 49.32 163.188 ; 
        RECT 48.784 158.814 48.888 163.188 ; 
        RECT 48.352 158.814 48.456 163.188 ; 
        RECT 47.92 158.814 48.024 163.188 ; 
        RECT 47.488 158.814 47.592 163.188 ; 
        RECT 47.056 158.814 47.16 163.188 ; 
        RECT 46.624 158.814 46.728 163.188 ; 
        RECT 46.192 158.814 46.296 163.188 ; 
        RECT 45.76 158.814 45.864 163.188 ; 
        RECT 45.328 158.814 45.432 163.188 ; 
        RECT 44.896 158.814 45 163.188 ; 
        RECT 44.464 158.814 44.568 163.188 ; 
        RECT 44.032 158.814 44.136 163.188 ; 
        RECT 43.6 158.814 43.704 163.188 ; 
        RECT 43.168 158.814 43.272 163.188 ; 
        RECT 42.736 158.814 42.84 163.188 ; 
        RECT 42.304 158.814 42.408 163.188 ; 
        RECT 41.872 158.814 41.976 163.188 ; 
        RECT 41.44 158.814 41.544 163.188 ; 
        RECT 41.008 158.814 41.112 163.188 ; 
        RECT 40.576 158.814 40.68 163.188 ; 
        RECT 40.144 158.814 40.248 163.188 ; 
        RECT 39.712 158.814 39.816 163.188 ; 
        RECT 39.28 158.814 39.384 163.188 ; 
        RECT 38.848 158.814 38.952 163.188 ; 
        RECT 38.416 158.814 38.52 163.188 ; 
        RECT 37.984 158.814 38.088 163.188 ; 
        RECT 37.552 158.814 37.656 163.188 ; 
        RECT 37.12 158.814 37.224 163.188 ; 
        RECT 36.688 158.814 36.792 163.188 ; 
        RECT 36.256 158.814 36.36 163.188 ; 
        RECT 35.824 158.814 35.928 163.188 ; 
        RECT 35.392 158.814 35.496 163.188 ; 
        RECT 34.96 158.814 35.064 163.188 ; 
        RECT 34.528 158.814 34.632 163.188 ; 
        RECT 34.096 158.814 34.2 163.188 ; 
        RECT 33.664 158.814 33.768 163.188 ; 
        RECT 33.232 158.814 33.336 163.188 ; 
        RECT 32.8 158.814 32.904 163.188 ; 
        RECT 32.368 158.814 32.472 163.188 ; 
        RECT 31.936 158.814 32.04 163.188 ; 
        RECT 31.504 158.814 31.608 163.188 ; 
        RECT 31.072 158.814 31.176 163.188 ; 
        RECT 30.64 158.814 30.744 163.188 ; 
        RECT 30.208 158.814 30.312 163.188 ; 
        RECT 29.776 158.814 29.88 163.188 ; 
        RECT 29.344 158.814 29.448 163.188 ; 
        RECT 28.912 158.814 29.016 163.188 ; 
        RECT 28.48 158.814 28.584 163.188 ; 
        RECT 28.048 158.814 28.152 163.188 ; 
        RECT 27.616 158.814 27.72 163.188 ; 
        RECT 27.184 158.814 27.288 163.188 ; 
        RECT 26.752 158.814 26.856 163.188 ; 
        RECT 26.32 158.814 26.424 163.188 ; 
        RECT 25.888 158.814 25.992 163.188 ; 
        RECT 25.456 158.814 25.56 163.188 ; 
        RECT 25.024 158.814 25.128 163.188 ; 
        RECT 24.592 158.814 24.696 163.188 ; 
        RECT 24.16 158.814 24.264 163.188 ; 
        RECT 23.728 158.814 23.832 163.188 ; 
        RECT 23.296 158.814 23.4 163.188 ; 
        RECT 22.864 158.814 22.968 163.188 ; 
        RECT 22.432 158.814 22.536 163.188 ; 
        RECT 22 158.814 22.104 163.188 ; 
        RECT 21.568 158.814 21.672 163.188 ; 
        RECT 21.136 158.814 21.24 163.188 ; 
        RECT 20.704 158.814 20.808 163.188 ; 
        RECT 20.272 158.814 20.376 163.188 ; 
        RECT 19.84 158.814 19.944 163.188 ; 
        RECT 19.408 158.814 19.512 163.188 ; 
        RECT 18.976 158.814 19.08 163.188 ; 
        RECT 18.544 158.814 18.648 163.188 ; 
        RECT 18.112 158.814 18.216 163.188 ; 
        RECT 17.68 158.814 17.784 163.188 ; 
        RECT 17.248 158.814 17.352 163.188 ; 
        RECT 16.816 158.814 16.92 163.188 ; 
        RECT 16.384 158.814 16.488 163.188 ; 
        RECT 15.952 158.814 16.056 163.188 ; 
        RECT 15.52 158.814 15.624 163.188 ; 
        RECT 15.088 158.814 15.192 163.188 ; 
        RECT 14.656 158.814 14.76 163.188 ; 
        RECT 14.224 158.814 14.328 163.188 ; 
        RECT 13.792 158.814 13.896 163.188 ; 
        RECT 13.36 158.814 13.464 163.188 ; 
        RECT 12.928 158.814 13.032 163.188 ; 
        RECT 12.496 158.814 12.6 163.188 ; 
        RECT 12.064 158.814 12.168 163.188 ; 
        RECT 11.632 158.814 11.736 163.188 ; 
        RECT 11.2 158.814 11.304 163.188 ; 
        RECT 10.768 158.814 10.872 163.188 ; 
        RECT 10.336 158.814 10.44 163.188 ; 
        RECT 9.904 158.814 10.008 163.188 ; 
        RECT 9.472 158.814 9.576 163.188 ; 
        RECT 9.04 158.814 9.144 163.188 ; 
        RECT 8.608 158.814 8.712 163.188 ; 
        RECT 8.176 158.814 8.28 163.188 ; 
        RECT 7.744 158.814 7.848 163.188 ; 
        RECT 7.312 158.814 7.416 163.188 ; 
        RECT 6.88 158.814 6.984 163.188 ; 
        RECT 6.448 158.814 6.552 163.188 ; 
        RECT 6.016 158.814 6.12 163.188 ; 
        RECT 5.584 158.814 5.688 163.188 ; 
        RECT 5.152 158.814 5.256 163.188 ; 
        RECT 4.72 158.814 4.824 163.188 ; 
        RECT 4.288 158.814 4.392 163.188 ; 
        RECT 3.856 158.814 3.96 163.188 ; 
        RECT 3.424 158.814 3.528 163.188 ; 
        RECT 2.992 158.814 3.096 163.188 ; 
        RECT 2.56 158.814 2.664 163.188 ; 
        RECT 2.128 158.814 2.232 163.188 ; 
        RECT 1.696 158.814 1.8 163.188 ; 
        RECT 1.264 158.814 1.368 163.188 ; 
        RECT 0.832 158.814 0.936 163.188 ; 
        RECT 0.02 158.814 0.36 163.188 ; 
        RECT 62.212 163.134 62.724 167.508 ; 
        RECT 62.156 165.796 62.724 167.086 ; 
        RECT 61.276 164.704 61.812 167.508 ; 
        RECT 61.184 166.044 61.812 167.076 ; 
        RECT 61.276 163.134 61.668 167.508 ; 
        RECT 61.276 163.618 61.724 164.576 ; 
        RECT 61.276 163.134 61.812 163.49 ; 
        RECT 60.376 164.936 60.912 167.508 ; 
        RECT 60.376 163.134 60.768 167.508 ; 
        RECT 58.708 163.134 59.04 167.508 ; 
        RECT 58.708 163.488 59.096 167.23 ; 
        RECT 121.072 163.134 121.412 167.508 ; 
        RECT 120.496 163.134 120.6 167.508 ; 
        RECT 120.064 163.134 120.168 167.508 ; 
        RECT 119.632 163.134 119.736 167.508 ; 
        RECT 119.2 163.134 119.304 167.508 ; 
        RECT 118.768 163.134 118.872 167.508 ; 
        RECT 118.336 163.134 118.44 167.508 ; 
        RECT 117.904 163.134 118.008 167.508 ; 
        RECT 117.472 163.134 117.576 167.508 ; 
        RECT 117.04 163.134 117.144 167.508 ; 
        RECT 116.608 163.134 116.712 167.508 ; 
        RECT 116.176 163.134 116.28 167.508 ; 
        RECT 115.744 163.134 115.848 167.508 ; 
        RECT 115.312 163.134 115.416 167.508 ; 
        RECT 114.88 163.134 114.984 167.508 ; 
        RECT 114.448 163.134 114.552 167.508 ; 
        RECT 114.016 163.134 114.12 167.508 ; 
        RECT 113.584 163.134 113.688 167.508 ; 
        RECT 113.152 163.134 113.256 167.508 ; 
        RECT 112.72 163.134 112.824 167.508 ; 
        RECT 112.288 163.134 112.392 167.508 ; 
        RECT 111.856 163.134 111.96 167.508 ; 
        RECT 111.424 163.134 111.528 167.508 ; 
        RECT 110.992 163.134 111.096 167.508 ; 
        RECT 110.56 163.134 110.664 167.508 ; 
        RECT 110.128 163.134 110.232 167.508 ; 
        RECT 109.696 163.134 109.8 167.508 ; 
        RECT 109.264 163.134 109.368 167.508 ; 
        RECT 108.832 163.134 108.936 167.508 ; 
        RECT 108.4 163.134 108.504 167.508 ; 
        RECT 107.968 163.134 108.072 167.508 ; 
        RECT 107.536 163.134 107.64 167.508 ; 
        RECT 107.104 163.134 107.208 167.508 ; 
        RECT 106.672 163.134 106.776 167.508 ; 
        RECT 106.24 163.134 106.344 167.508 ; 
        RECT 105.808 163.134 105.912 167.508 ; 
        RECT 105.376 163.134 105.48 167.508 ; 
        RECT 104.944 163.134 105.048 167.508 ; 
        RECT 104.512 163.134 104.616 167.508 ; 
        RECT 104.08 163.134 104.184 167.508 ; 
        RECT 103.648 163.134 103.752 167.508 ; 
        RECT 103.216 163.134 103.32 167.508 ; 
        RECT 102.784 163.134 102.888 167.508 ; 
        RECT 102.352 163.134 102.456 167.508 ; 
        RECT 101.92 163.134 102.024 167.508 ; 
        RECT 101.488 163.134 101.592 167.508 ; 
        RECT 101.056 163.134 101.16 167.508 ; 
        RECT 100.624 163.134 100.728 167.508 ; 
        RECT 100.192 163.134 100.296 167.508 ; 
        RECT 99.76 163.134 99.864 167.508 ; 
        RECT 99.328 163.134 99.432 167.508 ; 
        RECT 98.896 163.134 99 167.508 ; 
        RECT 98.464 163.134 98.568 167.508 ; 
        RECT 98.032 163.134 98.136 167.508 ; 
        RECT 97.6 163.134 97.704 167.508 ; 
        RECT 97.168 163.134 97.272 167.508 ; 
        RECT 96.736 163.134 96.84 167.508 ; 
        RECT 96.304 163.134 96.408 167.508 ; 
        RECT 95.872 163.134 95.976 167.508 ; 
        RECT 95.44 163.134 95.544 167.508 ; 
        RECT 95.008 163.134 95.112 167.508 ; 
        RECT 94.576 163.134 94.68 167.508 ; 
        RECT 94.144 163.134 94.248 167.508 ; 
        RECT 93.712 163.134 93.816 167.508 ; 
        RECT 93.28 163.134 93.384 167.508 ; 
        RECT 92.848 163.134 92.952 167.508 ; 
        RECT 92.416 163.134 92.52 167.508 ; 
        RECT 91.984 163.134 92.088 167.508 ; 
        RECT 91.552 163.134 91.656 167.508 ; 
        RECT 91.12 163.134 91.224 167.508 ; 
        RECT 90.688 163.134 90.792 167.508 ; 
        RECT 90.256 163.134 90.36 167.508 ; 
        RECT 89.824 163.134 89.928 167.508 ; 
        RECT 89.392 163.134 89.496 167.508 ; 
        RECT 88.96 163.134 89.064 167.508 ; 
        RECT 88.528 163.134 88.632 167.508 ; 
        RECT 88.096 163.134 88.2 167.508 ; 
        RECT 87.664 163.134 87.768 167.508 ; 
        RECT 87.232 163.134 87.336 167.508 ; 
        RECT 86.8 163.134 86.904 167.508 ; 
        RECT 86.368 163.134 86.472 167.508 ; 
        RECT 85.936 163.134 86.04 167.508 ; 
        RECT 85.504 163.134 85.608 167.508 ; 
        RECT 85.072 163.134 85.176 167.508 ; 
        RECT 84.64 163.134 84.744 167.508 ; 
        RECT 84.208 163.134 84.312 167.508 ; 
        RECT 83.776 163.134 83.88 167.508 ; 
        RECT 83.344 163.134 83.448 167.508 ; 
        RECT 82.912 163.134 83.016 167.508 ; 
        RECT 82.48 163.134 82.584 167.508 ; 
        RECT 82.048 163.134 82.152 167.508 ; 
        RECT 81.616 163.134 81.72 167.508 ; 
        RECT 81.184 163.134 81.288 167.508 ; 
        RECT 80.752 163.134 80.856 167.508 ; 
        RECT 80.32 163.134 80.424 167.508 ; 
        RECT 79.888 163.134 79.992 167.508 ; 
        RECT 79.456 163.134 79.56 167.508 ; 
        RECT 79.024 163.134 79.128 167.508 ; 
        RECT 78.592 163.134 78.696 167.508 ; 
        RECT 78.16 163.134 78.264 167.508 ; 
        RECT 77.728 163.134 77.832 167.508 ; 
        RECT 77.296 163.134 77.4 167.508 ; 
        RECT 76.864 163.134 76.968 167.508 ; 
        RECT 76.432 163.134 76.536 167.508 ; 
        RECT 76 163.134 76.104 167.508 ; 
        RECT 75.568 163.134 75.672 167.508 ; 
        RECT 75.136 163.134 75.24 167.508 ; 
        RECT 74.704 163.134 74.808 167.508 ; 
        RECT 74.272 163.134 74.376 167.508 ; 
        RECT 73.84 163.134 73.944 167.508 ; 
        RECT 73.408 163.134 73.512 167.508 ; 
        RECT 72.976 163.134 73.08 167.508 ; 
        RECT 72.544 163.134 72.648 167.508 ; 
        RECT 72.112 163.134 72.216 167.508 ; 
        RECT 71.68 163.134 71.784 167.508 ; 
        RECT 71.248 163.134 71.352 167.508 ; 
        RECT 70.816 163.134 70.92 167.508 ; 
        RECT 70.384 163.134 70.488 167.508 ; 
        RECT 69.952 163.134 70.056 167.508 ; 
        RECT 69.52 163.134 69.624 167.508 ; 
        RECT 69.088 163.134 69.192 167.508 ; 
        RECT 68.656 163.134 68.76 167.508 ; 
        RECT 68.224 163.134 68.328 167.508 ; 
        RECT 67.792 163.134 67.896 167.508 ; 
        RECT 67.36 163.134 67.464 167.508 ; 
        RECT 66.928 163.134 67.032 167.508 ; 
        RECT 66.496 163.134 66.6 167.508 ; 
        RECT 66.064 163.134 66.168 167.508 ; 
        RECT 65.632 163.134 65.736 167.508 ; 
        RECT 65.2 163.134 65.304 167.508 ; 
        RECT 64.348 163.134 64.656 167.508 ; 
        RECT 56.776 163.134 57.084 167.508 ; 
        RECT 56.128 163.134 56.232 167.508 ; 
        RECT 55.696 163.134 55.8 167.508 ; 
        RECT 55.264 163.134 55.368 167.508 ; 
        RECT 54.832 163.134 54.936 167.508 ; 
        RECT 54.4 163.134 54.504 167.508 ; 
        RECT 53.968 163.134 54.072 167.508 ; 
        RECT 53.536 163.134 53.64 167.508 ; 
        RECT 53.104 163.134 53.208 167.508 ; 
        RECT 52.672 163.134 52.776 167.508 ; 
        RECT 52.24 163.134 52.344 167.508 ; 
        RECT 51.808 163.134 51.912 167.508 ; 
        RECT 51.376 163.134 51.48 167.508 ; 
        RECT 50.944 163.134 51.048 167.508 ; 
        RECT 50.512 163.134 50.616 167.508 ; 
        RECT 50.08 163.134 50.184 167.508 ; 
        RECT 49.648 163.134 49.752 167.508 ; 
        RECT 49.216 163.134 49.32 167.508 ; 
        RECT 48.784 163.134 48.888 167.508 ; 
        RECT 48.352 163.134 48.456 167.508 ; 
        RECT 47.92 163.134 48.024 167.508 ; 
        RECT 47.488 163.134 47.592 167.508 ; 
        RECT 47.056 163.134 47.16 167.508 ; 
        RECT 46.624 163.134 46.728 167.508 ; 
        RECT 46.192 163.134 46.296 167.508 ; 
        RECT 45.76 163.134 45.864 167.508 ; 
        RECT 45.328 163.134 45.432 167.508 ; 
        RECT 44.896 163.134 45 167.508 ; 
        RECT 44.464 163.134 44.568 167.508 ; 
        RECT 44.032 163.134 44.136 167.508 ; 
        RECT 43.6 163.134 43.704 167.508 ; 
        RECT 43.168 163.134 43.272 167.508 ; 
        RECT 42.736 163.134 42.84 167.508 ; 
        RECT 42.304 163.134 42.408 167.508 ; 
        RECT 41.872 163.134 41.976 167.508 ; 
        RECT 41.44 163.134 41.544 167.508 ; 
        RECT 41.008 163.134 41.112 167.508 ; 
        RECT 40.576 163.134 40.68 167.508 ; 
        RECT 40.144 163.134 40.248 167.508 ; 
        RECT 39.712 163.134 39.816 167.508 ; 
        RECT 39.28 163.134 39.384 167.508 ; 
        RECT 38.848 163.134 38.952 167.508 ; 
        RECT 38.416 163.134 38.52 167.508 ; 
        RECT 37.984 163.134 38.088 167.508 ; 
        RECT 37.552 163.134 37.656 167.508 ; 
        RECT 37.12 163.134 37.224 167.508 ; 
        RECT 36.688 163.134 36.792 167.508 ; 
        RECT 36.256 163.134 36.36 167.508 ; 
        RECT 35.824 163.134 35.928 167.508 ; 
        RECT 35.392 163.134 35.496 167.508 ; 
        RECT 34.96 163.134 35.064 167.508 ; 
        RECT 34.528 163.134 34.632 167.508 ; 
        RECT 34.096 163.134 34.2 167.508 ; 
        RECT 33.664 163.134 33.768 167.508 ; 
        RECT 33.232 163.134 33.336 167.508 ; 
        RECT 32.8 163.134 32.904 167.508 ; 
        RECT 32.368 163.134 32.472 167.508 ; 
        RECT 31.936 163.134 32.04 167.508 ; 
        RECT 31.504 163.134 31.608 167.508 ; 
        RECT 31.072 163.134 31.176 167.508 ; 
        RECT 30.64 163.134 30.744 167.508 ; 
        RECT 30.208 163.134 30.312 167.508 ; 
        RECT 29.776 163.134 29.88 167.508 ; 
        RECT 29.344 163.134 29.448 167.508 ; 
        RECT 28.912 163.134 29.016 167.508 ; 
        RECT 28.48 163.134 28.584 167.508 ; 
        RECT 28.048 163.134 28.152 167.508 ; 
        RECT 27.616 163.134 27.72 167.508 ; 
        RECT 27.184 163.134 27.288 167.508 ; 
        RECT 26.752 163.134 26.856 167.508 ; 
        RECT 26.32 163.134 26.424 167.508 ; 
        RECT 25.888 163.134 25.992 167.508 ; 
        RECT 25.456 163.134 25.56 167.508 ; 
        RECT 25.024 163.134 25.128 167.508 ; 
        RECT 24.592 163.134 24.696 167.508 ; 
        RECT 24.16 163.134 24.264 167.508 ; 
        RECT 23.728 163.134 23.832 167.508 ; 
        RECT 23.296 163.134 23.4 167.508 ; 
        RECT 22.864 163.134 22.968 167.508 ; 
        RECT 22.432 163.134 22.536 167.508 ; 
        RECT 22 163.134 22.104 167.508 ; 
        RECT 21.568 163.134 21.672 167.508 ; 
        RECT 21.136 163.134 21.24 167.508 ; 
        RECT 20.704 163.134 20.808 167.508 ; 
        RECT 20.272 163.134 20.376 167.508 ; 
        RECT 19.84 163.134 19.944 167.508 ; 
        RECT 19.408 163.134 19.512 167.508 ; 
        RECT 18.976 163.134 19.08 167.508 ; 
        RECT 18.544 163.134 18.648 167.508 ; 
        RECT 18.112 163.134 18.216 167.508 ; 
        RECT 17.68 163.134 17.784 167.508 ; 
        RECT 17.248 163.134 17.352 167.508 ; 
        RECT 16.816 163.134 16.92 167.508 ; 
        RECT 16.384 163.134 16.488 167.508 ; 
        RECT 15.952 163.134 16.056 167.508 ; 
        RECT 15.52 163.134 15.624 167.508 ; 
        RECT 15.088 163.134 15.192 167.508 ; 
        RECT 14.656 163.134 14.76 167.508 ; 
        RECT 14.224 163.134 14.328 167.508 ; 
        RECT 13.792 163.134 13.896 167.508 ; 
        RECT 13.36 163.134 13.464 167.508 ; 
        RECT 12.928 163.134 13.032 167.508 ; 
        RECT 12.496 163.134 12.6 167.508 ; 
        RECT 12.064 163.134 12.168 167.508 ; 
        RECT 11.632 163.134 11.736 167.508 ; 
        RECT 11.2 163.134 11.304 167.508 ; 
        RECT 10.768 163.134 10.872 167.508 ; 
        RECT 10.336 163.134 10.44 167.508 ; 
        RECT 9.904 163.134 10.008 167.508 ; 
        RECT 9.472 163.134 9.576 167.508 ; 
        RECT 9.04 163.134 9.144 167.508 ; 
        RECT 8.608 163.134 8.712 167.508 ; 
        RECT 8.176 163.134 8.28 167.508 ; 
        RECT 7.744 163.134 7.848 167.508 ; 
        RECT 7.312 163.134 7.416 167.508 ; 
        RECT 6.88 163.134 6.984 167.508 ; 
        RECT 6.448 163.134 6.552 167.508 ; 
        RECT 6.016 163.134 6.12 167.508 ; 
        RECT 5.584 163.134 5.688 167.508 ; 
        RECT 5.152 163.134 5.256 167.508 ; 
        RECT 4.72 163.134 4.824 167.508 ; 
        RECT 4.288 163.134 4.392 167.508 ; 
        RECT 3.856 163.134 3.96 167.508 ; 
        RECT 3.424 163.134 3.528 167.508 ; 
        RECT 2.992 163.134 3.096 167.508 ; 
        RECT 2.56 163.134 2.664 167.508 ; 
        RECT 2.128 163.134 2.232 167.508 ; 
        RECT 1.696 163.134 1.8 167.508 ; 
        RECT 1.264 163.134 1.368 167.508 ; 
        RECT 0.832 163.134 0.936 167.508 ; 
        RECT 0.02 163.134 0.36 167.508 ; 
        RECT 62.212 167.454 62.724 171.828 ; 
        RECT 62.156 170.116 62.724 171.406 ; 
        RECT 61.276 169.024 61.812 171.828 ; 
        RECT 61.184 170.364 61.812 171.396 ; 
        RECT 61.276 167.454 61.668 171.828 ; 
        RECT 61.276 167.938 61.724 168.896 ; 
        RECT 61.276 167.454 61.812 167.81 ; 
        RECT 60.376 169.256 60.912 171.828 ; 
        RECT 60.376 167.454 60.768 171.828 ; 
        RECT 58.708 167.454 59.04 171.828 ; 
        RECT 58.708 167.808 59.096 171.55 ; 
        RECT 121.072 167.454 121.412 171.828 ; 
        RECT 120.496 167.454 120.6 171.828 ; 
        RECT 120.064 167.454 120.168 171.828 ; 
        RECT 119.632 167.454 119.736 171.828 ; 
        RECT 119.2 167.454 119.304 171.828 ; 
        RECT 118.768 167.454 118.872 171.828 ; 
        RECT 118.336 167.454 118.44 171.828 ; 
        RECT 117.904 167.454 118.008 171.828 ; 
        RECT 117.472 167.454 117.576 171.828 ; 
        RECT 117.04 167.454 117.144 171.828 ; 
        RECT 116.608 167.454 116.712 171.828 ; 
        RECT 116.176 167.454 116.28 171.828 ; 
        RECT 115.744 167.454 115.848 171.828 ; 
        RECT 115.312 167.454 115.416 171.828 ; 
        RECT 114.88 167.454 114.984 171.828 ; 
        RECT 114.448 167.454 114.552 171.828 ; 
        RECT 114.016 167.454 114.12 171.828 ; 
        RECT 113.584 167.454 113.688 171.828 ; 
        RECT 113.152 167.454 113.256 171.828 ; 
        RECT 112.72 167.454 112.824 171.828 ; 
        RECT 112.288 167.454 112.392 171.828 ; 
        RECT 111.856 167.454 111.96 171.828 ; 
        RECT 111.424 167.454 111.528 171.828 ; 
        RECT 110.992 167.454 111.096 171.828 ; 
        RECT 110.56 167.454 110.664 171.828 ; 
        RECT 110.128 167.454 110.232 171.828 ; 
        RECT 109.696 167.454 109.8 171.828 ; 
        RECT 109.264 167.454 109.368 171.828 ; 
        RECT 108.832 167.454 108.936 171.828 ; 
        RECT 108.4 167.454 108.504 171.828 ; 
        RECT 107.968 167.454 108.072 171.828 ; 
        RECT 107.536 167.454 107.64 171.828 ; 
        RECT 107.104 167.454 107.208 171.828 ; 
        RECT 106.672 167.454 106.776 171.828 ; 
        RECT 106.24 167.454 106.344 171.828 ; 
        RECT 105.808 167.454 105.912 171.828 ; 
        RECT 105.376 167.454 105.48 171.828 ; 
        RECT 104.944 167.454 105.048 171.828 ; 
        RECT 104.512 167.454 104.616 171.828 ; 
        RECT 104.08 167.454 104.184 171.828 ; 
        RECT 103.648 167.454 103.752 171.828 ; 
        RECT 103.216 167.454 103.32 171.828 ; 
        RECT 102.784 167.454 102.888 171.828 ; 
        RECT 102.352 167.454 102.456 171.828 ; 
        RECT 101.92 167.454 102.024 171.828 ; 
        RECT 101.488 167.454 101.592 171.828 ; 
        RECT 101.056 167.454 101.16 171.828 ; 
        RECT 100.624 167.454 100.728 171.828 ; 
        RECT 100.192 167.454 100.296 171.828 ; 
        RECT 99.76 167.454 99.864 171.828 ; 
        RECT 99.328 167.454 99.432 171.828 ; 
        RECT 98.896 167.454 99 171.828 ; 
        RECT 98.464 167.454 98.568 171.828 ; 
        RECT 98.032 167.454 98.136 171.828 ; 
        RECT 97.6 167.454 97.704 171.828 ; 
        RECT 97.168 167.454 97.272 171.828 ; 
        RECT 96.736 167.454 96.84 171.828 ; 
        RECT 96.304 167.454 96.408 171.828 ; 
        RECT 95.872 167.454 95.976 171.828 ; 
        RECT 95.44 167.454 95.544 171.828 ; 
        RECT 95.008 167.454 95.112 171.828 ; 
        RECT 94.576 167.454 94.68 171.828 ; 
        RECT 94.144 167.454 94.248 171.828 ; 
        RECT 93.712 167.454 93.816 171.828 ; 
        RECT 93.28 167.454 93.384 171.828 ; 
        RECT 92.848 167.454 92.952 171.828 ; 
        RECT 92.416 167.454 92.52 171.828 ; 
        RECT 91.984 167.454 92.088 171.828 ; 
        RECT 91.552 167.454 91.656 171.828 ; 
        RECT 91.12 167.454 91.224 171.828 ; 
        RECT 90.688 167.454 90.792 171.828 ; 
        RECT 90.256 167.454 90.36 171.828 ; 
        RECT 89.824 167.454 89.928 171.828 ; 
        RECT 89.392 167.454 89.496 171.828 ; 
        RECT 88.96 167.454 89.064 171.828 ; 
        RECT 88.528 167.454 88.632 171.828 ; 
        RECT 88.096 167.454 88.2 171.828 ; 
        RECT 87.664 167.454 87.768 171.828 ; 
        RECT 87.232 167.454 87.336 171.828 ; 
        RECT 86.8 167.454 86.904 171.828 ; 
        RECT 86.368 167.454 86.472 171.828 ; 
        RECT 85.936 167.454 86.04 171.828 ; 
        RECT 85.504 167.454 85.608 171.828 ; 
        RECT 85.072 167.454 85.176 171.828 ; 
        RECT 84.64 167.454 84.744 171.828 ; 
        RECT 84.208 167.454 84.312 171.828 ; 
        RECT 83.776 167.454 83.88 171.828 ; 
        RECT 83.344 167.454 83.448 171.828 ; 
        RECT 82.912 167.454 83.016 171.828 ; 
        RECT 82.48 167.454 82.584 171.828 ; 
        RECT 82.048 167.454 82.152 171.828 ; 
        RECT 81.616 167.454 81.72 171.828 ; 
        RECT 81.184 167.454 81.288 171.828 ; 
        RECT 80.752 167.454 80.856 171.828 ; 
        RECT 80.32 167.454 80.424 171.828 ; 
        RECT 79.888 167.454 79.992 171.828 ; 
        RECT 79.456 167.454 79.56 171.828 ; 
        RECT 79.024 167.454 79.128 171.828 ; 
        RECT 78.592 167.454 78.696 171.828 ; 
        RECT 78.16 167.454 78.264 171.828 ; 
        RECT 77.728 167.454 77.832 171.828 ; 
        RECT 77.296 167.454 77.4 171.828 ; 
        RECT 76.864 167.454 76.968 171.828 ; 
        RECT 76.432 167.454 76.536 171.828 ; 
        RECT 76 167.454 76.104 171.828 ; 
        RECT 75.568 167.454 75.672 171.828 ; 
        RECT 75.136 167.454 75.24 171.828 ; 
        RECT 74.704 167.454 74.808 171.828 ; 
        RECT 74.272 167.454 74.376 171.828 ; 
        RECT 73.84 167.454 73.944 171.828 ; 
        RECT 73.408 167.454 73.512 171.828 ; 
        RECT 72.976 167.454 73.08 171.828 ; 
        RECT 72.544 167.454 72.648 171.828 ; 
        RECT 72.112 167.454 72.216 171.828 ; 
        RECT 71.68 167.454 71.784 171.828 ; 
        RECT 71.248 167.454 71.352 171.828 ; 
        RECT 70.816 167.454 70.92 171.828 ; 
        RECT 70.384 167.454 70.488 171.828 ; 
        RECT 69.952 167.454 70.056 171.828 ; 
        RECT 69.52 167.454 69.624 171.828 ; 
        RECT 69.088 167.454 69.192 171.828 ; 
        RECT 68.656 167.454 68.76 171.828 ; 
        RECT 68.224 167.454 68.328 171.828 ; 
        RECT 67.792 167.454 67.896 171.828 ; 
        RECT 67.36 167.454 67.464 171.828 ; 
        RECT 66.928 167.454 67.032 171.828 ; 
        RECT 66.496 167.454 66.6 171.828 ; 
        RECT 66.064 167.454 66.168 171.828 ; 
        RECT 65.632 167.454 65.736 171.828 ; 
        RECT 65.2 167.454 65.304 171.828 ; 
        RECT 64.348 167.454 64.656 171.828 ; 
        RECT 56.776 167.454 57.084 171.828 ; 
        RECT 56.128 167.454 56.232 171.828 ; 
        RECT 55.696 167.454 55.8 171.828 ; 
        RECT 55.264 167.454 55.368 171.828 ; 
        RECT 54.832 167.454 54.936 171.828 ; 
        RECT 54.4 167.454 54.504 171.828 ; 
        RECT 53.968 167.454 54.072 171.828 ; 
        RECT 53.536 167.454 53.64 171.828 ; 
        RECT 53.104 167.454 53.208 171.828 ; 
        RECT 52.672 167.454 52.776 171.828 ; 
        RECT 52.24 167.454 52.344 171.828 ; 
        RECT 51.808 167.454 51.912 171.828 ; 
        RECT 51.376 167.454 51.48 171.828 ; 
        RECT 50.944 167.454 51.048 171.828 ; 
        RECT 50.512 167.454 50.616 171.828 ; 
        RECT 50.08 167.454 50.184 171.828 ; 
        RECT 49.648 167.454 49.752 171.828 ; 
        RECT 49.216 167.454 49.32 171.828 ; 
        RECT 48.784 167.454 48.888 171.828 ; 
        RECT 48.352 167.454 48.456 171.828 ; 
        RECT 47.92 167.454 48.024 171.828 ; 
        RECT 47.488 167.454 47.592 171.828 ; 
        RECT 47.056 167.454 47.16 171.828 ; 
        RECT 46.624 167.454 46.728 171.828 ; 
        RECT 46.192 167.454 46.296 171.828 ; 
        RECT 45.76 167.454 45.864 171.828 ; 
        RECT 45.328 167.454 45.432 171.828 ; 
        RECT 44.896 167.454 45 171.828 ; 
        RECT 44.464 167.454 44.568 171.828 ; 
        RECT 44.032 167.454 44.136 171.828 ; 
        RECT 43.6 167.454 43.704 171.828 ; 
        RECT 43.168 167.454 43.272 171.828 ; 
        RECT 42.736 167.454 42.84 171.828 ; 
        RECT 42.304 167.454 42.408 171.828 ; 
        RECT 41.872 167.454 41.976 171.828 ; 
        RECT 41.44 167.454 41.544 171.828 ; 
        RECT 41.008 167.454 41.112 171.828 ; 
        RECT 40.576 167.454 40.68 171.828 ; 
        RECT 40.144 167.454 40.248 171.828 ; 
        RECT 39.712 167.454 39.816 171.828 ; 
        RECT 39.28 167.454 39.384 171.828 ; 
        RECT 38.848 167.454 38.952 171.828 ; 
        RECT 38.416 167.454 38.52 171.828 ; 
        RECT 37.984 167.454 38.088 171.828 ; 
        RECT 37.552 167.454 37.656 171.828 ; 
        RECT 37.12 167.454 37.224 171.828 ; 
        RECT 36.688 167.454 36.792 171.828 ; 
        RECT 36.256 167.454 36.36 171.828 ; 
        RECT 35.824 167.454 35.928 171.828 ; 
        RECT 35.392 167.454 35.496 171.828 ; 
        RECT 34.96 167.454 35.064 171.828 ; 
        RECT 34.528 167.454 34.632 171.828 ; 
        RECT 34.096 167.454 34.2 171.828 ; 
        RECT 33.664 167.454 33.768 171.828 ; 
        RECT 33.232 167.454 33.336 171.828 ; 
        RECT 32.8 167.454 32.904 171.828 ; 
        RECT 32.368 167.454 32.472 171.828 ; 
        RECT 31.936 167.454 32.04 171.828 ; 
        RECT 31.504 167.454 31.608 171.828 ; 
        RECT 31.072 167.454 31.176 171.828 ; 
        RECT 30.64 167.454 30.744 171.828 ; 
        RECT 30.208 167.454 30.312 171.828 ; 
        RECT 29.776 167.454 29.88 171.828 ; 
        RECT 29.344 167.454 29.448 171.828 ; 
        RECT 28.912 167.454 29.016 171.828 ; 
        RECT 28.48 167.454 28.584 171.828 ; 
        RECT 28.048 167.454 28.152 171.828 ; 
        RECT 27.616 167.454 27.72 171.828 ; 
        RECT 27.184 167.454 27.288 171.828 ; 
        RECT 26.752 167.454 26.856 171.828 ; 
        RECT 26.32 167.454 26.424 171.828 ; 
        RECT 25.888 167.454 25.992 171.828 ; 
        RECT 25.456 167.454 25.56 171.828 ; 
        RECT 25.024 167.454 25.128 171.828 ; 
        RECT 24.592 167.454 24.696 171.828 ; 
        RECT 24.16 167.454 24.264 171.828 ; 
        RECT 23.728 167.454 23.832 171.828 ; 
        RECT 23.296 167.454 23.4 171.828 ; 
        RECT 22.864 167.454 22.968 171.828 ; 
        RECT 22.432 167.454 22.536 171.828 ; 
        RECT 22 167.454 22.104 171.828 ; 
        RECT 21.568 167.454 21.672 171.828 ; 
        RECT 21.136 167.454 21.24 171.828 ; 
        RECT 20.704 167.454 20.808 171.828 ; 
        RECT 20.272 167.454 20.376 171.828 ; 
        RECT 19.84 167.454 19.944 171.828 ; 
        RECT 19.408 167.454 19.512 171.828 ; 
        RECT 18.976 167.454 19.08 171.828 ; 
        RECT 18.544 167.454 18.648 171.828 ; 
        RECT 18.112 167.454 18.216 171.828 ; 
        RECT 17.68 167.454 17.784 171.828 ; 
        RECT 17.248 167.454 17.352 171.828 ; 
        RECT 16.816 167.454 16.92 171.828 ; 
        RECT 16.384 167.454 16.488 171.828 ; 
        RECT 15.952 167.454 16.056 171.828 ; 
        RECT 15.52 167.454 15.624 171.828 ; 
        RECT 15.088 167.454 15.192 171.828 ; 
        RECT 14.656 167.454 14.76 171.828 ; 
        RECT 14.224 167.454 14.328 171.828 ; 
        RECT 13.792 167.454 13.896 171.828 ; 
        RECT 13.36 167.454 13.464 171.828 ; 
        RECT 12.928 167.454 13.032 171.828 ; 
        RECT 12.496 167.454 12.6 171.828 ; 
        RECT 12.064 167.454 12.168 171.828 ; 
        RECT 11.632 167.454 11.736 171.828 ; 
        RECT 11.2 167.454 11.304 171.828 ; 
        RECT 10.768 167.454 10.872 171.828 ; 
        RECT 10.336 167.454 10.44 171.828 ; 
        RECT 9.904 167.454 10.008 171.828 ; 
        RECT 9.472 167.454 9.576 171.828 ; 
        RECT 9.04 167.454 9.144 171.828 ; 
        RECT 8.608 167.454 8.712 171.828 ; 
        RECT 8.176 167.454 8.28 171.828 ; 
        RECT 7.744 167.454 7.848 171.828 ; 
        RECT 7.312 167.454 7.416 171.828 ; 
        RECT 6.88 167.454 6.984 171.828 ; 
        RECT 6.448 167.454 6.552 171.828 ; 
        RECT 6.016 167.454 6.12 171.828 ; 
        RECT 5.584 167.454 5.688 171.828 ; 
        RECT 5.152 167.454 5.256 171.828 ; 
        RECT 4.72 167.454 4.824 171.828 ; 
        RECT 4.288 167.454 4.392 171.828 ; 
        RECT 3.856 167.454 3.96 171.828 ; 
        RECT 3.424 167.454 3.528 171.828 ; 
        RECT 2.992 167.454 3.096 171.828 ; 
        RECT 2.56 167.454 2.664 171.828 ; 
        RECT 2.128 167.454 2.232 171.828 ; 
        RECT 1.696 167.454 1.8 171.828 ; 
        RECT 1.264 167.454 1.368 171.828 ; 
        RECT 0.832 167.454 0.936 171.828 ; 
        RECT 0.02 167.454 0.36 171.828 ; 
        RECT 62.212 171.774 62.724 176.148 ; 
        RECT 62.156 174.436 62.724 175.726 ; 
        RECT 61.276 173.344 61.812 176.148 ; 
        RECT 61.184 174.684 61.812 175.716 ; 
        RECT 61.276 171.774 61.668 176.148 ; 
        RECT 61.276 172.258 61.724 173.216 ; 
        RECT 61.276 171.774 61.812 172.13 ; 
        RECT 60.376 173.576 60.912 176.148 ; 
        RECT 60.376 171.774 60.768 176.148 ; 
        RECT 58.708 171.774 59.04 176.148 ; 
        RECT 58.708 172.128 59.096 175.87 ; 
        RECT 121.072 171.774 121.412 176.148 ; 
        RECT 120.496 171.774 120.6 176.148 ; 
        RECT 120.064 171.774 120.168 176.148 ; 
        RECT 119.632 171.774 119.736 176.148 ; 
        RECT 119.2 171.774 119.304 176.148 ; 
        RECT 118.768 171.774 118.872 176.148 ; 
        RECT 118.336 171.774 118.44 176.148 ; 
        RECT 117.904 171.774 118.008 176.148 ; 
        RECT 117.472 171.774 117.576 176.148 ; 
        RECT 117.04 171.774 117.144 176.148 ; 
        RECT 116.608 171.774 116.712 176.148 ; 
        RECT 116.176 171.774 116.28 176.148 ; 
        RECT 115.744 171.774 115.848 176.148 ; 
        RECT 115.312 171.774 115.416 176.148 ; 
        RECT 114.88 171.774 114.984 176.148 ; 
        RECT 114.448 171.774 114.552 176.148 ; 
        RECT 114.016 171.774 114.12 176.148 ; 
        RECT 113.584 171.774 113.688 176.148 ; 
        RECT 113.152 171.774 113.256 176.148 ; 
        RECT 112.72 171.774 112.824 176.148 ; 
        RECT 112.288 171.774 112.392 176.148 ; 
        RECT 111.856 171.774 111.96 176.148 ; 
        RECT 111.424 171.774 111.528 176.148 ; 
        RECT 110.992 171.774 111.096 176.148 ; 
        RECT 110.56 171.774 110.664 176.148 ; 
        RECT 110.128 171.774 110.232 176.148 ; 
        RECT 109.696 171.774 109.8 176.148 ; 
        RECT 109.264 171.774 109.368 176.148 ; 
        RECT 108.832 171.774 108.936 176.148 ; 
        RECT 108.4 171.774 108.504 176.148 ; 
        RECT 107.968 171.774 108.072 176.148 ; 
        RECT 107.536 171.774 107.64 176.148 ; 
        RECT 107.104 171.774 107.208 176.148 ; 
        RECT 106.672 171.774 106.776 176.148 ; 
        RECT 106.24 171.774 106.344 176.148 ; 
        RECT 105.808 171.774 105.912 176.148 ; 
        RECT 105.376 171.774 105.48 176.148 ; 
        RECT 104.944 171.774 105.048 176.148 ; 
        RECT 104.512 171.774 104.616 176.148 ; 
        RECT 104.08 171.774 104.184 176.148 ; 
        RECT 103.648 171.774 103.752 176.148 ; 
        RECT 103.216 171.774 103.32 176.148 ; 
        RECT 102.784 171.774 102.888 176.148 ; 
        RECT 102.352 171.774 102.456 176.148 ; 
        RECT 101.92 171.774 102.024 176.148 ; 
        RECT 101.488 171.774 101.592 176.148 ; 
        RECT 101.056 171.774 101.16 176.148 ; 
        RECT 100.624 171.774 100.728 176.148 ; 
        RECT 100.192 171.774 100.296 176.148 ; 
        RECT 99.76 171.774 99.864 176.148 ; 
        RECT 99.328 171.774 99.432 176.148 ; 
        RECT 98.896 171.774 99 176.148 ; 
        RECT 98.464 171.774 98.568 176.148 ; 
        RECT 98.032 171.774 98.136 176.148 ; 
        RECT 97.6 171.774 97.704 176.148 ; 
        RECT 97.168 171.774 97.272 176.148 ; 
        RECT 96.736 171.774 96.84 176.148 ; 
        RECT 96.304 171.774 96.408 176.148 ; 
        RECT 95.872 171.774 95.976 176.148 ; 
        RECT 95.44 171.774 95.544 176.148 ; 
        RECT 95.008 171.774 95.112 176.148 ; 
        RECT 94.576 171.774 94.68 176.148 ; 
        RECT 94.144 171.774 94.248 176.148 ; 
        RECT 93.712 171.774 93.816 176.148 ; 
        RECT 93.28 171.774 93.384 176.148 ; 
        RECT 92.848 171.774 92.952 176.148 ; 
        RECT 92.416 171.774 92.52 176.148 ; 
        RECT 91.984 171.774 92.088 176.148 ; 
        RECT 91.552 171.774 91.656 176.148 ; 
        RECT 91.12 171.774 91.224 176.148 ; 
        RECT 90.688 171.774 90.792 176.148 ; 
        RECT 90.256 171.774 90.36 176.148 ; 
        RECT 89.824 171.774 89.928 176.148 ; 
        RECT 89.392 171.774 89.496 176.148 ; 
        RECT 88.96 171.774 89.064 176.148 ; 
        RECT 88.528 171.774 88.632 176.148 ; 
        RECT 88.096 171.774 88.2 176.148 ; 
        RECT 87.664 171.774 87.768 176.148 ; 
        RECT 87.232 171.774 87.336 176.148 ; 
        RECT 86.8 171.774 86.904 176.148 ; 
        RECT 86.368 171.774 86.472 176.148 ; 
        RECT 85.936 171.774 86.04 176.148 ; 
        RECT 85.504 171.774 85.608 176.148 ; 
        RECT 85.072 171.774 85.176 176.148 ; 
        RECT 84.64 171.774 84.744 176.148 ; 
        RECT 84.208 171.774 84.312 176.148 ; 
        RECT 83.776 171.774 83.88 176.148 ; 
        RECT 83.344 171.774 83.448 176.148 ; 
        RECT 82.912 171.774 83.016 176.148 ; 
        RECT 82.48 171.774 82.584 176.148 ; 
        RECT 82.048 171.774 82.152 176.148 ; 
        RECT 81.616 171.774 81.72 176.148 ; 
        RECT 81.184 171.774 81.288 176.148 ; 
        RECT 80.752 171.774 80.856 176.148 ; 
        RECT 80.32 171.774 80.424 176.148 ; 
        RECT 79.888 171.774 79.992 176.148 ; 
        RECT 79.456 171.774 79.56 176.148 ; 
        RECT 79.024 171.774 79.128 176.148 ; 
        RECT 78.592 171.774 78.696 176.148 ; 
        RECT 78.16 171.774 78.264 176.148 ; 
        RECT 77.728 171.774 77.832 176.148 ; 
        RECT 77.296 171.774 77.4 176.148 ; 
        RECT 76.864 171.774 76.968 176.148 ; 
        RECT 76.432 171.774 76.536 176.148 ; 
        RECT 76 171.774 76.104 176.148 ; 
        RECT 75.568 171.774 75.672 176.148 ; 
        RECT 75.136 171.774 75.24 176.148 ; 
        RECT 74.704 171.774 74.808 176.148 ; 
        RECT 74.272 171.774 74.376 176.148 ; 
        RECT 73.84 171.774 73.944 176.148 ; 
        RECT 73.408 171.774 73.512 176.148 ; 
        RECT 72.976 171.774 73.08 176.148 ; 
        RECT 72.544 171.774 72.648 176.148 ; 
        RECT 72.112 171.774 72.216 176.148 ; 
        RECT 71.68 171.774 71.784 176.148 ; 
        RECT 71.248 171.774 71.352 176.148 ; 
        RECT 70.816 171.774 70.92 176.148 ; 
        RECT 70.384 171.774 70.488 176.148 ; 
        RECT 69.952 171.774 70.056 176.148 ; 
        RECT 69.52 171.774 69.624 176.148 ; 
        RECT 69.088 171.774 69.192 176.148 ; 
        RECT 68.656 171.774 68.76 176.148 ; 
        RECT 68.224 171.774 68.328 176.148 ; 
        RECT 67.792 171.774 67.896 176.148 ; 
        RECT 67.36 171.774 67.464 176.148 ; 
        RECT 66.928 171.774 67.032 176.148 ; 
        RECT 66.496 171.774 66.6 176.148 ; 
        RECT 66.064 171.774 66.168 176.148 ; 
        RECT 65.632 171.774 65.736 176.148 ; 
        RECT 65.2 171.774 65.304 176.148 ; 
        RECT 64.348 171.774 64.656 176.148 ; 
        RECT 56.776 171.774 57.084 176.148 ; 
        RECT 56.128 171.774 56.232 176.148 ; 
        RECT 55.696 171.774 55.8 176.148 ; 
        RECT 55.264 171.774 55.368 176.148 ; 
        RECT 54.832 171.774 54.936 176.148 ; 
        RECT 54.4 171.774 54.504 176.148 ; 
        RECT 53.968 171.774 54.072 176.148 ; 
        RECT 53.536 171.774 53.64 176.148 ; 
        RECT 53.104 171.774 53.208 176.148 ; 
        RECT 52.672 171.774 52.776 176.148 ; 
        RECT 52.24 171.774 52.344 176.148 ; 
        RECT 51.808 171.774 51.912 176.148 ; 
        RECT 51.376 171.774 51.48 176.148 ; 
        RECT 50.944 171.774 51.048 176.148 ; 
        RECT 50.512 171.774 50.616 176.148 ; 
        RECT 50.08 171.774 50.184 176.148 ; 
        RECT 49.648 171.774 49.752 176.148 ; 
        RECT 49.216 171.774 49.32 176.148 ; 
        RECT 48.784 171.774 48.888 176.148 ; 
        RECT 48.352 171.774 48.456 176.148 ; 
        RECT 47.92 171.774 48.024 176.148 ; 
        RECT 47.488 171.774 47.592 176.148 ; 
        RECT 47.056 171.774 47.16 176.148 ; 
        RECT 46.624 171.774 46.728 176.148 ; 
        RECT 46.192 171.774 46.296 176.148 ; 
        RECT 45.76 171.774 45.864 176.148 ; 
        RECT 45.328 171.774 45.432 176.148 ; 
        RECT 44.896 171.774 45 176.148 ; 
        RECT 44.464 171.774 44.568 176.148 ; 
        RECT 44.032 171.774 44.136 176.148 ; 
        RECT 43.6 171.774 43.704 176.148 ; 
        RECT 43.168 171.774 43.272 176.148 ; 
        RECT 42.736 171.774 42.84 176.148 ; 
        RECT 42.304 171.774 42.408 176.148 ; 
        RECT 41.872 171.774 41.976 176.148 ; 
        RECT 41.44 171.774 41.544 176.148 ; 
        RECT 41.008 171.774 41.112 176.148 ; 
        RECT 40.576 171.774 40.68 176.148 ; 
        RECT 40.144 171.774 40.248 176.148 ; 
        RECT 39.712 171.774 39.816 176.148 ; 
        RECT 39.28 171.774 39.384 176.148 ; 
        RECT 38.848 171.774 38.952 176.148 ; 
        RECT 38.416 171.774 38.52 176.148 ; 
        RECT 37.984 171.774 38.088 176.148 ; 
        RECT 37.552 171.774 37.656 176.148 ; 
        RECT 37.12 171.774 37.224 176.148 ; 
        RECT 36.688 171.774 36.792 176.148 ; 
        RECT 36.256 171.774 36.36 176.148 ; 
        RECT 35.824 171.774 35.928 176.148 ; 
        RECT 35.392 171.774 35.496 176.148 ; 
        RECT 34.96 171.774 35.064 176.148 ; 
        RECT 34.528 171.774 34.632 176.148 ; 
        RECT 34.096 171.774 34.2 176.148 ; 
        RECT 33.664 171.774 33.768 176.148 ; 
        RECT 33.232 171.774 33.336 176.148 ; 
        RECT 32.8 171.774 32.904 176.148 ; 
        RECT 32.368 171.774 32.472 176.148 ; 
        RECT 31.936 171.774 32.04 176.148 ; 
        RECT 31.504 171.774 31.608 176.148 ; 
        RECT 31.072 171.774 31.176 176.148 ; 
        RECT 30.64 171.774 30.744 176.148 ; 
        RECT 30.208 171.774 30.312 176.148 ; 
        RECT 29.776 171.774 29.88 176.148 ; 
        RECT 29.344 171.774 29.448 176.148 ; 
        RECT 28.912 171.774 29.016 176.148 ; 
        RECT 28.48 171.774 28.584 176.148 ; 
        RECT 28.048 171.774 28.152 176.148 ; 
        RECT 27.616 171.774 27.72 176.148 ; 
        RECT 27.184 171.774 27.288 176.148 ; 
        RECT 26.752 171.774 26.856 176.148 ; 
        RECT 26.32 171.774 26.424 176.148 ; 
        RECT 25.888 171.774 25.992 176.148 ; 
        RECT 25.456 171.774 25.56 176.148 ; 
        RECT 25.024 171.774 25.128 176.148 ; 
        RECT 24.592 171.774 24.696 176.148 ; 
        RECT 24.16 171.774 24.264 176.148 ; 
        RECT 23.728 171.774 23.832 176.148 ; 
        RECT 23.296 171.774 23.4 176.148 ; 
        RECT 22.864 171.774 22.968 176.148 ; 
        RECT 22.432 171.774 22.536 176.148 ; 
        RECT 22 171.774 22.104 176.148 ; 
        RECT 21.568 171.774 21.672 176.148 ; 
        RECT 21.136 171.774 21.24 176.148 ; 
        RECT 20.704 171.774 20.808 176.148 ; 
        RECT 20.272 171.774 20.376 176.148 ; 
        RECT 19.84 171.774 19.944 176.148 ; 
        RECT 19.408 171.774 19.512 176.148 ; 
        RECT 18.976 171.774 19.08 176.148 ; 
        RECT 18.544 171.774 18.648 176.148 ; 
        RECT 18.112 171.774 18.216 176.148 ; 
        RECT 17.68 171.774 17.784 176.148 ; 
        RECT 17.248 171.774 17.352 176.148 ; 
        RECT 16.816 171.774 16.92 176.148 ; 
        RECT 16.384 171.774 16.488 176.148 ; 
        RECT 15.952 171.774 16.056 176.148 ; 
        RECT 15.52 171.774 15.624 176.148 ; 
        RECT 15.088 171.774 15.192 176.148 ; 
        RECT 14.656 171.774 14.76 176.148 ; 
        RECT 14.224 171.774 14.328 176.148 ; 
        RECT 13.792 171.774 13.896 176.148 ; 
        RECT 13.36 171.774 13.464 176.148 ; 
        RECT 12.928 171.774 13.032 176.148 ; 
        RECT 12.496 171.774 12.6 176.148 ; 
        RECT 12.064 171.774 12.168 176.148 ; 
        RECT 11.632 171.774 11.736 176.148 ; 
        RECT 11.2 171.774 11.304 176.148 ; 
        RECT 10.768 171.774 10.872 176.148 ; 
        RECT 10.336 171.774 10.44 176.148 ; 
        RECT 9.904 171.774 10.008 176.148 ; 
        RECT 9.472 171.774 9.576 176.148 ; 
        RECT 9.04 171.774 9.144 176.148 ; 
        RECT 8.608 171.774 8.712 176.148 ; 
        RECT 8.176 171.774 8.28 176.148 ; 
        RECT 7.744 171.774 7.848 176.148 ; 
        RECT 7.312 171.774 7.416 176.148 ; 
        RECT 6.88 171.774 6.984 176.148 ; 
        RECT 6.448 171.774 6.552 176.148 ; 
        RECT 6.016 171.774 6.12 176.148 ; 
        RECT 5.584 171.774 5.688 176.148 ; 
        RECT 5.152 171.774 5.256 176.148 ; 
        RECT 4.72 171.774 4.824 176.148 ; 
        RECT 4.288 171.774 4.392 176.148 ; 
        RECT 3.856 171.774 3.96 176.148 ; 
        RECT 3.424 171.774 3.528 176.148 ; 
        RECT 2.992 171.774 3.096 176.148 ; 
        RECT 2.56 171.774 2.664 176.148 ; 
        RECT 2.128 171.774 2.232 176.148 ; 
        RECT 1.696 171.774 1.8 176.148 ; 
        RECT 1.264 171.774 1.368 176.148 ; 
        RECT 0.832 171.774 0.936 176.148 ; 
        RECT 0.02 171.774 0.36 176.148 ; 
        RECT 62.212 176.094 62.724 180.468 ; 
        RECT 62.156 178.756 62.724 180.046 ; 
        RECT 61.276 177.664 61.812 180.468 ; 
        RECT 61.184 179.004 61.812 180.036 ; 
        RECT 61.276 176.094 61.668 180.468 ; 
        RECT 61.276 176.578 61.724 177.536 ; 
        RECT 61.276 176.094 61.812 176.45 ; 
        RECT 60.376 177.896 60.912 180.468 ; 
        RECT 60.376 176.094 60.768 180.468 ; 
        RECT 58.708 176.094 59.04 180.468 ; 
        RECT 58.708 176.448 59.096 180.19 ; 
        RECT 121.072 176.094 121.412 180.468 ; 
        RECT 120.496 176.094 120.6 180.468 ; 
        RECT 120.064 176.094 120.168 180.468 ; 
        RECT 119.632 176.094 119.736 180.468 ; 
        RECT 119.2 176.094 119.304 180.468 ; 
        RECT 118.768 176.094 118.872 180.468 ; 
        RECT 118.336 176.094 118.44 180.468 ; 
        RECT 117.904 176.094 118.008 180.468 ; 
        RECT 117.472 176.094 117.576 180.468 ; 
        RECT 117.04 176.094 117.144 180.468 ; 
        RECT 116.608 176.094 116.712 180.468 ; 
        RECT 116.176 176.094 116.28 180.468 ; 
        RECT 115.744 176.094 115.848 180.468 ; 
        RECT 115.312 176.094 115.416 180.468 ; 
        RECT 114.88 176.094 114.984 180.468 ; 
        RECT 114.448 176.094 114.552 180.468 ; 
        RECT 114.016 176.094 114.12 180.468 ; 
        RECT 113.584 176.094 113.688 180.468 ; 
        RECT 113.152 176.094 113.256 180.468 ; 
        RECT 112.72 176.094 112.824 180.468 ; 
        RECT 112.288 176.094 112.392 180.468 ; 
        RECT 111.856 176.094 111.96 180.468 ; 
        RECT 111.424 176.094 111.528 180.468 ; 
        RECT 110.992 176.094 111.096 180.468 ; 
        RECT 110.56 176.094 110.664 180.468 ; 
        RECT 110.128 176.094 110.232 180.468 ; 
        RECT 109.696 176.094 109.8 180.468 ; 
        RECT 109.264 176.094 109.368 180.468 ; 
        RECT 108.832 176.094 108.936 180.468 ; 
        RECT 108.4 176.094 108.504 180.468 ; 
        RECT 107.968 176.094 108.072 180.468 ; 
        RECT 107.536 176.094 107.64 180.468 ; 
        RECT 107.104 176.094 107.208 180.468 ; 
        RECT 106.672 176.094 106.776 180.468 ; 
        RECT 106.24 176.094 106.344 180.468 ; 
        RECT 105.808 176.094 105.912 180.468 ; 
        RECT 105.376 176.094 105.48 180.468 ; 
        RECT 104.944 176.094 105.048 180.468 ; 
        RECT 104.512 176.094 104.616 180.468 ; 
        RECT 104.08 176.094 104.184 180.468 ; 
        RECT 103.648 176.094 103.752 180.468 ; 
        RECT 103.216 176.094 103.32 180.468 ; 
        RECT 102.784 176.094 102.888 180.468 ; 
        RECT 102.352 176.094 102.456 180.468 ; 
        RECT 101.92 176.094 102.024 180.468 ; 
        RECT 101.488 176.094 101.592 180.468 ; 
        RECT 101.056 176.094 101.16 180.468 ; 
        RECT 100.624 176.094 100.728 180.468 ; 
        RECT 100.192 176.094 100.296 180.468 ; 
        RECT 99.76 176.094 99.864 180.468 ; 
        RECT 99.328 176.094 99.432 180.468 ; 
        RECT 98.896 176.094 99 180.468 ; 
        RECT 98.464 176.094 98.568 180.468 ; 
        RECT 98.032 176.094 98.136 180.468 ; 
        RECT 97.6 176.094 97.704 180.468 ; 
        RECT 97.168 176.094 97.272 180.468 ; 
        RECT 96.736 176.094 96.84 180.468 ; 
        RECT 96.304 176.094 96.408 180.468 ; 
        RECT 95.872 176.094 95.976 180.468 ; 
        RECT 95.44 176.094 95.544 180.468 ; 
        RECT 95.008 176.094 95.112 180.468 ; 
        RECT 94.576 176.094 94.68 180.468 ; 
        RECT 94.144 176.094 94.248 180.468 ; 
        RECT 93.712 176.094 93.816 180.468 ; 
        RECT 93.28 176.094 93.384 180.468 ; 
        RECT 92.848 176.094 92.952 180.468 ; 
        RECT 92.416 176.094 92.52 180.468 ; 
        RECT 91.984 176.094 92.088 180.468 ; 
        RECT 91.552 176.094 91.656 180.468 ; 
        RECT 91.12 176.094 91.224 180.468 ; 
        RECT 90.688 176.094 90.792 180.468 ; 
        RECT 90.256 176.094 90.36 180.468 ; 
        RECT 89.824 176.094 89.928 180.468 ; 
        RECT 89.392 176.094 89.496 180.468 ; 
        RECT 88.96 176.094 89.064 180.468 ; 
        RECT 88.528 176.094 88.632 180.468 ; 
        RECT 88.096 176.094 88.2 180.468 ; 
        RECT 87.664 176.094 87.768 180.468 ; 
        RECT 87.232 176.094 87.336 180.468 ; 
        RECT 86.8 176.094 86.904 180.468 ; 
        RECT 86.368 176.094 86.472 180.468 ; 
        RECT 85.936 176.094 86.04 180.468 ; 
        RECT 85.504 176.094 85.608 180.468 ; 
        RECT 85.072 176.094 85.176 180.468 ; 
        RECT 84.64 176.094 84.744 180.468 ; 
        RECT 84.208 176.094 84.312 180.468 ; 
        RECT 83.776 176.094 83.88 180.468 ; 
        RECT 83.344 176.094 83.448 180.468 ; 
        RECT 82.912 176.094 83.016 180.468 ; 
        RECT 82.48 176.094 82.584 180.468 ; 
        RECT 82.048 176.094 82.152 180.468 ; 
        RECT 81.616 176.094 81.72 180.468 ; 
        RECT 81.184 176.094 81.288 180.468 ; 
        RECT 80.752 176.094 80.856 180.468 ; 
        RECT 80.32 176.094 80.424 180.468 ; 
        RECT 79.888 176.094 79.992 180.468 ; 
        RECT 79.456 176.094 79.56 180.468 ; 
        RECT 79.024 176.094 79.128 180.468 ; 
        RECT 78.592 176.094 78.696 180.468 ; 
        RECT 78.16 176.094 78.264 180.468 ; 
        RECT 77.728 176.094 77.832 180.468 ; 
        RECT 77.296 176.094 77.4 180.468 ; 
        RECT 76.864 176.094 76.968 180.468 ; 
        RECT 76.432 176.094 76.536 180.468 ; 
        RECT 76 176.094 76.104 180.468 ; 
        RECT 75.568 176.094 75.672 180.468 ; 
        RECT 75.136 176.094 75.24 180.468 ; 
        RECT 74.704 176.094 74.808 180.468 ; 
        RECT 74.272 176.094 74.376 180.468 ; 
        RECT 73.84 176.094 73.944 180.468 ; 
        RECT 73.408 176.094 73.512 180.468 ; 
        RECT 72.976 176.094 73.08 180.468 ; 
        RECT 72.544 176.094 72.648 180.468 ; 
        RECT 72.112 176.094 72.216 180.468 ; 
        RECT 71.68 176.094 71.784 180.468 ; 
        RECT 71.248 176.094 71.352 180.468 ; 
        RECT 70.816 176.094 70.92 180.468 ; 
        RECT 70.384 176.094 70.488 180.468 ; 
        RECT 69.952 176.094 70.056 180.468 ; 
        RECT 69.52 176.094 69.624 180.468 ; 
        RECT 69.088 176.094 69.192 180.468 ; 
        RECT 68.656 176.094 68.76 180.468 ; 
        RECT 68.224 176.094 68.328 180.468 ; 
        RECT 67.792 176.094 67.896 180.468 ; 
        RECT 67.36 176.094 67.464 180.468 ; 
        RECT 66.928 176.094 67.032 180.468 ; 
        RECT 66.496 176.094 66.6 180.468 ; 
        RECT 66.064 176.094 66.168 180.468 ; 
        RECT 65.632 176.094 65.736 180.468 ; 
        RECT 65.2 176.094 65.304 180.468 ; 
        RECT 64.348 176.094 64.656 180.468 ; 
        RECT 56.776 176.094 57.084 180.468 ; 
        RECT 56.128 176.094 56.232 180.468 ; 
        RECT 55.696 176.094 55.8 180.468 ; 
        RECT 55.264 176.094 55.368 180.468 ; 
        RECT 54.832 176.094 54.936 180.468 ; 
        RECT 54.4 176.094 54.504 180.468 ; 
        RECT 53.968 176.094 54.072 180.468 ; 
        RECT 53.536 176.094 53.64 180.468 ; 
        RECT 53.104 176.094 53.208 180.468 ; 
        RECT 52.672 176.094 52.776 180.468 ; 
        RECT 52.24 176.094 52.344 180.468 ; 
        RECT 51.808 176.094 51.912 180.468 ; 
        RECT 51.376 176.094 51.48 180.468 ; 
        RECT 50.944 176.094 51.048 180.468 ; 
        RECT 50.512 176.094 50.616 180.468 ; 
        RECT 50.08 176.094 50.184 180.468 ; 
        RECT 49.648 176.094 49.752 180.468 ; 
        RECT 49.216 176.094 49.32 180.468 ; 
        RECT 48.784 176.094 48.888 180.468 ; 
        RECT 48.352 176.094 48.456 180.468 ; 
        RECT 47.92 176.094 48.024 180.468 ; 
        RECT 47.488 176.094 47.592 180.468 ; 
        RECT 47.056 176.094 47.16 180.468 ; 
        RECT 46.624 176.094 46.728 180.468 ; 
        RECT 46.192 176.094 46.296 180.468 ; 
        RECT 45.76 176.094 45.864 180.468 ; 
        RECT 45.328 176.094 45.432 180.468 ; 
        RECT 44.896 176.094 45 180.468 ; 
        RECT 44.464 176.094 44.568 180.468 ; 
        RECT 44.032 176.094 44.136 180.468 ; 
        RECT 43.6 176.094 43.704 180.468 ; 
        RECT 43.168 176.094 43.272 180.468 ; 
        RECT 42.736 176.094 42.84 180.468 ; 
        RECT 42.304 176.094 42.408 180.468 ; 
        RECT 41.872 176.094 41.976 180.468 ; 
        RECT 41.44 176.094 41.544 180.468 ; 
        RECT 41.008 176.094 41.112 180.468 ; 
        RECT 40.576 176.094 40.68 180.468 ; 
        RECT 40.144 176.094 40.248 180.468 ; 
        RECT 39.712 176.094 39.816 180.468 ; 
        RECT 39.28 176.094 39.384 180.468 ; 
        RECT 38.848 176.094 38.952 180.468 ; 
        RECT 38.416 176.094 38.52 180.468 ; 
        RECT 37.984 176.094 38.088 180.468 ; 
        RECT 37.552 176.094 37.656 180.468 ; 
        RECT 37.12 176.094 37.224 180.468 ; 
        RECT 36.688 176.094 36.792 180.468 ; 
        RECT 36.256 176.094 36.36 180.468 ; 
        RECT 35.824 176.094 35.928 180.468 ; 
        RECT 35.392 176.094 35.496 180.468 ; 
        RECT 34.96 176.094 35.064 180.468 ; 
        RECT 34.528 176.094 34.632 180.468 ; 
        RECT 34.096 176.094 34.2 180.468 ; 
        RECT 33.664 176.094 33.768 180.468 ; 
        RECT 33.232 176.094 33.336 180.468 ; 
        RECT 32.8 176.094 32.904 180.468 ; 
        RECT 32.368 176.094 32.472 180.468 ; 
        RECT 31.936 176.094 32.04 180.468 ; 
        RECT 31.504 176.094 31.608 180.468 ; 
        RECT 31.072 176.094 31.176 180.468 ; 
        RECT 30.64 176.094 30.744 180.468 ; 
        RECT 30.208 176.094 30.312 180.468 ; 
        RECT 29.776 176.094 29.88 180.468 ; 
        RECT 29.344 176.094 29.448 180.468 ; 
        RECT 28.912 176.094 29.016 180.468 ; 
        RECT 28.48 176.094 28.584 180.468 ; 
        RECT 28.048 176.094 28.152 180.468 ; 
        RECT 27.616 176.094 27.72 180.468 ; 
        RECT 27.184 176.094 27.288 180.468 ; 
        RECT 26.752 176.094 26.856 180.468 ; 
        RECT 26.32 176.094 26.424 180.468 ; 
        RECT 25.888 176.094 25.992 180.468 ; 
        RECT 25.456 176.094 25.56 180.468 ; 
        RECT 25.024 176.094 25.128 180.468 ; 
        RECT 24.592 176.094 24.696 180.468 ; 
        RECT 24.16 176.094 24.264 180.468 ; 
        RECT 23.728 176.094 23.832 180.468 ; 
        RECT 23.296 176.094 23.4 180.468 ; 
        RECT 22.864 176.094 22.968 180.468 ; 
        RECT 22.432 176.094 22.536 180.468 ; 
        RECT 22 176.094 22.104 180.468 ; 
        RECT 21.568 176.094 21.672 180.468 ; 
        RECT 21.136 176.094 21.24 180.468 ; 
        RECT 20.704 176.094 20.808 180.468 ; 
        RECT 20.272 176.094 20.376 180.468 ; 
        RECT 19.84 176.094 19.944 180.468 ; 
        RECT 19.408 176.094 19.512 180.468 ; 
        RECT 18.976 176.094 19.08 180.468 ; 
        RECT 18.544 176.094 18.648 180.468 ; 
        RECT 18.112 176.094 18.216 180.468 ; 
        RECT 17.68 176.094 17.784 180.468 ; 
        RECT 17.248 176.094 17.352 180.468 ; 
        RECT 16.816 176.094 16.92 180.468 ; 
        RECT 16.384 176.094 16.488 180.468 ; 
        RECT 15.952 176.094 16.056 180.468 ; 
        RECT 15.52 176.094 15.624 180.468 ; 
        RECT 15.088 176.094 15.192 180.468 ; 
        RECT 14.656 176.094 14.76 180.468 ; 
        RECT 14.224 176.094 14.328 180.468 ; 
        RECT 13.792 176.094 13.896 180.468 ; 
        RECT 13.36 176.094 13.464 180.468 ; 
        RECT 12.928 176.094 13.032 180.468 ; 
        RECT 12.496 176.094 12.6 180.468 ; 
        RECT 12.064 176.094 12.168 180.468 ; 
        RECT 11.632 176.094 11.736 180.468 ; 
        RECT 11.2 176.094 11.304 180.468 ; 
        RECT 10.768 176.094 10.872 180.468 ; 
        RECT 10.336 176.094 10.44 180.468 ; 
        RECT 9.904 176.094 10.008 180.468 ; 
        RECT 9.472 176.094 9.576 180.468 ; 
        RECT 9.04 176.094 9.144 180.468 ; 
        RECT 8.608 176.094 8.712 180.468 ; 
        RECT 8.176 176.094 8.28 180.468 ; 
        RECT 7.744 176.094 7.848 180.468 ; 
        RECT 7.312 176.094 7.416 180.468 ; 
        RECT 6.88 176.094 6.984 180.468 ; 
        RECT 6.448 176.094 6.552 180.468 ; 
        RECT 6.016 176.094 6.12 180.468 ; 
        RECT 5.584 176.094 5.688 180.468 ; 
        RECT 5.152 176.094 5.256 180.468 ; 
        RECT 4.72 176.094 4.824 180.468 ; 
        RECT 4.288 176.094 4.392 180.468 ; 
        RECT 3.856 176.094 3.96 180.468 ; 
        RECT 3.424 176.094 3.528 180.468 ; 
        RECT 2.992 176.094 3.096 180.468 ; 
        RECT 2.56 176.094 2.664 180.468 ; 
        RECT 2.128 176.094 2.232 180.468 ; 
        RECT 1.696 176.094 1.8 180.468 ; 
        RECT 1.264 176.094 1.368 180.468 ; 
        RECT 0.832 176.094 0.936 180.468 ; 
        RECT 0.02 176.094 0.36 180.468 ; 
        RECT 62.212 180.414 62.724 184.788 ; 
        RECT 62.156 183.076 62.724 184.366 ; 
        RECT 61.276 181.984 61.812 184.788 ; 
        RECT 61.184 183.324 61.812 184.356 ; 
        RECT 61.276 180.414 61.668 184.788 ; 
        RECT 61.276 180.898 61.724 181.856 ; 
        RECT 61.276 180.414 61.812 180.77 ; 
        RECT 60.376 182.216 60.912 184.788 ; 
        RECT 60.376 180.414 60.768 184.788 ; 
        RECT 58.708 180.414 59.04 184.788 ; 
        RECT 58.708 180.768 59.096 184.51 ; 
        RECT 121.072 180.414 121.412 184.788 ; 
        RECT 120.496 180.414 120.6 184.788 ; 
        RECT 120.064 180.414 120.168 184.788 ; 
        RECT 119.632 180.414 119.736 184.788 ; 
        RECT 119.2 180.414 119.304 184.788 ; 
        RECT 118.768 180.414 118.872 184.788 ; 
        RECT 118.336 180.414 118.44 184.788 ; 
        RECT 117.904 180.414 118.008 184.788 ; 
        RECT 117.472 180.414 117.576 184.788 ; 
        RECT 117.04 180.414 117.144 184.788 ; 
        RECT 116.608 180.414 116.712 184.788 ; 
        RECT 116.176 180.414 116.28 184.788 ; 
        RECT 115.744 180.414 115.848 184.788 ; 
        RECT 115.312 180.414 115.416 184.788 ; 
        RECT 114.88 180.414 114.984 184.788 ; 
        RECT 114.448 180.414 114.552 184.788 ; 
        RECT 114.016 180.414 114.12 184.788 ; 
        RECT 113.584 180.414 113.688 184.788 ; 
        RECT 113.152 180.414 113.256 184.788 ; 
        RECT 112.72 180.414 112.824 184.788 ; 
        RECT 112.288 180.414 112.392 184.788 ; 
        RECT 111.856 180.414 111.96 184.788 ; 
        RECT 111.424 180.414 111.528 184.788 ; 
        RECT 110.992 180.414 111.096 184.788 ; 
        RECT 110.56 180.414 110.664 184.788 ; 
        RECT 110.128 180.414 110.232 184.788 ; 
        RECT 109.696 180.414 109.8 184.788 ; 
        RECT 109.264 180.414 109.368 184.788 ; 
        RECT 108.832 180.414 108.936 184.788 ; 
        RECT 108.4 180.414 108.504 184.788 ; 
        RECT 107.968 180.414 108.072 184.788 ; 
        RECT 107.536 180.414 107.64 184.788 ; 
        RECT 107.104 180.414 107.208 184.788 ; 
        RECT 106.672 180.414 106.776 184.788 ; 
        RECT 106.24 180.414 106.344 184.788 ; 
        RECT 105.808 180.414 105.912 184.788 ; 
        RECT 105.376 180.414 105.48 184.788 ; 
        RECT 104.944 180.414 105.048 184.788 ; 
        RECT 104.512 180.414 104.616 184.788 ; 
        RECT 104.08 180.414 104.184 184.788 ; 
        RECT 103.648 180.414 103.752 184.788 ; 
        RECT 103.216 180.414 103.32 184.788 ; 
        RECT 102.784 180.414 102.888 184.788 ; 
        RECT 102.352 180.414 102.456 184.788 ; 
        RECT 101.92 180.414 102.024 184.788 ; 
        RECT 101.488 180.414 101.592 184.788 ; 
        RECT 101.056 180.414 101.16 184.788 ; 
        RECT 100.624 180.414 100.728 184.788 ; 
        RECT 100.192 180.414 100.296 184.788 ; 
        RECT 99.76 180.414 99.864 184.788 ; 
        RECT 99.328 180.414 99.432 184.788 ; 
        RECT 98.896 180.414 99 184.788 ; 
        RECT 98.464 180.414 98.568 184.788 ; 
        RECT 98.032 180.414 98.136 184.788 ; 
        RECT 97.6 180.414 97.704 184.788 ; 
        RECT 97.168 180.414 97.272 184.788 ; 
        RECT 96.736 180.414 96.84 184.788 ; 
        RECT 96.304 180.414 96.408 184.788 ; 
        RECT 95.872 180.414 95.976 184.788 ; 
        RECT 95.44 180.414 95.544 184.788 ; 
        RECT 95.008 180.414 95.112 184.788 ; 
        RECT 94.576 180.414 94.68 184.788 ; 
        RECT 94.144 180.414 94.248 184.788 ; 
        RECT 93.712 180.414 93.816 184.788 ; 
        RECT 93.28 180.414 93.384 184.788 ; 
        RECT 92.848 180.414 92.952 184.788 ; 
        RECT 92.416 180.414 92.52 184.788 ; 
        RECT 91.984 180.414 92.088 184.788 ; 
        RECT 91.552 180.414 91.656 184.788 ; 
        RECT 91.12 180.414 91.224 184.788 ; 
        RECT 90.688 180.414 90.792 184.788 ; 
        RECT 90.256 180.414 90.36 184.788 ; 
        RECT 89.824 180.414 89.928 184.788 ; 
        RECT 89.392 180.414 89.496 184.788 ; 
        RECT 88.96 180.414 89.064 184.788 ; 
        RECT 88.528 180.414 88.632 184.788 ; 
        RECT 88.096 180.414 88.2 184.788 ; 
        RECT 87.664 180.414 87.768 184.788 ; 
        RECT 87.232 180.414 87.336 184.788 ; 
        RECT 86.8 180.414 86.904 184.788 ; 
        RECT 86.368 180.414 86.472 184.788 ; 
        RECT 85.936 180.414 86.04 184.788 ; 
        RECT 85.504 180.414 85.608 184.788 ; 
        RECT 85.072 180.414 85.176 184.788 ; 
        RECT 84.64 180.414 84.744 184.788 ; 
        RECT 84.208 180.414 84.312 184.788 ; 
        RECT 83.776 180.414 83.88 184.788 ; 
        RECT 83.344 180.414 83.448 184.788 ; 
        RECT 82.912 180.414 83.016 184.788 ; 
        RECT 82.48 180.414 82.584 184.788 ; 
        RECT 82.048 180.414 82.152 184.788 ; 
        RECT 81.616 180.414 81.72 184.788 ; 
        RECT 81.184 180.414 81.288 184.788 ; 
        RECT 80.752 180.414 80.856 184.788 ; 
        RECT 80.32 180.414 80.424 184.788 ; 
        RECT 79.888 180.414 79.992 184.788 ; 
        RECT 79.456 180.414 79.56 184.788 ; 
        RECT 79.024 180.414 79.128 184.788 ; 
        RECT 78.592 180.414 78.696 184.788 ; 
        RECT 78.16 180.414 78.264 184.788 ; 
        RECT 77.728 180.414 77.832 184.788 ; 
        RECT 77.296 180.414 77.4 184.788 ; 
        RECT 76.864 180.414 76.968 184.788 ; 
        RECT 76.432 180.414 76.536 184.788 ; 
        RECT 76 180.414 76.104 184.788 ; 
        RECT 75.568 180.414 75.672 184.788 ; 
        RECT 75.136 180.414 75.24 184.788 ; 
        RECT 74.704 180.414 74.808 184.788 ; 
        RECT 74.272 180.414 74.376 184.788 ; 
        RECT 73.84 180.414 73.944 184.788 ; 
        RECT 73.408 180.414 73.512 184.788 ; 
        RECT 72.976 180.414 73.08 184.788 ; 
        RECT 72.544 180.414 72.648 184.788 ; 
        RECT 72.112 180.414 72.216 184.788 ; 
        RECT 71.68 180.414 71.784 184.788 ; 
        RECT 71.248 180.414 71.352 184.788 ; 
        RECT 70.816 180.414 70.92 184.788 ; 
        RECT 70.384 180.414 70.488 184.788 ; 
        RECT 69.952 180.414 70.056 184.788 ; 
        RECT 69.52 180.414 69.624 184.788 ; 
        RECT 69.088 180.414 69.192 184.788 ; 
        RECT 68.656 180.414 68.76 184.788 ; 
        RECT 68.224 180.414 68.328 184.788 ; 
        RECT 67.792 180.414 67.896 184.788 ; 
        RECT 67.36 180.414 67.464 184.788 ; 
        RECT 66.928 180.414 67.032 184.788 ; 
        RECT 66.496 180.414 66.6 184.788 ; 
        RECT 66.064 180.414 66.168 184.788 ; 
        RECT 65.632 180.414 65.736 184.788 ; 
        RECT 65.2 180.414 65.304 184.788 ; 
        RECT 64.348 180.414 64.656 184.788 ; 
        RECT 56.776 180.414 57.084 184.788 ; 
        RECT 56.128 180.414 56.232 184.788 ; 
        RECT 55.696 180.414 55.8 184.788 ; 
        RECT 55.264 180.414 55.368 184.788 ; 
        RECT 54.832 180.414 54.936 184.788 ; 
        RECT 54.4 180.414 54.504 184.788 ; 
        RECT 53.968 180.414 54.072 184.788 ; 
        RECT 53.536 180.414 53.64 184.788 ; 
        RECT 53.104 180.414 53.208 184.788 ; 
        RECT 52.672 180.414 52.776 184.788 ; 
        RECT 52.24 180.414 52.344 184.788 ; 
        RECT 51.808 180.414 51.912 184.788 ; 
        RECT 51.376 180.414 51.48 184.788 ; 
        RECT 50.944 180.414 51.048 184.788 ; 
        RECT 50.512 180.414 50.616 184.788 ; 
        RECT 50.08 180.414 50.184 184.788 ; 
        RECT 49.648 180.414 49.752 184.788 ; 
        RECT 49.216 180.414 49.32 184.788 ; 
        RECT 48.784 180.414 48.888 184.788 ; 
        RECT 48.352 180.414 48.456 184.788 ; 
        RECT 47.92 180.414 48.024 184.788 ; 
        RECT 47.488 180.414 47.592 184.788 ; 
        RECT 47.056 180.414 47.16 184.788 ; 
        RECT 46.624 180.414 46.728 184.788 ; 
        RECT 46.192 180.414 46.296 184.788 ; 
        RECT 45.76 180.414 45.864 184.788 ; 
        RECT 45.328 180.414 45.432 184.788 ; 
        RECT 44.896 180.414 45 184.788 ; 
        RECT 44.464 180.414 44.568 184.788 ; 
        RECT 44.032 180.414 44.136 184.788 ; 
        RECT 43.6 180.414 43.704 184.788 ; 
        RECT 43.168 180.414 43.272 184.788 ; 
        RECT 42.736 180.414 42.84 184.788 ; 
        RECT 42.304 180.414 42.408 184.788 ; 
        RECT 41.872 180.414 41.976 184.788 ; 
        RECT 41.44 180.414 41.544 184.788 ; 
        RECT 41.008 180.414 41.112 184.788 ; 
        RECT 40.576 180.414 40.68 184.788 ; 
        RECT 40.144 180.414 40.248 184.788 ; 
        RECT 39.712 180.414 39.816 184.788 ; 
        RECT 39.28 180.414 39.384 184.788 ; 
        RECT 38.848 180.414 38.952 184.788 ; 
        RECT 38.416 180.414 38.52 184.788 ; 
        RECT 37.984 180.414 38.088 184.788 ; 
        RECT 37.552 180.414 37.656 184.788 ; 
        RECT 37.12 180.414 37.224 184.788 ; 
        RECT 36.688 180.414 36.792 184.788 ; 
        RECT 36.256 180.414 36.36 184.788 ; 
        RECT 35.824 180.414 35.928 184.788 ; 
        RECT 35.392 180.414 35.496 184.788 ; 
        RECT 34.96 180.414 35.064 184.788 ; 
        RECT 34.528 180.414 34.632 184.788 ; 
        RECT 34.096 180.414 34.2 184.788 ; 
        RECT 33.664 180.414 33.768 184.788 ; 
        RECT 33.232 180.414 33.336 184.788 ; 
        RECT 32.8 180.414 32.904 184.788 ; 
        RECT 32.368 180.414 32.472 184.788 ; 
        RECT 31.936 180.414 32.04 184.788 ; 
        RECT 31.504 180.414 31.608 184.788 ; 
        RECT 31.072 180.414 31.176 184.788 ; 
        RECT 30.64 180.414 30.744 184.788 ; 
        RECT 30.208 180.414 30.312 184.788 ; 
        RECT 29.776 180.414 29.88 184.788 ; 
        RECT 29.344 180.414 29.448 184.788 ; 
        RECT 28.912 180.414 29.016 184.788 ; 
        RECT 28.48 180.414 28.584 184.788 ; 
        RECT 28.048 180.414 28.152 184.788 ; 
        RECT 27.616 180.414 27.72 184.788 ; 
        RECT 27.184 180.414 27.288 184.788 ; 
        RECT 26.752 180.414 26.856 184.788 ; 
        RECT 26.32 180.414 26.424 184.788 ; 
        RECT 25.888 180.414 25.992 184.788 ; 
        RECT 25.456 180.414 25.56 184.788 ; 
        RECT 25.024 180.414 25.128 184.788 ; 
        RECT 24.592 180.414 24.696 184.788 ; 
        RECT 24.16 180.414 24.264 184.788 ; 
        RECT 23.728 180.414 23.832 184.788 ; 
        RECT 23.296 180.414 23.4 184.788 ; 
        RECT 22.864 180.414 22.968 184.788 ; 
        RECT 22.432 180.414 22.536 184.788 ; 
        RECT 22 180.414 22.104 184.788 ; 
        RECT 21.568 180.414 21.672 184.788 ; 
        RECT 21.136 180.414 21.24 184.788 ; 
        RECT 20.704 180.414 20.808 184.788 ; 
        RECT 20.272 180.414 20.376 184.788 ; 
        RECT 19.84 180.414 19.944 184.788 ; 
        RECT 19.408 180.414 19.512 184.788 ; 
        RECT 18.976 180.414 19.08 184.788 ; 
        RECT 18.544 180.414 18.648 184.788 ; 
        RECT 18.112 180.414 18.216 184.788 ; 
        RECT 17.68 180.414 17.784 184.788 ; 
        RECT 17.248 180.414 17.352 184.788 ; 
        RECT 16.816 180.414 16.92 184.788 ; 
        RECT 16.384 180.414 16.488 184.788 ; 
        RECT 15.952 180.414 16.056 184.788 ; 
        RECT 15.52 180.414 15.624 184.788 ; 
        RECT 15.088 180.414 15.192 184.788 ; 
        RECT 14.656 180.414 14.76 184.788 ; 
        RECT 14.224 180.414 14.328 184.788 ; 
        RECT 13.792 180.414 13.896 184.788 ; 
        RECT 13.36 180.414 13.464 184.788 ; 
        RECT 12.928 180.414 13.032 184.788 ; 
        RECT 12.496 180.414 12.6 184.788 ; 
        RECT 12.064 180.414 12.168 184.788 ; 
        RECT 11.632 180.414 11.736 184.788 ; 
        RECT 11.2 180.414 11.304 184.788 ; 
        RECT 10.768 180.414 10.872 184.788 ; 
        RECT 10.336 180.414 10.44 184.788 ; 
        RECT 9.904 180.414 10.008 184.788 ; 
        RECT 9.472 180.414 9.576 184.788 ; 
        RECT 9.04 180.414 9.144 184.788 ; 
        RECT 8.608 180.414 8.712 184.788 ; 
        RECT 8.176 180.414 8.28 184.788 ; 
        RECT 7.744 180.414 7.848 184.788 ; 
        RECT 7.312 180.414 7.416 184.788 ; 
        RECT 6.88 180.414 6.984 184.788 ; 
        RECT 6.448 180.414 6.552 184.788 ; 
        RECT 6.016 180.414 6.12 184.788 ; 
        RECT 5.584 180.414 5.688 184.788 ; 
        RECT 5.152 180.414 5.256 184.788 ; 
        RECT 4.72 180.414 4.824 184.788 ; 
        RECT 4.288 180.414 4.392 184.788 ; 
        RECT 3.856 180.414 3.96 184.788 ; 
        RECT 3.424 180.414 3.528 184.788 ; 
        RECT 2.992 180.414 3.096 184.788 ; 
        RECT 2.56 180.414 2.664 184.788 ; 
        RECT 2.128 180.414 2.232 184.788 ; 
        RECT 1.696 180.414 1.8 184.788 ; 
        RECT 1.264 180.414 1.368 184.788 ; 
        RECT 0.832 180.414 0.936 184.788 ; 
        RECT 0.02 180.414 0.36 184.788 ; 
        RECT 62.212 184.734 62.724 189.108 ; 
        RECT 62.156 187.396 62.724 188.686 ; 
        RECT 61.276 186.304 61.812 189.108 ; 
        RECT 61.184 187.644 61.812 188.676 ; 
        RECT 61.276 184.734 61.668 189.108 ; 
        RECT 61.276 185.218 61.724 186.176 ; 
        RECT 61.276 184.734 61.812 185.09 ; 
        RECT 60.376 186.536 60.912 189.108 ; 
        RECT 60.376 184.734 60.768 189.108 ; 
        RECT 58.708 184.734 59.04 189.108 ; 
        RECT 58.708 185.088 59.096 188.83 ; 
        RECT 121.072 184.734 121.412 189.108 ; 
        RECT 120.496 184.734 120.6 189.108 ; 
        RECT 120.064 184.734 120.168 189.108 ; 
        RECT 119.632 184.734 119.736 189.108 ; 
        RECT 119.2 184.734 119.304 189.108 ; 
        RECT 118.768 184.734 118.872 189.108 ; 
        RECT 118.336 184.734 118.44 189.108 ; 
        RECT 117.904 184.734 118.008 189.108 ; 
        RECT 117.472 184.734 117.576 189.108 ; 
        RECT 117.04 184.734 117.144 189.108 ; 
        RECT 116.608 184.734 116.712 189.108 ; 
        RECT 116.176 184.734 116.28 189.108 ; 
        RECT 115.744 184.734 115.848 189.108 ; 
        RECT 115.312 184.734 115.416 189.108 ; 
        RECT 114.88 184.734 114.984 189.108 ; 
        RECT 114.448 184.734 114.552 189.108 ; 
        RECT 114.016 184.734 114.12 189.108 ; 
        RECT 113.584 184.734 113.688 189.108 ; 
        RECT 113.152 184.734 113.256 189.108 ; 
        RECT 112.72 184.734 112.824 189.108 ; 
        RECT 112.288 184.734 112.392 189.108 ; 
        RECT 111.856 184.734 111.96 189.108 ; 
        RECT 111.424 184.734 111.528 189.108 ; 
        RECT 110.992 184.734 111.096 189.108 ; 
        RECT 110.56 184.734 110.664 189.108 ; 
        RECT 110.128 184.734 110.232 189.108 ; 
        RECT 109.696 184.734 109.8 189.108 ; 
        RECT 109.264 184.734 109.368 189.108 ; 
        RECT 108.832 184.734 108.936 189.108 ; 
        RECT 108.4 184.734 108.504 189.108 ; 
        RECT 107.968 184.734 108.072 189.108 ; 
        RECT 107.536 184.734 107.64 189.108 ; 
        RECT 107.104 184.734 107.208 189.108 ; 
        RECT 106.672 184.734 106.776 189.108 ; 
        RECT 106.24 184.734 106.344 189.108 ; 
        RECT 105.808 184.734 105.912 189.108 ; 
        RECT 105.376 184.734 105.48 189.108 ; 
        RECT 104.944 184.734 105.048 189.108 ; 
        RECT 104.512 184.734 104.616 189.108 ; 
        RECT 104.08 184.734 104.184 189.108 ; 
        RECT 103.648 184.734 103.752 189.108 ; 
        RECT 103.216 184.734 103.32 189.108 ; 
        RECT 102.784 184.734 102.888 189.108 ; 
        RECT 102.352 184.734 102.456 189.108 ; 
        RECT 101.92 184.734 102.024 189.108 ; 
        RECT 101.488 184.734 101.592 189.108 ; 
        RECT 101.056 184.734 101.16 189.108 ; 
        RECT 100.624 184.734 100.728 189.108 ; 
        RECT 100.192 184.734 100.296 189.108 ; 
        RECT 99.76 184.734 99.864 189.108 ; 
        RECT 99.328 184.734 99.432 189.108 ; 
        RECT 98.896 184.734 99 189.108 ; 
        RECT 98.464 184.734 98.568 189.108 ; 
        RECT 98.032 184.734 98.136 189.108 ; 
        RECT 97.6 184.734 97.704 189.108 ; 
        RECT 97.168 184.734 97.272 189.108 ; 
        RECT 96.736 184.734 96.84 189.108 ; 
        RECT 96.304 184.734 96.408 189.108 ; 
        RECT 95.872 184.734 95.976 189.108 ; 
        RECT 95.44 184.734 95.544 189.108 ; 
        RECT 95.008 184.734 95.112 189.108 ; 
        RECT 94.576 184.734 94.68 189.108 ; 
        RECT 94.144 184.734 94.248 189.108 ; 
        RECT 93.712 184.734 93.816 189.108 ; 
        RECT 93.28 184.734 93.384 189.108 ; 
        RECT 92.848 184.734 92.952 189.108 ; 
        RECT 92.416 184.734 92.52 189.108 ; 
        RECT 91.984 184.734 92.088 189.108 ; 
        RECT 91.552 184.734 91.656 189.108 ; 
        RECT 91.12 184.734 91.224 189.108 ; 
        RECT 90.688 184.734 90.792 189.108 ; 
        RECT 90.256 184.734 90.36 189.108 ; 
        RECT 89.824 184.734 89.928 189.108 ; 
        RECT 89.392 184.734 89.496 189.108 ; 
        RECT 88.96 184.734 89.064 189.108 ; 
        RECT 88.528 184.734 88.632 189.108 ; 
        RECT 88.096 184.734 88.2 189.108 ; 
        RECT 87.664 184.734 87.768 189.108 ; 
        RECT 87.232 184.734 87.336 189.108 ; 
        RECT 86.8 184.734 86.904 189.108 ; 
        RECT 86.368 184.734 86.472 189.108 ; 
        RECT 85.936 184.734 86.04 189.108 ; 
        RECT 85.504 184.734 85.608 189.108 ; 
        RECT 85.072 184.734 85.176 189.108 ; 
        RECT 84.64 184.734 84.744 189.108 ; 
        RECT 84.208 184.734 84.312 189.108 ; 
        RECT 83.776 184.734 83.88 189.108 ; 
        RECT 83.344 184.734 83.448 189.108 ; 
        RECT 82.912 184.734 83.016 189.108 ; 
        RECT 82.48 184.734 82.584 189.108 ; 
        RECT 82.048 184.734 82.152 189.108 ; 
        RECT 81.616 184.734 81.72 189.108 ; 
        RECT 81.184 184.734 81.288 189.108 ; 
        RECT 80.752 184.734 80.856 189.108 ; 
        RECT 80.32 184.734 80.424 189.108 ; 
        RECT 79.888 184.734 79.992 189.108 ; 
        RECT 79.456 184.734 79.56 189.108 ; 
        RECT 79.024 184.734 79.128 189.108 ; 
        RECT 78.592 184.734 78.696 189.108 ; 
        RECT 78.16 184.734 78.264 189.108 ; 
        RECT 77.728 184.734 77.832 189.108 ; 
        RECT 77.296 184.734 77.4 189.108 ; 
        RECT 76.864 184.734 76.968 189.108 ; 
        RECT 76.432 184.734 76.536 189.108 ; 
        RECT 76 184.734 76.104 189.108 ; 
        RECT 75.568 184.734 75.672 189.108 ; 
        RECT 75.136 184.734 75.24 189.108 ; 
        RECT 74.704 184.734 74.808 189.108 ; 
        RECT 74.272 184.734 74.376 189.108 ; 
        RECT 73.84 184.734 73.944 189.108 ; 
        RECT 73.408 184.734 73.512 189.108 ; 
        RECT 72.976 184.734 73.08 189.108 ; 
        RECT 72.544 184.734 72.648 189.108 ; 
        RECT 72.112 184.734 72.216 189.108 ; 
        RECT 71.68 184.734 71.784 189.108 ; 
        RECT 71.248 184.734 71.352 189.108 ; 
        RECT 70.816 184.734 70.92 189.108 ; 
        RECT 70.384 184.734 70.488 189.108 ; 
        RECT 69.952 184.734 70.056 189.108 ; 
        RECT 69.52 184.734 69.624 189.108 ; 
        RECT 69.088 184.734 69.192 189.108 ; 
        RECT 68.656 184.734 68.76 189.108 ; 
        RECT 68.224 184.734 68.328 189.108 ; 
        RECT 67.792 184.734 67.896 189.108 ; 
        RECT 67.36 184.734 67.464 189.108 ; 
        RECT 66.928 184.734 67.032 189.108 ; 
        RECT 66.496 184.734 66.6 189.108 ; 
        RECT 66.064 184.734 66.168 189.108 ; 
        RECT 65.632 184.734 65.736 189.108 ; 
        RECT 65.2 184.734 65.304 189.108 ; 
        RECT 64.348 184.734 64.656 189.108 ; 
        RECT 56.776 184.734 57.084 189.108 ; 
        RECT 56.128 184.734 56.232 189.108 ; 
        RECT 55.696 184.734 55.8 189.108 ; 
        RECT 55.264 184.734 55.368 189.108 ; 
        RECT 54.832 184.734 54.936 189.108 ; 
        RECT 54.4 184.734 54.504 189.108 ; 
        RECT 53.968 184.734 54.072 189.108 ; 
        RECT 53.536 184.734 53.64 189.108 ; 
        RECT 53.104 184.734 53.208 189.108 ; 
        RECT 52.672 184.734 52.776 189.108 ; 
        RECT 52.24 184.734 52.344 189.108 ; 
        RECT 51.808 184.734 51.912 189.108 ; 
        RECT 51.376 184.734 51.48 189.108 ; 
        RECT 50.944 184.734 51.048 189.108 ; 
        RECT 50.512 184.734 50.616 189.108 ; 
        RECT 50.08 184.734 50.184 189.108 ; 
        RECT 49.648 184.734 49.752 189.108 ; 
        RECT 49.216 184.734 49.32 189.108 ; 
        RECT 48.784 184.734 48.888 189.108 ; 
        RECT 48.352 184.734 48.456 189.108 ; 
        RECT 47.92 184.734 48.024 189.108 ; 
        RECT 47.488 184.734 47.592 189.108 ; 
        RECT 47.056 184.734 47.16 189.108 ; 
        RECT 46.624 184.734 46.728 189.108 ; 
        RECT 46.192 184.734 46.296 189.108 ; 
        RECT 45.76 184.734 45.864 189.108 ; 
        RECT 45.328 184.734 45.432 189.108 ; 
        RECT 44.896 184.734 45 189.108 ; 
        RECT 44.464 184.734 44.568 189.108 ; 
        RECT 44.032 184.734 44.136 189.108 ; 
        RECT 43.6 184.734 43.704 189.108 ; 
        RECT 43.168 184.734 43.272 189.108 ; 
        RECT 42.736 184.734 42.84 189.108 ; 
        RECT 42.304 184.734 42.408 189.108 ; 
        RECT 41.872 184.734 41.976 189.108 ; 
        RECT 41.44 184.734 41.544 189.108 ; 
        RECT 41.008 184.734 41.112 189.108 ; 
        RECT 40.576 184.734 40.68 189.108 ; 
        RECT 40.144 184.734 40.248 189.108 ; 
        RECT 39.712 184.734 39.816 189.108 ; 
        RECT 39.28 184.734 39.384 189.108 ; 
        RECT 38.848 184.734 38.952 189.108 ; 
        RECT 38.416 184.734 38.52 189.108 ; 
        RECT 37.984 184.734 38.088 189.108 ; 
        RECT 37.552 184.734 37.656 189.108 ; 
        RECT 37.12 184.734 37.224 189.108 ; 
        RECT 36.688 184.734 36.792 189.108 ; 
        RECT 36.256 184.734 36.36 189.108 ; 
        RECT 35.824 184.734 35.928 189.108 ; 
        RECT 35.392 184.734 35.496 189.108 ; 
        RECT 34.96 184.734 35.064 189.108 ; 
        RECT 34.528 184.734 34.632 189.108 ; 
        RECT 34.096 184.734 34.2 189.108 ; 
        RECT 33.664 184.734 33.768 189.108 ; 
        RECT 33.232 184.734 33.336 189.108 ; 
        RECT 32.8 184.734 32.904 189.108 ; 
        RECT 32.368 184.734 32.472 189.108 ; 
        RECT 31.936 184.734 32.04 189.108 ; 
        RECT 31.504 184.734 31.608 189.108 ; 
        RECT 31.072 184.734 31.176 189.108 ; 
        RECT 30.64 184.734 30.744 189.108 ; 
        RECT 30.208 184.734 30.312 189.108 ; 
        RECT 29.776 184.734 29.88 189.108 ; 
        RECT 29.344 184.734 29.448 189.108 ; 
        RECT 28.912 184.734 29.016 189.108 ; 
        RECT 28.48 184.734 28.584 189.108 ; 
        RECT 28.048 184.734 28.152 189.108 ; 
        RECT 27.616 184.734 27.72 189.108 ; 
        RECT 27.184 184.734 27.288 189.108 ; 
        RECT 26.752 184.734 26.856 189.108 ; 
        RECT 26.32 184.734 26.424 189.108 ; 
        RECT 25.888 184.734 25.992 189.108 ; 
        RECT 25.456 184.734 25.56 189.108 ; 
        RECT 25.024 184.734 25.128 189.108 ; 
        RECT 24.592 184.734 24.696 189.108 ; 
        RECT 24.16 184.734 24.264 189.108 ; 
        RECT 23.728 184.734 23.832 189.108 ; 
        RECT 23.296 184.734 23.4 189.108 ; 
        RECT 22.864 184.734 22.968 189.108 ; 
        RECT 22.432 184.734 22.536 189.108 ; 
        RECT 22 184.734 22.104 189.108 ; 
        RECT 21.568 184.734 21.672 189.108 ; 
        RECT 21.136 184.734 21.24 189.108 ; 
        RECT 20.704 184.734 20.808 189.108 ; 
        RECT 20.272 184.734 20.376 189.108 ; 
        RECT 19.84 184.734 19.944 189.108 ; 
        RECT 19.408 184.734 19.512 189.108 ; 
        RECT 18.976 184.734 19.08 189.108 ; 
        RECT 18.544 184.734 18.648 189.108 ; 
        RECT 18.112 184.734 18.216 189.108 ; 
        RECT 17.68 184.734 17.784 189.108 ; 
        RECT 17.248 184.734 17.352 189.108 ; 
        RECT 16.816 184.734 16.92 189.108 ; 
        RECT 16.384 184.734 16.488 189.108 ; 
        RECT 15.952 184.734 16.056 189.108 ; 
        RECT 15.52 184.734 15.624 189.108 ; 
        RECT 15.088 184.734 15.192 189.108 ; 
        RECT 14.656 184.734 14.76 189.108 ; 
        RECT 14.224 184.734 14.328 189.108 ; 
        RECT 13.792 184.734 13.896 189.108 ; 
        RECT 13.36 184.734 13.464 189.108 ; 
        RECT 12.928 184.734 13.032 189.108 ; 
        RECT 12.496 184.734 12.6 189.108 ; 
        RECT 12.064 184.734 12.168 189.108 ; 
        RECT 11.632 184.734 11.736 189.108 ; 
        RECT 11.2 184.734 11.304 189.108 ; 
        RECT 10.768 184.734 10.872 189.108 ; 
        RECT 10.336 184.734 10.44 189.108 ; 
        RECT 9.904 184.734 10.008 189.108 ; 
        RECT 9.472 184.734 9.576 189.108 ; 
        RECT 9.04 184.734 9.144 189.108 ; 
        RECT 8.608 184.734 8.712 189.108 ; 
        RECT 8.176 184.734 8.28 189.108 ; 
        RECT 7.744 184.734 7.848 189.108 ; 
        RECT 7.312 184.734 7.416 189.108 ; 
        RECT 6.88 184.734 6.984 189.108 ; 
        RECT 6.448 184.734 6.552 189.108 ; 
        RECT 6.016 184.734 6.12 189.108 ; 
        RECT 5.584 184.734 5.688 189.108 ; 
        RECT 5.152 184.734 5.256 189.108 ; 
        RECT 4.72 184.734 4.824 189.108 ; 
        RECT 4.288 184.734 4.392 189.108 ; 
        RECT 3.856 184.734 3.96 189.108 ; 
        RECT 3.424 184.734 3.528 189.108 ; 
        RECT 2.992 184.734 3.096 189.108 ; 
        RECT 2.56 184.734 2.664 189.108 ; 
        RECT 2.128 184.734 2.232 189.108 ; 
        RECT 1.696 184.734 1.8 189.108 ; 
        RECT 1.264 184.734 1.368 189.108 ; 
        RECT 0.832 184.734 0.936 189.108 ; 
        RECT 0.02 184.734 0.36 189.108 ; 
        RECT 62.212 189.054 62.724 193.428 ; 
        RECT 62.156 191.716 62.724 193.006 ; 
        RECT 61.276 190.624 61.812 193.428 ; 
        RECT 61.184 191.964 61.812 192.996 ; 
        RECT 61.276 189.054 61.668 193.428 ; 
        RECT 61.276 189.538 61.724 190.496 ; 
        RECT 61.276 189.054 61.812 189.41 ; 
        RECT 60.376 190.856 60.912 193.428 ; 
        RECT 60.376 189.054 60.768 193.428 ; 
        RECT 58.708 189.054 59.04 193.428 ; 
        RECT 58.708 189.408 59.096 193.15 ; 
        RECT 121.072 189.054 121.412 193.428 ; 
        RECT 120.496 189.054 120.6 193.428 ; 
        RECT 120.064 189.054 120.168 193.428 ; 
        RECT 119.632 189.054 119.736 193.428 ; 
        RECT 119.2 189.054 119.304 193.428 ; 
        RECT 118.768 189.054 118.872 193.428 ; 
        RECT 118.336 189.054 118.44 193.428 ; 
        RECT 117.904 189.054 118.008 193.428 ; 
        RECT 117.472 189.054 117.576 193.428 ; 
        RECT 117.04 189.054 117.144 193.428 ; 
        RECT 116.608 189.054 116.712 193.428 ; 
        RECT 116.176 189.054 116.28 193.428 ; 
        RECT 115.744 189.054 115.848 193.428 ; 
        RECT 115.312 189.054 115.416 193.428 ; 
        RECT 114.88 189.054 114.984 193.428 ; 
        RECT 114.448 189.054 114.552 193.428 ; 
        RECT 114.016 189.054 114.12 193.428 ; 
        RECT 113.584 189.054 113.688 193.428 ; 
        RECT 113.152 189.054 113.256 193.428 ; 
        RECT 112.72 189.054 112.824 193.428 ; 
        RECT 112.288 189.054 112.392 193.428 ; 
        RECT 111.856 189.054 111.96 193.428 ; 
        RECT 111.424 189.054 111.528 193.428 ; 
        RECT 110.992 189.054 111.096 193.428 ; 
        RECT 110.56 189.054 110.664 193.428 ; 
        RECT 110.128 189.054 110.232 193.428 ; 
        RECT 109.696 189.054 109.8 193.428 ; 
        RECT 109.264 189.054 109.368 193.428 ; 
        RECT 108.832 189.054 108.936 193.428 ; 
        RECT 108.4 189.054 108.504 193.428 ; 
        RECT 107.968 189.054 108.072 193.428 ; 
        RECT 107.536 189.054 107.64 193.428 ; 
        RECT 107.104 189.054 107.208 193.428 ; 
        RECT 106.672 189.054 106.776 193.428 ; 
        RECT 106.24 189.054 106.344 193.428 ; 
        RECT 105.808 189.054 105.912 193.428 ; 
        RECT 105.376 189.054 105.48 193.428 ; 
        RECT 104.944 189.054 105.048 193.428 ; 
        RECT 104.512 189.054 104.616 193.428 ; 
        RECT 104.08 189.054 104.184 193.428 ; 
        RECT 103.648 189.054 103.752 193.428 ; 
        RECT 103.216 189.054 103.32 193.428 ; 
        RECT 102.784 189.054 102.888 193.428 ; 
        RECT 102.352 189.054 102.456 193.428 ; 
        RECT 101.92 189.054 102.024 193.428 ; 
        RECT 101.488 189.054 101.592 193.428 ; 
        RECT 101.056 189.054 101.16 193.428 ; 
        RECT 100.624 189.054 100.728 193.428 ; 
        RECT 100.192 189.054 100.296 193.428 ; 
        RECT 99.76 189.054 99.864 193.428 ; 
        RECT 99.328 189.054 99.432 193.428 ; 
        RECT 98.896 189.054 99 193.428 ; 
        RECT 98.464 189.054 98.568 193.428 ; 
        RECT 98.032 189.054 98.136 193.428 ; 
        RECT 97.6 189.054 97.704 193.428 ; 
        RECT 97.168 189.054 97.272 193.428 ; 
        RECT 96.736 189.054 96.84 193.428 ; 
        RECT 96.304 189.054 96.408 193.428 ; 
        RECT 95.872 189.054 95.976 193.428 ; 
        RECT 95.44 189.054 95.544 193.428 ; 
        RECT 95.008 189.054 95.112 193.428 ; 
        RECT 94.576 189.054 94.68 193.428 ; 
        RECT 94.144 189.054 94.248 193.428 ; 
        RECT 93.712 189.054 93.816 193.428 ; 
        RECT 93.28 189.054 93.384 193.428 ; 
        RECT 92.848 189.054 92.952 193.428 ; 
        RECT 92.416 189.054 92.52 193.428 ; 
        RECT 91.984 189.054 92.088 193.428 ; 
        RECT 91.552 189.054 91.656 193.428 ; 
        RECT 91.12 189.054 91.224 193.428 ; 
        RECT 90.688 189.054 90.792 193.428 ; 
        RECT 90.256 189.054 90.36 193.428 ; 
        RECT 89.824 189.054 89.928 193.428 ; 
        RECT 89.392 189.054 89.496 193.428 ; 
        RECT 88.96 189.054 89.064 193.428 ; 
        RECT 88.528 189.054 88.632 193.428 ; 
        RECT 88.096 189.054 88.2 193.428 ; 
        RECT 87.664 189.054 87.768 193.428 ; 
        RECT 87.232 189.054 87.336 193.428 ; 
        RECT 86.8 189.054 86.904 193.428 ; 
        RECT 86.368 189.054 86.472 193.428 ; 
        RECT 85.936 189.054 86.04 193.428 ; 
        RECT 85.504 189.054 85.608 193.428 ; 
        RECT 85.072 189.054 85.176 193.428 ; 
        RECT 84.64 189.054 84.744 193.428 ; 
        RECT 84.208 189.054 84.312 193.428 ; 
        RECT 83.776 189.054 83.88 193.428 ; 
        RECT 83.344 189.054 83.448 193.428 ; 
        RECT 82.912 189.054 83.016 193.428 ; 
        RECT 82.48 189.054 82.584 193.428 ; 
        RECT 82.048 189.054 82.152 193.428 ; 
        RECT 81.616 189.054 81.72 193.428 ; 
        RECT 81.184 189.054 81.288 193.428 ; 
        RECT 80.752 189.054 80.856 193.428 ; 
        RECT 80.32 189.054 80.424 193.428 ; 
        RECT 79.888 189.054 79.992 193.428 ; 
        RECT 79.456 189.054 79.56 193.428 ; 
        RECT 79.024 189.054 79.128 193.428 ; 
        RECT 78.592 189.054 78.696 193.428 ; 
        RECT 78.16 189.054 78.264 193.428 ; 
        RECT 77.728 189.054 77.832 193.428 ; 
        RECT 77.296 189.054 77.4 193.428 ; 
        RECT 76.864 189.054 76.968 193.428 ; 
        RECT 76.432 189.054 76.536 193.428 ; 
        RECT 76 189.054 76.104 193.428 ; 
        RECT 75.568 189.054 75.672 193.428 ; 
        RECT 75.136 189.054 75.24 193.428 ; 
        RECT 74.704 189.054 74.808 193.428 ; 
        RECT 74.272 189.054 74.376 193.428 ; 
        RECT 73.84 189.054 73.944 193.428 ; 
        RECT 73.408 189.054 73.512 193.428 ; 
        RECT 72.976 189.054 73.08 193.428 ; 
        RECT 72.544 189.054 72.648 193.428 ; 
        RECT 72.112 189.054 72.216 193.428 ; 
        RECT 71.68 189.054 71.784 193.428 ; 
        RECT 71.248 189.054 71.352 193.428 ; 
        RECT 70.816 189.054 70.92 193.428 ; 
        RECT 70.384 189.054 70.488 193.428 ; 
        RECT 69.952 189.054 70.056 193.428 ; 
        RECT 69.52 189.054 69.624 193.428 ; 
        RECT 69.088 189.054 69.192 193.428 ; 
        RECT 68.656 189.054 68.76 193.428 ; 
        RECT 68.224 189.054 68.328 193.428 ; 
        RECT 67.792 189.054 67.896 193.428 ; 
        RECT 67.36 189.054 67.464 193.428 ; 
        RECT 66.928 189.054 67.032 193.428 ; 
        RECT 66.496 189.054 66.6 193.428 ; 
        RECT 66.064 189.054 66.168 193.428 ; 
        RECT 65.632 189.054 65.736 193.428 ; 
        RECT 65.2 189.054 65.304 193.428 ; 
        RECT 64.348 189.054 64.656 193.428 ; 
        RECT 56.776 189.054 57.084 193.428 ; 
        RECT 56.128 189.054 56.232 193.428 ; 
        RECT 55.696 189.054 55.8 193.428 ; 
        RECT 55.264 189.054 55.368 193.428 ; 
        RECT 54.832 189.054 54.936 193.428 ; 
        RECT 54.4 189.054 54.504 193.428 ; 
        RECT 53.968 189.054 54.072 193.428 ; 
        RECT 53.536 189.054 53.64 193.428 ; 
        RECT 53.104 189.054 53.208 193.428 ; 
        RECT 52.672 189.054 52.776 193.428 ; 
        RECT 52.24 189.054 52.344 193.428 ; 
        RECT 51.808 189.054 51.912 193.428 ; 
        RECT 51.376 189.054 51.48 193.428 ; 
        RECT 50.944 189.054 51.048 193.428 ; 
        RECT 50.512 189.054 50.616 193.428 ; 
        RECT 50.08 189.054 50.184 193.428 ; 
        RECT 49.648 189.054 49.752 193.428 ; 
        RECT 49.216 189.054 49.32 193.428 ; 
        RECT 48.784 189.054 48.888 193.428 ; 
        RECT 48.352 189.054 48.456 193.428 ; 
        RECT 47.92 189.054 48.024 193.428 ; 
        RECT 47.488 189.054 47.592 193.428 ; 
        RECT 47.056 189.054 47.16 193.428 ; 
        RECT 46.624 189.054 46.728 193.428 ; 
        RECT 46.192 189.054 46.296 193.428 ; 
        RECT 45.76 189.054 45.864 193.428 ; 
        RECT 45.328 189.054 45.432 193.428 ; 
        RECT 44.896 189.054 45 193.428 ; 
        RECT 44.464 189.054 44.568 193.428 ; 
        RECT 44.032 189.054 44.136 193.428 ; 
        RECT 43.6 189.054 43.704 193.428 ; 
        RECT 43.168 189.054 43.272 193.428 ; 
        RECT 42.736 189.054 42.84 193.428 ; 
        RECT 42.304 189.054 42.408 193.428 ; 
        RECT 41.872 189.054 41.976 193.428 ; 
        RECT 41.44 189.054 41.544 193.428 ; 
        RECT 41.008 189.054 41.112 193.428 ; 
        RECT 40.576 189.054 40.68 193.428 ; 
        RECT 40.144 189.054 40.248 193.428 ; 
        RECT 39.712 189.054 39.816 193.428 ; 
        RECT 39.28 189.054 39.384 193.428 ; 
        RECT 38.848 189.054 38.952 193.428 ; 
        RECT 38.416 189.054 38.52 193.428 ; 
        RECT 37.984 189.054 38.088 193.428 ; 
        RECT 37.552 189.054 37.656 193.428 ; 
        RECT 37.12 189.054 37.224 193.428 ; 
        RECT 36.688 189.054 36.792 193.428 ; 
        RECT 36.256 189.054 36.36 193.428 ; 
        RECT 35.824 189.054 35.928 193.428 ; 
        RECT 35.392 189.054 35.496 193.428 ; 
        RECT 34.96 189.054 35.064 193.428 ; 
        RECT 34.528 189.054 34.632 193.428 ; 
        RECT 34.096 189.054 34.2 193.428 ; 
        RECT 33.664 189.054 33.768 193.428 ; 
        RECT 33.232 189.054 33.336 193.428 ; 
        RECT 32.8 189.054 32.904 193.428 ; 
        RECT 32.368 189.054 32.472 193.428 ; 
        RECT 31.936 189.054 32.04 193.428 ; 
        RECT 31.504 189.054 31.608 193.428 ; 
        RECT 31.072 189.054 31.176 193.428 ; 
        RECT 30.64 189.054 30.744 193.428 ; 
        RECT 30.208 189.054 30.312 193.428 ; 
        RECT 29.776 189.054 29.88 193.428 ; 
        RECT 29.344 189.054 29.448 193.428 ; 
        RECT 28.912 189.054 29.016 193.428 ; 
        RECT 28.48 189.054 28.584 193.428 ; 
        RECT 28.048 189.054 28.152 193.428 ; 
        RECT 27.616 189.054 27.72 193.428 ; 
        RECT 27.184 189.054 27.288 193.428 ; 
        RECT 26.752 189.054 26.856 193.428 ; 
        RECT 26.32 189.054 26.424 193.428 ; 
        RECT 25.888 189.054 25.992 193.428 ; 
        RECT 25.456 189.054 25.56 193.428 ; 
        RECT 25.024 189.054 25.128 193.428 ; 
        RECT 24.592 189.054 24.696 193.428 ; 
        RECT 24.16 189.054 24.264 193.428 ; 
        RECT 23.728 189.054 23.832 193.428 ; 
        RECT 23.296 189.054 23.4 193.428 ; 
        RECT 22.864 189.054 22.968 193.428 ; 
        RECT 22.432 189.054 22.536 193.428 ; 
        RECT 22 189.054 22.104 193.428 ; 
        RECT 21.568 189.054 21.672 193.428 ; 
        RECT 21.136 189.054 21.24 193.428 ; 
        RECT 20.704 189.054 20.808 193.428 ; 
        RECT 20.272 189.054 20.376 193.428 ; 
        RECT 19.84 189.054 19.944 193.428 ; 
        RECT 19.408 189.054 19.512 193.428 ; 
        RECT 18.976 189.054 19.08 193.428 ; 
        RECT 18.544 189.054 18.648 193.428 ; 
        RECT 18.112 189.054 18.216 193.428 ; 
        RECT 17.68 189.054 17.784 193.428 ; 
        RECT 17.248 189.054 17.352 193.428 ; 
        RECT 16.816 189.054 16.92 193.428 ; 
        RECT 16.384 189.054 16.488 193.428 ; 
        RECT 15.952 189.054 16.056 193.428 ; 
        RECT 15.52 189.054 15.624 193.428 ; 
        RECT 15.088 189.054 15.192 193.428 ; 
        RECT 14.656 189.054 14.76 193.428 ; 
        RECT 14.224 189.054 14.328 193.428 ; 
        RECT 13.792 189.054 13.896 193.428 ; 
        RECT 13.36 189.054 13.464 193.428 ; 
        RECT 12.928 189.054 13.032 193.428 ; 
        RECT 12.496 189.054 12.6 193.428 ; 
        RECT 12.064 189.054 12.168 193.428 ; 
        RECT 11.632 189.054 11.736 193.428 ; 
        RECT 11.2 189.054 11.304 193.428 ; 
        RECT 10.768 189.054 10.872 193.428 ; 
        RECT 10.336 189.054 10.44 193.428 ; 
        RECT 9.904 189.054 10.008 193.428 ; 
        RECT 9.472 189.054 9.576 193.428 ; 
        RECT 9.04 189.054 9.144 193.428 ; 
        RECT 8.608 189.054 8.712 193.428 ; 
        RECT 8.176 189.054 8.28 193.428 ; 
        RECT 7.744 189.054 7.848 193.428 ; 
        RECT 7.312 189.054 7.416 193.428 ; 
        RECT 6.88 189.054 6.984 193.428 ; 
        RECT 6.448 189.054 6.552 193.428 ; 
        RECT 6.016 189.054 6.12 193.428 ; 
        RECT 5.584 189.054 5.688 193.428 ; 
        RECT 5.152 189.054 5.256 193.428 ; 
        RECT 4.72 189.054 4.824 193.428 ; 
        RECT 4.288 189.054 4.392 193.428 ; 
        RECT 3.856 189.054 3.96 193.428 ; 
        RECT 3.424 189.054 3.528 193.428 ; 
        RECT 2.992 189.054 3.096 193.428 ; 
        RECT 2.56 189.054 2.664 193.428 ; 
        RECT 2.128 189.054 2.232 193.428 ; 
        RECT 1.696 189.054 1.8 193.428 ; 
        RECT 1.264 189.054 1.368 193.428 ; 
        RECT 0.832 189.054 0.936 193.428 ; 
        RECT 0.02 189.054 0.36 193.428 ; 
        RECT 62.212 193.374 62.724 197.748 ; 
        RECT 62.156 196.036 62.724 197.326 ; 
        RECT 61.276 194.944 61.812 197.748 ; 
        RECT 61.184 196.284 61.812 197.316 ; 
        RECT 61.276 193.374 61.668 197.748 ; 
        RECT 61.276 193.858 61.724 194.816 ; 
        RECT 61.276 193.374 61.812 193.73 ; 
        RECT 60.376 195.176 60.912 197.748 ; 
        RECT 60.376 193.374 60.768 197.748 ; 
        RECT 58.708 193.374 59.04 197.748 ; 
        RECT 58.708 193.728 59.096 197.47 ; 
        RECT 121.072 193.374 121.412 197.748 ; 
        RECT 120.496 193.374 120.6 197.748 ; 
        RECT 120.064 193.374 120.168 197.748 ; 
        RECT 119.632 193.374 119.736 197.748 ; 
        RECT 119.2 193.374 119.304 197.748 ; 
        RECT 118.768 193.374 118.872 197.748 ; 
        RECT 118.336 193.374 118.44 197.748 ; 
        RECT 117.904 193.374 118.008 197.748 ; 
        RECT 117.472 193.374 117.576 197.748 ; 
        RECT 117.04 193.374 117.144 197.748 ; 
        RECT 116.608 193.374 116.712 197.748 ; 
        RECT 116.176 193.374 116.28 197.748 ; 
        RECT 115.744 193.374 115.848 197.748 ; 
        RECT 115.312 193.374 115.416 197.748 ; 
        RECT 114.88 193.374 114.984 197.748 ; 
        RECT 114.448 193.374 114.552 197.748 ; 
        RECT 114.016 193.374 114.12 197.748 ; 
        RECT 113.584 193.374 113.688 197.748 ; 
        RECT 113.152 193.374 113.256 197.748 ; 
        RECT 112.72 193.374 112.824 197.748 ; 
        RECT 112.288 193.374 112.392 197.748 ; 
        RECT 111.856 193.374 111.96 197.748 ; 
        RECT 111.424 193.374 111.528 197.748 ; 
        RECT 110.992 193.374 111.096 197.748 ; 
        RECT 110.56 193.374 110.664 197.748 ; 
        RECT 110.128 193.374 110.232 197.748 ; 
        RECT 109.696 193.374 109.8 197.748 ; 
        RECT 109.264 193.374 109.368 197.748 ; 
        RECT 108.832 193.374 108.936 197.748 ; 
        RECT 108.4 193.374 108.504 197.748 ; 
        RECT 107.968 193.374 108.072 197.748 ; 
        RECT 107.536 193.374 107.64 197.748 ; 
        RECT 107.104 193.374 107.208 197.748 ; 
        RECT 106.672 193.374 106.776 197.748 ; 
        RECT 106.24 193.374 106.344 197.748 ; 
        RECT 105.808 193.374 105.912 197.748 ; 
        RECT 105.376 193.374 105.48 197.748 ; 
        RECT 104.944 193.374 105.048 197.748 ; 
        RECT 104.512 193.374 104.616 197.748 ; 
        RECT 104.08 193.374 104.184 197.748 ; 
        RECT 103.648 193.374 103.752 197.748 ; 
        RECT 103.216 193.374 103.32 197.748 ; 
        RECT 102.784 193.374 102.888 197.748 ; 
        RECT 102.352 193.374 102.456 197.748 ; 
        RECT 101.92 193.374 102.024 197.748 ; 
        RECT 101.488 193.374 101.592 197.748 ; 
        RECT 101.056 193.374 101.16 197.748 ; 
        RECT 100.624 193.374 100.728 197.748 ; 
        RECT 100.192 193.374 100.296 197.748 ; 
        RECT 99.76 193.374 99.864 197.748 ; 
        RECT 99.328 193.374 99.432 197.748 ; 
        RECT 98.896 193.374 99 197.748 ; 
        RECT 98.464 193.374 98.568 197.748 ; 
        RECT 98.032 193.374 98.136 197.748 ; 
        RECT 97.6 193.374 97.704 197.748 ; 
        RECT 97.168 193.374 97.272 197.748 ; 
        RECT 96.736 193.374 96.84 197.748 ; 
        RECT 96.304 193.374 96.408 197.748 ; 
        RECT 95.872 193.374 95.976 197.748 ; 
        RECT 95.44 193.374 95.544 197.748 ; 
        RECT 95.008 193.374 95.112 197.748 ; 
        RECT 94.576 193.374 94.68 197.748 ; 
        RECT 94.144 193.374 94.248 197.748 ; 
        RECT 93.712 193.374 93.816 197.748 ; 
        RECT 93.28 193.374 93.384 197.748 ; 
        RECT 92.848 193.374 92.952 197.748 ; 
        RECT 92.416 193.374 92.52 197.748 ; 
        RECT 91.984 193.374 92.088 197.748 ; 
        RECT 91.552 193.374 91.656 197.748 ; 
        RECT 91.12 193.374 91.224 197.748 ; 
        RECT 90.688 193.374 90.792 197.748 ; 
        RECT 90.256 193.374 90.36 197.748 ; 
        RECT 89.824 193.374 89.928 197.748 ; 
        RECT 89.392 193.374 89.496 197.748 ; 
        RECT 88.96 193.374 89.064 197.748 ; 
        RECT 88.528 193.374 88.632 197.748 ; 
        RECT 88.096 193.374 88.2 197.748 ; 
        RECT 87.664 193.374 87.768 197.748 ; 
        RECT 87.232 193.374 87.336 197.748 ; 
        RECT 86.8 193.374 86.904 197.748 ; 
        RECT 86.368 193.374 86.472 197.748 ; 
        RECT 85.936 193.374 86.04 197.748 ; 
        RECT 85.504 193.374 85.608 197.748 ; 
        RECT 85.072 193.374 85.176 197.748 ; 
        RECT 84.64 193.374 84.744 197.748 ; 
        RECT 84.208 193.374 84.312 197.748 ; 
        RECT 83.776 193.374 83.88 197.748 ; 
        RECT 83.344 193.374 83.448 197.748 ; 
        RECT 82.912 193.374 83.016 197.748 ; 
        RECT 82.48 193.374 82.584 197.748 ; 
        RECT 82.048 193.374 82.152 197.748 ; 
        RECT 81.616 193.374 81.72 197.748 ; 
        RECT 81.184 193.374 81.288 197.748 ; 
        RECT 80.752 193.374 80.856 197.748 ; 
        RECT 80.32 193.374 80.424 197.748 ; 
        RECT 79.888 193.374 79.992 197.748 ; 
        RECT 79.456 193.374 79.56 197.748 ; 
        RECT 79.024 193.374 79.128 197.748 ; 
        RECT 78.592 193.374 78.696 197.748 ; 
        RECT 78.16 193.374 78.264 197.748 ; 
        RECT 77.728 193.374 77.832 197.748 ; 
        RECT 77.296 193.374 77.4 197.748 ; 
        RECT 76.864 193.374 76.968 197.748 ; 
        RECT 76.432 193.374 76.536 197.748 ; 
        RECT 76 193.374 76.104 197.748 ; 
        RECT 75.568 193.374 75.672 197.748 ; 
        RECT 75.136 193.374 75.24 197.748 ; 
        RECT 74.704 193.374 74.808 197.748 ; 
        RECT 74.272 193.374 74.376 197.748 ; 
        RECT 73.84 193.374 73.944 197.748 ; 
        RECT 73.408 193.374 73.512 197.748 ; 
        RECT 72.976 193.374 73.08 197.748 ; 
        RECT 72.544 193.374 72.648 197.748 ; 
        RECT 72.112 193.374 72.216 197.748 ; 
        RECT 71.68 193.374 71.784 197.748 ; 
        RECT 71.248 193.374 71.352 197.748 ; 
        RECT 70.816 193.374 70.92 197.748 ; 
        RECT 70.384 193.374 70.488 197.748 ; 
        RECT 69.952 193.374 70.056 197.748 ; 
        RECT 69.52 193.374 69.624 197.748 ; 
        RECT 69.088 193.374 69.192 197.748 ; 
        RECT 68.656 193.374 68.76 197.748 ; 
        RECT 68.224 193.374 68.328 197.748 ; 
        RECT 67.792 193.374 67.896 197.748 ; 
        RECT 67.36 193.374 67.464 197.748 ; 
        RECT 66.928 193.374 67.032 197.748 ; 
        RECT 66.496 193.374 66.6 197.748 ; 
        RECT 66.064 193.374 66.168 197.748 ; 
        RECT 65.632 193.374 65.736 197.748 ; 
        RECT 65.2 193.374 65.304 197.748 ; 
        RECT 64.348 193.374 64.656 197.748 ; 
        RECT 56.776 193.374 57.084 197.748 ; 
        RECT 56.128 193.374 56.232 197.748 ; 
        RECT 55.696 193.374 55.8 197.748 ; 
        RECT 55.264 193.374 55.368 197.748 ; 
        RECT 54.832 193.374 54.936 197.748 ; 
        RECT 54.4 193.374 54.504 197.748 ; 
        RECT 53.968 193.374 54.072 197.748 ; 
        RECT 53.536 193.374 53.64 197.748 ; 
        RECT 53.104 193.374 53.208 197.748 ; 
        RECT 52.672 193.374 52.776 197.748 ; 
        RECT 52.24 193.374 52.344 197.748 ; 
        RECT 51.808 193.374 51.912 197.748 ; 
        RECT 51.376 193.374 51.48 197.748 ; 
        RECT 50.944 193.374 51.048 197.748 ; 
        RECT 50.512 193.374 50.616 197.748 ; 
        RECT 50.08 193.374 50.184 197.748 ; 
        RECT 49.648 193.374 49.752 197.748 ; 
        RECT 49.216 193.374 49.32 197.748 ; 
        RECT 48.784 193.374 48.888 197.748 ; 
        RECT 48.352 193.374 48.456 197.748 ; 
        RECT 47.92 193.374 48.024 197.748 ; 
        RECT 47.488 193.374 47.592 197.748 ; 
        RECT 47.056 193.374 47.16 197.748 ; 
        RECT 46.624 193.374 46.728 197.748 ; 
        RECT 46.192 193.374 46.296 197.748 ; 
        RECT 45.76 193.374 45.864 197.748 ; 
        RECT 45.328 193.374 45.432 197.748 ; 
        RECT 44.896 193.374 45 197.748 ; 
        RECT 44.464 193.374 44.568 197.748 ; 
        RECT 44.032 193.374 44.136 197.748 ; 
        RECT 43.6 193.374 43.704 197.748 ; 
        RECT 43.168 193.374 43.272 197.748 ; 
        RECT 42.736 193.374 42.84 197.748 ; 
        RECT 42.304 193.374 42.408 197.748 ; 
        RECT 41.872 193.374 41.976 197.748 ; 
        RECT 41.44 193.374 41.544 197.748 ; 
        RECT 41.008 193.374 41.112 197.748 ; 
        RECT 40.576 193.374 40.68 197.748 ; 
        RECT 40.144 193.374 40.248 197.748 ; 
        RECT 39.712 193.374 39.816 197.748 ; 
        RECT 39.28 193.374 39.384 197.748 ; 
        RECT 38.848 193.374 38.952 197.748 ; 
        RECT 38.416 193.374 38.52 197.748 ; 
        RECT 37.984 193.374 38.088 197.748 ; 
        RECT 37.552 193.374 37.656 197.748 ; 
        RECT 37.12 193.374 37.224 197.748 ; 
        RECT 36.688 193.374 36.792 197.748 ; 
        RECT 36.256 193.374 36.36 197.748 ; 
        RECT 35.824 193.374 35.928 197.748 ; 
        RECT 35.392 193.374 35.496 197.748 ; 
        RECT 34.96 193.374 35.064 197.748 ; 
        RECT 34.528 193.374 34.632 197.748 ; 
        RECT 34.096 193.374 34.2 197.748 ; 
        RECT 33.664 193.374 33.768 197.748 ; 
        RECT 33.232 193.374 33.336 197.748 ; 
        RECT 32.8 193.374 32.904 197.748 ; 
        RECT 32.368 193.374 32.472 197.748 ; 
        RECT 31.936 193.374 32.04 197.748 ; 
        RECT 31.504 193.374 31.608 197.748 ; 
        RECT 31.072 193.374 31.176 197.748 ; 
        RECT 30.64 193.374 30.744 197.748 ; 
        RECT 30.208 193.374 30.312 197.748 ; 
        RECT 29.776 193.374 29.88 197.748 ; 
        RECT 29.344 193.374 29.448 197.748 ; 
        RECT 28.912 193.374 29.016 197.748 ; 
        RECT 28.48 193.374 28.584 197.748 ; 
        RECT 28.048 193.374 28.152 197.748 ; 
        RECT 27.616 193.374 27.72 197.748 ; 
        RECT 27.184 193.374 27.288 197.748 ; 
        RECT 26.752 193.374 26.856 197.748 ; 
        RECT 26.32 193.374 26.424 197.748 ; 
        RECT 25.888 193.374 25.992 197.748 ; 
        RECT 25.456 193.374 25.56 197.748 ; 
        RECT 25.024 193.374 25.128 197.748 ; 
        RECT 24.592 193.374 24.696 197.748 ; 
        RECT 24.16 193.374 24.264 197.748 ; 
        RECT 23.728 193.374 23.832 197.748 ; 
        RECT 23.296 193.374 23.4 197.748 ; 
        RECT 22.864 193.374 22.968 197.748 ; 
        RECT 22.432 193.374 22.536 197.748 ; 
        RECT 22 193.374 22.104 197.748 ; 
        RECT 21.568 193.374 21.672 197.748 ; 
        RECT 21.136 193.374 21.24 197.748 ; 
        RECT 20.704 193.374 20.808 197.748 ; 
        RECT 20.272 193.374 20.376 197.748 ; 
        RECT 19.84 193.374 19.944 197.748 ; 
        RECT 19.408 193.374 19.512 197.748 ; 
        RECT 18.976 193.374 19.08 197.748 ; 
        RECT 18.544 193.374 18.648 197.748 ; 
        RECT 18.112 193.374 18.216 197.748 ; 
        RECT 17.68 193.374 17.784 197.748 ; 
        RECT 17.248 193.374 17.352 197.748 ; 
        RECT 16.816 193.374 16.92 197.748 ; 
        RECT 16.384 193.374 16.488 197.748 ; 
        RECT 15.952 193.374 16.056 197.748 ; 
        RECT 15.52 193.374 15.624 197.748 ; 
        RECT 15.088 193.374 15.192 197.748 ; 
        RECT 14.656 193.374 14.76 197.748 ; 
        RECT 14.224 193.374 14.328 197.748 ; 
        RECT 13.792 193.374 13.896 197.748 ; 
        RECT 13.36 193.374 13.464 197.748 ; 
        RECT 12.928 193.374 13.032 197.748 ; 
        RECT 12.496 193.374 12.6 197.748 ; 
        RECT 12.064 193.374 12.168 197.748 ; 
        RECT 11.632 193.374 11.736 197.748 ; 
        RECT 11.2 193.374 11.304 197.748 ; 
        RECT 10.768 193.374 10.872 197.748 ; 
        RECT 10.336 193.374 10.44 197.748 ; 
        RECT 9.904 193.374 10.008 197.748 ; 
        RECT 9.472 193.374 9.576 197.748 ; 
        RECT 9.04 193.374 9.144 197.748 ; 
        RECT 8.608 193.374 8.712 197.748 ; 
        RECT 8.176 193.374 8.28 197.748 ; 
        RECT 7.744 193.374 7.848 197.748 ; 
        RECT 7.312 193.374 7.416 197.748 ; 
        RECT 6.88 193.374 6.984 197.748 ; 
        RECT 6.448 193.374 6.552 197.748 ; 
        RECT 6.016 193.374 6.12 197.748 ; 
        RECT 5.584 193.374 5.688 197.748 ; 
        RECT 5.152 193.374 5.256 197.748 ; 
        RECT 4.72 193.374 4.824 197.748 ; 
        RECT 4.288 193.374 4.392 197.748 ; 
        RECT 3.856 193.374 3.96 197.748 ; 
        RECT 3.424 193.374 3.528 197.748 ; 
        RECT 2.992 193.374 3.096 197.748 ; 
        RECT 2.56 193.374 2.664 197.748 ; 
        RECT 2.128 193.374 2.232 197.748 ; 
        RECT 1.696 193.374 1.8 197.748 ; 
        RECT 1.264 193.374 1.368 197.748 ; 
        RECT 0.832 193.374 0.936 197.748 ; 
        RECT 0.02 193.374 0.36 197.748 ; 
        RECT 62.212 197.694 62.724 202.068 ; 
        RECT 62.156 200.356 62.724 201.646 ; 
        RECT 61.276 199.264 61.812 202.068 ; 
        RECT 61.184 200.604 61.812 201.636 ; 
        RECT 61.276 197.694 61.668 202.068 ; 
        RECT 61.276 198.178 61.724 199.136 ; 
        RECT 61.276 197.694 61.812 198.05 ; 
        RECT 60.376 199.496 60.912 202.068 ; 
        RECT 60.376 197.694 60.768 202.068 ; 
        RECT 58.708 197.694 59.04 202.068 ; 
        RECT 58.708 198.048 59.096 201.79 ; 
        RECT 121.072 197.694 121.412 202.068 ; 
        RECT 120.496 197.694 120.6 202.068 ; 
        RECT 120.064 197.694 120.168 202.068 ; 
        RECT 119.632 197.694 119.736 202.068 ; 
        RECT 119.2 197.694 119.304 202.068 ; 
        RECT 118.768 197.694 118.872 202.068 ; 
        RECT 118.336 197.694 118.44 202.068 ; 
        RECT 117.904 197.694 118.008 202.068 ; 
        RECT 117.472 197.694 117.576 202.068 ; 
        RECT 117.04 197.694 117.144 202.068 ; 
        RECT 116.608 197.694 116.712 202.068 ; 
        RECT 116.176 197.694 116.28 202.068 ; 
        RECT 115.744 197.694 115.848 202.068 ; 
        RECT 115.312 197.694 115.416 202.068 ; 
        RECT 114.88 197.694 114.984 202.068 ; 
        RECT 114.448 197.694 114.552 202.068 ; 
        RECT 114.016 197.694 114.12 202.068 ; 
        RECT 113.584 197.694 113.688 202.068 ; 
        RECT 113.152 197.694 113.256 202.068 ; 
        RECT 112.72 197.694 112.824 202.068 ; 
        RECT 112.288 197.694 112.392 202.068 ; 
        RECT 111.856 197.694 111.96 202.068 ; 
        RECT 111.424 197.694 111.528 202.068 ; 
        RECT 110.992 197.694 111.096 202.068 ; 
        RECT 110.56 197.694 110.664 202.068 ; 
        RECT 110.128 197.694 110.232 202.068 ; 
        RECT 109.696 197.694 109.8 202.068 ; 
        RECT 109.264 197.694 109.368 202.068 ; 
        RECT 108.832 197.694 108.936 202.068 ; 
        RECT 108.4 197.694 108.504 202.068 ; 
        RECT 107.968 197.694 108.072 202.068 ; 
        RECT 107.536 197.694 107.64 202.068 ; 
        RECT 107.104 197.694 107.208 202.068 ; 
        RECT 106.672 197.694 106.776 202.068 ; 
        RECT 106.24 197.694 106.344 202.068 ; 
        RECT 105.808 197.694 105.912 202.068 ; 
        RECT 105.376 197.694 105.48 202.068 ; 
        RECT 104.944 197.694 105.048 202.068 ; 
        RECT 104.512 197.694 104.616 202.068 ; 
        RECT 104.08 197.694 104.184 202.068 ; 
        RECT 103.648 197.694 103.752 202.068 ; 
        RECT 103.216 197.694 103.32 202.068 ; 
        RECT 102.784 197.694 102.888 202.068 ; 
        RECT 102.352 197.694 102.456 202.068 ; 
        RECT 101.92 197.694 102.024 202.068 ; 
        RECT 101.488 197.694 101.592 202.068 ; 
        RECT 101.056 197.694 101.16 202.068 ; 
        RECT 100.624 197.694 100.728 202.068 ; 
        RECT 100.192 197.694 100.296 202.068 ; 
        RECT 99.76 197.694 99.864 202.068 ; 
        RECT 99.328 197.694 99.432 202.068 ; 
        RECT 98.896 197.694 99 202.068 ; 
        RECT 98.464 197.694 98.568 202.068 ; 
        RECT 98.032 197.694 98.136 202.068 ; 
        RECT 97.6 197.694 97.704 202.068 ; 
        RECT 97.168 197.694 97.272 202.068 ; 
        RECT 96.736 197.694 96.84 202.068 ; 
        RECT 96.304 197.694 96.408 202.068 ; 
        RECT 95.872 197.694 95.976 202.068 ; 
        RECT 95.44 197.694 95.544 202.068 ; 
        RECT 95.008 197.694 95.112 202.068 ; 
        RECT 94.576 197.694 94.68 202.068 ; 
        RECT 94.144 197.694 94.248 202.068 ; 
        RECT 93.712 197.694 93.816 202.068 ; 
        RECT 93.28 197.694 93.384 202.068 ; 
        RECT 92.848 197.694 92.952 202.068 ; 
        RECT 92.416 197.694 92.52 202.068 ; 
        RECT 91.984 197.694 92.088 202.068 ; 
        RECT 91.552 197.694 91.656 202.068 ; 
        RECT 91.12 197.694 91.224 202.068 ; 
        RECT 90.688 197.694 90.792 202.068 ; 
        RECT 90.256 197.694 90.36 202.068 ; 
        RECT 89.824 197.694 89.928 202.068 ; 
        RECT 89.392 197.694 89.496 202.068 ; 
        RECT 88.96 197.694 89.064 202.068 ; 
        RECT 88.528 197.694 88.632 202.068 ; 
        RECT 88.096 197.694 88.2 202.068 ; 
        RECT 87.664 197.694 87.768 202.068 ; 
        RECT 87.232 197.694 87.336 202.068 ; 
        RECT 86.8 197.694 86.904 202.068 ; 
        RECT 86.368 197.694 86.472 202.068 ; 
        RECT 85.936 197.694 86.04 202.068 ; 
        RECT 85.504 197.694 85.608 202.068 ; 
        RECT 85.072 197.694 85.176 202.068 ; 
        RECT 84.64 197.694 84.744 202.068 ; 
        RECT 84.208 197.694 84.312 202.068 ; 
        RECT 83.776 197.694 83.88 202.068 ; 
        RECT 83.344 197.694 83.448 202.068 ; 
        RECT 82.912 197.694 83.016 202.068 ; 
        RECT 82.48 197.694 82.584 202.068 ; 
        RECT 82.048 197.694 82.152 202.068 ; 
        RECT 81.616 197.694 81.72 202.068 ; 
        RECT 81.184 197.694 81.288 202.068 ; 
        RECT 80.752 197.694 80.856 202.068 ; 
        RECT 80.32 197.694 80.424 202.068 ; 
        RECT 79.888 197.694 79.992 202.068 ; 
        RECT 79.456 197.694 79.56 202.068 ; 
        RECT 79.024 197.694 79.128 202.068 ; 
        RECT 78.592 197.694 78.696 202.068 ; 
        RECT 78.16 197.694 78.264 202.068 ; 
        RECT 77.728 197.694 77.832 202.068 ; 
        RECT 77.296 197.694 77.4 202.068 ; 
        RECT 76.864 197.694 76.968 202.068 ; 
        RECT 76.432 197.694 76.536 202.068 ; 
        RECT 76 197.694 76.104 202.068 ; 
        RECT 75.568 197.694 75.672 202.068 ; 
        RECT 75.136 197.694 75.24 202.068 ; 
        RECT 74.704 197.694 74.808 202.068 ; 
        RECT 74.272 197.694 74.376 202.068 ; 
        RECT 73.84 197.694 73.944 202.068 ; 
        RECT 73.408 197.694 73.512 202.068 ; 
        RECT 72.976 197.694 73.08 202.068 ; 
        RECT 72.544 197.694 72.648 202.068 ; 
        RECT 72.112 197.694 72.216 202.068 ; 
        RECT 71.68 197.694 71.784 202.068 ; 
        RECT 71.248 197.694 71.352 202.068 ; 
        RECT 70.816 197.694 70.92 202.068 ; 
        RECT 70.384 197.694 70.488 202.068 ; 
        RECT 69.952 197.694 70.056 202.068 ; 
        RECT 69.52 197.694 69.624 202.068 ; 
        RECT 69.088 197.694 69.192 202.068 ; 
        RECT 68.656 197.694 68.76 202.068 ; 
        RECT 68.224 197.694 68.328 202.068 ; 
        RECT 67.792 197.694 67.896 202.068 ; 
        RECT 67.36 197.694 67.464 202.068 ; 
        RECT 66.928 197.694 67.032 202.068 ; 
        RECT 66.496 197.694 66.6 202.068 ; 
        RECT 66.064 197.694 66.168 202.068 ; 
        RECT 65.632 197.694 65.736 202.068 ; 
        RECT 65.2 197.694 65.304 202.068 ; 
        RECT 64.348 197.694 64.656 202.068 ; 
        RECT 56.776 197.694 57.084 202.068 ; 
        RECT 56.128 197.694 56.232 202.068 ; 
        RECT 55.696 197.694 55.8 202.068 ; 
        RECT 55.264 197.694 55.368 202.068 ; 
        RECT 54.832 197.694 54.936 202.068 ; 
        RECT 54.4 197.694 54.504 202.068 ; 
        RECT 53.968 197.694 54.072 202.068 ; 
        RECT 53.536 197.694 53.64 202.068 ; 
        RECT 53.104 197.694 53.208 202.068 ; 
        RECT 52.672 197.694 52.776 202.068 ; 
        RECT 52.24 197.694 52.344 202.068 ; 
        RECT 51.808 197.694 51.912 202.068 ; 
        RECT 51.376 197.694 51.48 202.068 ; 
        RECT 50.944 197.694 51.048 202.068 ; 
        RECT 50.512 197.694 50.616 202.068 ; 
        RECT 50.08 197.694 50.184 202.068 ; 
        RECT 49.648 197.694 49.752 202.068 ; 
        RECT 49.216 197.694 49.32 202.068 ; 
        RECT 48.784 197.694 48.888 202.068 ; 
        RECT 48.352 197.694 48.456 202.068 ; 
        RECT 47.92 197.694 48.024 202.068 ; 
        RECT 47.488 197.694 47.592 202.068 ; 
        RECT 47.056 197.694 47.16 202.068 ; 
        RECT 46.624 197.694 46.728 202.068 ; 
        RECT 46.192 197.694 46.296 202.068 ; 
        RECT 45.76 197.694 45.864 202.068 ; 
        RECT 45.328 197.694 45.432 202.068 ; 
        RECT 44.896 197.694 45 202.068 ; 
        RECT 44.464 197.694 44.568 202.068 ; 
        RECT 44.032 197.694 44.136 202.068 ; 
        RECT 43.6 197.694 43.704 202.068 ; 
        RECT 43.168 197.694 43.272 202.068 ; 
        RECT 42.736 197.694 42.84 202.068 ; 
        RECT 42.304 197.694 42.408 202.068 ; 
        RECT 41.872 197.694 41.976 202.068 ; 
        RECT 41.44 197.694 41.544 202.068 ; 
        RECT 41.008 197.694 41.112 202.068 ; 
        RECT 40.576 197.694 40.68 202.068 ; 
        RECT 40.144 197.694 40.248 202.068 ; 
        RECT 39.712 197.694 39.816 202.068 ; 
        RECT 39.28 197.694 39.384 202.068 ; 
        RECT 38.848 197.694 38.952 202.068 ; 
        RECT 38.416 197.694 38.52 202.068 ; 
        RECT 37.984 197.694 38.088 202.068 ; 
        RECT 37.552 197.694 37.656 202.068 ; 
        RECT 37.12 197.694 37.224 202.068 ; 
        RECT 36.688 197.694 36.792 202.068 ; 
        RECT 36.256 197.694 36.36 202.068 ; 
        RECT 35.824 197.694 35.928 202.068 ; 
        RECT 35.392 197.694 35.496 202.068 ; 
        RECT 34.96 197.694 35.064 202.068 ; 
        RECT 34.528 197.694 34.632 202.068 ; 
        RECT 34.096 197.694 34.2 202.068 ; 
        RECT 33.664 197.694 33.768 202.068 ; 
        RECT 33.232 197.694 33.336 202.068 ; 
        RECT 32.8 197.694 32.904 202.068 ; 
        RECT 32.368 197.694 32.472 202.068 ; 
        RECT 31.936 197.694 32.04 202.068 ; 
        RECT 31.504 197.694 31.608 202.068 ; 
        RECT 31.072 197.694 31.176 202.068 ; 
        RECT 30.64 197.694 30.744 202.068 ; 
        RECT 30.208 197.694 30.312 202.068 ; 
        RECT 29.776 197.694 29.88 202.068 ; 
        RECT 29.344 197.694 29.448 202.068 ; 
        RECT 28.912 197.694 29.016 202.068 ; 
        RECT 28.48 197.694 28.584 202.068 ; 
        RECT 28.048 197.694 28.152 202.068 ; 
        RECT 27.616 197.694 27.72 202.068 ; 
        RECT 27.184 197.694 27.288 202.068 ; 
        RECT 26.752 197.694 26.856 202.068 ; 
        RECT 26.32 197.694 26.424 202.068 ; 
        RECT 25.888 197.694 25.992 202.068 ; 
        RECT 25.456 197.694 25.56 202.068 ; 
        RECT 25.024 197.694 25.128 202.068 ; 
        RECT 24.592 197.694 24.696 202.068 ; 
        RECT 24.16 197.694 24.264 202.068 ; 
        RECT 23.728 197.694 23.832 202.068 ; 
        RECT 23.296 197.694 23.4 202.068 ; 
        RECT 22.864 197.694 22.968 202.068 ; 
        RECT 22.432 197.694 22.536 202.068 ; 
        RECT 22 197.694 22.104 202.068 ; 
        RECT 21.568 197.694 21.672 202.068 ; 
        RECT 21.136 197.694 21.24 202.068 ; 
        RECT 20.704 197.694 20.808 202.068 ; 
        RECT 20.272 197.694 20.376 202.068 ; 
        RECT 19.84 197.694 19.944 202.068 ; 
        RECT 19.408 197.694 19.512 202.068 ; 
        RECT 18.976 197.694 19.08 202.068 ; 
        RECT 18.544 197.694 18.648 202.068 ; 
        RECT 18.112 197.694 18.216 202.068 ; 
        RECT 17.68 197.694 17.784 202.068 ; 
        RECT 17.248 197.694 17.352 202.068 ; 
        RECT 16.816 197.694 16.92 202.068 ; 
        RECT 16.384 197.694 16.488 202.068 ; 
        RECT 15.952 197.694 16.056 202.068 ; 
        RECT 15.52 197.694 15.624 202.068 ; 
        RECT 15.088 197.694 15.192 202.068 ; 
        RECT 14.656 197.694 14.76 202.068 ; 
        RECT 14.224 197.694 14.328 202.068 ; 
        RECT 13.792 197.694 13.896 202.068 ; 
        RECT 13.36 197.694 13.464 202.068 ; 
        RECT 12.928 197.694 13.032 202.068 ; 
        RECT 12.496 197.694 12.6 202.068 ; 
        RECT 12.064 197.694 12.168 202.068 ; 
        RECT 11.632 197.694 11.736 202.068 ; 
        RECT 11.2 197.694 11.304 202.068 ; 
        RECT 10.768 197.694 10.872 202.068 ; 
        RECT 10.336 197.694 10.44 202.068 ; 
        RECT 9.904 197.694 10.008 202.068 ; 
        RECT 9.472 197.694 9.576 202.068 ; 
        RECT 9.04 197.694 9.144 202.068 ; 
        RECT 8.608 197.694 8.712 202.068 ; 
        RECT 8.176 197.694 8.28 202.068 ; 
        RECT 7.744 197.694 7.848 202.068 ; 
        RECT 7.312 197.694 7.416 202.068 ; 
        RECT 6.88 197.694 6.984 202.068 ; 
        RECT 6.448 197.694 6.552 202.068 ; 
        RECT 6.016 197.694 6.12 202.068 ; 
        RECT 5.584 197.694 5.688 202.068 ; 
        RECT 5.152 197.694 5.256 202.068 ; 
        RECT 4.72 197.694 4.824 202.068 ; 
        RECT 4.288 197.694 4.392 202.068 ; 
        RECT 3.856 197.694 3.96 202.068 ; 
        RECT 3.424 197.694 3.528 202.068 ; 
        RECT 2.992 197.694 3.096 202.068 ; 
        RECT 2.56 197.694 2.664 202.068 ; 
        RECT 2.128 197.694 2.232 202.068 ; 
        RECT 1.696 197.694 1.8 202.068 ; 
        RECT 1.264 197.694 1.368 202.068 ; 
        RECT 0.832 197.694 0.936 202.068 ; 
        RECT 0.02 197.694 0.36 202.068 ; 
        RECT 62.212 202.014 62.724 206.388 ; 
        RECT 62.156 204.676 62.724 205.966 ; 
        RECT 61.276 203.584 61.812 206.388 ; 
        RECT 61.184 204.924 61.812 205.956 ; 
        RECT 61.276 202.014 61.668 206.388 ; 
        RECT 61.276 202.498 61.724 203.456 ; 
        RECT 61.276 202.014 61.812 202.37 ; 
        RECT 60.376 203.816 60.912 206.388 ; 
        RECT 60.376 202.014 60.768 206.388 ; 
        RECT 58.708 202.014 59.04 206.388 ; 
        RECT 58.708 202.368 59.096 206.11 ; 
        RECT 121.072 202.014 121.412 206.388 ; 
        RECT 120.496 202.014 120.6 206.388 ; 
        RECT 120.064 202.014 120.168 206.388 ; 
        RECT 119.632 202.014 119.736 206.388 ; 
        RECT 119.2 202.014 119.304 206.388 ; 
        RECT 118.768 202.014 118.872 206.388 ; 
        RECT 118.336 202.014 118.44 206.388 ; 
        RECT 117.904 202.014 118.008 206.388 ; 
        RECT 117.472 202.014 117.576 206.388 ; 
        RECT 117.04 202.014 117.144 206.388 ; 
        RECT 116.608 202.014 116.712 206.388 ; 
        RECT 116.176 202.014 116.28 206.388 ; 
        RECT 115.744 202.014 115.848 206.388 ; 
        RECT 115.312 202.014 115.416 206.388 ; 
        RECT 114.88 202.014 114.984 206.388 ; 
        RECT 114.448 202.014 114.552 206.388 ; 
        RECT 114.016 202.014 114.12 206.388 ; 
        RECT 113.584 202.014 113.688 206.388 ; 
        RECT 113.152 202.014 113.256 206.388 ; 
        RECT 112.72 202.014 112.824 206.388 ; 
        RECT 112.288 202.014 112.392 206.388 ; 
        RECT 111.856 202.014 111.96 206.388 ; 
        RECT 111.424 202.014 111.528 206.388 ; 
        RECT 110.992 202.014 111.096 206.388 ; 
        RECT 110.56 202.014 110.664 206.388 ; 
        RECT 110.128 202.014 110.232 206.388 ; 
        RECT 109.696 202.014 109.8 206.388 ; 
        RECT 109.264 202.014 109.368 206.388 ; 
        RECT 108.832 202.014 108.936 206.388 ; 
        RECT 108.4 202.014 108.504 206.388 ; 
        RECT 107.968 202.014 108.072 206.388 ; 
        RECT 107.536 202.014 107.64 206.388 ; 
        RECT 107.104 202.014 107.208 206.388 ; 
        RECT 106.672 202.014 106.776 206.388 ; 
        RECT 106.24 202.014 106.344 206.388 ; 
        RECT 105.808 202.014 105.912 206.388 ; 
        RECT 105.376 202.014 105.48 206.388 ; 
        RECT 104.944 202.014 105.048 206.388 ; 
        RECT 104.512 202.014 104.616 206.388 ; 
        RECT 104.08 202.014 104.184 206.388 ; 
        RECT 103.648 202.014 103.752 206.388 ; 
        RECT 103.216 202.014 103.32 206.388 ; 
        RECT 102.784 202.014 102.888 206.388 ; 
        RECT 102.352 202.014 102.456 206.388 ; 
        RECT 101.92 202.014 102.024 206.388 ; 
        RECT 101.488 202.014 101.592 206.388 ; 
        RECT 101.056 202.014 101.16 206.388 ; 
        RECT 100.624 202.014 100.728 206.388 ; 
        RECT 100.192 202.014 100.296 206.388 ; 
        RECT 99.76 202.014 99.864 206.388 ; 
        RECT 99.328 202.014 99.432 206.388 ; 
        RECT 98.896 202.014 99 206.388 ; 
        RECT 98.464 202.014 98.568 206.388 ; 
        RECT 98.032 202.014 98.136 206.388 ; 
        RECT 97.6 202.014 97.704 206.388 ; 
        RECT 97.168 202.014 97.272 206.388 ; 
        RECT 96.736 202.014 96.84 206.388 ; 
        RECT 96.304 202.014 96.408 206.388 ; 
        RECT 95.872 202.014 95.976 206.388 ; 
        RECT 95.44 202.014 95.544 206.388 ; 
        RECT 95.008 202.014 95.112 206.388 ; 
        RECT 94.576 202.014 94.68 206.388 ; 
        RECT 94.144 202.014 94.248 206.388 ; 
        RECT 93.712 202.014 93.816 206.388 ; 
        RECT 93.28 202.014 93.384 206.388 ; 
        RECT 92.848 202.014 92.952 206.388 ; 
        RECT 92.416 202.014 92.52 206.388 ; 
        RECT 91.984 202.014 92.088 206.388 ; 
        RECT 91.552 202.014 91.656 206.388 ; 
        RECT 91.12 202.014 91.224 206.388 ; 
        RECT 90.688 202.014 90.792 206.388 ; 
        RECT 90.256 202.014 90.36 206.388 ; 
        RECT 89.824 202.014 89.928 206.388 ; 
        RECT 89.392 202.014 89.496 206.388 ; 
        RECT 88.96 202.014 89.064 206.388 ; 
        RECT 88.528 202.014 88.632 206.388 ; 
        RECT 88.096 202.014 88.2 206.388 ; 
        RECT 87.664 202.014 87.768 206.388 ; 
        RECT 87.232 202.014 87.336 206.388 ; 
        RECT 86.8 202.014 86.904 206.388 ; 
        RECT 86.368 202.014 86.472 206.388 ; 
        RECT 85.936 202.014 86.04 206.388 ; 
        RECT 85.504 202.014 85.608 206.388 ; 
        RECT 85.072 202.014 85.176 206.388 ; 
        RECT 84.64 202.014 84.744 206.388 ; 
        RECT 84.208 202.014 84.312 206.388 ; 
        RECT 83.776 202.014 83.88 206.388 ; 
        RECT 83.344 202.014 83.448 206.388 ; 
        RECT 82.912 202.014 83.016 206.388 ; 
        RECT 82.48 202.014 82.584 206.388 ; 
        RECT 82.048 202.014 82.152 206.388 ; 
        RECT 81.616 202.014 81.72 206.388 ; 
        RECT 81.184 202.014 81.288 206.388 ; 
        RECT 80.752 202.014 80.856 206.388 ; 
        RECT 80.32 202.014 80.424 206.388 ; 
        RECT 79.888 202.014 79.992 206.388 ; 
        RECT 79.456 202.014 79.56 206.388 ; 
        RECT 79.024 202.014 79.128 206.388 ; 
        RECT 78.592 202.014 78.696 206.388 ; 
        RECT 78.16 202.014 78.264 206.388 ; 
        RECT 77.728 202.014 77.832 206.388 ; 
        RECT 77.296 202.014 77.4 206.388 ; 
        RECT 76.864 202.014 76.968 206.388 ; 
        RECT 76.432 202.014 76.536 206.388 ; 
        RECT 76 202.014 76.104 206.388 ; 
        RECT 75.568 202.014 75.672 206.388 ; 
        RECT 75.136 202.014 75.24 206.388 ; 
        RECT 74.704 202.014 74.808 206.388 ; 
        RECT 74.272 202.014 74.376 206.388 ; 
        RECT 73.84 202.014 73.944 206.388 ; 
        RECT 73.408 202.014 73.512 206.388 ; 
        RECT 72.976 202.014 73.08 206.388 ; 
        RECT 72.544 202.014 72.648 206.388 ; 
        RECT 72.112 202.014 72.216 206.388 ; 
        RECT 71.68 202.014 71.784 206.388 ; 
        RECT 71.248 202.014 71.352 206.388 ; 
        RECT 70.816 202.014 70.92 206.388 ; 
        RECT 70.384 202.014 70.488 206.388 ; 
        RECT 69.952 202.014 70.056 206.388 ; 
        RECT 69.52 202.014 69.624 206.388 ; 
        RECT 69.088 202.014 69.192 206.388 ; 
        RECT 68.656 202.014 68.76 206.388 ; 
        RECT 68.224 202.014 68.328 206.388 ; 
        RECT 67.792 202.014 67.896 206.388 ; 
        RECT 67.36 202.014 67.464 206.388 ; 
        RECT 66.928 202.014 67.032 206.388 ; 
        RECT 66.496 202.014 66.6 206.388 ; 
        RECT 66.064 202.014 66.168 206.388 ; 
        RECT 65.632 202.014 65.736 206.388 ; 
        RECT 65.2 202.014 65.304 206.388 ; 
        RECT 64.348 202.014 64.656 206.388 ; 
        RECT 56.776 202.014 57.084 206.388 ; 
        RECT 56.128 202.014 56.232 206.388 ; 
        RECT 55.696 202.014 55.8 206.388 ; 
        RECT 55.264 202.014 55.368 206.388 ; 
        RECT 54.832 202.014 54.936 206.388 ; 
        RECT 54.4 202.014 54.504 206.388 ; 
        RECT 53.968 202.014 54.072 206.388 ; 
        RECT 53.536 202.014 53.64 206.388 ; 
        RECT 53.104 202.014 53.208 206.388 ; 
        RECT 52.672 202.014 52.776 206.388 ; 
        RECT 52.24 202.014 52.344 206.388 ; 
        RECT 51.808 202.014 51.912 206.388 ; 
        RECT 51.376 202.014 51.48 206.388 ; 
        RECT 50.944 202.014 51.048 206.388 ; 
        RECT 50.512 202.014 50.616 206.388 ; 
        RECT 50.08 202.014 50.184 206.388 ; 
        RECT 49.648 202.014 49.752 206.388 ; 
        RECT 49.216 202.014 49.32 206.388 ; 
        RECT 48.784 202.014 48.888 206.388 ; 
        RECT 48.352 202.014 48.456 206.388 ; 
        RECT 47.92 202.014 48.024 206.388 ; 
        RECT 47.488 202.014 47.592 206.388 ; 
        RECT 47.056 202.014 47.16 206.388 ; 
        RECT 46.624 202.014 46.728 206.388 ; 
        RECT 46.192 202.014 46.296 206.388 ; 
        RECT 45.76 202.014 45.864 206.388 ; 
        RECT 45.328 202.014 45.432 206.388 ; 
        RECT 44.896 202.014 45 206.388 ; 
        RECT 44.464 202.014 44.568 206.388 ; 
        RECT 44.032 202.014 44.136 206.388 ; 
        RECT 43.6 202.014 43.704 206.388 ; 
        RECT 43.168 202.014 43.272 206.388 ; 
        RECT 42.736 202.014 42.84 206.388 ; 
        RECT 42.304 202.014 42.408 206.388 ; 
        RECT 41.872 202.014 41.976 206.388 ; 
        RECT 41.44 202.014 41.544 206.388 ; 
        RECT 41.008 202.014 41.112 206.388 ; 
        RECT 40.576 202.014 40.68 206.388 ; 
        RECT 40.144 202.014 40.248 206.388 ; 
        RECT 39.712 202.014 39.816 206.388 ; 
        RECT 39.28 202.014 39.384 206.388 ; 
        RECT 38.848 202.014 38.952 206.388 ; 
        RECT 38.416 202.014 38.52 206.388 ; 
        RECT 37.984 202.014 38.088 206.388 ; 
        RECT 37.552 202.014 37.656 206.388 ; 
        RECT 37.12 202.014 37.224 206.388 ; 
        RECT 36.688 202.014 36.792 206.388 ; 
        RECT 36.256 202.014 36.36 206.388 ; 
        RECT 35.824 202.014 35.928 206.388 ; 
        RECT 35.392 202.014 35.496 206.388 ; 
        RECT 34.96 202.014 35.064 206.388 ; 
        RECT 34.528 202.014 34.632 206.388 ; 
        RECT 34.096 202.014 34.2 206.388 ; 
        RECT 33.664 202.014 33.768 206.388 ; 
        RECT 33.232 202.014 33.336 206.388 ; 
        RECT 32.8 202.014 32.904 206.388 ; 
        RECT 32.368 202.014 32.472 206.388 ; 
        RECT 31.936 202.014 32.04 206.388 ; 
        RECT 31.504 202.014 31.608 206.388 ; 
        RECT 31.072 202.014 31.176 206.388 ; 
        RECT 30.64 202.014 30.744 206.388 ; 
        RECT 30.208 202.014 30.312 206.388 ; 
        RECT 29.776 202.014 29.88 206.388 ; 
        RECT 29.344 202.014 29.448 206.388 ; 
        RECT 28.912 202.014 29.016 206.388 ; 
        RECT 28.48 202.014 28.584 206.388 ; 
        RECT 28.048 202.014 28.152 206.388 ; 
        RECT 27.616 202.014 27.72 206.388 ; 
        RECT 27.184 202.014 27.288 206.388 ; 
        RECT 26.752 202.014 26.856 206.388 ; 
        RECT 26.32 202.014 26.424 206.388 ; 
        RECT 25.888 202.014 25.992 206.388 ; 
        RECT 25.456 202.014 25.56 206.388 ; 
        RECT 25.024 202.014 25.128 206.388 ; 
        RECT 24.592 202.014 24.696 206.388 ; 
        RECT 24.16 202.014 24.264 206.388 ; 
        RECT 23.728 202.014 23.832 206.388 ; 
        RECT 23.296 202.014 23.4 206.388 ; 
        RECT 22.864 202.014 22.968 206.388 ; 
        RECT 22.432 202.014 22.536 206.388 ; 
        RECT 22 202.014 22.104 206.388 ; 
        RECT 21.568 202.014 21.672 206.388 ; 
        RECT 21.136 202.014 21.24 206.388 ; 
        RECT 20.704 202.014 20.808 206.388 ; 
        RECT 20.272 202.014 20.376 206.388 ; 
        RECT 19.84 202.014 19.944 206.388 ; 
        RECT 19.408 202.014 19.512 206.388 ; 
        RECT 18.976 202.014 19.08 206.388 ; 
        RECT 18.544 202.014 18.648 206.388 ; 
        RECT 18.112 202.014 18.216 206.388 ; 
        RECT 17.68 202.014 17.784 206.388 ; 
        RECT 17.248 202.014 17.352 206.388 ; 
        RECT 16.816 202.014 16.92 206.388 ; 
        RECT 16.384 202.014 16.488 206.388 ; 
        RECT 15.952 202.014 16.056 206.388 ; 
        RECT 15.52 202.014 15.624 206.388 ; 
        RECT 15.088 202.014 15.192 206.388 ; 
        RECT 14.656 202.014 14.76 206.388 ; 
        RECT 14.224 202.014 14.328 206.388 ; 
        RECT 13.792 202.014 13.896 206.388 ; 
        RECT 13.36 202.014 13.464 206.388 ; 
        RECT 12.928 202.014 13.032 206.388 ; 
        RECT 12.496 202.014 12.6 206.388 ; 
        RECT 12.064 202.014 12.168 206.388 ; 
        RECT 11.632 202.014 11.736 206.388 ; 
        RECT 11.2 202.014 11.304 206.388 ; 
        RECT 10.768 202.014 10.872 206.388 ; 
        RECT 10.336 202.014 10.44 206.388 ; 
        RECT 9.904 202.014 10.008 206.388 ; 
        RECT 9.472 202.014 9.576 206.388 ; 
        RECT 9.04 202.014 9.144 206.388 ; 
        RECT 8.608 202.014 8.712 206.388 ; 
        RECT 8.176 202.014 8.28 206.388 ; 
        RECT 7.744 202.014 7.848 206.388 ; 
        RECT 7.312 202.014 7.416 206.388 ; 
        RECT 6.88 202.014 6.984 206.388 ; 
        RECT 6.448 202.014 6.552 206.388 ; 
        RECT 6.016 202.014 6.12 206.388 ; 
        RECT 5.584 202.014 5.688 206.388 ; 
        RECT 5.152 202.014 5.256 206.388 ; 
        RECT 4.72 202.014 4.824 206.388 ; 
        RECT 4.288 202.014 4.392 206.388 ; 
        RECT 3.856 202.014 3.96 206.388 ; 
        RECT 3.424 202.014 3.528 206.388 ; 
        RECT 2.992 202.014 3.096 206.388 ; 
        RECT 2.56 202.014 2.664 206.388 ; 
        RECT 2.128 202.014 2.232 206.388 ; 
        RECT 1.696 202.014 1.8 206.388 ; 
        RECT 1.264 202.014 1.368 206.388 ; 
        RECT 0.832 202.014 0.936 206.388 ; 
        RECT 0.02 202.014 0.36 206.388 ; 
        RECT 62.212 206.334 62.724 210.708 ; 
        RECT 62.156 208.996 62.724 210.286 ; 
        RECT 61.276 207.904 61.812 210.708 ; 
        RECT 61.184 209.244 61.812 210.276 ; 
        RECT 61.276 206.334 61.668 210.708 ; 
        RECT 61.276 206.818 61.724 207.776 ; 
        RECT 61.276 206.334 61.812 206.69 ; 
        RECT 60.376 208.136 60.912 210.708 ; 
        RECT 60.376 206.334 60.768 210.708 ; 
        RECT 58.708 206.334 59.04 210.708 ; 
        RECT 58.708 206.688 59.096 210.43 ; 
        RECT 121.072 206.334 121.412 210.708 ; 
        RECT 120.496 206.334 120.6 210.708 ; 
        RECT 120.064 206.334 120.168 210.708 ; 
        RECT 119.632 206.334 119.736 210.708 ; 
        RECT 119.2 206.334 119.304 210.708 ; 
        RECT 118.768 206.334 118.872 210.708 ; 
        RECT 118.336 206.334 118.44 210.708 ; 
        RECT 117.904 206.334 118.008 210.708 ; 
        RECT 117.472 206.334 117.576 210.708 ; 
        RECT 117.04 206.334 117.144 210.708 ; 
        RECT 116.608 206.334 116.712 210.708 ; 
        RECT 116.176 206.334 116.28 210.708 ; 
        RECT 115.744 206.334 115.848 210.708 ; 
        RECT 115.312 206.334 115.416 210.708 ; 
        RECT 114.88 206.334 114.984 210.708 ; 
        RECT 114.448 206.334 114.552 210.708 ; 
        RECT 114.016 206.334 114.12 210.708 ; 
        RECT 113.584 206.334 113.688 210.708 ; 
        RECT 113.152 206.334 113.256 210.708 ; 
        RECT 112.72 206.334 112.824 210.708 ; 
        RECT 112.288 206.334 112.392 210.708 ; 
        RECT 111.856 206.334 111.96 210.708 ; 
        RECT 111.424 206.334 111.528 210.708 ; 
        RECT 110.992 206.334 111.096 210.708 ; 
        RECT 110.56 206.334 110.664 210.708 ; 
        RECT 110.128 206.334 110.232 210.708 ; 
        RECT 109.696 206.334 109.8 210.708 ; 
        RECT 109.264 206.334 109.368 210.708 ; 
        RECT 108.832 206.334 108.936 210.708 ; 
        RECT 108.4 206.334 108.504 210.708 ; 
        RECT 107.968 206.334 108.072 210.708 ; 
        RECT 107.536 206.334 107.64 210.708 ; 
        RECT 107.104 206.334 107.208 210.708 ; 
        RECT 106.672 206.334 106.776 210.708 ; 
        RECT 106.24 206.334 106.344 210.708 ; 
        RECT 105.808 206.334 105.912 210.708 ; 
        RECT 105.376 206.334 105.48 210.708 ; 
        RECT 104.944 206.334 105.048 210.708 ; 
        RECT 104.512 206.334 104.616 210.708 ; 
        RECT 104.08 206.334 104.184 210.708 ; 
        RECT 103.648 206.334 103.752 210.708 ; 
        RECT 103.216 206.334 103.32 210.708 ; 
        RECT 102.784 206.334 102.888 210.708 ; 
        RECT 102.352 206.334 102.456 210.708 ; 
        RECT 101.92 206.334 102.024 210.708 ; 
        RECT 101.488 206.334 101.592 210.708 ; 
        RECT 101.056 206.334 101.16 210.708 ; 
        RECT 100.624 206.334 100.728 210.708 ; 
        RECT 100.192 206.334 100.296 210.708 ; 
        RECT 99.76 206.334 99.864 210.708 ; 
        RECT 99.328 206.334 99.432 210.708 ; 
        RECT 98.896 206.334 99 210.708 ; 
        RECT 98.464 206.334 98.568 210.708 ; 
        RECT 98.032 206.334 98.136 210.708 ; 
        RECT 97.6 206.334 97.704 210.708 ; 
        RECT 97.168 206.334 97.272 210.708 ; 
        RECT 96.736 206.334 96.84 210.708 ; 
        RECT 96.304 206.334 96.408 210.708 ; 
        RECT 95.872 206.334 95.976 210.708 ; 
        RECT 95.44 206.334 95.544 210.708 ; 
        RECT 95.008 206.334 95.112 210.708 ; 
        RECT 94.576 206.334 94.68 210.708 ; 
        RECT 94.144 206.334 94.248 210.708 ; 
        RECT 93.712 206.334 93.816 210.708 ; 
        RECT 93.28 206.334 93.384 210.708 ; 
        RECT 92.848 206.334 92.952 210.708 ; 
        RECT 92.416 206.334 92.52 210.708 ; 
        RECT 91.984 206.334 92.088 210.708 ; 
        RECT 91.552 206.334 91.656 210.708 ; 
        RECT 91.12 206.334 91.224 210.708 ; 
        RECT 90.688 206.334 90.792 210.708 ; 
        RECT 90.256 206.334 90.36 210.708 ; 
        RECT 89.824 206.334 89.928 210.708 ; 
        RECT 89.392 206.334 89.496 210.708 ; 
        RECT 88.96 206.334 89.064 210.708 ; 
        RECT 88.528 206.334 88.632 210.708 ; 
        RECT 88.096 206.334 88.2 210.708 ; 
        RECT 87.664 206.334 87.768 210.708 ; 
        RECT 87.232 206.334 87.336 210.708 ; 
        RECT 86.8 206.334 86.904 210.708 ; 
        RECT 86.368 206.334 86.472 210.708 ; 
        RECT 85.936 206.334 86.04 210.708 ; 
        RECT 85.504 206.334 85.608 210.708 ; 
        RECT 85.072 206.334 85.176 210.708 ; 
        RECT 84.64 206.334 84.744 210.708 ; 
        RECT 84.208 206.334 84.312 210.708 ; 
        RECT 83.776 206.334 83.88 210.708 ; 
        RECT 83.344 206.334 83.448 210.708 ; 
        RECT 82.912 206.334 83.016 210.708 ; 
        RECT 82.48 206.334 82.584 210.708 ; 
        RECT 82.048 206.334 82.152 210.708 ; 
        RECT 81.616 206.334 81.72 210.708 ; 
        RECT 81.184 206.334 81.288 210.708 ; 
        RECT 80.752 206.334 80.856 210.708 ; 
        RECT 80.32 206.334 80.424 210.708 ; 
        RECT 79.888 206.334 79.992 210.708 ; 
        RECT 79.456 206.334 79.56 210.708 ; 
        RECT 79.024 206.334 79.128 210.708 ; 
        RECT 78.592 206.334 78.696 210.708 ; 
        RECT 78.16 206.334 78.264 210.708 ; 
        RECT 77.728 206.334 77.832 210.708 ; 
        RECT 77.296 206.334 77.4 210.708 ; 
        RECT 76.864 206.334 76.968 210.708 ; 
        RECT 76.432 206.334 76.536 210.708 ; 
        RECT 76 206.334 76.104 210.708 ; 
        RECT 75.568 206.334 75.672 210.708 ; 
        RECT 75.136 206.334 75.24 210.708 ; 
        RECT 74.704 206.334 74.808 210.708 ; 
        RECT 74.272 206.334 74.376 210.708 ; 
        RECT 73.84 206.334 73.944 210.708 ; 
        RECT 73.408 206.334 73.512 210.708 ; 
        RECT 72.976 206.334 73.08 210.708 ; 
        RECT 72.544 206.334 72.648 210.708 ; 
        RECT 72.112 206.334 72.216 210.708 ; 
        RECT 71.68 206.334 71.784 210.708 ; 
        RECT 71.248 206.334 71.352 210.708 ; 
        RECT 70.816 206.334 70.92 210.708 ; 
        RECT 70.384 206.334 70.488 210.708 ; 
        RECT 69.952 206.334 70.056 210.708 ; 
        RECT 69.52 206.334 69.624 210.708 ; 
        RECT 69.088 206.334 69.192 210.708 ; 
        RECT 68.656 206.334 68.76 210.708 ; 
        RECT 68.224 206.334 68.328 210.708 ; 
        RECT 67.792 206.334 67.896 210.708 ; 
        RECT 67.36 206.334 67.464 210.708 ; 
        RECT 66.928 206.334 67.032 210.708 ; 
        RECT 66.496 206.334 66.6 210.708 ; 
        RECT 66.064 206.334 66.168 210.708 ; 
        RECT 65.632 206.334 65.736 210.708 ; 
        RECT 65.2 206.334 65.304 210.708 ; 
        RECT 64.348 206.334 64.656 210.708 ; 
        RECT 56.776 206.334 57.084 210.708 ; 
        RECT 56.128 206.334 56.232 210.708 ; 
        RECT 55.696 206.334 55.8 210.708 ; 
        RECT 55.264 206.334 55.368 210.708 ; 
        RECT 54.832 206.334 54.936 210.708 ; 
        RECT 54.4 206.334 54.504 210.708 ; 
        RECT 53.968 206.334 54.072 210.708 ; 
        RECT 53.536 206.334 53.64 210.708 ; 
        RECT 53.104 206.334 53.208 210.708 ; 
        RECT 52.672 206.334 52.776 210.708 ; 
        RECT 52.24 206.334 52.344 210.708 ; 
        RECT 51.808 206.334 51.912 210.708 ; 
        RECT 51.376 206.334 51.48 210.708 ; 
        RECT 50.944 206.334 51.048 210.708 ; 
        RECT 50.512 206.334 50.616 210.708 ; 
        RECT 50.08 206.334 50.184 210.708 ; 
        RECT 49.648 206.334 49.752 210.708 ; 
        RECT 49.216 206.334 49.32 210.708 ; 
        RECT 48.784 206.334 48.888 210.708 ; 
        RECT 48.352 206.334 48.456 210.708 ; 
        RECT 47.92 206.334 48.024 210.708 ; 
        RECT 47.488 206.334 47.592 210.708 ; 
        RECT 47.056 206.334 47.16 210.708 ; 
        RECT 46.624 206.334 46.728 210.708 ; 
        RECT 46.192 206.334 46.296 210.708 ; 
        RECT 45.76 206.334 45.864 210.708 ; 
        RECT 45.328 206.334 45.432 210.708 ; 
        RECT 44.896 206.334 45 210.708 ; 
        RECT 44.464 206.334 44.568 210.708 ; 
        RECT 44.032 206.334 44.136 210.708 ; 
        RECT 43.6 206.334 43.704 210.708 ; 
        RECT 43.168 206.334 43.272 210.708 ; 
        RECT 42.736 206.334 42.84 210.708 ; 
        RECT 42.304 206.334 42.408 210.708 ; 
        RECT 41.872 206.334 41.976 210.708 ; 
        RECT 41.44 206.334 41.544 210.708 ; 
        RECT 41.008 206.334 41.112 210.708 ; 
        RECT 40.576 206.334 40.68 210.708 ; 
        RECT 40.144 206.334 40.248 210.708 ; 
        RECT 39.712 206.334 39.816 210.708 ; 
        RECT 39.28 206.334 39.384 210.708 ; 
        RECT 38.848 206.334 38.952 210.708 ; 
        RECT 38.416 206.334 38.52 210.708 ; 
        RECT 37.984 206.334 38.088 210.708 ; 
        RECT 37.552 206.334 37.656 210.708 ; 
        RECT 37.12 206.334 37.224 210.708 ; 
        RECT 36.688 206.334 36.792 210.708 ; 
        RECT 36.256 206.334 36.36 210.708 ; 
        RECT 35.824 206.334 35.928 210.708 ; 
        RECT 35.392 206.334 35.496 210.708 ; 
        RECT 34.96 206.334 35.064 210.708 ; 
        RECT 34.528 206.334 34.632 210.708 ; 
        RECT 34.096 206.334 34.2 210.708 ; 
        RECT 33.664 206.334 33.768 210.708 ; 
        RECT 33.232 206.334 33.336 210.708 ; 
        RECT 32.8 206.334 32.904 210.708 ; 
        RECT 32.368 206.334 32.472 210.708 ; 
        RECT 31.936 206.334 32.04 210.708 ; 
        RECT 31.504 206.334 31.608 210.708 ; 
        RECT 31.072 206.334 31.176 210.708 ; 
        RECT 30.64 206.334 30.744 210.708 ; 
        RECT 30.208 206.334 30.312 210.708 ; 
        RECT 29.776 206.334 29.88 210.708 ; 
        RECT 29.344 206.334 29.448 210.708 ; 
        RECT 28.912 206.334 29.016 210.708 ; 
        RECT 28.48 206.334 28.584 210.708 ; 
        RECT 28.048 206.334 28.152 210.708 ; 
        RECT 27.616 206.334 27.72 210.708 ; 
        RECT 27.184 206.334 27.288 210.708 ; 
        RECT 26.752 206.334 26.856 210.708 ; 
        RECT 26.32 206.334 26.424 210.708 ; 
        RECT 25.888 206.334 25.992 210.708 ; 
        RECT 25.456 206.334 25.56 210.708 ; 
        RECT 25.024 206.334 25.128 210.708 ; 
        RECT 24.592 206.334 24.696 210.708 ; 
        RECT 24.16 206.334 24.264 210.708 ; 
        RECT 23.728 206.334 23.832 210.708 ; 
        RECT 23.296 206.334 23.4 210.708 ; 
        RECT 22.864 206.334 22.968 210.708 ; 
        RECT 22.432 206.334 22.536 210.708 ; 
        RECT 22 206.334 22.104 210.708 ; 
        RECT 21.568 206.334 21.672 210.708 ; 
        RECT 21.136 206.334 21.24 210.708 ; 
        RECT 20.704 206.334 20.808 210.708 ; 
        RECT 20.272 206.334 20.376 210.708 ; 
        RECT 19.84 206.334 19.944 210.708 ; 
        RECT 19.408 206.334 19.512 210.708 ; 
        RECT 18.976 206.334 19.08 210.708 ; 
        RECT 18.544 206.334 18.648 210.708 ; 
        RECT 18.112 206.334 18.216 210.708 ; 
        RECT 17.68 206.334 17.784 210.708 ; 
        RECT 17.248 206.334 17.352 210.708 ; 
        RECT 16.816 206.334 16.92 210.708 ; 
        RECT 16.384 206.334 16.488 210.708 ; 
        RECT 15.952 206.334 16.056 210.708 ; 
        RECT 15.52 206.334 15.624 210.708 ; 
        RECT 15.088 206.334 15.192 210.708 ; 
        RECT 14.656 206.334 14.76 210.708 ; 
        RECT 14.224 206.334 14.328 210.708 ; 
        RECT 13.792 206.334 13.896 210.708 ; 
        RECT 13.36 206.334 13.464 210.708 ; 
        RECT 12.928 206.334 13.032 210.708 ; 
        RECT 12.496 206.334 12.6 210.708 ; 
        RECT 12.064 206.334 12.168 210.708 ; 
        RECT 11.632 206.334 11.736 210.708 ; 
        RECT 11.2 206.334 11.304 210.708 ; 
        RECT 10.768 206.334 10.872 210.708 ; 
        RECT 10.336 206.334 10.44 210.708 ; 
        RECT 9.904 206.334 10.008 210.708 ; 
        RECT 9.472 206.334 9.576 210.708 ; 
        RECT 9.04 206.334 9.144 210.708 ; 
        RECT 8.608 206.334 8.712 210.708 ; 
        RECT 8.176 206.334 8.28 210.708 ; 
        RECT 7.744 206.334 7.848 210.708 ; 
        RECT 7.312 206.334 7.416 210.708 ; 
        RECT 6.88 206.334 6.984 210.708 ; 
        RECT 6.448 206.334 6.552 210.708 ; 
        RECT 6.016 206.334 6.12 210.708 ; 
        RECT 5.584 206.334 5.688 210.708 ; 
        RECT 5.152 206.334 5.256 210.708 ; 
        RECT 4.72 206.334 4.824 210.708 ; 
        RECT 4.288 206.334 4.392 210.708 ; 
        RECT 3.856 206.334 3.96 210.708 ; 
        RECT 3.424 206.334 3.528 210.708 ; 
        RECT 2.992 206.334 3.096 210.708 ; 
        RECT 2.56 206.334 2.664 210.708 ; 
        RECT 2.128 206.334 2.232 210.708 ; 
        RECT 1.696 206.334 1.8 210.708 ; 
        RECT 1.264 206.334 1.368 210.708 ; 
        RECT 0.832 206.334 0.936 210.708 ; 
        RECT 0.02 206.334 0.36 210.708 ; 
        RECT 62.212 210.654 62.724 215.028 ; 
        RECT 62.156 213.316 62.724 214.606 ; 
        RECT 61.276 212.224 61.812 215.028 ; 
        RECT 61.184 213.564 61.812 214.596 ; 
        RECT 61.276 210.654 61.668 215.028 ; 
        RECT 61.276 211.138 61.724 212.096 ; 
        RECT 61.276 210.654 61.812 211.01 ; 
        RECT 60.376 212.456 60.912 215.028 ; 
        RECT 60.376 210.654 60.768 215.028 ; 
        RECT 58.708 210.654 59.04 215.028 ; 
        RECT 58.708 211.008 59.096 214.75 ; 
        RECT 121.072 210.654 121.412 215.028 ; 
        RECT 120.496 210.654 120.6 215.028 ; 
        RECT 120.064 210.654 120.168 215.028 ; 
        RECT 119.632 210.654 119.736 215.028 ; 
        RECT 119.2 210.654 119.304 215.028 ; 
        RECT 118.768 210.654 118.872 215.028 ; 
        RECT 118.336 210.654 118.44 215.028 ; 
        RECT 117.904 210.654 118.008 215.028 ; 
        RECT 117.472 210.654 117.576 215.028 ; 
        RECT 117.04 210.654 117.144 215.028 ; 
        RECT 116.608 210.654 116.712 215.028 ; 
        RECT 116.176 210.654 116.28 215.028 ; 
        RECT 115.744 210.654 115.848 215.028 ; 
        RECT 115.312 210.654 115.416 215.028 ; 
        RECT 114.88 210.654 114.984 215.028 ; 
        RECT 114.448 210.654 114.552 215.028 ; 
        RECT 114.016 210.654 114.12 215.028 ; 
        RECT 113.584 210.654 113.688 215.028 ; 
        RECT 113.152 210.654 113.256 215.028 ; 
        RECT 112.72 210.654 112.824 215.028 ; 
        RECT 112.288 210.654 112.392 215.028 ; 
        RECT 111.856 210.654 111.96 215.028 ; 
        RECT 111.424 210.654 111.528 215.028 ; 
        RECT 110.992 210.654 111.096 215.028 ; 
        RECT 110.56 210.654 110.664 215.028 ; 
        RECT 110.128 210.654 110.232 215.028 ; 
        RECT 109.696 210.654 109.8 215.028 ; 
        RECT 109.264 210.654 109.368 215.028 ; 
        RECT 108.832 210.654 108.936 215.028 ; 
        RECT 108.4 210.654 108.504 215.028 ; 
        RECT 107.968 210.654 108.072 215.028 ; 
        RECT 107.536 210.654 107.64 215.028 ; 
        RECT 107.104 210.654 107.208 215.028 ; 
        RECT 106.672 210.654 106.776 215.028 ; 
        RECT 106.24 210.654 106.344 215.028 ; 
        RECT 105.808 210.654 105.912 215.028 ; 
        RECT 105.376 210.654 105.48 215.028 ; 
        RECT 104.944 210.654 105.048 215.028 ; 
        RECT 104.512 210.654 104.616 215.028 ; 
        RECT 104.08 210.654 104.184 215.028 ; 
        RECT 103.648 210.654 103.752 215.028 ; 
        RECT 103.216 210.654 103.32 215.028 ; 
        RECT 102.784 210.654 102.888 215.028 ; 
        RECT 102.352 210.654 102.456 215.028 ; 
        RECT 101.92 210.654 102.024 215.028 ; 
        RECT 101.488 210.654 101.592 215.028 ; 
        RECT 101.056 210.654 101.16 215.028 ; 
        RECT 100.624 210.654 100.728 215.028 ; 
        RECT 100.192 210.654 100.296 215.028 ; 
        RECT 99.76 210.654 99.864 215.028 ; 
        RECT 99.328 210.654 99.432 215.028 ; 
        RECT 98.896 210.654 99 215.028 ; 
        RECT 98.464 210.654 98.568 215.028 ; 
        RECT 98.032 210.654 98.136 215.028 ; 
        RECT 97.6 210.654 97.704 215.028 ; 
        RECT 97.168 210.654 97.272 215.028 ; 
        RECT 96.736 210.654 96.84 215.028 ; 
        RECT 96.304 210.654 96.408 215.028 ; 
        RECT 95.872 210.654 95.976 215.028 ; 
        RECT 95.44 210.654 95.544 215.028 ; 
        RECT 95.008 210.654 95.112 215.028 ; 
        RECT 94.576 210.654 94.68 215.028 ; 
        RECT 94.144 210.654 94.248 215.028 ; 
        RECT 93.712 210.654 93.816 215.028 ; 
        RECT 93.28 210.654 93.384 215.028 ; 
        RECT 92.848 210.654 92.952 215.028 ; 
        RECT 92.416 210.654 92.52 215.028 ; 
        RECT 91.984 210.654 92.088 215.028 ; 
        RECT 91.552 210.654 91.656 215.028 ; 
        RECT 91.12 210.654 91.224 215.028 ; 
        RECT 90.688 210.654 90.792 215.028 ; 
        RECT 90.256 210.654 90.36 215.028 ; 
        RECT 89.824 210.654 89.928 215.028 ; 
        RECT 89.392 210.654 89.496 215.028 ; 
        RECT 88.96 210.654 89.064 215.028 ; 
        RECT 88.528 210.654 88.632 215.028 ; 
        RECT 88.096 210.654 88.2 215.028 ; 
        RECT 87.664 210.654 87.768 215.028 ; 
        RECT 87.232 210.654 87.336 215.028 ; 
        RECT 86.8 210.654 86.904 215.028 ; 
        RECT 86.368 210.654 86.472 215.028 ; 
        RECT 85.936 210.654 86.04 215.028 ; 
        RECT 85.504 210.654 85.608 215.028 ; 
        RECT 85.072 210.654 85.176 215.028 ; 
        RECT 84.64 210.654 84.744 215.028 ; 
        RECT 84.208 210.654 84.312 215.028 ; 
        RECT 83.776 210.654 83.88 215.028 ; 
        RECT 83.344 210.654 83.448 215.028 ; 
        RECT 82.912 210.654 83.016 215.028 ; 
        RECT 82.48 210.654 82.584 215.028 ; 
        RECT 82.048 210.654 82.152 215.028 ; 
        RECT 81.616 210.654 81.72 215.028 ; 
        RECT 81.184 210.654 81.288 215.028 ; 
        RECT 80.752 210.654 80.856 215.028 ; 
        RECT 80.32 210.654 80.424 215.028 ; 
        RECT 79.888 210.654 79.992 215.028 ; 
        RECT 79.456 210.654 79.56 215.028 ; 
        RECT 79.024 210.654 79.128 215.028 ; 
        RECT 78.592 210.654 78.696 215.028 ; 
        RECT 78.16 210.654 78.264 215.028 ; 
        RECT 77.728 210.654 77.832 215.028 ; 
        RECT 77.296 210.654 77.4 215.028 ; 
        RECT 76.864 210.654 76.968 215.028 ; 
        RECT 76.432 210.654 76.536 215.028 ; 
        RECT 76 210.654 76.104 215.028 ; 
        RECT 75.568 210.654 75.672 215.028 ; 
        RECT 75.136 210.654 75.24 215.028 ; 
        RECT 74.704 210.654 74.808 215.028 ; 
        RECT 74.272 210.654 74.376 215.028 ; 
        RECT 73.84 210.654 73.944 215.028 ; 
        RECT 73.408 210.654 73.512 215.028 ; 
        RECT 72.976 210.654 73.08 215.028 ; 
        RECT 72.544 210.654 72.648 215.028 ; 
        RECT 72.112 210.654 72.216 215.028 ; 
        RECT 71.68 210.654 71.784 215.028 ; 
        RECT 71.248 210.654 71.352 215.028 ; 
        RECT 70.816 210.654 70.92 215.028 ; 
        RECT 70.384 210.654 70.488 215.028 ; 
        RECT 69.952 210.654 70.056 215.028 ; 
        RECT 69.52 210.654 69.624 215.028 ; 
        RECT 69.088 210.654 69.192 215.028 ; 
        RECT 68.656 210.654 68.76 215.028 ; 
        RECT 68.224 210.654 68.328 215.028 ; 
        RECT 67.792 210.654 67.896 215.028 ; 
        RECT 67.36 210.654 67.464 215.028 ; 
        RECT 66.928 210.654 67.032 215.028 ; 
        RECT 66.496 210.654 66.6 215.028 ; 
        RECT 66.064 210.654 66.168 215.028 ; 
        RECT 65.632 210.654 65.736 215.028 ; 
        RECT 65.2 210.654 65.304 215.028 ; 
        RECT 64.348 210.654 64.656 215.028 ; 
        RECT 56.776 210.654 57.084 215.028 ; 
        RECT 56.128 210.654 56.232 215.028 ; 
        RECT 55.696 210.654 55.8 215.028 ; 
        RECT 55.264 210.654 55.368 215.028 ; 
        RECT 54.832 210.654 54.936 215.028 ; 
        RECT 54.4 210.654 54.504 215.028 ; 
        RECT 53.968 210.654 54.072 215.028 ; 
        RECT 53.536 210.654 53.64 215.028 ; 
        RECT 53.104 210.654 53.208 215.028 ; 
        RECT 52.672 210.654 52.776 215.028 ; 
        RECT 52.24 210.654 52.344 215.028 ; 
        RECT 51.808 210.654 51.912 215.028 ; 
        RECT 51.376 210.654 51.48 215.028 ; 
        RECT 50.944 210.654 51.048 215.028 ; 
        RECT 50.512 210.654 50.616 215.028 ; 
        RECT 50.08 210.654 50.184 215.028 ; 
        RECT 49.648 210.654 49.752 215.028 ; 
        RECT 49.216 210.654 49.32 215.028 ; 
        RECT 48.784 210.654 48.888 215.028 ; 
        RECT 48.352 210.654 48.456 215.028 ; 
        RECT 47.92 210.654 48.024 215.028 ; 
        RECT 47.488 210.654 47.592 215.028 ; 
        RECT 47.056 210.654 47.16 215.028 ; 
        RECT 46.624 210.654 46.728 215.028 ; 
        RECT 46.192 210.654 46.296 215.028 ; 
        RECT 45.76 210.654 45.864 215.028 ; 
        RECT 45.328 210.654 45.432 215.028 ; 
        RECT 44.896 210.654 45 215.028 ; 
        RECT 44.464 210.654 44.568 215.028 ; 
        RECT 44.032 210.654 44.136 215.028 ; 
        RECT 43.6 210.654 43.704 215.028 ; 
        RECT 43.168 210.654 43.272 215.028 ; 
        RECT 42.736 210.654 42.84 215.028 ; 
        RECT 42.304 210.654 42.408 215.028 ; 
        RECT 41.872 210.654 41.976 215.028 ; 
        RECT 41.44 210.654 41.544 215.028 ; 
        RECT 41.008 210.654 41.112 215.028 ; 
        RECT 40.576 210.654 40.68 215.028 ; 
        RECT 40.144 210.654 40.248 215.028 ; 
        RECT 39.712 210.654 39.816 215.028 ; 
        RECT 39.28 210.654 39.384 215.028 ; 
        RECT 38.848 210.654 38.952 215.028 ; 
        RECT 38.416 210.654 38.52 215.028 ; 
        RECT 37.984 210.654 38.088 215.028 ; 
        RECT 37.552 210.654 37.656 215.028 ; 
        RECT 37.12 210.654 37.224 215.028 ; 
        RECT 36.688 210.654 36.792 215.028 ; 
        RECT 36.256 210.654 36.36 215.028 ; 
        RECT 35.824 210.654 35.928 215.028 ; 
        RECT 35.392 210.654 35.496 215.028 ; 
        RECT 34.96 210.654 35.064 215.028 ; 
        RECT 34.528 210.654 34.632 215.028 ; 
        RECT 34.096 210.654 34.2 215.028 ; 
        RECT 33.664 210.654 33.768 215.028 ; 
        RECT 33.232 210.654 33.336 215.028 ; 
        RECT 32.8 210.654 32.904 215.028 ; 
        RECT 32.368 210.654 32.472 215.028 ; 
        RECT 31.936 210.654 32.04 215.028 ; 
        RECT 31.504 210.654 31.608 215.028 ; 
        RECT 31.072 210.654 31.176 215.028 ; 
        RECT 30.64 210.654 30.744 215.028 ; 
        RECT 30.208 210.654 30.312 215.028 ; 
        RECT 29.776 210.654 29.88 215.028 ; 
        RECT 29.344 210.654 29.448 215.028 ; 
        RECT 28.912 210.654 29.016 215.028 ; 
        RECT 28.48 210.654 28.584 215.028 ; 
        RECT 28.048 210.654 28.152 215.028 ; 
        RECT 27.616 210.654 27.72 215.028 ; 
        RECT 27.184 210.654 27.288 215.028 ; 
        RECT 26.752 210.654 26.856 215.028 ; 
        RECT 26.32 210.654 26.424 215.028 ; 
        RECT 25.888 210.654 25.992 215.028 ; 
        RECT 25.456 210.654 25.56 215.028 ; 
        RECT 25.024 210.654 25.128 215.028 ; 
        RECT 24.592 210.654 24.696 215.028 ; 
        RECT 24.16 210.654 24.264 215.028 ; 
        RECT 23.728 210.654 23.832 215.028 ; 
        RECT 23.296 210.654 23.4 215.028 ; 
        RECT 22.864 210.654 22.968 215.028 ; 
        RECT 22.432 210.654 22.536 215.028 ; 
        RECT 22 210.654 22.104 215.028 ; 
        RECT 21.568 210.654 21.672 215.028 ; 
        RECT 21.136 210.654 21.24 215.028 ; 
        RECT 20.704 210.654 20.808 215.028 ; 
        RECT 20.272 210.654 20.376 215.028 ; 
        RECT 19.84 210.654 19.944 215.028 ; 
        RECT 19.408 210.654 19.512 215.028 ; 
        RECT 18.976 210.654 19.08 215.028 ; 
        RECT 18.544 210.654 18.648 215.028 ; 
        RECT 18.112 210.654 18.216 215.028 ; 
        RECT 17.68 210.654 17.784 215.028 ; 
        RECT 17.248 210.654 17.352 215.028 ; 
        RECT 16.816 210.654 16.92 215.028 ; 
        RECT 16.384 210.654 16.488 215.028 ; 
        RECT 15.952 210.654 16.056 215.028 ; 
        RECT 15.52 210.654 15.624 215.028 ; 
        RECT 15.088 210.654 15.192 215.028 ; 
        RECT 14.656 210.654 14.76 215.028 ; 
        RECT 14.224 210.654 14.328 215.028 ; 
        RECT 13.792 210.654 13.896 215.028 ; 
        RECT 13.36 210.654 13.464 215.028 ; 
        RECT 12.928 210.654 13.032 215.028 ; 
        RECT 12.496 210.654 12.6 215.028 ; 
        RECT 12.064 210.654 12.168 215.028 ; 
        RECT 11.632 210.654 11.736 215.028 ; 
        RECT 11.2 210.654 11.304 215.028 ; 
        RECT 10.768 210.654 10.872 215.028 ; 
        RECT 10.336 210.654 10.44 215.028 ; 
        RECT 9.904 210.654 10.008 215.028 ; 
        RECT 9.472 210.654 9.576 215.028 ; 
        RECT 9.04 210.654 9.144 215.028 ; 
        RECT 8.608 210.654 8.712 215.028 ; 
        RECT 8.176 210.654 8.28 215.028 ; 
        RECT 7.744 210.654 7.848 215.028 ; 
        RECT 7.312 210.654 7.416 215.028 ; 
        RECT 6.88 210.654 6.984 215.028 ; 
        RECT 6.448 210.654 6.552 215.028 ; 
        RECT 6.016 210.654 6.12 215.028 ; 
        RECT 5.584 210.654 5.688 215.028 ; 
        RECT 5.152 210.654 5.256 215.028 ; 
        RECT 4.72 210.654 4.824 215.028 ; 
        RECT 4.288 210.654 4.392 215.028 ; 
        RECT 3.856 210.654 3.96 215.028 ; 
        RECT 3.424 210.654 3.528 215.028 ; 
        RECT 2.992 210.654 3.096 215.028 ; 
        RECT 2.56 210.654 2.664 215.028 ; 
        RECT 2.128 210.654 2.232 215.028 ; 
        RECT 1.696 210.654 1.8 215.028 ; 
        RECT 1.264 210.654 1.368 215.028 ; 
        RECT 0.832 210.654 0.936 215.028 ; 
        RECT 0.02 210.654 0.36 215.028 ; 
        RECT 62.212 214.974 62.724 219.348 ; 
        RECT 62.156 217.636 62.724 218.926 ; 
        RECT 61.276 216.544 61.812 219.348 ; 
        RECT 61.184 217.884 61.812 218.916 ; 
        RECT 61.276 214.974 61.668 219.348 ; 
        RECT 61.276 215.458 61.724 216.416 ; 
        RECT 61.276 214.974 61.812 215.33 ; 
        RECT 60.376 216.776 60.912 219.348 ; 
        RECT 60.376 214.974 60.768 219.348 ; 
        RECT 58.708 214.974 59.04 219.348 ; 
        RECT 58.708 215.328 59.096 219.07 ; 
        RECT 121.072 214.974 121.412 219.348 ; 
        RECT 120.496 214.974 120.6 219.348 ; 
        RECT 120.064 214.974 120.168 219.348 ; 
        RECT 119.632 214.974 119.736 219.348 ; 
        RECT 119.2 214.974 119.304 219.348 ; 
        RECT 118.768 214.974 118.872 219.348 ; 
        RECT 118.336 214.974 118.44 219.348 ; 
        RECT 117.904 214.974 118.008 219.348 ; 
        RECT 117.472 214.974 117.576 219.348 ; 
        RECT 117.04 214.974 117.144 219.348 ; 
        RECT 116.608 214.974 116.712 219.348 ; 
        RECT 116.176 214.974 116.28 219.348 ; 
        RECT 115.744 214.974 115.848 219.348 ; 
        RECT 115.312 214.974 115.416 219.348 ; 
        RECT 114.88 214.974 114.984 219.348 ; 
        RECT 114.448 214.974 114.552 219.348 ; 
        RECT 114.016 214.974 114.12 219.348 ; 
        RECT 113.584 214.974 113.688 219.348 ; 
        RECT 113.152 214.974 113.256 219.348 ; 
        RECT 112.72 214.974 112.824 219.348 ; 
        RECT 112.288 214.974 112.392 219.348 ; 
        RECT 111.856 214.974 111.96 219.348 ; 
        RECT 111.424 214.974 111.528 219.348 ; 
        RECT 110.992 214.974 111.096 219.348 ; 
        RECT 110.56 214.974 110.664 219.348 ; 
        RECT 110.128 214.974 110.232 219.348 ; 
        RECT 109.696 214.974 109.8 219.348 ; 
        RECT 109.264 214.974 109.368 219.348 ; 
        RECT 108.832 214.974 108.936 219.348 ; 
        RECT 108.4 214.974 108.504 219.348 ; 
        RECT 107.968 214.974 108.072 219.348 ; 
        RECT 107.536 214.974 107.64 219.348 ; 
        RECT 107.104 214.974 107.208 219.348 ; 
        RECT 106.672 214.974 106.776 219.348 ; 
        RECT 106.24 214.974 106.344 219.348 ; 
        RECT 105.808 214.974 105.912 219.348 ; 
        RECT 105.376 214.974 105.48 219.348 ; 
        RECT 104.944 214.974 105.048 219.348 ; 
        RECT 104.512 214.974 104.616 219.348 ; 
        RECT 104.08 214.974 104.184 219.348 ; 
        RECT 103.648 214.974 103.752 219.348 ; 
        RECT 103.216 214.974 103.32 219.348 ; 
        RECT 102.784 214.974 102.888 219.348 ; 
        RECT 102.352 214.974 102.456 219.348 ; 
        RECT 101.92 214.974 102.024 219.348 ; 
        RECT 101.488 214.974 101.592 219.348 ; 
        RECT 101.056 214.974 101.16 219.348 ; 
        RECT 100.624 214.974 100.728 219.348 ; 
        RECT 100.192 214.974 100.296 219.348 ; 
        RECT 99.76 214.974 99.864 219.348 ; 
        RECT 99.328 214.974 99.432 219.348 ; 
        RECT 98.896 214.974 99 219.348 ; 
        RECT 98.464 214.974 98.568 219.348 ; 
        RECT 98.032 214.974 98.136 219.348 ; 
        RECT 97.6 214.974 97.704 219.348 ; 
        RECT 97.168 214.974 97.272 219.348 ; 
        RECT 96.736 214.974 96.84 219.348 ; 
        RECT 96.304 214.974 96.408 219.348 ; 
        RECT 95.872 214.974 95.976 219.348 ; 
        RECT 95.44 214.974 95.544 219.348 ; 
        RECT 95.008 214.974 95.112 219.348 ; 
        RECT 94.576 214.974 94.68 219.348 ; 
        RECT 94.144 214.974 94.248 219.348 ; 
        RECT 93.712 214.974 93.816 219.348 ; 
        RECT 93.28 214.974 93.384 219.348 ; 
        RECT 92.848 214.974 92.952 219.348 ; 
        RECT 92.416 214.974 92.52 219.348 ; 
        RECT 91.984 214.974 92.088 219.348 ; 
        RECT 91.552 214.974 91.656 219.348 ; 
        RECT 91.12 214.974 91.224 219.348 ; 
        RECT 90.688 214.974 90.792 219.348 ; 
        RECT 90.256 214.974 90.36 219.348 ; 
        RECT 89.824 214.974 89.928 219.348 ; 
        RECT 89.392 214.974 89.496 219.348 ; 
        RECT 88.96 214.974 89.064 219.348 ; 
        RECT 88.528 214.974 88.632 219.348 ; 
        RECT 88.096 214.974 88.2 219.348 ; 
        RECT 87.664 214.974 87.768 219.348 ; 
        RECT 87.232 214.974 87.336 219.348 ; 
        RECT 86.8 214.974 86.904 219.348 ; 
        RECT 86.368 214.974 86.472 219.348 ; 
        RECT 85.936 214.974 86.04 219.348 ; 
        RECT 85.504 214.974 85.608 219.348 ; 
        RECT 85.072 214.974 85.176 219.348 ; 
        RECT 84.64 214.974 84.744 219.348 ; 
        RECT 84.208 214.974 84.312 219.348 ; 
        RECT 83.776 214.974 83.88 219.348 ; 
        RECT 83.344 214.974 83.448 219.348 ; 
        RECT 82.912 214.974 83.016 219.348 ; 
        RECT 82.48 214.974 82.584 219.348 ; 
        RECT 82.048 214.974 82.152 219.348 ; 
        RECT 81.616 214.974 81.72 219.348 ; 
        RECT 81.184 214.974 81.288 219.348 ; 
        RECT 80.752 214.974 80.856 219.348 ; 
        RECT 80.32 214.974 80.424 219.348 ; 
        RECT 79.888 214.974 79.992 219.348 ; 
        RECT 79.456 214.974 79.56 219.348 ; 
        RECT 79.024 214.974 79.128 219.348 ; 
        RECT 78.592 214.974 78.696 219.348 ; 
        RECT 78.16 214.974 78.264 219.348 ; 
        RECT 77.728 214.974 77.832 219.348 ; 
        RECT 77.296 214.974 77.4 219.348 ; 
        RECT 76.864 214.974 76.968 219.348 ; 
        RECT 76.432 214.974 76.536 219.348 ; 
        RECT 76 214.974 76.104 219.348 ; 
        RECT 75.568 214.974 75.672 219.348 ; 
        RECT 75.136 214.974 75.24 219.348 ; 
        RECT 74.704 214.974 74.808 219.348 ; 
        RECT 74.272 214.974 74.376 219.348 ; 
        RECT 73.84 214.974 73.944 219.348 ; 
        RECT 73.408 214.974 73.512 219.348 ; 
        RECT 72.976 214.974 73.08 219.348 ; 
        RECT 72.544 214.974 72.648 219.348 ; 
        RECT 72.112 214.974 72.216 219.348 ; 
        RECT 71.68 214.974 71.784 219.348 ; 
        RECT 71.248 214.974 71.352 219.348 ; 
        RECT 70.816 214.974 70.92 219.348 ; 
        RECT 70.384 214.974 70.488 219.348 ; 
        RECT 69.952 214.974 70.056 219.348 ; 
        RECT 69.52 214.974 69.624 219.348 ; 
        RECT 69.088 214.974 69.192 219.348 ; 
        RECT 68.656 214.974 68.76 219.348 ; 
        RECT 68.224 214.974 68.328 219.348 ; 
        RECT 67.792 214.974 67.896 219.348 ; 
        RECT 67.36 214.974 67.464 219.348 ; 
        RECT 66.928 214.974 67.032 219.348 ; 
        RECT 66.496 214.974 66.6 219.348 ; 
        RECT 66.064 214.974 66.168 219.348 ; 
        RECT 65.632 214.974 65.736 219.348 ; 
        RECT 65.2 214.974 65.304 219.348 ; 
        RECT 64.348 214.974 64.656 219.348 ; 
        RECT 56.776 214.974 57.084 219.348 ; 
        RECT 56.128 214.974 56.232 219.348 ; 
        RECT 55.696 214.974 55.8 219.348 ; 
        RECT 55.264 214.974 55.368 219.348 ; 
        RECT 54.832 214.974 54.936 219.348 ; 
        RECT 54.4 214.974 54.504 219.348 ; 
        RECT 53.968 214.974 54.072 219.348 ; 
        RECT 53.536 214.974 53.64 219.348 ; 
        RECT 53.104 214.974 53.208 219.348 ; 
        RECT 52.672 214.974 52.776 219.348 ; 
        RECT 52.24 214.974 52.344 219.348 ; 
        RECT 51.808 214.974 51.912 219.348 ; 
        RECT 51.376 214.974 51.48 219.348 ; 
        RECT 50.944 214.974 51.048 219.348 ; 
        RECT 50.512 214.974 50.616 219.348 ; 
        RECT 50.08 214.974 50.184 219.348 ; 
        RECT 49.648 214.974 49.752 219.348 ; 
        RECT 49.216 214.974 49.32 219.348 ; 
        RECT 48.784 214.974 48.888 219.348 ; 
        RECT 48.352 214.974 48.456 219.348 ; 
        RECT 47.92 214.974 48.024 219.348 ; 
        RECT 47.488 214.974 47.592 219.348 ; 
        RECT 47.056 214.974 47.16 219.348 ; 
        RECT 46.624 214.974 46.728 219.348 ; 
        RECT 46.192 214.974 46.296 219.348 ; 
        RECT 45.76 214.974 45.864 219.348 ; 
        RECT 45.328 214.974 45.432 219.348 ; 
        RECT 44.896 214.974 45 219.348 ; 
        RECT 44.464 214.974 44.568 219.348 ; 
        RECT 44.032 214.974 44.136 219.348 ; 
        RECT 43.6 214.974 43.704 219.348 ; 
        RECT 43.168 214.974 43.272 219.348 ; 
        RECT 42.736 214.974 42.84 219.348 ; 
        RECT 42.304 214.974 42.408 219.348 ; 
        RECT 41.872 214.974 41.976 219.348 ; 
        RECT 41.44 214.974 41.544 219.348 ; 
        RECT 41.008 214.974 41.112 219.348 ; 
        RECT 40.576 214.974 40.68 219.348 ; 
        RECT 40.144 214.974 40.248 219.348 ; 
        RECT 39.712 214.974 39.816 219.348 ; 
        RECT 39.28 214.974 39.384 219.348 ; 
        RECT 38.848 214.974 38.952 219.348 ; 
        RECT 38.416 214.974 38.52 219.348 ; 
        RECT 37.984 214.974 38.088 219.348 ; 
        RECT 37.552 214.974 37.656 219.348 ; 
        RECT 37.12 214.974 37.224 219.348 ; 
        RECT 36.688 214.974 36.792 219.348 ; 
        RECT 36.256 214.974 36.36 219.348 ; 
        RECT 35.824 214.974 35.928 219.348 ; 
        RECT 35.392 214.974 35.496 219.348 ; 
        RECT 34.96 214.974 35.064 219.348 ; 
        RECT 34.528 214.974 34.632 219.348 ; 
        RECT 34.096 214.974 34.2 219.348 ; 
        RECT 33.664 214.974 33.768 219.348 ; 
        RECT 33.232 214.974 33.336 219.348 ; 
        RECT 32.8 214.974 32.904 219.348 ; 
        RECT 32.368 214.974 32.472 219.348 ; 
        RECT 31.936 214.974 32.04 219.348 ; 
        RECT 31.504 214.974 31.608 219.348 ; 
        RECT 31.072 214.974 31.176 219.348 ; 
        RECT 30.64 214.974 30.744 219.348 ; 
        RECT 30.208 214.974 30.312 219.348 ; 
        RECT 29.776 214.974 29.88 219.348 ; 
        RECT 29.344 214.974 29.448 219.348 ; 
        RECT 28.912 214.974 29.016 219.348 ; 
        RECT 28.48 214.974 28.584 219.348 ; 
        RECT 28.048 214.974 28.152 219.348 ; 
        RECT 27.616 214.974 27.72 219.348 ; 
        RECT 27.184 214.974 27.288 219.348 ; 
        RECT 26.752 214.974 26.856 219.348 ; 
        RECT 26.32 214.974 26.424 219.348 ; 
        RECT 25.888 214.974 25.992 219.348 ; 
        RECT 25.456 214.974 25.56 219.348 ; 
        RECT 25.024 214.974 25.128 219.348 ; 
        RECT 24.592 214.974 24.696 219.348 ; 
        RECT 24.16 214.974 24.264 219.348 ; 
        RECT 23.728 214.974 23.832 219.348 ; 
        RECT 23.296 214.974 23.4 219.348 ; 
        RECT 22.864 214.974 22.968 219.348 ; 
        RECT 22.432 214.974 22.536 219.348 ; 
        RECT 22 214.974 22.104 219.348 ; 
        RECT 21.568 214.974 21.672 219.348 ; 
        RECT 21.136 214.974 21.24 219.348 ; 
        RECT 20.704 214.974 20.808 219.348 ; 
        RECT 20.272 214.974 20.376 219.348 ; 
        RECT 19.84 214.974 19.944 219.348 ; 
        RECT 19.408 214.974 19.512 219.348 ; 
        RECT 18.976 214.974 19.08 219.348 ; 
        RECT 18.544 214.974 18.648 219.348 ; 
        RECT 18.112 214.974 18.216 219.348 ; 
        RECT 17.68 214.974 17.784 219.348 ; 
        RECT 17.248 214.974 17.352 219.348 ; 
        RECT 16.816 214.974 16.92 219.348 ; 
        RECT 16.384 214.974 16.488 219.348 ; 
        RECT 15.952 214.974 16.056 219.348 ; 
        RECT 15.52 214.974 15.624 219.348 ; 
        RECT 15.088 214.974 15.192 219.348 ; 
        RECT 14.656 214.974 14.76 219.348 ; 
        RECT 14.224 214.974 14.328 219.348 ; 
        RECT 13.792 214.974 13.896 219.348 ; 
        RECT 13.36 214.974 13.464 219.348 ; 
        RECT 12.928 214.974 13.032 219.348 ; 
        RECT 12.496 214.974 12.6 219.348 ; 
        RECT 12.064 214.974 12.168 219.348 ; 
        RECT 11.632 214.974 11.736 219.348 ; 
        RECT 11.2 214.974 11.304 219.348 ; 
        RECT 10.768 214.974 10.872 219.348 ; 
        RECT 10.336 214.974 10.44 219.348 ; 
        RECT 9.904 214.974 10.008 219.348 ; 
        RECT 9.472 214.974 9.576 219.348 ; 
        RECT 9.04 214.974 9.144 219.348 ; 
        RECT 8.608 214.974 8.712 219.348 ; 
        RECT 8.176 214.974 8.28 219.348 ; 
        RECT 7.744 214.974 7.848 219.348 ; 
        RECT 7.312 214.974 7.416 219.348 ; 
        RECT 6.88 214.974 6.984 219.348 ; 
        RECT 6.448 214.974 6.552 219.348 ; 
        RECT 6.016 214.974 6.12 219.348 ; 
        RECT 5.584 214.974 5.688 219.348 ; 
        RECT 5.152 214.974 5.256 219.348 ; 
        RECT 4.72 214.974 4.824 219.348 ; 
        RECT 4.288 214.974 4.392 219.348 ; 
        RECT 3.856 214.974 3.96 219.348 ; 
        RECT 3.424 214.974 3.528 219.348 ; 
        RECT 2.992 214.974 3.096 219.348 ; 
        RECT 2.56 214.974 2.664 219.348 ; 
        RECT 2.128 214.974 2.232 219.348 ; 
        RECT 1.696 214.974 1.8 219.348 ; 
        RECT 1.264 214.974 1.368 219.348 ; 
        RECT 0.832 214.974 0.936 219.348 ; 
        RECT 0.02 214.974 0.36 219.348 ; 
        RECT 62.212 219.294 62.724 223.668 ; 
        RECT 62.156 221.956 62.724 223.246 ; 
        RECT 61.276 220.864 61.812 223.668 ; 
        RECT 61.184 222.204 61.812 223.236 ; 
        RECT 61.276 219.294 61.668 223.668 ; 
        RECT 61.276 219.778 61.724 220.736 ; 
        RECT 61.276 219.294 61.812 219.65 ; 
        RECT 60.376 221.096 60.912 223.668 ; 
        RECT 60.376 219.294 60.768 223.668 ; 
        RECT 58.708 219.294 59.04 223.668 ; 
        RECT 58.708 219.648 59.096 223.39 ; 
        RECT 121.072 219.294 121.412 223.668 ; 
        RECT 120.496 219.294 120.6 223.668 ; 
        RECT 120.064 219.294 120.168 223.668 ; 
        RECT 119.632 219.294 119.736 223.668 ; 
        RECT 119.2 219.294 119.304 223.668 ; 
        RECT 118.768 219.294 118.872 223.668 ; 
        RECT 118.336 219.294 118.44 223.668 ; 
        RECT 117.904 219.294 118.008 223.668 ; 
        RECT 117.472 219.294 117.576 223.668 ; 
        RECT 117.04 219.294 117.144 223.668 ; 
        RECT 116.608 219.294 116.712 223.668 ; 
        RECT 116.176 219.294 116.28 223.668 ; 
        RECT 115.744 219.294 115.848 223.668 ; 
        RECT 115.312 219.294 115.416 223.668 ; 
        RECT 114.88 219.294 114.984 223.668 ; 
        RECT 114.448 219.294 114.552 223.668 ; 
        RECT 114.016 219.294 114.12 223.668 ; 
        RECT 113.584 219.294 113.688 223.668 ; 
        RECT 113.152 219.294 113.256 223.668 ; 
        RECT 112.72 219.294 112.824 223.668 ; 
        RECT 112.288 219.294 112.392 223.668 ; 
        RECT 111.856 219.294 111.96 223.668 ; 
        RECT 111.424 219.294 111.528 223.668 ; 
        RECT 110.992 219.294 111.096 223.668 ; 
        RECT 110.56 219.294 110.664 223.668 ; 
        RECT 110.128 219.294 110.232 223.668 ; 
        RECT 109.696 219.294 109.8 223.668 ; 
        RECT 109.264 219.294 109.368 223.668 ; 
        RECT 108.832 219.294 108.936 223.668 ; 
        RECT 108.4 219.294 108.504 223.668 ; 
        RECT 107.968 219.294 108.072 223.668 ; 
        RECT 107.536 219.294 107.64 223.668 ; 
        RECT 107.104 219.294 107.208 223.668 ; 
        RECT 106.672 219.294 106.776 223.668 ; 
        RECT 106.24 219.294 106.344 223.668 ; 
        RECT 105.808 219.294 105.912 223.668 ; 
        RECT 105.376 219.294 105.48 223.668 ; 
        RECT 104.944 219.294 105.048 223.668 ; 
        RECT 104.512 219.294 104.616 223.668 ; 
        RECT 104.08 219.294 104.184 223.668 ; 
        RECT 103.648 219.294 103.752 223.668 ; 
        RECT 103.216 219.294 103.32 223.668 ; 
        RECT 102.784 219.294 102.888 223.668 ; 
        RECT 102.352 219.294 102.456 223.668 ; 
        RECT 101.92 219.294 102.024 223.668 ; 
        RECT 101.488 219.294 101.592 223.668 ; 
        RECT 101.056 219.294 101.16 223.668 ; 
        RECT 100.624 219.294 100.728 223.668 ; 
        RECT 100.192 219.294 100.296 223.668 ; 
        RECT 99.76 219.294 99.864 223.668 ; 
        RECT 99.328 219.294 99.432 223.668 ; 
        RECT 98.896 219.294 99 223.668 ; 
        RECT 98.464 219.294 98.568 223.668 ; 
        RECT 98.032 219.294 98.136 223.668 ; 
        RECT 97.6 219.294 97.704 223.668 ; 
        RECT 97.168 219.294 97.272 223.668 ; 
        RECT 96.736 219.294 96.84 223.668 ; 
        RECT 96.304 219.294 96.408 223.668 ; 
        RECT 95.872 219.294 95.976 223.668 ; 
        RECT 95.44 219.294 95.544 223.668 ; 
        RECT 95.008 219.294 95.112 223.668 ; 
        RECT 94.576 219.294 94.68 223.668 ; 
        RECT 94.144 219.294 94.248 223.668 ; 
        RECT 93.712 219.294 93.816 223.668 ; 
        RECT 93.28 219.294 93.384 223.668 ; 
        RECT 92.848 219.294 92.952 223.668 ; 
        RECT 92.416 219.294 92.52 223.668 ; 
        RECT 91.984 219.294 92.088 223.668 ; 
        RECT 91.552 219.294 91.656 223.668 ; 
        RECT 91.12 219.294 91.224 223.668 ; 
        RECT 90.688 219.294 90.792 223.668 ; 
        RECT 90.256 219.294 90.36 223.668 ; 
        RECT 89.824 219.294 89.928 223.668 ; 
        RECT 89.392 219.294 89.496 223.668 ; 
        RECT 88.96 219.294 89.064 223.668 ; 
        RECT 88.528 219.294 88.632 223.668 ; 
        RECT 88.096 219.294 88.2 223.668 ; 
        RECT 87.664 219.294 87.768 223.668 ; 
        RECT 87.232 219.294 87.336 223.668 ; 
        RECT 86.8 219.294 86.904 223.668 ; 
        RECT 86.368 219.294 86.472 223.668 ; 
        RECT 85.936 219.294 86.04 223.668 ; 
        RECT 85.504 219.294 85.608 223.668 ; 
        RECT 85.072 219.294 85.176 223.668 ; 
        RECT 84.64 219.294 84.744 223.668 ; 
        RECT 84.208 219.294 84.312 223.668 ; 
        RECT 83.776 219.294 83.88 223.668 ; 
        RECT 83.344 219.294 83.448 223.668 ; 
        RECT 82.912 219.294 83.016 223.668 ; 
        RECT 82.48 219.294 82.584 223.668 ; 
        RECT 82.048 219.294 82.152 223.668 ; 
        RECT 81.616 219.294 81.72 223.668 ; 
        RECT 81.184 219.294 81.288 223.668 ; 
        RECT 80.752 219.294 80.856 223.668 ; 
        RECT 80.32 219.294 80.424 223.668 ; 
        RECT 79.888 219.294 79.992 223.668 ; 
        RECT 79.456 219.294 79.56 223.668 ; 
        RECT 79.024 219.294 79.128 223.668 ; 
        RECT 78.592 219.294 78.696 223.668 ; 
        RECT 78.16 219.294 78.264 223.668 ; 
        RECT 77.728 219.294 77.832 223.668 ; 
        RECT 77.296 219.294 77.4 223.668 ; 
        RECT 76.864 219.294 76.968 223.668 ; 
        RECT 76.432 219.294 76.536 223.668 ; 
        RECT 76 219.294 76.104 223.668 ; 
        RECT 75.568 219.294 75.672 223.668 ; 
        RECT 75.136 219.294 75.24 223.668 ; 
        RECT 74.704 219.294 74.808 223.668 ; 
        RECT 74.272 219.294 74.376 223.668 ; 
        RECT 73.84 219.294 73.944 223.668 ; 
        RECT 73.408 219.294 73.512 223.668 ; 
        RECT 72.976 219.294 73.08 223.668 ; 
        RECT 72.544 219.294 72.648 223.668 ; 
        RECT 72.112 219.294 72.216 223.668 ; 
        RECT 71.68 219.294 71.784 223.668 ; 
        RECT 71.248 219.294 71.352 223.668 ; 
        RECT 70.816 219.294 70.92 223.668 ; 
        RECT 70.384 219.294 70.488 223.668 ; 
        RECT 69.952 219.294 70.056 223.668 ; 
        RECT 69.52 219.294 69.624 223.668 ; 
        RECT 69.088 219.294 69.192 223.668 ; 
        RECT 68.656 219.294 68.76 223.668 ; 
        RECT 68.224 219.294 68.328 223.668 ; 
        RECT 67.792 219.294 67.896 223.668 ; 
        RECT 67.36 219.294 67.464 223.668 ; 
        RECT 66.928 219.294 67.032 223.668 ; 
        RECT 66.496 219.294 66.6 223.668 ; 
        RECT 66.064 219.294 66.168 223.668 ; 
        RECT 65.632 219.294 65.736 223.668 ; 
        RECT 65.2 219.294 65.304 223.668 ; 
        RECT 64.348 219.294 64.656 223.668 ; 
        RECT 56.776 219.294 57.084 223.668 ; 
        RECT 56.128 219.294 56.232 223.668 ; 
        RECT 55.696 219.294 55.8 223.668 ; 
        RECT 55.264 219.294 55.368 223.668 ; 
        RECT 54.832 219.294 54.936 223.668 ; 
        RECT 54.4 219.294 54.504 223.668 ; 
        RECT 53.968 219.294 54.072 223.668 ; 
        RECT 53.536 219.294 53.64 223.668 ; 
        RECT 53.104 219.294 53.208 223.668 ; 
        RECT 52.672 219.294 52.776 223.668 ; 
        RECT 52.24 219.294 52.344 223.668 ; 
        RECT 51.808 219.294 51.912 223.668 ; 
        RECT 51.376 219.294 51.48 223.668 ; 
        RECT 50.944 219.294 51.048 223.668 ; 
        RECT 50.512 219.294 50.616 223.668 ; 
        RECT 50.08 219.294 50.184 223.668 ; 
        RECT 49.648 219.294 49.752 223.668 ; 
        RECT 49.216 219.294 49.32 223.668 ; 
        RECT 48.784 219.294 48.888 223.668 ; 
        RECT 48.352 219.294 48.456 223.668 ; 
        RECT 47.92 219.294 48.024 223.668 ; 
        RECT 47.488 219.294 47.592 223.668 ; 
        RECT 47.056 219.294 47.16 223.668 ; 
        RECT 46.624 219.294 46.728 223.668 ; 
        RECT 46.192 219.294 46.296 223.668 ; 
        RECT 45.76 219.294 45.864 223.668 ; 
        RECT 45.328 219.294 45.432 223.668 ; 
        RECT 44.896 219.294 45 223.668 ; 
        RECT 44.464 219.294 44.568 223.668 ; 
        RECT 44.032 219.294 44.136 223.668 ; 
        RECT 43.6 219.294 43.704 223.668 ; 
        RECT 43.168 219.294 43.272 223.668 ; 
        RECT 42.736 219.294 42.84 223.668 ; 
        RECT 42.304 219.294 42.408 223.668 ; 
        RECT 41.872 219.294 41.976 223.668 ; 
        RECT 41.44 219.294 41.544 223.668 ; 
        RECT 41.008 219.294 41.112 223.668 ; 
        RECT 40.576 219.294 40.68 223.668 ; 
        RECT 40.144 219.294 40.248 223.668 ; 
        RECT 39.712 219.294 39.816 223.668 ; 
        RECT 39.28 219.294 39.384 223.668 ; 
        RECT 38.848 219.294 38.952 223.668 ; 
        RECT 38.416 219.294 38.52 223.668 ; 
        RECT 37.984 219.294 38.088 223.668 ; 
        RECT 37.552 219.294 37.656 223.668 ; 
        RECT 37.12 219.294 37.224 223.668 ; 
        RECT 36.688 219.294 36.792 223.668 ; 
        RECT 36.256 219.294 36.36 223.668 ; 
        RECT 35.824 219.294 35.928 223.668 ; 
        RECT 35.392 219.294 35.496 223.668 ; 
        RECT 34.96 219.294 35.064 223.668 ; 
        RECT 34.528 219.294 34.632 223.668 ; 
        RECT 34.096 219.294 34.2 223.668 ; 
        RECT 33.664 219.294 33.768 223.668 ; 
        RECT 33.232 219.294 33.336 223.668 ; 
        RECT 32.8 219.294 32.904 223.668 ; 
        RECT 32.368 219.294 32.472 223.668 ; 
        RECT 31.936 219.294 32.04 223.668 ; 
        RECT 31.504 219.294 31.608 223.668 ; 
        RECT 31.072 219.294 31.176 223.668 ; 
        RECT 30.64 219.294 30.744 223.668 ; 
        RECT 30.208 219.294 30.312 223.668 ; 
        RECT 29.776 219.294 29.88 223.668 ; 
        RECT 29.344 219.294 29.448 223.668 ; 
        RECT 28.912 219.294 29.016 223.668 ; 
        RECT 28.48 219.294 28.584 223.668 ; 
        RECT 28.048 219.294 28.152 223.668 ; 
        RECT 27.616 219.294 27.72 223.668 ; 
        RECT 27.184 219.294 27.288 223.668 ; 
        RECT 26.752 219.294 26.856 223.668 ; 
        RECT 26.32 219.294 26.424 223.668 ; 
        RECT 25.888 219.294 25.992 223.668 ; 
        RECT 25.456 219.294 25.56 223.668 ; 
        RECT 25.024 219.294 25.128 223.668 ; 
        RECT 24.592 219.294 24.696 223.668 ; 
        RECT 24.16 219.294 24.264 223.668 ; 
        RECT 23.728 219.294 23.832 223.668 ; 
        RECT 23.296 219.294 23.4 223.668 ; 
        RECT 22.864 219.294 22.968 223.668 ; 
        RECT 22.432 219.294 22.536 223.668 ; 
        RECT 22 219.294 22.104 223.668 ; 
        RECT 21.568 219.294 21.672 223.668 ; 
        RECT 21.136 219.294 21.24 223.668 ; 
        RECT 20.704 219.294 20.808 223.668 ; 
        RECT 20.272 219.294 20.376 223.668 ; 
        RECT 19.84 219.294 19.944 223.668 ; 
        RECT 19.408 219.294 19.512 223.668 ; 
        RECT 18.976 219.294 19.08 223.668 ; 
        RECT 18.544 219.294 18.648 223.668 ; 
        RECT 18.112 219.294 18.216 223.668 ; 
        RECT 17.68 219.294 17.784 223.668 ; 
        RECT 17.248 219.294 17.352 223.668 ; 
        RECT 16.816 219.294 16.92 223.668 ; 
        RECT 16.384 219.294 16.488 223.668 ; 
        RECT 15.952 219.294 16.056 223.668 ; 
        RECT 15.52 219.294 15.624 223.668 ; 
        RECT 15.088 219.294 15.192 223.668 ; 
        RECT 14.656 219.294 14.76 223.668 ; 
        RECT 14.224 219.294 14.328 223.668 ; 
        RECT 13.792 219.294 13.896 223.668 ; 
        RECT 13.36 219.294 13.464 223.668 ; 
        RECT 12.928 219.294 13.032 223.668 ; 
        RECT 12.496 219.294 12.6 223.668 ; 
        RECT 12.064 219.294 12.168 223.668 ; 
        RECT 11.632 219.294 11.736 223.668 ; 
        RECT 11.2 219.294 11.304 223.668 ; 
        RECT 10.768 219.294 10.872 223.668 ; 
        RECT 10.336 219.294 10.44 223.668 ; 
        RECT 9.904 219.294 10.008 223.668 ; 
        RECT 9.472 219.294 9.576 223.668 ; 
        RECT 9.04 219.294 9.144 223.668 ; 
        RECT 8.608 219.294 8.712 223.668 ; 
        RECT 8.176 219.294 8.28 223.668 ; 
        RECT 7.744 219.294 7.848 223.668 ; 
        RECT 7.312 219.294 7.416 223.668 ; 
        RECT 6.88 219.294 6.984 223.668 ; 
        RECT 6.448 219.294 6.552 223.668 ; 
        RECT 6.016 219.294 6.12 223.668 ; 
        RECT 5.584 219.294 5.688 223.668 ; 
        RECT 5.152 219.294 5.256 223.668 ; 
        RECT 4.72 219.294 4.824 223.668 ; 
        RECT 4.288 219.294 4.392 223.668 ; 
        RECT 3.856 219.294 3.96 223.668 ; 
        RECT 3.424 219.294 3.528 223.668 ; 
        RECT 2.992 219.294 3.096 223.668 ; 
        RECT 2.56 219.294 2.664 223.668 ; 
        RECT 2.128 219.294 2.232 223.668 ; 
        RECT 1.696 219.294 1.8 223.668 ; 
        RECT 1.264 219.294 1.368 223.668 ; 
        RECT 0.832 219.294 0.936 223.668 ; 
        RECT 0.02 219.294 0.36 223.668 ; 
        RECT 62.212 223.614 62.724 227.988 ; 
        RECT 62.156 226.276 62.724 227.566 ; 
        RECT 61.276 225.184 61.812 227.988 ; 
        RECT 61.184 226.524 61.812 227.556 ; 
        RECT 61.276 223.614 61.668 227.988 ; 
        RECT 61.276 224.098 61.724 225.056 ; 
        RECT 61.276 223.614 61.812 223.97 ; 
        RECT 60.376 225.416 60.912 227.988 ; 
        RECT 60.376 223.614 60.768 227.988 ; 
        RECT 58.708 223.614 59.04 227.988 ; 
        RECT 58.708 223.968 59.096 227.71 ; 
        RECT 121.072 223.614 121.412 227.988 ; 
        RECT 120.496 223.614 120.6 227.988 ; 
        RECT 120.064 223.614 120.168 227.988 ; 
        RECT 119.632 223.614 119.736 227.988 ; 
        RECT 119.2 223.614 119.304 227.988 ; 
        RECT 118.768 223.614 118.872 227.988 ; 
        RECT 118.336 223.614 118.44 227.988 ; 
        RECT 117.904 223.614 118.008 227.988 ; 
        RECT 117.472 223.614 117.576 227.988 ; 
        RECT 117.04 223.614 117.144 227.988 ; 
        RECT 116.608 223.614 116.712 227.988 ; 
        RECT 116.176 223.614 116.28 227.988 ; 
        RECT 115.744 223.614 115.848 227.988 ; 
        RECT 115.312 223.614 115.416 227.988 ; 
        RECT 114.88 223.614 114.984 227.988 ; 
        RECT 114.448 223.614 114.552 227.988 ; 
        RECT 114.016 223.614 114.12 227.988 ; 
        RECT 113.584 223.614 113.688 227.988 ; 
        RECT 113.152 223.614 113.256 227.988 ; 
        RECT 112.72 223.614 112.824 227.988 ; 
        RECT 112.288 223.614 112.392 227.988 ; 
        RECT 111.856 223.614 111.96 227.988 ; 
        RECT 111.424 223.614 111.528 227.988 ; 
        RECT 110.992 223.614 111.096 227.988 ; 
        RECT 110.56 223.614 110.664 227.988 ; 
        RECT 110.128 223.614 110.232 227.988 ; 
        RECT 109.696 223.614 109.8 227.988 ; 
        RECT 109.264 223.614 109.368 227.988 ; 
        RECT 108.832 223.614 108.936 227.988 ; 
        RECT 108.4 223.614 108.504 227.988 ; 
        RECT 107.968 223.614 108.072 227.988 ; 
        RECT 107.536 223.614 107.64 227.988 ; 
        RECT 107.104 223.614 107.208 227.988 ; 
        RECT 106.672 223.614 106.776 227.988 ; 
        RECT 106.24 223.614 106.344 227.988 ; 
        RECT 105.808 223.614 105.912 227.988 ; 
        RECT 105.376 223.614 105.48 227.988 ; 
        RECT 104.944 223.614 105.048 227.988 ; 
        RECT 104.512 223.614 104.616 227.988 ; 
        RECT 104.08 223.614 104.184 227.988 ; 
        RECT 103.648 223.614 103.752 227.988 ; 
        RECT 103.216 223.614 103.32 227.988 ; 
        RECT 102.784 223.614 102.888 227.988 ; 
        RECT 102.352 223.614 102.456 227.988 ; 
        RECT 101.92 223.614 102.024 227.988 ; 
        RECT 101.488 223.614 101.592 227.988 ; 
        RECT 101.056 223.614 101.16 227.988 ; 
        RECT 100.624 223.614 100.728 227.988 ; 
        RECT 100.192 223.614 100.296 227.988 ; 
        RECT 99.76 223.614 99.864 227.988 ; 
        RECT 99.328 223.614 99.432 227.988 ; 
        RECT 98.896 223.614 99 227.988 ; 
        RECT 98.464 223.614 98.568 227.988 ; 
        RECT 98.032 223.614 98.136 227.988 ; 
        RECT 97.6 223.614 97.704 227.988 ; 
        RECT 97.168 223.614 97.272 227.988 ; 
        RECT 96.736 223.614 96.84 227.988 ; 
        RECT 96.304 223.614 96.408 227.988 ; 
        RECT 95.872 223.614 95.976 227.988 ; 
        RECT 95.44 223.614 95.544 227.988 ; 
        RECT 95.008 223.614 95.112 227.988 ; 
        RECT 94.576 223.614 94.68 227.988 ; 
        RECT 94.144 223.614 94.248 227.988 ; 
        RECT 93.712 223.614 93.816 227.988 ; 
        RECT 93.28 223.614 93.384 227.988 ; 
        RECT 92.848 223.614 92.952 227.988 ; 
        RECT 92.416 223.614 92.52 227.988 ; 
        RECT 91.984 223.614 92.088 227.988 ; 
        RECT 91.552 223.614 91.656 227.988 ; 
        RECT 91.12 223.614 91.224 227.988 ; 
        RECT 90.688 223.614 90.792 227.988 ; 
        RECT 90.256 223.614 90.36 227.988 ; 
        RECT 89.824 223.614 89.928 227.988 ; 
        RECT 89.392 223.614 89.496 227.988 ; 
        RECT 88.96 223.614 89.064 227.988 ; 
        RECT 88.528 223.614 88.632 227.988 ; 
        RECT 88.096 223.614 88.2 227.988 ; 
        RECT 87.664 223.614 87.768 227.988 ; 
        RECT 87.232 223.614 87.336 227.988 ; 
        RECT 86.8 223.614 86.904 227.988 ; 
        RECT 86.368 223.614 86.472 227.988 ; 
        RECT 85.936 223.614 86.04 227.988 ; 
        RECT 85.504 223.614 85.608 227.988 ; 
        RECT 85.072 223.614 85.176 227.988 ; 
        RECT 84.64 223.614 84.744 227.988 ; 
        RECT 84.208 223.614 84.312 227.988 ; 
        RECT 83.776 223.614 83.88 227.988 ; 
        RECT 83.344 223.614 83.448 227.988 ; 
        RECT 82.912 223.614 83.016 227.988 ; 
        RECT 82.48 223.614 82.584 227.988 ; 
        RECT 82.048 223.614 82.152 227.988 ; 
        RECT 81.616 223.614 81.72 227.988 ; 
        RECT 81.184 223.614 81.288 227.988 ; 
        RECT 80.752 223.614 80.856 227.988 ; 
        RECT 80.32 223.614 80.424 227.988 ; 
        RECT 79.888 223.614 79.992 227.988 ; 
        RECT 79.456 223.614 79.56 227.988 ; 
        RECT 79.024 223.614 79.128 227.988 ; 
        RECT 78.592 223.614 78.696 227.988 ; 
        RECT 78.16 223.614 78.264 227.988 ; 
        RECT 77.728 223.614 77.832 227.988 ; 
        RECT 77.296 223.614 77.4 227.988 ; 
        RECT 76.864 223.614 76.968 227.988 ; 
        RECT 76.432 223.614 76.536 227.988 ; 
        RECT 76 223.614 76.104 227.988 ; 
        RECT 75.568 223.614 75.672 227.988 ; 
        RECT 75.136 223.614 75.24 227.988 ; 
        RECT 74.704 223.614 74.808 227.988 ; 
        RECT 74.272 223.614 74.376 227.988 ; 
        RECT 73.84 223.614 73.944 227.988 ; 
        RECT 73.408 223.614 73.512 227.988 ; 
        RECT 72.976 223.614 73.08 227.988 ; 
        RECT 72.544 223.614 72.648 227.988 ; 
        RECT 72.112 223.614 72.216 227.988 ; 
        RECT 71.68 223.614 71.784 227.988 ; 
        RECT 71.248 223.614 71.352 227.988 ; 
        RECT 70.816 223.614 70.92 227.988 ; 
        RECT 70.384 223.614 70.488 227.988 ; 
        RECT 69.952 223.614 70.056 227.988 ; 
        RECT 69.52 223.614 69.624 227.988 ; 
        RECT 69.088 223.614 69.192 227.988 ; 
        RECT 68.656 223.614 68.76 227.988 ; 
        RECT 68.224 223.614 68.328 227.988 ; 
        RECT 67.792 223.614 67.896 227.988 ; 
        RECT 67.36 223.614 67.464 227.988 ; 
        RECT 66.928 223.614 67.032 227.988 ; 
        RECT 66.496 223.614 66.6 227.988 ; 
        RECT 66.064 223.614 66.168 227.988 ; 
        RECT 65.632 223.614 65.736 227.988 ; 
        RECT 65.2 223.614 65.304 227.988 ; 
        RECT 64.348 223.614 64.656 227.988 ; 
        RECT 56.776 223.614 57.084 227.988 ; 
        RECT 56.128 223.614 56.232 227.988 ; 
        RECT 55.696 223.614 55.8 227.988 ; 
        RECT 55.264 223.614 55.368 227.988 ; 
        RECT 54.832 223.614 54.936 227.988 ; 
        RECT 54.4 223.614 54.504 227.988 ; 
        RECT 53.968 223.614 54.072 227.988 ; 
        RECT 53.536 223.614 53.64 227.988 ; 
        RECT 53.104 223.614 53.208 227.988 ; 
        RECT 52.672 223.614 52.776 227.988 ; 
        RECT 52.24 223.614 52.344 227.988 ; 
        RECT 51.808 223.614 51.912 227.988 ; 
        RECT 51.376 223.614 51.48 227.988 ; 
        RECT 50.944 223.614 51.048 227.988 ; 
        RECT 50.512 223.614 50.616 227.988 ; 
        RECT 50.08 223.614 50.184 227.988 ; 
        RECT 49.648 223.614 49.752 227.988 ; 
        RECT 49.216 223.614 49.32 227.988 ; 
        RECT 48.784 223.614 48.888 227.988 ; 
        RECT 48.352 223.614 48.456 227.988 ; 
        RECT 47.92 223.614 48.024 227.988 ; 
        RECT 47.488 223.614 47.592 227.988 ; 
        RECT 47.056 223.614 47.16 227.988 ; 
        RECT 46.624 223.614 46.728 227.988 ; 
        RECT 46.192 223.614 46.296 227.988 ; 
        RECT 45.76 223.614 45.864 227.988 ; 
        RECT 45.328 223.614 45.432 227.988 ; 
        RECT 44.896 223.614 45 227.988 ; 
        RECT 44.464 223.614 44.568 227.988 ; 
        RECT 44.032 223.614 44.136 227.988 ; 
        RECT 43.6 223.614 43.704 227.988 ; 
        RECT 43.168 223.614 43.272 227.988 ; 
        RECT 42.736 223.614 42.84 227.988 ; 
        RECT 42.304 223.614 42.408 227.988 ; 
        RECT 41.872 223.614 41.976 227.988 ; 
        RECT 41.44 223.614 41.544 227.988 ; 
        RECT 41.008 223.614 41.112 227.988 ; 
        RECT 40.576 223.614 40.68 227.988 ; 
        RECT 40.144 223.614 40.248 227.988 ; 
        RECT 39.712 223.614 39.816 227.988 ; 
        RECT 39.28 223.614 39.384 227.988 ; 
        RECT 38.848 223.614 38.952 227.988 ; 
        RECT 38.416 223.614 38.52 227.988 ; 
        RECT 37.984 223.614 38.088 227.988 ; 
        RECT 37.552 223.614 37.656 227.988 ; 
        RECT 37.12 223.614 37.224 227.988 ; 
        RECT 36.688 223.614 36.792 227.988 ; 
        RECT 36.256 223.614 36.36 227.988 ; 
        RECT 35.824 223.614 35.928 227.988 ; 
        RECT 35.392 223.614 35.496 227.988 ; 
        RECT 34.96 223.614 35.064 227.988 ; 
        RECT 34.528 223.614 34.632 227.988 ; 
        RECT 34.096 223.614 34.2 227.988 ; 
        RECT 33.664 223.614 33.768 227.988 ; 
        RECT 33.232 223.614 33.336 227.988 ; 
        RECT 32.8 223.614 32.904 227.988 ; 
        RECT 32.368 223.614 32.472 227.988 ; 
        RECT 31.936 223.614 32.04 227.988 ; 
        RECT 31.504 223.614 31.608 227.988 ; 
        RECT 31.072 223.614 31.176 227.988 ; 
        RECT 30.64 223.614 30.744 227.988 ; 
        RECT 30.208 223.614 30.312 227.988 ; 
        RECT 29.776 223.614 29.88 227.988 ; 
        RECT 29.344 223.614 29.448 227.988 ; 
        RECT 28.912 223.614 29.016 227.988 ; 
        RECT 28.48 223.614 28.584 227.988 ; 
        RECT 28.048 223.614 28.152 227.988 ; 
        RECT 27.616 223.614 27.72 227.988 ; 
        RECT 27.184 223.614 27.288 227.988 ; 
        RECT 26.752 223.614 26.856 227.988 ; 
        RECT 26.32 223.614 26.424 227.988 ; 
        RECT 25.888 223.614 25.992 227.988 ; 
        RECT 25.456 223.614 25.56 227.988 ; 
        RECT 25.024 223.614 25.128 227.988 ; 
        RECT 24.592 223.614 24.696 227.988 ; 
        RECT 24.16 223.614 24.264 227.988 ; 
        RECT 23.728 223.614 23.832 227.988 ; 
        RECT 23.296 223.614 23.4 227.988 ; 
        RECT 22.864 223.614 22.968 227.988 ; 
        RECT 22.432 223.614 22.536 227.988 ; 
        RECT 22 223.614 22.104 227.988 ; 
        RECT 21.568 223.614 21.672 227.988 ; 
        RECT 21.136 223.614 21.24 227.988 ; 
        RECT 20.704 223.614 20.808 227.988 ; 
        RECT 20.272 223.614 20.376 227.988 ; 
        RECT 19.84 223.614 19.944 227.988 ; 
        RECT 19.408 223.614 19.512 227.988 ; 
        RECT 18.976 223.614 19.08 227.988 ; 
        RECT 18.544 223.614 18.648 227.988 ; 
        RECT 18.112 223.614 18.216 227.988 ; 
        RECT 17.68 223.614 17.784 227.988 ; 
        RECT 17.248 223.614 17.352 227.988 ; 
        RECT 16.816 223.614 16.92 227.988 ; 
        RECT 16.384 223.614 16.488 227.988 ; 
        RECT 15.952 223.614 16.056 227.988 ; 
        RECT 15.52 223.614 15.624 227.988 ; 
        RECT 15.088 223.614 15.192 227.988 ; 
        RECT 14.656 223.614 14.76 227.988 ; 
        RECT 14.224 223.614 14.328 227.988 ; 
        RECT 13.792 223.614 13.896 227.988 ; 
        RECT 13.36 223.614 13.464 227.988 ; 
        RECT 12.928 223.614 13.032 227.988 ; 
        RECT 12.496 223.614 12.6 227.988 ; 
        RECT 12.064 223.614 12.168 227.988 ; 
        RECT 11.632 223.614 11.736 227.988 ; 
        RECT 11.2 223.614 11.304 227.988 ; 
        RECT 10.768 223.614 10.872 227.988 ; 
        RECT 10.336 223.614 10.44 227.988 ; 
        RECT 9.904 223.614 10.008 227.988 ; 
        RECT 9.472 223.614 9.576 227.988 ; 
        RECT 9.04 223.614 9.144 227.988 ; 
        RECT 8.608 223.614 8.712 227.988 ; 
        RECT 8.176 223.614 8.28 227.988 ; 
        RECT 7.744 223.614 7.848 227.988 ; 
        RECT 7.312 223.614 7.416 227.988 ; 
        RECT 6.88 223.614 6.984 227.988 ; 
        RECT 6.448 223.614 6.552 227.988 ; 
        RECT 6.016 223.614 6.12 227.988 ; 
        RECT 5.584 223.614 5.688 227.988 ; 
        RECT 5.152 223.614 5.256 227.988 ; 
        RECT 4.72 223.614 4.824 227.988 ; 
        RECT 4.288 223.614 4.392 227.988 ; 
        RECT 3.856 223.614 3.96 227.988 ; 
        RECT 3.424 223.614 3.528 227.988 ; 
        RECT 2.992 223.614 3.096 227.988 ; 
        RECT 2.56 223.614 2.664 227.988 ; 
        RECT 2.128 223.614 2.232 227.988 ; 
        RECT 1.696 223.614 1.8 227.988 ; 
        RECT 1.264 223.614 1.368 227.988 ; 
        RECT 0.832 223.614 0.936 227.988 ; 
        RECT 0.02 223.614 0.36 227.988 ; 
        RECT 62.212 227.934 62.724 232.308 ; 
        RECT 62.156 230.596 62.724 231.886 ; 
        RECT 61.276 229.504 61.812 232.308 ; 
        RECT 61.184 230.844 61.812 231.876 ; 
        RECT 61.276 227.934 61.668 232.308 ; 
        RECT 61.276 228.418 61.724 229.376 ; 
        RECT 61.276 227.934 61.812 228.29 ; 
        RECT 60.376 229.736 60.912 232.308 ; 
        RECT 60.376 227.934 60.768 232.308 ; 
        RECT 58.708 227.934 59.04 232.308 ; 
        RECT 58.708 228.288 59.096 232.03 ; 
        RECT 121.072 227.934 121.412 232.308 ; 
        RECT 120.496 227.934 120.6 232.308 ; 
        RECT 120.064 227.934 120.168 232.308 ; 
        RECT 119.632 227.934 119.736 232.308 ; 
        RECT 119.2 227.934 119.304 232.308 ; 
        RECT 118.768 227.934 118.872 232.308 ; 
        RECT 118.336 227.934 118.44 232.308 ; 
        RECT 117.904 227.934 118.008 232.308 ; 
        RECT 117.472 227.934 117.576 232.308 ; 
        RECT 117.04 227.934 117.144 232.308 ; 
        RECT 116.608 227.934 116.712 232.308 ; 
        RECT 116.176 227.934 116.28 232.308 ; 
        RECT 115.744 227.934 115.848 232.308 ; 
        RECT 115.312 227.934 115.416 232.308 ; 
        RECT 114.88 227.934 114.984 232.308 ; 
        RECT 114.448 227.934 114.552 232.308 ; 
        RECT 114.016 227.934 114.12 232.308 ; 
        RECT 113.584 227.934 113.688 232.308 ; 
        RECT 113.152 227.934 113.256 232.308 ; 
        RECT 112.72 227.934 112.824 232.308 ; 
        RECT 112.288 227.934 112.392 232.308 ; 
        RECT 111.856 227.934 111.96 232.308 ; 
        RECT 111.424 227.934 111.528 232.308 ; 
        RECT 110.992 227.934 111.096 232.308 ; 
        RECT 110.56 227.934 110.664 232.308 ; 
        RECT 110.128 227.934 110.232 232.308 ; 
        RECT 109.696 227.934 109.8 232.308 ; 
        RECT 109.264 227.934 109.368 232.308 ; 
        RECT 108.832 227.934 108.936 232.308 ; 
        RECT 108.4 227.934 108.504 232.308 ; 
        RECT 107.968 227.934 108.072 232.308 ; 
        RECT 107.536 227.934 107.64 232.308 ; 
        RECT 107.104 227.934 107.208 232.308 ; 
        RECT 106.672 227.934 106.776 232.308 ; 
        RECT 106.24 227.934 106.344 232.308 ; 
        RECT 105.808 227.934 105.912 232.308 ; 
        RECT 105.376 227.934 105.48 232.308 ; 
        RECT 104.944 227.934 105.048 232.308 ; 
        RECT 104.512 227.934 104.616 232.308 ; 
        RECT 104.08 227.934 104.184 232.308 ; 
        RECT 103.648 227.934 103.752 232.308 ; 
        RECT 103.216 227.934 103.32 232.308 ; 
        RECT 102.784 227.934 102.888 232.308 ; 
        RECT 102.352 227.934 102.456 232.308 ; 
        RECT 101.92 227.934 102.024 232.308 ; 
        RECT 101.488 227.934 101.592 232.308 ; 
        RECT 101.056 227.934 101.16 232.308 ; 
        RECT 100.624 227.934 100.728 232.308 ; 
        RECT 100.192 227.934 100.296 232.308 ; 
        RECT 99.76 227.934 99.864 232.308 ; 
        RECT 99.328 227.934 99.432 232.308 ; 
        RECT 98.896 227.934 99 232.308 ; 
        RECT 98.464 227.934 98.568 232.308 ; 
        RECT 98.032 227.934 98.136 232.308 ; 
        RECT 97.6 227.934 97.704 232.308 ; 
        RECT 97.168 227.934 97.272 232.308 ; 
        RECT 96.736 227.934 96.84 232.308 ; 
        RECT 96.304 227.934 96.408 232.308 ; 
        RECT 95.872 227.934 95.976 232.308 ; 
        RECT 95.44 227.934 95.544 232.308 ; 
        RECT 95.008 227.934 95.112 232.308 ; 
        RECT 94.576 227.934 94.68 232.308 ; 
        RECT 94.144 227.934 94.248 232.308 ; 
        RECT 93.712 227.934 93.816 232.308 ; 
        RECT 93.28 227.934 93.384 232.308 ; 
        RECT 92.848 227.934 92.952 232.308 ; 
        RECT 92.416 227.934 92.52 232.308 ; 
        RECT 91.984 227.934 92.088 232.308 ; 
        RECT 91.552 227.934 91.656 232.308 ; 
        RECT 91.12 227.934 91.224 232.308 ; 
        RECT 90.688 227.934 90.792 232.308 ; 
        RECT 90.256 227.934 90.36 232.308 ; 
        RECT 89.824 227.934 89.928 232.308 ; 
        RECT 89.392 227.934 89.496 232.308 ; 
        RECT 88.96 227.934 89.064 232.308 ; 
        RECT 88.528 227.934 88.632 232.308 ; 
        RECT 88.096 227.934 88.2 232.308 ; 
        RECT 87.664 227.934 87.768 232.308 ; 
        RECT 87.232 227.934 87.336 232.308 ; 
        RECT 86.8 227.934 86.904 232.308 ; 
        RECT 86.368 227.934 86.472 232.308 ; 
        RECT 85.936 227.934 86.04 232.308 ; 
        RECT 85.504 227.934 85.608 232.308 ; 
        RECT 85.072 227.934 85.176 232.308 ; 
        RECT 84.64 227.934 84.744 232.308 ; 
        RECT 84.208 227.934 84.312 232.308 ; 
        RECT 83.776 227.934 83.88 232.308 ; 
        RECT 83.344 227.934 83.448 232.308 ; 
        RECT 82.912 227.934 83.016 232.308 ; 
        RECT 82.48 227.934 82.584 232.308 ; 
        RECT 82.048 227.934 82.152 232.308 ; 
        RECT 81.616 227.934 81.72 232.308 ; 
        RECT 81.184 227.934 81.288 232.308 ; 
        RECT 80.752 227.934 80.856 232.308 ; 
        RECT 80.32 227.934 80.424 232.308 ; 
        RECT 79.888 227.934 79.992 232.308 ; 
        RECT 79.456 227.934 79.56 232.308 ; 
        RECT 79.024 227.934 79.128 232.308 ; 
        RECT 78.592 227.934 78.696 232.308 ; 
        RECT 78.16 227.934 78.264 232.308 ; 
        RECT 77.728 227.934 77.832 232.308 ; 
        RECT 77.296 227.934 77.4 232.308 ; 
        RECT 76.864 227.934 76.968 232.308 ; 
        RECT 76.432 227.934 76.536 232.308 ; 
        RECT 76 227.934 76.104 232.308 ; 
        RECT 75.568 227.934 75.672 232.308 ; 
        RECT 75.136 227.934 75.24 232.308 ; 
        RECT 74.704 227.934 74.808 232.308 ; 
        RECT 74.272 227.934 74.376 232.308 ; 
        RECT 73.84 227.934 73.944 232.308 ; 
        RECT 73.408 227.934 73.512 232.308 ; 
        RECT 72.976 227.934 73.08 232.308 ; 
        RECT 72.544 227.934 72.648 232.308 ; 
        RECT 72.112 227.934 72.216 232.308 ; 
        RECT 71.68 227.934 71.784 232.308 ; 
        RECT 71.248 227.934 71.352 232.308 ; 
        RECT 70.816 227.934 70.92 232.308 ; 
        RECT 70.384 227.934 70.488 232.308 ; 
        RECT 69.952 227.934 70.056 232.308 ; 
        RECT 69.52 227.934 69.624 232.308 ; 
        RECT 69.088 227.934 69.192 232.308 ; 
        RECT 68.656 227.934 68.76 232.308 ; 
        RECT 68.224 227.934 68.328 232.308 ; 
        RECT 67.792 227.934 67.896 232.308 ; 
        RECT 67.36 227.934 67.464 232.308 ; 
        RECT 66.928 227.934 67.032 232.308 ; 
        RECT 66.496 227.934 66.6 232.308 ; 
        RECT 66.064 227.934 66.168 232.308 ; 
        RECT 65.632 227.934 65.736 232.308 ; 
        RECT 65.2 227.934 65.304 232.308 ; 
        RECT 64.348 227.934 64.656 232.308 ; 
        RECT 56.776 227.934 57.084 232.308 ; 
        RECT 56.128 227.934 56.232 232.308 ; 
        RECT 55.696 227.934 55.8 232.308 ; 
        RECT 55.264 227.934 55.368 232.308 ; 
        RECT 54.832 227.934 54.936 232.308 ; 
        RECT 54.4 227.934 54.504 232.308 ; 
        RECT 53.968 227.934 54.072 232.308 ; 
        RECT 53.536 227.934 53.64 232.308 ; 
        RECT 53.104 227.934 53.208 232.308 ; 
        RECT 52.672 227.934 52.776 232.308 ; 
        RECT 52.24 227.934 52.344 232.308 ; 
        RECT 51.808 227.934 51.912 232.308 ; 
        RECT 51.376 227.934 51.48 232.308 ; 
        RECT 50.944 227.934 51.048 232.308 ; 
        RECT 50.512 227.934 50.616 232.308 ; 
        RECT 50.08 227.934 50.184 232.308 ; 
        RECT 49.648 227.934 49.752 232.308 ; 
        RECT 49.216 227.934 49.32 232.308 ; 
        RECT 48.784 227.934 48.888 232.308 ; 
        RECT 48.352 227.934 48.456 232.308 ; 
        RECT 47.92 227.934 48.024 232.308 ; 
        RECT 47.488 227.934 47.592 232.308 ; 
        RECT 47.056 227.934 47.16 232.308 ; 
        RECT 46.624 227.934 46.728 232.308 ; 
        RECT 46.192 227.934 46.296 232.308 ; 
        RECT 45.76 227.934 45.864 232.308 ; 
        RECT 45.328 227.934 45.432 232.308 ; 
        RECT 44.896 227.934 45 232.308 ; 
        RECT 44.464 227.934 44.568 232.308 ; 
        RECT 44.032 227.934 44.136 232.308 ; 
        RECT 43.6 227.934 43.704 232.308 ; 
        RECT 43.168 227.934 43.272 232.308 ; 
        RECT 42.736 227.934 42.84 232.308 ; 
        RECT 42.304 227.934 42.408 232.308 ; 
        RECT 41.872 227.934 41.976 232.308 ; 
        RECT 41.44 227.934 41.544 232.308 ; 
        RECT 41.008 227.934 41.112 232.308 ; 
        RECT 40.576 227.934 40.68 232.308 ; 
        RECT 40.144 227.934 40.248 232.308 ; 
        RECT 39.712 227.934 39.816 232.308 ; 
        RECT 39.28 227.934 39.384 232.308 ; 
        RECT 38.848 227.934 38.952 232.308 ; 
        RECT 38.416 227.934 38.52 232.308 ; 
        RECT 37.984 227.934 38.088 232.308 ; 
        RECT 37.552 227.934 37.656 232.308 ; 
        RECT 37.12 227.934 37.224 232.308 ; 
        RECT 36.688 227.934 36.792 232.308 ; 
        RECT 36.256 227.934 36.36 232.308 ; 
        RECT 35.824 227.934 35.928 232.308 ; 
        RECT 35.392 227.934 35.496 232.308 ; 
        RECT 34.96 227.934 35.064 232.308 ; 
        RECT 34.528 227.934 34.632 232.308 ; 
        RECT 34.096 227.934 34.2 232.308 ; 
        RECT 33.664 227.934 33.768 232.308 ; 
        RECT 33.232 227.934 33.336 232.308 ; 
        RECT 32.8 227.934 32.904 232.308 ; 
        RECT 32.368 227.934 32.472 232.308 ; 
        RECT 31.936 227.934 32.04 232.308 ; 
        RECT 31.504 227.934 31.608 232.308 ; 
        RECT 31.072 227.934 31.176 232.308 ; 
        RECT 30.64 227.934 30.744 232.308 ; 
        RECT 30.208 227.934 30.312 232.308 ; 
        RECT 29.776 227.934 29.88 232.308 ; 
        RECT 29.344 227.934 29.448 232.308 ; 
        RECT 28.912 227.934 29.016 232.308 ; 
        RECT 28.48 227.934 28.584 232.308 ; 
        RECT 28.048 227.934 28.152 232.308 ; 
        RECT 27.616 227.934 27.72 232.308 ; 
        RECT 27.184 227.934 27.288 232.308 ; 
        RECT 26.752 227.934 26.856 232.308 ; 
        RECT 26.32 227.934 26.424 232.308 ; 
        RECT 25.888 227.934 25.992 232.308 ; 
        RECT 25.456 227.934 25.56 232.308 ; 
        RECT 25.024 227.934 25.128 232.308 ; 
        RECT 24.592 227.934 24.696 232.308 ; 
        RECT 24.16 227.934 24.264 232.308 ; 
        RECT 23.728 227.934 23.832 232.308 ; 
        RECT 23.296 227.934 23.4 232.308 ; 
        RECT 22.864 227.934 22.968 232.308 ; 
        RECT 22.432 227.934 22.536 232.308 ; 
        RECT 22 227.934 22.104 232.308 ; 
        RECT 21.568 227.934 21.672 232.308 ; 
        RECT 21.136 227.934 21.24 232.308 ; 
        RECT 20.704 227.934 20.808 232.308 ; 
        RECT 20.272 227.934 20.376 232.308 ; 
        RECT 19.84 227.934 19.944 232.308 ; 
        RECT 19.408 227.934 19.512 232.308 ; 
        RECT 18.976 227.934 19.08 232.308 ; 
        RECT 18.544 227.934 18.648 232.308 ; 
        RECT 18.112 227.934 18.216 232.308 ; 
        RECT 17.68 227.934 17.784 232.308 ; 
        RECT 17.248 227.934 17.352 232.308 ; 
        RECT 16.816 227.934 16.92 232.308 ; 
        RECT 16.384 227.934 16.488 232.308 ; 
        RECT 15.952 227.934 16.056 232.308 ; 
        RECT 15.52 227.934 15.624 232.308 ; 
        RECT 15.088 227.934 15.192 232.308 ; 
        RECT 14.656 227.934 14.76 232.308 ; 
        RECT 14.224 227.934 14.328 232.308 ; 
        RECT 13.792 227.934 13.896 232.308 ; 
        RECT 13.36 227.934 13.464 232.308 ; 
        RECT 12.928 227.934 13.032 232.308 ; 
        RECT 12.496 227.934 12.6 232.308 ; 
        RECT 12.064 227.934 12.168 232.308 ; 
        RECT 11.632 227.934 11.736 232.308 ; 
        RECT 11.2 227.934 11.304 232.308 ; 
        RECT 10.768 227.934 10.872 232.308 ; 
        RECT 10.336 227.934 10.44 232.308 ; 
        RECT 9.904 227.934 10.008 232.308 ; 
        RECT 9.472 227.934 9.576 232.308 ; 
        RECT 9.04 227.934 9.144 232.308 ; 
        RECT 8.608 227.934 8.712 232.308 ; 
        RECT 8.176 227.934 8.28 232.308 ; 
        RECT 7.744 227.934 7.848 232.308 ; 
        RECT 7.312 227.934 7.416 232.308 ; 
        RECT 6.88 227.934 6.984 232.308 ; 
        RECT 6.448 227.934 6.552 232.308 ; 
        RECT 6.016 227.934 6.12 232.308 ; 
        RECT 5.584 227.934 5.688 232.308 ; 
        RECT 5.152 227.934 5.256 232.308 ; 
        RECT 4.72 227.934 4.824 232.308 ; 
        RECT 4.288 227.934 4.392 232.308 ; 
        RECT 3.856 227.934 3.96 232.308 ; 
        RECT 3.424 227.934 3.528 232.308 ; 
        RECT 2.992 227.934 3.096 232.308 ; 
        RECT 2.56 227.934 2.664 232.308 ; 
        RECT 2.128 227.934 2.232 232.308 ; 
        RECT 1.696 227.934 1.8 232.308 ; 
        RECT 1.264 227.934 1.368 232.308 ; 
        RECT 0.832 227.934 0.936 232.308 ; 
        RECT 0.02 227.934 0.36 232.308 ; 
        RECT 62.212 232.254 62.724 236.628 ; 
        RECT 62.156 234.916 62.724 236.206 ; 
        RECT 61.276 233.824 61.812 236.628 ; 
        RECT 61.184 235.164 61.812 236.196 ; 
        RECT 61.276 232.254 61.668 236.628 ; 
        RECT 61.276 232.738 61.724 233.696 ; 
        RECT 61.276 232.254 61.812 232.61 ; 
        RECT 60.376 234.056 60.912 236.628 ; 
        RECT 60.376 232.254 60.768 236.628 ; 
        RECT 58.708 232.254 59.04 236.628 ; 
        RECT 58.708 232.608 59.096 236.35 ; 
        RECT 121.072 232.254 121.412 236.628 ; 
        RECT 120.496 232.254 120.6 236.628 ; 
        RECT 120.064 232.254 120.168 236.628 ; 
        RECT 119.632 232.254 119.736 236.628 ; 
        RECT 119.2 232.254 119.304 236.628 ; 
        RECT 118.768 232.254 118.872 236.628 ; 
        RECT 118.336 232.254 118.44 236.628 ; 
        RECT 117.904 232.254 118.008 236.628 ; 
        RECT 117.472 232.254 117.576 236.628 ; 
        RECT 117.04 232.254 117.144 236.628 ; 
        RECT 116.608 232.254 116.712 236.628 ; 
        RECT 116.176 232.254 116.28 236.628 ; 
        RECT 115.744 232.254 115.848 236.628 ; 
        RECT 115.312 232.254 115.416 236.628 ; 
        RECT 114.88 232.254 114.984 236.628 ; 
        RECT 114.448 232.254 114.552 236.628 ; 
        RECT 114.016 232.254 114.12 236.628 ; 
        RECT 113.584 232.254 113.688 236.628 ; 
        RECT 113.152 232.254 113.256 236.628 ; 
        RECT 112.72 232.254 112.824 236.628 ; 
        RECT 112.288 232.254 112.392 236.628 ; 
        RECT 111.856 232.254 111.96 236.628 ; 
        RECT 111.424 232.254 111.528 236.628 ; 
        RECT 110.992 232.254 111.096 236.628 ; 
        RECT 110.56 232.254 110.664 236.628 ; 
        RECT 110.128 232.254 110.232 236.628 ; 
        RECT 109.696 232.254 109.8 236.628 ; 
        RECT 109.264 232.254 109.368 236.628 ; 
        RECT 108.832 232.254 108.936 236.628 ; 
        RECT 108.4 232.254 108.504 236.628 ; 
        RECT 107.968 232.254 108.072 236.628 ; 
        RECT 107.536 232.254 107.64 236.628 ; 
        RECT 107.104 232.254 107.208 236.628 ; 
        RECT 106.672 232.254 106.776 236.628 ; 
        RECT 106.24 232.254 106.344 236.628 ; 
        RECT 105.808 232.254 105.912 236.628 ; 
        RECT 105.376 232.254 105.48 236.628 ; 
        RECT 104.944 232.254 105.048 236.628 ; 
        RECT 104.512 232.254 104.616 236.628 ; 
        RECT 104.08 232.254 104.184 236.628 ; 
        RECT 103.648 232.254 103.752 236.628 ; 
        RECT 103.216 232.254 103.32 236.628 ; 
        RECT 102.784 232.254 102.888 236.628 ; 
        RECT 102.352 232.254 102.456 236.628 ; 
        RECT 101.92 232.254 102.024 236.628 ; 
        RECT 101.488 232.254 101.592 236.628 ; 
        RECT 101.056 232.254 101.16 236.628 ; 
        RECT 100.624 232.254 100.728 236.628 ; 
        RECT 100.192 232.254 100.296 236.628 ; 
        RECT 99.76 232.254 99.864 236.628 ; 
        RECT 99.328 232.254 99.432 236.628 ; 
        RECT 98.896 232.254 99 236.628 ; 
        RECT 98.464 232.254 98.568 236.628 ; 
        RECT 98.032 232.254 98.136 236.628 ; 
        RECT 97.6 232.254 97.704 236.628 ; 
        RECT 97.168 232.254 97.272 236.628 ; 
        RECT 96.736 232.254 96.84 236.628 ; 
        RECT 96.304 232.254 96.408 236.628 ; 
        RECT 95.872 232.254 95.976 236.628 ; 
        RECT 95.44 232.254 95.544 236.628 ; 
        RECT 95.008 232.254 95.112 236.628 ; 
        RECT 94.576 232.254 94.68 236.628 ; 
        RECT 94.144 232.254 94.248 236.628 ; 
        RECT 93.712 232.254 93.816 236.628 ; 
        RECT 93.28 232.254 93.384 236.628 ; 
        RECT 92.848 232.254 92.952 236.628 ; 
        RECT 92.416 232.254 92.52 236.628 ; 
        RECT 91.984 232.254 92.088 236.628 ; 
        RECT 91.552 232.254 91.656 236.628 ; 
        RECT 91.12 232.254 91.224 236.628 ; 
        RECT 90.688 232.254 90.792 236.628 ; 
        RECT 90.256 232.254 90.36 236.628 ; 
        RECT 89.824 232.254 89.928 236.628 ; 
        RECT 89.392 232.254 89.496 236.628 ; 
        RECT 88.96 232.254 89.064 236.628 ; 
        RECT 88.528 232.254 88.632 236.628 ; 
        RECT 88.096 232.254 88.2 236.628 ; 
        RECT 87.664 232.254 87.768 236.628 ; 
        RECT 87.232 232.254 87.336 236.628 ; 
        RECT 86.8 232.254 86.904 236.628 ; 
        RECT 86.368 232.254 86.472 236.628 ; 
        RECT 85.936 232.254 86.04 236.628 ; 
        RECT 85.504 232.254 85.608 236.628 ; 
        RECT 85.072 232.254 85.176 236.628 ; 
        RECT 84.64 232.254 84.744 236.628 ; 
        RECT 84.208 232.254 84.312 236.628 ; 
        RECT 83.776 232.254 83.88 236.628 ; 
        RECT 83.344 232.254 83.448 236.628 ; 
        RECT 82.912 232.254 83.016 236.628 ; 
        RECT 82.48 232.254 82.584 236.628 ; 
        RECT 82.048 232.254 82.152 236.628 ; 
        RECT 81.616 232.254 81.72 236.628 ; 
        RECT 81.184 232.254 81.288 236.628 ; 
        RECT 80.752 232.254 80.856 236.628 ; 
        RECT 80.32 232.254 80.424 236.628 ; 
        RECT 79.888 232.254 79.992 236.628 ; 
        RECT 79.456 232.254 79.56 236.628 ; 
        RECT 79.024 232.254 79.128 236.628 ; 
        RECT 78.592 232.254 78.696 236.628 ; 
        RECT 78.16 232.254 78.264 236.628 ; 
        RECT 77.728 232.254 77.832 236.628 ; 
        RECT 77.296 232.254 77.4 236.628 ; 
        RECT 76.864 232.254 76.968 236.628 ; 
        RECT 76.432 232.254 76.536 236.628 ; 
        RECT 76 232.254 76.104 236.628 ; 
        RECT 75.568 232.254 75.672 236.628 ; 
        RECT 75.136 232.254 75.24 236.628 ; 
        RECT 74.704 232.254 74.808 236.628 ; 
        RECT 74.272 232.254 74.376 236.628 ; 
        RECT 73.84 232.254 73.944 236.628 ; 
        RECT 73.408 232.254 73.512 236.628 ; 
        RECT 72.976 232.254 73.08 236.628 ; 
        RECT 72.544 232.254 72.648 236.628 ; 
        RECT 72.112 232.254 72.216 236.628 ; 
        RECT 71.68 232.254 71.784 236.628 ; 
        RECT 71.248 232.254 71.352 236.628 ; 
        RECT 70.816 232.254 70.92 236.628 ; 
        RECT 70.384 232.254 70.488 236.628 ; 
        RECT 69.952 232.254 70.056 236.628 ; 
        RECT 69.52 232.254 69.624 236.628 ; 
        RECT 69.088 232.254 69.192 236.628 ; 
        RECT 68.656 232.254 68.76 236.628 ; 
        RECT 68.224 232.254 68.328 236.628 ; 
        RECT 67.792 232.254 67.896 236.628 ; 
        RECT 67.36 232.254 67.464 236.628 ; 
        RECT 66.928 232.254 67.032 236.628 ; 
        RECT 66.496 232.254 66.6 236.628 ; 
        RECT 66.064 232.254 66.168 236.628 ; 
        RECT 65.632 232.254 65.736 236.628 ; 
        RECT 65.2 232.254 65.304 236.628 ; 
        RECT 64.348 232.254 64.656 236.628 ; 
        RECT 56.776 232.254 57.084 236.628 ; 
        RECT 56.128 232.254 56.232 236.628 ; 
        RECT 55.696 232.254 55.8 236.628 ; 
        RECT 55.264 232.254 55.368 236.628 ; 
        RECT 54.832 232.254 54.936 236.628 ; 
        RECT 54.4 232.254 54.504 236.628 ; 
        RECT 53.968 232.254 54.072 236.628 ; 
        RECT 53.536 232.254 53.64 236.628 ; 
        RECT 53.104 232.254 53.208 236.628 ; 
        RECT 52.672 232.254 52.776 236.628 ; 
        RECT 52.24 232.254 52.344 236.628 ; 
        RECT 51.808 232.254 51.912 236.628 ; 
        RECT 51.376 232.254 51.48 236.628 ; 
        RECT 50.944 232.254 51.048 236.628 ; 
        RECT 50.512 232.254 50.616 236.628 ; 
        RECT 50.08 232.254 50.184 236.628 ; 
        RECT 49.648 232.254 49.752 236.628 ; 
        RECT 49.216 232.254 49.32 236.628 ; 
        RECT 48.784 232.254 48.888 236.628 ; 
        RECT 48.352 232.254 48.456 236.628 ; 
        RECT 47.92 232.254 48.024 236.628 ; 
        RECT 47.488 232.254 47.592 236.628 ; 
        RECT 47.056 232.254 47.16 236.628 ; 
        RECT 46.624 232.254 46.728 236.628 ; 
        RECT 46.192 232.254 46.296 236.628 ; 
        RECT 45.76 232.254 45.864 236.628 ; 
        RECT 45.328 232.254 45.432 236.628 ; 
        RECT 44.896 232.254 45 236.628 ; 
        RECT 44.464 232.254 44.568 236.628 ; 
        RECT 44.032 232.254 44.136 236.628 ; 
        RECT 43.6 232.254 43.704 236.628 ; 
        RECT 43.168 232.254 43.272 236.628 ; 
        RECT 42.736 232.254 42.84 236.628 ; 
        RECT 42.304 232.254 42.408 236.628 ; 
        RECT 41.872 232.254 41.976 236.628 ; 
        RECT 41.44 232.254 41.544 236.628 ; 
        RECT 41.008 232.254 41.112 236.628 ; 
        RECT 40.576 232.254 40.68 236.628 ; 
        RECT 40.144 232.254 40.248 236.628 ; 
        RECT 39.712 232.254 39.816 236.628 ; 
        RECT 39.28 232.254 39.384 236.628 ; 
        RECT 38.848 232.254 38.952 236.628 ; 
        RECT 38.416 232.254 38.52 236.628 ; 
        RECT 37.984 232.254 38.088 236.628 ; 
        RECT 37.552 232.254 37.656 236.628 ; 
        RECT 37.12 232.254 37.224 236.628 ; 
        RECT 36.688 232.254 36.792 236.628 ; 
        RECT 36.256 232.254 36.36 236.628 ; 
        RECT 35.824 232.254 35.928 236.628 ; 
        RECT 35.392 232.254 35.496 236.628 ; 
        RECT 34.96 232.254 35.064 236.628 ; 
        RECT 34.528 232.254 34.632 236.628 ; 
        RECT 34.096 232.254 34.2 236.628 ; 
        RECT 33.664 232.254 33.768 236.628 ; 
        RECT 33.232 232.254 33.336 236.628 ; 
        RECT 32.8 232.254 32.904 236.628 ; 
        RECT 32.368 232.254 32.472 236.628 ; 
        RECT 31.936 232.254 32.04 236.628 ; 
        RECT 31.504 232.254 31.608 236.628 ; 
        RECT 31.072 232.254 31.176 236.628 ; 
        RECT 30.64 232.254 30.744 236.628 ; 
        RECT 30.208 232.254 30.312 236.628 ; 
        RECT 29.776 232.254 29.88 236.628 ; 
        RECT 29.344 232.254 29.448 236.628 ; 
        RECT 28.912 232.254 29.016 236.628 ; 
        RECT 28.48 232.254 28.584 236.628 ; 
        RECT 28.048 232.254 28.152 236.628 ; 
        RECT 27.616 232.254 27.72 236.628 ; 
        RECT 27.184 232.254 27.288 236.628 ; 
        RECT 26.752 232.254 26.856 236.628 ; 
        RECT 26.32 232.254 26.424 236.628 ; 
        RECT 25.888 232.254 25.992 236.628 ; 
        RECT 25.456 232.254 25.56 236.628 ; 
        RECT 25.024 232.254 25.128 236.628 ; 
        RECT 24.592 232.254 24.696 236.628 ; 
        RECT 24.16 232.254 24.264 236.628 ; 
        RECT 23.728 232.254 23.832 236.628 ; 
        RECT 23.296 232.254 23.4 236.628 ; 
        RECT 22.864 232.254 22.968 236.628 ; 
        RECT 22.432 232.254 22.536 236.628 ; 
        RECT 22 232.254 22.104 236.628 ; 
        RECT 21.568 232.254 21.672 236.628 ; 
        RECT 21.136 232.254 21.24 236.628 ; 
        RECT 20.704 232.254 20.808 236.628 ; 
        RECT 20.272 232.254 20.376 236.628 ; 
        RECT 19.84 232.254 19.944 236.628 ; 
        RECT 19.408 232.254 19.512 236.628 ; 
        RECT 18.976 232.254 19.08 236.628 ; 
        RECT 18.544 232.254 18.648 236.628 ; 
        RECT 18.112 232.254 18.216 236.628 ; 
        RECT 17.68 232.254 17.784 236.628 ; 
        RECT 17.248 232.254 17.352 236.628 ; 
        RECT 16.816 232.254 16.92 236.628 ; 
        RECT 16.384 232.254 16.488 236.628 ; 
        RECT 15.952 232.254 16.056 236.628 ; 
        RECT 15.52 232.254 15.624 236.628 ; 
        RECT 15.088 232.254 15.192 236.628 ; 
        RECT 14.656 232.254 14.76 236.628 ; 
        RECT 14.224 232.254 14.328 236.628 ; 
        RECT 13.792 232.254 13.896 236.628 ; 
        RECT 13.36 232.254 13.464 236.628 ; 
        RECT 12.928 232.254 13.032 236.628 ; 
        RECT 12.496 232.254 12.6 236.628 ; 
        RECT 12.064 232.254 12.168 236.628 ; 
        RECT 11.632 232.254 11.736 236.628 ; 
        RECT 11.2 232.254 11.304 236.628 ; 
        RECT 10.768 232.254 10.872 236.628 ; 
        RECT 10.336 232.254 10.44 236.628 ; 
        RECT 9.904 232.254 10.008 236.628 ; 
        RECT 9.472 232.254 9.576 236.628 ; 
        RECT 9.04 232.254 9.144 236.628 ; 
        RECT 8.608 232.254 8.712 236.628 ; 
        RECT 8.176 232.254 8.28 236.628 ; 
        RECT 7.744 232.254 7.848 236.628 ; 
        RECT 7.312 232.254 7.416 236.628 ; 
        RECT 6.88 232.254 6.984 236.628 ; 
        RECT 6.448 232.254 6.552 236.628 ; 
        RECT 6.016 232.254 6.12 236.628 ; 
        RECT 5.584 232.254 5.688 236.628 ; 
        RECT 5.152 232.254 5.256 236.628 ; 
        RECT 4.72 232.254 4.824 236.628 ; 
        RECT 4.288 232.254 4.392 236.628 ; 
        RECT 3.856 232.254 3.96 236.628 ; 
        RECT 3.424 232.254 3.528 236.628 ; 
        RECT 2.992 232.254 3.096 236.628 ; 
        RECT 2.56 232.254 2.664 236.628 ; 
        RECT 2.128 232.254 2.232 236.628 ; 
        RECT 1.696 232.254 1.8 236.628 ; 
        RECT 1.264 232.254 1.368 236.628 ; 
        RECT 0.832 232.254 0.936 236.628 ; 
        RECT 0.02 232.254 0.36 236.628 ; 
        RECT 62.212 236.574 62.724 240.948 ; 
        RECT 62.156 239.236 62.724 240.526 ; 
        RECT 61.276 238.144 61.812 240.948 ; 
        RECT 61.184 239.484 61.812 240.516 ; 
        RECT 61.276 236.574 61.668 240.948 ; 
        RECT 61.276 237.058 61.724 238.016 ; 
        RECT 61.276 236.574 61.812 236.93 ; 
        RECT 60.376 238.376 60.912 240.948 ; 
        RECT 60.376 236.574 60.768 240.948 ; 
        RECT 58.708 236.574 59.04 240.948 ; 
        RECT 58.708 236.928 59.096 240.67 ; 
        RECT 121.072 236.574 121.412 240.948 ; 
        RECT 120.496 236.574 120.6 240.948 ; 
        RECT 120.064 236.574 120.168 240.948 ; 
        RECT 119.632 236.574 119.736 240.948 ; 
        RECT 119.2 236.574 119.304 240.948 ; 
        RECT 118.768 236.574 118.872 240.948 ; 
        RECT 118.336 236.574 118.44 240.948 ; 
        RECT 117.904 236.574 118.008 240.948 ; 
        RECT 117.472 236.574 117.576 240.948 ; 
        RECT 117.04 236.574 117.144 240.948 ; 
        RECT 116.608 236.574 116.712 240.948 ; 
        RECT 116.176 236.574 116.28 240.948 ; 
        RECT 115.744 236.574 115.848 240.948 ; 
        RECT 115.312 236.574 115.416 240.948 ; 
        RECT 114.88 236.574 114.984 240.948 ; 
        RECT 114.448 236.574 114.552 240.948 ; 
        RECT 114.016 236.574 114.12 240.948 ; 
        RECT 113.584 236.574 113.688 240.948 ; 
        RECT 113.152 236.574 113.256 240.948 ; 
        RECT 112.72 236.574 112.824 240.948 ; 
        RECT 112.288 236.574 112.392 240.948 ; 
        RECT 111.856 236.574 111.96 240.948 ; 
        RECT 111.424 236.574 111.528 240.948 ; 
        RECT 110.992 236.574 111.096 240.948 ; 
        RECT 110.56 236.574 110.664 240.948 ; 
        RECT 110.128 236.574 110.232 240.948 ; 
        RECT 109.696 236.574 109.8 240.948 ; 
        RECT 109.264 236.574 109.368 240.948 ; 
        RECT 108.832 236.574 108.936 240.948 ; 
        RECT 108.4 236.574 108.504 240.948 ; 
        RECT 107.968 236.574 108.072 240.948 ; 
        RECT 107.536 236.574 107.64 240.948 ; 
        RECT 107.104 236.574 107.208 240.948 ; 
        RECT 106.672 236.574 106.776 240.948 ; 
        RECT 106.24 236.574 106.344 240.948 ; 
        RECT 105.808 236.574 105.912 240.948 ; 
        RECT 105.376 236.574 105.48 240.948 ; 
        RECT 104.944 236.574 105.048 240.948 ; 
        RECT 104.512 236.574 104.616 240.948 ; 
        RECT 104.08 236.574 104.184 240.948 ; 
        RECT 103.648 236.574 103.752 240.948 ; 
        RECT 103.216 236.574 103.32 240.948 ; 
        RECT 102.784 236.574 102.888 240.948 ; 
        RECT 102.352 236.574 102.456 240.948 ; 
        RECT 101.92 236.574 102.024 240.948 ; 
        RECT 101.488 236.574 101.592 240.948 ; 
        RECT 101.056 236.574 101.16 240.948 ; 
        RECT 100.624 236.574 100.728 240.948 ; 
        RECT 100.192 236.574 100.296 240.948 ; 
        RECT 99.76 236.574 99.864 240.948 ; 
        RECT 99.328 236.574 99.432 240.948 ; 
        RECT 98.896 236.574 99 240.948 ; 
        RECT 98.464 236.574 98.568 240.948 ; 
        RECT 98.032 236.574 98.136 240.948 ; 
        RECT 97.6 236.574 97.704 240.948 ; 
        RECT 97.168 236.574 97.272 240.948 ; 
        RECT 96.736 236.574 96.84 240.948 ; 
        RECT 96.304 236.574 96.408 240.948 ; 
        RECT 95.872 236.574 95.976 240.948 ; 
        RECT 95.44 236.574 95.544 240.948 ; 
        RECT 95.008 236.574 95.112 240.948 ; 
        RECT 94.576 236.574 94.68 240.948 ; 
        RECT 94.144 236.574 94.248 240.948 ; 
        RECT 93.712 236.574 93.816 240.948 ; 
        RECT 93.28 236.574 93.384 240.948 ; 
        RECT 92.848 236.574 92.952 240.948 ; 
        RECT 92.416 236.574 92.52 240.948 ; 
        RECT 91.984 236.574 92.088 240.948 ; 
        RECT 91.552 236.574 91.656 240.948 ; 
        RECT 91.12 236.574 91.224 240.948 ; 
        RECT 90.688 236.574 90.792 240.948 ; 
        RECT 90.256 236.574 90.36 240.948 ; 
        RECT 89.824 236.574 89.928 240.948 ; 
        RECT 89.392 236.574 89.496 240.948 ; 
        RECT 88.96 236.574 89.064 240.948 ; 
        RECT 88.528 236.574 88.632 240.948 ; 
        RECT 88.096 236.574 88.2 240.948 ; 
        RECT 87.664 236.574 87.768 240.948 ; 
        RECT 87.232 236.574 87.336 240.948 ; 
        RECT 86.8 236.574 86.904 240.948 ; 
        RECT 86.368 236.574 86.472 240.948 ; 
        RECT 85.936 236.574 86.04 240.948 ; 
        RECT 85.504 236.574 85.608 240.948 ; 
        RECT 85.072 236.574 85.176 240.948 ; 
        RECT 84.64 236.574 84.744 240.948 ; 
        RECT 84.208 236.574 84.312 240.948 ; 
        RECT 83.776 236.574 83.88 240.948 ; 
        RECT 83.344 236.574 83.448 240.948 ; 
        RECT 82.912 236.574 83.016 240.948 ; 
        RECT 82.48 236.574 82.584 240.948 ; 
        RECT 82.048 236.574 82.152 240.948 ; 
        RECT 81.616 236.574 81.72 240.948 ; 
        RECT 81.184 236.574 81.288 240.948 ; 
        RECT 80.752 236.574 80.856 240.948 ; 
        RECT 80.32 236.574 80.424 240.948 ; 
        RECT 79.888 236.574 79.992 240.948 ; 
        RECT 79.456 236.574 79.56 240.948 ; 
        RECT 79.024 236.574 79.128 240.948 ; 
        RECT 78.592 236.574 78.696 240.948 ; 
        RECT 78.16 236.574 78.264 240.948 ; 
        RECT 77.728 236.574 77.832 240.948 ; 
        RECT 77.296 236.574 77.4 240.948 ; 
        RECT 76.864 236.574 76.968 240.948 ; 
        RECT 76.432 236.574 76.536 240.948 ; 
        RECT 76 236.574 76.104 240.948 ; 
        RECT 75.568 236.574 75.672 240.948 ; 
        RECT 75.136 236.574 75.24 240.948 ; 
        RECT 74.704 236.574 74.808 240.948 ; 
        RECT 74.272 236.574 74.376 240.948 ; 
        RECT 73.84 236.574 73.944 240.948 ; 
        RECT 73.408 236.574 73.512 240.948 ; 
        RECT 72.976 236.574 73.08 240.948 ; 
        RECT 72.544 236.574 72.648 240.948 ; 
        RECT 72.112 236.574 72.216 240.948 ; 
        RECT 71.68 236.574 71.784 240.948 ; 
        RECT 71.248 236.574 71.352 240.948 ; 
        RECT 70.816 236.574 70.92 240.948 ; 
        RECT 70.384 236.574 70.488 240.948 ; 
        RECT 69.952 236.574 70.056 240.948 ; 
        RECT 69.52 236.574 69.624 240.948 ; 
        RECT 69.088 236.574 69.192 240.948 ; 
        RECT 68.656 236.574 68.76 240.948 ; 
        RECT 68.224 236.574 68.328 240.948 ; 
        RECT 67.792 236.574 67.896 240.948 ; 
        RECT 67.36 236.574 67.464 240.948 ; 
        RECT 66.928 236.574 67.032 240.948 ; 
        RECT 66.496 236.574 66.6 240.948 ; 
        RECT 66.064 236.574 66.168 240.948 ; 
        RECT 65.632 236.574 65.736 240.948 ; 
        RECT 65.2 236.574 65.304 240.948 ; 
        RECT 64.348 236.574 64.656 240.948 ; 
        RECT 56.776 236.574 57.084 240.948 ; 
        RECT 56.128 236.574 56.232 240.948 ; 
        RECT 55.696 236.574 55.8 240.948 ; 
        RECT 55.264 236.574 55.368 240.948 ; 
        RECT 54.832 236.574 54.936 240.948 ; 
        RECT 54.4 236.574 54.504 240.948 ; 
        RECT 53.968 236.574 54.072 240.948 ; 
        RECT 53.536 236.574 53.64 240.948 ; 
        RECT 53.104 236.574 53.208 240.948 ; 
        RECT 52.672 236.574 52.776 240.948 ; 
        RECT 52.24 236.574 52.344 240.948 ; 
        RECT 51.808 236.574 51.912 240.948 ; 
        RECT 51.376 236.574 51.48 240.948 ; 
        RECT 50.944 236.574 51.048 240.948 ; 
        RECT 50.512 236.574 50.616 240.948 ; 
        RECT 50.08 236.574 50.184 240.948 ; 
        RECT 49.648 236.574 49.752 240.948 ; 
        RECT 49.216 236.574 49.32 240.948 ; 
        RECT 48.784 236.574 48.888 240.948 ; 
        RECT 48.352 236.574 48.456 240.948 ; 
        RECT 47.92 236.574 48.024 240.948 ; 
        RECT 47.488 236.574 47.592 240.948 ; 
        RECT 47.056 236.574 47.16 240.948 ; 
        RECT 46.624 236.574 46.728 240.948 ; 
        RECT 46.192 236.574 46.296 240.948 ; 
        RECT 45.76 236.574 45.864 240.948 ; 
        RECT 45.328 236.574 45.432 240.948 ; 
        RECT 44.896 236.574 45 240.948 ; 
        RECT 44.464 236.574 44.568 240.948 ; 
        RECT 44.032 236.574 44.136 240.948 ; 
        RECT 43.6 236.574 43.704 240.948 ; 
        RECT 43.168 236.574 43.272 240.948 ; 
        RECT 42.736 236.574 42.84 240.948 ; 
        RECT 42.304 236.574 42.408 240.948 ; 
        RECT 41.872 236.574 41.976 240.948 ; 
        RECT 41.44 236.574 41.544 240.948 ; 
        RECT 41.008 236.574 41.112 240.948 ; 
        RECT 40.576 236.574 40.68 240.948 ; 
        RECT 40.144 236.574 40.248 240.948 ; 
        RECT 39.712 236.574 39.816 240.948 ; 
        RECT 39.28 236.574 39.384 240.948 ; 
        RECT 38.848 236.574 38.952 240.948 ; 
        RECT 38.416 236.574 38.52 240.948 ; 
        RECT 37.984 236.574 38.088 240.948 ; 
        RECT 37.552 236.574 37.656 240.948 ; 
        RECT 37.12 236.574 37.224 240.948 ; 
        RECT 36.688 236.574 36.792 240.948 ; 
        RECT 36.256 236.574 36.36 240.948 ; 
        RECT 35.824 236.574 35.928 240.948 ; 
        RECT 35.392 236.574 35.496 240.948 ; 
        RECT 34.96 236.574 35.064 240.948 ; 
        RECT 34.528 236.574 34.632 240.948 ; 
        RECT 34.096 236.574 34.2 240.948 ; 
        RECT 33.664 236.574 33.768 240.948 ; 
        RECT 33.232 236.574 33.336 240.948 ; 
        RECT 32.8 236.574 32.904 240.948 ; 
        RECT 32.368 236.574 32.472 240.948 ; 
        RECT 31.936 236.574 32.04 240.948 ; 
        RECT 31.504 236.574 31.608 240.948 ; 
        RECT 31.072 236.574 31.176 240.948 ; 
        RECT 30.64 236.574 30.744 240.948 ; 
        RECT 30.208 236.574 30.312 240.948 ; 
        RECT 29.776 236.574 29.88 240.948 ; 
        RECT 29.344 236.574 29.448 240.948 ; 
        RECT 28.912 236.574 29.016 240.948 ; 
        RECT 28.48 236.574 28.584 240.948 ; 
        RECT 28.048 236.574 28.152 240.948 ; 
        RECT 27.616 236.574 27.72 240.948 ; 
        RECT 27.184 236.574 27.288 240.948 ; 
        RECT 26.752 236.574 26.856 240.948 ; 
        RECT 26.32 236.574 26.424 240.948 ; 
        RECT 25.888 236.574 25.992 240.948 ; 
        RECT 25.456 236.574 25.56 240.948 ; 
        RECT 25.024 236.574 25.128 240.948 ; 
        RECT 24.592 236.574 24.696 240.948 ; 
        RECT 24.16 236.574 24.264 240.948 ; 
        RECT 23.728 236.574 23.832 240.948 ; 
        RECT 23.296 236.574 23.4 240.948 ; 
        RECT 22.864 236.574 22.968 240.948 ; 
        RECT 22.432 236.574 22.536 240.948 ; 
        RECT 22 236.574 22.104 240.948 ; 
        RECT 21.568 236.574 21.672 240.948 ; 
        RECT 21.136 236.574 21.24 240.948 ; 
        RECT 20.704 236.574 20.808 240.948 ; 
        RECT 20.272 236.574 20.376 240.948 ; 
        RECT 19.84 236.574 19.944 240.948 ; 
        RECT 19.408 236.574 19.512 240.948 ; 
        RECT 18.976 236.574 19.08 240.948 ; 
        RECT 18.544 236.574 18.648 240.948 ; 
        RECT 18.112 236.574 18.216 240.948 ; 
        RECT 17.68 236.574 17.784 240.948 ; 
        RECT 17.248 236.574 17.352 240.948 ; 
        RECT 16.816 236.574 16.92 240.948 ; 
        RECT 16.384 236.574 16.488 240.948 ; 
        RECT 15.952 236.574 16.056 240.948 ; 
        RECT 15.52 236.574 15.624 240.948 ; 
        RECT 15.088 236.574 15.192 240.948 ; 
        RECT 14.656 236.574 14.76 240.948 ; 
        RECT 14.224 236.574 14.328 240.948 ; 
        RECT 13.792 236.574 13.896 240.948 ; 
        RECT 13.36 236.574 13.464 240.948 ; 
        RECT 12.928 236.574 13.032 240.948 ; 
        RECT 12.496 236.574 12.6 240.948 ; 
        RECT 12.064 236.574 12.168 240.948 ; 
        RECT 11.632 236.574 11.736 240.948 ; 
        RECT 11.2 236.574 11.304 240.948 ; 
        RECT 10.768 236.574 10.872 240.948 ; 
        RECT 10.336 236.574 10.44 240.948 ; 
        RECT 9.904 236.574 10.008 240.948 ; 
        RECT 9.472 236.574 9.576 240.948 ; 
        RECT 9.04 236.574 9.144 240.948 ; 
        RECT 8.608 236.574 8.712 240.948 ; 
        RECT 8.176 236.574 8.28 240.948 ; 
        RECT 7.744 236.574 7.848 240.948 ; 
        RECT 7.312 236.574 7.416 240.948 ; 
        RECT 6.88 236.574 6.984 240.948 ; 
        RECT 6.448 236.574 6.552 240.948 ; 
        RECT 6.016 236.574 6.12 240.948 ; 
        RECT 5.584 236.574 5.688 240.948 ; 
        RECT 5.152 236.574 5.256 240.948 ; 
        RECT 4.72 236.574 4.824 240.948 ; 
        RECT 4.288 236.574 4.392 240.948 ; 
        RECT 3.856 236.574 3.96 240.948 ; 
        RECT 3.424 236.574 3.528 240.948 ; 
        RECT 2.992 236.574 3.096 240.948 ; 
        RECT 2.56 236.574 2.664 240.948 ; 
        RECT 2.128 236.574 2.232 240.948 ; 
        RECT 1.696 236.574 1.8 240.948 ; 
        RECT 1.264 236.574 1.368 240.948 ; 
        RECT 0.832 236.574 0.936 240.948 ; 
        RECT 0.02 236.574 0.36 240.948 ; 
  LAYER V3 SPACING 0.072 ; 
      RECT 0.02 4.88 121.412 5.4 ; 
      RECT 120.944 1.026 121.412 5.4 ; 
      RECT 64.856 4.496 120.872 5.4 ; 
      RECT 59.528 4.496 64.784 5.4 ; 
      RECT 56.648 1.026 59.168 5.4 ; 
      RECT 0.56 4.496 56.576 5.4 ; 
      RECT 0.02 1.026 0.488 5.4 ; 
      RECT 120.8 1.026 121.412 4.688 ; 
      RECT 65.072 1.026 120.728 5.4 ; 
      RECT 62.084 1.026 65 4.688 ; 
      RECT 61.148 1.808 61.94 5.4 ; 
      RECT 56.432 1.424 61.04 4.688 ; 
      RECT 0.704 1.026 56.36 5.4 ; 
      RECT 0.02 1.026 0.632 4.688 ; 
      RECT 61.868 1.026 121.412 4.304 ; 
      RECT 0.02 1.424 61.796 4.304 ; 
      RECT 60.968 1.026 121.412 1.712 ; 
      RECT 0.02 1.026 60.896 4.304 ; 
      RECT 0.02 1.026 121.412 1.328 ; 
      RECT 0.02 9.2 121.412 9.72 ; 
      RECT 120.944 5.346 121.412 9.72 ; 
      RECT 64.856 8.816 120.872 9.72 ; 
      RECT 59.528 8.816 64.784 9.72 ; 
      RECT 56.648 5.346 59.168 9.72 ; 
      RECT 0.56 8.816 56.576 9.72 ; 
      RECT 0.02 5.346 0.488 9.72 ; 
      RECT 120.8 5.346 121.412 9.008 ; 
      RECT 65.072 5.346 120.728 9.72 ; 
      RECT 62.084 5.346 65 9.008 ; 
      RECT 61.148 6.128 61.94 9.72 ; 
      RECT 56.432 5.744 61.04 9.008 ; 
      RECT 0.704 5.346 56.36 9.72 ; 
      RECT 0.02 5.346 0.632 9.008 ; 
      RECT 61.868 5.346 121.412 8.624 ; 
      RECT 0.02 5.744 61.796 8.624 ; 
      RECT 60.968 5.346 121.412 6.032 ; 
      RECT 0.02 5.346 60.896 8.624 ; 
      RECT 0.02 5.346 121.412 5.648 ; 
      RECT 0.02 13.52 121.412 14.04 ; 
      RECT 120.944 9.666 121.412 14.04 ; 
      RECT 64.856 13.136 120.872 14.04 ; 
      RECT 59.528 13.136 64.784 14.04 ; 
      RECT 56.648 9.666 59.168 14.04 ; 
      RECT 0.56 13.136 56.576 14.04 ; 
      RECT 0.02 9.666 0.488 14.04 ; 
      RECT 120.8 9.666 121.412 13.328 ; 
      RECT 65.072 9.666 120.728 14.04 ; 
      RECT 62.084 9.666 65 13.328 ; 
      RECT 61.148 10.448 61.94 14.04 ; 
      RECT 56.432 10.064 61.04 13.328 ; 
      RECT 0.704 9.666 56.36 14.04 ; 
      RECT 0.02 9.666 0.632 13.328 ; 
      RECT 61.868 9.666 121.412 12.944 ; 
      RECT 0.02 10.064 61.796 12.944 ; 
      RECT 60.968 9.666 121.412 10.352 ; 
      RECT 0.02 9.666 60.896 12.944 ; 
      RECT 0.02 9.666 121.412 9.968 ; 
      RECT 0.02 17.84 121.412 18.36 ; 
      RECT 120.944 13.986 121.412 18.36 ; 
      RECT 64.856 17.456 120.872 18.36 ; 
      RECT 59.528 17.456 64.784 18.36 ; 
      RECT 56.648 13.986 59.168 18.36 ; 
      RECT 0.56 17.456 56.576 18.36 ; 
      RECT 0.02 13.986 0.488 18.36 ; 
      RECT 120.8 13.986 121.412 17.648 ; 
      RECT 65.072 13.986 120.728 18.36 ; 
      RECT 62.084 13.986 65 17.648 ; 
      RECT 61.148 14.768 61.94 18.36 ; 
      RECT 56.432 14.384 61.04 17.648 ; 
      RECT 0.704 13.986 56.36 18.36 ; 
      RECT 0.02 13.986 0.632 17.648 ; 
      RECT 61.868 13.986 121.412 17.264 ; 
      RECT 0.02 14.384 61.796 17.264 ; 
      RECT 60.968 13.986 121.412 14.672 ; 
      RECT 0.02 13.986 60.896 17.264 ; 
      RECT 0.02 13.986 121.412 14.288 ; 
      RECT 0.02 22.16 121.412 22.68 ; 
      RECT 120.944 18.306 121.412 22.68 ; 
      RECT 64.856 21.776 120.872 22.68 ; 
      RECT 59.528 21.776 64.784 22.68 ; 
      RECT 56.648 18.306 59.168 22.68 ; 
      RECT 0.56 21.776 56.576 22.68 ; 
      RECT 0.02 18.306 0.488 22.68 ; 
      RECT 120.8 18.306 121.412 21.968 ; 
      RECT 65.072 18.306 120.728 22.68 ; 
      RECT 62.084 18.306 65 21.968 ; 
      RECT 61.148 19.088 61.94 22.68 ; 
      RECT 56.432 18.704 61.04 21.968 ; 
      RECT 0.704 18.306 56.36 22.68 ; 
      RECT 0.02 18.306 0.632 21.968 ; 
      RECT 61.868 18.306 121.412 21.584 ; 
      RECT 0.02 18.704 61.796 21.584 ; 
      RECT 60.968 18.306 121.412 18.992 ; 
      RECT 0.02 18.306 60.896 21.584 ; 
      RECT 0.02 18.306 121.412 18.608 ; 
      RECT 0.02 26.48 121.412 27 ; 
      RECT 120.944 22.626 121.412 27 ; 
      RECT 64.856 26.096 120.872 27 ; 
      RECT 59.528 26.096 64.784 27 ; 
      RECT 56.648 22.626 59.168 27 ; 
      RECT 0.56 26.096 56.576 27 ; 
      RECT 0.02 22.626 0.488 27 ; 
      RECT 120.8 22.626 121.412 26.288 ; 
      RECT 65.072 22.626 120.728 27 ; 
      RECT 62.084 22.626 65 26.288 ; 
      RECT 61.148 23.408 61.94 27 ; 
      RECT 56.432 23.024 61.04 26.288 ; 
      RECT 0.704 22.626 56.36 27 ; 
      RECT 0.02 22.626 0.632 26.288 ; 
      RECT 61.868 22.626 121.412 25.904 ; 
      RECT 0.02 23.024 61.796 25.904 ; 
      RECT 60.968 22.626 121.412 23.312 ; 
      RECT 0.02 22.626 60.896 25.904 ; 
      RECT 0.02 22.626 121.412 22.928 ; 
      RECT 0.02 30.8 121.412 31.32 ; 
      RECT 120.944 26.946 121.412 31.32 ; 
      RECT 64.856 30.416 120.872 31.32 ; 
      RECT 59.528 30.416 64.784 31.32 ; 
      RECT 56.648 26.946 59.168 31.32 ; 
      RECT 0.56 30.416 56.576 31.32 ; 
      RECT 0.02 26.946 0.488 31.32 ; 
      RECT 120.8 26.946 121.412 30.608 ; 
      RECT 65.072 26.946 120.728 31.32 ; 
      RECT 62.084 26.946 65 30.608 ; 
      RECT 61.148 27.728 61.94 31.32 ; 
      RECT 56.432 27.344 61.04 30.608 ; 
      RECT 0.704 26.946 56.36 31.32 ; 
      RECT 0.02 26.946 0.632 30.608 ; 
      RECT 61.868 26.946 121.412 30.224 ; 
      RECT 0.02 27.344 61.796 30.224 ; 
      RECT 60.968 26.946 121.412 27.632 ; 
      RECT 0.02 26.946 60.896 30.224 ; 
      RECT 0.02 26.946 121.412 27.248 ; 
      RECT 0.02 35.12 121.412 35.64 ; 
      RECT 120.944 31.266 121.412 35.64 ; 
      RECT 64.856 34.736 120.872 35.64 ; 
      RECT 59.528 34.736 64.784 35.64 ; 
      RECT 56.648 31.266 59.168 35.64 ; 
      RECT 0.56 34.736 56.576 35.64 ; 
      RECT 0.02 31.266 0.488 35.64 ; 
      RECT 120.8 31.266 121.412 34.928 ; 
      RECT 65.072 31.266 120.728 35.64 ; 
      RECT 62.084 31.266 65 34.928 ; 
      RECT 61.148 32.048 61.94 35.64 ; 
      RECT 56.432 31.664 61.04 34.928 ; 
      RECT 0.704 31.266 56.36 35.64 ; 
      RECT 0.02 31.266 0.632 34.928 ; 
      RECT 61.868 31.266 121.412 34.544 ; 
      RECT 0.02 31.664 61.796 34.544 ; 
      RECT 60.968 31.266 121.412 31.952 ; 
      RECT 0.02 31.266 60.896 34.544 ; 
      RECT 0.02 31.266 121.412 31.568 ; 
      RECT 0.02 39.44 121.412 39.96 ; 
      RECT 120.944 35.586 121.412 39.96 ; 
      RECT 64.856 39.056 120.872 39.96 ; 
      RECT 59.528 39.056 64.784 39.96 ; 
      RECT 56.648 35.586 59.168 39.96 ; 
      RECT 0.56 39.056 56.576 39.96 ; 
      RECT 0.02 35.586 0.488 39.96 ; 
      RECT 120.8 35.586 121.412 39.248 ; 
      RECT 65.072 35.586 120.728 39.96 ; 
      RECT 62.084 35.586 65 39.248 ; 
      RECT 61.148 36.368 61.94 39.96 ; 
      RECT 56.432 35.984 61.04 39.248 ; 
      RECT 0.704 35.586 56.36 39.96 ; 
      RECT 0.02 35.586 0.632 39.248 ; 
      RECT 61.868 35.586 121.412 38.864 ; 
      RECT 0.02 35.984 61.796 38.864 ; 
      RECT 60.968 35.586 121.412 36.272 ; 
      RECT 0.02 35.586 60.896 38.864 ; 
      RECT 0.02 35.586 121.412 35.888 ; 
      RECT 0.02 43.76 121.412 44.28 ; 
      RECT 120.944 39.906 121.412 44.28 ; 
      RECT 64.856 43.376 120.872 44.28 ; 
      RECT 59.528 43.376 64.784 44.28 ; 
      RECT 56.648 39.906 59.168 44.28 ; 
      RECT 0.56 43.376 56.576 44.28 ; 
      RECT 0.02 39.906 0.488 44.28 ; 
      RECT 120.8 39.906 121.412 43.568 ; 
      RECT 65.072 39.906 120.728 44.28 ; 
      RECT 62.084 39.906 65 43.568 ; 
      RECT 61.148 40.688 61.94 44.28 ; 
      RECT 56.432 40.304 61.04 43.568 ; 
      RECT 0.704 39.906 56.36 44.28 ; 
      RECT 0.02 39.906 0.632 43.568 ; 
      RECT 61.868 39.906 121.412 43.184 ; 
      RECT 0.02 40.304 61.796 43.184 ; 
      RECT 60.968 39.906 121.412 40.592 ; 
      RECT 0.02 39.906 60.896 43.184 ; 
      RECT 0.02 39.906 121.412 40.208 ; 
      RECT 0.02 48.08 121.412 48.6 ; 
      RECT 120.944 44.226 121.412 48.6 ; 
      RECT 64.856 47.696 120.872 48.6 ; 
      RECT 59.528 47.696 64.784 48.6 ; 
      RECT 56.648 44.226 59.168 48.6 ; 
      RECT 0.56 47.696 56.576 48.6 ; 
      RECT 0.02 44.226 0.488 48.6 ; 
      RECT 120.8 44.226 121.412 47.888 ; 
      RECT 65.072 44.226 120.728 48.6 ; 
      RECT 62.084 44.226 65 47.888 ; 
      RECT 61.148 45.008 61.94 48.6 ; 
      RECT 56.432 44.624 61.04 47.888 ; 
      RECT 0.704 44.226 56.36 48.6 ; 
      RECT 0.02 44.226 0.632 47.888 ; 
      RECT 61.868 44.226 121.412 47.504 ; 
      RECT 0.02 44.624 61.796 47.504 ; 
      RECT 60.968 44.226 121.412 44.912 ; 
      RECT 0.02 44.226 60.896 47.504 ; 
      RECT 0.02 44.226 121.412 44.528 ; 
      RECT 0.02 52.4 121.412 52.92 ; 
      RECT 120.944 48.546 121.412 52.92 ; 
      RECT 64.856 52.016 120.872 52.92 ; 
      RECT 59.528 52.016 64.784 52.92 ; 
      RECT 56.648 48.546 59.168 52.92 ; 
      RECT 0.56 52.016 56.576 52.92 ; 
      RECT 0.02 48.546 0.488 52.92 ; 
      RECT 120.8 48.546 121.412 52.208 ; 
      RECT 65.072 48.546 120.728 52.92 ; 
      RECT 62.084 48.546 65 52.208 ; 
      RECT 61.148 49.328 61.94 52.92 ; 
      RECT 56.432 48.944 61.04 52.208 ; 
      RECT 0.704 48.546 56.36 52.92 ; 
      RECT 0.02 48.546 0.632 52.208 ; 
      RECT 61.868 48.546 121.412 51.824 ; 
      RECT 0.02 48.944 61.796 51.824 ; 
      RECT 60.968 48.546 121.412 49.232 ; 
      RECT 0.02 48.546 60.896 51.824 ; 
      RECT 0.02 48.546 121.412 48.848 ; 
      RECT 0.02 56.72 121.412 57.24 ; 
      RECT 120.944 52.866 121.412 57.24 ; 
      RECT 64.856 56.336 120.872 57.24 ; 
      RECT 59.528 56.336 64.784 57.24 ; 
      RECT 56.648 52.866 59.168 57.24 ; 
      RECT 0.56 56.336 56.576 57.24 ; 
      RECT 0.02 52.866 0.488 57.24 ; 
      RECT 120.8 52.866 121.412 56.528 ; 
      RECT 65.072 52.866 120.728 57.24 ; 
      RECT 62.084 52.866 65 56.528 ; 
      RECT 61.148 53.648 61.94 57.24 ; 
      RECT 56.432 53.264 61.04 56.528 ; 
      RECT 0.704 52.866 56.36 57.24 ; 
      RECT 0.02 52.866 0.632 56.528 ; 
      RECT 61.868 52.866 121.412 56.144 ; 
      RECT 0.02 53.264 61.796 56.144 ; 
      RECT 60.968 52.866 121.412 53.552 ; 
      RECT 0.02 52.866 60.896 56.144 ; 
      RECT 0.02 52.866 121.412 53.168 ; 
      RECT 0.02 61.04 121.412 61.56 ; 
      RECT 120.944 57.186 121.412 61.56 ; 
      RECT 64.856 60.656 120.872 61.56 ; 
      RECT 59.528 60.656 64.784 61.56 ; 
      RECT 56.648 57.186 59.168 61.56 ; 
      RECT 0.56 60.656 56.576 61.56 ; 
      RECT 0.02 57.186 0.488 61.56 ; 
      RECT 120.8 57.186 121.412 60.848 ; 
      RECT 65.072 57.186 120.728 61.56 ; 
      RECT 62.084 57.186 65 60.848 ; 
      RECT 61.148 57.968 61.94 61.56 ; 
      RECT 56.432 57.584 61.04 60.848 ; 
      RECT 0.704 57.186 56.36 61.56 ; 
      RECT 0.02 57.186 0.632 60.848 ; 
      RECT 61.868 57.186 121.412 60.464 ; 
      RECT 0.02 57.584 61.796 60.464 ; 
      RECT 60.968 57.186 121.412 57.872 ; 
      RECT 0.02 57.186 60.896 60.464 ; 
      RECT 0.02 57.186 121.412 57.488 ; 
      RECT 0.02 65.36 121.412 65.88 ; 
      RECT 120.944 61.506 121.412 65.88 ; 
      RECT 64.856 64.976 120.872 65.88 ; 
      RECT 59.528 64.976 64.784 65.88 ; 
      RECT 56.648 61.506 59.168 65.88 ; 
      RECT 0.56 64.976 56.576 65.88 ; 
      RECT 0.02 61.506 0.488 65.88 ; 
      RECT 120.8 61.506 121.412 65.168 ; 
      RECT 65.072 61.506 120.728 65.88 ; 
      RECT 62.084 61.506 65 65.168 ; 
      RECT 61.148 62.288 61.94 65.88 ; 
      RECT 56.432 61.904 61.04 65.168 ; 
      RECT 0.704 61.506 56.36 65.88 ; 
      RECT 0.02 61.506 0.632 65.168 ; 
      RECT 61.868 61.506 121.412 64.784 ; 
      RECT 0.02 61.904 61.796 64.784 ; 
      RECT 60.968 61.506 121.412 62.192 ; 
      RECT 0.02 61.506 60.896 64.784 ; 
      RECT 0.02 61.506 121.412 61.808 ; 
      RECT 0.02 69.68 121.412 70.2 ; 
      RECT 120.944 65.826 121.412 70.2 ; 
      RECT 64.856 69.296 120.872 70.2 ; 
      RECT 59.528 69.296 64.784 70.2 ; 
      RECT 56.648 65.826 59.168 70.2 ; 
      RECT 0.56 69.296 56.576 70.2 ; 
      RECT 0.02 65.826 0.488 70.2 ; 
      RECT 120.8 65.826 121.412 69.488 ; 
      RECT 65.072 65.826 120.728 70.2 ; 
      RECT 62.084 65.826 65 69.488 ; 
      RECT 61.148 66.608 61.94 70.2 ; 
      RECT 56.432 66.224 61.04 69.488 ; 
      RECT 0.704 65.826 56.36 70.2 ; 
      RECT 0.02 65.826 0.632 69.488 ; 
      RECT 61.868 65.826 121.412 69.104 ; 
      RECT 0.02 66.224 61.796 69.104 ; 
      RECT 60.968 65.826 121.412 66.512 ; 
      RECT 0.02 65.826 60.896 69.104 ; 
      RECT 0.02 65.826 121.412 66.128 ; 
      RECT 0.02 74 121.412 74.52 ; 
      RECT 120.944 70.146 121.412 74.52 ; 
      RECT 64.856 73.616 120.872 74.52 ; 
      RECT 59.528 73.616 64.784 74.52 ; 
      RECT 56.648 70.146 59.168 74.52 ; 
      RECT 0.56 73.616 56.576 74.52 ; 
      RECT 0.02 70.146 0.488 74.52 ; 
      RECT 120.8 70.146 121.412 73.808 ; 
      RECT 65.072 70.146 120.728 74.52 ; 
      RECT 62.084 70.146 65 73.808 ; 
      RECT 61.148 70.928 61.94 74.52 ; 
      RECT 56.432 70.544 61.04 73.808 ; 
      RECT 0.704 70.146 56.36 74.52 ; 
      RECT 0.02 70.146 0.632 73.808 ; 
      RECT 61.868 70.146 121.412 73.424 ; 
      RECT 0.02 70.544 61.796 73.424 ; 
      RECT 60.968 70.146 121.412 70.832 ; 
      RECT 0.02 70.146 60.896 73.424 ; 
      RECT 0.02 70.146 121.412 70.448 ; 
      RECT 0.02 78.32 121.412 78.84 ; 
      RECT 120.944 74.466 121.412 78.84 ; 
      RECT 64.856 77.936 120.872 78.84 ; 
      RECT 59.528 77.936 64.784 78.84 ; 
      RECT 56.648 74.466 59.168 78.84 ; 
      RECT 0.56 77.936 56.576 78.84 ; 
      RECT 0.02 74.466 0.488 78.84 ; 
      RECT 120.8 74.466 121.412 78.128 ; 
      RECT 65.072 74.466 120.728 78.84 ; 
      RECT 62.084 74.466 65 78.128 ; 
      RECT 61.148 75.248 61.94 78.84 ; 
      RECT 56.432 74.864 61.04 78.128 ; 
      RECT 0.704 74.466 56.36 78.84 ; 
      RECT 0.02 74.466 0.632 78.128 ; 
      RECT 61.868 74.466 121.412 77.744 ; 
      RECT 0.02 74.864 61.796 77.744 ; 
      RECT 60.968 74.466 121.412 75.152 ; 
      RECT 0.02 74.466 60.896 77.744 ; 
      RECT 0.02 74.466 121.412 74.768 ; 
      RECT 0.02 82.64 121.412 83.16 ; 
      RECT 120.944 78.786 121.412 83.16 ; 
      RECT 64.856 82.256 120.872 83.16 ; 
      RECT 59.528 82.256 64.784 83.16 ; 
      RECT 56.648 78.786 59.168 83.16 ; 
      RECT 0.56 82.256 56.576 83.16 ; 
      RECT 0.02 78.786 0.488 83.16 ; 
      RECT 120.8 78.786 121.412 82.448 ; 
      RECT 65.072 78.786 120.728 83.16 ; 
      RECT 62.084 78.786 65 82.448 ; 
      RECT 61.148 79.568 61.94 83.16 ; 
      RECT 56.432 79.184 61.04 82.448 ; 
      RECT 0.704 78.786 56.36 83.16 ; 
      RECT 0.02 78.786 0.632 82.448 ; 
      RECT 61.868 78.786 121.412 82.064 ; 
      RECT 0.02 79.184 61.796 82.064 ; 
      RECT 60.968 78.786 121.412 79.472 ; 
      RECT 0.02 78.786 60.896 82.064 ; 
      RECT 0.02 78.786 121.412 79.088 ; 
      RECT 0.02 86.96 121.412 87.48 ; 
      RECT 120.944 83.106 121.412 87.48 ; 
      RECT 64.856 86.576 120.872 87.48 ; 
      RECT 59.528 86.576 64.784 87.48 ; 
      RECT 56.648 83.106 59.168 87.48 ; 
      RECT 0.56 86.576 56.576 87.48 ; 
      RECT 0.02 83.106 0.488 87.48 ; 
      RECT 120.8 83.106 121.412 86.768 ; 
      RECT 65.072 83.106 120.728 87.48 ; 
      RECT 62.084 83.106 65 86.768 ; 
      RECT 61.148 83.888 61.94 87.48 ; 
      RECT 56.432 83.504 61.04 86.768 ; 
      RECT 0.704 83.106 56.36 87.48 ; 
      RECT 0.02 83.106 0.632 86.768 ; 
      RECT 61.868 83.106 121.412 86.384 ; 
      RECT 0.02 83.504 61.796 86.384 ; 
      RECT 60.968 83.106 121.412 83.792 ; 
      RECT 0.02 83.106 60.896 86.384 ; 
      RECT 0.02 83.106 121.412 83.408 ; 
      RECT 0.02 91.28 121.412 91.8 ; 
      RECT 120.944 87.426 121.412 91.8 ; 
      RECT 64.856 90.896 120.872 91.8 ; 
      RECT 59.528 90.896 64.784 91.8 ; 
      RECT 56.648 87.426 59.168 91.8 ; 
      RECT 0.56 90.896 56.576 91.8 ; 
      RECT 0.02 87.426 0.488 91.8 ; 
      RECT 120.8 87.426 121.412 91.088 ; 
      RECT 65.072 87.426 120.728 91.8 ; 
      RECT 62.084 87.426 65 91.088 ; 
      RECT 61.148 88.208 61.94 91.8 ; 
      RECT 56.432 87.824 61.04 91.088 ; 
      RECT 0.704 87.426 56.36 91.8 ; 
      RECT 0.02 87.426 0.632 91.088 ; 
      RECT 61.868 87.426 121.412 90.704 ; 
      RECT 0.02 87.824 61.796 90.704 ; 
      RECT 60.968 87.426 121.412 88.112 ; 
      RECT 0.02 87.426 60.896 90.704 ; 
      RECT 0.02 87.426 121.412 87.728 ; 
      RECT 0.02 95.6 121.412 96.12 ; 
      RECT 120.944 91.746 121.412 96.12 ; 
      RECT 64.856 95.216 120.872 96.12 ; 
      RECT 59.528 95.216 64.784 96.12 ; 
      RECT 56.648 91.746 59.168 96.12 ; 
      RECT 0.56 95.216 56.576 96.12 ; 
      RECT 0.02 91.746 0.488 96.12 ; 
      RECT 120.8 91.746 121.412 95.408 ; 
      RECT 65.072 91.746 120.728 96.12 ; 
      RECT 62.084 91.746 65 95.408 ; 
      RECT 61.148 92.528 61.94 96.12 ; 
      RECT 56.432 92.144 61.04 95.408 ; 
      RECT 0.704 91.746 56.36 96.12 ; 
      RECT 0.02 91.746 0.632 95.408 ; 
      RECT 61.868 91.746 121.412 95.024 ; 
      RECT 0.02 92.144 61.796 95.024 ; 
      RECT 60.968 91.746 121.412 92.432 ; 
      RECT 0.02 91.746 60.896 95.024 ; 
      RECT 0.02 91.746 121.412 92.048 ; 
      RECT 0.02 99.92 121.412 100.44 ; 
      RECT 120.944 96.066 121.412 100.44 ; 
      RECT 64.856 99.536 120.872 100.44 ; 
      RECT 59.528 99.536 64.784 100.44 ; 
      RECT 56.648 96.066 59.168 100.44 ; 
      RECT 0.56 99.536 56.576 100.44 ; 
      RECT 0.02 96.066 0.488 100.44 ; 
      RECT 120.8 96.066 121.412 99.728 ; 
      RECT 65.072 96.066 120.728 100.44 ; 
      RECT 62.084 96.066 65 99.728 ; 
      RECT 61.148 96.848 61.94 100.44 ; 
      RECT 56.432 96.464 61.04 99.728 ; 
      RECT 0.704 96.066 56.36 100.44 ; 
      RECT 0.02 96.066 0.632 99.728 ; 
      RECT 61.868 96.066 121.412 99.344 ; 
      RECT 0.02 96.464 61.796 99.344 ; 
      RECT 60.968 96.066 121.412 96.752 ; 
      RECT 0.02 96.066 60.896 99.344 ; 
      RECT 0.02 96.066 121.412 96.368 ; 
      RECT 0.02 104.24 121.412 104.76 ; 
      RECT 120.944 100.386 121.412 104.76 ; 
      RECT 64.856 103.856 120.872 104.76 ; 
      RECT 59.528 103.856 64.784 104.76 ; 
      RECT 56.648 100.386 59.168 104.76 ; 
      RECT 0.56 103.856 56.576 104.76 ; 
      RECT 0.02 100.386 0.488 104.76 ; 
      RECT 120.8 100.386 121.412 104.048 ; 
      RECT 65.072 100.386 120.728 104.76 ; 
      RECT 62.084 100.386 65 104.048 ; 
      RECT 61.148 101.168 61.94 104.76 ; 
      RECT 56.432 100.784 61.04 104.048 ; 
      RECT 0.704 100.386 56.36 104.76 ; 
      RECT 0.02 100.386 0.632 104.048 ; 
      RECT 61.868 100.386 121.412 103.664 ; 
      RECT 0.02 100.784 61.796 103.664 ; 
      RECT 60.968 100.386 121.412 101.072 ; 
      RECT 0.02 100.386 60.896 103.664 ; 
      RECT 0.02 100.386 121.412 100.688 ; 
      RECT 0 134.134 121.392 139.468 ; 
      RECT 70.884 104.854 121.392 139.468 ; 
      RECT 62.084 110.71 121.392 139.468 ; 
      RECT 65.7 109.942 121.392 139.468 ; 
      RECT 61.876 104.854 62.012 139.468 ; 
      RECT 61.668 104.854 61.804 139.468 ; 
      RECT 61.46 104.854 61.596 139.468 ; 
      RECT 61.252 104.854 61.388 139.468 ; 
      RECT 0 111.094 61.18 139.468 ; 
      RECT 0 121.462 121.392 133.27 ; 
      RECT 56.628 108.79 63.324 120.598 ; 
      RECT 0 109.942 56.556 139.468 ; 
      RECT 0 110.326 65.628 110.998 ; 
      RECT 64.836 109.942 121.392 110.614 ; 
      RECT 0 109.942 64.764 110.998 ; 
      RECT 70.02 104.854 70.812 139.468 ; 
      RECT 54.9 109.174 69.948 110.23 ; 
      RECT 51.444 107.638 54.828 139.468 ; 
      RECT 0 104.854 51.372 139.468 ; 
      RECT 69.156 104.854 121.392 109.846 ; 
      RECT 68.292 107.638 121.392 109.846 ; 
      RECT 63.396 108.79 68.22 110.23 ; 
      RECT 0 108.79 63.324 109.846 ; 
      RECT 67.428 104.854 69.084 109.078 ; 
      RECT 65.052 107.638 121.392 109.078 ; 
      RECT 62.084 107.638 64.98 109.078 ; 
      RECT 56.412 107.638 61.18 110.998 ; 
      RECT 0 107.638 56.34 109.846 ; 
      RECT 62.244 107.446 67.356 107.926 ; 
      RECT 57.492 107.446 62.172 107.926 ; 
      RECT 54.036 107.446 57.42 107.926 ; 
      RECT 52.308 107.446 53.964 139.468 ; 
      RECT 0 104.854 52.236 109.846 ; 
      RECT 66.564 104.854 121.392 107.542 ; 
      RECT 60.66 104.854 66.492 107.542 ; 
      RECT 56.772 104.854 60.588 107.542 ; 
      RECT 53.172 104.854 56.7 107.542 ; 
      RECT 0 104.854 53.1 107.542 ; 
      RECT 0 104.854 121.392 107.35 ; 
        RECT 0.02 141.068 121.412 141.588 ; 
        RECT 120.944 137.214 121.412 141.588 ; 
        RECT 64.856 140.684 120.872 141.588 ; 
        RECT 59.528 140.684 64.784 141.588 ; 
        RECT 56.648 137.214 59.168 141.588 ; 
        RECT 0.56 140.684 56.576 141.588 ; 
        RECT 0.02 137.214 0.488 141.588 ; 
        RECT 120.8 137.214 121.412 140.876 ; 
        RECT 65.072 137.214 120.728 141.588 ; 
        RECT 62.084 137.214 65 140.876 ; 
        RECT 61.148 137.996 61.94 141.588 ; 
        RECT 56.432 137.612 61.04 140.876 ; 
        RECT 0.704 137.214 56.36 141.588 ; 
        RECT 0.02 137.214 0.632 140.876 ; 
        RECT 61.868 137.214 121.412 140.492 ; 
        RECT 0.02 137.612 61.796 140.492 ; 
        RECT 60.968 137.214 121.412 137.9 ; 
        RECT 0.02 137.214 60.896 140.492 ; 
        RECT 0.02 137.214 121.412 137.516 ; 
        RECT 0.02 145.388 121.412 145.908 ; 
        RECT 120.944 141.534 121.412 145.908 ; 
        RECT 64.856 145.004 120.872 145.908 ; 
        RECT 59.528 145.004 64.784 145.908 ; 
        RECT 56.648 141.534 59.168 145.908 ; 
        RECT 0.56 145.004 56.576 145.908 ; 
        RECT 0.02 141.534 0.488 145.908 ; 
        RECT 120.8 141.534 121.412 145.196 ; 
        RECT 65.072 141.534 120.728 145.908 ; 
        RECT 62.084 141.534 65 145.196 ; 
        RECT 61.148 142.316 61.94 145.908 ; 
        RECT 56.432 141.932 61.04 145.196 ; 
        RECT 0.704 141.534 56.36 145.908 ; 
        RECT 0.02 141.534 0.632 145.196 ; 
        RECT 61.868 141.534 121.412 144.812 ; 
        RECT 0.02 141.932 61.796 144.812 ; 
        RECT 60.968 141.534 121.412 142.22 ; 
        RECT 0.02 141.534 60.896 144.812 ; 
        RECT 0.02 141.534 121.412 141.836 ; 
        RECT 0.02 149.708 121.412 150.228 ; 
        RECT 120.944 145.854 121.412 150.228 ; 
        RECT 64.856 149.324 120.872 150.228 ; 
        RECT 59.528 149.324 64.784 150.228 ; 
        RECT 56.648 145.854 59.168 150.228 ; 
        RECT 0.56 149.324 56.576 150.228 ; 
        RECT 0.02 145.854 0.488 150.228 ; 
        RECT 120.8 145.854 121.412 149.516 ; 
        RECT 65.072 145.854 120.728 150.228 ; 
        RECT 62.084 145.854 65 149.516 ; 
        RECT 61.148 146.636 61.94 150.228 ; 
        RECT 56.432 146.252 61.04 149.516 ; 
        RECT 0.704 145.854 56.36 150.228 ; 
        RECT 0.02 145.854 0.632 149.516 ; 
        RECT 61.868 145.854 121.412 149.132 ; 
        RECT 0.02 146.252 61.796 149.132 ; 
        RECT 60.968 145.854 121.412 146.54 ; 
        RECT 0.02 145.854 60.896 149.132 ; 
        RECT 0.02 145.854 121.412 146.156 ; 
        RECT 0.02 154.028 121.412 154.548 ; 
        RECT 120.944 150.174 121.412 154.548 ; 
        RECT 64.856 153.644 120.872 154.548 ; 
        RECT 59.528 153.644 64.784 154.548 ; 
        RECT 56.648 150.174 59.168 154.548 ; 
        RECT 0.56 153.644 56.576 154.548 ; 
        RECT 0.02 150.174 0.488 154.548 ; 
        RECT 120.8 150.174 121.412 153.836 ; 
        RECT 65.072 150.174 120.728 154.548 ; 
        RECT 62.084 150.174 65 153.836 ; 
        RECT 61.148 150.956 61.94 154.548 ; 
        RECT 56.432 150.572 61.04 153.836 ; 
        RECT 0.704 150.174 56.36 154.548 ; 
        RECT 0.02 150.174 0.632 153.836 ; 
        RECT 61.868 150.174 121.412 153.452 ; 
        RECT 0.02 150.572 61.796 153.452 ; 
        RECT 60.968 150.174 121.412 150.86 ; 
        RECT 0.02 150.174 60.896 153.452 ; 
        RECT 0.02 150.174 121.412 150.476 ; 
        RECT 0.02 158.348 121.412 158.868 ; 
        RECT 120.944 154.494 121.412 158.868 ; 
        RECT 64.856 157.964 120.872 158.868 ; 
        RECT 59.528 157.964 64.784 158.868 ; 
        RECT 56.648 154.494 59.168 158.868 ; 
        RECT 0.56 157.964 56.576 158.868 ; 
        RECT 0.02 154.494 0.488 158.868 ; 
        RECT 120.8 154.494 121.412 158.156 ; 
        RECT 65.072 154.494 120.728 158.868 ; 
        RECT 62.084 154.494 65 158.156 ; 
        RECT 61.148 155.276 61.94 158.868 ; 
        RECT 56.432 154.892 61.04 158.156 ; 
        RECT 0.704 154.494 56.36 158.868 ; 
        RECT 0.02 154.494 0.632 158.156 ; 
        RECT 61.868 154.494 121.412 157.772 ; 
        RECT 0.02 154.892 61.796 157.772 ; 
        RECT 60.968 154.494 121.412 155.18 ; 
        RECT 0.02 154.494 60.896 157.772 ; 
        RECT 0.02 154.494 121.412 154.796 ; 
        RECT 0.02 162.668 121.412 163.188 ; 
        RECT 120.944 158.814 121.412 163.188 ; 
        RECT 64.856 162.284 120.872 163.188 ; 
        RECT 59.528 162.284 64.784 163.188 ; 
        RECT 56.648 158.814 59.168 163.188 ; 
        RECT 0.56 162.284 56.576 163.188 ; 
        RECT 0.02 158.814 0.488 163.188 ; 
        RECT 120.8 158.814 121.412 162.476 ; 
        RECT 65.072 158.814 120.728 163.188 ; 
        RECT 62.084 158.814 65 162.476 ; 
        RECT 61.148 159.596 61.94 163.188 ; 
        RECT 56.432 159.212 61.04 162.476 ; 
        RECT 0.704 158.814 56.36 163.188 ; 
        RECT 0.02 158.814 0.632 162.476 ; 
        RECT 61.868 158.814 121.412 162.092 ; 
        RECT 0.02 159.212 61.796 162.092 ; 
        RECT 60.968 158.814 121.412 159.5 ; 
        RECT 0.02 158.814 60.896 162.092 ; 
        RECT 0.02 158.814 121.412 159.116 ; 
        RECT 0.02 166.988 121.412 167.508 ; 
        RECT 120.944 163.134 121.412 167.508 ; 
        RECT 64.856 166.604 120.872 167.508 ; 
        RECT 59.528 166.604 64.784 167.508 ; 
        RECT 56.648 163.134 59.168 167.508 ; 
        RECT 0.56 166.604 56.576 167.508 ; 
        RECT 0.02 163.134 0.488 167.508 ; 
        RECT 120.8 163.134 121.412 166.796 ; 
        RECT 65.072 163.134 120.728 167.508 ; 
        RECT 62.084 163.134 65 166.796 ; 
        RECT 61.148 163.916 61.94 167.508 ; 
        RECT 56.432 163.532 61.04 166.796 ; 
        RECT 0.704 163.134 56.36 167.508 ; 
        RECT 0.02 163.134 0.632 166.796 ; 
        RECT 61.868 163.134 121.412 166.412 ; 
        RECT 0.02 163.532 61.796 166.412 ; 
        RECT 60.968 163.134 121.412 163.82 ; 
        RECT 0.02 163.134 60.896 166.412 ; 
        RECT 0.02 163.134 121.412 163.436 ; 
        RECT 0.02 171.308 121.412 171.828 ; 
        RECT 120.944 167.454 121.412 171.828 ; 
        RECT 64.856 170.924 120.872 171.828 ; 
        RECT 59.528 170.924 64.784 171.828 ; 
        RECT 56.648 167.454 59.168 171.828 ; 
        RECT 0.56 170.924 56.576 171.828 ; 
        RECT 0.02 167.454 0.488 171.828 ; 
        RECT 120.8 167.454 121.412 171.116 ; 
        RECT 65.072 167.454 120.728 171.828 ; 
        RECT 62.084 167.454 65 171.116 ; 
        RECT 61.148 168.236 61.94 171.828 ; 
        RECT 56.432 167.852 61.04 171.116 ; 
        RECT 0.704 167.454 56.36 171.828 ; 
        RECT 0.02 167.454 0.632 171.116 ; 
        RECT 61.868 167.454 121.412 170.732 ; 
        RECT 0.02 167.852 61.796 170.732 ; 
        RECT 60.968 167.454 121.412 168.14 ; 
        RECT 0.02 167.454 60.896 170.732 ; 
        RECT 0.02 167.454 121.412 167.756 ; 
        RECT 0.02 175.628 121.412 176.148 ; 
        RECT 120.944 171.774 121.412 176.148 ; 
        RECT 64.856 175.244 120.872 176.148 ; 
        RECT 59.528 175.244 64.784 176.148 ; 
        RECT 56.648 171.774 59.168 176.148 ; 
        RECT 0.56 175.244 56.576 176.148 ; 
        RECT 0.02 171.774 0.488 176.148 ; 
        RECT 120.8 171.774 121.412 175.436 ; 
        RECT 65.072 171.774 120.728 176.148 ; 
        RECT 62.084 171.774 65 175.436 ; 
        RECT 61.148 172.556 61.94 176.148 ; 
        RECT 56.432 172.172 61.04 175.436 ; 
        RECT 0.704 171.774 56.36 176.148 ; 
        RECT 0.02 171.774 0.632 175.436 ; 
        RECT 61.868 171.774 121.412 175.052 ; 
        RECT 0.02 172.172 61.796 175.052 ; 
        RECT 60.968 171.774 121.412 172.46 ; 
        RECT 0.02 171.774 60.896 175.052 ; 
        RECT 0.02 171.774 121.412 172.076 ; 
        RECT 0.02 179.948 121.412 180.468 ; 
        RECT 120.944 176.094 121.412 180.468 ; 
        RECT 64.856 179.564 120.872 180.468 ; 
        RECT 59.528 179.564 64.784 180.468 ; 
        RECT 56.648 176.094 59.168 180.468 ; 
        RECT 0.56 179.564 56.576 180.468 ; 
        RECT 0.02 176.094 0.488 180.468 ; 
        RECT 120.8 176.094 121.412 179.756 ; 
        RECT 65.072 176.094 120.728 180.468 ; 
        RECT 62.084 176.094 65 179.756 ; 
        RECT 61.148 176.876 61.94 180.468 ; 
        RECT 56.432 176.492 61.04 179.756 ; 
        RECT 0.704 176.094 56.36 180.468 ; 
        RECT 0.02 176.094 0.632 179.756 ; 
        RECT 61.868 176.094 121.412 179.372 ; 
        RECT 0.02 176.492 61.796 179.372 ; 
        RECT 60.968 176.094 121.412 176.78 ; 
        RECT 0.02 176.094 60.896 179.372 ; 
        RECT 0.02 176.094 121.412 176.396 ; 
        RECT 0.02 184.268 121.412 184.788 ; 
        RECT 120.944 180.414 121.412 184.788 ; 
        RECT 64.856 183.884 120.872 184.788 ; 
        RECT 59.528 183.884 64.784 184.788 ; 
        RECT 56.648 180.414 59.168 184.788 ; 
        RECT 0.56 183.884 56.576 184.788 ; 
        RECT 0.02 180.414 0.488 184.788 ; 
        RECT 120.8 180.414 121.412 184.076 ; 
        RECT 65.072 180.414 120.728 184.788 ; 
        RECT 62.084 180.414 65 184.076 ; 
        RECT 61.148 181.196 61.94 184.788 ; 
        RECT 56.432 180.812 61.04 184.076 ; 
        RECT 0.704 180.414 56.36 184.788 ; 
        RECT 0.02 180.414 0.632 184.076 ; 
        RECT 61.868 180.414 121.412 183.692 ; 
        RECT 0.02 180.812 61.796 183.692 ; 
        RECT 60.968 180.414 121.412 181.1 ; 
        RECT 0.02 180.414 60.896 183.692 ; 
        RECT 0.02 180.414 121.412 180.716 ; 
        RECT 0.02 188.588 121.412 189.108 ; 
        RECT 120.944 184.734 121.412 189.108 ; 
        RECT 64.856 188.204 120.872 189.108 ; 
        RECT 59.528 188.204 64.784 189.108 ; 
        RECT 56.648 184.734 59.168 189.108 ; 
        RECT 0.56 188.204 56.576 189.108 ; 
        RECT 0.02 184.734 0.488 189.108 ; 
        RECT 120.8 184.734 121.412 188.396 ; 
        RECT 65.072 184.734 120.728 189.108 ; 
        RECT 62.084 184.734 65 188.396 ; 
        RECT 61.148 185.516 61.94 189.108 ; 
        RECT 56.432 185.132 61.04 188.396 ; 
        RECT 0.704 184.734 56.36 189.108 ; 
        RECT 0.02 184.734 0.632 188.396 ; 
        RECT 61.868 184.734 121.412 188.012 ; 
        RECT 0.02 185.132 61.796 188.012 ; 
        RECT 60.968 184.734 121.412 185.42 ; 
        RECT 0.02 184.734 60.896 188.012 ; 
        RECT 0.02 184.734 121.412 185.036 ; 
        RECT 0.02 192.908 121.412 193.428 ; 
        RECT 120.944 189.054 121.412 193.428 ; 
        RECT 64.856 192.524 120.872 193.428 ; 
        RECT 59.528 192.524 64.784 193.428 ; 
        RECT 56.648 189.054 59.168 193.428 ; 
        RECT 0.56 192.524 56.576 193.428 ; 
        RECT 0.02 189.054 0.488 193.428 ; 
        RECT 120.8 189.054 121.412 192.716 ; 
        RECT 65.072 189.054 120.728 193.428 ; 
        RECT 62.084 189.054 65 192.716 ; 
        RECT 61.148 189.836 61.94 193.428 ; 
        RECT 56.432 189.452 61.04 192.716 ; 
        RECT 0.704 189.054 56.36 193.428 ; 
        RECT 0.02 189.054 0.632 192.716 ; 
        RECT 61.868 189.054 121.412 192.332 ; 
        RECT 0.02 189.452 61.796 192.332 ; 
        RECT 60.968 189.054 121.412 189.74 ; 
        RECT 0.02 189.054 60.896 192.332 ; 
        RECT 0.02 189.054 121.412 189.356 ; 
        RECT 0.02 197.228 121.412 197.748 ; 
        RECT 120.944 193.374 121.412 197.748 ; 
        RECT 64.856 196.844 120.872 197.748 ; 
        RECT 59.528 196.844 64.784 197.748 ; 
        RECT 56.648 193.374 59.168 197.748 ; 
        RECT 0.56 196.844 56.576 197.748 ; 
        RECT 0.02 193.374 0.488 197.748 ; 
        RECT 120.8 193.374 121.412 197.036 ; 
        RECT 65.072 193.374 120.728 197.748 ; 
        RECT 62.084 193.374 65 197.036 ; 
        RECT 61.148 194.156 61.94 197.748 ; 
        RECT 56.432 193.772 61.04 197.036 ; 
        RECT 0.704 193.374 56.36 197.748 ; 
        RECT 0.02 193.374 0.632 197.036 ; 
        RECT 61.868 193.374 121.412 196.652 ; 
        RECT 0.02 193.772 61.796 196.652 ; 
        RECT 60.968 193.374 121.412 194.06 ; 
        RECT 0.02 193.374 60.896 196.652 ; 
        RECT 0.02 193.374 121.412 193.676 ; 
        RECT 0.02 201.548 121.412 202.068 ; 
        RECT 120.944 197.694 121.412 202.068 ; 
        RECT 64.856 201.164 120.872 202.068 ; 
        RECT 59.528 201.164 64.784 202.068 ; 
        RECT 56.648 197.694 59.168 202.068 ; 
        RECT 0.56 201.164 56.576 202.068 ; 
        RECT 0.02 197.694 0.488 202.068 ; 
        RECT 120.8 197.694 121.412 201.356 ; 
        RECT 65.072 197.694 120.728 202.068 ; 
        RECT 62.084 197.694 65 201.356 ; 
        RECT 61.148 198.476 61.94 202.068 ; 
        RECT 56.432 198.092 61.04 201.356 ; 
        RECT 0.704 197.694 56.36 202.068 ; 
        RECT 0.02 197.694 0.632 201.356 ; 
        RECT 61.868 197.694 121.412 200.972 ; 
        RECT 0.02 198.092 61.796 200.972 ; 
        RECT 60.968 197.694 121.412 198.38 ; 
        RECT 0.02 197.694 60.896 200.972 ; 
        RECT 0.02 197.694 121.412 197.996 ; 
        RECT 0.02 205.868 121.412 206.388 ; 
        RECT 120.944 202.014 121.412 206.388 ; 
        RECT 64.856 205.484 120.872 206.388 ; 
        RECT 59.528 205.484 64.784 206.388 ; 
        RECT 56.648 202.014 59.168 206.388 ; 
        RECT 0.56 205.484 56.576 206.388 ; 
        RECT 0.02 202.014 0.488 206.388 ; 
        RECT 120.8 202.014 121.412 205.676 ; 
        RECT 65.072 202.014 120.728 206.388 ; 
        RECT 62.084 202.014 65 205.676 ; 
        RECT 61.148 202.796 61.94 206.388 ; 
        RECT 56.432 202.412 61.04 205.676 ; 
        RECT 0.704 202.014 56.36 206.388 ; 
        RECT 0.02 202.014 0.632 205.676 ; 
        RECT 61.868 202.014 121.412 205.292 ; 
        RECT 0.02 202.412 61.796 205.292 ; 
        RECT 60.968 202.014 121.412 202.7 ; 
        RECT 0.02 202.014 60.896 205.292 ; 
        RECT 0.02 202.014 121.412 202.316 ; 
        RECT 0.02 210.188 121.412 210.708 ; 
        RECT 120.944 206.334 121.412 210.708 ; 
        RECT 64.856 209.804 120.872 210.708 ; 
        RECT 59.528 209.804 64.784 210.708 ; 
        RECT 56.648 206.334 59.168 210.708 ; 
        RECT 0.56 209.804 56.576 210.708 ; 
        RECT 0.02 206.334 0.488 210.708 ; 
        RECT 120.8 206.334 121.412 209.996 ; 
        RECT 65.072 206.334 120.728 210.708 ; 
        RECT 62.084 206.334 65 209.996 ; 
        RECT 61.148 207.116 61.94 210.708 ; 
        RECT 56.432 206.732 61.04 209.996 ; 
        RECT 0.704 206.334 56.36 210.708 ; 
        RECT 0.02 206.334 0.632 209.996 ; 
        RECT 61.868 206.334 121.412 209.612 ; 
        RECT 0.02 206.732 61.796 209.612 ; 
        RECT 60.968 206.334 121.412 207.02 ; 
        RECT 0.02 206.334 60.896 209.612 ; 
        RECT 0.02 206.334 121.412 206.636 ; 
        RECT 0.02 214.508 121.412 215.028 ; 
        RECT 120.944 210.654 121.412 215.028 ; 
        RECT 64.856 214.124 120.872 215.028 ; 
        RECT 59.528 214.124 64.784 215.028 ; 
        RECT 56.648 210.654 59.168 215.028 ; 
        RECT 0.56 214.124 56.576 215.028 ; 
        RECT 0.02 210.654 0.488 215.028 ; 
        RECT 120.8 210.654 121.412 214.316 ; 
        RECT 65.072 210.654 120.728 215.028 ; 
        RECT 62.084 210.654 65 214.316 ; 
        RECT 61.148 211.436 61.94 215.028 ; 
        RECT 56.432 211.052 61.04 214.316 ; 
        RECT 0.704 210.654 56.36 215.028 ; 
        RECT 0.02 210.654 0.632 214.316 ; 
        RECT 61.868 210.654 121.412 213.932 ; 
        RECT 0.02 211.052 61.796 213.932 ; 
        RECT 60.968 210.654 121.412 211.34 ; 
        RECT 0.02 210.654 60.896 213.932 ; 
        RECT 0.02 210.654 121.412 210.956 ; 
        RECT 0.02 218.828 121.412 219.348 ; 
        RECT 120.944 214.974 121.412 219.348 ; 
        RECT 64.856 218.444 120.872 219.348 ; 
        RECT 59.528 218.444 64.784 219.348 ; 
        RECT 56.648 214.974 59.168 219.348 ; 
        RECT 0.56 218.444 56.576 219.348 ; 
        RECT 0.02 214.974 0.488 219.348 ; 
        RECT 120.8 214.974 121.412 218.636 ; 
        RECT 65.072 214.974 120.728 219.348 ; 
        RECT 62.084 214.974 65 218.636 ; 
        RECT 61.148 215.756 61.94 219.348 ; 
        RECT 56.432 215.372 61.04 218.636 ; 
        RECT 0.704 214.974 56.36 219.348 ; 
        RECT 0.02 214.974 0.632 218.636 ; 
        RECT 61.868 214.974 121.412 218.252 ; 
        RECT 0.02 215.372 61.796 218.252 ; 
        RECT 60.968 214.974 121.412 215.66 ; 
        RECT 0.02 214.974 60.896 218.252 ; 
        RECT 0.02 214.974 121.412 215.276 ; 
        RECT 0.02 223.148 121.412 223.668 ; 
        RECT 120.944 219.294 121.412 223.668 ; 
        RECT 64.856 222.764 120.872 223.668 ; 
        RECT 59.528 222.764 64.784 223.668 ; 
        RECT 56.648 219.294 59.168 223.668 ; 
        RECT 0.56 222.764 56.576 223.668 ; 
        RECT 0.02 219.294 0.488 223.668 ; 
        RECT 120.8 219.294 121.412 222.956 ; 
        RECT 65.072 219.294 120.728 223.668 ; 
        RECT 62.084 219.294 65 222.956 ; 
        RECT 61.148 220.076 61.94 223.668 ; 
        RECT 56.432 219.692 61.04 222.956 ; 
        RECT 0.704 219.294 56.36 223.668 ; 
        RECT 0.02 219.294 0.632 222.956 ; 
        RECT 61.868 219.294 121.412 222.572 ; 
        RECT 0.02 219.692 61.796 222.572 ; 
        RECT 60.968 219.294 121.412 219.98 ; 
        RECT 0.02 219.294 60.896 222.572 ; 
        RECT 0.02 219.294 121.412 219.596 ; 
        RECT 0.02 227.468 121.412 227.988 ; 
        RECT 120.944 223.614 121.412 227.988 ; 
        RECT 64.856 227.084 120.872 227.988 ; 
        RECT 59.528 227.084 64.784 227.988 ; 
        RECT 56.648 223.614 59.168 227.988 ; 
        RECT 0.56 227.084 56.576 227.988 ; 
        RECT 0.02 223.614 0.488 227.988 ; 
        RECT 120.8 223.614 121.412 227.276 ; 
        RECT 65.072 223.614 120.728 227.988 ; 
        RECT 62.084 223.614 65 227.276 ; 
        RECT 61.148 224.396 61.94 227.988 ; 
        RECT 56.432 224.012 61.04 227.276 ; 
        RECT 0.704 223.614 56.36 227.988 ; 
        RECT 0.02 223.614 0.632 227.276 ; 
        RECT 61.868 223.614 121.412 226.892 ; 
        RECT 0.02 224.012 61.796 226.892 ; 
        RECT 60.968 223.614 121.412 224.3 ; 
        RECT 0.02 223.614 60.896 226.892 ; 
        RECT 0.02 223.614 121.412 223.916 ; 
        RECT 0.02 231.788 121.412 232.308 ; 
        RECT 120.944 227.934 121.412 232.308 ; 
        RECT 64.856 231.404 120.872 232.308 ; 
        RECT 59.528 231.404 64.784 232.308 ; 
        RECT 56.648 227.934 59.168 232.308 ; 
        RECT 0.56 231.404 56.576 232.308 ; 
        RECT 0.02 227.934 0.488 232.308 ; 
        RECT 120.8 227.934 121.412 231.596 ; 
        RECT 65.072 227.934 120.728 232.308 ; 
        RECT 62.084 227.934 65 231.596 ; 
        RECT 61.148 228.716 61.94 232.308 ; 
        RECT 56.432 228.332 61.04 231.596 ; 
        RECT 0.704 227.934 56.36 232.308 ; 
        RECT 0.02 227.934 0.632 231.596 ; 
        RECT 61.868 227.934 121.412 231.212 ; 
        RECT 0.02 228.332 61.796 231.212 ; 
        RECT 60.968 227.934 121.412 228.62 ; 
        RECT 0.02 227.934 60.896 231.212 ; 
        RECT 0.02 227.934 121.412 228.236 ; 
        RECT 0.02 236.108 121.412 236.628 ; 
        RECT 120.944 232.254 121.412 236.628 ; 
        RECT 64.856 235.724 120.872 236.628 ; 
        RECT 59.528 235.724 64.784 236.628 ; 
        RECT 56.648 232.254 59.168 236.628 ; 
        RECT 0.56 235.724 56.576 236.628 ; 
        RECT 0.02 232.254 0.488 236.628 ; 
        RECT 120.8 232.254 121.412 235.916 ; 
        RECT 65.072 232.254 120.728 236.628 ; 
        RECT 62.084 232.254 65 235.916 ; 
        RECT 61.148 233.036 61.94 236.628 ; 
        RECT 56.432 232.652 61.04 235.916 ; 
        RECT 0.704 232.254 56.36 236.628 ; 
        RECT 0.02 232.254 0.632 235.916 ; 
        RECT 61.868 232.254 121.412 235.532 ; 
        RECT 0.02 232.652 61.796 235.532 ; 
        RECT 60.968 232.254 121.412 232.94 ; 
        RECT 0.02 232.254 60.896 235.532 ; 
        RECT 0.02 232.254 121.412 232.556 ; 
        RECT 0.02 240.428 121.412 240.948 ; 
        RECT 120.944 236.574 121.412 240.948 ; 
        RECT 64.856 240.044 120.872 240.948 ; 
        RECT 59.528 240.044 64.784 240.948 ; 
        RECT 56.648 236.574 59.168 240.948 ; 
        RECT 0.56 240.044 56.576 240.948 ; 
        RECT 0.02 236.574 0.488 240.948 ; 
        RECT 120.8 236.574 121.412 240.236 ; 
        RECT 65.072 236.574 120.728 240.948 ; 
        RECT 62.084 236.574 65 240.236 ; 
        RECT 61.148 237.356 61.94 240.948 ; 
        RECT 56.432 236.972 61.04 240.236 ; 
        RECT 0.704 236.574 56.36 240.948 ; 
        RECT 0.02 236.574 0.632 240.236 ; 
        RECT 61.868 236.574 121.412 239.852 ; 
        RECT 0.02 236.972 61.796 239.852 ; 
        RECT 60.968 236.574 121.412 237.26 ; 
        RECT 0.02 236.574 60.896 239.852 ; 
        RECT 0.02 236.574 121.412 236.876 ; 
  LAYER M4 ; 
      RECT 6.4 111.706 115.342 111.802 ; 
      RECT 6.4 112.858 115.342 112.954 ; 
      RECT 6.4 114.394 115.342 114.49 ; 
      RECT 6.4 114.778 115.342 114.874 ; 
      RECT 6.4 116.122 115.342 116.218 ; 
      RECT 6.4 117.658 115.342 117.754 ; 
      RECT 6.4 118.042 115.342 118.138 ; 
      RECT 41.904 106.198 79.488 107.062 ; 
      RECT 71.468 107.542 71.804 107.638 ; 
      RECT 70.714 109.27 71.234 109.366 ; 
      RECT 70.748 113.05 71.216 113.146 ; 
      RECT 70.746 111.9 71.214 111.996 ; 
      RECT 68.15 109.27 70.434 109.366 ; 
      RECT 68.39 112.33 68.822 112.426 ; 
      RECT 63.1 113.878 67.472 113.974 ; 
      RECT 65.852 112.15 66.188 112.246 ; 
      RECT 62.716 116.95 66.188 117.046 ; 
      RECT 65.852 117.334 66.188 117.43 ; 
      RECT 65.14 110.23 65.476 110.326 ; 
      RECT 64.988 115.606 65.324 115.702 ; 
      RECT 64.988 118.486 65.324 118.582 ; 
      RECT 63.912 105.078 64.964 105.174 ; 
      RECT 64.436 120.214 64.884 120.31 ; 
      RECT 64.276 109.846 64.612 109.942 ; 
      RECT 63.42 104.694 64.472 104.79 ; 
      RECT 63.42 139.114 64.472 139.21 ; 
      RECT 63.484 115.798 64.46 115.894 ; 
      RECT 64.124 116.374 64.46 116.47 ; 
      RECT 58.3 117.334 64.46 117.43 ; 
      RECT 64.124 118.486 64.46 118.582 ; 
      RECT 63.188 138.73 64.24 138.826 ; 
      RECT 63.184 104.31 64.236 104.406 ; 
      RECT 57.24 118.87 64.152 119.734 ; 
      RECT 57.24 131.542 64.152 132.406 ; 
      RECT 63.032 103.926 64.084 104.022 ; 
      RECT 63.032 137.962 64.084 138.058 ; 
      RECT 63.692 120.214 64.028 120.31 ; 
      RECT 60.604 121.75 64.028 121.846 ; 
      RECT 62.14 130.774 64.028 130.87 ; 
      RECT 63.692 131.158 64.028 131.254 ; 
      RECT 62.84 103.542 63.892 103.638 ; 
      RECT 62.84 137.578 63.892 137.674 ; 
      RECT 61.948 127.126 63.728 127.222 ; 
      RECT 62.664 103.158 63.716 103.254 ; 
      RECT 62.664 138.922 63.716 139.018 ; 
      RECT 62.468 104.502 63.52 104.598 ; 
      RECT 62.468 138.538 63.52 138.634 ; 
      RECT 62.992 116.374 63.476 116.47 ; 
      RECT 62.908 124.822 63.44 124.918 ; 
      RECT 62.28 104.118 63.332 104.214 ; 
      RECT 62.28 138.154 63.332 138.25 ; 
      RECT 62.14 102.966 63.192 103.062 ; 
      RECT 62.14 137.77 63.192 137.866 ; 
      RECT 58.876 131.158 63.152 131.254 ; 
      RECT 62.816 135.766 63.152 135.862 ; 
      RECT 61.916 102.39 62.968 102.486 ; 
      RECT 61.916 137.386 62.968 137.482 ; 
      RECT 62.524 120.214 62.864 120.31 ; 
      RECT 58.108 122.518 62.576 122.614 ; 
      RECT 60.688 113.878 62.516 113.974 ; 
      RECT 59.996 105.27 61.064 105.366 ; 
      RECT 59.996 136.81 61.064 136.906 ; 
      RECT 60.544 120.022 60.98 120.118 ; 
      RECT 59.904 104.886 60.872 104.982 ; 
      RECT 59.904 139.306 60.872 139.402 ; 
      RECT 59.68 102.966 60.648 103.062 ; 
      RECT 59.796 139.69 60.648 139.786 ; 
      RECT 60.26 118.486 60.596 118.582 ; 
      RECT 59.464 103.35 60.456 103.446 ; 
      RECT 59.464 139.114 60.456 139.21 ; 
      RECT 58.528 128.854 60.212 128.95 ; 
      RECT 58.4 104.694 59.468 104.79 ; 
      RECT 58.4 139.69 59.468 139.786 ; 
      RECT 58.96 123.094 59.444 123.19 ; 
      RECT 58.928 135.766 59.264 135.862 ; 
      RECT 58.264 104.31 59.252 104.406 ; 
      RECT 57.996 137.962 59.252 138.058 ; 
      RECT 58.16 103.926 59.08 104.022 ; 
      RECT 58.112 139.306 59.08 139.402 ; 
      RECT 57.948 103.542 58.868 103.638 ; 
      RECT 58.532 129.43 58.868 129.526 ; 
      RECT 57.748 137.578 58.868 137.674 ; 
      RECT 57.768 103.158 58.688 103.254 ; 
      RECT 57.768 138.922 58.688 139.018 ; 
      RECT 53.92 118.486 58.676 118.582 ; 
      RECT 57.616 104.118 58.536 104.214 ; 
      RECT 57.616 138.538 58.536 138.634 ; 
      RECT 57.544 103.734 58.316 103.83 ; 
      RECT 57.544 138.154 58.316 138.25 ; 
      RECT 57.348 103.35 58.12 103.446 ; 
      RECT 57.348 137.77 58.12 137.866 ; 
      RECT 57.364 122.134 58.1 122.23 ; 
      RECT 57.14 102.966 57.912 103.062 ; 
      RECT 57.14 137.386 57.912 137.482 ; 
      RECT 55.204 111.382 57.908 111.478 ; 
      RECT 57.364 122.518 57.7 122.614 ; 
      RECT 56.288 105.078 57.34 105.174 ; 
      RECT 56.78 113.878 57.116 113.974 ; 
      RECT 56.504 120.214 56.952 120.31 ; 
      RECT 55.052 112.15 55.388 112.246 ; 
  LAYER V4 ; 
      RECT 71.664 107.542 71.76 107.638 ; 
      RECT 71.664 111.706 71.76 111.802 ; 
      RECT 70.992 111.9 71.088 111.996 ; 
      RECT 70.992 113.05 71.088 113.146 ; 
      RECT 70.99 109.27 71.086 109.366 ; 
      RECT 68.454 109.27 68.55 109.366 ; 
      RECT 68.454 112.33 68.55 112.426 ; 
      RECT 66.048 112.15 66.144 112.246 ; 
      RECT 66.048 112.858 66.144 112.954 ; 
      RECT 66.048 116.95 66.144 117.046 ; 
      RECT 66.048 117.334 66.144 117.43 ; 
      RECT 65.184 110.23 65.28 110.326 ; 
      RECT 65.184 114.394 65.28 114.49 ; 
      RECT 65.184 115.606 65.28 115.702 ; 
      RECT 65.184 116.122 65.28 116.218 ; 
      RECT 65.184 117.658 65.28 117.754 ; 
      RECT 65.184 118.486 65.28 118.582 ; 
      RECT 64.508 105.078 64.604 105.174 ; 
      RECT 64.512 106.198 64.604 107.062 ; 
      RECT 64.508 120.214 64.604 120.31 ; 
      RECT 64.32 109.846 64.416 109.942 ; 
      RECT 64.32 114.778 64.416 114.874 ; 
      RECT 64.32 115.798 64.416 115.894 ; 
      RECT 64.32 116.374 64.416 116.47 ; 
      RECT 64.32 117.334 64.416 117.43 ; 
      RECT 64.32 118.486 64.416 118.582 ; 
      RECT 63.888 120.214 63.984 120.31 ; 
      RECT 63.888 121.75 63.984 121.846 ; 
      RECT 63.888 130.774 63.984 130.87 ; 
      RECT 63.888 131.158 63.984 131.254 ; 
      RECT 63.528 104.694 63.624 104.79 ; 
      RECT 63.528 115.798 63.624 115.894 ; 
      RECT 63.528 139.114 63.624 139.21 ; 
      RECT 63.336 104.31 63.432 104.406 ; 
      RECT 63.336 116.374 63.432 116.47 ; 
      RECT 63.336 138.73 63.432 138.826 ; 
      RECT 63.144 103.926 63.24 104.022 ; 
      RECT 63.144 113.878 63.24 113.974 ; 
      RECT 63.144 137.962 63.24 138.058 ; 
      RECT 62.952 103.542 63.048 103.638 ; 
      RECT 62.952 124.822 63.048 124.918 ; 
      RECT 62.952 135.766 63.048 135.862 ; 
      RECT 62.952 137.578 63.048 137.674 ; 
      RECT 62.76 103.158 62.856 103.254 ; 
      RECT 62.76 116.95 62.856 117.046 ; 
      RECT 62.76 138.922 62.856 139.018 ; 
      RECT 62.568 104.502 62.664 104.598 ; 
      RECT 62.568 120.214 62.664 120.31 ; 
      RECT 62.568 138.538 62.664 138.634 ; 
      RECT 62.376 104.118 62.472 104.214 ; 
      RECT 62.376 113.878 62.472 113.974 ; 
      RECT 62.376 138.154 62.472 138.25 ; 
      RECT 62.184 102.966 62.28 103.062 ; 
      RECT 62.184 130.774 62.28 130.87 ; 
      RECT 62.184 137.77 62.28 137.866 ; 
      RECT 61.992 102.39 62.088 102.486 ; 
      RECT 61.992 127.126 62.088 127.222 ; 
      RECT 61.992 137.386 62.088 137.482 ; 
      RECT 60.84 105.27 60.936 105.366 ; 
      RECT 60.84 120.022 60.936 120.118 ; 
      RECT 60.84 136.81 60.936 136.906 ; 
      RECT 60.648 104.886 60.744 104.982 ; 
      RECT 60.648 121.75 60.744 121.846 ; 
      RECT 60.648 139.306 60.744 139.402 ; 
      RECT 60.456 102.966 60.552 103.062 ; 
      RECT 60.456 118.486 60.552 118.582 ; 
      RECT 60.456 139.69 60.552 139.786 ; 
      RECT 60.072 103.35 60.168 103.446 ; 
      RECT 60.072 128.854 60.168 128.95 ; 
      RECT 60.072 139.114 60.168 139.21 ; 
      RECT 59.304 104.694 59.4 104.79 ; 
      RECT 59.304 123.094 59.4 123.19 ; 
      RECT 59.304 139.69 59.4 139.786 ; 
      RECT 59.112 104.31 59.208 104.406 ; 
      RECT 59.112 135.766 59.208 135.862 ; 
      RECT 59.112 137.962 59.208 138.058 ; 
      RECT 58.92 103.926 59.016 104.022 ; 
      RECT 58.92 131.158 59.016 131.254 ; 
      RECT 58.92 139.306 59.016 139.402 ; 
      RECT 58.728 103.542 58.824 103.638 ; 
      RECT 58.728 129.43 58.824 129.526 ; 
      RECT 58.728 137.578 58.824 137.674 ; 
      RECT 58.536 103.158 58.632 103.254 ; 
      RECT 58.536 118.486 58.632 118.582 ; 
      RECT 58.536 138.922 58.632 139.018 ; 
      RECT 58.344 104.118 58.44 104.214 ; 
      RECT 58.344 117.334 58.44 117.43 ; 
      RECT 58.344 138.538 58.44 138.634 ; 
      RECT 58.152 103.734 58.248 103.83 ; 
      RECT 58.152 122.518 58.248 122.614 ; 
      RECT 58.152 138.154 58.248 138.25 ; 
      RECT 57.96 103.35 58.056 103.446 ; 
      RECT 57.96 122.134 58.056 122.23 ; 
      RECT 57.96 137.77 58.056 137.866 ; 
      RECT 57.768 102.966 57.864 103.062 ; 
      RECT 57.768 111.382 57.864 111.478 ; 
      RECT 57.768 137.386 57.864 137.482 ; 
      RECT 57.408 122.134 57.504 122.23 ; 
      RECT 57.408 122.518 57.504 122.614 ; 
      RECT 56.976 113.878 57.072 113.974 ; 
      RECT 56.976 118.042 57.072 118.138 ; 
      RECT 56.736 105.078 56.832 105.174 ; 
      RECT 56.74 106.198 56.832 107.062 ; 
      RECT 56.736 120.214 56.832 120.31 ; 
      RECT 55.248 111.382 55.344 111.478 ; 
      RECT 55.248 112.15 55.344 112.246 ; 
  LAYER M5 ; 
      RECT 71.664 107.498 71.76 111.846 ; 
      RECT 70.99 109.088 71.086 113.33 ; 
      RECT 68.454 109.104 68.55 112.588 ; 
      RECT 66.048 112.106 66.144 112.998 ; 
      RECT 66.048 116.906 66.144 117.474 ; 
      RECT 65.184 110.186 65.28 114.534 ; 
      RECT 65.184 115.562 65.28 116.262 ; 
      RECT 65.184 117.614 65.28 118.626 ; 
      RECT 64.508 105.006 64.604 120.382 ; 
      RECT 64.32 109.802 64.416 114.918 ; 
      RECT 64.32 115.754 64.416 116.514 ; 
      RECT 64.32 117.29 64.416 118.626 ; 
      RECT 63.888 120.17 63.984 121.89 ; 
      RECT 63.888 130.73 63.984 131.298 ; 
      RECT 63.528 102.084 63.624 140.09 ; 
      RECT 63.336 102.084 63.432 140.086 ; 
      RECT 63.144 102.084 63.24 140.086 ; 
      RECT 62.952 102.084 63.048 139.97 ; 
      RECT 62.76 102.084 62.856 139.958 ; 
      RECT 62.568 102.084 62.664 139.966 ; 
      RECT 62.376 102.084 62.472 139.938 ; 
      RECT 62.184 102.084 62.28 140.002 ; 
      RECT 61.992 102.084 62.088 139.998 ; 
      RECT 60.84 102.906 60.936 140.222 ; 
      RECT 60.648 102.91 60.744 140.226 ; 
      RECT 60.456 102.906 60.552 140.222 ; 
      RECT 60.072 102.97 60.168 140.226 ; 
      RECT 59.304 102.966 59.4 140.038 ; 
      RECT 59.112 102.966 59.208 140.038 ; 
      RECT 58.92 102.966 59.016 140.038 ; 
      RECT 58.728 102.966 58.824 140.038 ; 
      RECT 58.536 102.966 58.632 140.038 ; 
      RECT 58.344 102.85 58.44 140.038 ; 
      RECT 58.152 102.674 58.248 138.894 ; 
      RECT 57.96 102.526 58.056 138.71 ; 
      RECT 57.768 102.31 57.864 138.494 ; 
      RECT 57.408 122.09 57.504 122.658 ; 
      RECT 56.976 113.834 57.072 118.182 ; 
      RECT 56.736 105.006 56.832 120.382 ; 
      RECT 55.248 111.338 55.344 112.29 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 120.96 241.776 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 120.96 241.776 ; 
  END 
END srambank_256x4x48_6t122 
