VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_64x4x48_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_64x4x48_6t122 0 0 ; 
  SIZE 38.448 BY 241.92 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.688 38.036 4.88 ; 
        RECT 0.404 9.008 38.036 9.2 ; 
        RECT 0.404 13.328 38.036 13.52 ; 
        RECT 0.404 17.648 38.036 17.84 ; 
        RECT 0.404 21.968 38.036 22.16 ; 
        RECT 0.404 26.288 38.036 26.48 ; 
        RECT 0.404 30.608 38.036 30.8 ; 
        RECT 0.404 34.928 38.036 35.12 ; 
        RECT 0.404 39.248 38.036 39.44 ; 
        RECT 0.404 43.568 38.036 43.76 ; 
        RECT 0.404 47.888 38.036 48.08 ; 
        RECT 0.404 52.208 38.036 52.4 ; 
        RECT 0.404 56.528 38.036 56.72 ; 
        RECT 0.404 60.848 38.036 61.04 ; 
        RECT 0.404 65.168 38.036 65.36 ; 
        RECT 0.404 69.488 38.036 69.68 ; 
        RECT 0.404 73.808 38.036 74 ; 
        RECT 0.404 78.128 38.036 78.32 ; 
        RECT 0.404 82.448 38.036 82.64 ; 
        RECT 0.404 86.768 38.036 86.96 ; 
        RECT 0.404 91.088 38.036 91.28 ; 
        RECT 0.404 95.408 38.036 95.6 ; 
        RECT 0.404 99.728 38.036 99.92 ; 
        RECT 0.404 104.048 38.036 104.24 ; 
        RECT 0.432 105.996 38.016 106.86 ; 
        RECT 22.44 104.876 23.492 104.972 ; 
        RECT 22.964 120.012 23.412 120.108 ; 
        RECT 15.768 118.668 22.68 119.532 ; 
        RECT 15.768 131.34 22.68 132.204 ; 
        RECT 0.404 140.876 38.036 141.068 ; 
        RECT 0.404 145.196 38.036 145.388 ; 
        RECT 0.404 149.516 38.036 149.708 ; 
        RECT 0.404 153.836 38.036 154.028 ; 
        RECT 0.404 158.156 38.036 158.348 ; 
        RECT 0.404 162.476 38.036 162.668 ; 
        RECT 0.404 166.796 38.036 166.988 ; 
        RECT 0.404 171.116 38.036 171.308 ; 
        RECT 0.404 175.436 38.036 175.628 ; 
        RECT 0.404 179.756 38.036 179.948 ; 
        RECT 0.404 184.076 38.036 184.268 ; 
        RECT 0.404 188.396 38.036 188.588 ; 
        RECT 0.404 192.716 38.036 192.908 ; 
        RECT 0.404 197.036 38.036 197.228 ; 
        RECT 0.404 201.356 38.036 201.548 ; 
        RECT 0.404 205.676 38.036 205.868 ; 
        RECT 0.404 209.996 38.036 210.188 ; 
        RECT 0.404 214.316 38.036 214.508 ; 
        RECT 0.404 218.636 38.036 218.828 ; 
        RECT 0.404 222.956 38.036 223.148 ; 
        RECT 0.404 227.276 38.036 227.468 ; 
        RECT 0.404 231.596 38.036 231.788 ; 
        RECT 0.404 235.916 38.036 236.108 ; 
        RECT 0.404 240.236 38.036 240.428 ; 
      LAYER M3 ; 
        RECT 37.908 0.866 37.98 5.506 ; 
        RECT 23.292 0.868 23.364 5.504 ; 
        RECT 17.676 1.012 18.036 5.468 ; 
        RECT 15.084 0.868 15.156 5.504 ; 
        RECT 0.468 0.866 0.54 5.506 ; 
        RECT 37.908 5.186 37.98 9.826 ; 
        RECT 23.292 5.188 23.364 9.824 ; 
        RECT 17.676 5.332 18.036 9.788 ; 
        RECT 15.084 5.188 15.156 9.824 ; 
        RECT 0.468 5.186 0.54 9.826 ; 
        RECT 37.908 9.506 37.98 14.146 ; 
        RECT 23.292 9.508 23.364 14.144 ; 
        RECT 17.676 9.652 18.036 14.108 ; 
        RECT 15.084 9.508 15.156 14.144 ; 
        RECT 0.468 9.506 0.54 14.146 ; 
        RECT 37.908 13.826 37.98 18.466 ; 
        RECT 23.292 13.828 23.364 18.464 ; 
        RECT 17.676 13.972 18.036 18.428 ; 
        RECT 15.084 13.828 15.156 18.464 ; 
        RECT 0.468 13.826 0.54 18.466 ; 
        RECT 37.908 18.146 37.98 22.786 ; 
        RECT 23.292 18.148 23.364 22.784 ; 
        RECT 17.676 18.292 18.036 22.748 ; 
        RECT 15.084 18.148 15.156 22.784 ; 
        RECT 0.468 18.146 0.54 22.786 ; 
        RECT 37.908 22.466 37.98 27.106 ; 
        RECT 23.292 22.468 23.364 27.104 ; 
        RECT 17.676 22.612 18.036 27.068 ; 
        RECT 15.084 22.468 15.156 27.104 ; 
        RECT 0.468 22.466 0.54 27.106 ; 
        RECT 37.908 26.786 37.98 31.426 ; 
        RECT 23.292 26.788 23.364 31.424 ; 
        RECT 17.676 26.932 18.036 31.388 ; 
        RECT 15.084 26.788 15.156 31.424 ; 
        RECT 0.468 26.786 0.54 31.426 ; 
        RECT 37.908 31.106 37.98 35.746 ; 
        RECT 23.292 31.108 23.364 35.744 ; 
        RECT 17.676 31.252 18.036 35.708 ; 
        RECT 15.084 31.108 15.156 35.744 ; 
        RECT 0.468 31.106 0.54 35.746 ; 
        RECT 37.908 35.426 37.98 40.066 ; 
        RECT 23.292 35.428 23.364 40.064 ; 
        RECT 17.676 35.572 18.036 40.028 ; 
        RECT 15.084 35.428 15.156 40.064 ; 
        RECT 0.468 35.426 0.54 40.066 ; 
        RECT 37.908 39.746 37.98 44.386 ; 
        RECT 23.292 39.748 23.364 44.384 ; 
        RECT 17.676 39.892 18.036 44.348 ; 
        RECT 15.084 39.748 15.156 44.384 ; 
        RECT 0.468 39.746 0.54 44.386 ; 
        RECT 37.908 44.066 37.98 48.706 ; 
        RECT 23.292 44.068 23.364 48.704 ; 
        RECT 17.676 44.212 18.036 48.668 ; 
        RECT 15.084 44.068 15.156 48.704 ; 
        RECT 0.468 44.066 0.54 48.706 ; 
        RECT 37.908 48.386 37.98 53.026 ; 
        RECT 23.292 48.388 23.364 53.024 ; 
        RECT 17.676 48.532 18.036 52.988 ; 
        RECT 15.084 48.388 15.156 53.024 ; 
        RECT 0.468 48.386 0.54 53.026 ; 
        RECT 37.908 52.706 37.98 57.346 ; 
        RECT 23.292 52.708 23.364 57.344 ; 
        RECT 17.676 52.852 18.036 57.308 ; 
        RECT 15.084 52.708 15.156 57.344 ; 
        RECT 0.468 52.706 0.54 57.346 ; 
        RECT 37.908 57.026 37.98 61.666 ; 
        RECT 23.292 57.028 23.364 61.664 ; 
        RECT 17.676 57.172 18.036 61.628 ; 
        RECT 15.084 57.028 15.156 61.664 ; 
        RECT 0.468 57.026 0.54 61.666 ; 
        RECT 37.908 61.346 37.98 65.986 ; 
        RECT 23.292 61.348 23.364 65.984 ; 
        RECT 17.676 61.492 18.036 65.948 ; 
        RECT 15.084 61.348 15.156 65.984 ; 
        RECT 0.468 61.346 0.54 65.986 ; 
        RECT 37.908 65.666 37.98 70.306 ; 
        RECT 23.292 65.668 23.364 70.304 ; 
        RECT 17.676 65.812 18.036 70.268 ; 
        RECT 15.084 65.668 15.156 70.304 ; 
        RECT 0.468 65.666 0.54 70.306 ; 
        RECT 37.908 69.986 37.98 74.626 ; 
        RECT 23.292 69.988 23.364 74.624 ; 
        RECT 17.676 70.132 18.036 74.588 ; 
        RECT 15.084 69.988 15.156 74.624 ; 
        RECT 0.468 69.986 0.54 74.626 ; 
        RECT 37.908 74.306 37.98 78.946 ; 
        RECT 23.292 74.308 23.364 78.944 ; 
        RECT 17.676 74.452 18.036 78.908 ; 
        RECT 15.084 74.308 15.156 78.944 ; 
        RECT 0.468 74.306 0.54 78.946 ; 
        RECT 37.908 78.626 37.98 83.266 ; 
        RECT 23.292 78.628 23.364 83.264 ; 
        RECT 17.676 78.772 18.036 83.228 ; 
        RECT 15.084 78.628 15.156 83.264 ; 
        RECT 0.468 78.626 0.54 83.266 ; 
        RECT 37.908 82.946 37.98 87.586 ; 
        RECT 23.292 82.948 23.364 87.584 ; 
        RECT 17.676 83.092 18.036 87.548 ; 
        RECT 15.084 82.948 15.156 87.584 ; 
        RECT 0.468 82.946 0.54 87.586 ; 
        RECT 37.908 87.266 37.98 91.906 ; 
        RECT 23.292 87.268 23.364 91.904 ; 
        RECT 17.676 87.412 18.036 91.868 ; 
        RECT 15.084 87.268 15.156 91.904 ; 
        RECT 0.468 87.266 0.54 91.906 ; 
        RECT 37.908 91.586 37.98 96.226 ; 
        RECT 23.292 91.588 23.364 96.224 ; 
        RECT 17.676 91.732 18.036 96.188 ; 
        RECT 15.084 91.588 15.156 96.224 ; 
        RECT 0.468 91.586 0.54 96.226 ; 
        RECT 37.908 95.906 37.98 100.546 ; 
        RECT 23.292 95.908 23.364 100.544 ; 
        RECT 17.676 96.052 18.036 100.508 ; 
        RECT 15.084 95.908 15.156 100.544 ; 
        RECT 0.468 95.906 0.54 100.546 ; 
        RECT 37.908 100.226 37.98 104.866 ; 
        RECT 23.292 100.228 23.364 104.864 ; 
        RECT 17.676 100.372 18.036 104.828 ; 
        RECT 15.084 100.228 15.156 104.864 ; 
        RECT 0.468 100.226 0.54 104.866 ; 
        RECT 37.908 104.546 37.98 137.374 ; 
        RECT 23.292 104.864 23.364 105.23 ; 
        RECT 23.292 119.824 23.364 137.264 ; 
        RECT 17.82 105.84 18.756 136.172 ; 
        RECT 17.676 135.828 18.036 137.968 ; 
        RECT 17.676 104.72 18.036 106.86 ; 
        RECT 0.468 104.546 0.54 137.374 ; 
        RECT 37.908 137.054 37.98 141.694 ; 
        RECT 23.292 137.056 23.364 141.692 ; 
        RECT 17.676 137.2 18.036 141.656 ; 
        RECT 15.084 137.056 15.156 141.692 ; 
        RECT 0.468 137.054 0.54 141.694 ; 
        RECT 37.908 141.374 37.98 146.014 ; 
        RECT 23.292 141.376 23.364 146.012 ; 
        RECT 17.676 141.52 18.036 145.976 ; 
        RECT 15.084 141.376 15.156 146.012 ; 
        RECT 0.468 141.374 0.54 146.014 ; 
        RECT 37.908 145.694 37.98 150.334 ; 
        RECT 23.292 145.696 23.364 150.332 ; 
        RECT 17.676 145.84 18.036 150.296 ; 
        RECT 15.084 145.696 15.156 150.332 ; 
        RECT 0.468 145.694 0.54 150.334 ; 
        RECT 37.908 150.014 37.98 154.654 ; 
        RECT 23.292 150.016 23.364 154.652 ; 
        RECT 17.676 150.16 18.036 154.616 ; 
        RECT 15.084 150.016 15.156 154.652 ; 
        RECT 0.468 150.014 0.54 154.654 ; 
        RECT 37.908 154.334 37.98 158.974 ; 
        RECT 23.292 154.336 23.364 158.972 ; 
        RECT 17.676 154.48 18.036 158.936 ; 
        RECT 15.084 154.336 15.156 158.972 ; 
        RECT 0.468 154.334 0.54 158.974 ; 
        RECT 37.908 158.654 37.98 163.294 ; 
        RECT 23.292 158.656 23.364 163.292 ; 
        RECT 17.676 158.8 18.036 163.256 ; 
        RECT 15.084 158.656 15.156 163.292 ; 
        RECT 0.468 158.654 0.54 163.294 ; 
        RECT 37.908 162.974 37.98 167.614 ; 
        RECT 23.292 162.976 23.364 167.612 ; 
        RECT 17.676 163.12 18.036 167.576 ; 
        RECT 15.084 162.976 15.156 167.612 ; 
        RECT 0.468 162.974 0.54 167.614 ; 
        RECT 37.908 167.294 37.98 171.934 ; 
        RECT 23.292 167.296 23.364 171.932 ; 
        RECT 17.676 167.44 18.036 171.896 ; 
        RECT 15.084 167.296 15.156 171.932 ; 
        RECT 0.468 167.294 0.54 171.934 ; 
        RECT 37.908 171.614 37.98 176.254 ; 
        RECT 23.292 171.616 23.364 176.252 ; 
        RECT 17.676 171.76 18.036 176.216 ; 
        RECT 15.084 171.616 15.156 176.252 ; 
        RECT 0.468 171.614 0.54 176.254 ; 
        RECT 37.908 175.934 37.98 180.574 ; 
        RECT 23.292 175.936 23.364 180.572 ; 
        RECT 17.676 176.08 18.036 180.536 ; 
        RECT 15.084 175.936 15.156 180.572 ; 
        RECT 0.468 175.934 0.54 180.574 ; 
        RECT 37.908 180.254 37.98 184.894 ; 
        RECT 23.292 180.256 23.364 184.892 ; 
        RECT 17.676 180.4 18.036 184.856 ; 
        RECT 15.084 180.256 15.156 184.892 ; 
        RECT 0.468 180.254 0.54 184.894 ; 
        RECT 37.908 184.574 37.98 189.214 ; 
        RECT 23.292 184.576 23.364 189.212 ; 
        RECT 17.676 184.72 18.036 189.176 ; 
        RECT 15.084 184.576 15.156 189.212 ; 
        RECT 0.468 184.574 0.54 189.214 ; 
        RECT 37.908 188.894 37.98 193.534 ; 
        RECT 23.292 188.896 23.364 193.532 ; 
        RECT 17.676 189.04 18.036 193.496 ; 
        RECT 15.084 188.896 15.156 193.532 ; 
        RECT 0.468 188.894 0.54 193.534 ; 
        RECT 37.908 193.214 37.98 197.854 ; 
        RECT 23.292 193.216 23.364 197.852 ; 
        RECT 17.676 193.36 18.036 197.816 ; 
        RECT 15.084 193.216 15.156 197.852 ; 
        RECT 0.468 193.214 0.54 197.854 ; 
        RECT 37.908 197.534 37.98 202.174 ; 
        RECT 23.292 197.536 23.364 202.172 ; 
        RECT 17.676 197.68 18.036 202.136 ; 
        RECT 15.084 197.536 15.156 202.172 ; 
        RECT 0.468 197.534 0.54 202.174 ; 
        RECT 37.908 201.854 37.98 206.494 ; 
        RECT 23.292 201.856 23.364 206.492 ; 
        RECT 17.676 202 18.036 206.456 ; 
        RECT 15.084 201.856 15.156 206.492 ; 
        RECT 0.468 201.854 0.54 206.494 ; 
        RECT 37.908 206.174 37.98 210.814 ; 
        RECT 23.292 206.176 23.364 210.812 ; 
        RECT 17.676 206.32 18.036 210.776 ; 
        RECT 15.084 206.176 15.156 210.812 ; 
        RECT 0.468 206.174 0.54 210.814 ; 
        RECT 37.908 210.494 37.98 215.134 ; 
        RECT 23.292 210.496 23.364 215.132 ; 
        RECT 17.676 210.64 18.036 215.096 ; 
        RECT 15.084 210.496 15.156 215.132 ; 
        RECT 0.468 210.494 0.54 215.134 ; 
        RECT 37.908 214.814 37.98 219.454 ; 
        RECT 23.292 214.816 23.364 219.452 ; 
        RECT 17.676 214.96 18.036 219.416 ; 
        RECT 15.084 214.816 15.156 219.452 ; 
        RECT 0.468 214.814 0.54 219.454 ; 
        RECT 37.908 219.134 37.98 223.774 ; 
        RECT 23.292 219.136 23.364 223.772 ; 
        RECT 17.676 219.28 18.036 223.736 ; 
        RECT 15.084 219.136 15.156 223.772 ; 
        RECT 0.468 219.134 0.54 223.774 ; 
        RECT 37.908 223.454 37.98 228.094 ; 
        RECT 23.292 223.456 23.364 228.092 ; 
        RECT 17.676 223.6 18.036 228.056 ; 
        RECT 15.084 223.456 15.156 228.092 ; 
        RECT 0.468 223.454 0.54 228.094 ; 
        RECT 37.908 227.774 37.98 232.414 ; 
        RECT 23.292 227.776 23.364 232.412 ; 
        RECT 17.676 227.92 18.036 232.376 ; 
        RECT 15.084 227.776 15.156 232.412 ; 
        RECT 0.468 227.774 0.54 232.414 ; 
        RECT 37.908 232.094 37.98 236.734 ; 
        RECT 23.292 232.096 23.364 236.732 ; 
        RECT 17.676 232.24 18.036 236.696 ; 
        RECT 15.084 232.096 15.156 236.732 ; 
        RECT 0.468 232.094 0.54 236.734 ; 
        RECT 37.908 236.414 37.98 241.054 ; 
        RECT 23.292 236.416 23.364 241.052 ; 
        RECT 17.676 236.56 18.036 241.016 ; 
        RECT 15.084 236.416 15.156 241.052 ; 
        RECT 0.468 236.414 0.54 241.054 ; 
      LAYER V3 ; 
        RECT 0.468 4.688 0.54 4.88 ; 
        RECT 15.084 4.688 15.156 4.88 ; 
        RECT 17.676 4.688 18.036 4.88 ; 
        RECT 23.292 4.688 23.364 4.88 ; 
        RECT 37.908 4.688 37.98 4.88 ; 
        RECT 0.468 9.008 0.54 9.2 ; 
        RECT 15.084 9.008 15.156 9.2 ; 
        RECT 17.676 9.008 18.036 9.2 ; 
        RECT 23.292 9.008 23.364 9.2 ; 
        RECT 37.908 9.008 37.98 9.2 ; 
        RECT 0.468 13.328 0.54 13.52 ; 
        RECT 15.084 13.328 15.156 13.52 ; 
        RECT 17.676 13.328 18.036 13.52 ; 
        RECT 23.292 13.328 23.364 13.52 ; 
        RECT 37.908 13.328 37.98 13.52 ; 
        RECT 0.468 17.648 0.54 17.84 ; 
        RECT 15.084 17.648 15.156 17.84 ; 
        RECT 17.676 17.648 18.036 17.84 ; 
        RECT 23.292 17.648 23.364 17.84 ; 
        RECT 37.908 17.648 37.98 17.84 ; 
        RECT 0.468 21.968 0.54 22.16 ; 
        RECT 15.084 21.968 15.156 22.16 ; 
        RECT 17.676 21.968 18.036 22.16 ; 
        RECT 23.292 21.968 23.364 22.16 ; 
        RECT 37.908 21.968 37.98 22.16 ; 
        RECT 0.468 26.288 0.54 26.48 ; 
        RECT 15.084 26.288 15.156 26.48 ; 
        RECT 17.676 26.288 18.036 26.48 ; 
        RECT 23.292 26.288 23.364 26.48 ; 
        RECT 37.908 26.288 37.98 26.48 ; 
        RECT 0.468 30.608 0.54 30.8 ; 
        RECT 15.084 30.608 15.156 30.8 ; 
        RECT 17.676 30.608 18.036 30.8 ; 
        RECT 23.292 30.608 23.364 30.8 ; 
        RECT 37.908 30.608 37.98 30.8 ; 
        RECT 0.468 34.928 0.54 35.12 ; 
        RECT 15.084 34.928 15.156 35.12 ; 
        RECT 17.676 34.928 18.036 35.12 ; 
        RECT 23.292 34.928 23.364 35.12 ; 
        RECT 37.908 34.928 37.98 35.12 ; 
        RECT 0.468 39.248 0.54 39.44 ; 
        RECT 15.084 39.248 15.156 39.44 ; 
        RECT 17.676 39.248 18.036 39.44 ; 
        RECT 23.292 39.248 23.364 39.44 ; 
        RECT 37.908 39.248 37.98 39.44 ; 
        RECT 0.468 43.568 0.54 43.76 ; 
        RECT 15.084 43.568 15.156 43.76 ; 
        RECT 17.676 43.568 18.036 43.76 ; 
        RECT 23.292 43.568 23.364 43.76 ; 
        RECT 37.908 43.568 37.98 43.76 ; 
        RECT 0.468 47.888 0.54 48.08 ; 
        RECT 15.084 47.888 15.156 48.08 ; 
        RECT 17.676 47.888 18.036 48.08 ; 
        RECT 23.292 47.888 23.364 48.08 ; 
        RECT 37.908 47.888 37.98 48.08 ; 
        RECT 0.468 52.208 0.54 52.4 ; 
        RECT 15.084 52.208 15.156 52.4 ; 
        RECT 17.676 52.208 18.036 52.4 ; 
        RECT 23.292 52.208 23.364 52.4 ; 
        RECT 37.908 52.208 37.98 52.4 ; 
        RECT 0.468 56.528 0.54 56.72 ; 
        RECT 15.084 56.528 15.156 56.72 ; 
        RECT 17.676 56.528 18.036 56.72 ; 
        RECT 23.292 56.528 23.364 56.72 ; 
        RECT 37.908 56.528 37.98 56.72 ; 
        RECT 0.468 60.848 0.54 61.04 ; 
        RECT 15.084 60.848 15.156 61.04 ; 
        RECT 17.676 60.848 18.036 61.04 ; 
        RECT 23.292 60.848 23.364 61.04 ; 
        RECT 37.908 60.848 37.98 61.04 ; 
        RECT 0.468 65.168 0.54 65.36 ; 
        RECT 15.084 65.168 15.156 65.36 ; 
        RECT 17.676 65.168 18.036 65.36 ; 
        RECT 23.292 65.168 23.364 65.36 ; 
        RECT 37.908 65.168 37.98 65.36 ; 
        RECT 0.468 69.488 0.54 69.68 ; 
        RECT 15.084 69.488 15.156 69.68 ; 
        RECT 17.676 69.488 18.036 69.68 ; 
        RECT 23.292 69.488 23.364 69.68 ; 
        RECT 37.908 69.488 37.98 69.68 ; 
        RECT 0.468 73.808 0.54 74 ; 
        RECT 15.084 73.808 15.156 74 ; 
        RECT 17.676 73.808 18.036 74 ; 
        RECT 23.292 73.808 23.364 74 ; 
        RECT 37.908 73.808 37.98 74 ; 
        RECT 0.468 78.128 0.54 78.32 ; 
        RECT 15.084 78.128 15.156 78.32 ; 
        RECT 17.676 78.128 18.036 78.32 ; 
        RECT 23.292 78.128 23.364 78.32 ; 
        RECT 37.908 78.128 37.98 78.32 ; 
        RECT 0.468 82.448 0.54 82.64 ; 
        RECT 15.084 82.448 15.156 82.64 ; 
        RECT 17.676 82.448 18.036 82.64 ; 
        RECT 23.292 82.448 23.364 82.64 ; 
        RECT 37.908 82.448 37.98 82.64 ; 
        RECT 0.468 86.768 0.54 86.96 ; 
        RECT 15.084 86.768 15.156 86.96 ; 
        RECT 17.676 86.768 18.036 86.96 ; 
        RECT 23.292 86.768 23.364 86.96 ; 
        RECT 37.908 86.768 37.98 86.96 ; 
        RECT 0.468 91.088 0.54 91.28 ; 
        RECT 15.084 91.088 15.156 91.28 ; 
        RECT 17.676 91.088 18.036 91.28 ; 
        RECT 23.292 91.088 23.364 91.28 ; 
        RECT 37.908 91.088 37.98 91.28 ; 
        RECT 0.468 95.408 0.54 95.6 ; 
        RECT 15.084 95.408 15.156 95.6 ; 
        RECT 17.676 95.408 18.036 95.6 ; 
        RECT 23.292 95.408 23.364 95.6 ; 
        RECT 37.908 95.408 37.98 95.6 ; 
        RECT 0.468 99.728 0.54 99.92 ; 
        RECT 15.084 99.728 15.156 99.92 ; 
        RECT 17.676 99.728 18.036 99.92 ; 
        RECT 23.292 99.728 23.364 99.92 ; 
        RECT 37.908 99.728 37.98 99.92 ; 
        RECT 0.468 104.048 0.54 104.24 ; 
        RECT 15.084 104.048 15.156 104.24 ; 
        RECT 17.676 104.048 18.036 104.24 ; 
        RECT 23.292 104.048 23.364 104.24 ; 
        RECT 37.908 104.048 37.98 104.24 ; 
        RECT 0.468 105.996 0.54 106.86 ; 
        RECT 17.836 131.34 17.908 132.204 ; 
        RECT 17.836 118.668 17.908 119.532 ; 
        RECT 17.836 105.996 17.908 106.86 ; 
        RECT 18.044 131.34 18.116 132.204 ; 
        RECT 18.044 118.668 18.116 119.532 ; 
        RECT 18.044 105.996 18.116 106.86 ; 
        RECT 18.252 131.34 18.324 132.204 ; 
        RECT 18.252 118.668 18.324 119.532 ; 
        RECT 18.252 105.996 18.324 106.86 ; 
        RECT 18.46 131.34 18.532 132.204 ; 
        RECT 18.46 118.668 18.532 119.532 ; 
        RECT 18.46 105.996 18.532 106.86 ; 
        RECT 18.668 131.34 18.74 132.204 ; 
        RECT 18.668 118.668 18.74 119.532 ; 
        RECT 18.668 105.996 18.74 106.86 ; 
        RECT 23.292 120.012 23.364 120.108 ; 
        RECT 23.292 104.876 23.364 104.972 ; 
        RECT 0.468 140.876 0.54 141.068 ; 
        RECT 15.084 140.876 15.156 141.068 ; 
        RECT 17.676 140.876 18.036 141.068 ; 
        RECT 23.292 140.876 23.364 141.068 ; 
        RECT 37.908 140.876 37.98 141.068 ; 
        RECT 0.468 145.196 0.54 145.388 ; 
        RECT 15.084 145.196 15.156 145.388 ; 
        RECT 17.676 145.196 18.036 145.388 ; 
        RECT 23.292 145.196 23.364 145.388 ; 
        RECT 37.908 145.196 37.98 145.388 ; 
        RECT 0.468 149.516 0.54 149.708 ; 
        RECT 15.084 149.516 15.156 149.708 ; 
        RECT 17.676 149.516 18.036 149.708 ; 
        RECT 23.292 149.516 23.364 149.708 ; 
        RECT 37.908 149.516 37.98 149.708 ; 
        RECT 0.468 153.836 0.54 154.028 ; 
        RECT 15.084 153.836 15.156 154.028 ; 
        RECT 17.676 153.836 18.036 154.028 ; 
        RECT 23.292 153.836 23.364 154.028 ; 
        RECT 37.908 153.836 37.98 154.028 ; 
        RECT 0.468 158.156 0.54 158.348 ; 
        RECT 15.084 158.156 15.156 158.348 ; 
        RECT 17.676 158.156 18.036 158.348 ; 
        RECT 23.292 158.156 23.364 158.348 ; 
        RECT 37.908 158.156 37.98 158.348 ; 
        RECT 0.468 162.476 0.54 162.668 ; 
        RECT 15.084 162.476 15.156 162.668 ; 
        RECT 17.676 162.476 18.036 162.668 ; 
        RECT 23.292 162.476 23.364 162.668 ; 
        RECT 37.908 162.476 37.98 162.668 ; 
        RECT 0.468 166.796 0.54 166.988 ; 
        RECT 15.084 166.796 15.156 166.988 ; 
        RECT 17.676 166.796 18.036 166.988 ; 
        RECT 23.292 166.796 23.364 166.988 ; 
        RECT 37.908 166.796 37.98 166.988 ; 
        RECT 0.468 171.116 0.54 171.308 ; 
        RECT 15.084 171.116 15.156 171.308 ; 
        RECT 17.676 171.116 18.036 171.308 ; 
        RECT 23.292 171.116 23.364 171.308 ; 
        RECT 37.908 171.116 37.98 171.308 ; 
        RECT 0.468 175.436 0.54 175.628 ; 
        RECT 15.084 175.436 15.156 175.628 ; 
        RECT 17.676 175.436 18.036 175.628 ; 
        RECT 23.292 175.436 23.364 175.628 ; 
        RECT 37.908 175.436 37.98 175.628 ; 
        RECT 0.468 179.756 0.54 179.948 ; 
        RECT 15.084 179.756 15.156 179.948 ; 
        RECT 17.676 179.756 18.036 179.948 ; 
        RECT 23.292 179.756 23.364 179.948 ; 
        RECT 37.908 179.756 37.98 179.948 ; 
        RECT 0.468 184.076 0.54 184.268 ; 
        RECT 15.084 184.076 15.156 184.268 ; 
        RECT 17.676 184.076 18.036 184.268 ; 
        RECT 23.292 184.076 23.364 184.268 ; 
        RECT 37.908 184.076 37.98 184.268 ; 
        RECT 0.468 188.396 0.54 188.588 ; 
        RECT 15.084 188.396 15.156 188.588 ; 
        RECT 17.676 188.396 18.036 188.588 ; 
        RECT 23.292 188.396 23.364 188.588 ; 
        RECT 37.908 188.396 37.98 188.588 ; 
        RECT 0.468 192.716 0.54 192.908 ; 
        RECT 15.084 192.716 15.156 192.908 ; 
        RECT 17.676 192.716 18.036 192.908 ; 
        RECT 23.292 192.716 23.364 192.908 ; 
        RECT 37.908 192.716 37.98 192.908 ; 
        RECT 0.468 197.036 0.54 197.228 ; 
        RECT 15.084 197.036 15.156 197.228 ; 
        RECT 17.676 197.036 18.036 197.228 ; 
        RECT 23.292 197.036 23.364 197.228 ; 
        RECT 37.908 197.036 37.98 197.228 ; 
        RECT 0.468 201.356 0.54 201.548 ; 
        RECT 15.084 201.356 15.156 201.548 ; 
        RECT 17.676 201.356 18.036 201.548 ; 
        RECT 23.292 201.356 23.364 201.548 ; 
        RECT 37.908 201.356 37.98 201.548 ; 
        RECT 0.468 205.676 0.54 205.868 ; 
        RECT 15.084 205.676 15.156 205.868 ; 
        RECT 17.676 205.676 18.036 205.868 ; 
        RECT 23.292 205.676 23.364 205.868 ; 
        RECT 37.908 205.676 37.98 205.868 ; 
        RECT 0.468 209.996 0.54 210.188 ; 
        RECT 15.084 209.996 15.156 210.188 ; 
        RECT 17.676 209.996 18.036 210.188 ; 
        RECT 23.292 209.996 23.364 210.188 ; 
        RECT 37.908 209.996 37.98 210.188 ; 
        RECT 0.468 214.316 0.54 214.508 ; 
        RECT 15.084 214.316 15.156 214.508 ; 
        RECT 17.676 214.316 18.036 214.508 ; 
        RECT 23.292 214.316 23.364 214.508 ; 
        RECT 37.908 214.316 37.98 214.508 ; 
        RECT 0.468 218.636 0.54 218.828 ; 
        RECT 15.084 218.636 15.156 218.828 ; 
        RECT 17.676 218.636 18.036 218.828 ; 
        RECT 23.292 218.636 23.364 218.828 ; 
        RECT 37.908 218.636 37.98 218.828 ; 
        RECT 0.468 222.956 0.54 223.148 ; 
        RECT 15.084 222.956 15.156 223.148 ; 
        RECT 17.676 222.956 18.036 223.148 ; 
        RECT 23.292 222.956 23.364 223.148 ; 
        RECT 37.908 222.956 37.98 223.148 ; 
        RECT 0.468 227.276 0.54 227.468 ; 
        RECT 15.084 227.276 15.156 227.468 ; 
        RECT 17.676 227.276 18.036 227.468 ; 
        RECT 23.292 227.276 23.364 227.468 ; 
        RECT 37.908 227.276 37.98 227.468 ; 
        RECT 0.468 231.596 0.54 231.788 ; 
        RECT 15.084 231.596 15.156 231.788 ; 
        RECT 17.676 231.596 18.036 231.788 ; 
        RECT 23.292 231.596 23.364 231.788 ; 
        RECT 37.908 231.596 37.98 231.788 ; 
        RECT 0.468 235.916 0.54 236.108 ; 
        RECT 15.084 235.916 15.156 236.108 ; 
        RECT 17.676 235.916 18.036 236.108 ; 
        RECT 23.292 235.916 23.364 236.108 ; 
        RECT 37.908 235.916 37.98 236.108 ; 
        RECT 0.468 240.236 0.54 240.428 ; 
        RECT 15.084 240.236 15.156 240.428 ; 
        RECT 17.676 240.236 18.036 240.428 ; 
        RECT 23.292 240.236 23.364 240.428 ; 
        RECT 37.908 240.236 37.98 240.428 ; 
      LAYER M5 ; 
        RECT 23.036 104.804 23.132 120.18 ; 
      LAYER V4 ; 
        RECT 23.036 120.012 23.132 120.108 ; 
        RECT 23.036 104.876 23.132 104.972 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.304 38.016 4.496 ; 
        RECT 0.404 8.624 38.016 8.816 ; 
        RECT 0.404 12.944 38.016 13.136 ; 
        RECT 0.404 17.264 38.016 17.456 ; 
        RECT 0.404 21.584 38.016 21.776 ; 
        RECT 0.404 25.904 38.016 26.096 ; 
        RECT 0.404 30.224 38.016 30.416 ; 
        RECT 0.404 34.544 38.016 34.736 ; 
        RECT 0.404 38.864 38.016 39.056 ; 
        RECT 0.404 43.184 38.016 43.376 ; 
        RECT 0.404 47.504 38.016 47.696 ; 
        RECT 0.404 51.824 38.016 52.016 ; 
        RECT 0.404 56.144 38.016 56.336 ; 
        RECT 0.404 60.464 38.016 60.656 ; 
        RECT 0.404 64.784 38.016 64.976 ; 
        RECT 0.404 69.104 38.016 69.296 ; 
        RECT 0.404 73.424 38.016 73.616 ; 
        RECT 0.404 77.744 38.016 77.936 ; 
        RECT 0.404 82.064 38.016 82.256 ; 
        RECT 0.404 86.384 38.016 86.576 ; 
        RECT 0.404 90.704 38.016 90.896 ; 
        RECT 0.404 95.024 38.016 95.216 ; 
        RECT 0.404 99.344 38.016 99.536 ; 
        RECT 0.404 103.664 38.016 103.856 ; 
        RECT 0.432 107.724 38.016 108.588 ; 
        RECT 15.768 120.396 22.68 121.26 ; 
        RECT 15.768 133.068 22.68 133.932 ; 
        RECT 0.404 140.492 38.016 140.684 ; 
        RECT 0.404 144.812 38.016 145.004 ; 
        RECT 0.404 149.132 38.016 149.324 ; 
        RECT 0.404 153.452 38.016 153.644 ; 
        RECT 0.404 157.772 38.016 157.964 ; 
        RECT 0.404 162.092 38.016 162.284 ; 
        RECT 0.404 166.412 38.016 166.604 ; 
        RECT 0.404 170.732 38.016 170.924 ; 
        RECT 0.404 175.052 38.016 175.244 ; 
        RECT 0.404 179.372 38.016 179.564 ; 
        RECT 0.404 183.692 38.016 183.884 ; 
        RECT 0.404 188.012 38.016 188.204 ; 
        RECT 0.404 192.332 38.016 192.524 ; 
        RECT 0.404 196.652 38.016 196.844 ; 
        RECT 0.404 200.972 38.016 201.164 ; 
        RECT 0.404 205.292 38.016 205.484 ; 
        RECT 0.404 209.612 38.016 209.804 ; 
        RECT 0.404 213.932 38.016 214.124 ; 
        RECT 0.404 218.252 38.016 218.444 ; 
        RECT 0.404 222.572 38.016 222.764 ; 
        RECT 0.404 226.892 38.016 227.084 ; 
        RECT 0.404 231.212 38.016 231.404 ; 
        RECT 0.404 235.532 38.016 235.724 ; 
        RECT 0.404 239.852 38.016 240.044 ; 
      LAYER M3 ; 
        RECT 37.764 0.866 37.836 5.506 ; 
        RECT 23.508 0.866 23.58 5.506 ; 
        RECT 20.448 1.012 20.592 5.468 ; 
        RECT 19.836 1.012 19.944 5.468 ; 
        RECT 14.868 0.866 14.94 5.506 ; 
        RECT 0.612 0.866 0.684 5.506 ; 
        RECT 37.764 5.186 37.836 9.826 ; 
        RECT 23.508 5.186 23.58 9.826 ; 
        RECT 20.448 5.332 20.592 9.788 ; 
        RECT 19.836 5.332 19.944 9.788 ; 
        RECT 14.868 5.186 14.94 9.826 ; 
        RECT 0.612 5.186 0.684 9.826 ; 
        RECT 37.764 9.506 37.836 14.146 ; 
        RECT 23.508 9.506 23.58 14.146 ; 
        RECT 20.448 9.652 20.592 14.108 ; 
        RECT 19.836 9.652 19.944 14.108 ; 
        RECT 14.868 9.506 14.94 14.146 ; 
        RECT 0.612 9.506 0.684 14.146 ; 
        RECT 37.764 13.826 37.836 18.466 ; 
        RECT 23.508 13.826 23.58 18.466 ; 
        RECT 20.448 13.972 20.592 18.428 ; 
        RECT 19.836 13.972 19.944 18.428 ; 
        RECT 14.868 13.826 14.94 18.466 ; 
        RECT 0.612 13.826 0.684 18.466 ; 
        RECT 37.764 18.146 37.836 22.786 ; 
        RECT 23.508 18.146 23.58 22.786 ; 
        RECT 20.448 18.292 20.592 22.748 ; 
        RECT 19.836 18.292 19.944 22.748 ; 
        RECT 14.868 18.146 14.94 22.786 ; 
        RECT 0.612 18.146 0.684 22.786 ; 
        RECT 37.764 22.466 37.836 27.106 ; 
        RECT 23.508 22.466 23.58 27.106 ; 
        RECT 20.448 22.612 20.592 27.068 ; 
        RECT 19.836 22.612 19.944 27.068 ; 
        RECT 14.868 22.466 14.94 27.106 ; 
        RECT 0.612 22.466 0.684 27.106 ; 
        RECT 37.764 26.786 37.836 31.426 ; 
        RECT 23.508 26.786 23.58 31.426 ; 
        RECT 20.448 26.932 20.592 31.388 ; 
        RECT 19.836 26.932 19.944 31.388 ; 
        RECT 14.868 26.786 14.94 31.426 ; 
        RECT 0.612 26.786 0.684 31.426 ; 
        RECT 37.764 31.106 37.836 35.746 ; 
        RECT 23.508 31.106 23.58 35.746 ; 
        RECT 20.448 31.252 20.592 35.708 ; 
        RECT 19.836 31.252 19.944 35.708 ; 
        RECT 14.868 31.106 14.94 35.746 ; 
        RECT 0.612 31.106 0.684 35.746 ; 
        RECT 37.764 35.426 37.836 40.066 ; 
        RECT 23.508 35.426 23.58 40.066 ; 
        RECT 20.448 35.572 20.592 40.028 ; 
        RECT 19.836 35.572 19.944 40.028 ; 
        RECT 14.868 35.426 14.94 40.066 ; 
        RECT 0.612 35.426 0.684 40.066 ; 
        RECT 37.764 39.746 37.836 44.386 ; 
        RECT 23.508 39.746 23.58 44.386 ; 
        RECT 20.448 39.892 20.592 44.348 ; 
        RECT 19.836 39.892 19.944 44.348 ; 
        RECT 14.868 39.746 14.94 44.386 ; 
        RECT 0.612 39.746 0.684 44.386 ; 
        RECT 37.764 44.066 37.836 48.706 ; 
        RECT 23.508 44.066 23.58 48.706 ; 
        RECT 20.448 44.212 20.592 48.668 ; 
        RECT 19.836 44.212 19.944 48.668 ; 
        RECT 14.868 44.066 14.94 48.706 ; 
        RECT 0.612 44.066 0.684 48.706 ; 
        RECT 37.764 48.386 37.836 53.026 ; 
        RECT 23.508 48.386 23.58 53.026 ; 
        RECT 20.448 48.532 20.592 52.988 ; 
        RECT 19.836 48.532 19.944 52.988 ; 
        RECT 14.868 48.386 14.94 53.026 ; 
        RECT 0.612 48.386 0.684 53.026 ; 
        RECT 37.764 52.706 37.836 57.346 ; 
        RECT 23.508 52.706 23.58 57.346 ; 
        RECT 20.448 52.852 20.592 57.308 ; 
        RECT 19.836 52.852 19.944 57.308 ; 
        RECT 14.868 52.706 14.94 57.346 ; 
        RECT 0.612 52.706 0.684 57.346 ; 
        RECT 37.764 57.026 37.836 61.666 ; 
        RECT 23.508 57.026 23.58 61.666 ; 
        RECT 20.448 57.172 20.592 61.628 ; 
        RECT 19.836 57.172 19.944 61.628 ; 
        RECT 14.868 57.026 14.94 61.666 ; 
        RECT 0.612 57.026 0.684 61.666 ; 
        RECT 37.764 61.346 37.836 65.986 ; 
        RECT 23.508 61.346 23.58 65.986 ; 
        RECT 20.448 61.492 20.592 65.948 ; 
        RECT 19.836 61.492 19.944 65.948 ; 
        RECT 14.868 61.346 14.94 65.986 ; 
        RECT 0.612 61.346 0.684 65.986 ; 
        RECT 37.764 65.666 37.836 70.306 ; 
        RECT 23.508 65.666 23.58 70.306 ; 
        RECT 20.448 65.812 20.592 70.268 ; 
        RECT 19.836 65.812 19.944 70.268 ; 
        RECT 14.868 65.666 14.94 70.306 ; 
        RECT 0.612 65.666 0.684 70.306 ; 
        RECT 37.764 69.986 37.836 74.626 ; 
        RECT 23.508 69.986 23.58 74.626 ; 
        RECT 20.448 70.132 20.592 74.588 ; 
        RECT 19.836 70.132 19.944 74.588 ; 
        RECT 14.868 69.986 14.94 74.626 ; 
        RECT 0.612 69.986 0.684 74.626 ; 
        RECT 37.764 74.306 37.836 78.946 ; 
        RECT 23.508 74.306 23.58 78.946 ; 
        RECT 20.448 74.452 20.592 78.908 ; 
        RECT 19.836 74.452 19.944 78.908 ; 
        RECT 14.868 74.306 14.94 78.946 ; 
        RECT 0.612 74.306 0.684 78.946 ; 
        RECT 37.764 78.626 37.836 83.266 ; 
        RECT 23.508 78.626 23.58 83.266 ; 
        RECT 20.448 78.772 20.592 83.228 ; 
        RECT 19.836 78.772 19.944 83.228 ; 
        RECT 14.868 78.626 14.94 83.266 ; 
        RECT 0.612 78.626 0.684 83.266 ; 
        RECT 37.764 82.946 37.836 87.586 ; 
        RECT 23.508 82.946 23.58 87.586 ; 
        RECT 20.448 83.092 20.592 87.548 ; 
        RECT 19.836 83.092 19.944 87.548 ; 
        RECT 14.868 82.946 14.94 87.586 ; 
        RECT 0.612 82.946 0.684 87.586 ; 
        RECT 37.764 87.266 37.836 91.906 ; 
        RECT 23.508 87.266 23.58 91.906 ; 
        RECT 20.448 87.412 20.592 91.868 ; 
        RECT 19.836 87.412 19.944 91.868 ; 
        RECT 14.868 87.266 14.94 91.906 ; 
        RECT 0.612 87.266 0.684 91.906 ; 
        RECT 37.764 91.586 37.836 96.226 ; 
        RECT 23.508 91.586 23.58 96.226 ; 
        RECT 20.448 91.732 20.592 96.188 ; 
        RECT 19.836 91.732 19.944 96.188 ; 
        RECT 14.868 91.586 14.94 96.226 ; 
        RECT 0.612 91.586 0.684 96.226 ; 
        RECT 37.764 95.906 37.836 100.546 ; 
        RECT 23.508 95.906 23.58 100.546 ; 
        RECT 20.448 96.052 20.592 100.508 ; 
        RECT 19.836 96.052 19.944 100.508 ; 
        RECT 14.868 95.906 14.94 100.546 ; 
        RECT 0.612 95.906 0.684 100.546 ; 
        RECT 37.764 100.226 37.836 104.866 ; 
        RECT 23.508 100.226 23.58 104.866 ; 
        RECT 20.448 100.372 20.592 104.828 ; 
        RECT 19.836 100.372 19.944 104.828 ; 
        RECT 14.868 100.226 14.94 104.866 ; 
        RECT 0.612 100.226 0.684 104.866 ; 
        RECT 37.764 104.546 37.836 137.374 ; 
        RECT 23.508 104.546 23.58 137.374 ; 
        RECT 19.692 105.44 20.628 136.172 ; 
        RECT 20.448 104.72 20.592 137.268 ; 
        RECT 19.836 104.72 19.944 137.256 ; 
        RECT 14.868 104.546 14.94 137.374 ; 
        RECT 0.612 104.546 0.684 137.374 ; 
        RECT 37.764 137.054 37.836 141.694 ; 
        RECT 23.508 137.054 23.58 141.694 ; 
        RECT 20.448 137.2 20.592 141.656 ; 
        RECT 19.836 137.2 19.944 141.656 ; 
        RECT 14.868 137.054 14.94 141.694 ; 
        RECT 0.612 137.054 0.684 141.694 ; 
        RECT 37.764 141.374 37.836 146.014 ; 
        RECT 23.508 141.374 23.58 146.014 ; 
        RECT 20.448 141.52 20.592 145.976 ; 
        RECT 19.836 141.52 19.944 145.976 ; 
        RECT 14.868 141.374 14.94 146.014 ; 
        RECT 0.612 141.374 0.684 146.014 ; 
        RECT 37.764 145.694 37.836 150.334 ; 
        RECT 23.508 145.694 23.58 150.334 ; 
        RECT 20.448 145.84 20.592 150.296 ; 
        RECT 19.836 145.84 19.944 150.296 ; 
        RECT 14.868 145.694 14.94 150.334 ; 
        RECT 0.612 145.694 0.684 150.334 ; 
        RECT 37.764 150.014 37.836 154.654 ; 
        RECT 23.508 150.014 23.58 154.654 ; 
        RECT 20.448 150.16 20.592 154.616 ; 
        RECT 19.836 150.16 19.944 154.616 ; 
        RECT 14.868 150.014 14.94 154.654 ; 
        RECT 0.612 150.014 0.684 154.654 ; 
        RECT 37.764 154.334 37.836 158.974 ; 
        RECT 23.508 154.334 23.58 158.974 ; 
        RECT 20.448 154.48 20.592 158.936 ; 
        RECT 19.836 154.48 19.944 158.936 ; 
        RECT 14.868 154.334 14.94 158.974 ; 
        RECT 0.612 154.334 0.684 158.974 ; 
        RECT 37.764 158.654 37.836 163.294 ; 
        RECT 23.508 158.654 23.58 163.294 ; 
        RECT 20.448 158.8 20.592 163.256 ; 
        RECT 19.836 158.8 19.944 163.256 ; 
        RECT 14.868 158.654 14.94 163.294 ; 
        RECT 0.612 158.654 0.684 163.294 ; 
        RECT 37.764 162.974 37.836 167.614 ; 
        RECT 23.508 162.974 23.58 167.614 ; 
        RECT 20.448 163.12 20.592 167.576 ; 
        RECT 19.836 163.12 19.944 167.576 ; 
        RECT 14.868 162.974 14.94 167.614 ; 
        RECT 0.612 162.974 0.684 167.614 ; 
        RECT 37.764 167.294 37.836 171.934 ; 
        RECT 23.508 167.294 23.58 171.934 ; 
        RECT 20.448 167.44 20.592 171.896 ; 
        RECT 19.836 167.44 19.944 171.896 ; 
        RECT 14.868 167.294 14.94 171.934 ; 
        RECT 0.612 167.294 0.684 171.934 ; 
        RECT 37.764 171.614 37.836 176.254 ; 
        RECT 23.508 171.614 23.58 176.254 ; 
        RECT 20.448 171.76 20.592 176.216 ; 
        RECT 19.836 171.76 19.944 176.216 ; 
        RECT 14.868 171.614 14.94 176.254 ; 
        RECT 0.612 171.614 0.684 176.254 ; 
        RECT 37.764 175.934 37.836 180.574 ; 
        RECT 23.508 175.934 23.58 180.574 ; 
        RECT 20.448 176.08 20.592 180.536 ; 
        RECT 19.836 176.08 19.944 180.536 ; 
        RECT 14.868 175.934 14.94 180.574 ; 
        RECT 0.612 175.934 0.684 180.574 ; 
        RECT 37.764 180.254 37.836 184.894 ; 
        RECT 23.508 180.254 23.58 184.894 ; 
        RECT 20.448 180.4 20.592 184.856 ; 
        RECT 19.836 180.4 19.944 184.856 ; 
        RECT 14.868 180.254 14.94 184.894 ; 
        RECT 0.612 180.254 0.684 184.894 ; 
        RECT 37.764 184.574 37.836 189.214 ; 
        RECT 23.508 184.574 23.58 189.214 ; 
        RECT 20.448 184.72 20.592 189.176 ; 
        RECT 19.836 184.72 19.944 189.176 ; 
        RECT 14.868 184.574 14.94 189.214 ; 
        RECT 0.612 184.574 0.684 189.214 ; 
        RECT 37.764 188.894 37.836 193.534 ; 
        RECT 23.508 188.894 23.58 193.534 ; 
        RECT 20.448 189.04 20.592 193.496 ; 
        RECT 19.836 189.04 19.944 193.496 ; 
        RECT 14.868 188.894 14.94 193.534 ; 
        RECT 0.612 188.894 0.684 193.534 ; 
        RECT 37.764 193.214 37.836 197.854 ; 
        RECT 23.508 193.214 23.58 197.854 ; 
        RECT 20.448 193.36 20.592 197.816 ; 
        RECT 19.836 193.36 19.944 197.816 ; 
        RECT 14.868 193.214 14.94 197.854 ; 
        RECT 0.612 193.214 0.684 197.854 ; 
        RECT 37.764 197.534 37.836 202.174 ; 
        RECT 23.508 197.534 23.58 202.174 ; 
        RECT 20.448 197.68 20.592 202.136 ; 
        RECT 19.836 197.68 19.944 202.136 ; 
        RECT 14.868 197.534 14.94 202.174 ; 
        RECT 0.612 197.534 0.684 202.174 ; 
        RECT 37.764 201.854 37.836 206.494 ; 
        RECT 23.508 201.854 23.58 206.494 ; 
        RECT 20.448 202 20.592 206.456 ; 
        RECT 19.836 202 19.944 206.456 ; 
        RECT 14.868 201.854 14.94 206.494 ; 
        RECT 0.612 201.854 0.684 206.494 ; 
        RECT 37.764 206.174 37.836 210.814 ; 
        RECT 23.508 206.174 23.58 210.814 ; 
        RECT 20.448 206.32 20.592 210.776 ; 
        RECT 19.836 206.32 19.944 210.776 ; 
        RECT 14.868 206.174 14.94 210.814 ; 
        RECT 0.612 206.174 0.684 210.814 ; 
        RECT 37.764 210.494 37.836 215.134 ; 
        RECT 23.508 210.494 23.58 215.134 ; 
        RECT 20.448 210.64 20.592 215.096 ; 
        RECT 19.836 210.64 19.944 215.096 ; 
        RECT 14.868 210.494 14.94 215.134 ; 
        RECT 0.612 210.494 0.684 215.134 ; 
        RECT 37.764 214.814 37.836 219.454 ; 
        RECT 23.508 214.814 23.58 219.454 ; 
        RECT 20.448 214.96 20.592 219.416 ; 
        RECT 19.836 214.96 19.944 219.416 ; 
        RECT 14.868 214.814 14.94 219.454 ; 
        RECT 0.612 214.814 0.684 219.454 ; 
        RECT 37.764 219.134 37.836 223.774 ; 
        RECT 23.508 219.134 23.58 223.774 ; 
        RECT 20.448 219.28 20.592 223.736 ; 
        RECT 19.836 219.28 19.944 223.736 ; 
        RECT 14.868 219.134 14.94 223.774 ; 
        RECT 0.612 219.134 0.684 223.774 ; 
        RECT 37.764 223.454 37.836 228.094 ; 
        RECT 23.508 223.454 23.58 228.094 ; 
        RECT 20.448 223.6 20.592 228.056 ; 
        RECT 19.836 223.6 19.944 228.056 ; 
        RECT 14.868 223.454 14.94 228.094 ; 
        RECT 0.612 223.454 0.684 228.094 ; 
        RECT 37.764 227.774 37.836 232.414 ; 
        RECT 23.508 227.774 23.58 232.414 ; 
        RECT 20.448 227.92 20.592 232.376 ; 
        RECT 19.836 227.92 19.944 232.376 ; 
        RECT 14.868 227.774 14.94 232.414 ; 
        RECT 0.612 227.774 0.684 232.414 ; 
        RECT 37.764 232.094 37.836 236.734 ; 
        RECT 23.508 232.094 23.58 236.734 ; 
        RECT 20.448 232.24 20.592 236.696 ; 
        RECT 19.836 232.24 19.944 236.696 ; 
        RECT 14.868 232.094 14.94 236.734 ; 
        RECT 0.612 232.094 0.684 236.734 ; 
        RECT 37.764 236.414 37.836 241.054 ; 
        RECT 23.508 236.414 23.58 241.054 ; 
        RECT 20.448 236.56 20.592 241.016 ; 
        RECT 19.836 236.56 19.944 241.016 ; 
        RECT 14.868 236.414 14.94 241.054 ; 
        RECT 0.612 236.414 0.684 241.054 ; 
      LAYER V3 ; 
        RECT 0.612 4.304 0.684 4.496 ; 
        RECT 14.868 4.304 14.94 4.496 ; 
        RECT 19.836 4.304 19.944 4.496 ; 
        RECT 20.448 4.304 20.592 4.496 ; 
        RECT 23.508 4.304 23.58 4.496 ; 
        RECT 37.764 4.304 37.836 4.496 ; 
        RECT 0.612 8.624 0.684 8.816 ; 
        RECT 14.868 8.624 14.94 8.816 ; 
        RECT 19.836 8.624 19.944 8.816 ; 
        RECT 20.448 8.624 20.592 8.816 ; 
        RECT 23.508 8.624 23.58 8.816 ; 
        RECT 37.764 8.624 37.836 8.816 ; 
        RECT 0.612 12.944 0.684 13.136 ; 
        RECT 14.868 12.944 14.94 13.136 ; 
        RECT 19.836 12.944 19.944 13.136 ; 
        RECT 20.448 12.944 20.592 13.136 ; 
        RECT 23.508 12.944 23.58 13.136 ; 
        RECT 37.764 12.944 37.836 13.136 ; 
        RECT 0.612 17.264 0.684 17.456 ; 
        RECT 14.868 17.264 14.94 17.456 ; 
        RECT 19.836 17.264 19.944 17.456 ; 
        RECT 20.448 17.264 20.592 17.456 ; 
        RECT 23.508 17.264 23.58 17.456 ; 
        RECT 37.764 17.264 37.836 17.456 ; 
        RECT 0.612 21.584 0.684 21.776 ; 
        RECT 14.868 21.584 14.94 21.776 ; 
        RECT 19.836 21.584 19.944 21.776 ; 
        RECT 20.448 21.584 20.592 21.776 ; 
        RECT 23.508 21.584 23.58 21.776 ; 
        RECT 37.764 21.584 37.836 21.776 ; 
        RECT 0.612 25.904 0.684 26.096 ; 
        RECT 14.868 25.904 14.94 26.096 ; 
        RECT 19.836 25.904 19.944 26.096 ; 
        RECT 20.448 25.904 20.592 26.096 ; 
        RECT 23.508 25.904 23.58 26.096 ; 
        RECT 37.764 25.904 37.836 26.096 ; 
        RECT 0.612 30.224 0.684 30.416 ; 
        RECT 14.868 30.224 14.94 30.416 ; 
        RECT 19.836 30.224 19.944 30.416 ; 
        RECT 20.448 30.224 20.592 30.416 ; 
        RECT 23.508 30.224 23.58 30.416 ; 
        RECT 37.764 30.224 37.836 30.416 ; 
        RECT 0.612 34.544 0.684 34.736 ; 
        RECT 14.868 34.544 14.94 34.736 ; 
        RECT 19.836 34.544 19.944 34.736 ; 
        RECT 20.448 34.544 20.592 34.736 ; 
        RECT 23.508 34.544 23.58 34.736 ; 
        RECT 37.764 34.544 37.836 34.736 ; 
        RECT 0.612 38.864 0.684 39.056 ; 
        RECT 14.868 38.864 14.94 39.056 ; 
        RECT 19.836 38.864 19.944 39.056 ; 
        RECT 20.448 38.864 20.592 39.056 ; 
        RECT 23.508 38.864 23.58 39.056 ; 
        RECT 37.764 38.864 37.836 39.056 ; 
        RECT 0.612 43.184 0.684 43.376 ; 
        RECT 14.868 43.184 14.94 43.376 ; 
        RECT 19.836 43.184 19.944 43.376 ; 
        RECT 20.448 43.184 20.592 43.376 ; 
        RECT 23.508 43.184 23.58 43.376 ; 
        RECT 37.764 43.184 37.836 43.376 ; 
        RECT 0.612 47.504 0.684 47.696 ; 
        RECT 14.868 47.504 14.94 47.696 ; 
        RECT 19.836 47.504 19.944 47.696 ; 
        RECT 20.448 47.504 20.592 47.696 ; 
        RECT 23.508 47.504 23.58 47.696 ; 
        RECT 37.764 47.504 37.836 47.696 ; 
        RECT 0.612 51.824 0.684 52.016 ; 
        RECT 14.868 51.824 14.94 52.016 ; 
        RECT 19.836 51.824 19.944 52.016 ; 
        RECT 20.448 51.824 20.592 52.016 ; 
        RECT 23.508 51.824 23.58 52.016 ; 
        RECT 37.764 51.824 37.836 52.016 ; 
        RECT 0.612 56.144 0.684 56.336 ; 
        RECT 14.868 56.144 14.94 56.336 ; 
        RECT 19.836 56.144 19.944 56.336 ; 
        RECT 20.448 56.144 20.592 56.336 ; 
        RECT 23.508 56.144 23.58 56.336 ; 
        RECT 37.764 56.144 37.836 56.336 ; 
        RECT 0.612 60.464 0.684 60.656 ; 
        RECT 14.868 60.464 14.94 60.656 ; 
        RECT 19.836 60.464 19.944 60.656 ; 
        RECT 20.448 60.464 20.592 60.656 ; 
        RECT 23.508 60.464 23.58 60.656 ; 
        RECT 37.764 60.464 37.836 60.656 ; 
        RECT 0.612 64.784 0.684 64.976 ; 
        RECT 14.868 64.784 14.94 64.976 ; 
        RECT 19.836 64.784 19.944 64.976 ; 
        RECT 20.448 64.784 20.592 64.976 ; 
        RECT 23.508 64.784 23.58 64.976 ; 
        RECT 37.764 64.784 37.836 64.976 ; 
        RECT 0.612 69.104 0.684 69.296 ; 
        RECT 14.868 69.104 14.94 69.296 ; 
        RECT 19.836 69.104 19.944 69.296 ; 
        RECT 20.448 69.104 20.592 69.296 ; 
        RECT 23.508 69.104 23.58 69.296 ; 
        RECT 37.764 69.104 37.836 69.296 ; 
        RECT 0.612 73.424 0.684 73.616 ; 
        RECT 14.868 73.424 14.94 73.616 ; 
        RECT 19.836 73.424 19.944 73.616 ; 
        RECT 20.448 73.424 20.592 73.616 ; 
        RECT 23.508 73.424 23.58 73.616 ; 
        RECT 37.764 73.424 37.836 73.616 ; 
        RECT 0.612 77.744 0.684 77.936 ; 
        RECT 14.868 77.744 14.94 77.936 ; 
        RECT 19.836 77.744 19.944 77.936 ; 
        RECT 20.448 77.744 20.592 77.936 ; 
        RECT 23.508 77.744 23.58 77.936 ; 
        RECT 37.764 77.744 37.836 77.936 ; 
        RECT 0.612 82.064 0.684 82.256 ; 
        RECT 14.868 82.064 14.94 82.256 ; 
        RECT 19.836 82.064 19.944 82.256 ; 
        RECT 20.448 82.064 20.592 82.256 ; 
        RECT 23.508 82.064 23.58 82.256 ; 
        RECT 37.764 82.064 37.836 82.256 ; 
        RECT 0.612 86.384 0.684 86.576 ; 
        RECT 14.868 86.384 14.94 86.576 ; 
        RECT 19.836 86.384 19.944 86.576 ; 
        RECT 20.448 86.384 20.592 86.576 ; 
        RECT 23.508 86.384 23.58 86.576 ; 
        RECT 37.764 86.384 37.836 86.576 ; 
        RECT 0.612 90.704 0.684 90.896 ; 
        RECT 14.868 90.704 14.94 90.896 ; 
        RECT 19.836 90.704 19.944 90.896 ; 
        RECT 20.448 90.704 20.592 90.896 ; 
        RECT 23.508 90.704 23.58 90.896 ; 
        RECT 37.764 90.704 37.836 90.896 ; 
        RECT 0.612 95.024 0.684 95.216 ; 
        RECT 14.868 95.024 14.94 95.216 ; 
        RECT 19.836 95.024 19.944 95.216 ; 
        RECT 20.448 95.024 20.592 95.216 ; 
        RECT 23.508 95.024 23.58 95.216 ; 
        RECT 37.764 95.024 37.836 95.216 ; 
        RECT 0.612 99.344 0.684 99.536 ; 
        RECT 14.868 99.344 14.94 99.536 ; 
        RECT 19.836 99.344 19.944 99.536 ; 
        RECT 20.448 99.344 20.592 99.536 ; 
        RECT 23.508 99.344 23.58 99.536 ; 
        RECT 37.764 99.344 37.836 99.536 ; 
        RECT 0.612 103.664 0.684 103.856 ; 
        RECT 14.868 103.664 14.94 103.856 ; 
        RECT 19.836 103.664 19.944 103.856 ; 
        RECT 20.448 103.664 20.592 103.856 ; 
        RECT 23.508 103.664 23.58 103.856 ; 
        RECT 37.764 103.664 37.836 103.856 ; 
        RECT 0.612 107.724 0.684 108.588 ; 
        RECT 19.708 133.068 19.78 133.932 ; 
        RECT 19.708 120.396 19.78 121.26 ; 
        RECT 19.708 107.724 19.78 108.588 ; 
        RECT 19.916 133.068 19.988 133.932 ; 
        RECT 19.916 120.396 19.988 121.26 ; 
        RECT 19.916 107.724 19.988 108.588 ; 
        RECT 20.124 133.068 20.196 133.932 ; 
        RECT 20.124 120.396 20.196 121.26 ; 
        RECT 20.124 107.724 20.196 108.588 ; 
        RECT 20.332 133.068 20.404 133.932 ; 
        RECT 20.332 120.396 20.404 121.26 ; 
        RECT 20.332 107.724 20.404 108.588 ; 
        RECT 20.54 133.068 20.612 133.932 ; 
        RECT 20.54 120.396 20.612 121.26 ; 
        RECT 20.54 107.724 20.612 108.588 ; 
        RECT 0.612 140.492 0.684 140.684 ; 
        RECT 14.868 140.492 14.94 140.684 ; 
        RECT 19.836 140.492 19.944 140.684 ; 
        RECT 20.448 140.492 20.592 140.684 ; 
        RECT 23.508 140.492 23.58 140.684 ; 
        RECT 37.764 140.492 37.836 140.684 ; 
        RECT 0.612 144.812 0.684 145.004 ; 
        RECT 14.868 144.812 14.94 145.004 ; 
        RECT 19.836 144.812 19.944 145.004 ; 
        RECT 20.448 144.812 20.592 145.004 ; 
        RECT 23.508 144.812 23.58 145.004 ; 
        RECT 37.764 144.812 37.836 145.004 ; 
        RECT 0.612 149.132 0.684 149.324 ; 
        RECT 14.868 149.132 14.94 149.324 ; 
        RECT 19.836 149.132 19.944 149.324 ; 
        RECT 20.448 149.132 20.592 149.324 ; 
        RECT 23.508 149.132 23.58 149.324 ; 
        RECT 37.764 149.132 37.836 149.324 ; 
        RECT 0.612 153.452 0.684 153.644 ; 
        RECT 14.868 153.452 14.94 153.644 ; 
        RECT 19.836 153.452 19.944 153.644 ; 
        RECT 20.448 153.452 20.592 153.644 ; 
        RECT 23.508 153.452 23.58 153.644 ; 
        RECT 37.764 153.452 37.836 153.644 ; 
        RECT 0.612 157.772 0.684 157.964 ; 
        RECT 14.868 157.772 14.94 157.964 ; 
        RECT 19.836 157.772 19.944 157.964 ; 
        RECT 20.448 157.772 20.592 157.964 ; 
        RECT 23.508 157.772 23.58 157.964 ; 
        RECT 37.764 157.772 37.836 157.964 ; 
        RECT 0.612 162.092 0.684 162.284 ; 
        RECT 14.868 162.092 14.94 162.284 ; 
        RECT 19.836 162.092 19.944 162.284 ; 
        RECT 20.448 162.092 20.592 162.284 ; 
        RECT 23.508 162.092 23.58 162.284 ; 
        RECT 37.764 162.092 37.836 162.284 ; 
        RECT 0.612 166.412 0.684 166.604 ; 
        RECT 14.868 166.412 14.94 166.604 ; 
        RECT 19.836 166.412 19.944 166.604 ; 
        RECT 20.448 166.412 20.592 166.604 ; 
        RECT 23.508 166.412 23.58 166.604 ; 
        RECT 37.764 166.412 37.836 166.604 ; 
        RECT 0.612 170.732 0.684 170.924 ; 
        RECT 14.868 170.732 14.94 170.924 ; 
        RECT 19.836 170.732 19.944 170.924 ; 
        RECT 20.448 170.732 20.592 170.924 ; 
        RECT 23.508 170.732 23.58 170.924 ; 
        RECT 37.764 170.732 37.836 170.924 ; 
        RECT 0.612 175.052 0.684 175.244 ; 
        RECT 14.868 175.052 14.94 175.244 ; 
        RECT 19.836 175.052 19.944 175.244 ; 
        RECT 20.448 175.052 20.592 175.244 ; 
        RECT 23.508 175.052 23.58 175.244 ; 
        RECT 37.764 175.052 37.836 175.244 ; 
        RECT 0.612 179.372 0.684 179.564 ; 
        RECT 14.868 179.372 14.94 179.564 ; 
        RECT 19.836 179.372 19.944 179.564 ; 
        RECT 20.448 179.372 20.592 179.564 ; 
        RECT 23.508 179.372 23.58 179.564 ; 
        RECT 37.764 179.372 37.836 179.564 ; 
        RECT 0.612 183.692 0.684 183.884 ; 
        RECT 14.868 183.692 14.94 183.884 ; 
        RECT 19.836 183.692 19.944 183.884 ; 
        RECT 20.448 183.692 20.592 183.884 ; 
        RECT 23.508 183.692 23.58 183.884 ; 
        RECT 37.764 183.692 37.836 183.884 ; 
        RECT 0.612 188.012 0.684 188.204 ; 
        RECT 14.868 188.012 14.94 188.204 ; 
        RECT 19.836 188.012 19.944 188.204 ; 
        RECT 20.448 188.012 20.592 188.204 ; 
        RECT 23.508 188.012 23.58 188.204 ; 
        RECT 37.764 188.012 37.836 188.204 ; 
        RECT 0.612 192.332 0.684 192.524 ; 
        RECT 14.868 192.332 14.94 192.524 ; 
        RECT 19.836 192.332 19.944 192.524 ; 
        RECT 20.448 192.332 20.592 192.524 ; 
        RECT 23.508 192.332 23.58 192.524 ; 
        RECT 37.764 192.332 37.836 192.524 ; 
        RECT 0.612 196.652 0.684 196.844 ; 
        RECT 14.868 196.652 14.94 196.844 ; 
        RECT 19.836 196.652 19.944 196.844 ; 
        RECT 20.448 196.652 20.592 196.844 ; 
        RECT 23.508 196.652 23.58 196.844 ; 
        RECT 37.764 196.652 37.836 196.844 ; 
        RECT 0.612 200.972 0.684 201.164 ; 
        RECT 14.868 200.972 14.94 201.164 ; 
        RECT 19.836 200.972 19.944 201.164 ; 
        RECT 20.448 200.972 20.592 201.164 ; 
        RECT 23.508 200.972 23.58 201.164 ; 
        RECT 37.764 200.972 37.836 201.164 ; 
        RECT 0.612 205.292 0.684 205.484 ; 
        RECT 14.868 205.292 14.94 205.484 ; 
        RECT 19.836 205.292 19.944 205.484 ; 
        RECT 20.448 205.292 20.592 205.484 ; 
        RECT 23.508 205.292 23.58 205.484 ; 
        RECT 37.764 205.292 37.836 205.484 ; 
        RECT 0.612 209.612 0.684 209.804 ; 
        RECT 14.868 209.612 14.94 209.804 ; 
        RECT 19.836 209.612 19.944 209.804 ; 
        RECT 20.448 209.612 20.592 209.804 ; 
        RECT 23.508 209.612 23.58 209.804 ; 
        RECT 37.764 209.612 37.836 209.804 ; 
        RECT 0.612 213.932 0.684 214.124 ; 
        RECT 14.868 213.932 14.94 214.124 ; 
        RECT 19.836 213.932 19.944 214.124 ; 
        RECT 20.448 213.932 20.592 214.124 ; 
        RECT 23.508 213.932 23.58 214.124 ; 
        RECT 37.764 213.932 37.836 214.124 ; 
        RECT 0.612 218.252 0.684 218.444 ; 
        RECT 14.868 218.252 14.94 218.444 ; 
        RECT 19.836 218.252 19.944 218.444 ; 
        RECT 20.448 218.252 20.592 218.444 ; 
        RECT 23.508 218.252 23.58 218.444 ; 
        RECT 37.764 218.252 37.836 218.444 ; 
        RECT 0.612 222.572 0.684 222.764 ; 
        RECT 14.868 222.572 14.94 222.764 ; 
        RECT 19.836 222.572 19.944 222.764 ; 
        RECT 20.448 222.572 20.592 222.764 ; 
        RECT 23.508 222.572 23.58 222.764 ; 
        RECT 37.764 222.572 37.836 222.764 ; 
        RECT 0.612 226.892 0.684 227.084 ; 
        RECT 14.868 226.892 14.94 227.084 ; 
        RECT 19.836 226.892 19.944 227.084 ; 
        RECT 20.448 226.892 20.592 227.084 ; 
        RECT 23.508 226.892 23.58 227.084 ; 
        RECT 37.764 226.892 37.836 227.084 ; 
        RECT 0.612 231.212 0.684 231.404 ; 
        RECT 14.868 231.212 14.94 231.404 ; 
        RECT 19.836 231.212 19.944 231.404 ; 
        RECT 20.448 231.212 20.592 231.404 ; 
        RECT 23.508 231.212 23.58 231.404 ; 
        RECT 37.764 231.212 37.836 231.404 ; 
        RECT 0.612 235.532 0.684 235.724 ; 
        RECT 14.868 235.532 14.94 235.724 ; 
        RECT 19.836 235.532 19.944 235.724 ; 
        RECT 20.448 235.532 20.592 235.724 ; 
        RECT 23.508 235.532 23.58 235.724 ; 
        RECT 37.764 235.532 37.836 235.724 ; 
        RECT 0.612 239.852 0.684 240.044 ; 
        RECT 14.868 239.852 14.94 240.044 ; 
        RECT 19.836 239.852 19.944 240.044 ; 
        RECT 20.448 239.852 20.592 240.044 ; 
        RECT 23.508 239.852 23.58 240.044 ; 
        RECT 37.764 239.852 37.836 240.044 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.34 109.612 29.412 109.76 ; 
      LAYER M4 ; 
        RECT 29.132 109.644 29.468 109.74 ; 
      LAYER M5 ; 
        RECT 29.328 105.84 29.424 118.8 ; 
      LAYER V3 ; 
        RECT 29.34 109.644 29.412 109.74 ; 
      LAYER V4 ; 
        RECT 29.328 109.644 29.424 109.74 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.476 109.624 28.548 109.772 ; 
      LAYER M4 ; 
        RECT 28.268 109.644 28.604 109.74 ; 
      LAYER M5 ; 
        RECT 28.464 105.84 28.56 118.8 ; 
      LAYER V3 ; 
        RECT 28.476 109.644 28.548 109.74 ; 
      LAYER V4 ; 
        RECT 28.464 109.644 28.56 109.74 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.612 107.308 27.684 107.456 ; 
      LAYER M4 ; 
        RECT 27.404 107.34 27.74 107.436 ; 
      LAYER M5 ; 
        RECT 27.6 105.84 27.696 118.8 ; 
      LAYER V3 ; 
        RECT 27.612 107.34 27.684 107.436 ; 
      LAYER V4 ; 
        RECT 27.6 107.34 27.696 107.436 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.748 108.268 26.82 108.992 ; 
      LAYER M4 ; 
        RECT 26.54 108.876 26.876 108.972 ; 
      LAYER M5 ; 
        RECT 26.736 105.84 26.832 118.8 ; 
      LAYER V3 ; 
        RECT 26.748 108.876 26.82 108.972 ; 
      LAYER V4 ; 
        RECT 26.736 108.876 26.832 108.972 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.884 107.32 25.956 107.588 ; 
      LAYER M4 ; 
        RECT 25.676 107.34 26.012 107.436 ; 
      LAYER M5 ; 
        RECT 25.872 105.84 25.968 118.8 ; 
      LAYER V3 ; 
        RECT 25.884 107.34 25.956 107.436 ; 
      LAYER V4 ; 
        RECT 25.872 107.34 25.968 107.436 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.02 106.252 25.092 107.264 ; 
      LAYER M4 ; 
        RECT 24.812 107.148 25.148 107.244 ; 
      LAYER M5 ; 
        RECT 25.008 105.84 25.104 118.8 ; 
      LAYER V3 ; 
        RECT 25.02 107.148 25.092 107.244 ; 
      LAYER V4 ; 
        RECT 25.008 107.148 25.104 107.244 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.156 110.392 24.228 110.54 ; 
      LAYER M4 ; 
        RECT 23.948 110.412 24.284 110.508 ; 
      LAYER M5 ; 
        RECT 24.144 105.84 24.24 118.8 ; 
      LAYER V3 ; 
        RECT 24.156 110.412 24.228 110.508 ; 
      LAYER V4 ; 
        RECT 24.144 110.412 24.24 110.508 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 20.7 107.32 20.772 107.588 ; 
      LAYER M4 ; 
        RECT 19.564 107.34 20.816 107.436 ; 
      LAYER M5 ; 
        RECT 19.608 105.84 19.704 118.8 ; 
      LAYER V3 ; 
        RECT 20.7 107.34 20.772 107.436 ; 
      LAYER V4 ; 
        RECT 19.608 107.34 19.704 107.436 ; 
    END 
  END ADDRESS[7] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 19.116 106.252 19.188 107.264 ; 
      LAYER M4 ; 
        RECT 18.268 107.148 19.232 107.244 ; 
      LAYER M5 ; 
        RECT 18.312 105.84 18.408 118.8 ; 
      LAYER V3 ; 
        RECT 19.116 107.148 19.188 107.244 ; 
      LAYER V4 ; 
        RECT 18.312 107.148 18.408 107.244 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.948 107.32 16.02 107.588 ; 
      LAYER M4 ; 
        RECT 15.74 107.34 16.076 107.436 ; 
      LAYER M5 ; 
        RECT 15.936 105.84 16.032 118.8 ; 
      LAYER V3 ; 
        RECT 15.948 107.34 16.02 107.436 ; 
      LAYER V4 ; 
        RECT 15.936 107.34 16.032 107.436 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.084 110.776 15.156 110.972 ; 
      LAYER M4 ; 
        RECT 14.876 110.796 15.212 110.892 ; 
      LAYER M5 ; 
        RECT 15.072 105.84 15.168 118.8 ; 
      LAYER V3 ; 
        RECT 15.084 110.796 15.156 110.892 ; 
      LAYER V4 ; 
        RECT 15.072 110.796 15.168 110.892 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.228 106.252 15.3 107.264 ; 
      LAYER M4 ; 
        RECT 14.164 107.148 15.344 107.244 ; 
      LAYER M5 ; 
        RECT 14.208 105.84 14.304 118.8 ; 
      LAYER V3 ; 
        RECT 15.228 107.148 15.3 107.244 ; 
      LAYER V4 ; 
        RECT 14.208 107.148 14.304 107.244 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 13.356 109.612 13.428 109.76 ; 
      LAYER M4 ; 
        RECT 13.148 109.644 13.484 109.74 ; 
      LAYER M5 ; 
        RECT 13.344 105.84 13.44 118.8 ; 
      LAYER V3 ; 
        RECT 13.356 109.644 13.428 109.74 ; 
      LAYER V4 ; 
        RECT 13.344 109.644 13.44 109.74 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 12.492 107.32 12.564 108.236 ; 
      LAYER M4 ; 
        RECT 12.284 107.34 12.62 107.436 ; 
      LAYER M5 ; 
        RECT 12.48 105.84 12.576 118.8 ; 
      LAYER V3 ; 
        RECT 12.492 107.34 12.564 107.436 ; 
      LAYER V4 ; 
        RECT 12.48 107.34 12.576 107.436 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 11.628 106.252 11.7 107.264 ; 
      LAYER M4 ; 
        RECT 11.42 107.148 11.756 107.244 ; 
      LAYER M5 ; 
        RECT 11.616 105.84 11.712 118.8 ; 
      LAYER V3 ; 
        RECT 11.628 107.148 11.7 107.244 ; 
      LAYER V4 ; 
        RECT 11.616 107.148 11.712 107.244 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 10.764 107.308 10.836 107.456 ; 
      LAYER M4 ; 
        RECT 10.556 107.34 10.892 107.436 ; 
      LAYER M5 ; 
        RECT 10.752 105.84 10.848 118.8 ; 
      LAYER V3 ; 
        RECT 10.764 107.34 10.836 107.436 ; 
      LAYER V4 ; 
        RECT 10.752 107.34 10.848 107.436 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 9.9 109.612 9.972 109.76 ; 
      LAYER M4 ; 
        RECT 9.692 109.644 10.028 109.74 ; 
      LAYER M5 ; 
        RECT 9.888 105.84 9.984 118.8 ; 
      LAYER V3 ; 
        RECT 9.9 109.644 9.972 109.74 ; 
      LAYER V4 ; 
        RECT 9.888 109.644 9.984 109.74 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.712 20.544 1.808 ; 
      LAYER M3 ; 
        RECT 20.304 1.51 20.376 2.468 ; 
      LAYER V3 ; 
        RECT 20.304 1.712 20.376 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.328 20.816 1.424 ; 
      LAYER M3 ; 
        RECT 19.404 1.08 19.476 2.7 ; 
      LAYER V3 ; 
        RECT 19.404 1.328 19.476 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 6.032 20.544 6.128 ; 
      LAYER M3 ; 
        RECT 20.304 5.83 20.376 6.788 ; 
      LAYER V3 ; 
        RECT 20.304 6.032 20.376 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 5.648 20.816 5.744 ; 
      LAYER M3 ; 
        RECT 19.404 5.4 19.476 7.02 ; 
      LAYER V3 ; 
        RECT 19.404 5.648 19.476 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 10.352 20.544 10.448 ; 
      LAYER M3 ; 
        RECT 20.304 10.15 20.376 11.108 ; 
      LAYER V3 ; 
        RECT 20.304 10.352 20.376 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 9.968 20.816 10.064 ; 
      LAYER M3 ; 
        RECT 19.404 9.72 19.476 11.34 ; 
      LAYER V3 ; 
        RECT 19.404 9.968 19.476 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.672 20.544 14.768 ; 
      LAYER M3 ; 
        RECT 20.304 14.47 20.376 15.428 ; 
      LAYER V3 ; 
        RECT 20.304 14.672 20.376 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.288 20.816 14.384 ; 
      LAYER M3 ; 
        RECT 19.404 14.04 19.476 15.66 ; 
      LAYER V3 ; 
        RECT 19.404 14.288 19.476 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.992 20.544 19.088 ; 
      LAYER M3 ; 
        RECT 20.304 18.79 20.376 19.748 ; 
      LAYER V3 ; 
        RECT 20.304 18.992 20.376 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.608 20.816 18.704 ; 
      LAYER M3 ; 
        RECT 19.404 18.36 19.476 19.98 ; 
      LAYER V3 ; 
        RECT 19.404 18.608 19.476 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 23.312 20.544 23.408 ; 
      LAYER M3 ; 
        RECT 20.304 23.11 20.376 24.068 ; 
      LAYER V3 ; 
        RECT 20.304 23.312 20.376 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 22.928 20.816 23.024 ; 
      LAYER M3 ; 
        RECT 19.404 22.68 19.476 24.3 ; 
      LAYER V3 ; 
        RECT 19.404 22.928 19.476 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.632 20.544 27.728 ; 
      LAYER M3 ; 
        RECT 20.304 27.43 20.376 28.388 ; 
      LAYER V3 ; 
        RECT 20.304 27.632 20.376 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.248 20.816 27.344 ; 
      LAYER M3 ; 
        RECT 19.404 27 19.476 28.62 ; 
      LAYER V3 ; 
        RECT 19.404 27.248 19.476 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.952 20.544 32.048 ; 
      LAYER M3 ; 
        RECT 20.304 31.75 20.376 32.708 ; 
      LAYER V3 ; 
        RECT 20.304 31.952 20.376 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.568 20.816 31.664 ; 
      LAYER M3 ; 
        RECT 19.404 31.32 19.476 32.94 ; 
      LAYER V3 ; 
        RECT 19.404 31.568 19.476 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 36.272 20.544 36.368 ; 
      LAYER M3 ; 
        RECT 20.304 36.07 20.376 37.028 ; 
      LAYER V3 ; 
        RECT 20.304 36.272 20.376 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 35.888 20.816 35.984 ; 
      LAYER M3 ; 
        RECT 19.404 35.64 19.476 37.26 ; 
      LAYER V3 ; 
        RECT 19.404 35.888 19.476 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 40.592 20.544 40.688 ; 
      LAYER M3 ; 
        RECT 20.304 40.39 20.376 41.348 ; 
      LAYER V3 ; 
        RECT 20.304 40.592 20.376 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 40.208 20.816 40.304 ; 
      LAYER M3 ; 
        RECT 19.404 39.96 19.476 41.58 ; 
      LAYER V3 ; 
        RECT 19.404 40.208 19.476 40.304 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 44.912 20.544 45.008 ; 
      LAYER M3 ; 
        RECT 20.304 44.71 20.376 45.668 ; 
      LAYER V3 ; 
        RECT 20.304 44.912 20.376 45.008 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 44.528 20.816 44.624 ; 
      LAYER M3 ; 
        RECT 19.404 44.28 19.476 45.9 ; 
      LAYER V3 ; 
        RECT 19.404 44.528 19.476 44.624 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 49.232 20.544 49.328 ; 
      LAYER M3 ; 
        RECT 20.304 49.03 20.376 49.988 ; 
      LAYER V3 ; 
        RECT 20.304 49.232 20.376 49.328 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 48.848 20.816 48.944 ; 
      LAYER M3 ; 
        RECT 19.404 48.6 19.476 50.22 ; 
      LAYER V3 ; 
        RECT 19.404 48.848 19.476 48.944 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 53.552 20.544 53.648 ; 
      LAYER M3 ; 
        RECT 20.304 53.35 20.376 54.308 ; 
      LAYER V3 ; 
        RECT 20.304 53.552 20.376 53.648 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 53.168 20.816 53.264 ; 
      LAYER M3 ; 
        RECT 19.404 52.92 19.476 54.54 ; 
      LAYER V3 ; 
        RECT 19.404 53.168 19.476 53.264 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 57.872 20.544 57.968 ; 
      LAYER M3 ; 
        RECT 20.304 57.67 20.376 58.628 ; 
      LAYER V3 ; 
        RECT 20.304 57.872 20.376 57.968 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 57.488 20.816 57.584 ; 
      LAYER M3 ; 
        RECT 19.404 57.24 19.476 58.86 ; 
      LAYER V3 ; 
        RECT 19.404 57.488 19.476 57.584 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 62.192 20.544 62.288 ; 
      LAYER M3 ; 
        RECT 20.304 61.99 20.376 62.948 ; 
      LAYER V3 ; 
        RECT 20.304 62.192 20.376 62.288 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 61.808 20.816 61.904 ; 
      LAYER M3 ; 
        RECT 19.404 61.56 19.476 63.18 ; 
      LAYER V3 ; 
        RECT 19.404 61.808 19.476 61.904 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 66.512 20.544 66.608 ; 
      LAYER M3 ; 
        RECT 20.304 66.31 20.376 67.268 ; 
      LAYER V3 ; 
        RECT 20.304 66.512 20.376 66.608 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 66.128 20.816 66.224 ; 
      LAYER M3 ; 
        RECT 19.404 65.88 19.476 67.5 ; 
      LAYER V3 ; 
        RECT 19.404 66.128 19.476 66.224 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 70.832 20.544 70.928 ; 
      LAYER M3 ; 
        RECT 20.304 70.63 20.376 71.588 ; 
      LAYER V3 ; 
        RECT 20.304 70.832 20.376 70.928 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 70.448 20.816 70.544 ; 
      LAYER M3 ; 
        RECT 19.404 70.2 19.476 71.82 ; 
      LAYER V3 ; 
        RECT 19.404 70.448 19.476 70.544 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 75.152 20.544 75.248 ; 
      LAYER M3 ; 
        RECT 20.304 74.95 20.376 75.908 ; 
      LAYER V3 ; 
        RECT 20.304 75.152 20.376 75.248 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 74.768 20.816 74.864 ; 
      LAYER M3 ; 
        RECT 19.404 74.52 19.476 76.14 ; 
      LAYER V3 ; 
        RECT 19.404 74.768 19.476 74.864 ; 
    END 
  END wd[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 79.472 20.544 79.568 ; 
      LAYER M3 ; 
        RECT 20.304 79.27 20.376 80.228 ; 
      LAYER V3 ; 
        RECT 20.304 79.472 20.376 79.568 ; 
    END 
  END dataout[18] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 79.088 20.816 79.184 ; 
      LAYER M3 ; 
        RECT 19.404 78.84 19.476 80.46 ; 
      LAYER V3 ; 
        RECT 19.404 79.088 19.476 79.184 ; 
    END 
  END wd[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 83.792 20.544 83.888 ; 
      LAYER M3 ; 
        RECT 20.304 83.59 20.376 84.548 ; 
      LAYER V3 ; 
        RECT 20.304 83.792 20.376 83.888 ; 
    END 
  END dataout[19] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 83.408 20.816 83.504 ; 
      LAYER M3 ; 
        RECT 19.404 83.16 19.476 84.78 ; 
      LAYER V3 ; 
        RECT 19.404 83.408 19.476 83.504 ; 
    END 
  END wd[19] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 88.112 20.544 88.208 ; 
      LAYER M3 ; 
        RECT 20.304 87.91 20.376 88.868 ; 
      LAYER V3 ; 
        RECT 20.304 88.112 20.376 88.208 ; 
    END 
  END dataout[20] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 87.728 20.816 87.824 ; 
      LAYER M3 ; 
        RECT 19.404 87.48 19.476 89.1 ; 
      LAYER V3 ; 
        RECT 19.404 87.728 19.476 87.824 ; 
    END 
  END wd[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 92.432 20.544 92.528 ; 
      LAYER M3 ; 
        RECT 20.304 92.23 20.376 93.188 ; 
      LAYER V3 ; 
        RECT 20.304 92.432 20.376 92.528 ; 
    END 
  END dataout[21] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 92.048 20.816 92.144 ; 
      LAYER M3 ; 
        RECT 19.404 91.8 19.476 93.42 ; 
      LAYER V3 ; 
        RECT 19.404 92.048 19.476 92.144 ; 
    END 
  END wd[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 96.752 20.544 96.848 ; 
      LAYER M3 ; 
        RECT 20.304 96.55 20.376 97.508 ; 
      LAYER V3 ; 
        RECT 20.304 96.752 20.376 96.848 ; 
    END 
  END dataout[22] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 96.368 20.816 96.464 ; 
      LAYER M3 ; 
        RECT 19.404 96.12 19.476 97.74 ; 
      LAYER V3 ; 
        RECT 19.404 96.368 19.476 96.464 ; 
    END 
  END wd[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 101.072 20.544 101.168 ; 
      LAYER M3 ; 
        RECT 20.304 100.87 20.376 101.828 ; 
      LAYER V3 ; 
        RECT 20.304 101.072 20.376 101.168 ; 
    END 
  END dataout[23] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 100.688 20.816 100.784 ; 
      LAYER M3 ; 
        RECT 19.404 100.44 19.476 102.06 ; 
      LAYER V3 ; 
        RECT 19.404 100.688 19.476 100.784 ; 
    END 
  END wd[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 137.9 20.544 137.996 ; 
      LAYER M3 ; 
        RECT 20.304 137.698 20.376 138.656 ; 
      LAYER V3 ; 
        RECT 20.304 137.9 20.376 137.996 ; 
    END 
  END dataout[24] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 137.516 20.816 137.612 ; 
      LAYER M3 ; 
        RECT 19.404 137.268 19.476 138.888 ; 
      LAYER V3 ; 
        RECT 19.404 137.516 19.476 137.612 ; 
    END 
  END wd[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 142.22 20.544 142.316 ; 
      LAYER M3 ; 
        RECT 20.304 142.018 20.376 142.976 ; 
      LAYER V3 ; 
        RECT 20.304 142.22 20.376 142.316 ; 
    END 
  END dataout[25] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 141.836 20.816 141.932 ; 
      LAYER M3 ; 
        RECT 19.404 141.588 19.476 143.208 ; 
      LAYER V3 ; 
        RECT 19.404 141.836 19.476 141.932 ; 
    END 
  END wd[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 146.54 20.544 146.636 ; 
      LAYER M3 ; 
        RECT 20.304 146.338 20.376 147.296 ; 
      LAYER V3 ; 
        RECT 20.304 146.54 20.376 146.636 ; 
    END 
  END dataout[26] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 146.156 20.816 146.252 ; 
      LAYER M3 ; 
        RECT 19.404 145.908 19.476 147.528 ; 
      LAYER V3 ; 
        RECT 19.404 146.156 19.476 146.252 ; 
    END 
  END wd[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 150.86 20.544 150.956 ; 
      LAYER M3 ; 
        RECT 20.304 150.658 20.376 151.616 ; 
      LAYER V3 ; 
        RECT 20.304 150.86 20.376 150.956 ; 
    END 
  END dataout[27] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 150.476 20.816 150.572 ; 
      LAYER M3 ; 
        RECT 19.404 150.228 19.476 151.848 ; 
      LAYER V3 ; 
        RECT 19.404 150.476 19.476 150.572 ; 
    END 
  END wd[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 155.18 20.544 155.276 ; 
      LAYER M3 ; 
        RECT 20.304 154.978 20.376 155.936 ; 
      LAYER V3 ; 
        RECT 20.304 155.18 20.376 155.276 ; 
    END 
  END dataout[28] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 154.796 20.816 154.892 ; 
      LAYER M3 ; 
        RECT 19.404 154.548 19.476 156.168 ; 
      LAYER V3 ; 
        RECT 19.404 154.796 19.476 154.892 ; 
    END 
  END wd[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 159.5 20.544 159.596 ; 
      LAYER M3 ; 
        RECT 20.304 159.298 20.376 160.256 ; 
      LAYER V3 ; 
        RECT 20.304 159.5 20.376 159.596 ; 
    END 
  END dataout[29] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 159.116 20.816 159.212 ; 
      LAYER M3 ; 
        RECT 19.404 158.868 19.476 160.488 ; 
      LAYER V3 ; 
        RECT 19.404 159.116 19.476 159.212 ; 
    END 
  END wd[29] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 163.82 20.544 163.916 ; 
      LAYER M3 ; 
        RECT 20.304 163.618 20.376 164.576 ; 
      LAYER V3 ; 
        RECT 20.304 163.82 20.376 163.916 ; 
    END 
  END dataout[30] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 163.436 20.816 163.532 ; 
      LAYER M3 ; 
        RECT 19.404 163.188 19.476 164.808 ; 
      LAYER V3 ; 
        RECT 19.404 163.436 19.476 163.532 ; 
    END 
  END wd[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 168.14 20.544 168.236 ; 
      LAYER M3 ; 
        RECT 20.304 167.938 20.376 168.896 ; 
      LAYER V3 ; 
        RECT 20.304 168.14 20.376 168.236 ; 
    END 
  END dataout[31] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 167.756 20.816 167.852 ; 
      LAYER M3 ; 
        RECT 19.404 167.508 19.476 169.128 ; 
      LAYER V3 ; 
        RECT 19.404 167.756 19.476 167.852 ; 
    END 
  END wd[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 172.46 20.544 172.556 ; 
      LAYER M3 ; 
        RECT 20.304 172.258 20.376 173.216 ; 
      LAYER V3 ; 
        RECT 20.304 172.46 20.376 172.556 ; 
    END 
  END dataout[32] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 172.076 20.816 172.172 ; 
      LAYER M3 ; 
        RECT 19.404 171.828 19.476 173.448 ; 
      LAYER V3 ; 
        RECT 19.404 172.076 19.476 172.172 ; 
    END 
  END wd[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 176.78 20.544 176.876 ; 
      LAYER M3 ; 
        RECT 20.304 176.578 20.376 177.536 ; 
      LAYER V3 ; 
        RECT 20.304 176.78 20.376 176.876 ; 
    END 
  END dataout[33] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 176.396 20.816 176.492 ; 
      LAYER M3 ; 
        RECT 19.404 176.148 19.476 177.768 ; 
      LAYER V3 ; 
        RECT 19.404 176.396 19.476 176.492 ; 
    END 
  END wd[33] 
  PIN dataout[34] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 181.1 20.544 181.196 ; 
      LAYER M3 ; 
        RECT 20.304 180.898 20.376 181.856 ; 
      LAYER V3 ; 
        RECT 20.304 181.1 20.376 181.196 ; 
    END 
  END dataout[34] 
  PIN wd[34] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 180.716 20.816 180.812 ; 
      LAYER M3 ; 
        RECT 19.404 180.468 19.476 182.088 ; 
      LAYER V3 ; 
        RECT 19.404 180.716 19.476 180.812 ; 
    END 
  END wd[34] 
  PIN dataout[35] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 185.42 20.544 185.516 ; 
      LAYER M3 ; 
        RECT 20.304 185.218 20.376 186.176 ; 
      LAYER V3 ; 
        RECT 20.304 185.42 20.376 185.516 ; 
    END 
  END dataout[35] 
  PIN wd[35] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 185.036 20.816 185.132 ; 
      LAYER M3 ; 
        RECT 19.404 184.788 19.476 186.408 ; 
      LAYER V3 ; 
        RECT 19.404 185.036 19.476 185.132 ; 
    END 
  END wd[35] 
  PIN dataout[36] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 189.74 20.544 189.836 ; 
      LAYER M3 ; 
        RECT 20.304 189.538 20.376 190.496 ; 
      LAYER V3 ; 
        RECT 20.304 189.74 20.376 189.836 ; 
    END 
  END dataout[36] 
  PIN wd[36] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 189.356 20.816 189.452 ; 
      LAYER M3 ; 
        RECT 19.404 189.108 19.476 190.728 ; 
      LAYER V3 ; 
        RECT 19.404 189.356 19.476 189.452 ; 
    END 
  END wd[36] 
  PIN dataout[37] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 194.06 20.544 194.156 ; 
      LAYER M3 ; 
        RECT 20.304 193.858 20.376 194.816 ; 
      LAYER V3 ; 
        RECT 20.304 194.06 20.376 194.156 ; 
    END 
  END dataout[37] 
  PIN wd[37] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 193.676 20.816 193.772 ; 
      LAYER M3 ; 
        RECT 19.404 193.428 19.476 195.048 ; 
      LAYER V3 ; 
        RECT 19.404 193.676 19.476 193.772 ; 
    END 
  END wd[37] 
  PIN dataout[38] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 198.38 20.544 198.476 ; 
      LAYER M3 ; 
        RECT 20.304 198.178 20.376 199.136 ; 
      LAYER V3 ; 
        RECT 20.304 198.38 20.376 198.476 ; 
    END 
  END dataout[38] 
  PIN wd[38] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 197.996 20.816 198.092 ; 
      LAYER M3 ; 
        RECT 19.404 197.748 19.476 199.368 ; 
      LAYER V3 ; 
        RECT 19.404 197.996 19.476 198.092 ; 
    END 
  END wd[38] 
  PIN dataout[39] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 202.7 20.544 202.796 ; 
      LAYER M3 ; 
        RECT 20.304 202.498 20.376 203.456 ; 
      LAYER V3 ; 
        RECT 20.304 202.7 20.376 202.796 ; 
    END 
  END dataout[39] 
  PIN wd[39] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 202.316 20.816 202.412 ; 
      LAYER M3 ; 
        RECT 19.404 202.068 19.476 203.688 ; 
      LAYER V3 ; 
        RECT 19.404 202.316 19.476 202.412 ; 
    END 
  END wd[39] 
  PIN dataout[40] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 207.02 20.544 207.116 ; 
      LAYER M3 ; 
        RECT 20.304 206.818 20.376 207.776 ; 
      LAYER V3 ; 
        RECT 20.304 207.02 20.376 207.116 ; 
    END 
  END dataout[40] 
  PIN wd[40] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 206.636 20.816 206.732 ; 
      LAYER M3 ; 
        RECT 19.404 206.388 19.476 208.008 ; 
      LAYER V3 ; 
        RECT 19.404 206.636 19.476 206.732 ; 
    END 
  END wd[40] 
  PIN dataout[41] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 211.34 20.544 211.436 ; 
      LAYER M3 ; 
        RECT 20.304 211.138 20.376 212.096 ; 
      LAYER V3 ; 
        RECT 20.304 211.34 20.376 211.436 ; 
    END 
  END dataout[41] 
  PIN wd[41] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 210.956 20.816 211.052 ; 
      LAYER M3 ; 
        RECT 19.404 210.708 19.476 212.328 ; 
      LAYER V3 ; 
        RECT 19.404 210.956 19.476 211.052 ; 
    END 
  END wd[41] 
  PIN dataout[42] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 215.66 20.544 215.756 ; 
      LAYER M3 ; 
        RECT 20.304 215.458 20.376 216.416 ; 
      LAYER V3 ; 
        RECT 20.304 215.66 20.376 215.756 ; 
    END 
  END dataout[42] 
  PIN wd[42] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 215.276 20.816 215.372 ; 
      LAYER M3 ; 
        RECT 19.404 215.028 19.476 216.648 ; 
      LAYER V3 ; 
        RECT 19.404 215.276 19.476 215.372 ; 
    END 
  END wd[42] 
  PIN dataout[43] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 219.98 20.544 220.076 ; 
      LAYER M3 ; 
        RECT 20.304 219.778 20.376 220.736 ; 
      LAYER V3 ; 
        RECT 20.304 219.98 20.376 220.076 ; 
    END 
  END dataout[43] 
  PIN wd[43] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 219.596 20.816 219.692 ; 
      LAYER M3 ; 
        RECT 19.404 219.348 19.476 220.968 ; 
      LAYER V3 ; 
        RECT 19.404 219.596 19.476 219.692 ; 
    END 
  END wd[43] 
  PIN dataout[44] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 224.3 20.544 224.396 ; 
      LAYER M3 ; 
        RECT 20.304 224.098 20.376 225.056 ; 
      LAYER V3 ; 
        RECT 20.304 224.3 20.376 224.396 ; 
    END 
  END dataout[44] 
  PIN wd[44] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 223.916 20.816 224.012 ; 
      LAYER M3 ; 
        RECT 19.404 223.668 19.476 225.288 ; 
      LAYER V3 ; 
        RECT 19.404 223.916 19.476 224.012 ; 
    END 
  END wd[44] 
  PIN dataout[45] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 228.62 20.544 228.716 ; 
      LAYER M3 ; 
        RECT 20.304 228.418 20.376 229.376 ; 
      LAYER V3 ; 
        RECT 20.304 228.62 20.376 228.716 ; 
    END 
  END dataout[45] 
  PIN wd[45] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 228.236 20.816 228.332 ; 
      LAYER M3 ; 
        RECT 19.404 227.988 19.476 229.608 ; 
      LAYER V3 ; 
        RECT 19.404 228.236 19.476 228.332 ; 
    END 
  END wd[45] 
  PIN dataout[46] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 232.94 20.544 233.036 ; 
      LAYER M3 ; 
        RECT 20.304 232.738 20.376 233.696 ; 
      LAYER V3 ; 
        RECT 20.304 232.94 20.376 233.036 ; 
    END 
  END dataout[46] 
  PIN wd[46] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 232.556 20.816 232.652 ; 
      LAYER M3 ; 
        RECT 19.404 232.308 19.476 233.928 ; 
      LAYER V3 ; 
        RECT 19.404 232.556 19.476 232.652 ; 
    END 
  END wd[46] 
  PIN dataout[47] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 237.26 20.544 237.356 ; 
      LAYER M3 ; 
        RECT 20.304 237.058 20.376 238.016 ; 
      LAYER V3 ; 
        RECT 20.304 237.26 20.376 237.356 ; 
    END 
  END dataout[47] 
  PIN wd[47] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 236.876 20.816 236.972 ; 
      LAYER M3 ; 
        RECT 19.404 236.628 19.476 238.248 ; 
      LAYER V3 ; 
        RECT 19.404 236.876 19.476 236.972 ; 
    END 
  END wd[47] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.652 38.448 139.266 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
        RECT 0 180.414 38.448 184.788 ; 
        RECT 0 184.734 38.448 189.108 ; 
        RECT 0 189.054 38.448 193.428 ; 
        RECT 0 193.374 38.448 197.748 ; 
        RECT 0 197.694 38.448 202.068 ; 
        RECT 0 202.014 38.448 206.388 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.652 38.448 139.266 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
        RECT 0 180.414 38.448 184.788 ; 
        RECT 0 184.734 38.448 189.108 ; 
        RECT 0 189.054 38.448 193.428 ; 
        RECT 0 193.374 38.448 197.748 ; 
        RECT 0 197.694 38.448 202.068 ; 
        RECT 0 202.014 38.448 206.388 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
  LAYER V1 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.652 38.448 139.266 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
        RECT 0 180.414 38.448 184.788 ; 
        RECT 0 184.734 38.448 189.108 ; 
        RECT 0 189.054 38.448 193.428 ; 
        RECT 0 193.374 38.448 197.748 ; 
        RECT 0 197.694 38.448 202.068 ; 
        RECT 0 202.014 38.448 206.388 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
  LAYER V2 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.652 38.448 139.266 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
        RECT 0 180.414 38.448 184.788 ; 
        RECT 0 184.734 38.448 189.108 ; 
        RECT 0 189.054 38.448 193.428 ; 
        RECT 0 193.374 38.448 197.748 ; 
        RECT 0 197.694 38.448 202.068 ; 
        RECT 0 202.014 38.448 206.388 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
  LAYER M3 ; 
      RECT 20.952 1.38 21.024 5.122 ; 
      RECT 20.808 1.38 20.88 5.122 ; 
      RECT 20.664 3.688 20.736 4.978 ; 
      RECT 20.196 4.476 20.268 4.914 ; 
      RECT 20.16 1.51 20.232 2.468 ; 
      RECT 20.016 3.834 20.088 4.448 ; 
      RECT 19.692 3.936 19.764 4.968 ; 
      RECT 17.532 1.38 17.604 5.122 ; 
      RECT 17.388 1.38 17.46 5.122 ; 
      RECT 17.244 2.104 17.316 4.376 ; 
      RECT 20.952 5.7 21.024 9.442 ; 
      RECT 20.808 5.7 20.88 9.442 ; 
      RECT 20.664 8.008 20.736 9.298 ; 
      RECT 20.196 8.796 20.268 9.234 ; 
      RECT 20.16 5.83 20.232 6.788 ; 
      RECT 20.016 8.154 20.088 8.768 ; 
      RECT 19.692 8.256 19.764 9.288 ; 
      RECT 17.532 5.7 17.604 9.442 ; 
      RECT 17.388 5.7 17.46 9.442 ; 
      RECT 17.244 6.424 17.316 8.696 ; 
      RECT 20.952 10.02 21.024 13.762 ; 
      RECT 20.808 10.02 20.88 13.762 ; 
      RECT 20.664 12.328 20.736 13.618 ; 
      RECT 20.196 13.116 20.268 13.554 ; 
      RECT 20.16 10.15 20.232 11.108 ; 
      RECT 20.016 12.474 20.088 13.088 ; 
      RECT 19.692 12.576 19.764 13.608 ; 
      RECT 17.532 10.02 17.604 13.762 ; 
      RECT 17.388 10.02 17.46 13.762 ; 
      RECT 17.244 10.744 17.316 13.016 ; 
      RECT 20.952 14.34 21.024 18.082 ; 
      RECT 20.808 14.34 20.88 18.082 ; 
      RECT 20.664 16.648 20.736 17.938 ; 
      RECT 20.196 17.436 20.268 17.874 ; 
      RECT 20.16 14.47 20.232 15.428 ; 
      RECT 20.016 16.794 20.088 17.408 ; 
      RECT 19.692 16.896 19.764 17.928 ; 
      RECT 17.532 14.34 17.604 18.082 ; 
      RECT 17.388 14.34 17.46 18.082 ; 
      RECT 17.244 15.064 17.316 17.336 ; 
      RECT 20.952 18.66 21.024 22.402 ; 
      RECT 20.808 18.66 20.88 22.402 ; 
      RECT 20.664 20.968 20.736 22.258 ; 
      RECT 20.196 21.756 20.268 22.194 ; 
      RECT 20.16 18.79 20.232 19.748 ; 
      RECT 20.016 21.114 20.088 21.728 ; 
      RECT 19.692 21.216 19.764 22.248 ; 
      RECT 17.532 18.66 17.604 22.402 ; 
      RECT 17.388 18.66 17.46 22.402 ; 
      RECT 17.244 19.384 17.316 21.656 ; 
      RECT 20.952 22.98 21.024 26.722 ; 
      RECT 20.808 22.98 20.88 26.722 ; 
      RECT 20.664 25.288 20.736 26.578 ; 
      RECT 20.196 26.076 20.268 26.514 ; 
      RECT 20.16 23.11 20.232 24.068 ; 
      RECT 20.016 25.434 20.088 26.048 ; 
      RECT 19.692 25.536 19.764 26.568 ; 
      RECT 17.532 22.98 17.604 26.722 ; 
      RECT 17.388 22.98 17.46 26.722 ; 
      RECT 17.244 23.704 17.316 25.976 ; 
      RECT 20.952 27.3 21.024 31.042 ; 
      RECT 20.808 27.3 20.88 31.042 ; 
      RECT 20.664 29.608 20.736 30.898 ; 
      RECT 20.196 30.396 20.268 30.834 ; 
      RECT 20.16 27.43 20.232 28.388 ; 
      RECT 20.016 29.754 20.088 30.368 ; 
      RECT 19.692 29.856 19.764 30.888 ; 
      RECT 17.532 27.3 17.604 31.042 ; 
      RECT 17.388 27.3 17.46 31.042 ; 
      RECT 17.244 28.024 17.316 30.296 ; 
      RECT 20.952 31.62 21.024 35.362 ; 
      RECT 20.808 31.62 20.88 35.362 ; 
      RECT 20.664 33.928 20.736 35.218 ; 
      RECT 20.196 34.716 20.268 35.154 ; 
      RECT 20.16 31.75 20.232 32.708 ; 
      RECT 20.016 34.074 20.088 34.688 ; 
      RECT 19.692 34.176 19.764 35.208 ; 
      RECT 17.532 31.62 17.604 35.362 ; 
      RECT 17.388 31.62 17.46 35.362 ; 
      RECT 17.244 32.344 17.316 34.616 ; 
      RECT 20.952 35.94 21.024 39.682 ; 
      RECT 20.808 35.94 20.88 39.682 ; 
      RECT 20.664 38.248 20.736 39.538 ; 
      RECT 20.196 39.036 20.268 39.474 ; 
      RECT 20.16 36.07 20.232 37.028 ; 
      RECT 20.016 38.394 20.088 39.008 ; 
      RECT 19.692 38.496 19.764 39.528 ; 
      RECT 17.532 35.94 17.604 39.682 ; 
      RECT 17.388 35.94 17.46 39.682 ; 
      RECT 17.244 36.664 17.316 38.936 ; 
      RECT 20.952 40.26 21.024 44.002 ; 
      RECT 20.808 40.26 20.88 44.002 ; 
      RECT 20.664 42.568 20.736 43.858 ; 
      RECT 20.196 43.356 20.268 43.794 ; 
      RECT 20.16 40.39 20.232 41.348 ; 
      RECT 20.016 42.714 20.088 43.328 ; 
      RECT 19.692 42.816 19.764 43.848 ; 
      RECT 17.532 40.26 17.604 44.002 ; 
      RECT 17.388 40.26 17.46 44.002 ; 
      RECT 17.244 40.984 17.316 43.256 ; 
      RECT 20.952 44.58 21.024 48.322 ; 
      RECT 20.808 44.58 20.88 48.322 ; 
      RECT 20.664 46.888 20.736 48.178 ; 
      RECT 20.196 47.676 20.268 48.114 ; 
      RECT 20.16 44.71 20.232 45.668 ; 
      RECT 20.016 47.034 20.088 47.648 ; 
      RECT 19.692 47.136 19.764 48.168 ; 
      RECT 17.532 44.58 17.604 48.322 ; 
      RECT 17.388 44.58 17.46 48.322 ; 
      RECT 17.244 45.304 17.316 47.576 ; 
      RECT 20.952 48.9 21.024 52.642 ; 
      RECT 20.808 48.9 20.88 52.642 ; 
      RECT 20.664 51.208 20.736 52.498 ; 
      RECT 20.196 51.996 20.268 52.434 ; 
      RECT 20.16 49.03 20.232 49.988 ; 
      RECT 20.016 51.354 20.088 51.968 ; 
      RECT 19.692 51.456 19.764 52.488 ; 
      RECT 17.532 48.9 17.604 52.642 ; 
      RECT 17.388 48.9 17.46 52.642 ; 
      RECT 17.244 49.624 17.316 51.896 ; 
      RECT 20.952 53.22 21.024 56.962 ; 
      RECT 20.808 53.22 20.88 56.962 ; 
      RECT 20.664 55.528 20.736 56.818 ; 
      RECT 20.196 56.316 20.268 56.754 ; 
      RECT 20.16 53.35 20.232 54.308 ; 
      RECT 20.016 55.674 20.088 56.288 ; 
      RECT 19.692 55.776 19.764 56.808 ; 
      RECT 17.532 53.22 17.604 56.962 ; 
      RECT 17.388 53.22 17.46 56.962 ; 
      RECT 17.244 53.944 17.316 56.216 ; 
      RECT 20.952 57.54 21.024 61.282 ; 
      RECT 20.808 57.54 20.88 61.282 ; 
      RECT 20.664 59.848 20.736 61.138 ; 
      RECT 20.196 60.636 20.268 61.074 ; 
      RECT 20.16 57.67 20.232 58.628 ; 
      RECT 20.016 59.994 20.088 60.608 ; 
      RECT 19.692 60.096 19.764 61.128 ; 
      RECT 17.532 57.54 17.604 61.282 ; 
      RECT 17.388 57.54 17.46 61.282 ; 
      RECT 17.244 58.264 17.316 60.536 ; 
      RECT 20.952 61.86 21.024 65.602 ; 
      RECT 20.808 61.86 20.88 65.602 ; 
      RECT 20.664 64.168 20.736 65.458 ; 
      RECT 20.196 64.956 20.268 65.394 ; 
      RECT 20.16 61.99 20.232 62.948 ; 
      RECT 20.016 64.314 20.088 64.928 ; 
      RECT 19.692 64.416 19.764 65.448 ; 
      RECT 17.532 61.86 17.604 65.602 ; 
      RECT 17.388 61.86 17.46 65.602 ; 
      RECT 17.244 62.584 17.316 64.856 ; 
      RECT 20.952 66.18 21.024 69.922 ; 
      RECT 20.808 66.18 20.88 69.922 ; 
      RECT 20.664 68.488 20.736 69.778 ; 
      RECT 20.196 69.276 20.268 69.714 ; 
      RECT 20.16 66.31 20.232 67.268 ; 
      RECT 20.016 68.634 20.088 69.248 ; 
      RECT 19.692 68.736 19.764 69.768 ; 
      RECT 17.532 66.18 17.604 69.922 ; 
      RECT 17.388 66.18 17.46 69.922 ; 
      RECT 17.244 66.904 17.316 69.176 ; 
      RECT 20.952 70.5 21.024 74.242 ; 
      RECT 20.808 70.5 20.88 74.242 ; 
      RECT 20.664 72.808 20.736 74.098 ; 
      RECT 20.196 73.596 20.268 74.034 ; 
      RECT 20.16 70.63 20.232 71.588 ; 
      RECT 20.016 72.954 20.088 73.568 ; 
      RECT 19.692 73.056 19.764 74.088 ; 
      RECT 17.532 70.5 17.604 74.242 ; 
      RECT 17.388 70.5 17.46 74.242 ; 
      RECT 17.244 71.224 17.316 73.496 ; 
      RECT 20.952 74.82 21.024 78.562 ; 
      RECT 20.808 74.82 20.88 78.562 ; 
      RECT 20.664 77.128 20.736 78.418 ; 
      RECT 20.196 77.916 20.268 78.354 ; 
      RECT 20.16 74.95 20.232 75.908 ; 
      RECT 20.016 77.274 20.088 77.888 ; 
      RECT 19.692 77.376 19.764 78.408 ; 
      RECT 17.532 74.82 17.604 78.562 ; 
      RECT 17.388 74.82 17.46 78.562 ; 
      RECT 17.244 75.544 17.316 77.816 ; 
      RECT 20.952 79.14 21.024 82.882 ; 
      RECT 20.808 79.14 20.88 82.882 ; 
      RECT 20.664 81.448 20.736 82.738 ; 
      RECT 20.196 82.236 20.268 82.674 ; 
      RECT 20.16 79.27 20.232 80.228 ; 
      RECT 20.016 81.594 20.088 82.208 ; 
      RECT 19.692 81.696 19.764 82.728 ; 
      RECT 17.532 79.14 17.604 82.882 ; 
      RECT 17.388 79.14 17.46 82.882 ; 
      RECT 17.244 79.864 17.316 82.136 ; 
      RECT 20.952 83.46 21.024 87.202 ; 
      RECT 20.808 83.46 20.88 87.202 ; 
      RECT 20.664 85.768 20.736 87.058 ; 
      RECT 20.196 86.556 20.268 86.994 ; 
      RECT 20.16 83.59 20.232 84.548 ; 
      RECT 20.016 85.914 20.088 86.528 ; 
      RECT 19.692 86.016 19.764 87.048 ; 
      RECT 17.532 83.46 17.604 87.202 ; 
      RECT 17.388 83.46 17.46 87.202 ; 
      RECT 17.244 84.184 17.316 86.456 ; 
      RECT 20.952 87.78 21.024 91.522 ; 
      RECT 20.808 87.78 20.88 91.522 ; 
      RECT 20.664 90.088 20.736 91.378 ; 
      RECT 20.196 90.876 20.268 91.314 ; 
      RECT 20.16 87.91 20.232 88.868 ; 
      RECT 20.016 90.234 20.088 90.848 ; 
      RECT 19.692 90.336 19.764 91.368 ; 
      RECT 17.532 87.78 17.604 91.522 ; 
      RECT 17.388 87.78 17.46 91.522 ; 
      RECT 17.244 88.504 17.316 90.776 ; 
      RECT 20.952 92.1 21.024 95.842 ; 
      RECT 20.808 92.1 20.88 95.842 ; 
      RECT 20.664 94.408 20.736 95.698 ; 
      RECT 20.196 95.196 20.268 95.634 ; 
      RECT 20.16 92.23 20.232 93.188 ; 
      RECT 20.016 94.554 20.088 95.168 ; 
      RECT 19.692 94.656 19.764 95.688 ; 
      RECT 17.532 92.1 17.604 95.842 ; 
      RECT 17.388 92.1 17.46 95.842 ; 
      RECT 17.244 92.824 17.316 95.096 ; 
      RECT 20.952 96.42 21.024 100.162 ; 
      RECT 20.808 96.42 20.88 100.162 ; 
      RECT 20.664 98.728 20.736 100.018 ; 
      RECT 20.196 99.516 20.268 99.954 ; 
      RECT 20.16 96.55 20.232 97.508 ; 
      RECT 20.016 98.874 20.088 99.488 ; 
      RECT 19.692 98.976 19.764 100.008 ; 
      RECT 17.532 96.42 17.604 100.162 ; 
      RECT 17.388 96.42 17.46 100.162 ; 
      RECT 17.244 97.144 17.316 99.416 ; 
      RECT 20.952 100.74 21.024 104.482 ; 
      RECT 20.808 100.74 20.88 104.482 ; 
      RECT 20.664 103.048 20.736 104.338 ; 
      RECT 20.196 103.836 20.268 104.274 ; 
      RECT 20.16 100.87 20.232 101.828 ; 
      RECT 20.016 103.194 20.088 103.808 ; 
      RECT 19.692 103.296 19.764 104.328 ; 
      RECT 17.532 100.74 17.604 104.482 ; 
      RECT 17.388 100.74 17.46 104.482 ; 
      RECT 17.244 101.464 17.316 103.736 ; 
      RECT 37.62 119.824 37.692 137.246 ; 
      RECT 37.476 114.564 37.548 114.84 ; 
      RECT 37.476 121.796 37.548 123.654 ; 
      RECT 37.332 104.546 37.404 137.374 ; 
      RECT 37.188 119.624 37.26 122.714 ; 
      RECT 37.188 122.9188 37.26 124.884 ; 
      RECT 37.188 125.084 37.26 126.57 ; 
      RECT 37.188 126.822 37.26 130.068 ; 
      RECT 37.044 119.966 37.116 122.534 ; 
      RECT 37.044 125.244 37.116 127.372 ; 
      RECT 36.9 104.546 36.972 105.946 ; 
      RECT 36.468 104.546 36.54 105.946 ; 
      RECT 36.036 104.546 36.108 105.946 ; 
      RECT 35.604 104.546 35.676 105.946 ; 
      RECT 35.172 104.546 35.244 105.946 ; 
      RECT 34.74 104.546 34.812 105.946 ; 
      RECT 34.308 104.546 34.38 105.946 ; 
      RECT 33.876 104.546 33.948 105.946 ; 
      RECT 33.444 104.546 33.516 105.946 ; 
      RECT 33.012 104.546 33.084 105.946 ; 
      RECT 32.58 104.546 32.652 105.946 ; 
      RECT 32.148 104.546 32.22 105.946 ; 
      RECT 31.716 104.546 31.788 105.946 ; 
      RECT 31.284 104.546 31.356 105.946 ; 
      RECT 30.852 104.546 30.924 105.946 ; 
      RECT 30.42 104.546 30.492 105.946 ; 
      RECT 29.988 104.546 30.06 105.946 ; 
      RECT 29.556 104.546 29.628 105.946 ; 
      RECT 29.124 104.546 29.196 105.946 ; 
      RECT 28.692 104.546 28.764 105.946 ; 
      RECT 28.26 104.546 28.332 105.946 ; 
      RECT 27.828 104.546 27.9 105.946 ; 
      RECT 27.396 104.546 27.468 105.946 ; 
      RECT 26.964 104.546 27.036 105.946 ; 
      RECT 26.532 104.546 26.604 105.946 ; 
      RECT 26.1 104.546 26.172 105.946 ; 
      RECT 25.668 104.546 25.74 105.946 ; 
      RECT 25.236 104.546 25.308 105.946 ; 
      RECT 24.804 104.546 24.876 105.946 ; 
      RECT 24.372 104.546 24.444 105.946 ; 
      RECT 24.228 119.7 24.3 122.5188 ; 
      RECT 24.228 125.488 24.3 130.212 ; 
      RECT 24.156 107.188 24.228 109.892 ; 
      RECT 24.156 112.876 24.228 114.068 ; 
      RECT 24.084 119.954 24.156 122.714 ; 
      RECT 24.084 122.918 24.156 126.884 ; 
      RECT 24.084 127.004 24.156 130.14 ; 
      RECT 23.94 104.546 24.012 137.374 ; 
      RECT 23.796 121.044 23.868 121.376 ; 
      RECT 23.724 107.62 23.796 110.144 ; 
      RECT 23.724 111.796 23.796 112.556 ; 
      RECT 23.724 115.324 23.796 115.52 ; 
      RECT 23.652 119.824 23.724 137.264 ; 
      RECT 23.292 106.108 23.364 109.316 ; 
      RECT 23.292 111.508 23.364 113.78 ; 
      RECT 23.148 111.796 23.22 113.276 ; 
      RECT 23.004 109.204 23.076 109.748 ; 
      RECT 23.004 113.164 23.076 114.068 ; 
      RECT 23.004 118.132 23.076 118.388 ; 
      RECT 22.86 109.612 22.932 109.76 ; 
      RECT 22.86 116.116 22.932 116.288 ; 
      RECT 22.86 118.252 22.932 118.4 ; 
      RECT 22.716 110.86 22.788 112.844 ; 
      RECT 22.716 113.02 22.788 113.78 ; 
      RECT 22.716 116.86 22.788 118.1 ; 
      RECT 22.572 125.98 22.644 128.9 ; 
      RECT 22.572 130.3 22.644 133.22 ; 
      RECT 21.276 109.348 21.348 110.54 ; 
      RECT 21.276 114.1 21.348 114.356 ; 
      RECT 21.276 115.18 21.348 117.02 ; 
      RECT 21.276 119.98 21.348 120.128 ; 
      RECT 21.276 128.14 21.348 129.332 ; 
      RECT 21.132 109.636 21.204 111.656 ; 
      RECT 21.132 112.732 21.204 115.94 ; 
      RECT 21.132 120.112 21.204 121.196 ; 
      RECT 21.132 121.516 21.204 122.42 ; 
      RECT 20.988 109.348 21.06 112.052 ; 
      RECT 20.988 112.444 21.06 113.78 ; 
      RECT 20.988 114.604 21.06 115.148 ; 
      RECT 20.988 117.34 21.06 120.548 ; 
      RECT 20.988 122.284 21.06 122.432 ; 
      RECT 20.988 130.948 21.06 132.284 ; 
      RECT 20.844 110.284 20.916 110.828 ; 
      RECT 20.844 117.844 20.916 121.772 ; 
      RECT 20.844 123.532 20.916 124.724 ; 
      RECT 20.844 130.3 20.916 131.348 ; 
      RECT 20.7 106.54 20.772 107.156 ; 
      RECT 20.7 109.78 20.772 116.924 ; 
      RECT 20.7 121.084 20.772 130.412 ; 
      RECT 20.7 131.236 20.772 135.668 ; 
      RECT 19.548 107.62 19.62 108.668 ; 
      RECT 19.548 109.204 19.62 109.46 ; 
      RECT 19.548 109.78 19.62 110.684 ; 
      RECT 19.548 110.86 19.62 111.62 ; 
      RECT 19.548 111.94 19.62 122.42 ; 
      RECT 19.548 122.596 19.62 127.82 ; 
      RECT 19.548 132.172 19.62 133.22 ; 
      RECT 19.404 111.616 19.476 112.7 ; 
      RECT 19.404 113.02 19.476 116.372 ; 
      RECT 19.404 117.052 19.476 120.404 ; 
      RECT 19.404 120.58 19.476 125.66 ; 
      RECT 19.404 126.484 19.476 127.172 ; 
      RECT 19.404 130.012 19.476 134.3 ; 
      RECT 19.26 111.94 19.332 113.024 ; 
      RECT 19.26 113.644 19.332 113.792 ; 
      RECT 19.26 116.764 19.332 120.692 ; 
      RECT 19.26 121.66 19.332 123.5 ; 
      RECT 19.26 124.9 19.332 127.856 ; 
      RECT 19.116 108.412 19.188 112.7 ; 
      RECT 19.116 119.068 19.188 119.936 ; 
      RECT 19.116 124.612 19.188 125.804 ; 
      RECT 18.972 111.004 19.044 112.844 ; 
      RECT 18.972 117.34 19.044 118.1 ; 
      RECT 18.972 118.264 19.044 118.412 ; 
      RECT 18.972 119.356 19.044 120.692 ; 
      RECT 18.972 121.228 19.044 126.596 ; 
      RECT 18.972 127.024 19.044 131.492 ; 
      RECT 18.828 108.7 18.9 109.46 ; 
      RECT 18.828 110.284 18.9 110.828 ; 
      RECT 18.828 111.94 18.9 124.58 ; 
      RECT 18.828 124.9 18.9 126.74 ; 
      RECT 18.828 129.22 18.9 131.06 ; 
      RECT 18.828 134.476 18.9 135.38 ; 
      RECT 18.684 104.652 18.756 105.268 ; 
      RECT 18.684 136.696 18.756 137.312 ; 
      RECT 18.54 104.652 18.612 104.852 ; 
      RECT 18.252 104.652 18.324 104.938 ; 
      RECT 18.252 136.974 18.324 137.374 ; 
      RECT 17.676 110.716 17.748 111.476 ; 
      RECT 17.676 113.668 17.748 115.148 ; 
      RECT 17.676 121.516 17.748 122.42 ; 
      RECT 17.676 123.676 17.748 128.252 ; 
      RECT 17.676 131.38 17.748 133.22 ; 
      RECT 17.676 135.532 17.748 135.68 ; 
      RECT 17.532 106.54 17.604 108.524 ; 
      RECT 17.532 122.86 17.604 123.008 ; 
      RECT 17.532 127.168 17.604 130.412 ; 
      RECT 17.388 108.412 17.46 109.46 ; 
      RECT 17.388 110.572 17.46 111.908 ; 
      RECT 17.388 112.732 17.46 113.132 ; 
      RECT 17.388 116.26 17.46 127.316 ; 
      RECT 17.388 127.852 17.46 128.756 ; 
      RECT 17.244 107.044 17.316 111.62 ; 
      RECT 17.244 125.98 17.316 126.74 ; 
      RECT 17.244 129.196 17.316 129.344 ; 
      RECT 17.244 130.3 17.316 133.508 ; 
      RECT 17.1 110.86 17.172 114.86 ; 
      RECT 17.1 128.62 17.172 128.768 ; 
      RECT 16.956 107.62 17.028 107.732 ; 
      RECT 15.66 109.204 15.732 110.828 ; 
      RECT 15.372 109.348 15.444 111.764 ; 
      RECT 15.228 108.7 15.3 108.956 ; 
      RECT 15.084 104.864 15.156 105.068 ; 
      RECT 15.084 117.34 15.156 118.1 ; 
      RECT 15.084 119.824 15.156 137.264 ; 
      RECT 14.724 119.824 14.796 137.264 ; 
      RECT 14.652 106.54 14.724 107.3 ; 
      RECT 14.652 109.636 14.724 118.676 ; 
      RECT 14.58 121.044 14.652 121.376 ; 
      RECT 14.436 104.546 14.508 137.374 ; 
      RECT 14.292 119.954 14.364 122.714 ; 
      RECT 14.292 122.918 14.364 126.884 ; 
      RECT 14.292 127.004 14.364 130.14 ; 
      RECT 14.22 106.54 14.292 108.524 ; 
      RECT 14.22 111.652 14.292 113.924 ; 
      RECT 14.22 115.18 14.292 118.1 ; 
      RECT 14.148 119.7 14.22 122.5188 ; 
      RECT 14.148 125.488 14.22 130.212 ; 
      RECT 14.004 104.546 14.076 105.946 ; 
      RECT 13.572 104.546 13.644 105.946 ; 
      RECT 13.14 104.546 13.212 105.946 ; 
      RECT 12.708 104.546 12.78 105.946 ; 
      RECT 12.276 104.546 12.348 105.946 ; 
      RECT 11.844 104.546 11.916 105.946 ; 
      RECT 11.412 104.546 11.484 105.946 ; 
      RECT 10.98 104.546 11.052 105.946 ; 
      RECT 10.548 104.546 10.62 105.946 ; 
      RECT 10.116 104.546 10.188 105.946 ; 
      RECT 9.684 104.546 9.756 105.946 ; 
      RECT 9.252 104.546 9.324 105.946 ; 
      RECT 8.82 104.546 8.892 105.946 ; 
      RECT 8.388 104.546 8.46 105.946 ; 
      RECT 7.956 104.546 8.028 105.946 ; 
      RECT 7.524 104.546 7.596 105.946 ; 
      RECT 7.092 104.546 7.164 105.946 ; 
      RECT 6.66 104.546 6.732 105.946 ; 
      RECT 6.228 104.546 6.3 105.946 ; 
      RECT 5.796 104.546 5.868 105.946 ; 
      RECT 5.364 104.546 5.436 105.946 ; 
      RECT 4.932 104.546 5.004 105.946 ; 
      RECT 4.5 104.546 4.572 105.946 ; 
      RECT 4.068 104.546 4.14 105.946 ; 
      RECT 3.636 104.546 3.708 105.946 ; 
      RECT 3.204 104.546 3.276 105.946 ; 
      RECT 2.772 104.546 2.844 105.946 ; 
      RECT 2.34 104.546 2.412 105.946 ; 
      RECT 1.908 104.546 1.98 105.946 ; 
      RECT 1.476 104.546 1.548 105.946 ; 
      RECT 1.332 119.966 1.404 122.534 ; 
      RECT 1.332 125.244 1.404 127.372 ; 
      RECT 1.26 108.7 1.332 109.604 ; 
      RECT 1.188 119.624 1.26 122.714 ; 
      RECT 1.188 122.9188 1.26 124.884 ; 
      RECT 1.188 125.084 1.26 126.57 ; 
      RECT 1.188 126.822 1.26 130.068 ; 
      RECT 1.044 104.546 1.116 137.374 ; 
      RECT 0.9 114.564 0.972 114.84 ; 
      RECT 0.9 121.796 0.972 123.654 ; 
      RECT 0.756 119.824 0.828 137.246 ; 
        RECT 20.952 137.568 21.024 141.31 ; 
        RECT 20.808 137.568 20.88 141.31 ; 
        RECT 20.664 139.876 20.736 141.166 ; 
        RECT 20.196 140.664 20.268 141.102 ; 
        RECT 20.16 137.698 20.232 138.656 ; 
        RECT 20.016 140.022 20.088 140.636 ; 
        RECT 19.692 140.124 19.764 141.156 ; 
        RECT 17.532 137.568 17.604 141.31 ; 
        RECT 17.388 137.568 17.46 141.31 ; 
        RECT 17.244 138.292 17.316 140.564 ; 
        RECT 20.952 141.888 21.024 145.63 ; 
        RECT 20.808 141.888 20.88 145.63 ; 
        RECT 20.664 144.196 20.736 145.486 ; 
        RECT 20.196 144.984 20.268 145.422 ; 
        RECT 20.16 142.018 20.232 142.976 ; 
        RECT 20.016 144.342 20.088 144.956 ; 
        RECT 19.692 144.444 19.764 145.476 ; 
        RECT 17.532 141.888 17.604 145.63 ; 
        RECT 17.388 141.888 17.46 145.63 ; 
        RECT 17.244 142.612 17.316 144.884 ; 
        RECT 20.952 146.208 21.024 149.95 ; 
        RECT 20.808 146.208 20.88 149.95 ; 
        RECT 20.664 148.516 20.736 149.806 ; 
        RECT 20.196 149.304 20.268 149.742 ; 
        RECT 20.16 146.338 20.232 147.296 ; 
        RECT 20.016 148.662 20.088 149.276 ; 
        RECT 19.692 148.764 19.764 149.796 ; 
        RECT 17.532 146.208 17.604 149.95 ; 
        RECT 17.388 146.208 17.46 149.95 ; 
        RECT 17.244 146.932 17.316 149.204 ; 
        RECT 20.952 150.528 21.024 154.27 ; 
        RECT 20.808 150.528 20.88 154.27 ; 
        RECT 20.664 152.836 20.736 154.126 ; 
        RECT 20.196 153.624 20.268 154.062 ; 
        RECT 20.16 150.658 20.232 151.616 ; 
        RECT 20.016 152.982 20.088 153.596 ; 
        RECT 19.692 153.084 19.764 154.116 ; 
        RECT 17.532 150.528 17.604 154.27 ; 
        RECT 17.388 150.528 17.46 154.27 ; 
        RECT 17.244 151.252 17.316 153.524 ; 
        RECT 20.952 154.848 21.024 158.59 ; 
        RECT 20.808 154.848 20.88 158.59 ; 
        RECT 20.664 157.156 20.736 158.446 ; 
        RECT 20.196 157.944 20.268 158.382 ; 
        RECT 20.16 154.978 20.232 155.936 ; 
        RECT 20.016 157.302 20.088 157.916 ; 
        RECT 19.692 157.404 19.764 158.436 ; 
        RECT 17.532 154.848 17.604 158.59 ; 
        RECT 17.388 154.848 17.46 158.59 ; 
        RECT 17.244 155.572 17.316 157.844 ; 
        RECT 20.952 159.168 21.024 162.91 ; 
        RECT 20.808 159.168 20.88 162.91 ; 
        RECT 20.664 161.476 20.736 162.766 ; 
        RECT 20.196 162.264 20.268 162.702 ; 
        RECT 20.16 159.298 20.232 160.256 ; 
        RECT 20.016 161.622 20.088 162.236 ; 
        RECT 19.692 161.724 19.764 162.756 ; 
        RECT 17.532 159.168 17.604 162.91 ; 
        RECT 17.388 159.168 17.46 162.91 ; 
        RECT 17.244 159.892 17.316 162.164 ; 
        RECT 20.952 163.488 21.024 167.23 ; 
        RECT 20.808 163.488 20.88 167.23 ; 
        RECT 20.664 165.796 20.736 167.086 ; 
        RECT 20.196 166.584 20.268 167.022 ; 
        RECT 20.16 163.618 20.232 164.576 ; 
        RECT 20.016 165.942 20.088 166.556 ; 
        RECT 19.692 166.044 19.764 167.076 ; 
        RECT 17.532 163.488 17.604 167.23 ; 
        RECT 17.388 163.488 17.46 167.23 ; 
        RECT 17.244 164.212 17.316 166.484 ; 
        RECT 20.952 167.808 21.024 171.55 ; 
        RECT 20.808 167.808 20.88 171.55 ; 
        RECT 20.664 170.116 20.736 171.406 ; 
        RECT 20.196 170.904 20.268 171.342 ; 
        RECT 20.16 167.938 20.232 168.896 ; 
        RECT 20.016 170.262 20.088 170.876 ; 
        RECT 19.692 170.364 19.764 171.396 ; 
        RECT 17.532 167.808 17.604 171.55 ; 
        RECT 17.388 167.808 17.46 171.55 ; 
        RECT 17.244 168.532 17.316 170.804 ; 
        RECT 20.952 172.128 21.024 175.87 ; 
        RECT 20.808 172.128 20.88 175.87 ; 
        RECT 20.664 174.436 20.736 175.726 ; 
        RECT 20.196 175.224 20.268 175.662 ; 
        RECT 20.16 172.258 20.232 173.216 ; 
        RECT 20.016 174.582 20.088 175.196 ; 
        RECT 19.692 174.684 19.764 175.716 ; 
        RECT 17.532 172.128 17.604 175.87 ; 
        RECT 17.388 172.128 17.46 175.87 ; 
        RECT 17.244 172.852 17.316 175.124 ; 
        RECT 20.952 176.448 21.024 180.19 ; 
        RECT 20.808 176.448 20.88 180.19 ; 
        RECT 20.664 178.756 20.736 180.046 ; 
        RECT 20.196 179.544 20.268 179.982 ; 
        RECT 20.16 176.578 20.232 177.536 ; 
        RECT 20.016 178.902 20.088 179.516 ; 
        RECT 19.692 179.004 19.764 180.036 ; 
        RECT 17.532 176.448 17.604 180.19 ; 
        RECT 17.388 176.448 17.46 180.19 ; 
        RECT 17.244 177.172 17.316 179.444 ; 
        RECT 20.952 180.768 21.024 184.51 ; 
        RECT 20.808 180.768 20.88 184.51 ; 
        RECT 20.664 183.076 20.736 184.366 ; 
        RECT 20.196 183.864 20.268 184.302 ; 
        RECT 20.16 180.898 20.232 181.856 ; 
        RECT 20.016 183.222 20.088 183.836 ; 
        RECT 19.692 183.324 19.764 184.356 ; 
        RECT 17.532 180.768 17.604 184.51 ; 
        RECT 17.388 180.768 17.46 184.51 ; 
        RECT 17.244 181.492 17.316 183.764 ; 
        RECT 20.952 185.088 21.024 188.83 ; 
        RECT 20.808 185.088 20.88 188.83 ; 
        RECT 20.664 187.396 20.736 188.686 ; 
        RECT 20.196 188.184 20.268 188.622 ; 
        RECT 20.16 185.218 20.232 186.176 ; 
        RECT 20.016 187.542 20.088 188.156 ; 
        RECT 19.692 187.644 19.764 188.676 ; 
        RECT 17.532 185.088 17.604 188.83 ; 
        RECT 17.388 185.088 17.46 188.83 ; 
        RECT 17.244 185.812 17.316 188.084 ; 
        RECT 20.952 189.408 21.024 193.15 ; 
        RECT 20.808 189.408 20.88 193.15 ; 
        RECT 20.664 191.716 20.736 193.006 ; 
        RECT 20.196 192.504 20.268 192.942 ; 
        RECT 20.16 189.538 20.232 190.496 ; 
        RECT 20.016 191.862 20.088 192.476 ; 
        RECT 19.692 191.964 19.764 192.996 ; 
        RECT 17.532 189.408 17.604 193.15 ; 
        RECT 17.388 189.408 17.46 193.15 ; 
        RECT 17.244 190.132 17.316 192.404 ; 
        RECT 20.952 193.728 21.024 197.47 ; 
        RECT 20.808 193.728 20.88 197.47 ; 
        RECT 20.664 196.036 20.736 197.326 ; 
        RECT 20.196 196.824 20.268 197.262 ; 
        RECT 20.16 193.858 20.232 194.816 ; 
        RECT 20.016 196.182 20.088 196.796 ; 
        RECT 19.692 196.284 19.764 197.316 ; 
        RECT 17.532 193.728 17.604 197.47 ; 
        RECT 17.388 193.728 17.46 197.47 ; 
        RECT 17.244 194.452 17.316 196.724 ; 
        RECT 20.952 198.048 21.024 201.79 ; 
        RECT 20.808 198.048 20.88 201.79 ; 
        RECT 20.664 200.356 20.736 201.646 ; 
        RECT 20.196 201.144 20.268 201.582 ; 
        RECT 20.16 198.178 20.232 199.136 ; 
        RECT 20.016 200.502 20.088 201.116 ; 
        RECT 19.692 200.604 19.764 201.636 ; 
        RECT 17.532 198.048 17.604 201.79 ; 
        RECT 17.388 198.048 17.46 201.79 ; 
        RECT 17.244 198.772 17.316 201.044 ; 
        RECT 20.952 202.368 21.024 206.11 ; 
        RECT 20.808 202.368 20.88 206.11 ; 
        RECT 20.664 204.676 20.736 205.966 ; 
        RECT 20.196 205.464 20.268 205.902 ; 
        RECT 20.16 202.498 20.232 203.456 ; 
        RECT 20.016 204.822 20.088 205.436 ; 
        RECT 19.692 204.924 19.764 205.956 ; 
        RECT 17.532 202.368 17.604 206.11 ; 
        RECT 17.388 202.368 17.46 206.11 ; 
        RECT 17.244 203.092 17.316 205.364 ; 
        RECT 20.952 206.688 21.024 210.43 ; 
        RECT 20.808 206.688 20.88 210.43 ; 
        RECT 20.664 208.996 20.736 210.286 ; 
        RECT 20.196 209.784 20.268 210.222 ; 
        RECT 20.16 206.818 20.232 207.776 ; 
        RECT 20.016 209.142 20.088 209.756 ; 
        RECT 19.692 209.244 19.764 210.276 ; 
        RECT 17.532 206.688 17.604 210.43 ; 
        RECT 17.388 206.688 17.46 210.43 ; 
        RECT 17.244 207.412 17.316 209.684 ; 
        RECT 20.952 211.008 21.024 214.75 ; 
        RECT 20.808 211.008 20.88 214.75 ; 
        RECT 20.664 213.316 20.736 214.606 ; 
        RECT 20.196 214.104 20.268 214.542 ; 
        RECT 20.16 211.138 20.232 212.096 ; 
        RECT 20.016 213.462 20.088 214.076 ; 
        RECT 19.692 213.564 19.764 214.596 ; 
        RECT 17.532 211.008 17.604 214.75 ; 
        RECT 17.388 211.008 17.46 214.75 ; 
        RECT 17.244 211.732 17.316 214.004 ; 
        RECT 20.952 215.328 21.024 219.07 ; 
        RECT 20.808 215.328 20.88 219.07 ; 
        RECT 20.664 217.636 20.736 218.926 ; 
        RECT 20.196 218.424 20.268 218.862 ; 
        RECT 20.16 215.458 20.232 216.416 ; 
        RECT 20.016 217.782 20.088 218.396 ; 
        RECT 19.692 217.884 19.764 218.916 ; 
        RECT 17.532 215.328 17.604 219.07 ; 
        RECT 17.388 215.328 17.46 219.07 ; 
        RECT 17.244 216.052 17.316 218.324 ; 
        RECT 20.952 219.648 21.024 223.39 ; 
        RECT 20.808 219.648 20.88 223.39 ; 
        RECT 20.664 221.956 20.736 223.246 ; 
        RECT 20.196 222.744 20.268 223.182 ; 
        RECT 20.16 219.778 20.232 220.736 ; 
        RECT 20.016 222.102 20.088 222.716 ; 
        RECT 19.692 222.204 19.764 223.236 ; 
        RECT 17.532 219.648 17.604 223.39 ; 
        RECT 17.388 219.648 17.46 223.39 ; 
        RECT 17.244 220.372 17.316 222.644 ; 
        RECT 20.952 223.968 21.024 227.71 ; 
        RECT 20.808 223.968 20.88 227.71 ; 
        RECT 20.664 226.276 20.736 227.566 ; 
        RECT 20.196 227.064 20.268 227.502 ; 
        RECT 20.16 224.098 20.232 225.056 ; 
        RECT 20.016 226.422 20.088 227.036 ; 
        RECT 19.692 226.524 19.764 227.556 ; 
        RECT 17.532 223.968 17.604 227.71 ; 
        RECT 17.388 223.968 17.46 227.71 ; 
        RECT 17.244 224.692 17.316 226.964 ; 
        RECT 20.952 228.288 21.024 232.03 ; 
        RECT 20.808 228.288 20.88 232.03 ; 
        RECT 20.664 230.596 20.736 231.886 ; 
        RECT 20.196 231.384 20.268 231.822 ; 
        RECT 20.16 228.418 20.232 229.376 ; 
        RECT 20.016 230.742 20.088 231.356 ; 
        RECT 19.692 230.844 19.764 231.876 ; 
        RECT 17.532 228.288 17.604 232.03 ; 
        RECT 17.388 228.288 17.46 232.03 ; 
        RECT 17.244 229.012 17.316 231.284 ; 
        RECT 20.952 232.608 21.024 236.35 ; 
        RECT 20.808 232.608 20.88 236.35 ; 
        RECT 20.664 234.916 20.736 236.206 ; 
        RECT 20.196 235.704 20.268 236.142 ; 
        RECT 20.16 232.738 20.232 233.696 ; 
        RECT 20.016 235.062 20.088 235.676 ; 
        RECT 19.692 235.164 19.764 236.196 ; 
        RECT 17.532 232.608 17.604 236.35 ; 
        RECT 17.388 232.608 17.46 236.35 ; 
        RECT 17.244 233.332 17.316 235.604 ; 
        RECT 20.952 236.928 21.024 240.67 ; 
        RECT 20.808 236.928 20.88 240.67 ; 
        RECT 20.664 239.236 20.736 240.526 ; 
        RECT 20.196 240.024 20.268 240.462 ; 
        RECT 20.16 237.058 20.232 238.016 ; 
        RECT 20.016 239.382 20.088 239.996 ; 
        RECT 19.692 239.484 19.764 240.516 ; 
        RECT 17.532 236.928 17.604 240.67 ; 
        RECT 17.388 236.928 17.46 240.67 ; 
        RECT 17.244 237.652 17.316 239.924 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 20.72 1.026 21.232 5.4 ; 
      RECT 20.664 3.688 21.232 4.978 ; 
      RECT 20.072 2.596 20.32 5.4 ; 
      RECT 20.016 3.834 20.32 4.448 ; 
      RECT 20.072 1.026 20.176 5.4 ; 
      RECT 20.072 1.51 20.232 2.468 ; 
      RECT 20.072 1.026 20.32 1.382 ; 
      RECT 18.884 2.828 19.708 5.4 ; 
      RECT 19.604 1.026 19.708 5.4 ; 
      RECT 18.884 3.936 19.764 4.968 ; 
      RECT 18.884 1.026 19.276 5.4 ; 
      RECT 17.216 1.026 17.548 5.4 ; 
      RECT 17.216 1.38 17.604 5.122 ; 
      RECT 38.108 1.026 38.448 5.4 ; 
      RECT 37.532 1.026 37.636 5.4 ; 
      RECT 37.1 1.026 37.204 5.4 ; 
      RECT 36.668 1.026 36.772 5.4 ; 
      RECT 36.236 1.026 36.34 5.4 ; 
      RECT 35.804 1.026 35.908 5.4 ; 
      RECT 35.372 1.026 35.476 5.4 ; 
      RECT 34.94 1.026 35.044 5.4 ; 
      RECT 34.508 1.026 34.612 5.4 ; 
      RECT 34.076 1.026 34.18 5.4 ; 
      RECT 33.644 1.026 33.748 5.4 ; 
      RECT 33.212 1.026 33.316 5.4 ; 
      RECT 32.78 1.026 32.884 5.4 ; 
      RECT 32.348 1.026 32.452 5.4 ; 
      RECT 31.916 1.026 32.02 5.4 ; 
      RECT 31.484 1.026 31.588 5.4 ; 
      RECT 31.052 1.026 31.156 5.4 ; 
      RECT 30.62 1.026 30.724 5.4 ; 
      RECT 30.188 1.026 30.292 5.4 ; 
      RECT 29.756 1.026 29.86 5.4 ; 
      RECT 29.324 1.026 29.428 5.4 ; 
      RECT 28.892 1.026 28.996 5.4 ; 
      RECT 28.46 1.026 28.564 5.4 ; 
      RECT 28.028 1.026 28.132 5.4 ; 
      RECT 27.596 1.026 27.7 5.4 ; 
      RECT 27.164 1.026 27.268 5.4 ; 
      RECT 26.732 1.026 26.836 5.4 ; 
      RECT 26.3 1.026 26.404 5.4 ; 
      RECT 25.868 1.026 25.972 5.4 ; 
      RECT 25.436 1.026 25.54 5.4 ; 
      RECT 25.004 1.026 25.108 5.4 ; 
      RECT 24.572 1.026 24.676 5.4 ; 
      RECT 24.14 1.026 24.244 5.4 ; 
      RECT 23.708 1.026 23.812 5.4 ; 
      RECT 22.856 1.026 23.164 5.4 ; 
      RECT 15.284 1.026 15.592 5.4 ; 
      RECT 14.636 1.026 14.74 5.4 ; 
      RECT 14.204 1.026 14.308 5.4 ; 
      RECT 13.772 1.026 13.876 5.4 ; 
      RECT 13.34 1.026 13.444 5.4 ; 
      RECT 12.908 1.026 13.012 5.4 ; 
      RECT 12.476 1.026 12.58 5.4 ; 
      RECT 12.044 1.026 12.148 5.4 ; 
      RECT 11.612 1.026 11.716 5.4 ; 
      RECT 11.18 1.026 11.284 5.4 ; 
      RECT 10.748 1.026 10.852 5.4 ; 
      RECT 10.316 1.026 10.42 5.4 ; 
      RECT 9.884 1.026 9.988 5.4 ; 
      RECT 9.452 1.026 9.556 5.4 ; 
      RECT 9.02 1.026 9.124 5.4 ; 
      RECT 8.588 1.026 8.692 5.4 ; 
      RECT 8.156 1.026 8.26 5.4 ; 
      RECT 7.724 1.026 7.828 5.4 ; 
      RECT 7.292 1.026 7.396 5.4 ; 
      RECT 6.86 1.026 6.964 5.4 ; 
      RECT 6.428 1.026 6.532 5.4 ; 
      RECT 5.996 1.026 6.1 5.4 ; 
      RECT 5.564 1.026 5.668 5.4 ; 
      RECT 5.132 1.026 5.236 5.4 ; 
      RECT 4.7 1.026 4.804 5.4 ; 
      RECT 4.268 1.026 4.372 5.4 ; 
      RECT 3.836 1.026 3.94 5.4 ; 
      RECT 3.404 1.026 3.508 5.4 ; 
      RECT 2.972 1.026 3.076 5.4 ; 
      RECT 2.54 1.026 2.644 5.4 ; 
      RECT 2.108 1.026 2.212 5.4 ; 
      RECT 1.676 1.026 1.78 5.4 ; 
      RECT 1.244 1.026 1.348 5.4 ; 
      RECT 0.812 1.026 0.916 5.4 ; 
      RECT 0 1.026 0.34 5.4 ; 
      RECT 20.72 5.346 21.232 9.72 ; 
      RECT 20.664 8.008 21.232 9.298 ; 
      RECT 20.072 6.916 20.32 9.72 ; 
      RECT 20.016 8.154 20.32 8.768 ; 
      RECT 20.072 5.346 20.176 9.72 ; 
      RECT 20.072 5.83 20.232 6.788 ; 
      RECT 20.072 5.346 20.32 5.702 ; 
      RECT 18.884 7.148 19.708 9.72 ; 
      RECT 19.604 5.346 19.708 9.72 ; 
      RECT 18.884 8.256 19.764 9.288 ; 
      RECT 18.884 5.346 19.276 9.72 ; 
      RECT 17.216 5.346 17.548 9.72 ; 
      RECT 17.216 5.7 17.604 9.442 ; 
      RECT 38.108 5.346 38.448 9.72 ; 
      RECT 37.532 5.346 37.636 9.72 ; 
      RECT 37.1 5.346 37.204 9.72 ; 
      RECT 36.668 5.346 36.772 9.72 ; 
      RECT 36.236 5.346 36.34 9.72 ; 
      RECT 35.804 5.346 35.908 9.72 ; 
      RECT 35.372 5.346 35.476 9.72 ; 
      RECT 34.94 5.346 35.044 9.72 ; 
      RECT 34.508 5.346 34.612 9.72 ; 
      RECT 34.076 5.346 34.18 9.72 ; 
      RECT 33.644 5.346 33.748 9.72 ; 
      RECT 33.212 5.346 33.316 9.72 ; 
      RECT 32.78 5.346 32.884 9.72 ; 
      RECT 32.348 5.346 32.452 9.72 ; 
      RECT 31.916 5.346 32.02 9.72 ; 
      RECT 31.484 5.346 31.588 9.72 ; 
      RECT 31.052 5.346 31.156 9.72 ; 
      RECT 30.62 5.346 30.724 9.72 ; 
      RECT 30.188 5.346 30.292 9.72 ; 
      RECT 29.756 5.346 29.86 9.72 ; 
      RECT 29.324 5.346 29.428 9.72 ; 
      RECT 28.892 5.346 28.996 9.72 ; 
      RECT 28.46 5.346 28.564 9.72 ; 
      RECT 28.028 5.346 28.132 9.72 ; 
      RECT 27.596 5.346 27.7 9.72 ; 
      RECT 27.164 5.346 27.268 9.72 ; 
      RECT 26.732 5.346 26.836 9.72 ; 
      RECT 26.3 5.346 26.404 9.72 ; 
      RECT 25.868 5.346 25.972 9.72 ; 
      RECT 25.436 5.346 25.54 9.72 ; 
      RECT 25.004 5.346 25.108 9.72 ; 
      RECT 24.572 5.346 24.676 9.72 ; 
      RECT 24.14 5.346 24.244 9.72 ; 
      RECT 23.708 5.346 23.812 9.72 ; 
      RECT 22.856 5.346 23.164 9.72 ; 
      RECT 15.284 5.346 15.592 9.72 ; 
      RECT 14.636 5.346 14.74 9.72 ; 
      RECT 14.204 5.346 14.308 9.72 ; 
      RECT 13.772 5.346 13.876 9.72 ; 
      RECT 13.34 5.346 13.444 9.72 ; 
      RECT 12.908 5.346 13.012 9.72 ; 
      RECT 12.476 5.346 12.58 9.72 ; 
      RECT 12.044 5.346 12.148 9.72 ; 
      RECT 11.612 5.346 11.716 9.72 ; 
      RECT 11.18 5.346 11.284 9.72 ; 
      RECT 10.748 5.346 10.852 9.72 ; 
      RECT 10.316 5.346 10.42 9.72 ; 
      RECT 9.884 5.346 9.988 9.72 ; 
      RECT 9.452 5.346 9.556 9.72 ; 
      RECT 9.02 5.346 9.124 9.72 ; 
      RECT 8.588 5.346 8.692 9.72 ; 
      RECT 8.156 5.346 8.26 9.72 ; 
      RECT 7.724 5.346 7.828 9.72 ; 
      RECT 7.292 5.346 7.396 9.72 ; 
      RECT 6.86 5.346 6.964 9.72 ; 
      RECT 6.428 5.346 6.532 9.72 ; 
      RECT 5.996 5.346 6.1 9.72 ; 
      RECT 5.564 5.346 5.668 9.72 ; 
      RECT 5.132 5.346 5.236 9.72 ; 
      RECT 4.7 5.346 4.804 9.72 ; 
      RECT 4.268 5.346 4.372 9.72 ; 
      RECT 3.836 5.346 3.94 9.72 ; 
      RECT 3.404 5.346 3.508 9.72 ; 
      RECT 2.972 5.346 3.076 9.72 ; 
      RECT 2.54 5.346 2.644 9.72 ; 
      RECT 2.108 5.346 2.212 9.72 ; 
      RECT 1.676 5.346 1.78 9.72 ; 
      RECT 1.244 5.346 1.348 9.72 ; 
      RECT 0.812 5.346 0.916 9.72 ; 
      RECT 0 5.346 0.34 9.72 ; 
      RECT 20.72 9.666 21.232 14.04 ; 
      RECT 20.664 12.328 21.232 13.618 ; 
      RECT 20.072 11.236 20.32 14.04 ; 
      RECT 20.016 12.474 20.32 13.088 ; 
      RECT 20.072 9.666 20.176 14.04 ; 
      RECT 20.072 10.15 20.232 11.108 ; 
      RECT 20.072 9.666 20.32 10.022 ; 
      RECT 18.884 11.468 19.708 14.04 ; 
      RECT 19.604 9.666 19.708 14.04 ; 
      RECT 18.884 12.576 19.764 13.608 ; 
      RECT 18.884 9.666 19.276 14.04 ; 
      RECT 17.216 9.666 17.548 14.04 ; 
      RECT 17.216 10.02 17.604 13.762 ; 
      RECT 38.108 9.666 38.448 14.04 ; 
      RECT 37.532 9.666 37.636 14.04 ; 
      RECT 37.1 9.666 37.204 14.04 ; 
      RECT 36.668 9.666 36.772 14.04 ; 
      RECT 36.236 9.666 36.34 14.04 ; 
      RECT 35.804 9.666 35.908 14.04 ; 
      RECT 35.372 9.666 35.476 14.04 ; 
      RECT 34.94 9.666 35.044 14.04 ; 
      RECT 34.508 9.666 34.612 14.04 ; 
      RECT 34.076 9.666 34.18 14.04 ; 
      RECT 33.644 9.666 33.748 14.04 ; 
      RECT 33.212 9.666 33.316 14.04 ; 
      RECT 32.78 9.666 32.884 14.04 ; 
      RECT 32.348 9.666 32.452 14.04 ; 
      RECT 31.916 9.666 32.02 14.04 ; 
      RECT 31.484 9.666 31.588 14.04 ; 
      RECT 31.052 9.666 31.156 14.04 ; 
      RECT 30.62 9.666 30.724 14.04 ; 
      RECT 30.188 9.666 30.292 14.04 ; 
      RECT 29.756 9.666 29.86 14.04 ; 
      RECT 29.324 9.666 29.428 14.04 ; 
      RECT 28.892 9.666 28.996 14.04 ; 
      RECT 28.46 9.666 28.564 14.04 ; 
      RECT 28.028 9.666 28.132 14.04 ; 
      RECT 27.596 9.666 27.7 14.04 ; 
      RECT 27.164 9.666 27.268 14.04 ; 
      RECT 26.732 9.666 26.836 14.04 ; 
      RECT 26.3 9.666 26.404 14.04 ; 
      RECT 25.868 9.666 25.972 14.04 ; 
      RECT 25.436 9.666 25.54 14.04 ; 
      RECT 25.004 9.666 25.108 14.04 ; 
      RECT 24.572 9.666 24.676 14.04 ; 
      RECT 24.14 9.666 24.244 14.04 ; 
      RECT 23.708 9.666 23.812 14.04 ; 
      RECT 22.856 9.666 23.164 14.04 ; 
      RECT 15.284 9.666 15.592 14.04 ; 
      RECT 14.636 9.666 14.74 14.04 ; 
      RECT 14.204 9.666 14.308 14.04 ; 
      RECT 13.772 9.666 13.876 14.04 ; 
      RECT 13.34 9.666 13.444 14.04 ; 
      RECT 12.908 9.666 13.012 14.04 ; 
      RECT 12.476 9.666 12.58 14.04 ; 
      RECT 12.044 9.666 12.148 14.04 ; 
      RECT 11.612 9.666 11.716 14.04 ; 
      RECT 11.18 9.666 11.284 14.04 ; 
      RECT 10.748 9.666 10.852 14.04 ; 
      RECT 10.316 9.666 10.42 14.04 ; 
      RECT 9.884 9.666 9.988 14.04 ; 
      RECT 9.452 9.666 9.556 14.04 ; 
      RECT 9.02 9.666 9.124 14.04 ; 
      RECT 8.588 9.666 8.692 14.04 ; 
      RECT 8.156 9.666 8.26 14.04 ; 
      RECT 7.724 9.666 7.828 14.04 ; 
      RECT 7.292 9.666 7.396 14.04 ; 
      RECT 6.86 9.666 6.964 14.04 ; 
      RECT 6.428 9.666 6.532 14.04 ; 
      RECT 5.996 9.666 6.1 14.04 ; 
      RECT 5.564 9.666 5.668 14.04 ; 
      RECT 5.132 9.666 5.236 14.04 ; 
      RECT 4.7 9.666 4.804 14.04 ; 
      RECT 4.268 9.666 4.372 14.04 ; 
      RECT 3.836 9.666 3.94 14.04 ; 
      RECT 3.404 9.666 3.508 14.04 ; 
      RECT 2.972 9.666 3.076 14.04 ; 
      RECT 2.54 9.666 2.644 14.04 ; 
      RECT 2.108 9.666 2.212 14.04 ; 
      RECT 1.676 9.666 1.78 14.04 ; 
      RECT 1.244 9.666 1.348 14.04 ; 
      RECT 0.812 9.666 0.916 14.04 ; 
      RECT 0 9.666 0.34 14.04 ; 
      RECT 20.72 13.986 21.232 18.36 ; 
      RECT 20.664 16.648 21.232 17.938 ; 
      RECT 20.072 15.556 20.32 18.36 ; 
      RECT 20.016 16.794 20.32 17.408 ; 
      RECT 20.072 13.986 20.176 18.36 ; 
      RECT 20.072 14.47 20.232 15.428 ; 
      RECT 20.072 13.986 20.32 14.342 ; 
      RECT 18.884 15.788 19.708 18.36 ; 
      RECT 19.604 13.986 19.708 18.36 ; 
      RECT 18.884 16.896 19.764 17.928 ; 
      RECT 18.884 13.986 19.276 18.36 ; 
      RECT 17.216 13.986 17.548 18.36 ; 
      RECT 17.216 14.34 17.604 18.082 ; 
      RECT 38.108 13.986 38.448 18.36 ; 
      RECT 37.532 13.986 37.636 18.36 ; 
      RECT 37.1 13.986 37.204 18.36 ; 
      RECT 36.668 13.986 36.772 18.36 ; 
      RECT 36.236 13.986 36.34 18.36 ; 
      RECT 35.804 13.986 35.908 18.36 ; 
      RECT 35.372 13.986 35.476 18.36 ; 
      RECT 34.94 13.986 35.044 18.36 ; 
      RECT 34.508 13.986 34.612 18.36 ; 
      RECT 34.076 13.986 34.18 18.36 ; 
      RECT 33.644 13.986 33.748 18.36 ; 
      RECT 33.212 13.986 33.316 18.36 ; 
      RECT 32.78 13.986 32.884 18.36 ; 
      RECT 32.348 13.986 32.452 18.36 ; 
      RECT 31.916 13.986 32.02 18.36 ; 
      RECT 31.484 13.986 31.588 18.36 ; 
      RECT 31.052 13.986 31.156 18.36 ; 
      RECT 30.62 13.986 30.724 18.36 ; 
      RECT 30.188 13.986 30.292 18.36 ; 
      RECT 29.756 13.986 29.86 18.36 ; 
      RECT 29.324 13.986 29.428 18.36 ; 
      RECT 28.892 13.986 28.996 18.36 ; 
      RECT 28.46 13.986 28.564 18.36 ; 
      RECT 28.028 13.986 28.132 18.36 ; 
      RECT 27.596 13.986 27.7 18.36 ; 
      RECT 27.164 13.986 27.268 18.36 ; 
      RECT 26.732 13.986 26.836 18.36 ; 
      RECT 26.3 13.986 26.404 18.36 ; 
      RECT 25.868 13.986 25.972 18.36 ; 
      RECT 25.436 13.986 25.54 18.36 ; 
      RECT 25.004 13.986 25.108 18.36 ; 
      RECT 24.572 13.986 24.676 18.36 ; 
      RECT 24.14 13.986 24.244 18.36 ; 
      RECT 23.708 13.986 23.812 18.36 ; 
      RECT 22.856 13.986 23.164 18.36 ; 
      RECT 15.284 13.986 15.592 18.36 ; 
      RECT 14.636 13.986 14.74 18.36 ; 
      RECT 14.204 13.986 14.308 18.36 ; 
      RECT 13.772 13.986 13.876 18.36 ; 
      RECT 13.34 13.986 13.444 18.36 ; 
      RECT 12.908 13.986 13.012 18.36 ; 
      RECT 12.476 13.986 12.58 18.36 ; 
      RECT 12.044 13.986 12.148 18.36 ; 
      RECT 11.612 13.986 11.716 18.36 ; 
      RECT 11.18 13.986 11.284 18.36 ; 
      RECT 10.748 13.986 10.852 18.36 ; 
      RECT 10.316 13.986 10.42 18.36 ; 
      RECT 9.884 13.986 9.988 18.36 ; 
      RECT 9.452 13.986 9.556 18.36 ; 
      RECT 9.02 13.986 9.124 18.36 ; 
      RECT 8.588 13.986 8.692 18.36 ; 
      RECT 8.156 13.986 8.26 18.36 ; 
      RECT 7.724 13.986 7.828 18.36 ; 
      RECT 7.292 13.986 7.396 18.36 ; 
      RECT 6.86 13.986 6.964 18.36 ; 
      RECT 6.428 13.986 6.532 18.36 ; 
      RECT 5.996 13.986 6.1 18.36 ; 
      RECT 5.564 13.986 5.668 18.36 ; 
      RECT 5.132 13.986 5.236 18.36 ; 
      RECT 4.7 13.986 4.804 18.36 ; 
      RECT 4.268 13.986 4.372 18.36 ; 
      RECT 3.836 13.986 3.94 18.36 ; 
      RECT 3.404 13.986 3.508 18.36 ; 
      RECT 2.972 13.986 3.076 18.36 ; 
      RECT 2.54 13.986 2.644 18.36 ; 
      RECT 2.108 13.986 2.212 18.36 ; 
      RECT 1.676 13.986 1.78 18.36 ; 
      RECT 1.244 13.986 1.348 18.36 ; 
      RECT 0.812 13.986 0.916 18.36 ; 
      RECT 0 13.986 0.34 18.36 ; 
      RECT 20.72 18.306 21.232 22.68 ; 
      RECT 20.664 20.968 21.232 22.258 ; 
      RECT 20.072 19.876 20.32 22.68 ; 
      RECT 20.016 21.114 20.32 21.728 ; 
      RECT 20.072 18.306 20.176 22.68 ; 
      RECT 20.072 18.79 20.232 19.748 ; 
      RECT 20.072 18.306 20.32 18.662 ; 
      RECT 18.884 20.108 19.708 22.68 ; 
      RECT 19.604 18.306 19.708 22.68 ; 
      RECT 18.884 21.216 19.764 22.248 ; 
      RECT 18.884 18.306 19.276 22.68 ; 
      RECT 17.216 18.306 17.548 22.68 ; 
      RECT 17.216 18.66 17.604 22.402 ; 
      RECT 38.108 18.306 38.448 22.68 ; 
      RECT 37.532 18.306 37.636 22.68 ; 
      RECT 37.1 18.306 37.204 22.68 ; 
      RECT 36.668 18.306 36.772 22.68 ; 
      RECT 36.236 18.306 36.34 22.68 ; 
      RECT 35.804 18.306 35.908 22.68 ; 
      RECT 35.372 18.306 35.476 22.68 ; 
      RECT 34.94 18.306 35.044 22.68 ; 
      RECT 34.508 18.306 34.612 22.68 ; 
      RECT 34.076 18.306 34.18 22.68 ; 
      RECT 33.644 18.306 33.748 22.68 ; 
      RECT 33.212 18.306 33.316 22.68 ; 
      RECT 32.78 18.306 32.884 22.68 ; 
      RECT 32.348 18.306 32.452 22.68 ; 
      RECT 31.916 18.306 32.02 22.68 ; 
      RECT 31.484 18.306 31.588 22.68 ; 
      RECT 31.052 18.306 31.156 22.68 ; 
      RECT 30.62 18.306 30.724 22.68 ; 
      RECT 30.188 18.306 30.292 22.68 ; 
      RECT 29.756 18.306 29.86 22.68 ; 
      RECT 29.324 18.306 29.428 22.68 ; 
      RECT 28.892 18.306 28.996 22.68 ; 
      RECT 28.46 18.306 28.564 22.68 ; 
      RECT 28.028 18.306 28.132 22.68 ; 
      RECT 27.596 18.306 27.7 22.68 ; 
      RECT 27.164 18.306 27.268 22.68 ; 
      RECT 26.732 18.306 26.836 22.68 ; 
      RECT 26.3 18.306 26.404 22.68 ; 
      RECT 25.868 18.306 25.972 22.68 ; 
      RECT 25.436 18.306 25.54 22.68 ; 
      RECT 25.004 18.306 25.108 22.68 ; 
      RECT 24.572 18.306 24.676 22.68 ; 
      RECT 24.14 18.306 24.244 22.68 ; 
      RECT 23.708 18.306 23.812 22.68 ; 
      RECT 22.856 18.306 23.164 22.68 ; 
      RECT 15.284 18.306 15.592 22.68 ; 
      RECT 14.636 18.306 14.74 22.68 ; 
      RECT 14.204 18.306 14.308 22.68 ; 
      RECT 13.772 18.306 13.876 22.68 ; 
      RECT 13.34 18.306 13.444 22.68 ; 
      RECT 12.908 18.306 13.012 22.68 ; 
      RECT 12.476 18.306 12.58 22.68 ; 
      RECT 12.044 18.306 12.148 22.68 ; 
      RECT 11.612 18.306 11.716 22.68 ; 
      RECT 11.18 18.306 11.284 22.68 ; 
      RECT 10.748 18.306 10.852 22.68 ; 
      RECT 10.316 18.306 10.42 22.68 ; 
      RECT 9.884 18.306 9.988 22.68 ; 
      RECT 9.452 18.306 9.556 22.68 ; 
      RECT 9.02 18.306 9.124 22.68 ; 
      RECT 8.588 18.306 8.692 22.68 ; 
      RECT 8.156 18.306 8.26 22.68 ; 
      RECT 7.724 18.306 7.828 22.68 ; 
      RECT 7.292 18.306 7.396 22.68 ; 
      RECT 6.86 18.306 6.964 22.68 ; 
      RECT 6.428 18.306 6.532 22.68 ; 
      RECT 5.996 18.306 6.1 22.68 ; 
      RECT 5.564 18.306 5.668 22.68 ; 
      RECT 5.132 18.306 5.236 22.68 ; 
      RECT 4.7 18.306 4.804 22.68 ; 
      RECT 4.268 18.306 4.372 22.68 ; 
      RECT 3.836 18.306 3.94 22.68 ; 
      RECT 3.404 18.306 3.508 22.68 ; 
      RECT 2.972 18.306 3.076 22.68 ; 
      RECT 2.54 18.306 2.644 22.68 ; 
      RECT 2.108 18.306 2.212 22.68 ; 
      RECT 1.676 18.306 1.78 22.68 ; 
      RECT 1.244 18.306 1.348 22.68 ; 
      RECT 0.812 18.306 0.916 22.68 ; 
      RECT 0 18.306 0.34 22.68 ; 
      RECT 20.72 22.626 21.232 27 ; 
      RECT 20.664 25.288 21.232 26.578 ; 
      RECT 20.072 24.196 20.32 27 ; 
      RECT 20.016 25.434 20.32 26.048 ; 
      RECT 20.072 22.626 20.176 27 ; 
      RECT 20.072 23.11 20.232 24.068 ; 
      RECT 20.072 22.626 20.32 22.982 ; 
      RECT 18.884 24.428 19.708 27 ; 
      RECT 19.604 22.626 19.708 27 ; 
      RECT 18.884 25.536 19.764 26.568 ; 
      RECT 18.884 22.626 19.276 27 ; 
      RECT 17.216 22.626 17.548 27 ; 
      RECT 17.216 22.98 17.604 26.722 ; 
      RECT 38.108 22.626 38.448 27 ; 
      RECT 37.532 22.626 37.636 27 ; 
      RECT 37.1 22.626 37.204 27 ; 
      RECT 36.668 22.626 36.772 27 ; 
      RECT 36.236 22.626 36.34 27 ; 
      RECT 35.804 22.626 35.908 27 ; 
      RECT 35.372 22.626 35.476 27 ; 
      RECT 34.94 22.626 35.044 27 ; 
      RECT 34.508 22.626 34.612 27 ; 
      RECT 34.076 22.626 34.18 27 ; 
      RECT 33.644 22.626 33.748 27 ; 
      RECT 33.212 22.626 33.316 27 ; 
      RECT 32.78 22.626 32.884 27 ; 
      RECT 32.348 22.626 32.452 27 ; 
      RECT 31.916 22.626 32.02 27 ; 
      RECT 31.484 22.626 31.588 27 ; 
      RECT 31.052 22.626 31.156 27 ; 
      RECT 30.62 22.626 30.724 27 ; 
      RECT 30.188 22.626 30.292 27 ; 
      RECT 29.756 22.626 29.86 27 ; 
      RECT 29.324 22.626 29.428 27 ; 
      RECT 28.892 22.626 28.996 27 ; 
      RECT 28.46 22.626 28.564 27 ; 
      RECT 28.028 22.626 28.132 27 ; 
      RECT 27.596 22.626 27.7 27 ; 
      RECT 27.164 22.626 27.268 27 ; 
      RECT 26.732 22.626 26.836 27 ; 
      RECT 26.3 22.626 26.404 27 ; 
      RECT 25.868 22.626 25.972 27 ; 
      RECT 25.436 22.626 25.54 27 ; 
      RECT 25.004 22.626 25.108 27 ; 
      RECT 24.572 22.626 24.676 27 ; 
      RECT 24.14 22.626 24.244 27 ; 
      RECT 23.708 22.626 23.812 27 ; 
      RECT 22.856 22.626 23.164 27 ; 
      RECT 15.284 22.626 15.592 27 ; 
      RECT 14.636 22.626 14.74 27 ; 
      RECT 14.204 22.626 14.308 27 ; 
      RECT 13.772 22.626 13.876 27 ; 
      RECT 13.34 22.626 13.444 27 ; 
      RECT 12.908 22.626 13.012 27 ; 
      RECT 12.476 22.626 12.58 27 ; 
      RECT 12.044 22.626 12.148 27 ; 
      RECT 11.612 22.626 11.716 27 ; 
      RECT 11.18 22.626 11.284 27 ; 
      RECT 10.748 22.626 10.852 27 ; 
      RECT 10.316 22.626 10.42 27 ; 
      RECT 9.884 22.626 9.988 27 ; 
      RECT 9.452 22.626 9.556 27 ; 
      RECT 9.02 22.626 9.124 27 ; 
      RECT 8.588 22.626 8.692 27 ; 
      RECT 8.156 22.626 8.26 27 ; 
      RECT 7.724 22.626 7.828 27 ; 
      RECT 7.292 22.626 7.396 27 ; 
      RECT 6.86 22.626 6.964 27 ; 
      RECT 6.428 22.626 6.532 27 ; 
      RECT 5.996 22.626 6.1 27 ; 
      RECT 5.564 22.626 5.668 27 ; 
      RECT 5.132 22.626 5.236 27 ; 
      RECT 4.7 22.626 4.804 27 ; 
      RECT 4.268 22.626 4.372 27 ; 
      RECT 3.836 22.626 3.94 27 ; 
      RECT 3.404 22.626 3.508 27 ; 
      RECT 2.972 22.626 3.076 27 ; 
      RECT 2.54 22.626 2.644 27 ; 
      RECT 2.108 22.626 2.212 27 ; 
      RECT 1.676 22.626 1.78 27 ; 
      RECT 1.244 22.626 1.348 27 ; 
      RECT 0.812 22.626 0.916 27 ; 
      RECT 0 22.626 0.34 27 ; 
      RECT 20.72 26.946 21.232 31.32 ; 
      RECT 20.664 29.608 21.232 30.898 ; 
      RECT 20.072 28.516 20.32 31.32 ; 
      RECT 20.016 29.754 20.32 30.368 ; 
      RECT 20.072 26.946 20.176 31.32 ; 
      RECT 20.072 27.43 20.232 28.388 ; 
      RECT 20.072 26.946 20.32 27.302 ; 
      RECT 18.884 28.748 19.708 31.32 ; 
      RECT 19.604 26.946 19.708 31.32 ; 
      RECT 18.884 29.856 19.764 30.888 ; 
      RECT 18.884 26.946 19.276 31.32 ; 
      RECT 17.216 26.946 17.548 31.32 ; 
      RECT 17.216 27.3 17.604 31.042 ; 
      RECT 38.108 26.946 38.448 31.32 ; 
      RECT 37.532 26.946 37.636 31.32 ; 
      RECT 37.1 26.946 37.204 31.32 ; 
      RECT 36.668 26.946 36.772 31.32 ; 
      RECT 36.236 26.946 36.34 31.32 ; 
      RECT 35.804 26.946 35.908 31.32 ; 
      RECT 35.372 26.946 35.476 31.32 ; 
      RECT 34.94 26.946 35.044 31.32 ; 
      RECT 34.508 26.946 34.612 31.32 ; 
      RECT 34.076 26.946 34.18 31.32 ; 
      RECT 33.644 26.946 33.748 31.32 ; 
      RECT 33.212 26.946 33.316 31.32 ; 
      RECT 32.78 26.946 32.884 31.32 ; 
      RECT 32.348 26.946 32.452 31.32 ; 
      RECT 31.916 26.946 32.02 31.32 ; 
      RECT 31.484 26.946 31.588 31.32 ; 
      RECT 31.052 26.946 31.156 31.32 ; 
      RECT 30.62 26.946 30.724 31.32 ; 
      RECT 30.188 26.946 30.292 31.32 ; 
      RECT 29.756 26.946 29.86 31.32 ; 
      RECT 29.324 26.946 29.428 31.32 ; 
      RECT 28.892 26.946 28.996 31.32 ; 
      RECT 28.46 26.946 28.564 31.32 ; 
      RECT 28.028 26.946 28.132 31.32 ; 
      RECT 27.596 26.946 27.7 31.32 ; 
      RECT 27.164 26.946 27.268 31.32 ; 
      RECT 26.732 26.946 26.836 31.32 ; 
      RECT 26.3 26.946 26.404 31.32 ; 
      RECT 25.868 26.946 25.972 31.32 ; 
      RECT 25.436 26.946 25.54 31.32 ; 
      RECT 25.004 26.946 25.108 31.32 ; 
      RECT 24.572 26.946 24.676 31.32 ; 
      RECT 24.14 26.946 24.244 31.32 ; 
      RECT 23.708 26.946 23.812 31.32 ; 
      RECT 22.856 26.946 23.164 31.32 ; 
      RECT 15.284 26.946 15.592 31.32 ; 
      RECT 14.636 26.946 14.74 31.32 ; 
      RECT 14.204 26.946 14.308 31.32 ; 
      RECT 13.772 26.946 13.876 31.32 ; 
      RECT 13.34 26.946 13.444 31.32 ; 
      RECT 12.908 26.946 13.012 31.32 ; 
      RECT 12.476 26.946 12.58 31.32 ; 
      RECT 12.044 26.946 12.148 31.32 ; 
      RECT 11.612 26.946 11.716 31.32 ; 
      RECT 11.18 26.946 11.284 31.32 ; 
      RECT 10.748 26.946 10.852 31.32 ; 
      RECT 10.316 26.946 10.42 31.32 ; 
      RECT 9.884 26.946 9.988 31.32 ; 
      RECT 9.452 26.946 9.556 31.32 ; 
      RECT 9.02 26.946 9.124 31.32 ; 
      RECT 8.588 26.946 8.692 31.32 ; 
      RECT 8.156 26.946 8.26 31.32 ; 
      RECT 7.724 26.946 7.828 31.32 ; 
      RECT 7.292 26.946 7.396 31.32 ; 
      RECT 6.86 26.946 6.964 31.32 ; 
      RECT 6.428 26.946 6.532 31.32 ; 
      RECT 5.996 26.946 6.1 31.32 ; 
      RECT 5.564 26.946 5.668 31.32 ; 
      RECT 5.132 26.946 5.236 31.32 ; 
      RECT 4.7 26.946 4.804 31.32 ; 
      RECT 4.268 26.946 4.372 31.32 ; 
      RECT 3.836 26.946 3.94 31.32 ; 
      RECT 3.404 26.946 3.508 31.32 ; 
      RECT 2.972 26.946 3.076 31.32 ; 
      RECT 2.54 26.946 2.644 31.32 ; 
      RECT 2.108 26.946 2.212 31.32 ; 
      RECT 1.676 26.946 1.78 31.32 ; 
      RECT 1.244 26.946 1.348 31.32 ; 
      RECT 0.812 26.946 0.916 31.32 ; 
      RECT 0 26.946 0.34 31.32 ; 
      RECT 20.72 31.266 21.232 35.64 ; 
      RECT 20.664 33.928 21.232 35.218 ; 
      RECT 20.072 32.836 20.32 35.64 ; 
      RECT 20.016 34.074 20.32 34.688 ; 
      RECT 20.072 31.266 20.176 35.64 ; 
      RECT 20.072 31.75 20.232 32.708 ; 
      RECT 20.072 31.266 20.32 31.622 ; 
      RECT 18.884 33.068 19.708 35.64 ; 
      RECT 19.604 31.266 19.708 35.64 ; 
      RECT 18.884 34.176 19.764 35.208 ; 
      RECT 18.884 31.266 19.276 35.64 ; 
      RECT 17.216 31.266 17.548 35.64 ; 
      RECT 17.216 31.62 17.604 35.362 ; 
      RECT 38.108 31.266 38.448 35.64 ; 
      RECT 37.532 31.266 37.636 35.64 ; 
      RECT 37.1 31.266 37.204 35.64 ; 
      RECT 36.668 31.266 36.772 35.64 ; 
      RECT 36.236 31.266 36.34 35.64 ; 
      RECT 35.804 31.266 35.908 35.64 ; 
      RECT 35.372 31.266 35.476 35.64 ; 
      RECT 34.94 31.266 35.044 35.64 ; 
      RECT 34.508 31.266 34.612 35.64 ; 
      RECT 34.076 31.266 34.18 35.64 ; 
      RECT 33.644 31.266 33.748 35.64 ; 
      RECT 33.212 31.266 33.316 35.64 ; 
      RECT 32.78 31.266 32.884 35.64 ; 
      RECT 32.348 31.266 32.452 35.64 ; 
      RECT 31.916 31.266 32.02 35.64 ; 
      RECT 31.484 31.266 31.588 35.64 ; 
      RECT 31.052 31.266 31.156 35.64 ; 
      RECT 30.62 31.266 30.724 35.64 ; 
      RECT 30.188 31.266 30.292 35.64 ; 
      RECT 29.756 31.266 29.86 35.64 ; 
      RECT 29.324 31.266 29.428 35.64 ; 
      RECT 28.892 31.266 28.996 35.64 ; 
      RECT 28.46 31.266 28.564 35.64 ; 
      RECT 28.028 31.266 28.132 35.64 ; 
      RECT 27.596 31.266 27.7 35.64 ; 
      RECT 27.164 31.266 27.268 35.64 ; 
      RECT 26.732 31.266 26.836 35.64 ; 
      RECT 26.3 31.266 26.404 35.64 ; 
      RECT 25.868 31.266 25.972 35.64 ; 
      RECT 25.436 31.266 25.54 35.64 ; 
      RECT 25.004 31.266 25.108 35.64 ; 
      RECT 24.572 31.266 24.676 35.64 ; 
      RECT 24.14 31.266 24.244 35.64 ; 
      RECT 23.708 31.266 23.812 35.64 ; 
      RECT 22.856 31.266 23.164 35.64 ; 
      RECT 15.284 31.266 15.592 35.64 ; 
      RECT 14.636 31.266 14.74 35.64 ; 
      RECT 14.204 31.266 14.308 35.64 ; 
      RECT 13.772 31.266 13.876 35.64 ; 
      RECT 13.34 31.266 13.444 35.64 ; 
      RECT 12.908 31.266 13.012 35.64 ; 
      RECT 12.476 31.266 12.58 35.64 ; 
      RECT 12.044 31.266 12.148 35.64 ; 
      RECT 11.612 31.266 11.716 35.64 ; 
      RECT 11.18 31.266 11.284 35.64 ; 
      RECT 10.748 31.266 10.852 35.64 ; 
      RECT 10.316 31.266 10.42 35.64 ; 
      RECT 9.884 31.266 9.988 35.64 ; 
      RECT 9.452 31.266 9.556 35.64 ; 
      RECT 9.02 31.266 9.124 35.64 ; 
      RECT 8.588 31.266 8.692 35.64 ; 
      RECT 8.156 31.266 8.26 35.64 ; 
      RECT 7.724 31.266 7.828 35.64 ; 
      RECT 7.292 31.266 7.396 35.64 ; 
      RECT 6.86 31.266 6.964 35.64 ; 
      RECT 6.428 31.266 6.532 35.64 ; 
      RECT 5.996 31.266 6.1 35.64 ; 
      RECT 5.564 31.266 5.668 35.64 ; 
      RECT 5.132 31.266 5.236 35.64 ; 
      RECT 4.7 31.266 4.804 35.64 ; 
      RECT 4.268 31.266 4.372 35.64 ; 
      RECT 3.836 31.266 3.94 35.64 ; 
      RECT 3.404 31.266 3.508 35.64 ; 
      RECT 2.972 31.266 3.076 35.64 ; 
      RECT 2.54 31.266 2.644 35.64 ; 
      RECT 2.108 31.266 2.212 35.64 ; 
      RECT 1.676 31.266 1.78 35.64 ; 
      RECT 1.244 31.266 1.348 35.64 ; 
      RECT 0.812 31.266 0.916 35.64 ; 
      RECT 0 31.266 0.34 35.64 ; 
      RECT 20.72 35.586 21.232 39.96 ; 
      RECT 20.664 38.248 21.232 39.538 ; 
      RECT 20.072 37.156 20.32 39.96 ; 
      RECT 20.016 38.394 20.32 39.008 ; 
      RECT 20.072 35.586 20.176 39.96 ; 
      RECT 20.072 36.07 20.232 37.028 ; 
      RECT 20.072 35.586 20.32 35.942 ; 
      RECT 18.884 37.388 19.708 39.96 ; 
      RECT 19.604 35.586 19.708 39.96 ; 
      RECT 18.884 38.496 19.764 39.528 ; 
      RECT 18.884 35.586 19.276 39.96 ; 
      RECT 17.216 35.586 17.548 39.96 ; 
      RECT 17.216 35.94 17.604 39.682 ; 
      RECT 38.108 35.586 38.448 39.96 ; 
      RECT 37.532 35.586 37.636 39.96 ; 
      RECT 37.1 35.586 37.204 39.96 ; 
      RECT 36.668 35.586 36.772 39.96 ; 
      RECT 36.236 35.586 36.34 39.96 ; 
      RECT 35.804 35.586 35.908 39.96 ; 
      RECT 35.372 35.586 35.476 39.96 ; 
      RECT 34.94 35.586 35.044 39.96 ; 
      RECT 34.508 35.586 34.612 39.96 ; 
      RECT 34.076 35.586 34.18 39.96 ; 
      RECT 33.644 35.586 33.748 39.96 ; 
      RECT 33.212 35.586 33.316 39.96 ; 
      RECT 32.78 35.586 32.884 39.96 ; 
      RECT 32.348 35.586 32.452 39.96 ; 
      RECT 31.916 35.586 32.02 39.96 ; 
      RECT 31.484 35.586 31.588 39.96 ; 
      RECT 31.052 35.586 31.156 39.96 ; 
      RECT 30.62 35.586 30.724 39.96 ; 
      RECT 30.188 35.586 30.292 39.96 ; 
      RECT 29.756 35.586 29.86 39.96 ; 
      RECT 29.324 35.586 29.428 39.96 ; 
      RECT 28.892 35.586 28.996 39.96 ; 
      RECT 28.46 35.586 28.564 39.96 ; 
      RECT 28.028 35.586 28.132 39.96 ; 
      RECT 27.596 35.586 27.7 39.96 ; 
      RECT 27.164 35.586 27.268 39.96 ; 
      RECT 26.732 35.586 26.836 39.96 ; 
      RECT 26.3 35.586 26.404 39.96 ; 
      RECT 25.868 35.586 25.972 39.96 ; 
      RECT 25.436 35.586 25.54 39.96 ; 
      RECT 25.004 35.586 25.108 39.96 ; 
      RECT 24.572 35.586 24.676 39.96 ; 
      RECT 24.14 35.586 24.244 39.96 ; 
      RECT 23.708 35.586 23.812 39.96 ; 
      RECT 22.856 35.586 23.164 39.96 ; 
      RECT 15.284 35.586 15.592 39.96 ; 
      RECT 14.636 35.586 14.74 39.96 ; 
      RECT 14.204 35.586 14.308 39.96 ; 
      RECT 13.772 35.586 13.876 39.96 ; 
      RECT 13.34 35.586 13.444 39.96 ; 
      RECT 12.908 35.586 13.012 39.96 ; 
      RECT 12.476 35.586 12.58 39.96 ; 
      RECT 12.044 35.586 12.148 39.96 ; 
      RECT 11.612 35.586 11.716 39.96 ; 
      RECT 11.18 35.586 11.284 39.96 ; 
      RECT 10.748 35.586 10.852 39.96 ; 
      RECT 10.316 35.586 10.42 39.96 ; 
      RECT 9.884 35.586 9.988 39.96 ; 
      RECT 9.452 35.586 9.556 39.96 ; 
      RECT 9.02 35.586 9.124 39.96 ; 
      RECT 8.588 35.586 8.692 39.96 ; 
      RECT 8.156 35.586 8.26 39.96 ; 
      RECT 7.724 35.586 7.828 39.96 ; 
      RECT 7.292 35.586 7.396 39.96 ; 
      RECT 6.86 35.586 6.964 39.96 ; 
      RECT 6.428 35.586 6.532 39.96 ; 
      RECT 5.996 35.586 6.1 39.96 ; 
      RECT 5.564 35.586 5.668 39.96 ; 
      RECT 5.132 35.586 5.236 39.96 ; 
      RECT 4.7 35.586 4.804 39.96 ; 
      RECT 4.268 35.586 4.372 39.96 ; 
      RECT 3.836 35.586 3.94 39.96 ; 
      RECT 3.404 35.586 3.508 39.96 ; 
      RECT 2.972 35.586 3.076 39.96 ; 
      RECT 2.54 35.586 2.644 39.96 ; 
      RECT 2.108 35.586 2.212 39.96 ; 
      RECT 1.676 35.586 1.78 39.96 ; 
      RECT 1.244 35.586 1.348 39.96 ; 
      RECT 0.812 35.586 0.916 39.96 ; 
      RECT 0 35.586 0.34 39.96 ; 
      RECT 20.72 39.906 21.232 44.28 ; 
      RECT 20.664 42.568 21.232 43.858 ; 
      RECT 20.072 41.476 20.32 44.28 ; 
      RECT 20.016 42.714 20.32 43.328 ; 
      RECT 20.072 39.906 20.176 44.28 ; 
      RECT 20.072 40.39 20.232 41.348 ; 
      RECT 20.072 39.906 20.32 40.262 ; 
      RECT 18.884 41.708 19.708 44.28 ; 
      RECT 19.604 39.906 19.708 44.28 ; 
      RECT 18.884 42.816 19.764 43.848 ; 
      RECT 18.884 39.906 19.276 44.28 ; 
      RECT 17.216 39.906 17.548 44.28 ; 
      RECT 17.216 40.26 17.604 44.002 ; 
      RECT 38.108 39.906 38.448 44.28 ; 
      RECT 37.532 39.906 37.636 44.28 ; 
      RECT 37.1 39.906 37.204 44.28 ; 
      RECT 36.668 39.906 36.772 44.28 ; 
      RECT 36.236 39.906 36.34 44.28 ; 
      RECT 35.804 39.906 35.908 44.28 ; 
      RECT 35.372 39.906 35.476 44.28 ; 
      RECT 34.94 39.906 35.044 44.28 ; 
      RECT 34.508 39.906 34.612 44.28 ; 
      RECT 34.076 39.906 34.18 44.28 ; 
      RECT 33.644 39.906 33.748 44.28 ; 
      RECT 33.212 39.906 33.316 44.28 ; 
      RECT 32.78 39.906 32.884 44.28 ; 
      RECT 32.348 39.906 32.452 44.28 ; 
      RECT 31.916 39.906 32.02 44.28 ; 
      RECT 31.484 39.906 31.588 44.28 ; 
      RECT 31.052 39.906 31.156 44.28 ; 
      RECT 30.62 39.906 30.724 44.28 ; 
      RECT 30.188 39.906 30.292 44.28 ; 
      RECT 29.756 39.906 29.86 44.28 ; 
      RECT 29.324 39.906 29.428 44.28 ; 
      RECT 28.892 39.906 28.996 44.28 ; 
      RECT 28.46 39.906 28.564 44.28 ; 
      RECT 28.028 39.906 28.132 44.28 ; 
      RECT 27.596 39.906 27.7 44.28 ; 
      RECT 27.164 39.906 27.268 44.28 ; 
      RECT 26.732 39.906 26.836 44.28 ; 
      RECT 26.3 39.906 26.404 44.28 ; 
      RECT 25.868 39.906 25.972 44.28 ; 
      RECT 25.436 39.906 25.54 44.28 ; 
      RECT 25.004 39.906 25.108 44.28 ; 
      RECT 24.572 39.906 24.676 44.28 ; 
      RECT 24.14 39.906 24.244 44.28 ; 
      RECT 23.708 39.906 23.812 44.28 ; 
      RECT 22.856 39.906 23.164 44.28 ; 
      RECT 15.284 39.906 15.592 44.28 ; 
      RECT 14.636 39.906 14.74 44.28 ; 
      RECT 14.204 39.906 14.308 44.28 ; 
      RECT 13.772 39.906 13.876 44.28 ; 
      RECT 13.34 39.906 13.444 44.28 ; 
      RECT 12.908 39.906 13.012 44.28 ; 
      RECT 12.476 39.906 12.58 44.28 ; 
      RECT 12.044 39.906 12.148 44.28 ; 
      RECT 11.612 39.906 11.716 44.28 ; 
      RECT 11.18 39.906 11.284 44.28 ; 
      RECT 10.748 39.906 10.852 44.28 ; 
      RECT 10.316 39.906 10.42 44.28 ; 
      RECT 9.884 39.906 9.988 44.28 ; 
      RECT 9.452 39.906 9.556 44.28 ; 
      RECT 9.02 39.906 9.124 44.28 ; 
      RECT 8.588 39.906 8.692 44.28 ; 
      RECT 8.156 39.906 8.26 44.28 ; 
      RECT 7.724 39.906 7.828 44.28 ; 
      RECT 7.292 39.906 7.396 44.28 ; 
      RECT 6.86 39.906 6.964 44.28 ; 
      RECT 6.428 39.906 6.532 44.28 ; 
      RECT 5.996 39.906 6.1 44.28 ; 
      RECT 5.564 39.906 5.668 44.28 ; 
      RECT 5.132 39.906 5.236 44.28 ; 
      RECT 4.7 39.906 4.804 44.28 ; 
      RECT 4.268 39.906 4.372 44.28 ; 
      RECT 3.836 39.906 3.94 44.28 ; 
      RECT 3.404 39.906 3.508 44.28 ; 
      RECT 2.972 39.906 3.076 44.28 ; 
      RECT 2.54 39.906 2.644 44.28 ; 
      RECT 2.108 39.906 2.212 44.28 ; 
      RECT 1.676 39.906 1.78 44.28 ; 
      RECT 1.244 39.906 1.348 44.28 ; 
      RECT 0.812 39.906 0.916 44.28 ; 
      RECT 0 39.906 0.34 44.28 ; 
      RECT 20.72 44.226 21.232 48.6 ; 
      RECT 20.664 46.888 21.232 48.178 ; 
      RECT 20.072 45.796 20.32 48.6 ; 
      RECT 20.016 47.034 20.32 47.648 ; 
      RECT 20.072 44.226 20.176 48.6 ; 
      RECT 20.072 44.71 20.232 45.668 ; 
      RECT 20.072 44.226 20.32 44.582 ; 
      RECT 18.884 46.028 19.708 48.6 ; 
      RECT 19.604 44.226 19.708 48.6 ; 
      RECT 18.884 47.136 19.764 48.168 ; 
      RECT 18.884 44.226 19.276 48.6 ; 
      RECT 17.216 44.226 17.548 48.6 ; 
      RECT 17.216 44.58 17.604 48.322 ; 
      RECT 38.108 44.226 38.448 48.6 ; 
      RECT 37.532 44.226 37.636 48.6 ; 
      RECT 37.1 44.226 37.204 48.6 ; 
      RECT 36.668 44.226 36.772 48.6 ; 
      RECT 36.236 44.226 36.34 48.6 ; 
      RECT 35.804 44.226 35.908 48.6 ; 
      RECT 35.372 44.226 35.476 48.6 ; 
      RECT 34.94 44.226 35.044 48.6 ; 
      RECT 34.508 44.226 34.612 48.6 ; 
      RECT 34.076 44.226 34.18 48.6 ; 
      RECT 33.644 44.226 33.748 48.6 ; 
      RECT 33.212 44.226 33.316 48.6 ; 
      RECT 32.78 44.226 32.884 48.6 ; 
      RECT 32.348 44.226 32.452 48.6 ; 
      RECT 31.916 44.226 32.02 48.6 ; 
      RECT 31.484 44.226 31.588 48.6 ; 
      RECT 31.052 44.226 31.156 48.6 ; 
      RECT 30.62 44.226 30.724 48.6 ; 
      RECT 30.188 44.226 30.292 48.6 ; 
      RECT 29.756 44.226 29.86 48.6 ; 
      RECT 29.324 44.226 29.428 48.6 ; 
      RECT 28.892 44.226 28.996 48.6 ; 
      RECT 28.46 44.226 28.564 48.6 ; 
      RECT 28.028 44.226 28.132 48.6 ; 
      RECT 27.596 44.226 27.7 48.6 ; 
      RECT 27.164 44.226 27.268 48.6 ; 
      RECT 26.732 44.226 26.836 48.6 ; 
      RECT 26.3 44.226 26.404 48.6 ; 
      RECT 25.868 44.226 25.972 48.6 ; 
      RECT 25.436 44.226 25.54 48.6 ; 
      RECT 25.004 44.226 25.108 48.6 ; 
      RECT 24.572 44.226 24.676 48.6 ; 
      RECT 24.14 44.226 24.244 48.6 ; 
      RECT 23.708 44.226 23.812 48.6 ; 
      RECT 22.856 44.226 23.164 48.6 ; 
      RECT 15.284 44.226 15.592 48.6 ; 
      RECT 14.636 44.226 14.74 48.6 ; 
      RECT 14.204 44.226 14.308 48.6 ; 
      RECT 13.772 44.226 13.876 48.6 ; 
      RECT 13.34 44.226 13.444 48.6 ; 
      RECT 12.908 44.226 13.012 48.6 ; 
      RECT 12.476 44.226 12.58 48.6 ; 
      RECT 12.044 44.226 12.148 48.6 ; 
      RECT 11.612 44.226 11.716 48.6 ; 
      RECT 11.18 44.226 11.284 48.6 ; 
      RECT 10.748 44.226 10.852 48.6 ; 
      RECT 10.316 44.226 10.42 48.6 ; 
      RECT 9.884 44.226 9.988 48.6 ; 
      RECT 9.452 44.226 9.556 48.6 ; 
      RECT 9.02 44.226 9.124 48.6 ; 
      RECT 8.588 44.226 8.692 48.6 ; 
      RECT 8.156 44.226 8.26 48.6 ; 
      RECT 7.724 44.226 7.828 48.6 ; 
      RECT 7.292 44.226 7.396 48.6 ; 
      RECT 6.86 44.226 6.964 48.6 ; 
      RECT 6.428 44.226 6.532 48.6 ; 
      RECT 5.996 44.226 6.1 48.6 ; 
      RECT 5.564 44.226 5.668 48.6 ; 
      RECT 5.132 44.226 5.236 48.6 ; 
      RECT 4.7 44.226 4.804 48.6 ; 
      RECT 4.268 44.226 4.372 48.6 ; 
      RECT 3.836 44.226 3.94 48.6 ; 
      RECT 3.404 44.226 3.508 48.6 ; 
      RECT 2.972 44.226 3.076 48.6 ; 
      RECT 2.54 44.226 2.644 48.6 ; 
      RECT 2.108 44.226 2.212 48.6 ; 
      RECT 1.676 44.226 1.78 48.6 ; 
      RECT 1.244 44.226 1.348 48.6 ; 
      RECT 0.812 44.226 0.916 48.6 ; 
      RECT 0 44.226 0.34 48.6 ; 
      RECT 20.72 48.546 21.232 52.92 ; 
      RECT 20.664 51.208 21.232 52.498 ; 
      RECT 20.072 50.116 20.32 52.92 ; 
      RECT 20.016 51.354 20.32 51.968 ; 
      RECT 20.072 48.546 20.176 52.92 ; 
      RECT 20.072 49.03 20.232 49.988 ; 
      RECT 20.072 48.546 20.32 48.902 ; 
      RECT 18.884 50.348 19.708 52.92 ; 
      RECT 19.604 48.546 19.708 52.92 ; 
      RECT 18.884 51.456 19.764 52.488 ; 
      RECT 18.884 48.546 19.276 52.92 ; 
      RECT 17.216 48.546 17.548 52.92 ; 
      RECT 17.216 48.9 17.604 52.642 ; 
      RECT 38.108 48.546 38.448 52.92 ; 
      RECT 37.532 48.546 37.636 52.92 ; 
      RECT 37.1 48.546 37.204 52.92 ; 
      RECT 36.668 48.546 36.772 52.92 ; 
      RECT 36.236 48.546 36.34 52.92 ; 
      RECT 35.804 48.546 35.908 52.92 ; 
      RECT 35.372 48.546 35.476 52.92 ; 
      RECT 34.94 48.546 35.044 52.92 ; 
      RECT 34.508 48.546 34.612 52.92 ; 
      RECT 34.076 48.546 34.18 52.92 ; 
      RECT 33.644 48.546 33.748 52.92 ; 
      RECT 33.212 48.546 33.316 52.92 ; 
      RECT 32.78 48.546 32.884 52.92 ; 
      RECT 32.348 48.546 32.452 52.92 ; 
      RECT 31.916 48.546 32.02 52.92 ; 
      RECT 31.484 48.546 31.588 52.92 ; 
      RECT 31.052 48.546 31.156 52.92 ; 
      RECT 30.62 48.546 30.724 52.92 ; 
      RECT 30.188 48.546 30.292 52.92 ; 
      RECT 29.756 48.546 29.86 52.92 ; 
      RECT 29.324 48.546 29.428 52.92 ; 
      RECT 28.892 48.546 28.996 52.92 ; 
      RECT 28.46 48.546 28.564 52.92 ; 
      RECT 28.028 48.546 28.132 52.92 ; 
      RECT 27.596 48.546 27.7 52.92 ; 
      RECT 27.164 48.546 27.268 52.92 ; 
      RECT 26.732 48.546 26.836 52.92 ; 
      RECT 26.3 48.546 26.404 52.92 ; 
      RECT 25.868 48.546 25.972 52.92 ; 
      RECT 25.436 48.546 25.54 52.92 ; 
      RECT 25.004 48.546 25.108 52.92 ; 
      RECT 24.572 48.546 24.676 52.92 ; 
      RECT 24.14 48.546 24.244 52.92 ; 
      RECT 23.708 48.546 23.812 52.92 ; 
      RECT 22.856 48.546 23.164 52.92 ; 
      RECT 15.284 48.546 15.592 52.92 ; 
      RECT 14.636 48.546 14.74 52.92 ; 
      RECT 14.204 48.546 14.308 52.92 ; 
      RECT 13.772 48.546 13.876 52.92 ; 
      RECT 13.34 48.546 13.444 52.92 ; 
      RECT 12.908 48.546 13.012 52.92 ; 
      RECT 12.476 48.546 12.58 52.92 ; 
      RECT 12.044 48.546 12.148 52.92 ; 
      RECT 11.612 48.546 11.716 52.92 ; 
      RECT 11.18 48.546 11.284 52.92 ; 
      RECT 10.748 48.546 10.852 52.92 ; 
      RECT 10.316 48.546 10.42 52.92 ; 
      RECT 9.884 48.546 9.988 52.92 ; 
      RECT 9.452 48.546 9.556 52.92 ; 
      RECT 9.02 48.546 9.124 52.92 ; 
      RECT 8.588 48.546 8.692 52.92 ; 
      RECT 8.156 48.546 8.26 52.92 ; 
      RECT 7.724 48.546 7.828 52.92 ; 
      RECT 7.292 48.546 7.396 52.92 ; 
      RECT 6.86 48.546 6.964 52.92 ; 
      RECT 6.428 48.546 6.532 52.92 ; 
      RECT 5.996 48.546 6.1 52.92 ; 
      RECT 5.564 48.546 5.668 52.92 ; 
      RECT 5.132 48.546 5.236 52.92 ; 
      RECT 4.7 48.546 4.804 52.92 ; 
      RECT 4.268 48.546 4.372 52.92 ; 
      RECT 3.836 48.546 3.94 52.92 ; 
      RECT 3.404 48.546 3.508 52.92 ; 
      RECT 2.972 48.546 3.076 52.92 ; 
      RECT 2.54 48.546 2.644 52.92 ; 
      RECT 2.108 48.546 2.212 52.92 ; 
      RECT 1.676 48.546 1.78 52.92 ; 
      RECT 1.244 48.546 1.348 52.92 ; 
      RECT 0.812 48.546 0.916 52.92 ; 
      RECT 0 48.546 0.34 52.92 ; 
      RECT 20.72 52.866 21.232 57.24 ; 
      RECT 20.664 55.528 21.232 56.818 ; 
      RECT 20.072 54.436 20.32 57.24 ; 
      RECT 20.016 55.674 20.32 56.288 ; 
      RECT 20.072 52.866 20.176 57.24 ; 
      RECT 20.072 53.35 20.232 54.308 ; 
      RECT 20.072 52.866 20.32 53.222 ; 
      RECT 18.884 54.668 19.708 57.24 ; 
      RECT 19.604 52.866 19.708 57.24 ; 
      RECT 18.884 55.776 19.764 56.808 ; 
      RECT 18.884 52.866 19.276 57.24 ; 
      RECT 17.216 52.866 17.548 57.24 ; 
      RECT 17.216 53.22 17.604 56.962 ; 
      RECT 38.108 52.866 38.448 57.24 ; 
      RECT 37.532 52.866 37.636 57.24 ; 
      RECT 37.1 52.866 37.204 57.24 ; 
      RECT 36.668 52.866 36.772 57.24 ; 
      RECT 36.236 52.866 36.34 57.24 ; 
      RECT 35.804 52.866 35.908 57.24 ; 
      RECT 35.372 52.866 35.476 57.24 ; 
      RECT 34.94 52.866 35.044 57.24 ; 
      RECT 34.508 52.866 34.612 57.24 ; 
      RECT 34.076 52.866 34.18 57.24 ; 
      RECT 33.644 52.866 33.748 57.24 ; 
      RECT 33.212 52.866 33.316 57.24 ; 
      RECT 32.78 52.866 32.884 57.24 ; 
      RECT 32.348 52.866 32.452 57.24 ; 
      RECT 31.916 52.866 32.02 57.24 ; 
      RECT 31.484 52.866 31.588 57.24 ; 
      RECT 31.052 52.866 31.156 57.24 ; 
      RECT 30.62 52.866 30.724 57.24 ; 
      RECT 30.188 52.866 30.292 57.24 ; 
      RECT 29.756 52.866 29.86 57.24 ; 
      RECT 29.324 52.866 29.428 57.24 ; 
      RECT 28.892 52.866 28.996 57.24 ; 
      RECT 28.46 52.866 28.564 57.24 ; 
      RECT 28.028 52.866 28.132 57.24 ; 
      RECT 27.596 52.866 27.7 57.24 ; 
      RECT 27.164 52.866 27.268 57.24 ; 
      RECT 26.732 52.866 26.836 57.24 ; 
      RECT 26.3 52.866 26.404 57.24 ; 
      RECT 25.868 52.866 25.972 57.24 ; 
      RECT 25.436 52.866 25.54 57.24 ; 
      RECT 25.004 52.866 25.108 57.24 ; 
      RECT 24.572 52.866 24.676 57.24 ; 
      RECT 24.14 52.866 24.244 57.24 ; 
      RECT 23.708 52.866 23.812 57.24 ; 
      RECT 22.856 52.866 23.164 57.24 ; 
      RECT 15.284 52.866 15.592 57.24 ; 
      RECT 14.636 52.866 14.74 57.24 ; 
      RECT 14.204 52.866 14.308 57.24 ; 
      RECT 13.772 52.866 13.876 57.24 ; 
      RECT 13.34 52.866 13.444 57.24 ; 
      RECT 12.908 52.866 13.012 57.24 ; 
      RECT 12.476 52.866 12.58 57.24 ; 
      RECT 12.044 52.866 12.148 57.24 ; 
      RECT 11.612 52.866 11.716 57.24 ; 
      RECT 11.18 52.866 11.284 57.24 ; 
      RECT 10.748 52.866 10.852 57.24 ; 
      RECT 10.316 52.866 10.42 57.24 ; 
      RECT 9.884 52.866 9.988 57.24 ; 
      RECT 9.452 52.866 9.556 57.24 ; 
      RECT 9.02 52.866 9.124 57.24 ; 
      RECT 8.588 52.866 8.692 57.24 ; 
      RECT 8.156 52.866 8.26 57.24 ; 
      RECT 7.724 52.866 7.828 57.24 ; 
      RECT 7.292 52.866 7.396 57.24 ; 
      RECT 6.86 52.866 6.964 57.24 ; 
      RECT 6.428 52.866 6.532 57.24 ; 
      RECT 5.996 52.866 6.1 57.24 ; 
      RECT 5.564 52.866 5.668 57.24 ; 
      RECT 5.132 52.866 5.236 57.24 ; 
      RECT 4.7 52.866 4.804 57.24 ; 
      RECT 4.268 52.866 4.372 57.24 ; 
      RECT 3.836 52.866 3.94 57.24 ; 
      RECT 3.404 52.866 3.508 57.24 ; 
      RECT 2.972 52.866 3.076 57.24 ; 
      RECT 2.54 52.866 2.644 57.24 ; 
      RECT 2.108 52.866 2.212 57.24 ; 
      RECT 1.676 52.866 1.78 57.24 ; 
      RECT 1.244 52.866 1.348 57.24 ; 
      RECT 0.812 52.866 0.916 57.24 ; 
      RECT 0 52.866 0.34 57.24 ; 
      RECT 20.72 57.186 21.232 61.56 ; 
      RECT 20.664 59.848 21.232 61.138 ; 
      RECT 20.072 58.756 20.32 61.56 ; 
      RECT 20.016 59.994 20.32 60.608 ; 
      RECT 20.072 57.186 20.176 61.56 ; 
      RECT 20.072 57.67 20.232 58.628 ; 
      RECT 20.072 57.186 20.32 57.542 ; 
      RECT 18.884 58.988 19.708 61.56 ; 
      RECT 19.604 57.186 19.708 61.56 ; 
      RECT 18.884 60.096 19.764 61.128 ; 
      RECT 18.884 57.186 19.276 61.56 ; 
      RECT 17.216 57.186 17.548 61.56 ; 
      RECT 17.216 57.54 17.604 61.282 ; 
      RECT 38.108 57.186 38.448 61.56 ; 
      RECT 37.532 57.186 37.636 61.56 ; 
      RECT 37.1 57.186 37.204 61.56 ; 
      RECT 36.668 57.186 36.772 61.56 ; 
      RECT 36.236 57.186 36.34 61.56 ; 
      RECT 35.804 57.186 35.908 61.56 ; 
      RECT 35.372 57.186 35.476 61.56 ; 
      RECT 34.94 57.186 35.044 61.56 ; 
      RECT 34.508 57.186 34.612 61.56 ; 
      RECT 34.076 57.186 34.18 61.56 ; 
      RECT 33.644 57.186 33.748 61.56 ; 
      RECT 33.212 57.186 33.316 61.56 ; 
      RECT 32.78 57.186 32.884 61.56 ; 
      RECT 32.348 57.186 32.452 61.56 ; 
      RECT 31.916 57.186 32.02 61.56 ; 
      RECT 31.484 57.186 31.588 61.56 ; 
      RECT 31.052 57.186 31.156 61.56 ; 
      RECT 30.62 57.186 30.724 61.56 ; 
      RECT 30.188 57.186 30.292 61.56 ; 
      RECT 29.756 57.186 29.86 61.56 ; 
      RECT 29.324 57.186 29.428 61.56 ; 
      RECT 28.892 57.186 28.996 61.56 ; 
      RECT 28.46 57.186 28.564 61.56 ; 
      RECT 28.028 57.186 28.132 61.56 ; 
      RECT 27.596 57.186 27.7 61.56 ; 
      RECT 27.164 57.186 27.268 61.56 ; 
      RECT 26.732 57.186 26.836 61.56 ; 
      RECT 26.3 57.186 26.404 61.56 ; 
      RECT 25.868 57.186 25.972 61.56 ; 
      RECT 25.436 57.186 25.54 61.56 ; 
      RECT 25.004 57.186 25.108 61.56 ; 
      RECT 24.572 57.186 24.676 61.56 ; 
      RECT 24.14 57.186 24.244 61.56 ; 
      RECT 23.708 57.186 23.812 61.56 ; 
      RECT 22.856 57.186 23.164 61.56 ; 
      RECT 15.284 57.186 15.592 61.56 ; 
      RECT 14.636 57.186 14.74 61.56 ; 
      RECT 14.204 57.186 14.308 61.56 ; 
      RECT 13.772 57.186 13.876 61.56 ; 
      RECT 13.34 57.186 13.444 61.56 ; 
      RECT 12.908 57.186 13.012 61.56 ; 
      RECT 12.476 57.186 12.58 61.56 ; 
      RECT 12.044 57.186 12.148 61.56 ; 
      RECT 11.612 57.186 11.716 61.56 ; 
      RECT 11.18 57.186 11.284 61.56 ; 
      RECT 10.748 57.186 10.852 61.56 ; 
      RECT 10.316 57.186 10.42 61.56 ; 
      RECT 9.884 57.186 9.988 61.56 ; 
      RECT 9.452 57.186 9.556 61.56 ; 
      RECT 9.02 57.186 9.124 61.56 ; 
      RECT 8.588 57.186 8.692 61.56 ; 
      RECT 8.156 57.186 8.26 61.56 ; 
      RECT 7.724 57.186 7.828 61.56 ; 
      RECT 7.292 57.186 7.396 61.56 ; 
      RECT 6.86 57.186 6.964 61.56 ; 
      RECT 6.428 57.186 6.532 61.56 ; 
      RECT 5.996 57.186 6.1 61.56 ; 
      RECT 5.564 57.186 5.668 61.56 ; 
      RECT 5.132 57.186 5.236 61.56 ; 
      RECT 4.7 57.186 4.804 61.56 ; 
      RECT 4.268 57.186 4.372 61.56 ; 
      RECT 3.836 57.186 3.94 61.56 ; 
      RECT 3.404 57.186 3.508 61.56 ; 
      RECT 2.972 57.186 3.076 61.56 ; 
      RECT 2.54 57.186 2.644 61.56 ; 
      RECT 2.108 57.186 2.212 61.56 ; 
      RECT 1.676 57.186 1.78 61.56 ; 
      RECT 1.244 57.186 1.348 61.56 ; 
      RECT 0.812 57.186 0.916 61.56 ; 
      RECT 0 57.186 0.34 61.56 ; 
      RECT 20.72 61.506 21.232 65.88 ; 
      RECT 20.664 64.168 21.232 65.458 ; 
      RECT 20.072 63.076 20.32 65.88 ; 
      RECT 20.016 64.314 20.32 64.928 ; 
      RECT 20.072 61.506 20.176 65.88 ; 
      RECT 20.072 61.99 20.232 62.948 ; 
      RECT 20.072 61.506 20.32 61.862 ; 
      RECT 18.884 63.308 19.708 65.88 ; 
      RECT 19.604 61.506 19.708 65.88 ; 
      RECT 18.884 64.416 19.764 65.448 ; 
      RECT 18.884 61.506 19.276 65.88 ; 
      RECT 17.216 61.506 17.548 65.88 ; 
      RECT 17.216 61.86 17.604 65.602 ; 
      RECT 38.108 61.506 38.448 65.88 ; 
      RECT 37.532 61.506 37.636 65.88 ; 
      RECT 37.1 61.506 37.204 65.88 ; 
      RECT 36.668 61.506 36.772 65.88 ; 
      RECT 36.236 61.506 36.34 65.88 ; 
      RECT 35.804 61.506 35.908 65.88 ; 
      RECT 35.372 61.506 35.476 65.88 ; 
      RECT 34.94 61.506 35.044 65.88 ; 
      RECT 34.508 61.506 34.612 65.88 ; 
      RECT 34.076 61.506 34.18 65.88 ; 
      RECT 33.644 61.506 33.748 65.88 ; 
      RECT 33.212 61.506 33.316 65.88 ; 
      RECT 32.78 61.506 32.884 65.88 ; 
      RECT 32.348 61.506 32.452 65.88 ; 
      RECT 31.916 61.506 32.02 65.88 ; 
      RECT 31.484 61.506 31.588 65.88 ; 
      RECT 31.052 61.506 31.156 65.88 ; 
      RECT 30.62 61.506 30.724 65.88 ; 
      RECT 30.188 61.506 30.292 65.88 ; 
      RECT 29.756 61.506 29.86 65.88 ; 
      RECT 29.324 61.506 29.428 65.88 ; 
      RECT 28.892 61.506 28.996 65.88 ; 
      RECT 28.46 61.506 28.564 65.88 ; 
      RECT 28.028 61.506 28.132 65.88 ; 
      RECT 27.596 61.506 27.7 65.88 ; 
      RECT 27.164 61.506 27.268 65.88 ; 
      RECT 26.732 61.506 26.836 65.88 ; 
      RECT 26.3 61.506 26.404 65.88 ; 
      RECT 25.868 61.506 25.972 65.88 ; 
      RECT 25.436 61.506 25.54 65.88 ; 
      RECT 25.004 61.506 25.108 65.88 ; 
      RECT 24.572 61.506 24.676 65.88 ; 
      RECT 24.14 61.506 24.244 65.88 ; 
      RECT 23.708 61.506 23.812 65.88 ; 
      RECT 22.856 61.506 23.164 65.88 ; 
      RECT 15.284 61.506 15.592 65.88 ; 
      RECT 14.636 61.506 14.74 65.88 ; 
      RECT 14.204 61.506 14.308 65.88 ; 
      RECT 13.772 61.506 13.876 65.88 ; 
      RECT 13.34 61.506 13.444 65.88 ; 
      RECT 12.908 61.506 13.012 65.88 ; 
      RECT 12.476 61.506 12.58 65.88 ; 
      RECT 12.044 61.506 12.148 65.88 ; 
      RECT 11.612 61.506 11.716 65.88 ; 
      RECT 11.18 61.506 11.284 65.88 ; 
      RECT 10.748 61.506 10.852 65.88 ; 
      RECT 10.316 61.506 10.42 65.88 ; 
      RECT 9.884 61.506 9.988 65.88 ; 
      RECT 9.452 61.506 9.556 65.88 ; 
      RECT 9.02 61.506 9.124 65.88 ; 
      RECT 8.588 61.506 8.692 65.88 ; 
      RECT 8.156 61.506 8.26 65.88 ; 
      RECT 7.724 61.506 7.828 65.88 ; 
      RECT 7.292 61.506 7.396 65.88 ; 
      RECT 6.86 61.506 6.964 65.88 ; 
      RECT 6.428 61.506 6.532 65.88 ; 
      RECT 5.996 61.506 6.1 65.88 ; 
      RECT 5.564 61.506 5.668 65.88 ; 
      RECT 5.132 61.506 5.236 65.88 ; 
      RECT 4.7 61.506 4.804 65.88 ; 
      RECT 4.268 61.506 4.372 65.88 ; 
      RECT 3.836 61.506 3.94 65.88 ; 
      RECT 3.404 61.506 3.508 65.88 ; 
      RECT 2.972 61.506 3.076 65.88 ; 
      RECT 2.54 61.506 2.644 65.88 ; 
      RECT 2.108 61.506 2.212 65.88 ; 
      RECT 1.676 61.506 1.78 65.88 ; 
      RECT 1.244 61.506 1.348 65.88 ; 
      RECT 0.812 61.506 0.916 65.88 ; 
      RECT 0 61.506 0.34 65.88 ; 
      RECT 20.72 65.826 21.232 70.2 ; 
      RECT 20.664 68.488 21.232 69.778 ; 
      RECT 20.072 67.396 20.32 70.2 ; 
      RECT 20.016 68.634 20.32 69.248 ; 
      RECT 20.072 65.826 20.176 70.2 ; 
      RECT 20.072 66.31 20.232 67.268 ; 
      RECT 20.072 65.826 20.32 66.182 ; 
      RECT 18.884 67.628 19.708 70.2 ; 
      RECT 19.604 65.826 19.708 70.2 ; 
      RECT 18.884 68.736 19.764 69.768 ; 
      RECT 18.884 65.826 19.276 70.2 ; 
      RECT 17.216 65.826 17.548 70.2 ; 
      RECT 17.216 66.18 17.604 69.922 ; 
      RECT 38.108 65.826 38.448 70.2 ; 
      RECT 37.532 65.826 37.636 70.2 ; 
      RECT 37.1 65.826 37.204 70.2 ; 
      RECT 36.668 65.826 36.772 70.2 ; 
      RECT 36.236 65.826 36.34 70.2 ; 
      RECT 35.804 65.826 35.908 70.2 ; 
      RECT 35.372 65.826 35.476 70.2 ; 
      RECT 34.94 65.826 35.044 70.2 ; 
      RECT 34.508 65.826 34.612 70.2 ; 
      RECT 34.076 65.826 34.18 70.2 ; 
      RECT 33.644 65.826 33.748 70.2 ; 
      RECT 33.212 65.826 33.316 70.2 ; 
      RECT 32.78 65.826 32.884 70.2 ; 
      RECT 32.348 65.826 32.452 70.2 ; 
      RECT 31.916 65.826 32.02 70.2 ; 
      RECT 31.484 65.826 31.588 70.2 ; 
      RECT 31.052 65.826 31.156 70.2 ; 
      RECT 30.62 65.826 30.724 70.2 ; 
      RECT 30.188 65.826 30.292 70.2 ; 
      RECT 29.756 65.826 29.86 70.2 ; 
      RECT 29.324 65.826 29.428 70.2 ; 
      RECT 28.892 65.826 28.996 70.2 ; 
      RECT 28.46 65.826 28.564 70.2 ; 
      RECT 28.028 65.826 28.132 70.2 ; 
      RECT 27.596 65.826 27.7 70.2 ; 
      RECT 27.164 65.826 27.268 70.2 ; 
      RECT 26.732 65.826 26.836 70.2 ; 
      RECT 26.3 65.826 26.404 70.2 ; 
      RECT 25.868 65.826 25.972 70.2 ; 
      RECT 25.436 65.826 25.54 70.2 ; 
      RECT 25.004 65.826 25.108 70.2 ; 
      RECT 24.572 65.826 24.676 70.2 ; 
      RECT 24.14 65.826 24.244 70.2 ; 
      RECT 23.708 65.826 23.812 70.2 ; 
      RECT 22.856 65.826 23.164 70.2 ; 
      RECT 15.284 65.826 15.592 70.2 ; 
      RECT 14.636 65.826 14.74 70.2 ; 
      RECT 14.204 65.826 14.308 70.2 ; 
      RECT 13.772 65.826 13.876 70.2 ; 
      RECT 13.34 65.826 13.444 70.2 ; 
      RECT 12.908 65.826 13.012 70.2 ; 
      RECT 12.476 65.826 12.58 70.2 ; 
      RECT 12.044 65.826 12.148 70.2 ; 
      RECT 11.612 65.826 11.716 70.2 ; 
      RECT 11.18 65.826 11.284 70.2 ; 
      RECT 10.748 65.826 10.852 70.2 ; 
      RECT 10.316 65.826 10.42 70.2 ; 
      RECT 9.884 65.826 9.988 70.2 ; 
      RECT 9.452 65.826 9.556 70.2 ; 
      RECT 9.02 65.826 9.124 70.2 ; 
      RECT 8.588 65.826 8.692 70.2 ; 
      RECT 8.156 65.826 8.26 70.2 ; 
      RECT 7.724 65.826 7.828 70.2 ; 
      RECT 7.292 65.826 7.396 70.2 ; 
      RECT 6.86 65.826 6.964 70.2 ; 
      RECT 6.428 65.826 6.532 70.2 ; 
      RECT 5.996 65.826 6.1 70.2 ; 
      RECT 5.564 65.826 5.668 70.2 ; 
      RECT 5.132 65.826 5.236 70.2 ; 
      RECT 4.7 65.826 4.804 70.2 ; 
      RECT 4.268 65.826 4.372 70.2 ; 
      RECT 3.836 65.826 3.94 70.2 ; 
      RECT 3.404 65.826 3.508 70.2 ; 
      RECT 2.972 65.826 3.076 70.2 ; 
      RECT 2.54 65.826 2.644 70.2 ; 
      RECT 2.108 65.826 2.212 70.2 ; 
      RECT 1.676 65.826 1.78 70.2 ; 
      RECT 1.244 65.826 1.348 70.2 ; 
      RECT 0.812 65.826 0.916 70.2 ; 
      RECT 0 65.826 0.34 70.2 ; 
      RECT 20.72 70.146 21.232 74.52 ; 
      RECT 20.664 72.808 21.232 74.098 ; 
      RECT 20.072 71.716 20.32 74.52 ; 
      RECT 20.016 72.954 20.32 73.568 ; 
      RECT 20.072 70.146 20.176 74.52 ; 
      RECT 20.072 70.63 20.232 71.588 ; 
      RECT 20.072 70.146 20.32 70.502 ; 
      RECT 18.884 71.948 19.708 74.52 ; 
      RECT 19.604 70.146 19.708 74.52 ; 
      RECT 18.884 73.056 19.764 74.088 ; 
      RECT 18.884 70.146 19.276 74.52 ; 
      RECT 17.216 70.146 17.548 74.52 ; 
      RECT 17.216 70.5 17.604 74.242 ; 
      RECT 38.108 70.146 38.448 74.52 ; 
      RECT 37.532 70.146 37.636 74.52 ; 
      RECT 37.1 70.146 37.204 74.52 ; 
      RECT 36.668 70.146 36.772 74.52 ; 
      RECT 36.236 70.146 36.34 74.52 ; 
      RECT 35.804 70.146 35.908 74.52 ; 
      RECT 35.372 70.146 35.476 74.52 ; 
      RECT 34.94 70.146 35.044 74.52 ; 
      RECT 34.508 70.146 34.612 74.52 ; 
      RECT 34.076 70.146 34.18 74.52 ; 
      RECT 33.644 70.146 33.748 74.52 ; 
      RECT 33.212 70.146 33.316 74.52 ; 
      RECT 32.78 70.146 32.884 74.52 ; 
      RECT 32.348 70.146 32.452 74.52 ; 
      RECT 31.916 70.146 32.02 74.52 ; 
      RECT 31.484 70.146 31.588 74.52 ; 
      RECT 31.052 70.146 31.156 74.52 ; 
      RECT 30.62 70.146 30.724 74.52 ; 
      RECT 30.188 70.146 30.292 74.52 ; 
      RECT 29.756 70.146 29.86 74.52 ; 
      RECT 29.324 70.146 29.428 74.52 ; 
      RECT 28.892 70.146 28.996 74.52 ; 
      RECT 28.46 70.146 28.564 74.52 ; 
      RECT 28.028 70.146 28.132 74.52 ; 
      RECT 27.596 70.146 27.7 74.52 ; 
      RECT 27.164 70.146 27.268 74.52 ; 
      RECT 26.732 70.146 26.836 74.52 ; 
      RECT 26.3 70.146 26.404 74.52 ; 
      RECT 25.868 70.146 25.972 74.52 ; 
      RECT 25.436 70.146 25.54 74.52 ; 
      RECT 25.004 70.146 25.108 74.52 ; 
      RECT 24.572 70.146 24.676 74.52 ; 
      RECT 24.14 70.146 24.244 74.52 ; 
      RECT 23.708 70.146 23.812 74.52 ; 
      RECT 22.856 70.146 23.164 74.52 ; 
      RECT 15.284 70.146 15.592 74.52 ; 
      RECT 14.636 70.146 14.74 74.52 ; 
      RECT 14.204 70.146 14.308 74.52 ; 
      RECT 13.772 70.146 13.876 74.52 ; 
      RECT 13.34 70.146 13.444 74.52 ; 
      RECT 12.908 70.146 13.012 74.52 ; 
      RECT 12.476 70.146 12.58 74.52 ; 
      RECT 12.044 70.146 12.148 74.52 ; 
      RECT 11.612 70.146 11.716 74.52 ; 
      RECT 11.18 70.146 11.284 74.52 ; 
      RECT 10.748 70.146 10.852 74.52 ; 
      RECT 10.316 70.146 10.42 74.52 ; 
      RECT 9.884 70.146 9.988 74.52 ; 
      RECT 9.452 70.146 9.556 74.52 ; 
      RECT 9.02 70.146 9.124 74.52 ; 
      RECT 8.588 70.146 8.692 74.52 ; 
      RECT 8.156 70.146 8.26 74.52 ; 
      RECT 7.724 70.146 7.828 74.52 ; 
      RECT 7.292 70.146 7.396 74.52 ; 
      RECT 6.86 70.146 6.964 74.52 ; 
      RECT 6.428 70.146 6.532 74.52 ; 
      RECT 5.996 70.146 6.1 74.52 ; 
      RECT 5.564 70.146 5.668 74.52 ; 
      RECT 5.132 70.146 5.236 74.52 ; 
      RECT 4.7 70.146 4.804 74.52 ; 
      RECT 4.268 70.146 4.372 74.52 ; 
      RECT 3.836 70.146 3.94 74.52 ; 
      RECT 3.404 70.146 3.508 74.52 ; 
      RECT 2.972 70.146 3.076 74.52 ; 
      RECT 2.54 70.146 2.644 74.52 ; 
      RECT 2.108 70.146 2.212 74.52 ; 
      RECT 1.676 70.146 1.78 74.52 ; 
      RECT 1.244 70.146 1.348 74.52 ; 
      RECT 0.812 70.146 0.916 74.52 ; 
      RECT 0 70.146 0.34 74.52 ; 
      RECT 20.72 74.466 21.232 78.84 ; 
      RECT 20.664 77.128 21.232 78.418 ; 
      RECT 20.072 76.036 20.32 78.84 ; 
      RECT 20.016 77.274 20.32 77.888 ; 
      RECT 20.072 74.466 20.176 78.84 ; 
      RECT 20.072 74.95 20.232 75.908 ; 
      RECT 20.072 74.466 20.32 74.822 ; 
      RECT 18.884 76.268 19.708 78.84 ; 
      RECT 19.604 74.466 19.708 78.84 ; 
      RECT 18.884 77.376 19.764 78.408 ; 
      RECT 18.884 74.466 19.276 78.84 ; 
      RECT 17.216 74.466 17.548 78.84 ; 
      RECT 17.216 74.82 17.604 78.562 ; 
      RECT 38.108 74.466 38.448 78.84 ; 
      RECT 37.532 74.466 37.636 78.84 ; 
      RECT 37.1 74.466 37.204 78.84 ; 
      RECT 36.668 74.466 36.772 78.84 ; 
      RECT 36.236 74.466 36.34 78.84 ; 
      RECT 35.804 74.466 35.908 78.84 ; 
      RECT 35.372 74.466 35.476 78.84 ; 
      RECT 34.94 74.466 35.044 78.84 ; 
      RECT 34.508 74.466 34.612 78.84 ; 
      RECT 34.076 74.466 34.18 78.84 ; 
      RECT 33.644 74.466 33.748 78.84 ; 
      RECT 33.212 74.466 33.316 78.84 ; 
      RECT 32.78 74.466 32.884 78.84 ; 
      RECT 32.348 74.466 32.452 78.84 ; 
      RECT 31.916 74.466 32.02 78.84 ; 
      RECT 31.484 74.466 31.588 78.84 ; 
      RECT 31.052 74.466 31.156 78.84 ; 
      RECT 30.62 74.466 30.724 78.84 ; 
      RECT 30.188 74.466 30.292 78.84 ; 
      RECT 29.756 74.466 29.86 78.84 ; 
      RECT 29.324 74.466 29.428 78.84 ; 
      RECT 28.892 74.466 28.996 78.84 ; 
      RECT 28.46 74.466 28.564 78.84 ; 
      RECT 28.028 74.466 28.132 78.84 ; 
      RECT 27.596 74.466 27.7 78.84 ; 
      RECT 27.164 74.466 27.268 78.84 ; 
      RECT 26.732 74.466 26.836 78.84 ; 
      RECT 26.3 74.466 26.404 78.84 ; 
      RECT 25.868 74.466 25.972 78.84 ; 
      RECT 25.436 74.466 25.54 78.84 ; 
      RECT 25.004 74.466 25.108 78.84 ; 
      RECT 24.572 74.466 24.676 78.84 ; 
      RECT 24.14 74.466 24.244 78.84 ; 
      RECT 23.708 74.466 23.812 78.84 ; 
      RECT 22.856 74.466 23.164 78.84 ; 
      RECT 15.284 74.466 15.592 78.84 ; 
      RECT 14.636 74.466 14.74 78.84 ; 
      RECT 14.204 74.466 14.308 78.84 ; 
      RECT 13.772 74.466 13.876 78.84 ; 
      RECT 13.34 74.466 13.444 78.84 ; 
      RECT 12.908 74.466 13.012 78.84 ; 
      RECT 12.476 74.466 12.58 78.84 ; 
      RECT 12.044 74.466 12.148 78.84 ; 
      RECT 11.612 74.466 11.716 78.84 ; 
      RECT 11.18 74.466 11.284 78.84 ; 
      RECT 10.748 74.466 10.852 78.84 ; 
      RECT 10.316 74.466 10.42 78.84 ; 
      RECT 9.884 74.466 9.988 78.84 ; 
      RECT 9.452 74.466 9.556 78.84 ; 
      RECT 9.02 74.466 9.124 78.84 ; 
      RECT 8.588 74.466 8.692 78.84 ; 
      RECT 8.156 74.466 8.26 78.84 ; 
      RECT 7.724 74.466 7.828 78.84 ; 
      RECT 7.292 74.466 7.396 78.84 ; 
      RECT 6.86 74.466 6.964 78.84 ; 
      RECT 6.428 74.466 6.532 78.84 ; 
      RECT 5.996 74.466 6.1 78.84 ; 
      RECT 5.564 74.466 5.668 78.84 ; 
      RECT 5.132 74.466 5.236 78.84 ; 
      RECT 4.7 74.466 4.804 78.84 ; 
      RECT 4.268 74.466 4.372 78.84 ; 
      RECT 3.836 74.466 3.94 78.84 ; 
      RECT 3.404 74.466 3.508 78.84 ; 
      RECT 2.972 74.466 3.076 78.84 ; 
      RECT 2.54 74.466 2.644 78.84 ; 
      RECT 2.108 74.466 2.212 78.84 ; 
      RECT 1.676 74.466 1.78 78.84 ; 
      RECT 1.244 74.466 1.348 78.84 ; 
      RECT 0.812 74.466 0.916 78.84 ; 
      RECT 0 74.466 0.34 78.84 ; 
      RECT 20.72 78.786 21.232 83.16 ; 
      RECT 20.664 81.448 21.232 82.738 ; 
      RECT 20.072 80.356 20.32 83.16 ; 
      RECT 20.016 81.594 20.32 82.208 ; 
      RECT 20.072 78.786 20.176 83.16 ; 
      RECT 20.072 79.27 20.232 80.228 ; 
      RECT 20.072 78.786 20.32 79.142 ; 
      RECT 18.884 80.588 19.708 83.16 ; 
      RECT 19.604 78.786 19.708 83.16 ; 
      RECT 18.884 81.696 19.764 82.728 ; 
      RECT 18.884 78.786 19.276 83.16 ; 
      RECT 17.216 78.786 17.548 83.16 ; 
      RECT 17.216 79.14 17.604 82.882 ; 
      RECT 38.108 78.786 38.448 83.16 ; 
      RECT 37.532 78.786 37.636 83.16 ; 
      RECT 37.1 78.786 37.204 83.16 ; 
      RECT 36.668 78.786 36.772 83.16 ; 
      RECT 36.236 78.786 36.34 83.16 ; 
      RECT 35.804 78.786 35.908 83.16 ; 
      RECT 35.372 78.786 35.476 83.16 ; 
      RECT 34.94 78.786 35.044 83.16 ; 
      RECT 34.508 78.786 34.612 83.16 ; 
      RECT 34.076 78.786 34.18 83.16 ; 
      RECT 33.644 78.786 33.748 83.16 ; 
      RECT 33.212 78.786 33.316 83.16 ; 
      RECT 32.78 78.786 32.884 83.16 ; 
      RECT 32.348 78.786 32.452 83.16 ; 
      RECT 31.916 78.786 32.02 83.16 ; 
      RECT 31.484 78.786 31.588 83.16 ; 
      RECT 31.052 78.786 31.156 83.16 ; 
      RECT 30.62 78.786 30.724 83.16 ; 
      RECT 30.188 78.786 30.292 83.16 ; 
      RECT 29.756 78.786 29.86 83.16 ; 
      RECT 29.324 78.786 29.428 83.16 ; 
      RECT 28.892 78.786 28.996 83.16 ; 
      RECT 28.46 78.786 28.564 83.16 ; 
      RECT 28.028 78.786 28.132 83.16 ; 
      RECT 27.596 78.786 27.7 83.16 ; 
      RECT 27.164 78.786 27.268 83.16 ; 
      RECT 26.732 78.786 26.836 83.16 ; 
      RECT 26.3 78.786 26.404 83.16 ; 
      RECT 25.868 78.786 25.972 83.16 ; 
      RECT 25.436 78.786 25.54 83.16 ; 
      RECT 25.004 78.786 25.108 83.16 ; 
      RECT 24.572 78.786 24.676 83.16 ; 
      RECT 24.14 78.786 24.244 83.16 ; 
      RECT 23.708 78.786 23.812 83.16 ; 
      RECT 22.856 78.786 23.164 83.16 ; 
      RECT 15.284 78.786 15.592 83.16 ; 
      RECT 14.636 78.786 14.74 83.16 ; 
      RECT 14.204 78.786 14.308 83.16 ; 
      RECT 13.772 78.786 13.876 83.16 ; 
      RECT 13.34 78.786 13.444 83.16 ; 
      RECT 12.908 78.786 13.012 83.16 ; 
      RECT 12.476 78.786 12.58 83.16 ; 
      RECT 12.044 78.786 12.148 83.16 ; 
      RECT 11.612 78.786 11.716 83.16 ; 
      RECT 11.18 78.786 11.284 83.16 ; 
      RECT 10.748 78.786 10.852 83.16 ; 
      RECT 10.316 78.786 10.42 83.16 ; 
      RECT 9.884 78.786 9.988 83.16 ; 
      RECT 9.452 78.786 9.556 83.16 ; 
      RECT 9.02 78.786 9.124 83.16 ; 
      RECT 8.588 78.786 8.692 83.16 ; 
      RECT 8.156 78.786 8.26 83.16 ; 
      RECT 7.724 78.786 7.828 83.16 ; 
      RECT 7.292 78.786 7.396 83.16 ; 
      RECT 6.86 78.786 6.964 83.16 ; 
      RECT 6.428 78.786 6.532 83.16 ; 
      RECT 5.996 78.786 6.1 83.16 ; 
      RECT 5.564 78.786 5.668 83.16 ; 
      RECT 5.132 78.786 5.236 83.16 ; 
      RECT 4.7 78.786 4.804 83.16 ; 
      RECT 4.268 78.786 4.372 83.16 ; 
      RECT 3.836 78.786 3.94 83.16 ; 
      RECT 3.404 78.786 3.508 83.16 ; 
      RECT 2.972 78.786 3.076 83.16 ; 
      RECT 2.54 78.786 2.644 83.16 ; 
      RECT 2.108 78.786 2.212 83.16 ; 
      RECT 1.676 78.786 1.78 83.16 ; 
      RECT 1.244 78.786 1.348 83.16 ; 
      RECT 0.812 78.786 0.916 83.16 ; 
      RECT 0 78.786 0.34 83.16 ; 
      RECT 20.72 83.106 21.232 87.48 ; 
      RECT 20.664 85.768 21.232 87.058 ; 
      RECT 20.072 84.676 20.32 87.48 ; 
      RECT 20.016 85.914 20.32 86.528 ; 
      RECT 20.072 83.106 20.176 87.48 ; 
      RECT 20.072 83.59 20.232 84.548 ; 
      RECT 20.072 83.106 20.32 83.462 ; 
      RECT 18.884 84.908 19.708 87.48 ; 
      RECT 19.604 83.106 19.708 87.48 ; 
      RECT 18.884 86.016 19.764 87.048 ; 
      RECT 18.884 83.106 19.276 87.48 ; 
      RECT 17.216 83.106 17.548 87.48 ; 
      RECT 17.216 83.46 17.604 87.202 ; 
      RECT 38.108 83.106 38.448 87.48 ; 
      RECT 37.532 83.106 37.636 87.48 ; 
      RECT 37.1 83.106 37.204 87.48 ; 
      RECT 36.668 83.106 36.772 87.48 ; 
      RECT 36.236 83.106 36.34 87.48 ; 
      RECT 35.804 83.106 35.908 87.48 ; 
      RECT 35.372 83.106 35.476 87.48 ; 
      RECT 34.94 83.106 35.044 87.48 ; 
      RECT 34.508 83.106 34.612 87.48 ; 
      RECT 34.076 83.106 34.18 87.48 ; 
      RECT 33.644 83.106 33.748 87.48 ; 
      RECT 33.212 83.106 33.316 87.48 ; 
      RECT 32.78 83.106 32.884 87.48 ; 
      RECT 32.348 83.106 32.452 87.48 ; 
      RECT 31.916 83.106 32.02 87.48 ; 
      RECT 31.484 83.106 31.588 87.48 ; 
      RECT 31.052 83.106 31.156 87.48 ; 
      RECT 30.62 83.106 30.724 87.48 ; 
      RECT 30.188 83.106 30.292 87.48 ; 
      RECT 29.756 83.106 29.86 87.48 ; 
      RECT 29.324 83.106 29.428 87.48 ; 
      RECT 28.892 83.106 28.996 87.48 ; 
      RECT 28.46 83.106 28.564 87.48 ; 
      RECT 28.028 83.106 28.132 87.48 ; 
      RECT 27.596 83.106 27.7 87.48 ; 
      RECT 27.164 83.106 27.268 87.48 ; 
      RECT 26.732 83.106 26.836 87.48 ; 
      RECT 26.3 83.106 26.404 87.48 ; 
      RECT 25.868 83.106 25.972 87.48 ; 
      RECT 25.436 83.106 25.54 87.48 ; 
      RECT 25.004 83.106 25.108 87.48 ; 
      RECT 24.572 83.106 24.676 87.48 ; 
      RECT 24.14 83.106 24.244 87.48 ; 
      RECT 23.708 83.106 23.812 87.48 ; 
      RECT 22.856 83.106 23.164 87.48 ; 
      RECT 15.284 83.106 15.592 87.48 ; 
      RECT 14.636 83.106 14.74 87.48 ; 
      RECT 14.204 83.106 14.308 87.48 ; 
      RECT 13.772 83.106 13.876 87.48 ; 
      RECT 13.34 83.106 13.444 87.48 ; 
      RECT 12.908 83.106 13.012 87.48 ; 
      RECT 12.476 83.106 12.58 87.48 ; 
      RECT 12.044 83.106 12.148 87.48 ; 
      RECT 11.612 83.106 11.716 87.48 ; 
      RECT 11.18 83.106 11.284 87.48 ; 
      RECT 10.748 83.106 10.852 87.48 ; 
      RECT 10.316 83.106 10.42 87.48 ; 
      RECT 9.884 83.106 9.988 87.48 ; 
      RECT 9.452 83.106 9.556 87.48 ; 
      RECT 9.02 83.106 9.124 87.48 ; 
      RECT 8.588 83.106 8.692 87.48 ; 
      RECT 8.156 83.106 8.26 87.48 ; 
      RECT 7.724 83.106 7.828 87.48 ; 
      RECT 7.292 83.106 7.396 87.48 ; 
      RECT 6.86 83.106 6.964 87.48 ; 
      RECT 6.428 83.106 6.532 87.48 ; 
      RECT 5.996 83.106 6.1 87.48 ; 
      RECT 5.564 83.106 5.668 87.48 ; 
      RECT 5.132 83.106 5.236 87.48 ; 
      RECT 4.7 83.106 4.804 87.48 ; 
      RECT 4.268 83.106 4.372 87.48 ; 
      RECT 3.836 83.106 3.94 87.48 ; 
      RECT 3.404 83.106 3.508 87.48 ; 
      RECT 2.972 83.106 3.076 87.48 ; 
      RECT 2.54 83.106 2.644 87.48 ; 
      RECT 2.108 83.106 2.212 87.48 ; 
      RECT 1.676 83.106 1.78 87.48 ; 
      RECT 1.244 83.106 1.348 87.48 ; 
      RECT 0.812 83.106 0.916 87.48 ; 
      RECT 0 83.106 0.34 87.48 ; 
      RECT 20.72 87.426 21.232 91.8 ; 
      RECT 20.664 90.088 21.232 91.378 ; 
      RECT 20.072 88.996 20.32 91.8 ; 
      RECT 20.016 90.234 20.32 90.848 ; 
      RECT 20.072 87.426 20.176 91.8 ; 
      RECT 20.072 87.91 20.232 88.868 ; 
      RECT 20.072 87.426 20.32 87.782 ; 
      RECT 18.884 89.228 19.708 91.8 ; 
      RECT 19.604 87.426 19.708 91.8 ; 
      RECT 18.884 90.336 19.764 91.368 ; 
      RECT 18.884 87.426 19.276 91.8 ; 
      RECT 17.216 87.426 17.548 91.8 ; 
      RECT 17.216 87.78 17.604 91.522 ; 
      RECT 38.108 87.426 38.448 91.8 ; 
      RECT 37.532 87.426 37.636 91.8 ; 
      RECT 37.1 87.426 37.204 91.8 ; 
      RECT 36.668 87.426 36.772 91.8 ; 
      RECT 36.236 87.426 36.34 91.8 ; 
      RECT 35.804 87.426 35.908 91.8 ; 
      RECT 35.372 87.426 35.476 91.8 ; 
      RECT 34.94 87.426 35.044 91.8 ; 
      RECT 34.508 87.426 34.612 91.8 ; 
      RECT 34.076 87.426 34.18 91.8 ; 
      RECT 33.644 87.426 33.748 91.8 ; 
      RECT 33.212 87.426 33.316 91.8 ; 
      RECT 32.78 87.426 32.884 91.8 ; 
      RECT 32.348 87.426 32.452 91.8 ; 
      RECT 31.916 87.426 32.02 91.8 ; 
      RECT 31.484 87.426 31.588 91.8 ; 
      RECT 31.052 87.426 31.156 91.8 ; 
      RECT 30.62 87.426 30.724 91.8 ; 
      RECT 30.188 87.426 30.292 91.8 ; 
      RECT 29.756 87.426 29.86 91.8 ; 
      RECT 29.324 87.426 29.428 91.8 ; 
      RECT 28.892 87.426 28.996 91.8 ; 
      RECT 28.46 87.426 28.564 91.8 ; 
      RECT 28.028 87.426 28.132 91.8 ; 
      RECT 27.596 87.426 27.7 91.8 ; 
      RECT 27.164 87.426 27.268 91.8 ; 
      RECT 26.732 87.426 26.836 91.8 ; 
      RECT 26.3 87.426 26.404 91.8 ; 
      RECT 25.868 87.426 25.972 91.8 ; 
      RECT 25.436 87.426 25.54 91.8 ; 
      RECT 25.004 87.426 25.108 91.8 ; 
      RECT 24.572 87.426 24.676 91.8 ; 
      RECT 24.14 87.426 24.244 91.8 ; 
      RECT 23.708 87.426 23.812 91.8 ; 
      RECT 22.856 87.426 23.164 91.8 ; 
      RECT 15.284 87.426 15.592 91.8 ; 
      RECT 14.636 87.426 14.74 91.8 ; 
      RECT 14.204 87.426 14.308 91.8 ; 
      RECT 13.772 87.426 13.876 91.8 ; 
      RECT 13.34 87.426 13.444 91.8 ; 
      RECT 12.908 87.426 13.012 91.8 ; 
      RECT 12.476 87.426 12.58 91.8 ; 
      RECT 12.044 87.426 12.148 91.8 ; 
      RECT 11.612 87.426 11.716 91.8 ; 
      RECT 11.18 87.426 11.284 91.8 ; 
      RECT 10.748 87.426 10.852 91.8 ; 
      RECT 10.316 87.426 10.42 91.8 ; 
      RECT 9.884 87.426 9.988 91.8 ; 
      RECT 9.452 87.426 9.556 91.8 ; 
      RECT 9.02 87.426 9.124 91.8 ; 
      RECT 8.588 87.426 8.692 91.8 ; 
      RECT 8.156 87.426 8.26 91.8 ; 
      RECT 7.724 87.426 7.828 91.8 ; 
      RECT 7.292 87.426 7.396 91.8 ; 
      RECT 6.86 87.426 6.964 91.8 ; 
      RECT 6.428 87.426 6.532 91.8 ; 
      RECT 5.996 87.426 6.1 91.8 ; 
      RECT 5.564 87.426 5.668 91.8 ; 
      RECT 5.132 87.426 5.236 91.8 ; 
      RECT 4.7 87.426 4.804 91.8 ; 
      RECT 4.268 87.426 4.372 91.8 ; 
      RECT 3.836 87.426 3.94 91.8 ; 
      RECT 3.404 87.426 3.508 91.8 ; 
      RECT 2.972 87.426 3.076 91.8 ; 
      RECT 2.54 87.426 2.644 91.8 ; 
      RECT 2.108 87.426 2.212 91.8 ; 
      RECT 1.676 87.426 1.78 91.8 ; 
      RECT 1.244 87.426 1.348 91.8 ; 
      RECT 0.812 87.426 0.916 91.8 ; 
      RECT 0 87.426 0.34 91.8 ; 
      RECT 20.72 91.746 21.232 96.12 ; 
      RECT 20.664 94.408 21.232 95.698 ; 
      RECT 20.072 93.316 20.32 96.12 ; 
      RECT 20.016 94.554 20.32 95.168 ; 
      RECT 20.072 91.746 20.176 96.12 ; 
      RECT 20.072 92.23 20.232 93.188 ; 
      RECT 20.072 91.746 20.32 92.102 ; 
      RECT 18.884 93.548 19.708 96.12 ; 
      RECT 19.604 91.746 19.708 96.12 ; 
      RECT 18.884 94.656 19.764 95.688 ; 
      RECT 18.884 91.746 19.276 96.12 ; 
      RECT 17.216 91.746 17.548 96.12 ; 
      RECT 17.216 92.1 17.604 95.842 ; 
      RECT 38.108 91.746 38.448 96.12 ; 
      RECT 37.532 91.746 37.636 96.12 ; 
      RECT 37.1 91.746 37.204 96.12 ; 
      RECT 36.668 91.746 36.772 96.12 ; 
      RECT 36.236 91.746 36.34 96.12 ; 
      RECT 35.804 91.746 35.908 96.12 ; 
      RECT 35.372 91.746 35.476 96.12 ; 
      RECT 34.94 91.746 35.044 96.12 ; 
      RECT 34.508 91.746 34.612 96.12 ; 
      RECT 34.076 91.746 34.18 96.12 ; 
      RECT 33.644 91.746 33.748 96.12 ; 
      RECT 33.212 91.746 33.316 96.12 ; 
      RECT 32.78 91.746 32.884 96.12 ; 
      RECT 32.348 91.746 32.452 96.12 ; 
      RECT 31.916 91.746 32.02 96.12 ; 
      RECT 31.484 91.746 31.588 96.12 ; 
      RECT 31.052 91.746 31.156 96.12 ; 
      RECT 30.62 91.746 30.724 96.12 ; 
      RECT 30.188 91.746 30.292 96.12 ; 
      RECT 29.756 91.746 29.86 96.12 ; 
      RECT 29.324 91.746 29.428 96.12 ; 
      RECT 28.892 91.746 28.996 96.12 ; 
      RECT 28.46 91.746 28.564 96.12 ; 
      RECT 28.028 91.746 28.132 96.12 ; 
      RECT 27.596 91.746 27.7 96.12 ; 
      RECT 27.164 91.746 27.268 96.12 ; 
      RECT 26.732 91.746 26.836 96.12 ; 
      RECT 26.3 91.746 26.404 96.12 ; 
      RECT 25.868 91.746 25.972 96.12 ; 
      RECT 25.436 91.746 25.54 96.12 ; 
      RECT 25.004 91.746 25.108 96.12 ; 
      RECT 24.572 91.746 24.676 96.12 ; 
      RECT 24.14 91.746 24.244 96.12 ; 
      RECT 23.708 91.746 23.812 96.12 ; 
      RECT 22.856 91.746 23.164 96.12 ; 
      RECT 15.284 91.746 15.592 96.12 ; 
      RECT 14.636 91.746 14.74 96.12 ; 
      RECT 14.204 91.746 14.308 96.12 ; 
      RECT 13.772 91.746 13.876 96.12 ; 
      RECT 13.34 91.746 13.444 96.12 ; 
      RECT 12.908 91.746 13.012 96.12 ; 
      RECT 12.476 91.746 12.58 96.12 ; 
      RECT 12.044 91.746 12.148 96.12 ; 
      RECT 11.612 91.746 11.716 96.12 ; 
      RECT 11.18 91.746 11.284 96.12 ; 
      RECT 10.748 91.746 10.852 96.12 ; 
      RECT 10.316 91.746 10.42 96.12 ; 
      RECT 9.884 91.746 9.988 96.12 ; 
      RECT 9.452 91.746 9.556 96.12 ; 
      RECT 9.02 91.746 9.124 96.12 ; 
      RECT 8.588 91.746 8.692 96.12 ; 
      RECT 8.156 91.746 8.26 96.12 ; 
      RECT 7.724 91.746 7.828 96.12 ; 
      RECT 7.292 91.746 7.396 96.12 ; 
      RECT 6.86 91.746 6.964 96.12 ; 
      RECT 6.428 91.746 6.532 96.12 ; 
      RECT 5.996 91.746 6.1 96.12 ; 
      RECT 5.564 91.746 5.668 96.12 ; 
      RECT 5.132 91.746 5.236 96.12 ; 
      RECT 4.7 91.746 4.804 96.12 ; 
      RECT 4.268 91.746 4.372 96.12 ; 
      RECT 3.836 91.746 3.94 96.12 ; 
      RECT 3.404 91.746 3.508 96.12 ; 
      RECT 2.972 91.746 3.076 96.12 ; 
      RECT 2.54 91.746 2.644 96.12 ; 
      RECT 2.108 91.746 2.212 96.12 ; 
      RECT 1.676 91.746 1.78 96.12 ; 
      RECT 1.244 91.746 1.348 96.12 ; 
      RECT 0.812 91.746 0.916 96.12 ; 
      RECT 0 91.746 0.34 96.12 ; 
      RECT 20.72 96.066 21.232 100.44 ; 
      RECT 20.664 98.728 21.232 100.018 ; 
      RECT 20.072 97.636 20.32 100.44 ; 
      RECT 20.016 98.874 20.32 99.488 ; 
      RECT 20.072 96.066 20.176 100.44 ; 
      RECT 20.072 96.55 20.232 97.508 ; 
      RECT 20.072 96.066 20.32 96.422 ; 
      RECT 18.884 97.868 19.708 100.44 ; 
      RECT 19.604 96.066 19.708 100.44 ; 
      RECT 18.884 98.976 19.764 100.008 ; 
      RECT 18.884 96.066 19.276 100.44 ; 
      RECT 17.216 96.066 17.548 100.44 ; 
      RECT 17.216 96.42 17.604 100.162 ; 
      RECT 38.108 96.066 38.448 100.44 ; 
      RECT 37.532 96.066 37.636 100.44 ; 
      RECT 37.1 96.066 37.204 100.44 ; 
      RECT 36.668 96.066 36.772 100.44 ; 
      RECT 36.236 96.066 36.34 100.44 ; 
      RECT 35.804 96.066 35.908 100.44 ; 
      RECT 35.372 96.066 35.476 100.44 ; 
      RECT 34.94 96.066 35.044 100.44 ; 
      RECT 34.508 96.066 34.612 100.44 ; 
      RECT 34.076 96.066 34.18 100.44 ; 
      RECT 33.644 96.066 33.748 100.44 ; 
      RECT 33.212 96.066 33.316 100.44 ; 
      RECT 32.78 96.066 32.884 100.44 ; 
      RECT 32.348 96.066 32.452 100.44 ; 
      RECT 31.916 96.066 32.02 100.44 ; 
      RECT 31.484 96.066 31.588 100.44 ; 
      RECT 31.052 96.066 31.156 100.44 ; 
      RECT 30.62 96.066 30.724 100.44 ; 
      RECT 30.188 96.066 30.292 100.44 ; 
      RECT 29.756 96.066 29.86 100.44 ; 
      RECT 29.324 96.066 29.428 100.44 ; 
      RECT 28.892 96.066 28.996 100.44 ; 
      RECT 28.46 96.066 28.564 100.44 ; 
      RECT 28.028 96.066 28.132 100.44 ; 
      RECT 27.596 96.066 27.7 100.44 ; 
      RECT 27.164 96.066 27.268 100.44 ; 
      RECT 26.732 96.066 26.836 100.44 ; 
      RECT 26.3 96.066 26.404 100.44 ; 
      RECT 25.868 96.066 25.972 100.44 ; 
      RECT 25.436 96.066 25.54 100.44 ; 
      RECT 25.004 96.066 25.108 100.44 ; 
      RECT 24.572 96.066 24.676 100.44 ; 
      RECT 24.14 96.066 24.244 100.44 ; 
      RECT 23.708 96.066 23.812 100.44 ; 
      RECT 22.856 96.066 23.164 100.44 ; 
      RECT 15.284 96.066 15.592 100.44 ; 
      RECT 14.636 96.066 14.74 100.44 ; 
      RECT 14.204 96.066 14.308 100.44 ; 
      RECT 13.772 96.066 13.876 100.44 ; 
      RECT 13.34 96.066 13.444 100.44 ; 
      RECT 12.908 96.066 13.012 100.44 ; 
      RECT 12.476 96.066 12.58 100.44 ; 
      RECT 12.044 96.066 12.148 100.44 ; 
      RECT 11.612 96.066 11.716 100.44 ; 
      RECT 11.18 96.066 11.284 100.44 ; 
      RECT 10.748 96.066 10.852 100.44 ; 
      RECT 10.316 96.066 10.42 100.44 ; 
      RECT 9.884 96.066 9.988 100.44 ; 
      RECT 9.452 96.066 9.556 100.44 ; 
      RECT 9.02 96.066 9.124 100.44 ; 
      RECT 8.588 96.066 8.692 100.44 ; 
      RECT 8.156 96.066 8.26 100.44 ; 
      RECT 7.724 96.066 7.828 100.44 ; 
      RECT 7.292 96.066 7.396 100.44 ; 
      RECT 6.86 96.066 6.964 100.44 ; 
      RECT 6.428 96.066 6.532 100.44 ; 
      RECT 5.996 96.066 6.1 100.44 ; 
      RECT 5.564 96.066 5.668 100.44 ; 
      RECT 5.132 96.066 5.236 100.44 ; 
      RECT 4.7 96.066 4.804 100.44 ; 
      RECT 4.268 96.066 4.372 100.44 ; 
      RECT 3.836 96.066 3.94 100.44 ; 
      RECT 3.404 96.066 3.508 100.44 ; 
      RECT 2.972 96.066 3.076 100.44 ; 
      RECT 2.54 96.066 2.644 100.44 ; 
      RECT 2.108 96.066 2.212 100.44 ; 
      RECT 1.676 96.066 1.78 100.44 ; 
      RECT 1.244 96.066 1.348 100.44 ; 
      RECT 0.812 96.066 0.916 100.44 ; 
      RECT 0 96.066 0.34 100.44 ; 
      RECT 20.72 100.386 21.232 104.76 ; 
      RECT 20.664 103.048 21.232 104.338 ; 
      RECT 20.072 101.956 20.32 104.76 ; 
      RECT 20.016 103.194 20.32 103.808 ; 
      RECT 20.072 100.386 20.176 104.76 ; 
      RECT 20.072 100.87 20.232 101.828 ; 
      RECT 20.072 100.386 20.32 100.742 ; 
      RECT 18.884 102.188 19.708 104.76 ; 
      RECT 19.604 100.386 19.708 104.76 ; 
      RECT 18.884 103.296 19.764 104.328 ; 
      RECT 18.884 100.386 19.276 104.76 ; 
      RECT 17.216 100.386 17.548 104.76 ; 
      RECT 17.216 100.74 17.604 104.482 ; 
      RECT 38.108 100.386 38.448 104.76 ; 
      RECT 37.532 100.386 37.636 104.76 ; 
      RECT 37.1 100.386 37.204 104.76 ; 
      RECT 36.668 100.386 36.772 104.76 ; 
      RECT 36.236 100.386 36.34 104.76 ; 
      RECT 35.804 100.386 35.908 104.76 ; 
      RECT 35.372 100.386 35.476 104.76 ; 
      RECT 34.94 100.386 35.044 104.76 ; 
      RECT 34.508 100.386 34.612 104.76 ; 
      RECT 34.076 100.386 34.18 104.76 ; 
      RECT 33.644 100.386 33.748 104.76 ; 
      RECT 33.212 100.386 33.316 104.76 ; 
      RECT 32.78 100.386 32.884 104.76 ; 
      RECT 32.348 100.386 32.452 104.76 ; 
      RECT 31.916 100.386 32.02 104.76 ; 
      RECT 31.484 100.386 31.588 104.76 ; 
      RECT 31.052 100.386 31.156 104.76 ; 
      RECT 30.62 100.386 30.724 104.76 ; 
      RECT 30.188 100.386 30.292 104.76 ; 
      RECT 29.756 100.386 29.86 104.76 ; 
      RECT 29.324 100.386 29.428 104.76 ; 
      RECT 28.892 100.386 28.996 104.76 ; 
      RECT 28.46 100.386 28.564 104.76 ; 
      RECT 28.028 100.386 28.132 104.76 ; 
      RECT 27.596 100.386 27.7 104.76 ; 
      RECT 27.164 100.386 27.268 104.76 ; 
      RECT 26.732 100.386 26.836 104.76 ; 
      RECT 26.3 100.386 26.404 104.76 ; 
      RECT 25.868 100.386 25.972 104.76 ; 
      RECT 25.436 100.386 25.54 104.76 ; 
      RECT 25.004 100.386 25.108 104.76 ; 
      RECT 24.572 100.386 24.676 104.76 ; 
      RECT 24.14 100.386 24.244 104.76 ; 
      RECT 23.708 100.386 23.812 104.76 ; 
      RECT 22.856 100.386 23.164 104.76 ; 
      RECT 15.284 100.386 15.592 104.76 ; 
      RECT 14.636 100.386 14.74 104.76 ; 
      RECT 14.204 100.386 14.308 104.76 ; 
      RECT 13.772 100.386 13.876 104.76 ; 
      RECT 13.34 100.386 13.444 104.76 ; 
      RECT 12.908 100.386 13.012 104.76 ; 
      RECT 12.476 100.386 12.58 104.76 ; 
      RECT 12.044 100.386 12.148 104.76 ; 
      RECT 11.612 100.386 11.716 104.76 ; 
      RECT 11.18 100.386 11.284 104.76 ; 
      RECT 10.748 100.386 10.852 104.76 ; 
      RECT 10.316 100.386 10.42 104.76 ; 
      RECT 9.884 100.386 9.988 104.76 ; 
      RECT 9.452 100.386 9.556 104.76 ; 
      RECT 9.02 100.386 9.124 104.76 ; 
      RECT 8.588 100.386 8.692 104.76 ; 
      RECT 8.156 100.386 8.26 104.76 ; 
      RECT 7.724 100.386 7.828 104.76 ; 
      RECT 7.292 100.386 7.396 104.76 ; 
      RECT 6.86 100.386 6.964 104.76 ; 
      RECT 6.428 100.386 6.532 104.76 ; 
      RECT 5.996 100.386 6.1 104.76 ; 
      RECT 5.564 100.386 5.668 104.76 ; 
      RECT 5.132 100.386 5.236 104.76 ; 
      RECT 4.7 100.386 4.804 104.76 ; 
      RECT 4.268 100.386 4.372 104.76 ; 
      RECT 3.836 100.386 3.94 104.76 ; 
      RECT 3.404 100.386 3.508 104.76 ; 
      RECT 2.972 100.386 3.076 104.76 ; 
      RECT 2.54 100.386 2.644 104.76 ; 
      RECT 2.108 100.386 2.212 104.76 ; 
      RECT 1.676 100.386 1.78 104.76 ; 
      RECT 1.244 100.386 1.348 104.76 ; 
      RECT 0.812 100.386 0.916 104.76 ; 
      RECT 0 100.386 0.34 104.76 ; 
      RECT 0 138.096 38.448 139.266 ; 
      RECT 38.108 104.652 38.448 139.266 ; 
      RECT 18.164 137.502 38.448 139.266 ; 
      RECT 0 137.502 17.548 139.266 ; 
      RECT 23.708 110.668 37.636 139.266 ; 
      RECT 29.54 104.652 37.636 139.266 ; 
      RECT 18.164 137.396 23.38 139.266 ; 
      RECT 20.72 137.392 23.38 139.266 ; 
      RECT 15.068 111.1 17.548 139.266 ; 
      RECT 15.284 107.716 17.548 139.266 ; 
      RECT 0.812 109.888 14.74 139.266 ; 
      RECT 13.556 104.652 14.74 139.266 ; 
      RECT 0 104.652 0.34 139.266 ; 
      RECT 18.164 137.384 20.32 139.266 ; 
      RECT 20.072 136.3 20.32 139.266 ; 
      RECT 20.72 136.3 23.164 139.266 ; 
      RECT 18.164 136.3 19.708 139.266 ; 
      RECT 23.652 119.824 37.636 137.264 ; 
      RECT 0.812 119.824 14.796 137.264 ; 
      RECT 23.652 119.824 37.692 137.246 ; 
      RECT 0.756 119.824 14.796 137.246 ; 
      RECT 20.756 107.716 23.164 139.266 ; 
      RECT 18.884 107.392 19.564 139.266 ; 
      RECT 19.316 104.652 19.564 139.266 ; 
      RECT 16.148 106.988 17.692 135.7 ; 
      RECT 15.068 135.532 17.748 135.68 ; 
      RECT 20.7 131.236 23.164 135.668 ; 
      RECT 18.828 134.476 19.564 135.38 ; 
      RECT 18.884 132.172 19.62 133.22 ; 
      RECT 15.068 131.38 17.748 133.22 ; 
      RECT 18.828 129.22 19.564 131.06 ; 
      RECT 20.7 121.084 23.164 130.412 ; 
      RECT 15.068 123.676 17.748 128.252 ; 
      RECT 18.884 122.596 19.62 127.82 ; 
      RECT 18.828 124.9 19.62 126.74 ; 
      RECT 18.828 111.94 19.564 124.58 ; 
      RECT 18.828 111.94 19.62 122.42 ; 
      RECT 15.068 121.516 17.748 122.42 ; 
      RECT 20.9 105.358 23.38 119.696 ; 
      RECT 20.7 109.78 23.38 116.924 ; 
      RECT 15.068 113.668 17.748 115.148 ; 
      RECT 18.884 110.86 19.62 111.62 ; 
      RECT 15.284 110.716 17.748 111.476 ; 
      RECT 18.828 110.284 19.564 110.828 ; 
      RECT 18.884 109.78 19.62 110.684 ; 
      RECT 24.356 109.9 37.636 139.266 ; 
      RECT 28.676 109.888 37.636 139.266 ; 
      RECT 23.708 104.652 24.028 139.266 ; 
      RECT 15.068 107.392 15.82 110.648 ; 
      RECT 23.708 104.652 24.892 110.264 ; 
      RECT 23.708 109.12 28.348 110.264 ; 
      RECT 28.676 104.652 29.212 139.266 ; 
      RECT 10.1 108.364 13.228 139.266 ; 
      RECT 0.812 104.652 9.772 139.266 ; 
      RECT 23.708 109.12 29.212 109.496 ; 
      RECT 27.812 104.652 37.636 109.484 ; 
      RECT 12.692 104.652 14.74 109.484 ; 
      RECT 18.828 109.204 19.62 109.46 ; 
      RECT 18.828 108.7 19.564 109.46 ; 
      RECT 26.948 107.584 37.636 109.484 ; 
      RECT 23.708 107.716 26.62 110.264 ; 
      RECT 18.884 107.62 19.62 108.668 ; 
      RECT 0.812 107.584 12.364 109.484 ; 
      RECT 11.828 104.652 12.364 139.266 ; 
      RECT 26.084 104.652 27.484 108.14 ; 
      RECT 23.708 107.392 25.756 110.264 ; 
      RECT 25.22 104.652 25.756 139.266 ; 
      RECT 10.964 107.392 12.364 139.266 ; 
      RECT 0.812 104.652 10.636 109.484 ; 
      RECT 18.884 104.652 18.988 139.266 ; 
      RECT 15.428 104.652 15.82 139.266 ; 
      RECT 10.964 104.652 11.5 139.266 ; 
      RECT 25.22 104.652 27.484 107.192 ; 
      RECT 20.756 104.652 23.164 107.192 ; 
      RECT 15.428 104.652 17.548 107.192 ; 
      RECT 11.828 104.652 14.74 107.192 ; 
      RECT 25.22 104.652 37.636 107.18 ; 
      RECT 0.812 104.652 11.5 107.18 ; 
      RECT 20.7 106.54 23.38 107.156 ; 
      RECT 15.428 106.54 17.604 107.192 ; 
      RECT 23.708 104.652 37.636 106.124 ; 
      RECT 18.884 104.652 19.564 106.124 ; 
      RECT 15.068 104.652 17.548 106.124 ; 
      RECT 0.812 104.652 14.74 106.124 ; 
      RECT 18.164 104.652 19.564 105.712 ; 
      RECT 20.72 104.652 23.164 105.312 ; 
      RECT 18.164 104.652 19.708 105.312 ; 
      RECT 20.72 104.652 23.38 104.736 ; 
      RECT 25.236 104.546 25.308 139.266 ; 
      RECT 24.804 104.546 24.876 139.266 ; 
      RECT 11.844 104.546 11.916 139.266 ; 
      RECT 11.412 104.546 11.484 139.266 ; 
      RECT 20.072 104.652 20.32 105.312 ; 
        RECT 20.72 137.214 21.232 141.588 ; 
        RECT 20.664 139.876 21.232 141.166 ; 
        RECT 20.072 138.784 20.32 141.588 ; 
        RECT 20.016 140.022 20.32 140.636 ; 
        RECT 20.072 137.214 20.176 141.588 ; 
        RECT 20.072 137.698 20.232 138.656 ; 
        RECT 20.072 137.214 20.32 137.57 ; 
        RECT 18.884 139.016 19.708 141.588 ; 
        RECT 19.604 137.214 19.708 141.588 ; 
        RECT 18.884 140.124 19.764 141.156 ; 
        RECT 18.884 137.214 19.276 141.588 ; 
        RECT 17.216 137.214 17.548 141.588 ; 
        RECT 17.216 137.568 17.604 141.31 ; 
        RECT 38.108 137.214 38.448 141.588 ; 
        RECT 37.532 137.214 37.636 141.588 ; 
        RECT 37.1 137.214 37.204 141.588 ; 
        RECT 36.668 137.214 36.772 141.588 ; 
        RECT 36.236 137.214 36.34 141.588 ; 
        RECT 35.804 137.214 35.908 141.588 ; 
        RECT 35.372 137.214 35.476 141.588 ; 
        RECT 34.94 137.214 35.044 141.588 ; 
        RECT 34.508 137.214 34.612 141.588 ; 
        RECT 34.076 137.214 34.18 141.588 ; 
        RECT 33.644 137.214 33.748 141.588 ; 
        RECT 33.212 137.214 33.316 141.588 ; 
        RECT 32.78 137.214 32.884 141.588 ; 
        RECT 32.348 137.214 32.452 141.588 ; 
        RECT 31.916 137.214 32.02 141.588 ; 
        RECT 31.484 137.214 31.588 141.588 ; 
        RECT 31.052 137.214 31.156 141.588 ; 
        RECT 30.62 137.214 30.724 141.588 ; 
        RECT 30.188 137.214 30.292 141.588 ; 
        RECT 29.756 137.214 29.86 141.588 ; 
        RECT 29.324 137.214 29.428 141.588 ; 
        RECT 28.892 137.214 28.996 141.588 ; 
        RECT 28.46 137.214 28.564 141.588 ; 
        RECT 28.028 137.214 28.132 141.588 ; 
        RECT 27.596 137.214 27.7 141.588 ; 
        RECT 27.164 137.214 27.268 141.588 ; 
        RECT 26.732 137.214 26.836 141.588 ; 
        RECT 26.3 137.214 26.404 141.588 ; 
        RECT 25.868 137.214 25.972 141.588 ; 
        RECT 25.436 137.214 25.54 141.588 ; 
        RECT 25.004 137.214 25.108 141.588 ; 
        RECT 24.572 137.214 24.676 141.588 ; 
        RECT 24.14 137.214 24.244 141.588 ; 
        RECT 23.708 137.214 23.812 141.588 ; 
        RECT 22.856 137.214 23.164 141.588 ; 
        RECT 15.284 137.214 15.592 141.588 ; 
        RECT 14.636 137.214 14.74 141.588 ; 
        RECT 14.204 137.214 14.308 141.588 ; 
        RECT 13.772 137.214 13.876 141.588 ; 
        RECT 13.34 137.214 13.444 141.588 ; 
        RECT 12.908 137.214 13.012 141.588 ; 
        RECT 12.476 137.214 12.58 141.588 ; 
        RECT 12.044 137.214 12.148 141.588 ; 
        RECT 11.612 137.214 11.716 141.588 ; 
        RECT 11.18 137.214 11.284 141.588 ; 
        RECT 10.748 137.214 10.852 141.588 ; 
        RECT 10.316 137.214 10.42 141.588 ; 
        RECT 9.884 137.214 9.988 141.588 ; 
        RECT 9.452 137.214 9.556 141.588 ; 
        RECT 9.02 137.214 9.124 141.588 ; 
        RECT 8.588 137.214 8.692 141.588 ; 
        RECT 8.156 137.214 8.26 141.588 ; 
        RECT 7.724 137.214 7.828 141.588 ; 
        RECT 7.292 137.214 7.396 141.588 ; 
        RECT 6.86 137.214 6.964 141.588 ; 
        RECT 6.428 137.214 6.532 141.588 ; 
        RECT 5.996 137.214 6.1 141.588 ; 
        RECT 5.564 137.214 5.668 141.588 ; 
        RECT 5.132 137.214 5.236 141.588 ; 
        RECT 4.7 137.214 4.804 141.588 ; 
        RECT 4.268 137.214 4.372 141.588 ; 
        RECT 3.836 137.214 3.94 141.588 ; 
        RECT 3.404 137.214 3.508 141.588 ; 
        RECT 2.972 137.214 3.076 141.588 ; 
        RECT 2.54 137.214 2.644 141.588 ; 
        RECT 2.108 137.214 2.212 141.588 ; 
        RECT 1.676 137.214 1.78 141.588 ; 
        RECT 1.244 137.214 1.348 141.588 ; 
        RECT 0.812 137.214 0.916 141.588 ; 
        RECT 0 137.214 0.34 141.588 ; 
        RECT 20.72 141.534 21.232 145.908 ; 
        RECT 20.664 144.196 21.232 145.486 ; 
        RECT 20.072 143.104 20.32 145.908 ; 
        RECT 20.016 144.342 20.32 144.956 ; 
        RECT 20.072 141.534 20.176 145.908 ; 
        RECT 20.072 142.018 20.232 142.976 ; 
        RECT 20.072 141.534 20.32 141.89 ; 
        RECT 18.884 143.336 19.708 145.908 ; 
        RECT 19.604 141.534 19.708 145.908 ; 
        RECT 18.884 144.444 19.764 145.476 ; 
        RECT 18.884 141.534 19.276 145.908 ; 
        RECT 17.216 141.534 17.548 145.908 ; 
        RECT 17.216 141.888 17.604 145.63 ; 
        RECT 38.108 141.534 38.448 145.908 ; 
        RECT 37.532 141.534 37.636 145.908 ; 
        RECT 37.1 141.534 37.204 145.908 ; 
        RECT 36.668 141.534 36.772 145.908 ; 
        RECT 36.236 141.534 36.34 145.908 ; 
        RECT 35.804 141.534 35.908 145.908 ; 
        RECT 35.372 141.534 35.476 145.908 ; 
        RECT 34.94 141.534 35.044 145.908 ; 
        RECT 34.508 141.534 34.612 145.908 ; 
        RECT 34.076 141.534 34.18 145.908 ; 
        RECT 33.644 141.534 33.748 145.908 ; 
        RECT 33.212 141.534 33.316 145.908 ; 
        RECT 32.78 141.534 32.884 145.908 ; 
        RECT 32.348 141.534 32.452 145.908 ; 
        RECT 31.916 141.534 32.02 145.908 ; 
        RECT 31.484 141.534 31.588 145.908 ; 
        RECT 31.052 141.534 31.156 145.908 ; 
        RECT 30.62 141.534 30.724 145.908 ; 
        RECT 30.188 141.534 30.292 145.908 ; 
        RECT 29.756 141.534 29.86 145.908 ; 
        RECT 29.324 141.534 29.428 145.908 ; 
        RECT 28.892 141.534 28.996 145.908 ; 
        RECT 28.46 141.534 28.564 145.908 ; 
        RECT 28.028 141.534 28.132 145.908 ; 
        RECT 27.596 141.534 27.7 145.908 ; 
        RECT 27.164 141.534 27.268 145.908 ; 
        RECT 26.732 141.534 26.836 145.908 ; 
        RECT 26.3 141.534 26.404 145.908 ; 
        RECT 25.868 141.534 25.972 145.908 ; 
        RECT 25.436 141.534 25.54 145.908 ; 
        RECT 25.004 141.534 25.108 145.908 ; 
        RECT 24.572 141.534 24.676 145.908 ; 
        RECT 24.14 141.534 24.244 145.908 ; 
        RECT 23.708 141.534 23.812 145.908 ; 
        RECT 22.856 141.534 23.164 145.908 ; 
        RECT 15.284 141.534 15.592 145.908 ; 
        RECT 14.636 141.534 14.74 145.908 ; 
        RECT 14.204 141.534 14.308 145.908 ; 
        RECT 13.772 141.534 13.876 145.908 ; 
        RECT 13.34 141.534 13.444 145.908 ; 
        RECT 12.908 141.534 13.012 145.908 ; 
        RECT 12.476 141.534 12.58 145.908 ; 
        RECT 12.044 141.534 12.148 145.908 ; 
        RECT 11.612 141.534 11.716 145.908 ; 
        RECT 11.18 141.534 11.284 145.908 ; 
        RECT 10.748 141.534 10.852 145.908 ; 
        RECT 10.316 141.534 10.42 145.908 ; 
        RECT 9.884 141.534 9.988 145.908 ; 
        RECT 9.452 141.534 9.556 145.908 ; 
        RECT 9.02 141.534 9.124 145.908 ; 
        RECT 8.588 141.534 8.692 145.908 ; 
        RECT 8.156 141.534 8.26 145.908 ; 
        RECT 7.724 141.534 7.828 145.908 ; 
        RECT 7.292 141.534 7.396 145.908 ; 
        RECT 6.86 141.534 6.964 145.908 ; 
        RECT 6.428 141.534 6.532 145.908 ; 
        RECT 5.996 141.534 6.1 145.908 ; 
        RECT 5.564 141.534 5.668 145.908 ; 
        RECT 5.132 141.534 5.236 145.908 ; 
        RECT 4.7 141.534 4.804 145.908 ; 
        RECT 4.268 141.534 4.372 145.908 ; 
        RECT 3.836 141.534 3.94 145.908 ; 
        RECT 3.404 141.534 3.508 145.908 ; 
        RECT 2.972 141.534 3.076 145.908 ; 
        RECT 2.54 141.534 2.644 145.908 ; 
        RECT 2.108 141.534 2.212 145.908 ; 
        RECT 1.676 141.534 1.78 145.908 ; 
        RECT 1.244 141.534 1.348 145.908 ; 
        RECT 0.812 141.534 0.916 145.908 ; 
        RECT 0 141.534 0.34 145.908 ; 
        RECT 20.72 145.854 21.232 150.228 ; 
        RECT 20.664 148.516 21.232 149.806 ; 
        RECT 20.072 147.424 20.32 150.228 ; 
        RECT 20.016 148.662 20.32 149.276 ; 
        RECT 20.072 145.854 20.176 150.228 ; 
        RECT 20.072 146.338 20.232 147.296 ; 
        RECT 20.072 145.854 20.32 146.21 ; 
        RECT 18.884 147.656 19.708 150.228 ; 
        RECT 19.604 145.854 19.708 150.228 ; 
        RECT 18.884 148.764 19.764 149.796 ; 
        RECT 18.884 145.854 19.276 150.228 ; 
        RECT 17.216 145.854 17.548 150.228 ; 
        RECT 17.216 146.208 17.604 149.95 ; 
        RECT 38.108 145.854 38.448 150.228 ; 
        RECT 37.532 145.854 37.636 150.228 ; 
        RECT 37.1 145.854 37.204 150.228 ; 
        RECT 36.668 145.854 36.772 150.228 ; 
        RECT 36.236 145.854 36.34 150.228 ; 
        RECT 35.804 145.854 35.908 150.228 ; 
        RECT 35.372 145.854 35.476 150.228 ; 
        RECT 34.94 145.854 35.044 150.228 ; 
        RECT 34.508 145.854 34.612 150.228 ; 
        RECT 34.076 145.854 34.18 150.228 ; 
        RECT 33.644 145.854 33.748 150.228 ; 
        RECT 33.212 145.854 33.316 150.228 ; 
        RECT 32.78 145.854 32.884 150.228 ; 
        RECT 32.348 145.854 32.452 150.228 ; 
        RECT 31.916 145.854 32.02 150.228 ; 
        RECT 31.484 145.854 31.588 150.228 ; 
        RECT 31.052 145.854 31.156 150.228 ; 
        RECT 30.62 145.854 30.724 150.228 ; 
        RECT 30.188 145.854 30.292 150.228 ; 
        RECT 29.756 145.854 29.86 150.228 ; 
        RECT 29.324 145.854 29.428 150.228 ; 
        RECT 28.892 145.854 28.996 150.228 ; 
        RECT 28.46 145.854 28.564 150.228 ; 
        RECT 28.028 145.854 28.132 150.228 ; 
        RECT 27.596 145.854 27.7 150.228 ; 
        RECT 27.164 145.854 27.268 150.228 ; 
        RECT 26.732 145.854 26.836 150.228 ; 
        RECT 26.3 145.854 26.404 150.228 ; 
        RECT 25.868 145.854 25.972 150.228 ; 
        RECT 25.436 145.854 25.54 150.228 ; 
        RECT 25.004 145.854 25.108 150.228 ; 
        RECT 24.572 145.854 24.676 150.228 ; 
        RECT 24.14 145.854 24.244 150.228 ; 
        RECT 23.708 145.854 23.812 150.228 ; 
        RECT 22.856 145.854 23.164 150.228 ; 
        RECT 15.284 145.854 15.592 150.228 ; 
        RECT 14.636 145.854 14.74 150.228 ; 
        RECT 14.204 145.854 14.308 150.228 ; 
        RECT 13.772 145.854 13.876 150.228 ; 
        RECT 13.34 145.854 13.444 150.228 ; 
        RECT 12.908 145.854 13.012 150.228 ; 
        RECT 12.476 145.854 12.58 150.228 ; 
        RECT 12.044 145.854 12.148 150.228 ; 
        RECT 11.612 145.854 11.716 150.228 ; 
        RECT 11.18 145.854 11.284 150.228 ; 
        RECT 10.748 145.854 10.852 150.228 ; 
        RECT 10.316 145.854 10.42 150.228 ; 
        RECT 9.884 145.854 9.988 150.228 ; 
        RECT 9.452 145.854 9.556 150.228 ; 
        RECT 9.02 145.854 9.124 150.228 ; 
        RECT 8.588 145.854 8.692 150.228 ; 
        RECT 8.156 145.854 8.26 150.228 ; 
        RECT 7.724 145.854 7.828 150.228 ; 
        RECT 7.292 145.854 7.396 150.228 ; 
        RECT 6.86 145.854 6.964 150.228 ; 
        RECT 6.428 145.854 6.532 150.228 ; 
        RECT 5.996 145.854 6.1 150.228 ; 
        RECT 5.564 145.854 5.668 150.228 ; 
        RECT 5.132 145.854 5.236 150.228 ; 
        RECT 4.7 145.854 4.804 150.228 ; 
        RECT 4.268 145.854 4.372 150.228 ; 
        RECT 3.836 145.854 3.94 150.228 ; 
        RECT 3.404 145.854 3.508 150.228 ; 
        RECT 2.972 145.854 3.076 150.228 ; 
        RECT 2.54 145.854 2.644 150.228 ; 
        RECT 2.108 145.854 2.212 150.228 ; 
        RECT 1.676 145.854 1.78 150.228 ; 
        RECT 1.244 145.854 1.348 150.228 ; 
        RECT 0.812 145.854 0.916 150.228 ; 
        RECT 0 145.854 0.34 150.228 ; 
        RECT 20.72 150.174 21.232 154.548 ; 
        RECT 20.664 152.836 21.232 154.126 ; 
        RECT 20.072 151.744 20.32 154.548 ; 
        RECT 20.016 152.982 20.32 153.596 ; 
        RECT 20.072 150.174 20.176 154.548 ; 
        RECT 20.072 150.658 20.232 151.616 ; 
        RECT 20.072 150.174 20.32 150.53 ; 
        RECT 18.884 151.976 19.708 154.548 ; 
        RECT 19.604 150.174 19.708 154.548 ; 
        RECT 18.884 153.084 19.764 154.116 ; 
        RECT 18.884 150.174 19.276 154.548 ; 
        RECT 17.216 150.174 17.548 154.548 ; 
        RECT 17.216 150.528 17.604 154.27 ; 
        RECT 38.108 150.174 38.448 154.548 ; 
        RECT 37.532 150.174 37.636 154.548 ; 
        RECT 37.1 150.174 37.204 154.548 ; 
        RECT 36.668 150.174 36.772 154.548 ; 
        RECT 36.236 150.174 36.34 154.548 ; 
        RECT 35.804 150.174 35.908 154.548 ; 
        RECT 35.372 150.174 35.476 154.548 ; 
        RECT 34.94 150.174 35.044 154.548 ; 
        RECT 34.508 150.174 34.612 154.548 ; 
        RECT 34.076 150.174 34.18 154.548 ; 
        RECT 33.644 150.174 33.748 154.548 ; 
        RECT 33.212 150.174 33.316 154.548 ; 
        RECT 32.78 150.174 32.884 154.548 ; 
        RECT 32.348 150.174 32.452 154.548 ; 
        RECT 31.916 150.174 32.02 154.548 ; 
        RECT 31.484 150.174 31.588 154.548 ; 
        RECT 31.052 150.174 31.156 154.548 ; 
        RECT 30.62 150.174 30.724 154.548 ; 
        RECT 30.188 150.174 30.292 154.548 ; 
        RECT 29.756 150.174 29.86 154.548 ; 
        RECT 29.324 150.174 29.428 154.548 ; 
        RECT 28.892 150.174 28.996 154.548 ; 
        RECT 28.46 150.174 28.564 154.548 ; 
        RECT 28.028 150.174 28.132 154.548 ; 
        RECT 27.596 150.174 27.7 154.548 ; 
        RECT 27.164 150.174 27.268 154.548 ; 
        RECT 26.732 150.174 26.836 154.548 ; 
        RECT 26.3 150.174 26.404 154.548 ; 
        RECT 25.868 150.174 25.972 154.548 ; 
        RECT 25.436 150.174 25.54 154.548 ; 
        RECT 25.004 150.174 25.108 154.548 ; 
        RECT 24.572 150.174 24.676 154.548 ; 
        RECT 24.14 150.174 24.244 154.548 ; 
        RECT 23.708 150.174 23.812 154.548 ; 
        RECT 22.856 150.174 23.164 154.548 ; 
        RECT 15.284 150.174 15.592 154.548 ; 
        RECT 14.636 150.174 14.74 154.548 ; 
        RECT 14.204 150.174 14.308 154.548 ; 
        RECT 13.772 150.174 13.876 154.548 ; 
        RECT 13.34 150.174 13.444 154.548 ; 
        RECT 12.908 150.174 13.012 154.548 ; 
        RECT 12.476 150.174 12.58 154.548 ; 
        RECT 12.044 150.174 12.148 154.548 ; 
        RECT 11.612 150.174 11.716 154.548 ; 
        RECT 11.18 150.174 11.284 154.548 ; 
        RECT 10.748 150.174 10.852 154.548 ; 
        RECT 10.316 150.174 10.42 154.548 ; 
        RECT 9.884 150.174 9.988 154.548 ; 
        RECT 9.452 150.174 9.556 154.548 ; 
        RECT 9.02 150.174 9.124 154.548 ; 
        RECT 8.588 150.174 8.692 154.548 ; 
        RECT 8.156 150.174 8.26 154.548 ; 
        RECT 7.724 150.174 7.828 154.548 ; 
        RECT 7.292 150.174 7.396 154.548 ; 
        RECT 6.86 150.174 6.964 154.548 ; 
        RECT 6.428 150.174 6.532 154.548 ; 
        RECT 5.996 150.174 6.1 154.548 ; 
        RECT 5.564 150.174 5.668 154.548 ; 
        RECT 5.132 150.174 5.236 154.548 ; 
        RECT 4.7 150.174 4.804 154.548 ; 
        RECT 4.268 150.174 4.372 154.548 ; 
        RECT 3.836 150.174 3.94 154.548 ; 
        RECT 3.404 150.174 3.508 154.548 ; 
        RECT 2.972 150.174 3.076 154.548 ; 
        RECT 2.54 150.174 2.644 154.548 ; 
        RECT 2.108 150.174 2.212 154.548 ; 
        RECT 1.676 150.174 1.78 154.548 ; 
        RECT 1.244 150.174 1.348 154.548 ; 
        RECT 0.812 150.174 0.916 154.548 ; 
        RECT 0 150.174 0.34 154.548 ; 
        RECT 20.72 154.494 21.232 158.868 ; 
        RECT 20.664 157.156 21.232 158.446 ; 
        RECT 20.072 156.064 20.32 158.868 ; 
        RECT 20.016 157.302 20.32 157.916 ; 
        RECT 20.072 154.494 20.176 158.868 ; 
        RECT 20.072 154.978 20.232 155.936 ; 
        RECT 20.072 154.494 20.32 154.85 ; 
        RECT 18.884 156.296 19.708 158.868 ; 
        RECT 19.604 154.494 19.708 158.868 ; 
        RECT 18.884 157.404 19.764 158.436 ; 
        RECT 18.884 154.494 19.276 158.868 ; 
        RECT 17.216 154.494 17.548 158.868 ; 
        RECT 17.216 154.848 17.604 158.59 ; 
        RECT 38.108 154.494 38.448 158.868 ; 
        RECT 37.532 154.494 37.636 158.868 ; 
        RECT 37.1 154.494 37.204 158.868 ; 
        RECT 36.668 154.494 36.772 158.868 ; 
        RECT 36.236 154.494 36.34 158.868 ; 
        RECT 35.804 154.494 35.908 158.868 ; 
        RECT 35.372 154.494 35.476 158.868 ; 
        RECT 34.94 154.494 35.044 158.868 ; 
        RECT 34.508 154.494 34.612 158.868 ; 
        RECT 34.076 154.494 34.18 158.868 ; 
        RECT 33.644 154.494 33.748 158.868 ; 
        RECT 33.212 154.494 33.316 158.868 ; 
        RECT 32.78 154.494 32.884 158.868 ; 
        RECT 32.348 154.494 32.452 158.868 ; 
        RECT 31.916 154.494 32.02 158.868 ; 
        RECT 31.484 154.494 31.588 158.868 ; 
        RECT 31.052 154.494 31.156 158.868 ; 
        RECT 30.62 154.494 30.724 158.868 ; 
        RECT 30.188 154.494 30.292 158.868 ; 
        RECT 29.756 154.494 29.86 158.868 ; 
        RECT 29.324 154.494 29.428 158.868 ; 
        RECT 28.892 154.494 28.996 158.868 ; 
        RECT 28.46 154.494 28.564 158.868 ; 
        RECT 28.028 154.494 28.132 158.868 ; 
        RECT 27.596 154.494 27.7 158.868 ; 
        RECT 27.164 154.494 27.268 158.868 ; 
        RECT 26.732 154.494 26.836 158.868 ; 
        RECT 26.3 154.494 26.404 158.868 ; 
        RECT 25.868 154.494 25.972 158.868 ; 
        RECT 25.436 154.494 25.54 158.868 ; 
        RECT 25.004 154.494 25.108 158.868 ; 
        RECT 24.572 154.494 24.676 158.868 ; 
        RECT 24.14 154.494 24.244 158.868 ; 
        RECT 23.708 154.494 23.812 158.868 ; 
        RECT 22.856 154.494 23.164 158.868 ; 
        RECT 15.284 154.494 15.592 158.868 ; 
        RECT 14.636 154.494 14.74 158.868 ; 
        RECT 14.204 154.494 14.308 158.868 ; 
        RECT 13.772 154.494 13.876 158.868 ; 
        RECT 13.34 154.494 13.444 158.868 ; 
        RECT 12.908 154.494 13.012 158.868 ; 
        RECT 12.476 154.494 12.58 158.868 ; 
        RECT 12.044 154.494 12.148 158.868 ; 
        RECT 11.612 154.494 11.716 158.868 ; 
        RECT 11.18 154.494 11.284 158.868 ; 
        RECT 10.748 154.494 10.852 158.868 ; 
        RECT 10.316 154.494 10.42 158.868 ; 
        RECT 9.884 154.494 9.988 158.868 ; 
        RECT 9.452 154.494 9.556 158.868 ; 
        RECT 9.02 154.494 9.124 158.868 ; 
        RECT 8.588 154.494 8.692 158.868 ; 
        RECT 8.156 154.494 8.26 158.868 ; 
        RECT 7.724 154.494 7.828 158.868 ; 
        RECT 7.292 154.494 7.396 158.868 ; 
        RECT 6.86 154.494 6.964 158.868 ; 
        RECT 6.428 154.494 6.532 158.868 ; 
        RECT 5.996 154.494 6.1 158.868 ; 
        RECT 5.564 154.494 5.668 158.868 ; 
        RECT 5.132 154.494 5.236 158.868 ; 
        RECT 4.7 154.494 4.804 158.868 ; 
        RECT 4.268 154.494 4.372 158.868 ; 
        RECT 3.836 154.494 3.94 158.868 ; 
        RECT 3.404 154.494 3.508 158.868 ; 
        RECT 2.972 154.494 3.076 158.868 ; 
        RECT 2.54 154.494 2.644 158.868 ; 
        RECT 2.108 154.494 2.212 158.868 ; 
        RECT 1.676 154.494 1.78 158.868 ; 
        RECT 1.244 154.494 1.348 158.868 ; 
        RECT 0.812 154.494 0.916 158.868 ; 
        RECT 0 154.494 0.34 158.868 ; 
        RECT 20.72 158.814 21.232 163.188 ; 
        RECT 20.664 161.476 21.232 162.766 ; 
        RECT 20.072 160.384 20.32 163.188 ; 
        RECT 20.016 161.622 20.32 162.236 ; 
        RECT 20.072 158.814 20.176 163.188 ; 
        RECT 20.072 159.298 20.232 160.256 ; 
        RECT 20.072 158.814 20.32 159.17 ; 
        RECT 18.884 160.616 19.708 163.188 ; 
        RECT 19.604 158.814 19.708 163.188 ; 
        RECT 18.884 161.724 19.764 162.756 ; 
        RECT 18.884 158.814 19.276 163.188 ; 
        RECT 17.216 158.814 17.548 163.188 ; 
        RECT 17.216 159.168 17.604 162.91 ; 
        RECT 38.108 158.814 38.448 163.188 ; 
        RECT 37.532 158.814 37.636 163.188 ; 
        RECT 37.1 158.814 37.204 163.188 ; 
        RECT 36.668 158.814 36.772 163.188 ; 
        RECT 36.236 158.814 36.34 163.188 ; 
        RECT 35.804 158.814 35.908 163.188 ; 
        RECT 35.372 158.814 35.476 163.188 ; 
        RECT 34.94 158.814 35.044 163.188 ; 
        RECT 34.508 158.814 34.612 163.188 ; 
        RECT 34.076 158.814 34.18 163.188 ; 
        RECT 33.644 158.814 33.748 163.188 ; 
        RECT 33.212 158.814 33.316 163.188 ; 
        RECT 32.78 158.814 32.884 163.188 ; 
        RECT 32.348 158.814 32.452 163.188 ; 
        RECT 31.916 158.814 32.02 163.188 ; 
        RECT 31.484 158.814 31.588 163.188 ; 
        RECT 31.052 158.814 31.156 163.188 ; 
        RECT 30.62 158.814 30.724 163.188 ; 
        RECT 30.188 158.814 30.292 163.188 ; 
        RECT 29.756 158.814 29.86 163.188 ; 
        RECT 29.324 158.814 29.428 163.188 ; 
        RECT 28.892 158.814 28.996 163.188 ; 
        RECT 28.46 158.814 28.564 163.188 ; 
        RECT 28.028 158.814 28.132 163.188 ; 
        RECT 27.596 158.814 27.7 163.188 ; 
        RECT 27.164 158.814 27.268 163.188 ; 
        RECT 26.732 158.814 26.836 163.188 ; 
        RECT 26.3 158.814 26.404 163.188 ; 
        RECT 25.868 158.814 25.972 163.188 ; 
        RECT 25.436 158.814 25.54 163.188 ; 
        RECT 25.004 158.814 25.108 163.188 ; 
        RECT 24.572 158.814 24.676 163.188 ; 
        RECT 24.14 158.814 24.244 163.188 ; 
        RECT 23.708 158.814 23.812 163.188 ; 
        RECT 22.856 158.814 23.164 163.188 ; 
        RECT 15.284 158.814 15.592 163.188 ; 
        RECT 14.636 158.814 14.74 163.188 ; 
        RECT 14.204 158.814 14.308 163.188 ; 
        RECT 13.772 158.814 13.876 163.188 ; 
        RECT 13.34 158.814 13.444 163.188 ; 
        RECT 12.908 158.814 13.012 163.188 ; 
        RECT 12.476 158.814 12.58 163.188 ; 
        RECT 12.044 158.814 12.148 163.188 ; 
        RECT 11.612 158.814 11.716 163.188 ; 
        RECT 11.18 158.814 11.284 163.188 ; 
        RECT 10.748 158.814 10.852 163.188 ; 
        RECT 10.316 158.814 10.42 163.188 ; 
        RECT 9.884 158.814 9.988 163.188 ; 
        RECT 9.452 158.814 9.556 163.188 ; 
        RECT 9.02 158.814 9.124 163.188 ; 
        RECT 8.588 158.814 8.692 163.188 ; 
        RECT 8.156 158.814 8.26 163.188 ; 
        RECT 7.724 158.814 7.828 163.188 ; 
        RECT 7.292 158.814 7.396 163.188 ; 
        RECT 6.86 158.814 6.964 163.188 ; 
        RECT 6.428 158.814 6.532 163.188 ; 
        RECT 5.996 158.814 6.1 163.188 ; 
        RECT 5.564 158.814 5.668 163.188 ; 
        RECT 5.132 158.814 5.236 163.188 ; 
        RECT 4.7 158.814 4.804 163.188 ; 
        RECT 4.268 158.814 4.372 163.188 ; 
        RECT 3.836 158.814 3.94 163.188 ; 
        RECT 3.404 158.814 3.508 163.188 ; 
        RECT 2.972 158.814 3.076 163.188 ; 
        RECT 2.54 158.814 2.644 163.188 ; 
        RECT 2.108 158.814 2.212 163.188 ; 
        RECT 1.676 158.814 1.78 163.188 ; 
        RECT 1.244 158.814 1.348 163.188 ; 
        RECT 0.812 158.814 0.916 163.188 ; 
        RECT 0 158.814 0.34 163.188 ; 
        RECT 20.72 163.134 21.232 167.508 ; 
        RECT 20.664 165.796 21.232 167.086 ; 
        RECT 20.072 164.704 20.32 167.508 ; 
        RECT 20.016 165.942 20.32 166.556 ; 
        RECT 20.072 163.134 20.176 167.508 ; 
        RECT 20.072 163.618 20.232 164.576 ; 
        RECT 20.072 163.134 20.32 163.49 ; 
        RECT 18.884 164.936 19.708 167.508 ; 
        RECT 19.604 163.134 19.708 167.508 ; 
        RECT 18.884 166.044 19.764 167.076 ; 
        RECT 18.884 163.134 19.276 167.508 ; 
        RECT 17.216 163.134 17.548 167.508 ; 
        RECT 17.216 163.488 17.604 167.23 ; 
        RECT 38.108 163.134 38.448 167.508 ; 
        RECT 37.532 163.134 37.636 167.508 ; 
        RECT 37.1 163.134 37.204 167.508 ; 
        RECT 36.668 163.134 36.772 167.508 ; 
        RECT 36.236 163.134 36.34 167.508 ; 
        RECT 35.804 163.134 35.908 167.508 ; 
        RECT 35.372 163.134 35.476 167.508 ; 
        RECT 34.94 163.134 35.044 167.508 ; 
        RECT 34.508 163.134 34.612 167.508 ; 
        RECT 34.076 163.134 34.18 167.508 ; 
        RECT 33.644 163.134 33.748 167.508 ; 
        RECT 33.212 163.134 33.316 167.508 ; 
        RECT 32.78 163.134 32.884 167.508 ; 
        RECT 32.348 163.134 32.452 167.508 ; 
        RECT 31.916 163.134 32.02 167.508 ; 
        RECT 31.484 163.134 31.588 167.508 ; 
        RECT 31.052 163.134 31.156 167.508 ; 
        RECT 30.62 163.134 30.724 167.508 ; 
        RECT 30.188 163.134 30.292 167.508 ; 
        RECT 29.756 163.134 29.86 167.508 ; 
        RECT 29.324 163.134 29.428 167.508 ; 
        RECT 28.892 163.134 28.996 167.508 ; 
        RECT 28.46 163.134 28.564 167.508 ; 
        RECT 28.028 163.134 28.132 167.508 ; 
        RECT 27.596 163.134 27.7 167.508 ; 
        RECT 27.164 163.134 27.268 167.508 ; 
        RECT 26.732 163.134 26.836 167.508 ; 
        RECT 26.3 163.134 26.404 167.508 ; 
        RECT 25.868 163.134 25.972 167.508 ; 
        RECT 25.436 163.134 25.54 167.508 ; 
        RECT 25.004 163.134 25.108 167.508 ; 
        RECT 24.572 163.134 24.676 167.508 ; 
        RECT 24.14 163.134 24.244 167.508 ; 
        RECT 23.708 163.134 23.812 167.508 ; 
        RECT 22.856 163.134 23.164 167.508 ; 
        RECT 15.284 163.134 15.592 167.508 ; 
        RECT 14.636 163.134 14.74 167.508 ; 
        RECT 14.204 163.134 14.308 167.508 ; 
        RECT 13.772 163.134 13.876 167.508 ; 
        RECT 13.34 163.134 13.444 167.508 ; 
        RECT 12.908 163.134 13.012 167.508 ; 
        RECT 12.476 163.134 12.58 167.508 ; 
        RECT 12.044 163.134 12.148 167.508 ; 
        RECT 11.612 163.134 11.716 167.508 ; 
        RECT 11.18 163.134 11.284 167.508 ; 
        RECT 10.748 163.134 10.852 167.508 ; 
        RECT 10.316 163.134 10.42 167.508 ; 
        RECT 9.884 163.134 9.988 167.508 ; 
        RECT 9.452 163.134 9.556 167.508 ; 
        RECT 9.02 163.134 9.124 167.508 ; 
        RECT 8.588 163.134 8.692 167.508 ; 
        RECT 8.156 163.134 8.26 167.508 ; 
        RECT 7.724 163.134 7.828 167.508 ; 
        RECT 7.292 163.134 7.396 167.508 ; 
        RECT 6.86 163.134 6.964 167.508 ; 
        RECT 6.428 163.134 6.532 167.508 ; 
        RECT 5.996 163.134 6.1 167.508 ; 
        RECT 5.564 163.134 5.668 167.508 ; 
        RECT 5.132 163.134 5.236 167.508 ; 
        RECT 4.7 163.134 4.804 167.508 ; 
        RECT 4.268 163.134 4.372 167.508 ; 
        RECT 3.836 163.134 3.94 167.508 ; 
        RECT 3.404 163.134 3.508 167.508 ; 
        RECT 2.972 163.134 3.076 167.508 ; 
        RECT 2.54 163.134 2.644 167.508 ; 
        RECT 2.108 163.134 2.212 167.508 ; 
        RECT 1.676 163.134 1.78 167.508 ; 
        RECT 1.244 163.134 1.348 167.508 ; 
        RECT 0.812 163.134 0.916 167.508 ; 
        RECT 0 163.134 0.34 167.508 ; 
        RECT 20.72 167.454 21.232 171.828 ; 
        RECT 20.664 170.116 21.232 171.406 ; 
        RECT 20.072 169.024 20.32 171.828 ; 
        RECT 20.016 170.262 20.32 170.876 ; 
        RECT 20.072 167.454 20.176 171.828 ; 
        RECT 20.072 167.938 20.232 168.896 ; 
        RECT 20.072 167.454 20.32 167.81 ; 
        RECT 18.884 169.256 19.708 171.828 ; 
        RECT 19.604 167.454 19.708 171.828 ; 
        RECT 18.884 170.364 19.764 171.396 ; 
        RECT 18.884 167.454 19.276 171.828 ; 
        RECT 17.216 167.454 17.548 171.828 ; 
        RECT 17.216 167.808 17.604 171.55 ; 
        RECT 38.108 167.454 38.448 171.828 ; 
        RECT 37.532 167.454 37.636 171.828 ; 
        RECT 37.1 167.454 37.204 171.828 ; 
        RECT 36.668 167.454 36.772 171.828 ; 
        RECT 36.236 167.454 36.34 171.828 ; 
        RECT 35.804 167.454 35.908 171.828 ; 
        RECT 35.372 167.454 35.476 171.828 ; 
        RECT 34.94 167.454 35.044 171.828 ; 
        RECT 34.508 167.454 34.612 171.828 ; 
        RECT 34.076 167.454 34.18 171.828 ; 
        RECT 33.644 167.454 33.748 171.828 ; 
        RECT 33.212 167.454 33.316 171.828 ; 
        RECT 32.78 167.454 32.884 171.828 ; 
        RECT 32.348 167.454 32.452 171.828 ; 
        RECT 31.916 167.454 32.02 171.828 ; 
        RECT 31.484 167.454 31.588 171.828 ; 
        RECT 31.052 167.454 31.156 171.828 ; 
        RECT 30.62 167.454 30.724 171.828 ; 
        RECT 30.188 167.454 30.292 171.828 ; 
        RECT 29.756 167.454 29.86 171.828 ; 
        RECT 29.324 167.454 29.428 171.828 ; 
        RECT 28.892 167.454 28.996 171.828 ; 
        RECT 28.46 167.454 28.564 171.828 ; 
        RECT 28.028 167.454 28.132 171.828 ; 
        RECT 27.596 167.454 27.7 171.828 ; 
        RECT 27.164 167.454 27.268 171.828 ; 
        RECT 26.732 167.454 26.836 171.828 ; 
        RECT 26.3 167.454 26.404 171.828 ; 
        RECT 25.868 167.454 25.972 171.828 ; 
        RECT 25.436 167.454 25.54 171.828 ; 
        RECT 25.004 167.454 25.108 171.828 ; 
        RECT 24.572 167.454 24.676 171.828 ; 
        RECT 24.14 167.454 24.244 171.828 ; 
        RECT 23.708 167.454 23.812 171.828 ; 
        RECT 22.856 167.454 23.164 171.828 ; 
        RECT 15.284 167.454 15.592 171.828 ; 
        RECT 14.636 167.454 14.74 171.828 ; 
        RECT 14.204 167.454 14.308 171.828 ; 
        RECT 13.772 167.454 13.876 171.828 ; 
        RECT 13.34 167.454 13.444 171.828 ; 
        RECT 12.908 167.454 13.012 171.828 ; 
        RECT 12.476 167.454 12.58 171.828 ; 
        RECT 12.044 167.454 12.148 171.828 ; 
        RECT 11.612 167.454 11.716 171.828 ; 
        RECT 11.18 167.454 11.284 171.828 ; 
        RECT 10.748 167.454 10.852 171.828 ; 
        RECT 10.316 167.454 10.42 171.828 ; 
        RECT 9.884 167.454 9.988 171.828 ; 
        RECT 9.452 167.454 9.556 171.828 ; 
        RECT 9.02 167.454 9.124 171.828 ; 
        RECT 8.588 167.454 8.692 171.828 ; 
        RECT 8.156 167.454 8.26 171.828 ; 
        RECT 7.724 167.454 7.828 171.828 ; 
        RECT 7.292 167.454 7.396 171.828 ; 
        RECT 6.86 167.454 6.964 171.828 ; 
        RECT 6.428 167.454 6.532 171.828 ; 
        RECT 5.996 167.454 6.1 171.828 ; 
        RECT 5.564 167.454 5.668 171.828 ; 
        RECT 5.132 167.454 5.236 171.828 ; 
        RECT 4.7 167.454 4.804 171.828 ; 
        RECT 4.268 167.454 4.372 171.828 ; 
        RECT 3.836 167.454 3.94 171.828 ; 
        RECT 3.404 167.454 3.508 171.828 ; 
        RECT 2.972 167.454 3.076 171.828 ; 
        RECT 2.54 167.454 2.644 171.828 ; 
        RECT 2.108 167.454 2.212 171.828 ; 
        RECT 1.676 167.454 1.78 171.828 ; 
        RECT 1.244 167.454 1.348 171.828 ; 
        RECT 0.812 167.454 0.916 171.828 ; 
        RECT 0 167.454 0.34 171.828 ; 
        RECT 20.72 171.774 21.232 176.148 ; 
        RECT 20.664 174.436 21.232 175.726 ; 
        RECT 20.072 173.344 20.32 176.148 ; 
        RECT 20.016 174.582 20.32 175.196 ; 
        RECT 20.072 171.774 20.176 176.148 ; 
        RECT 20.072 172.258 20.232 173.216 ; 
        RECT 20.072 171.774 20.32 172.13 ; 
        RECT 18.884 173.576 19.708 176.148 ; 
        RECT 19.604 171.774 19.708 176.148 ; 
        RECT 18.884 174.684 19.764 175.716 ; 
        RECT 18.884 171.774 19.276 176.148 ; 
        RECT 17.216 171.774 17.548 176.148 ; 
        RECT 17.216 172.128 17.604 175.87 ; 
        RECT 38.108 171.774 38.448 176.148 ; 
        RECT 37.532 171.774 37.636 176.148 ; 
        RECT 37.1 171.774 37.204 176.148 ; 
        RECT 36.668 171.774 36.772 176.148 ; 
        RECT 36.236 171.774 36.34 176.148 ; 
        RECT 35.804 171.774 35.908 176.148 ; 
        RECT 35.372 171.774 35.476 176.148 ; 
        RECT 34.94 171.774 35.044 176.148 ; 
        RECT 34.508 171.774 34.612 176.148 ; 
        RECT 34.076 171.774 34.18 176.148 ; 
        RECT 33.644 171.774 33.748 176.148 ; 
        RECT 33.212 171.774 33.316 176.148 ; 
        RECT 32.78 171.774 32.884 176.148 ; 
        RECT 32.348 171.774 32.452 176.148 ; 
        RECT 31.916 171.774 32.02 176.148 ; 
        RECT 31.484 171.774 31.588 176.148 ; 
        RECT 31.052 171.774 31.156 176.148 ; 
        RECT 30.62 171.774 30.724 176.148 ; 
        RECT 30.188 171.774 30.292 176.148 ; 
        RECT 29.756 171.774 29.86 176.148 ; 
        RECT 29.324 171.774 29.428 176.148 ; 
        RECT 28.892 171.774 28.996 176.148 ; 
        RECT 28.46 171.774 28.564 176.148 ; 
        RECT 28.028 171.774 28.132 176.148 ; 
        RECT 27.596 171.774 27.7 176.148 ; 
        RECT 27.164 171.774 27.268 176.148 ; 
        RECT 26.732 171.774 26.836 176.148 ; 
        RECT 26.3 171.774 26.404 176.148 ; 
        RECT 25.868 171.774 25.972 176.148 ; 
        RECT 25.436 171.774 25.54 176.148 ; 
        RECT 25.004 171.774 25.108 176.148 ; 
        RECT 24.572 171.774 24.676 176.148 ; 
        RECT 24.14 171.774 24.244 176.148 ; 
        RECT 23.708 171.774 23.812 176.148 ; 
        RECT 22.856 171.774 23.164 176.148 ; 
        RECT 15.284 171.774 15.592 176.148 ; 
        RECT 14.636 171.774 14.74 176.148 ; 
        RECT 14.204 171.774 14.308 176.148 ; 
        RECT 13.772 171.774 13.876 176.148 ; 
        RECT 13.34 171.774 13.444 176.148 ; 
        RECT 12.908 171.774 13.012 176.148 ; 
        RECT 12.476 171.774 12.58 176.148 ; 
        RECT 12.044 171.774 12.148 176.148 ; 
        RECT 11.612 171.774 11.716 176.148 ; 
        RECT 11.18 171.774 11.284 176.148 ; 
        RECT 10.748 171.774 10.852 176.148 ; 
        RECT 10.316 171.774 10.42 176.148 ; 
        RECT 9.884 171.774 9.988 176.148 ; 
        RECT 9.452 171.774 9.556 176.148 ; 
        RECT 9.02 171.774 9.124 176.148 ; 
        RECT 8.588 171.774 8.692 176.148 ; 
        RECT 8.156 171.774 8.26 176.148 ; 
        RECT 7.724 171.774 7.828 176.148 ; 
        RECT 7.292 171.774 7.396 176.148 ; 
        RECT 6.86 171.774 6.964 176.148 ; 
        RECT 6.428 171.774 6.532 176.148 ; 
        RECT 5.996 171.774 6.1 176.148 ; 
        RECT 5.564 171.774 5.668 176.148 ; 
        RECT 5.132 171.774 5.236 176.148 ; 
        RECT 4.7 171.774 4.804 176.148 ; 
        RECT 4.268 171.774 4.372 176.148 ; 
        RECT 3.836 171.774 3.94 176.148 ; 
        RECT 3.404 171.774 3.508 176.148 ; 
        RECT 2.972 171.774 3.076 176.148 ; 
        RECT 2.54 171.774 2.644 176.148 ; 
        RECT 2.108 171.774 2.212 176.148 ; 
        RECT 1.676 171.774 1.78 176.148 ; 
        RECT 1.244 171.774 1.348 176.148 ; 
        RECT 0.812 171.774 0.916 176.148 ; 
        RECT 0 171.774 0.34 176.148 ; 
        RECT 20.72 176.094 21.232 180.468 ; 
        RECT 20.664 178.756 21.232 180.046 ; 
        RECT 20.072 177.664 20.32 180.468 ; 
        RECT 20.016 178.902 20.32 179.516 ; 
        RECT 20.072 176.094 20.176 180.468 ; 
        RECT 20.072 176.578 20.232 177.536 ; 
        RECT 20.072 176.094 20.32 176.45 ; 
        RECT 18.884 177.896 19.708 180.468 ; 
        RECT 19.604 176.094 19.708 180.468 ; 
        RECT 18.884 179.004 19.764 180.036 ; 
        RECT 18.884 176.094 19.276 180.468 ; 
        RECT 17.216 176.094 17.548 180.468 ; 
        RECT 17.216 176.448 17.604 180.19 ; 
        RECT 38.108 176.094 38.448 180.468 ; 
        RECT 37.532 176.094 37.636 180.468 ; 
        RECT 37.1 176.094 37.204 180.468 ; 
        RECT 36.668 176.094 36.772 180.468 ; 
        RECT 36.236 176.094 36.34 180.468 ; 
        RECT 35.804 176.094 35.908 180.468 ; 
        RECT 35.372 176.094 35.476 180.468 ; 
        RECT 34.94 176.094 35.044 180.468 ; 
        RECT 34.508 176.094 34.612 180.468 ; 
        RECT 34.076 176.094 34.18 180.468 ; 
        RECT 33.644 176.094 33.748 180.468 ; 
        RECT 33.212 176.094 33.316 180.468 ; 
        RECT 32.78 176.094 32.884 180.468 ; 
        RECT 32.348 176.094 32.452 180.468 ; 
        RECT 31.916 176.094 32.02 180.468 ; 
        RECT 31.484 176.094 31.588 180.468 ; 
        RECT 31.052 176.094 31.156 180.468 ; 
        RECT 30.62 176.094 30.724 180.468 ; 
        RECT 30.188 176.094 30.292 180.468 ; 
        RECT 29.756 176.094 29.86 180.468 ; 
        RECT 29.324 176.094 29.428 180.468 ; 
        RECT 28.892 176.094 28.996 180.468 ; 
        RECT 28.46 176.094 28.564 180.468 ; 
        RECT 28.028 176.094 28.132 180.468 ; 
        RECT 27.596 176.094 27.7 180.468 ; 
        RECT 27.164 176.094 27.268 180.468 ; 
        RECT 26.732 176.094 26.836 180.468 ; 
        RECT 26.3 176.094 26.404 180.468 ; 
        RECT 25.868 176.094 25.972 180.468 ; 
        RECT 25.436 176.094 25.54 180.468 ; 
        RECT 25.004 176.094 25.108 180.468 ; 
        RECT 24.572 176.094 24.676 180.468 ; 
        RECT 24.14 176.094 24.244 180.468 ; 
        RECT 23.708 176.094 23.812 180.468 ; 
        RECT 22.856 176.094 23.164 180.468 ; 
        RECT 15.284 176.094 15.592 180.468 ; 
        RECT 14.636 176.094 14.74 180.468 ; 
        RECT 14.204 176.094 14.308 180.468 ; 
        RECT 13.772 176.094 13.876 180.468 ; 
        RECT 13.34 176.094 13.444 180.468 ; 
        RECT 12.908 176.094 13.012 180.468 ; 
        RECT 12.476 176.094 12.58 180.468 ; 
        RECT 12.044 176.094 12.148 180.468 ; 
        RECT 11.612 176.094 11.716 180.468 ; 
        RECT 11.18 176.094 11.284 180.468 ; 
        RECT 10.748 176.094 10.852 180.468 ; 
        RECT 10.316 176.094 10.42 180.468 ; 
        RECT 9.884 176.094 9.988 180.468 ; 
        RECT 9.452 176.094 9.556 180.468 ; 
        RECT 9.02 176.094 9.124 180.468 ; 
        RECT 8.588 176.094 8.692 180.468 ; 
        RECT 8.156 176.094 8.26 180.468 ; 
        RECT 7.724 176.094 7.828 180.468 ; 
        RECT 7.292 176.094 7.396 180.468 ; 
        RECT 6.86 176.094 6.964 180.468 ; 
        RECT 6.428 176.094 6.532 180.468 ; 
        RECT 5.996 176.094 6.1 180.468 ; 
        RECT 5.564 176.094 5.668 180.468 ; 
        RECT 5.132 176.094 5.236 180.468 ; 
        RECT 4.7 176.094 4.804 180.468 ; 
        RECT 4.268 176.094 4.372 180.468 ; 
        RECT 3.836 176.094 3.94 180.468 ; 
        RECT 3.404 176.094 3.508 180.468 ; 
        RECT 2.972 176.094 3.076 180.468 ; 
        RECT 2.54 176.094 2.644 180.468 ; 
        RECT 2.108 176.094 2.212 180.468 ; 
        RECT 1.676 176.094 1.78 180.468 ; 
        RECT 1.244 176.094 1.348 180.468 ; 
        RECT 0.812 176.094 0.916 180.468 ; 
        RECT 0 176.094 0.34 180.468 ; 
        RECT 20.72 180.414 21.232 184.788 ; 
        RECT 20.664 183.076 21.232 184.366 ; 
        RECT 20.072 181.984 20.32 184.788 ; 
        RECT 20.016 183.222 20.32 183.836 ; 
        RECT 20.072 180.414 20.176 184.788 ; 
        RECT 20.072 180.898 20.232 181.856 ; 
        RECT 20.072 180.414 20.32 180.77 ; 
        RECT 18.884 182.216 19.708 184.788 ; 
        RECT 19.604 180.414 19.708 184.788 ; 
        RECT 18.884 183.324 19.764 184.356 ; 
        RECT 18.884 180.414 19.276 184.788 ; 
        RECT 17.216 180.414 17.548 184.788 ; 
        RECT 17.216 180.768 17.604 184.51 ; 
        RECT 38.108 180.414 38.448 184.788 ; 
        RECT 37.532 180.414 37.636 184.788 ; 
        RECT 37.1 180.414 37.204 184.788 ; 
        RECT 36.668 180.414 36.772 184.788 ; 
        RECT 36.236 180.414 36.34 184.788 ; 
        RECT 35.804 180.414 35.908 184.788 ; 
        RECT 35.372 180.414 35.476 184.788 ; 
        RECT 34.94 180.414 35.044 184.788 ; 
        RECT 34.508 180.414 34.612 184.788 ; 
        RECT 34.076 180.414 34.18 184.788 ; 
        RECT 33.644 180.414 33.748 184.788 ; 
        RECT 33.212 180.414 33.316 184.788 ; 
        RECT 32.78 180.414 32.884 184.788 ; 
        RECT 32.348 180.414 32.452 184.788 ; 
        RECT 31.916 180.414 32.02 184.788 ; 
        RECT 31.484 180.414 31.588 184.788 ; 
        RECT 31.052 180.414 31.156 184.788 ; 
        RECT 30.62 180.414 30.724 184.788 ; 
        RECT 30.188 180.414 30.292 184.788 ; 
        RECT 29.756 180.414 29.86 184.788 ; 
        RECT 29.324 180.414 29.428 184.788 ; 
        RECT 28.892 180.414 28.996 184.788 ; 
        RECT 28.46 180.414 28.564 184.788 ; 
        RECT 28.028 180.414 28.132 184.788 ; 
        RECT 27.596 180.414 27.7 184.788 ; 
        RECT 27.164 180.414 27.268 184.788 ; 
        RECT 26.732 180.414 26.836 184.788 ; 
        RECT 26.3 180.414 26.404 184.788 ; 
        RECT 25.868 180.414 25.972 184.788 ; 
        RECT 25.436 180.414 25.54 184.788 ; 
        RECT 25.004 180.414 25.108 184.788 ; 
        RECT 24.572 180.414 24.676 184.788 ; 
        RECT 24.14 180.414 24.244 184.788 ; 
        RECT 23.708 180.414 23.812 184.788 ; 
        RECT 22.856 180.414 23.164 184.788 ; 
        RECT 15.284 180.414 15.592 184.788 ; 
        RECT 14.636 180.414 14.74 184.788 ; 
        RECT 14.204 180.414 14.308 184.788 ; 
        RECT 13.772 180.414 13.876 184.788 ; 
        RECT 13.34 180.414 13.444 184.788 ; 
        RECT 12.908 180.414 13.012 184.788 ; 
        RECT 12.476 180.414 12.58 184.788 ; 
        RECT 12.044 180.414 12.148 184.788 ; 
        RECT 11.612 180.414 11.716 184.788 ; 
        RECT 11.18 180.414 11.284 184.788 ; 
        RECT 10.748 180.414 10.852 184.788 ; 
        RECT 10.316 180.414 10.42 184.788 ; 
        RECT 9.884 180.414 9.988 184.788 ; 
        RECT 9.452 180.414 9.556 184.788 ; 
        RECT 9.02 180.414 9.124 184.788 ; 
        RECT 8.588 180.414 8.692 184.788 ; 
        RECT 8.156 180.414 8.26 184.788 ; 
        RECT 7.724 180.414 7.828 184.788 ; 
        RECT 7.292 180.414 7.396 184.788 ; 
        RECT 6.86 180.414 6.964 184.788 ; 
        RECT 6.428 180.414 6.532 184.788 ; 
        RECT 5.996 180.414 6.1 184.788 ; 
        RECT 5.564 180.414 5.668 184.788 ; 
        RECT 5.132 180.414 5.236 184.788 ; 
        RECT 4.7 180.414 4.804 184.788 ; 
        RECT 4.268 180.414 4.372 184.788 ; 
        RECT 3.836 180.414 3.94 184.788 ; 
        RECT 3.404 180.414 3.508 184.788 ; 
        RECT 2.972 180.414 3.076 184.788 ; 
        RECT 2.54 180.414 2.644 184.788 ; 
        RECT 2.108 180.414 2.212 184.788 ; 
        RECT 1.676 180.414 1.78 184.788 ; 
        RECT 1.244 180.414 1.348 184.788 ; 
        RECT 0.812 180.414 0.916 184.788 ; 
        RECT 0 180.414 0.34 184.788 ; 
        RECT 20.72 184.734 21.232 189.108 ; 
        RECT 20.664 187.396 21.232 188.686 ; 
        RECT 20.072 186.304 20.32 189.108 ; 
        RECT 20.016 187.542 20.32 188.156 ; 
        RECT 20.072 184.734 20.176 189.108 ; 
        RECT 20.072 185.218 20.232 186.176 ; 
        RECT 20.072 184.734 20.32 185.09 ; 
        RECT 18.884 186.536 19.708 189.108 ; 
        RECT 19.604 184.734 19.708 189.108 ; 
        RECT 18.884 187.644 19.764 188.676 ; 
        RECT 18.884 184.734 19.276 189.108 ; 
        RECT 17.216 184.734 17.548 189.108 ; 
        RECT 17.216 185.088 17.604 188.83 ; 
        RECT 38.108 184.734 38.448 189.108 ; 
        RECT 37.532 184.734 37.636 189.108 ; 
        RECT 37.1 184.734 37.204 189.108 ; 
        RECT 36.668 184.734 36.772 189.108 ; 
        RECT 36.236 184.734 36.34 189.108 ; 
        RECT 35.804 184.734 35.908 189.108 ; 
        RECT 35.372 184.734 35.476 189.108 ; 
        RECT 34.94 184.734 35.044 189.108 ; 
        RECT 34.508 184.734 34.612 189.108 ; 
        RECT 34.076 184.734 34.18 189.108 ; 
        RECT 33.644 184.734 33.748 189.108 ; 
        RECT 33.212 184.734 33.316 189.108 ; 
        RECT 32.78 184.734 32.884 189.108 ; 
        RECT 32.348 184.734 32.452 189.108 ; 
        RECT 31.916 184.734 32.02 189.108 ; 
        RECT 31.484 184.734 31.588 189.108 ; 
        RECT 31.052 184.734 31.156 189.108 ; 
        RECT 30.62 184.734 30.724 189.108 ; 
        RECT 30.188 184.734 30.292 189.108 ; 
        RECT 29.756 184.734 29.86 189.108 ; 
        RECT 29.324 184.734 29.428 189.108 ; 
        RECT 28.892 184.734 28.996 189.108 ; 
        RECT 28.46 184.734 28.564 189.108 ; 
        RECT 28.028 184.734 28.132 189.108 ; 
        RECT 27.596 184.734 27.7 189.108 ; 
        RECT 27.164 184.734 27.268 189.108 ; 
        RECT 26.732 184.734 26.836 189.108 ; 
        RECT 26.3 184.734 26.404 189.108 ; 
        RECT 25.868 184.734 25.972 189.108 ; 
        RECT 25.436 184.734 25.54 189.108 ; 
        RECT 25.004 184.734 25.108 189.108 ; 
        RECT 24.572 184.734 24.676 189.108 ; 
        RECT 24.14 184.734 24.244 189.108 ; 
        RECT 23.708 184.734 23.812 189.108 ; 
        RECT 22.856 184.734 23.164 189.108 ; 
        RECT 15.284 184.734 15.592 189.108 ; 
        RECT 14.636 184.734 14.74 189.108 ; 
        RECT 14.204 184.734 14.308 189.108 ; 
        RECT 13.772 184.734 13.876 189.108 ; 
        RECT 13.34 184.734 13.444 189.108 ; 
        RECT 12.908 184.734 13.012 189.108 ; 
        RECT 12.476 184.734 12.58 189.108 ; 
        RECT 12.044 184.734 12.148 189.108 ; 
        RECT 11.612 184.734 11.716 189.108 ; 
        RECT 11.18 184.734 11.284 189.108 ; 
        RECT 10.748 184.734 10.852 189.108 ; 
        RECT 10.316 184.734 10.42 189.108 ; 
        RECT 9.884 184.734 9.988 189.108 ; 
        RECT 9.452 184.734 9.556 189.108 ; 
        RECT 9.02 184.734 9.124 189.108 ; 
        RECT 8.588 184.734 8.692 189.108 ; 
        RECT 8.156 184.734 8.26 189.108 ; 
        RECT 7.724 184.734 7.828 189.108 ; 
        RECT 7.292 184.734 7.396 189.108 ; 
        RECT 6.86 184.734 6.964 189.108 ; 
        RECT 6.428 184.734 6.532 189.108 ; 
        RECT 5.996 184.734 6.1 189.108 ; 
        RECT 5.564 184.734 5.668 189.108 ; 
        RECT 5.132 184.734 5.236 189.108 ; 
        RECT 4.7 184.734 4.804 189.108 ; 
        RECT 4.268 184.734 4.372 189.108 ; 
        RECT 3.836 184.734 3.94 189.108 ; 
        RECT 3.404 184.734 3.508 189.108 ; 
        RECT 2.972 184.734 3.076 189.108 ; 
        RECT 2.54 184.734 2.644 189.108 ; 
        RECT 2.108 184.734 2.212 189.108 ; 
        RECT 1.676 184.734 1.78 189.108 ; 
        RECT 1.244 184.734 1.348 189.108 ; 
        RECT 0.812 184.734 0.916 189.108 ; 
        RECT 0 184.734 0.34 189.108 ; 
        RECT 20.72 189.054 21.232 193.428 ; 
        RECT 20.664 191.716 21.232 193.006 ; 
        RECT 20.072 190.624 20.32 193.428 ; 
        RECT 20.016 191.862 20.32 192.476 ; 
        RECT 20.072 189.054 20.176 193.428 ; 
        RECT 20.072 189.538 20.232 190.496 ; 
        RECT 20.072 189.054 20.32 189.41 ; 
        RECT 18.884 190.856 19.708 193.428 ; 
        RECT 19.604 189.054 19.708 193.428 ; 
        RECT 18.884 191.964 19.764 192.996 ; 
        RECT 18.884 189.054 19.276 193.428 ; 
        RECT 17.216 189.054 17.548 193.428 ; 
        RECT 17.216 189.408 17.604 193.15 ; 
        RECT 38.108 189.054 38.448 193.428 ; 
        RECT 37.532 189.054 37.636 193.428 ; 
        RECT 37.1 189.054 37.204 193.428 ; 
        RECT 36.668 189.054 36.772 193.428 ; 
        RECT 36.236 189.054 36.34 193.428 ; 
        RECT 35.804 189.054 35.908 193.428 ; 
        RECT 35.372 189.054 35.476 193.428 ; 
        RECT 34.94 189.054 35.044 193.428 ; 
        RECT 34.508 189.054 34.612 193.428 ; 
        RECT 34.076 189.054 34.18 193.428 ; 
        RECT 33.644 189.054 33.748 193.428 ; 
        RECT 33.212 189.054 33.316 193.428 ; 
        RECT 32.78 189.054 32.884 193.428 ; 
        RECT 32.348 189.054 32.452 193.428 ; 
        RECT 31.916 189.054 32.02 193.428 ; 
        RECT 31.484 189.054 31.588 193.428 ; 
        RECT 31.052 189.054 31.156 193.428 ; 
        RECT 30.62 189.054 30.724 193.428 ; 
        RECT 30.188 189.054 30.292 193.428 ; 
        RECT 29.756 189.054 29.86 193.428 ; 
        RECT 29.324 189.054 29.428 193.428 ; 
        RECT 28.892 189.054 28.996 193.428 ; 
        RECT 28.46 189.054 28.564 193.428 ; 
        RECT 28.028 189.054 28.132 193.428 ; 
        RECT 27.596 189.054 27.7 193.428 ; 
        RECT 27.164 189.054 27.268 193.428 ; 
        RECT 26.732 189.054 26.836 193.428 ; 
        RECT 26.3 189.054 26.404 193.428 ; 
        RECT 25.868 189.054 25.972 193.428 ; 
        RECT 25.436 189.054 25.54 193.428 ; 
        RECT 25.004 189.054 25.108 193.428 ; 
        RECT 24.572 189.054 24.676 193.428 ; 
        RECT 24.14 189.054 24.244 193.428 ; 
        RECT 23.708 189.054 23.812 193.428 ; 
        RECT 22.856 189.054 23.164 193.428 ; 
        RECT 15.284 189.054 15.592 193.428 ; 
        RECT 14.636 189.054 14.74 193.428 ; 
        RECT 14.204 189.054 14.308 193.428 ; 
        RECT 13.772 189.054 13.876 193.428 ; 
        RECT 13.34 189.054 13.444 193.428 ; 
        RECT 12.908 189.054 13.012 193.428 ; 
        RECT 12.476 189.054 12.58 193.428 ; 
        RECT 12.044 189.054 12.148 193.428 ; 
        RECT 11.612 189.054 11.716 193.428 ; 
        RECT 11.18 189.054 11.284 193.428 ; 
        RECT 10.748 189.054 10.852 193.428 ; 
        RECT 10.316 189.054 10.42 193.428 ; 
        RECT 9.884 189.054 9.988 193.428 ; 
        RECT 9.452 189.054 9.556 193.428 ; 
        RECT 9.02 189.054 9.124 193.428 ; 
        RECT 8.588 189.054 8.692 193.428 ; 
        RECT 8.156 189.054 8.26 193.428 ; 
        RECT 7.724 189.054 7.828 193.428 ; 
        RECT 7.292 189.054 7.396 193.428 ; 
        RECT 6.86 189.054 6.964 193.428 ; 
        RECT 6.428 189.054 6.532 193.428 ; 
        RECT 5.996 189.054 6.1 193.428 ; 
        RECT 5.564 189.054 5.668 193.428 ; 
        RECT 5.132 189.054 5.236 193.428 ; 
        RECT 4.7 189.054 4.804 193.428 ; 
        RECT 4.268 189.054 4.372 193.428 ; 
        RECT 3.836 189.054 3.94 193.428 ; 
        RECT 3.404 189.054 3.508 193.428 ; 
        RECT 2.972 189.054 3.076 193.428 ; 
        RECT 2.54 189.054 2.644 193.428 ; 
        RECT 2.108 189.054 2.212 193.428 ; 
        RECT 1.676 189.054 1.78 193.428 ; 
        RECT 1.244 189.054 1.348 193.428 ; 
        RECT 0.812 189.054 0.916 193.428 ; 
        RECT 0 189.054 0.34 193.428 ; 
        RECT 20.72 193.374 21.232 197.748 ; 
        RECT 20.664 196.036 21.232 197.326 ; 
        RECT 20.072 194.944 20.32 197.748 ; 
        RECT 20.016 196.182 20.32 196.796 ; 
        RECT 20.072 193.374 20.176 197.748 ; 
        RECT 20.072 193.858 20.232 194.816 ; 
        RECT 20.072 193.374 20.32 193.73 ; 
        RECT 18.884 195.176 19.708 197.748 ; 
        RECT 19.604 193.374 19.708 197.748 ; 
        RECT 18.884 196.284 19.764 197.316 ; 
        RECT 18.884 193.374 19.276 197.748 ; 
        RECT 17.216 193.374 17.548 197.748 ; 
        RECT 17.216 193.728 17.604 197.47 ; 
        RECT 38.108 193.374 38.448 197.748 ; 
        RECT 37.532 193.374 37.636 197.748 ; 
        RECT 37.1 193.374 37.204 197.748 ; 
        RECT 36.668 193.374 36.772 197.748 ; 
        RECT 36.236 193.374 36.34 197.748 ; 
        RECT 35.804 193.374 35.908 197.748 ; 
        RECT 35.372 193.374 35.476 197.748 ; 
        RECT 34.94 193.374 35.044 197.748 ; 
        RECT 34.508 193.374 34.612 197.748 ; 
        RECT 34.076 193.374 34.18 197.748 ; 
        RECT 33.644 193.374 33.748 197.748 ; 
        RECT 33.212 193.374 33.316 197.748 ; 
        RECT 32.78 193.374 32.884 197.748 ; 
        RECT 32.348 193.374 32.452 197.748 ; 
        RECT 31.916 193.374 32.02 197.748 ; 
        RECT 31.484 193.374 31.588 197.748 ; 
        RECT 31.052 193.374 31.156 197.748 ; 
        RECT 30.62 193.374 30.724 197.748 ; 
        RECT 30.188 193.374 30.292 197.748 ; 
        RECT 29.756 193.374 29.86 197.748 ; 
        RECT 29.324 193.374 29.428 197.748 ; 
        RECT 28.892 193.374 28.996 197.748 ; 
        RECT 28.46 193.374 28.564 197.748 ; 
        RECT 28.028 193.374 28.132 197.748 ; 
        RECT 27.596 193.374 27.7 197.748 ; 
        RECT 27.164 193.374 27.268 197.748 ; 
        RECT 26.732 193.374 26.836 197.748 ; 
        RECT 26.3 193.374 26.404 197.748 ; 
        RECT 25.868 193.374 25.972 197.748 ; 
        RECT 25.436 193.374 25.54 197.748 ; 
        RECT 25.004 193.374 25.108 197.748 ; 
        RECT 24.572 193.374 24.676 197.748 ; 
        RECT 24.14 193.374 24.244 197.748 ; 
        RECT 23.708 193.374 23.812 197.748 ; 
        RECT 22.856 193.374 23.164 197.748 ; 
        RECT 15.284 193.374 15.592 197.748 ; 
        RECT 14.636 193.374 14.74 197.748 ; 
        RECT 14.204 193.374 14.308 197.748 ; 
        RECT 13.772 193.374 13.876 197.748 ; 
        RECT 13.34 193.374 13.444 197.748 ; 
        RECT 12.908 193.374 13.012 197.748 ; 
        RECT 12.476 193.374 12.58 197.748 ; 
        RECT 12.044 193.374 12.148 197.748 ; 
        RECT 11.612 193.374 11.716 197.748 ; 
        RECT 11.18 193.374 11.284 197.748 ; 
        RECT 10.748 193.374 10.852 197.748 ; 
        RECT 10.316 193.374 10.42 197.748 ; 
        RECT 9.884 193.374 9.988 197.748 ; 
        RECT 9.452 193.374 9.556 197.748 ; 
        RECT 9.02 193.374 9.124 197.748 ; 
        RECT 8.588 193.374 8.692 197.748 ; 
        RECT 8.156 193.374 8.26 197.748 ; 
        RECT 7.724 193.374 7.828 197.748 ; 
        RECT 7.292 193.374 7.396 197.748 ; 
        RECT 6.86 193.374 6.964 197.748 ; 
        RECT 6.428 193.374 6.532 197.748 ; 
        RECT 5.996 193.374 6.1 197.748 ; 
        RECT 5.564 193.374 5.668 197.748 ; 
        RECT 5.132 193.374 5.236 197.748 ; 
        RECT 4.7 193.374 4.804 197.748 ; 
        RECT 4.268 193.374 4.372 197.748 ; 
        RECT 3.836 193.374 3.94 197.748 ; 
        RECT 3.404 193.374 3.508 197.748 ; 
        RECT 2.972 193.374 3.076 197.748 ; 
        RECT 2.54 193.374 2.644 197.748 ; 
        RECT 2.108 193.374 2.212 197.748 ; 
        RECT 1.676 193.374 1.78 197.748 ; 
        RECT 1.244 193.374 1.348 197.748 ; 
        RECT 0.812 193.374 0.916 197.748 ; 
        RECT 0 193.374 0.34 197.748 ; 
        RECT 20.72 197.694 21.232 202.068 ; 
        RECT 20.664 200.356 21.232 201.646 ; 
        RECT 20.072 199.264 20.32 202.068 ; 
        RECT 20.016 200.502 20.32 201.116 ; 
        RECT 20.072 197.694 20.176 202.068 ; 
        RECT 20.072 198.178 20.232 199.136 ; 
        RECT 20.072 197.694 20.32 198.05 ; 
        RECT 18.884 199.496 19.708 202.068 ; 
        RECT 19.604 197.694 19.708 202.068 ; 
        RECT 18.884 200.604 19.764 201.636 ; 
        RECT 18.884 197.694 19.276 202.068 ; 
        RECT 17.216 197.694 17.548 202.068 ; 
        RECT 17.216 198.048 17.604 201.79 ; 
        RECT 38.108 197.694 38.448 202.068 ; 
        RECT 37.532 197.694 37.636 202.068 ; 
        RECT 37.1 197.694 37.204 202.068 ; 
        RECT 36.668 197.694 36.772 202.068 ; 
        RECT 36.236 197.694 36.34 202.068 ; 
        RECT 35.804 197.694 35.908 202.068 ; 
        RECT 35.372 197.694 35.476 202.068 ; 
        RECT 34.94 197.694 35.044 202.068 ; 
        RECT 34.508 197.694 34.612 202.068 ; 
        RECT 34.076 197.694 34.18 202.068 ; 
        RECT 33.644 197.694 33.748 202.068 ; 
        RECT 33.212 197.694 33.316 202.068 ; 
        RECT 32.78 197.694 32.884 202.068 ; 
        RECT 32.348 197.694 32.452 202.068 ; 
        RECT 31.916 197.694 32.02 202.068 ; 
        RECT 31.484 197.694 31.588 202.068 ; 
        RECT 31.052 197.694 31.156 202.068 ; 
        RECT 30.62 197.694 30.724 202.068 ; 
        RECT 30.188 197.694 30.292 202.068 ; 
        RECT 29.756 197.694 29.86 202.068 ; 
        RECT 29.324 197.694 29.428 202.068 ; 
        RECT 28.892 197.694 28.996 202.068 ; 
        RECT 28.46 197.694 28.564 202.068 ; 
        RECT 28.028 197.694 28.132 202.068 ; 
        RECT 27.596 197.694 27.7 202.068 ; 
        RECT 27.164 197.694 27.268 202.068 ; 
        RECT 26.732 197.694 26.836 202.068 ; 
        RECT 26.3 197.694 26.404 202.068 ; 
        RECT 25.868 197.694 25.972 202.068 ; 
        RECT 25.436 197.694 25.54 202.068 ; 
        RECT 25.004 197.694 25.108 202.068 ; 
        RECT 24.572 197.694 24.676 202.068 ; 
        RECT 24.14 197.694 24.244 202.068 ; 
        RECT 23.708 197.694 23.812 202.068 ; 
        RECT 22.856 197.694 23.164 202.068 ; 
        RECT 15.284 197.694 15.592 202.068 ; 
        RECT 14.636 197.694 14.74 202.068 ; 
        RECT 14.204 197.694 14.308 202.068 ; 
        RECT 13.772 197.694 13.876 202.068 ; 
        RECT 13.34 197.694 13.444 202.068 ; 
        RECT 12.908 197.694 13.012 202.068 ; 
        RECT 12.476 197.694 12.58 202.068 ; 
        RECT 12.044 197.694 12.148 202.068 ; 
        RECT 11.612 197.694 11.716 202.068 ; 
        RECT 11.18 197.694 11.284 202.068 ; 
        RECT 10.748 197.694 10.852 202.068 ; 
        RECT 10.316 197.694 10.42 202.068 ; 
        RECT 9.884 197.694 9.988 202.068 ; 
        RECT 9.452 197.694 9.556 202.068 ; 
        RECT 9.02 197.694 9.124 202.068 ; 
        RECT 8.588 197.694 8.692 202.068 ; 
        RECT 8.156 197.694 8.26 202.068 ; 
        RECT 7.724 197.694 7.828 202.068 ; 
        RECT 7.292 197.694 7.396 202.068 ; 
        RECT 6.86 197.694 6.964 202.068 ; 
        RECT 6.428 197.694 6.532 202.068 ; 
        RECT 5.996 197.694 6.1 202.068 ; 
        RECT 5.564 197.694 5.668 202.068 ; 
        RECT 5.132 197.694 5.236 202.068 ; 
        RECT 4.7 197.694 4.804 202.068 ; 
        RECT 4.268 197.694 4.372 202.068 ; 
        RECT 3.836 197.694 3.94 202.068 ; 
        RECT 3.404 197.694 3.508 202.068 ; 
        RECT 2.972 197.694 3.076 202.068 ; 
        RECT 2.54 197.694 2.644 202.068 ; 
        RECT 2.108 197.694 2.212 202.068 ; 
        RECT 1.676 197.694 1.78 202.068 ; 
        RECT 1.244 197.694 1.348 202.068 ; 
        RECT 0.812 197.694 0.916 202.068 ; 
        RECT 0 197.694 0.34 202.068 ; 
        RECT 20.72 202.014 21.232 206.388 ; 
        RECT 20.664 204.676 21.232 205.966 ; 
        RECT 20.072 203.584 20.32 206.388 ; 
        RECT 20.016 204.822 20.32 205.436 ; 
        RECT 20.072 202.014 20.176 206.388 ; 
        RECT 20.072 202.498 20.232 203.456 ; 
        RECT 20.072 202.014 20.32 202.37 ; 
        RECT 18.884 203.816 19.708 206.388 ; 
        RECT 19.604 202.014 19.708 206.388 ; 
        RECT 18.884 204.924 19.764 205.956 ; 
        RECT 18.884 202.014 19.276 206.388 ; 
        RECT 17.216 202.014 17.548 206.388 ; 
        RECT 17.216 202.368 17.604 206.11 ; 
        RECT 38.108 202.014 38.448 206.388 ; 
        RECT 37.532 202.014 37.636 206.388 ; 
        RECT 37.1 202.014 37.204 206.388 ; 
        RECT 36.668 202.014 36.772 206.388 ; 
        RECT 36.236 202.014 36.34 206.388 ; 
        RECT 35.804 202.014 35.908 206.388 ; 
        RECT 35.372 202.014 35.476 206.388 ; 
        RECT 34.94 202.014 35.044 206.388 ; 
        RECT 34.508 202.014 34.612 206.388 ; 
        RECT 34.076 202.014 34.18 206.388 ; 
        RECT 33.644 202.014 33.748 206.388 ; 
        RECT 33.212 202.014 33.316 206.388 ; 
        RECT 32.78 202.014 32.884 206.388 ; 
        RECT 32.348 202.014 32.452 206.388 ; 
        RECT 31.916 202.014 32.02 206.388 ; 
        RECT 31.484 202.014 31.588 206.388 ; 
        RECT 31.052 202.014 31.156 206.388 ; 
        RECT 30.62 202.014 30.724 206.388 ; 
        RECT 30.188 202.014 30.292 206.388 ; 
        RECT 29.756 202.014 29.86 206.388 ; 
        RECT 29.324 202.014 29.428 206.388 ; 
        RECT 28.892 202.014 28.996 206.388 ; 
        RECT 28.46 202.014 28.564 206.388 ; 
        RECT 28.028 202.014 28.132 206.388 ; 
        RECT 27.596 202.014 27.7 206.388 ; 
        RECT 27.164 202.014 27.268 206.388 ; 
        RECT 26.732 202.014 26.836 206.388 ; 
        RECT 26.3 202.014 26.404 206.388 ; 
        RECT 25.868 202.014 25.972 206.388 ; 
        RECT 25.436 202.014 25.54 206.388 ; 
        RECT 25.004 202.014 25.108 206.388 ; 
        RECT 24.572 202.014 24.676 206.388 ; 
        RECT 24.14 202.014 24.244 206.388 ; 
        RECT 23.708 202.014 23.812 206.388 ; 
        RECT 22.856 202.014 23.164 206.388 ; 
        RECT 15.284 202.014 15.592 206.388 ; 
        RECT 14.636 202.014 14.74 206.388 ; 
        RECT 14.204 202.014 14.308 206.388 ; 
        RECT 13.772 202.014 13.876 206.388 ; 
        RECT 13.34 202.014 13.444 206.388 ; 
        RECT 12.908 202.014 13.012 206.388 ; 
        RECT 12.476 202.014 12.58 206.388 ; 
        RECT 12.044 202.014 12.148 206.388 ; 
        RECT 11.612 202.014 11.716 206.388 ; 
        RECT 11.18 202.014 11.284 206.388 ; 
        RECT 10.748 202.014 10.852 206.388 ; 
        RECT 10.316 202.014 10.42 206.388 ; 
        RECT 9.884 202.014 9.988 206.388 ; 
        RECT 9.452 202.014 9.556 206.388 ; 
        RECT 9.02 202.014 9.124 206.388 ; 
        RECT 8.588 202.014 8.692 206.388 ; 
        RECT 8.156 202.014 8.26 206.388 ; 
        RECT 7.724 202.014 7.828 206.388 ; 
        RECT 7.292 202.014 7.396 206.388 ; 
        RECT 6.86 202.014 6.964 206.388 ; 
        RECT 6.428 202.014 6.532 206.388 ; 
        RECT 5.996 202.014 6.1 206.388 ; 
        RECT 5.564 202.014 5.668 206.388 ; 
        RECT 5.132 202.014 5.236 206.388 ; 
        RECT 4.7 202.014 4.804 206.388 ; 
        RECT 4.268 202.014 4.372 206.388 ; 
        RECT 3.836 202.014 3.94 206.388 ; 
        RECT 3.404 202.014 3.508 206.388 ; 
        RECT 2.972 202.014 3.076 206.388 ; 
        RECT 2.54 202.014 2.644 206.388 ; 
        RECT 2.108 202.014 2.212 206.388 ; 
        RECT 1.676 202.014 1.78 206.388 ; 
        RECT 1.244 202.014 1.348 206.388 ; 
        RECT 0.812 202.014 0.916 206.388 ; 
        RECT 0 202.014 0.34 206.388 ; 
        RECT 20.72 206.334 21.232 210.708 ; 
        RECT 20.664 208.996 21.232 210.286 ; 
        RECT 20.072 207.904 20.32 210.708 ; 
        RECT 20.016 209.142 20.32 209.756 ; 
        RECT 20.072 206.334 20.176 210.708 ; 
        RECT 20.072 206.818 20.232 207.776 ; 
        RECT 20.072 206.334 20.32 206.69 ; 
        RECT 18.884 208.136 19.708 210.708 ; 
        RECT 19.604 206.334 19.708 210.708 ; 
        RECT 18.884 209.244 19.764 210.276 ; 
        RECT 18.884 206.334 19.276 210.708 ; 
        RECT 17.216 206.334 17.548 210.708 ; 
        RECT 17.216 206.688 17.604 210.43 ; 
        RECT 38.108 206.334 38.448 210.708 ; 
        RECT 37.532 206.334 37.636 210.708 ; 
        RECT 37.1 206.334 37.204 210.708 ; 
        RECT 36.668 206.334 36.772 210.708 ; 
        RECT 36.236 206.334 36.34 210.708 ; 
        RECT 35.804 206.334 35.908 210.708 ; 
        RECT 35.372 206.334 35.476 210.708 ; 
        RECT 34.94 206.334 35.044 210.708 ; 
        RECT 34.508 206.334 34.612 210.708 ; 
        RECT 34.076 206.334 34.18 210.708 ; 
        RECT 33.644 206.334 33.748 210.708 ; 
        RECT 33.212 206.334 33.316 210.708 ; 
        RECT 32.78 206.334 32.884 210.708 ; 
        RECT 32.348 206.334 32.452 210.708 ; 
        RECT 31.916 206.334 32.02 210.708 ; 
        RECT 31.484 206.334 31.588 210.708 ; 
        RECT 31.052 206.334 31.156 210.708 ; 
        RECT 30.62 206.334 30.724 210.708 ; 
        RECT 30.188 206.334 30.292 210.708 ; 
        RECT 29.756 206.334 29.86 210.708 ; 
        RECT 29.324 206.334 29.428 210.708 ; 
        RECT 28.892 206.334 28.996 210.708 ; 
        RECT 28.46 206.334 28.564 210.708 ; 
        RECT 28.028 206.334 28.132 210.708 ; 
        RECT 27.596 206.334 27.7 210.708 ; 
        RECT 27.164 206.334 27.268 210.708 ; 
        RECT 26.732 206.334 26.836 210.708 ; 
        RECT 26.3 206.334 26.404 210.708 ; 
        RECT 25.868 206.334 25.972 210.708 ; 
        RECT 25.436 206.334 25.54 210.708 ; 
        RECT 25.004 206.334 25.108 210.708 ; 
        RECT 24.572 206.334 24.676 210.708 ; 
        RECT 24.14 206.334 24.244 210.708 ; 
        RECT 23.708 206.334 23.812 210.708 ; 
        RECT 22.856 206.334 23.164 210.708 ; 
        RECT 15.284 206.334 15.592 210.708 ; 
        RECT 14.636 206.334 14.74 210.708 ; 
        RECT 14.204 206.334 14.308 210.708 ; 
        RECT 13.772 206.334 13.876 210.708 ; 
        RECT 13.34 206.334 13.444 210.708 ; 
        RECT 12.908 206.334 13.012 210.708 ; 
        RECT 12.476 206.334 12.58 210.708 ; 
        RECT 12.044 206.334 12.148 210.708 ; 
        RECT 11.612 206.334 11.716 210.708 ; 
        RECT 11.18 206.334 11.284 210.708 ; 
        RECT 10.748 206.334 10.852 210.708 ; 
        RECT 10.316 206.334 10.42 210.708 ; 
        RECT 9.884 206.334 9.988 210.708 ; 
        RECT 9.452 206.334 9.556 210.708 ; 
        RECT 9.02 206.334 9.124 210.708 ; 
        RECT 8.588 206.334 8.692 210.708 ; 
        RECT 8.156 206.334 8.26 210.708 ; 
        RECT 7.724 206.334 7.828 210.708 ; 
        RECT 7.292 206.334 7.396 210.708 ; 
        RECT 6.86 206.334 6.964 210.708 ; 
        RECT 6.428 206.334 6.532 210.708 ; 
        RECT 5.996 206.334 6.1 210.708 ; 
        RECT 5.564 206.334 5.668 210.708 ; 
        RECT 5.132 206.334 5.236 210.708 ; 
        RECT 4.7 206.334 4.804 210.708 ; 
        RECT 4.268 206.334 4.372 210.708 ; 
        RECT 3.836 206.334 3.94 210.708 ; 
        RECT 3.404 206.334 3.508 210.708 ; 
        RECT 2.972 206.334 3.076 210.708 ; 
        RECT 2.54 206.334 2.644 210.708 ; 
        RECT 2.108 206.334 2.212 210.708 ; 
        RECT 1.676 206.334 1.78 210.708 ; 
        RECT 1.244 206.334 1.348 210.708 ; 
        RECT 0.812 206.334 0.916 210.708 ; 
        RECT 0 206.334 0.34 210.708 ; 
        RECT 20.72 210.654 21.232 215.028 ; 
        RECT 20.664 213.316 21.232 214.606 ; 
        RECT 20.072 212.224 20.32 215.028 ; 
        RECT 20.016 213.462 20.32 214.076 ; 
        RECT 20.072 210.654 20.176 215.028 ; 
        RECT 20.072 211.138 20.232 212.096 ; 
        RECT 20.072 210.654 20.32 211.01 ; 
        RECT 18.884 212.456 19.708 215.028 ; 
        RECT 19.604 210.654 19.708 215.028 ; 
        RECT 18.884 213.564 19.764 214.596 ; 
        RECT 18.884 210.654 19.276 215.028 ; 
        RECT 17.216 210.654 17.548 215.028 ; 
        RECT 17.216 211.008 17.604 214.75 ; 
        RECT 38.108 210.654 38.448 215.028 ; 
        RECT 37.532 210.654 37.636 215.028 ; 
        RECT 37.1 210.654 37.204 215.028 ; 
        RECT 36.668 210.654 36.772 215.028 ; 
        RECT 36.236 210.654 36.34 215.028 ; 
        RECT 35.804 210.654 35.908 215.028 ; 
        RECT 35.372 210.654 35.476 215.028 ; 
        RECT 34.94 210.654 35.044 215.028 ; 
        RECT 34.508 210.654 34.612 215.028 ; 
        RECT 34.076 210.654 34.18 215.028 ; 
        RECT 33.644 210.654 33.748 215.028 ; 
        RECT 33.212 210.654 33.316 215.028 ; 
        RECT 32.78 210.654 32.884 215.028 ; 
        RECT 32.348 210.654 32.452 215.028 ; 
        RECT 31.916 210.654 32.02 215.028 ; 
        RECT 31.484 210.654 31.588 215.028 ; 
        RECT 31.052 210.654 31.156 215.028 ; 
        RECT 30.62 210.654 30.724 215.028 ; 
        RECT 30.188 210.654 30.292 215.028 ; 
        RECT 29.756 210.654 29.86 215.028 ; 
        RECT 29.324 210.654 29.428 215.028 ; 
        RECT 28.892 210.654 28.996 215.028 ; 
        RECT 28.46 210.654 28.564 215.028 ; 
        RECT 28.028 210.654 28.132 215.028 ; 
        RECT 27.596 210.654 27.7 215.028 ; 
        RECT 27.164 210.654 27.268 215.028 ; 
        RECT 26.732 210.654 26.836 215.028 ; 
        RECT 26.3 210.654 26.404 215.028 ; 
        RECT 25.868 210.654 25.972 215.028 ; 
        RECT 25.436 210.654 25.54 215.028 ; 
        RECT 25.004 210.654 25.108 215.028 ; 
        RECT 24.572 210.654 24.676 215.028 ; 
        RECT 24.14 210.654 24.244 215.028 ; 
        RECT 23.708 210.654 23.812 215.028 ; 
        RECT 22.856 210.654 23.164 215.028 ; 
        RECT 15.284 210.654 15.592 215.028 ; 
        RECT 14.636 210.654 14.74 215.028 ; 
        RECT 14.204 210.654 14.308 215.028 ; 
        RECT 13.772 210.654 13.876 215.028 ; 
        RECT 13.34 210.654 13.444 215.028 ; 
        RECT 12.908 210.654 13.012 215.028 ; 
        RECT 12.476 210.654 12.58 215.028 ; 
        RECT 12.044 210.654 12.148 215.028 ; 
        RECT 11.612 210.654 11.716 215.028 ; 
        RECT 11.18 210.654 11.284 215.028 ; 
        RECT 10.748 210.654 10.852 215.028 ; 
        RECT 10.316 210.654 10.42 215.028 ; 
        RECT 9.884 210.654 9.988 215.028 ; 
        RECT 9.452 210.654 9.556 215.028 ; 
        RECT 9.02 210.654 9.124 215.028 ; 
        RECT 8.588 210.654 8.692 215.028 ; 
        RECT 8.156 210.654 8.26 215.028 ; 
        RECT 7.724 210.654 7.828 215.028 ; 
        RECT 7.292 210.654 7.396 215.028 ; 
        RECT 6.86 210.654 6.964 215.028 ; 
        RECT 6.428 210.654 6.532 215.028 ; 
        RECT 5.996 210.654 6.1 215.028 ; 
        RECT 5.564 210.654 5.668 215.028 ; 
        RECT 5.132 210.654 5.236 215.028 ; 
        RECT 4.7 210.654 4.804 215.028 ; 
        RECT 4.268 210.654 4.372 215.028 ; 
        RECT 3.836 210.654 3.94 215.028 ; 
        RECT 3.404 210.654 3.508 215.028 ; 
        RECT 2.972 210.654 3.076 215.028 ; 
        RECT 2.54 210.654 2.644 215.028 ; 
        RECT 2.108 210.654 2.212 215.028 ; 
        RECT 1.676 210.654 1.78 215.028 ; 
        RECT 1.244 210.654 1.348 215.028 ; 
        RECT 0.812 210.654 0.916 215.028 ; 
        RECT 0 210.654 0.34 215.028 ; 
        RECT 20.72 214.974 21.232 219.348 ; 
        RECT 20.664 217.636 21.232 218.926 ; 
        RECT 20.072 216.544 20.32 219.348 ; 
        RECT 20.016 217.782 20.32 218.396 ; 
        RECT 20.072 214.974 20.176 219.348 ; 
        RECT 20.072 215.458 20.232 216.416 ; 
        RECT 20.072 214.974 20.32 215.33 ; 
        RECT 18.884 216.776 19.708 219.348 ; 
        RECT 19.604 214.974 19.708 219.348 ; 
        RECT 18.884 217.884 19.764 218.916 ; 
        RECT 18.884 214.974 19.276 219.348 ; 
        RECT 17.216 214.974 17.548 219.348 ; 
        RECT 17.216 215.328 17.604 219.07 ; 
        RECT 38.108 214.974 38.448 219.348 ; 
        RECT 37.532 214.974 37.636 219.348 ; 
        RECT 37.1 214.974 37.204 219.348 ; 
        RECT 36.668 214.974 36.772 219.348 ; 
        RECT 36.236 214.974 36.34 219.348 ; 
        RECT 35.804 214.974 35.908 219.348 ; 
        RECT 35.372 214.974 35.476 219.348 ; 
        RECT 34.94 214.974 35.044 219.348 ; 
        RECT 34.508 214.974 34.612 219.348 ; 
        RECT 34.076 214.974 34.18 219.348 ; 
        RECT 33.644 214.974 33.748 219.348 ; 
        RECT 33.212 214.974 33.316 219.348 ; 
        RECT 32.78 214.974 32.884 219.348 ; 
        RECT 32.348 214.974 32.452 219.348 ; 
        RECT 31.916 214.974 32.02 219.348 ; 
        RECT 31.484 214.974 31.588 219.348 ; 
        RECT 31.052 214.974 31.156 219.348 ; 
        RECT 30.62 214.974 30.724 219.348 ; 
        RECT 30.188 214.974 30.292 219.348 ; 
        RECT 29.756 214.974 29.86 219.348 ; 
        RECT 29.324 214.974 29.428 219.348 ; 
        RECT 28.892 214.974 28.996 219.348 ; 
        RECT 28.46 214.974 28.564 219.348 ; 
        RECT 28.028 214.974 28.132 219.348 ; 
        RECT 27.596 214.974 27.7 219.348 ; 
        RECT 27.164 214.974 27.268 219.348 ; 
        RECT 26.732 214.974 26.836 219.348 ; 
        RECT 26.3 214.974 26.404 219.348 ; 
        RECT 25.868 214.974 25.972 219.348 ; 
        RECT 25.436 214.974 25.54 219.348 ; 
        RECT 25.004 214.974 25.108 219.348 ; 
        RECT 24.572 214.974 24.676 219.348 ; 
        RECT 24.14 214.974 24.244 219.348 ; 
        RECT 23.708 214.974 23.812 219.348 ; 
        RECT 22.856 214.974 23.164 219.348 ; 
        RECT 15.284 214.974 15.592 219.348 ; 
        RECT 14.636 214.974 14.74 219.348 ; 
        RECT 14.204 214.974 14.308 219.348 ; 
        RECT 13.772 214.974 13.876 219.348 ; 
        RECT 13.34 214.974 13.444 219.348 ; 
        RECT 12.908 214.974 13.012 219.348 ; 
        RECT 12.476 214.974 12.58 219.348 ; 
        RECT 12.044 214.974 12.148 219.348 ; 
        RECT 11.612 214.974 11.716 219.348 ; 
        RECT 11.18 214.974 11.284 219.348 ; 
        RECT 10.748 214.974 10.852 219.348 ; 
        RECT 10.316 214.974 10.42 219.348 ; 
        RECT 9.884 214.974 9.988 219.348 ; 
        RECT 9.452 214.974 9.556 219.348 ; 
        RECT 9.02 214.974 9.124 219.348 ; 
        RECT 8.588 214.974 8.692 219.348 ; 
        RECT 8.156 214.974 8.26 219.348 ; 
        RECT 7.724 214.974 7.828 219.348 ; 
        RECT 7.292 214.974 7.396 219.348 ; 
        RECT 6.86 214.974 6.964 219.348 ; 
        RECT 6.428 214.974 6.532 219.348 ; 
        RECT 5.996 214.974 6.1 219.348 ; 
        RECT 5.564 214.974 5.668 219.348 ; 
        RECT 5.132 214.974 5.236 219.348 ; 
        RECT 4.7 214.974 4.804 219.348 ; 
        RECT 4.268 214.974 4.372 219.348 ; 
        RECT 3.836 214.974 3.94 219.348 ; 
        RECT 3.404 214.974 3.508 219.348 ; 
        RECT 2.972 214.974 3.076 219.348 ; 
        RECT 2.54 214.974 2.644 219.348 ; 
        RECT 2.108 214.974 2.212 219.348 ; 
        RECT 1.676 214.974 1.78 219.348 ; 
        RECT 1.244 214.974 1.348 219.348 ; 
        RECT 0.812 214.974 0.916 219.348 ; 
        RECT 0 214.974 0.34 219.348 ; 
        RECT 20.72 219.294 21.232 223.668 ; 
        RECT 20.664 221.956 21.232 223.246 ; 
        RECT 20.072 220.864 20.32 223.668 ; 
        RECT 20.016 222.102 20.32 222.716 ; 
        RECT 20.072 219.294 20.176 223.668 ; 
        RECT 20.072 219.778 20.232 220.736 ; 
        RECT 20.072 219.294 20.32 219.65 ; 
        RECT 18.884 221.096 19.708 223.668 ; 
        RECT 19.604 219.294 19.708 223.668 ; 
        RECT 18.884 222.204 19.764 223.236 ; 
        RECT 18.884 219.294 19.276 223.668 ; 
        RECT 17.216 219.294 17.548 223.668 ; 
        RECT 17.216 219.648 17.604 223.39 ; 
        RECT 38.108 219.294 38.448 223.668 ; 
        RECT 37.532 219.294 37.636 223.668 ; 
        RECT 37.1 219.294 37.204 223.668 ; 
        RECT 36.668 219.294 36.772 223.668 ; 
        RECT 36.236 219.294 36.34 223.668 ; 
        RECT 35.804 219.294 35.908 223.668 ; 
        RECT 35.372 219.294 35.476 223.668 ; 
        RECT 34.94 219.294 35.044 223.668 ; 
        RECT 34.508 219.294 34.612 223.668 ; 
        RECT 34.076 219.294 34.18 223.668 ; 
        RECT 33.644 219.294 33.748 223.668 ; 
        RECT 33.212 219.294 33.316 223.668 ; 
        RECT 32.78 219.294 32.884 223.668 ; 
        RECT 32.348 219.294 32.452 223.668 ; 
        RECT 31.916 219.294 32.02 223.668 ; 
        RECT 31.484 219.294 31.588 223.668 ; 
        RECT 31.052 219.294 31.156 223.668 ; 
        RECT 30.62 219.294 30.724 223.668 ; 
        RECT 30.188 219.294 30.292 223.668 ; 
        RECT 29.756 219.294 29.86 223.668 ; 
        RECT 29.324 219.294 29.428 223.668 ; 
        RECT 28.892 219.294 28.996 223.668 ; 
        RECT 28.46 219.294 28.564 223.668 ; 
        RECT 28.028 219.294 28.132 223.668 ; 
        RECT 27.596 219.294 27.7 223.668 ; 
        RECT 27.164 219.294 27.268 223.668 ; 
        RECT 26.732 219.294 26.836 223.668 ; 
        RECT 26.3 219.294 26.404 223.668 ; 
        RECT 25.868 219.294 25.972 223.668 ; 
        RECT 25.436 219.294 25.54 223.668 ; 
        RECT 25.004 219.294 25.108 223.668 ; 
        RECT 24.572 219.294 24.676 223.668 ; 
        RECT 24.14 219.294 24.244 223.668 ; 
        RECT 23.708 219.294 23.812 223.668 ; 
        RECT 22.856 219.294 23.164 223.668 ; 
        RECT 15.284 219.294 15.592 223.668 ; 
        RECT 14.636 219.294 14.74 223.668 ; 
        RECT 14.204 219.294 14.308 223.668 ; 
        RECT 13.772 219.294 13.876 223.668 ; 
        RECT 13.34 219.294 13.444 223.668 ; 
        RECT 12.908 219.294 13.012 223.668 ; 
        RECT 12.476 219.294 12.58 223.668 ; 
        RECT 12.044 219.294 12.148 223.668 ; 
        RECT 11.612 219.294 11.716 223.668 ; 
        RECT 11.18 219.294 11.284 223.668 ; 
        RECT 10.748 219.294 10.852 223.668 ; 
        RECT 10.316 219.294 10.42 223.668 ; 
        RECT 9.884 219.294 9.988 223.668 ; 
        RECT 9.452 219.294 9.556 223.668 ; 
        RECT 9.02 219.294 9.124 223.668 ; 
        RECT 8.588 219.294 8.692 223.668 ; 
        RECT 8.156 219.294 8.26 223.668 ; 
        RECT 7.724 219.294 7.828 223.668 ; 
        RECT 7.292 219.294 7.396 223.668 ; 
        RECT 6.86 219.294 6.964 223.668 ; 
        RECT 6.428 219.294 6.532 223.668 ; 
        RECT 5.996 219.294 6.1 223.668 ; 
        RECT 5.564 219.294 5.668 223.668 ; 
        RECT 5.132 219.294 5.236 223.668 ; 
        RECT 4.7 219.294 4.804 223.668 ; 
        RECT 4.268 219.294 4.372 223.668 ; 
        RECT 3.836 219.294 3.94 223.668 ; 
        RECT 3.404 219.294 3.508 223.668 ; 
        RECT 2.972 219.294 3.076 223.668 ; 
        RECT 2.54 219.294 2.644 223.668 ; 
        RECT 2.108 219.294 2.212 223.668 ; 
        RECT 1.676 219.294 1.78 223.668 ; 
        RECT 1.244 219.294 1.348 223.668 ; 
        RECT 0.812 219.294 0.916 223.668 ; 
        RECT 0 219.294 0.34 223.668 ; 
        RECT 20.72 223.614 21.232 227.988 ; 
        RECT 20.664 226.276 21.232 227.566 ; 
        RECT 20.072 225.184 20.32 227.988 ; 
        RECT 20.016 226.422 20.32 227.036 ; 
        RECT 20.072 223.614 20.176 227.988 ; 
        RECT 20.072 224.098 20.232 225.056 ; 
        RECT 20.072 223.614 20.32 223.97 ; 
        RECT 18.884 225.416 19.708 227.988 ; 
        RECT 19.604 223.614 19.708 227.988 ; 
        RECT 18.884 226.524 19.764 227.556 ; 
        RECT 18.884 223.614 19.276 227.988 ; 
        RECT 17.216 223.614 17.548 227.988 ; 
        RECT 17.216 223.968 17.604 227.71 ; 
        RECT 38.108 223.614 38.448 227.988 ; 
        RECT 37.532 223.614 37.636 227.988 ; 
        RECT 37.1 223.614 37.204 227.988 ; 
        RECT 36.668 223.614 36.772 227.988 ; 
        RECT 36.236 223.614 36.34 227.988 ; 
        RECT 35.804 223.614 35.908 227.988 ; 
        RECT 35.372 223.614 35.476 227.988 ; 
        RECT 34.94 223.614 35.044 227.988 ; 
        RECT 34.508 223.614 34.612 227.988 ; 
        RECT 34.076 223.614 34.18 227.988 ; 
        RECT 33.644 223.614 33.748 227.988 ; 
        RECT 33.212 223.614 33.316 227.988 ; 
        RECT 32.78 223.614 32.884 227.988 ; 
        RECT 32.348 223.614 32.452 227.988 ; 
        RECT 31.916 223.614 32.02 227.988 ; 
        RECT 31.484 223.614 31.588 227.988 ; 
        RECT 31.052 223.614 31.156 227.988 ; 
        RECT 30.62 223.614 30.724 227.988 ; 
        RECT 30.188 223.614 30.292 227.988 ; 
        RECT 29.756 223.614 29.86 227.988 ; 
        RECT 29.324 223.614 29.428 227.988 ; 
        RECT 28.892 223.614 28.996 227.988 ; 
        RECT 28.46 223.614 28.564 227.988 ; 
        RECT 28.028 223.614 28.132 227.988 ; 
        RECT 27.596 223.614 27.7 227.988 ; 
        RECT 27.164 223.614 27.268 227.988 ; 
        RECT 26.732 223.614 26.836 227.988 ; 
        RECT 26.3 223.614 26.404 227.988 ; 
        RECT 25.868 223.614 25.972 227.988 ; 
        RECT 25.436 223.614 25.54 227.988 ; 
        RECT 25.004 223.614 25.108 227.988 ; 
        RECT 24.572 223.614 24.676 227.988 ; 
        RECT 24.14 223.614 24.244 227.988 ; 
        RECT 23.708 223.614 23.812 227.988 ; 
        RECT 22.856 223.614 23.164 227.988 ; 
        RECT 15.284 223.614 15.592 227.988 ; 
        RECT 14.636 223.614 14.74 227.988 ; 
        RECT 14.204 223.614 14.308 227.988 ; 
        RECT 13.772 223.614 13.876 227.988 ; 
        RECT 13.34 223.614 13.444 227.988 ; 
        RECT 12.908 223.614 13.012 227.988 ; 
        RECT 12.476 223.614 12.58 227.988 ; 
        RECT 12.044 223.614 12.148 227.988 ; 
        RECT 11.612 223.614 11.716 227.988 ; 
        RECT 11.18 223.614 11.284 227.988 ; 
        RECT 10.748 223.614 10.852 227.988 ; 
        RECT 10.316 223.614 10.42 227.988 ; 
        RECT 9.884 223.614 9.988 227.988 ; 
        RECT 9.452 223.614 9.556 227.988 ; 
        RECT 9.02 223.614 9.124 227.988 ; 
        RECT 8.588 223.614 8.692 227.988 ; 
        RECT 8.156 223.614 8.26 227.988 ; 
        RECT 7.724 223.614 7.828 227.988 ; 
        RECT 7.292 223.614 7.396 227.988 ; 
        RECT 6.86 223.614 6.964 227.988 ; 
        RECT 6.428 223.614 6.532 227.988 ; 
        RECT 5.996 223.614 6.1 227.988 ; 
        RECT 5.564 223.614 5.668 227.988 ; 
        RECT 5.132 223.614 5.236 227.988 ; 
        RECT 4.7 223.614 4.804 227.988 ; 
        RECT 4.268 223.614 4.372 227.988 ; 
        RECT 3.836 223.614 3.94 227.988 ; 
        RECT 3.404 223.614 3.508 227.988 ; 
        RECT 2.972 223.614 3.076 227.988 ; 
        RECT 2.54 223.614 2.644 227.988 ; 
        RECT 2.108 223.614 2.212 227.988 ; 
        RECT 1.676 223.614 1.78 227.988 ; 
        RECT 1.244 223.614 1.348 227.988 ; 
        RECT 0.812 223.614 0.916 227.988 ; 
        RECT 0 223.614 0.34 227.988 ; 
        RECT 20.72 227.934 21.232 232.308 ; 
        RECT 20.664 230.596 21.232 231.886 ; 
        RECT 20.072 229.504 20.32 232.308 ; 
        RECT 20.016 230.742 20.32 231.356 ; 
        RECT 20.072 227.934 20.176 232.308 ; 
        RECT 20.072 228.418 20.232 229.376 ; 
        RECT 20.072 227.934 20.32 228.29 ; 
        RECT 18.884 229.736 19.708 232.308 ; 
        RECT 19.604 227.934 19.708 232.308 ; 
        RECT 18.884 230.844 19.764 231.876 ; 
        RECT 18.884 227.934 19.276 232.308 ; 
        RECT 17.216 227.934 17.548 232.308 ; 
        RECT 17.216 228.288 17.604 232.03 ; 
        RECT 38.108 227.934 38.448 232.308 ; 
        RECT 37.532 227.934 37.636 232.308 ; 
        RECT 37.1 227.934 37.204 232.308 ; 
        RECT 36.668 227.934 36.772 232.308 ; 
        RECT 36.236 227.934 36.34 232.308 ; 
        RECT 35.804 227.934 35.908 232.308 ; 
        RECT 35.372 227.934 35.476 232.308 ; 
        RECT 34.94 227.934 35.044 232.308 ; 
        RECT 34.508 227.934 34.612 232.308 ; 
        RECT 34.076 227.934 34.18 232.308 ; 
        RECT 33.644 227.934 33.748 232.308 ; 
        RECT 33.212 227.934 33.316 232.308 ; 
        RECT 32.78 227.934 32.884 232.308 ; 
        RECT 32.348 227.934 32.452 232.308 ; 
        RECT 31.916 227.934 32.02 232.308 ; 
        RECT 31.484 227.934 31.588 232.308 ; 
        RECT 31.052 227.934 31.156 232.308 ; 
        RECT 30.62 227.934 30.724 232.308 ; 
        RECT 30.188 227.934 30.292 232.308 ; 
        RECT 29.756 227.934 29.86 232.308 ; 
        RECT 29.324 227.934 29.428 232.308 ; 
        RECT 28.892 227.934 28.996 232.308 ; 
        RECT 28.46 227.934 28.564 232.308 ; 
        RECT 28.028 227.934 28.132 232.308 ; 
        RECT 27.596 227.934 27.7 232.308 ; 
        RECT 27.164 227.934 27.268 232.308 ; 
        RECT 26.732 227.934 26.836 232.308 ; 
        RECT 26.3 227.934 26.404 232.308 ; 
        RECT 25.868 227.934 25.972 232.308 ; 
        RECT 25.436 227.934 25.54 232.308 ; 
        RECT 25.004 227.934 25.108 232.308 ; 
        RECT 24.572 227.934 24.676 232.308 ; 
        RECT 24.14 227.934 24.244 232.308 ; 
        RECT 23.708 227.934 23.812 232.308 ; 
        RECT 22.856 227.934 23.164 232.308 ; 
        RECT 15.284 227.934 15.592 232.308 ; 
        RECT 14.636 227.934 14.74 232.308 ; 
        RECT 14.204 227.934 14.308 232.308 ; 
        RECT 13.772 227.934 13.876 232.308 ; 
        RECT 13.34 227.934 13.444 232.308 ; 
        RECT 12.908 227.934 13.012 232.308 ; 
        RECT 12.476 227.934 12.58 232.308 ; 
        RECT 12.044 227.934 12.148 232.308 ; 
        RECT 11.612 227.934 11.716 232.308 ; 
        RECT 11.18 227.934 11.284 232.308 ; 
        RECT 10.748 227.934 10.852 232.308 ; 
        RECT 10.316 227.934 10.42 232.308 ; 
        RECT 9.884 227.934 9.988 232.308 ; 
        RECT 9.452 227.934 9.556 232.308 ; 
        RECT 9.02 227.934 9.124 232.308 ; 
        RECT 8.588 227.934 8.692 232.308 ; 
        RECT 8.156 227.934 8.26 232.308 ; 
        RECT 7.724 227.934 7.828 232.308 ; 
        RECT 7.292 227.934 7.396 232.308 ; 
        RECT 6.86 227.934 6.964 232.308 ; 
        RECT 6.428 227.934 6.532 232.308 ; 
        RECT 5.996 227.934 6.1 232.308 ; 
        RECT 5.564 227.934 5.668 232.308 ; 
        RECT 5.132 227.934 5.236 232.308 ; 
        RECT 4.7 227.934 4.804 232.308 ; 
        RECT 4.268 227.934 4.372 232.308 ; 
        RECT 3.836 227.934 3.94 232.308 ; 
        RECT 3.404 227.934 3.508 232.308 ; 
        RECT 2.972 227.934 3.076 232.308 ; 
        RECT 2.54 227.934 2.644 232.308 ; 
        RECT 2.108 227.934 2.212 232.308 ; 
        RECT 1.676 227.934 1.78 232.308 ; 
        RECT 1.244 227.934 1.348 232.308 ; 
        RECT 0.812 227.934 0.916 232.308 ; 
        RECT 0 227.934 0.34 232.308 ; 
        RECT 20.72 232.254 21.232 236.628 ; 
        RECT 20.664 234.916 21.232 236.206 ; 
        RECT 20.072 233.824 20.32 236.628 ; 
        RECT 20.016 235.062 20.32 235.676 ; 
        RECT 20.072 232.254 20.176 236.628 ; 
        RECT 20.072 232.738 20.232 233.696 ; 
        RECT 20.072 232.254 20.32 232.61 ; 
        RECT 18.884 234.056 19.708 236.628 ; 
        RECT 19.604 232.254 19.708 236.628 ; 
        RECT 18.884 235.164 19.764 236.196 ; 
        RECT 18.884 232.254 19.276 236.628 ; 
        RECT 17.216 232.254 17.548 236.628 ; 
        RECT 17.216 232.608 17.604 236.35 ; 
        RECT 38.108 232.254 38.448 236.628 ; 
        RECT 37.532 232.254 37.636 236.628 ; 
        RECT 37.1 232.254 37.204 236.628 ; 
        RECT 36.668 232.254 36.772 236.628 ; 
        RECT 36.236 232.254 36.34 236.628 ; 
        RECT 35.804 232.254 35.908 236.628 ; 
        RECT 35.372 232.254 35.476 236.628 ; 
        RECT 34.94 232.254 35.044 236.628 ; 
        RECT 34.508 232.254 34.612 236.628 ; 
        RECT 34.076 232.254 34.18 236.628 ; 
        RECT 33.644 232.254 33.748 236.628 ; 
        RECT 33.212 232.254 33.316 236.628 ; 
        RECT 32.78 232.254 32.884 236.628 ; 
        RECT 32.348 232.254 32.452 236.628 ; 
        RECT 31.916 232.254 32.02 236.628 ; 
        RECT 31.484 232.254 31.588 236.628 ; 
        RECT 31.052 232.254 31.156 236.628 ; 
        RECT 30.62 232.254 30.724 236.628 ; 
        RECT 30.188 232.254 30.292 236.628 ; 
        RECT 29.756 232.254 29.86 236.628 ; 
        RECT 29.324 232.254 29.428 236.628 ; 
        RECT 28.892 232.254 28.996 236.628 ; 
        RECT 28.46 232.254 28.564 236.628 ; 
        RECT 28.028 232.254 28.132 236.628 ; 
        RECT 27.596 232.254 27.7 236.628 ; 
        RECT 27.164 232.254 27.268 236.628 ; 
        RECT 26.732 232.254 26.836 236.628 ; 
        RECT 26.3 232.254 26.404 236.628 ; 
        RECT 25.868 232.254 25.972 236.628 ; 
        RECT 25.436 232.254 25.54 236.628 ; 
        RECT 25.004 232.254 25.108 236.628 ; 
        RECT 24.572 232.254 24.676 236.628 ; 
        RECT 24.14 232.254 24.244 236.628 ; 
        RECT 23.708 232.254 23.812 236.628 ; 
        RECT 22.856 232.254 23.164 236.628 ; 
        RECT 15.284 232.254 15.592 236.628 ; 
        RECT 14.636 232.254 14.74 236.628 ; 
        RECT 14.204 232.254 14.308 236.628 ; 
        RECT 13.772 232.254 13.876 236.628 ; 
        RECT 13.34 232.254 13.444 236.628 ; 
        RECT 12.908 232.254 13.012 236.628 ; 
        RECT 12.476 232.254 12.58 236.628 ; 
        RECT 12.044 232.254 12.148 236.628 ; 
        RECT 11.612 232.254 11.716 236.628 ; 
        RECT 11.18 232.254 11.284 236.628 ; 
        RECT 10.748 232.254 10.852 236.628 ; 
        RECT 10.316 232.254 10.42 236.628 ; 
        RECT 9.884 232.254 9.988 236.628 ; 
        RECT 9.452 232.254 9.556 236.628 ; 
        RECT 9.02 232.254 9.124 236.628 ; 
        RECT 8.588 232.254 8.692 236.628 ; 
        RECT 8.156 232.254 8.26 236.628 ; 
        RECT 7.724 232.254 7.828 236.628 ; 
        RECT 7.292 232.254 7.396 236.628 ; 
        RECT 6.86 232.254 6.964 236.628 ; 
        RECT 6.428 232.254 6.532 236.628 ; 
        RECT 5.996 232.254 6.1 236.628 ; 
        RECT 5.564 232.254 5.668 236.628 ; 
        RECT 5.132 232.254 5.236 236.628 ; 
        RECT 4.7 232.254 4.804 236.628 ; 
        RECT 4.268 232.254 4.372 236.628 ; 
        RECT 3.836 232.254 3.94 236.628 ; 
        RECT 3.404 232.254 3.508 236.628 ; 
        RECT 2.972 232.254 3.076 236.628 ; 
        RECT 2.54 232.254 2.644 236.628 ; 
        RECT 2.108 232.254 2.212 236.628 ; 
        RECT 1.676 232.254 1.78 236.628 ; 
        RECT 1.244 232.254 1.348 236.628 ; 
        RECT 0.812 232.254 0.916 236.628 ; 
        RECT 0 232.254 0.34 236.628 ; 
        RECT 20.72 236.574 21.232 240.948 ; 
        RECT 20.664 239.236 21.232 240.526 ; 
        RECT 20.072 238.144 20.32 240.948 ; 
        RECT 20.016 239.382 20.32 239.996 ; 
        RECT 20.072 236.574 20.176 240.948 ; 
        RECT 20.072 237.058 20.232 238.016 ; 
        RECT 20.072 236.574 20.32 236.93 ; 
        RECT 18.884 238.376 19.708 240.948 ; 
        RECT 19.604 236.574 19.708 240.948 ; 
        RECT 18.884 239.484 19.764 240.516 ; 
        RECT 18.884 236.574 19.276 240.948 ; 
        RECT 17.216 236.574 17.548 240.948 ; 
        RECT 17.216 236.928 17.604 240.67 ; 
        RECT 38.108 236.574 38.448 240.948 ; 
        RECT 37.532 236.574 37.636 240.948 ; 
        RECT 37.1 236.574 37.204 240.948 ; 
        RECT 36.668 236.574 36.772 240.948 ; 
        RECT 36.236 236.574 36.34 240.948 ; 
        RECT 35.804 236.574 35.908 240.948 ; 
        RECT 35.372 236.574 35.476 240.948 ; 
        RECT 34.94 236.574 35.044 240.948 ; 
        RECT 34.508 236.574 34.612 240.948 ; 
        RECT 34.076 236.574 34.18 240.948 ; 
        RECT 33.644 236.574 33.748 240.948 ; 
        RECT 33.212 236.574 33.316 240.948 ; 
        RECT 32.78 236.574 32.884 240.948 ; 
        RECT 32.348 236.574 32.452 240.948 ; 
        RECT 31.916 236.574 32.02 240.948 ; 
        RECT 31.484 236.574 31.588 240.948 ; 
        RECT 31.052 236.574 31.156 240.948 ; 
        RECT 30.62 236.574 30.724 240.948 ; 
        RECT 30.188 236.574 30.292 240.948 ; 
        RECT 29.756 236.574 29.86 240.948 ; 
        RECT 29.324 236.574 29.428 240.948 ; 
        RECT 28.892 236.574 28.996 240.948 ; 
        RECT 28.46 236.574 28.564 240.948 ; 
        RECT 28.028 236.574 28.132 240.948 ; 
        RECT 27.596 236.574 27.7 240.948 ; 
        RECT 27.164 236.574 27.268 240.948 ; 
        RECT 26.732 236.574 26.836 240.948 ; 
        RECT 26.3 236.574 26.404 240.948 ; 
        RECT 25.868 236.574 25.972 240.948 ; 
        RECT 25.436 236.574 25.54 240.948 ; 
        RECT 25.004 236.574 25.108 240.948 ; 
        RECT 24.572 236.574 24.676 240.948 ; 
        RECT 24.14 236.574 24.244 240.948 ; 
        RECT 23.708 236.574 23.812 240.948 ; 
        RECT 22.856 236.574 23.164 240.948 ; 
        RECT 15.284 236.574 15.592 240.948 ; 
        RECT 14.636 236.574 14.74 240.948 ; 
        RECT 14.204 236.574 14.308 240.948 ; 
        RECT 13.772 236.574 13.876 240.948 ; 
        RECT 13.34 236.574 13.444 240.948 ; 
        RECT 12.908 236.574 13.012 240.948 ; 
        RECT 12.476 236.574 12.58 240.948 ; 
        RECT 12.044 236.574 12.148 240.948 ; 
        RECT 11.612 236.574 11.716 240.948 ; 
        RECT 11.18 236.574 11.284 240.948 ; 
        RECT 10.748 236.574 10.852 240.948 ; 
        RECT 10.316 236.574 10.42 240.948 ; 
        RECT 9.884 236.574 9.988 240.948 ; 
        RECT 9.452 236.574 9.556 240.948 ; 
        RECT 9.02 236.574 9.124 240.948 ; 
        RECT 8.588 236.574 8.692 240.948 ; 
        RECT 8.156 236.574 8.26 240.948 ; 
        RECT 7.724 236.574 7.828 240.948 ; 
        RECT 7.292 236.574 7.396 240.948 ; 
        RECT 6.86 236.574 6.964 240.948 ; 
        RECT 6.428 236.574 6.532 240.948 ; 
        RECT 5.996 236.574 6.1 240.948 ; 
        RECT 5.564 236.574 5.668 240.948 ; 
        RECT 5.132 236.574 5.236 240.948 ; 
        RECT 4.7 236.574 4.804 240.948 ; 
        RECT 4.268 236.574 4.372 240.948 ; 
        RECT 3.836 236.574 3.94 240.948 ; 
        RECT 3.404 236.574 3.508 240.948 ; 
        RECT 2.972 236.574 3.076 240.948 ; 
        RECT 2.54 236.574 2.644 240.948 ; 
        RECT 2.108 236.574 2.212 240.948 ; 
        RECT 1.676 236.574 1.78 240.948 ; 
        RECT 1.244 236.574 1.348 240.948 ; 
        RECT 0.812 236.574 0.916 240.948 ; 
        RECT 0 236.574 0.34 240.948 ; 
  LAYER V3 ; 
      RECT 0 4.88 38.448 5.4 ; 
      RECT 37.98 1.026 38.448 5.4 ; 
      RECT 23.364 4.496 37.908 5.4 ; 
      RECT 18.036 4.496 23.292 5.4 ; 
      RECT 15.156 1.026 17.676 5.4 ; 
      RECT 0.54 4.496 15.084 5.4 ; 
      RECT 0 1.026 0.468 5.4 ; 
      RECT 37.836 1.026 38.448 4.688 ; 
      RECT 23.58 1.026 37.764 5.4 ; 
      RECT 20.592 1.026 23.508 4.688 ; 
      RECT 19.944 1.808 20.448 5.4 ; 
      RECT 14.94 1.424 19.836 4.688 ; 
      RECT 0.684 1.026 14.868 5.4 ; 
      RECT 0 1.026 0.612 4.688 ; 
      RECT 20.376 1.026 38.448 4.304 ; 
      RECT 0 1.424 20.304 4.304 ; 
      RECT 19.476 1.026 38.448 1.712 ; 
      RECT 0 1.026 19.404 4.304 ; 
      RECT 0 1.026 38.448 1.328 ; 
      RECT 0 9.2 38.448 9.72 ; 
      RECT 37.98 5.346 38.448 9.72 ; 
      RECT 23.364 8.816 37.908 9.72 ; 
      RECT 18.036 8.816 23.292 9.72 ; 
      RECT 15.156 5.346 17.676 9.72 ; 
      RECT 0.54 8.816 15.084 9.72 ; 
      RECT 0 5.346 0.468 9.72 ; 
      RECT 37.836 5.346 38.448 9.008 ; 
      RECT 23.58 5.346 37.764 9.72 ; 
      RECT 20.592 5.346 23.508 9.008 ; 
      RECT 19.944 6.128 20.448 9.72 ; 
      RECT 14.94 5.744 19.836 9.008 ; 
      RECT 0.684 5.346 14.868 9.72 ; 
      RECT 0 5.346 0.612 9.008 ; 
      RECT 20.376 5.346 38.448 8.624 ; 
      RECT 0 5.744 20.304 8.624 ; 
      RECT 19.476 5.346 38.448 6.032 ; 
      RECT 0 5.346 19.404 8.624 ; 
      RECT 0 5.346 38.448 5.648 ; 
      RECT 0 13.52 38.448 14.04 ; 
      RECT 37.98 9.666 38.448 14.04 ; 
      RECT 23.364 13.136 37.908 14.04 ; 
      RECT 18.036 13.136 23.292 14.04 ; 
      RECT 15.156 9.666 17.676 14.04 ; 
      RECT 0.54 13.136 15.084 14.04 ; 
      RECT 0 9.666 0.468 14.04 ; 
      RECT 37.836 9.666 38.448 13.328 ; 
      RECT 23.58 9.666 37.764 14.04 ; 
      RECT 20.592 9.666 23.508 13.328 ; 
      RECT 19.944 10.448 20.448 14.04 ; 
      RECT 14.94 10.064 19.836 13.328 ; 
      RECT 0.684 9.666 14.868 14.04 ; 
      RECT 0 9.666 0.612 13.328 ; 
      RECT 20.376 9.666 38.448 12.944 ; 
      RECT 0 10.064 20.304 12.944 ; 
      RECT 19.476 9.666 38.448 10.352 ; 
      RECT 0 9.666 19.404 12.944 ; 
      RECT 0 9.666 38.448 9.968 ; 
      RECT 0 17.84 38.448 18.36 ; 
      RECT 37.98 13.986 38.448 18.36 ; 
      RECT 23.364 17.456 37.908 18.36 ; 
      RECT 18.036 17.456 23.292 18.36 ; 
      RECT 15.156 13.986 17.676 18.36 ; 
      RECT 0.54 17.456 15.084 18.36 ; 
      RECT 0 13.986 0.468 18.36 ; 
      RECT 37.836 13.986 38.448 17.648 ; 
      RECT 23.58 13.986 37.764 18.36 ; 
      RECT 20.592 13.986 23.508 17.648 ; 
      RECT 19.944 14.768 20.448 18.36 ; 
      RECT 14.94 14.384 19.836 17.648 ; 
      RECT 0.684 13.986 14.868 18.36 ; 
      RECT 0 13.986 0.612 17.648 ; 
      RECT 20.376 13.986 38.448 17.264 ; 
      RECT 0 14.384 20.304 17.264 ; 
      RECT 19.476 13.986 38.448 14.672 ; 
      RECT 0 13.986 19.404 17.264 ; 
      RECT 0 13.986 38.448 14.288 ; 
      RECT 0 22.16 38.448 22.68 ; 
      RECT 37.98 18.306 38.448 22.68 ; 
      RECT 23.364 21.776 37.908 22.68 ; 
      RECT 18.036 21.776 23.292 22.68 ; 
      RECT 15.156 18.306 17.676 22.68 ; 
      RECT 0.54 21.776 15.084 22.68 ; 
      RECT 0 18.306 0.468 22.68 ; 
      RECT 37.836 18.306 38.448 21.968 ; 
      RECT 23.58 18.306 37.764 22.68 ; 
      RECT 20.592 18.306 23.508 21.968 ; 
      RECT 19.944 19.088 20.448 22.68 ; 
      RECT 14.94 18.704 19.836 21.968 ; 
      RECT 0.684 18.306 14.868 22.68 ; 
      RECT 0 18.306 0.612 21.968 ; 
      RECT 20.376 18.306 38.448 21.584 ; 
      RECT 0 18.704 20.304 21.584 ; 
      RECT 19.476 18.306 38.448 18.992 ; 
      RECT 0 18.306 19.404 21.584 ; 
      RECT 0 18.306 38.448 18.608 ; 
      RECT 0 26.48 38.448 27 ; 
      RECT 37.98 22.626 38.448 27 ; 
      RECT 23.364 26.096 37.908 27 ; 
      RECT 18.036 26.096 23.292 27 ; 
      RECT 15.156 22.626 17.676 27 ; 
      RECT 0.54 26.096 15.084 27 ; 
      RECT 0 22.626 0.468 27 ; 
      RECT 37.836 22.626 38.448 26.288 ; 
      RECT 23.58 22.626 37.764 27 ; 
      RECT 20.592 22.626 23.508 26.288 ; 
      RECT 19.944 23.408 20.448 27 ; 
      RECT 14.94 23.024 19.836 26.288 ; 
      RECT 0.684 22.626 14.868 27 ; 
      RECT 0 22.626 0.612 26.288 ; 
      RECT 20.376 22.626 38.448 25.904 ; 
      RECT 0 23.024 20.304 25.904 ; 
      RECT 19.476 22.626 38.448 23.312 ; 
      RECT 0 22.626 19.404 25.904 ; 
      RECT 0 22.626 38.448 22.928 ; 
      RECT 0 30.8 38.448 31.32 ; 
      RECT 37.98 26.946 38.448 31.32 ; 
      RECT 23.364 30.416 37.908 31.32 ; 
      RECT 18.036 30.416 23.292 31.32 ; 
      RECT 15.156 26.946 17.676 31.32 ; 
      RECT 0.54 30.416 15.084 31.32 ; 
      RECT 0 26.946 0.468 31.32 ; 
      RECT 37.836 26.946 38.448 30.608 ; 
      RECT 23.58 26.946 37.764 31.32 ; 
      RECT 20.592 26.946 23.508 30.608 ; 
      RECT 19.944 27.728 20.448 31.32 ; 
      RECT 14.94 27.344 19.836 30.608 ; 
      RECT 0.684 26.946 14.868 31.32 ; 
      RECT 0 26.946 0.612 30.608 ; 
      RECT 20.376 26.946 38.448 30.224 ; 
      RECT 0 27.344 20.304 30.224 ; 
      RECT 19.476 26.946 38.448 27.632 ; 
      RECT 0 26.946 19.404 30.224 ; 
      RECT 0 26.946 38.448 27.248 ; 
      RECT 0 35.12 38.448 35.64 ; 
      RECT 37.98 31.266 38.448 35.64 ; 
      RECT 23.364 34.736 37.908 35.64 ; 
      RECT 18.036 34.736 23.292 35.64 ; 
      RECT 15.156 31.266 17.676 35.64 ; 
      RECT 0.54 34.736 15.084 35.64 ; 
      RECT 0 31.266 0.468 35.64 ; 
      RECT 37.836 31.266 38.448 34.928 ; 
      RECT 23.58 31.266 37.764 35.64 ; 
      RECT 20.592 31.266 23.508 34.928 ; 
      RECT 19.944 32.048 20.448 35.64 ; 
      RECT 14.94 31.664 19.836 34.928 ; 
      RECT 0.684 31.266 14.868 35.64 ; 
      RECT 0 31.266 0.612 34.928 ; 
      RECT 20.376 31.266 38.448 34.544 ; 
      RECT 0 31.664 20.304 34.544 ; 
      RECT 19.476 31.266 38.448 31.952 ; 
      RECT 0 31.266 19.404 34.544 ; 
      RECT 0 31.266 38.448 31.568 ; 
      RECT 0 39.44 38.448 39.96 ; 
      RECT 37.98 35.586 38.448 39.96 ; 
      RECT 23.364 39.056 37.908 39.96 ; 
      RECT 18.036 39.056 23.292 39.96 ; 
      RECT 15.156 35.586 17.676 39.96 ; 
      RECT 0.54 39.056 15.084 39.96 ; 
      RECT 0 35.586 0.468 39.96 ; 
      RECT 37.836 35.586 38.448 39.248 ; 
      RECT 23.58 35.586 37.764 39.96 ; 
      RECT 20.592 35.586 23.508 39.248 ; 
      RECT 19.944 36.368 20.448 39.96 ; 
      RECT 14.94 35.984 19.836 39.248 ; 
      RECT 0.684 35.586 14.868 39.96 ; 
      RECT 0 35.586 0.612 39.248 ; 
      RECT 20.376 35.586 38.448 38.864 ; 
      RECT 0 35.984 20.304 38.864 ; 
      RECT 19.476 35.586 38.448 36.272 ; 
      RECT 0 35.586 19.404 38.864 ; 
      RECT 0 35.586 38.448 35.888 ; 
      RECT 0 43.76 38.448 44.28 ; 
      RECT 37.98 39.906 38.448 44.28 ; 
      RECT 23.364 43.376 37.908 44.28 ; 
      RECT 18.036 43.376 23.292 44.28 ; 
      RECT 15.156 39.906 17.676 44.28 ; 
      RECT 0.54 43.376 15.084 44.28 ; 
      RECT 0 39.906 0.468 44.28 ; 
      RECT 37.836 39.906 38.448 43.568 ; 
      RECT 23.58 39.906 37.764 44.28 ; 
      RECT 20.592 39.906 23.508 43.568 ; 
      RECT 19.944 40.688 20.448 44.28 ; 
      RECT 14.94 40.304 19.836 43.568 ; 
      RECT 0.684 39.906 14.868 44.28 ; 
      RECT 0 39.906 0.612 43.568 ; 
      RECT 20.376 39.906 38.448 43.184 ; 
      RECT 0 40.304 20.304 43.184 ; 
      RECT 19.476 39.906 38.448 40.592 ; 
      RECT 0 39.906 19.404 43.184 ; 
      RECT 0 39.906 38.448 40.208 ; 
      RECT 0 48.08 38.448 48.6 ; 
      RECT 37.98 44.226 38.448 48.6 ; 
      RECT 23.364 47.696 37.908 48.6 ; 
      RECT 18.036 47.696 23.292 48.6 ; 
      RECT 15.156 44.226 17.676 48.6 ; 
      RECT 0.54 47.696 15.084 48.6 ; 
      RECT 0 44.226 0.468 48.6 ; 
      RECT 37.836 44.226 38.448 47.888 ; 
      RECT 23.58 44.226 37.764 48.6 ; 
      RECT 20.592 44.226 23.508 47.888 ; 
      RECT 19.944 45.008 20.448 48.6 ; 
      RECT 14.94 44.624 19.836 47.888 ; 
      RECT 0.684 44.226 14.868 48.6 ; 
      RECT 0 44.226 0.612 47.888 ; 
      RECT 20.376 44.226 38.448 47.504 ; 
      RECT 0 44.624 20.304 47.504 ; 
      RECT 19.476 44.226 38.448 44.912 ; 
      RECT 0 44.226 19.404 47.504 ; 
      RECT 0 44.226 38.448 44.528 ; 
      RECT 0 52.4 38.448 52.92 ; 
      RECT 37.98 48.546 38.448 52.92 ; 
      RECT 23.364 52.016 37.908 52.92 ; 
      RECT 18.036 52.016 23.292 52.92 ; 
      RECT 15.156 48.546 17.676 52.92 ; 
      RECT 0.54 52.016 15.084 52.92 ; 
      RECT 0 48.546 0.468 52.92 ; 
      RECT 37.836 48.546 38.448 52.208 ; 
      RECT 23.58 48.546 37.764 52.92 ; 
      RECT 20.592 48.546 23.508 52.208 ; 
      RECT 19.944 49.328 20.448 52.92 ; 
      RECT 14.94 48.944 19.836 52.208 ; 
      RECT 0.684 48.546 14.868 52.92 ; 
      RECT 0 48.546 0.612 52.208 ; 
      RECT 20.376 48.546 38.448 51.824 ; 
      RECT 0 48.944 20.304 51.824 ; 
      RECT 19.476 48.546 38.448 49.232 ; 
      RECT 0 48.546 19.404 51.824 ; 
      RECT 0 48.546 38.448 48.848 ; 
      RECT 0 56.72 38.448 57.24 ; 
      RECT 37.98 52.866 38.448 57.24 ; 
      RECT 23.364 56.336 37.908 57.24 ; 
      RECT 18.036 56.336 23.292 57.24 ; 
      RECT 15.156 52.866 17.676 57.24 ; 
      RECT 0.54 56.336 15.084 57.24 ; 
      RECT 0 52.866 0.468 57.24 ; 
      RECT 37.836 52.866 38.448 56.528 ; 
      RECT 23.58 52.866 37.764 57.24 ; 
      RECT 20.592 52.866 23.508 56.528 ; 
      RECT 19.944 53.648 20.448 57.24 ; 
      RECT 14.94 53.264 19.836 56.528 ; 
      RECT 0.684 52.866 14.868 57.24 ; 
      RECT 0 52.866 0.612 56.528 ; 
      RECT 20.376 52.866 38.448 56.144 ; 
      RECT 0 53.264 20.304 56.144 ; 
      RECT 19.476 52.866 38.448 53.552 ; 
      RECT 0 52.866 19.404 56.144 ; 
      RECT 0 52.866 38.448 53.168 ; 
      RECT 0 61.04 38.448 61.56 ; 
      RECT 37.98 57.186 38.448 61.56 ; 
      RECT 23.364 60.656 37.908 61.56 ; 
      RECT 18.036 60.656 23.292 61.56 ; 
      RECT 15.156 57.186 17.676 61.56 ; 
      RECT 0.54 60.656 15.084 61.56 ; 
      RECT 0 57.186 0.468 61.56 ; 
      RECT 37.836 57.186 38.448 60.848 ; 
      RECT 23.58 57.186 37.764 61.56 ; 
      RECT 20.592 57.186 23.508 60.848 ; 
      RECT 19.944 57.968 20.448 61.56 ; 
      RECT 14.94 57.584 19.836 60.848 ; 
      RECT 0.684 57.186 14.868 61.56 ; 
      RECT 0 57.186 0.612 60.848 ; 
      RECT 20.376 57.186 38.448 60.464 ; 
      RECT 0 57.584 20.304 60.464 ; 
      RECT 19.476 57.186 38.448 57.872 ; 
      RECT 0 57.186 19.404 60.464 ; 
      RECT 0 57.186 38.448 57.488 ; 
      RECT 0 65.36 38.448 65.88 ; 
      RECT 37.98 61.506 38.448 65.88 ; 
      RECT 23.364 64.976 37.908 65.88 ; 
      RECT 18.036 64.976 23.292 65.88 ; 
      RECT 15.156 61.506 17.676 65.88 ; 
      RECT 0.54 64.976 15.084 65.88 ; 
      RECT 0 61.506 0.468 65.88 ; 
      RECT 37.836 61.506 38.448 65.168 ; 
      RECT 23.58 61.506 37.764 65.88 ; 
      RECT 20.592 61.506 23.508 65.168 ; 
      RECT 19.944 62.288 20.448 65.88 ; 
      RECT 14.94 61.904 19.836 65.168 ; 
      RECT 0.684 61.506 14.868 65.88 ; 
      RECT 0 61.506 0.612 65.168 ; 
      RECT 20.376 61.506 38.448 64.784 ; 
      RECT 0 61.904 20.304 64.784 ; 
      RECT 19.476 61.506 38.448 62.192 ; 
      RECT 0 61.506 19.404 64.784 ; 
      RECT 0 61.506 38.448 61.808 ; 
      RECT 0 69.68 38.448 70.2 ; 
      RECT 37.98 65.826 38.448 70.2 ; 
      RECT 23.364 69.296 37.908 70.2 ; 
      RECT 18.036 69.296 23.292 70.2 ; 
      RECT 15.156 65.826 17.676 70.2 ; 
      RECT 0.54 69.296 15.084 70.2 ; 
      RECT 0 65.826 0.468 70.2 ; 
      RECT 37.836 65.826 38.448 69.488 ; 
      RECT 23.58 65.826 37.764 70.2 ; 
      RECT 20.592 65.826 23.508 69.488 ; 
      RECT 19.944 66.608 20.448 70.2 ; 
      RECT 14.94 66.224 19.836 69.488 ; 
      RECT 0.684 65.826 14.868 70.2 ; 
      RECT 0 65.826 0.612 69.488 ; 
      RECT 20.376 65.826 38.448 69.104 ; 
      RECT 0 66.224 20.304 69.104 ; 
      RECT 19.476 65.826 38.448 66.512 ; 
      RECT 0 65.826 19.404 69.104 ; 
      RECT 0 65.826 38.448 66.128 ; 
      RECT 0 74 38.448 74.52 ; 
      RECT 37.98 70.146 38.448 74.52 ; 
      RECT 23.364 73.616 37.908 74.52 ; 
      RECT 18.036 73.616 23.292 74.52 ; 
      RECT 15.156 70.146 17.676 74.52 ; 
      RECT 0.54 73.616 15.084 74.52 ; 
      RECT 0 70.146 0.468 74.52 ; 
      RECT 37.836 70.146 38.448 73.808 ; 
      RECT 23.58 70.146 37.764 74.52 ; 
      RECT 20.592 70.146 23.508 73.808 ; 
      RECT 19.944 70.928 20.448 74.52 ; 
      RECT 14.94 70.544 19.836 73.808 ; 
      RECT 0.684 70.146 14.868 74.52 ; 
      RECT 0 70.146 0.612 73.808 ; 
      RECT 20.376 70.146 38.448 73.424 ; 
      RECT 0 70.544 20.304 73.424 ; 
      RECT 19.476 70.146 38.448 70.832 ; 
      RECT 0 70.146 19.404 73.424 ; 
      RECT 0 70.146 38.448 70.448 ; 
      RECT 0 78.32 38.448 78.84 ; 
      RECT 37.98 74.466 38.448 78.84 ; 
      RECT 23.364 77.936 37.908 78.84 ; 
      RECT 18.036 77.936 23.292 78.84 ; 
      RECT 15.156 74.466 17.676 78.84 ; 
      RECT 0.54 77.936 15.084 78.84 ; 
      RECT 0 74.466 0.468 78.84 ; 
      RECT 37.836 74.466 38.448 78.128 ; 
      RECT 23.58 74.466 37.764 78.84 ; 
      RECT 20.592 74.466 23.508 78.128 ; 
      RECT 19.944 75.248 20.448 78.84 ; 
      RECT 14.94 74.864 19.836 78.128 ; 
      RECT 0.684 74.466 14.868 78.84 ; 
      RECT 0 74.466 0.612 78.128 ; 
      RECT 20.376 74.466 38.448 77.744 ; 
      RECT 0 74.864 20.304 77.744 ; 
      RECT 19.476 74.466 38.448 75.152 ; 
      RECT 0 74.466 19.404 77.744 ; 
      RECT 0 74.466 38.448 74.768 ; 
      RECT 0 82.64 38.448 83.16 ; 
      RECT 37.98 78.786 38.448 83.16 ; 
      RECT 23.364 82.256 37.908 83.16 ; 
      RECT 18.036 82.256 23.292 83.16 ; 
      RECT 15.156 78.786 17.676 83.16 ; 
      RECT 0.54 82.256 15.084 83.16 ; 
      RECT 0 78.786 0.468 83.16 ; 
      RECT 37.836 78.786 38.448 82.448 ; 
      RECT 23.58 78.786 37.764 83.16 ; 
      RECT 20.592 78.786 23.508 82.448 ; 
      RECT 19.944 79.568 20.448 83.16 ; 
      RECT 14.94 79.184 19.836 82.448 ; 
      RECT 0.684 78.786 14.868 83.16 ; 
      RECT 0 78.786 0.612 82.448 ; 
      RECT 20.376 78.786 38.448 82.064 ; 
      RECT 0 79.184 20.304 82.064 ; 
      RECT 19.476 78.786 38.448 79.472 ; 
      RECT 0 78.786 19.404 82.064 ; 
      RECT 0 78.786 38.448 79.088 ; 
      RECT 0 86.96 38.448 87.48 ; 
      RECT 37.98 83.106 38.448 87.48 ; 
      RECT 23.364 86.576 37.908 87.48 ; 
      RECT 18.036 86.576 23.292 87.48 ; 
      RECT 15.156 83.106 17.676 87.48 ; 
      RECT 0.54 86.576 15.084 87.48 ; 
      RECT 0 83.106 0.468 87.48 ; 
      RECT 37.836 83.106 38.448 86.768 ; 
      RECT 23.58 83.106 37.764 87.48 ; 
      RECT 20.592 83.106 23.508 86.768 ; 
      RECT 19.944 83.888 20.448 87.48 ; 
      RECT 14.94 83.504 19.836 86.768 ; 
      RECT 0.684 83.106 14.868 87.48 ; 
      RECT 0 83.106 0.612 86.768 ; 
      RECT 20.376 83.106 38.448 86.384 ; 
      RECT 0 83.504 20.304 86.384 ; 
      RECT 19.476 83.106 38.448 83.792 ; 
      RECT 0 83.106 19.404 86.384 ; 
      RECT 0 83.106 38.448 83.408 ; 
      RECT 0 91.28 38.448 91.8 ; 
      RECT 37.98 87.426 38.448 91.8 ; 
      RECT 23.364 90.896 37.908 91.8 ; 
      RECT 18.036 90.896 23.292 91.8 ; 
      RECT 15.156 87.426 17.676 91.8 ; 
      RECT 0.54 90.896 15.084 91.8 ; 
      RECT 0 87.426 0.468 91.8 ; 
      RECT 37.836 87.426 38.448 91.088 ; 
      RECT 23.58 87.426 37.764 91.8 ; 
      RECT 20.592 87.426 23.508 91.088 ; 
      RECT 19.944 88.208 20.448 91.8 ; 
      RECT 14.94 87.824 19.836 91.088 ; 
      RECT 0.684 87.426 14.868 91.8 ; 
      RECT 0 87.426 0.612 91.088 ; 
      RECT 20.376 87.426 38.448 90.704 ; 
      RECT 0 87.824 20.304 90.704 ; 
      RECT 19.476 87.426 38.448 88.112 ; 
      RECT 0 87.426 19.404 90.704 ; 
      RECT 0 87.426 38.448 87.728 ; 
      RECT 0 95.6 38.448 96.12 ; 
      RECT 37.98 91.746 38.448 96.12 ; 
      RECT 23.364 95.216 37.908 96.12 ; 
      RECT 18.036 95.216 23.292 96.12 ; 
      RECT 15.156 91.746 17.676 96.12 ; 
      RECT 0.54 95.216 15.084 96.12 ; 
      RECT 0 91.746 0.468 96.12 ; 
      RECT 37.836 91.746 38.448 95.408 ; 
      RECT 23.58 91.746 37.764 96.12 ; 
      RECT 20.592 91.746 23.508 95.408 ; 
      RECT 19.944 92.528 20.448 96.12 ; 
      RECT 14.94 92.144 19.836 95.408 ; 
      RECT 0.684 91.746 14.868 96.12 ; 
      RECT 0 91.746 0.612 95.408 ; 
      RECT 20.376 91.746 38.448 95.024 ; 
      RECT 0 92.144 20.304 95.024 ; 
      RECT 19.476 91.746 38.448 92.432 ; 
      RECT 0 91.746 19.404 95.024 ; 
      RECT 0 91.746 38.448 92.048 ; 
      RECT 0 99.92 38.448 100.44 ; 
      RECT 37.98 96.066 38.448 100.44 ; 
      RECT 23.364 99.536 37.908 100.44 ; 
      RECT 18.036 99.536 23.292 100.44 ; 
      RECT 15.156 96.066 17.676 100.44 ; 
      RECT 0.54 99.536 15.084 100.44 ; 
      RECT 0 96.066 0.468 100.44 ; 
      RECT 37.836 96.066 38.448 99.728 ; 
      RECT 23.58 96.066 37.764 100.44 ; 
      RECT 20.592 96.066 23.508 99.728 ; 
      RECT 19.944 96.848 20.448 100.44 ; 
      RECT 14.94 96.464 19.836 99.728 ; 
      RECT 0.684 96.066 14.868 100.44 ; 
      RECT 0 96.066 0.612 99.728 ; 
      RECT 20.376 96.066 38.448 99.344 ; 
      RECT 0 96.464 20.304 99.344 ; 
      RECT 19.476 96.066 38.448 96.752 ; 
      RECT 0 96.066 19.404 99.344 ; 
      RECT 0 96.066 38.448 96.368 ; 
      RECT 0 104.24 38.448 104.76 ; 
      RECT 37.98 100.386 38.448 104.76 ; 
      RECT 23.364 103.856 37.908 104.76 ; 
      RECT 18.036 103.856 23.292 104.76 ; 
      RECT 15.156 100.386 17.676 104.76 ; 
      RECT 0.54 103.856 15.084 104.76 ; 
      RECT 0 100.386 0.468 104.76 ; 
      RECT 37.836 100.386 38.448 104.048 ; 
      RECT 23.58 100.386 37.764 104.76 ; 
      RECT 20.592 100.386 23.508 104.048 ; 
      RECT 19.944 101.168 20.448 104.76 ; 
      RECT 14.94 100.784 19.836 104.048 ; 
      RECT 0.684 100.386 14.868 104.76 ; 
      RECT 0 100.386 0.612 104.048 ; 
      RECT 20.376 100.386 38.448 103.664 ; 
      RECT 0 100.784 20.304 103.664 ; 
      RECT 19.476 100.386 38.448 101.072 ; 
      RECT 0 100.386 19.404 103.664 ; 
      RECT 0 100.386 38.448 100.688 ; 
      RECT 0 133.932 38.448 139.266 ; 
      RECT 29.412 104.652 38.448 139.266 ; 
      RECT 20.612 120.108 38.448 139.266 ; 
      RECT 24.228 109.74 38.448 139.266 ; 
      RECT 20.404 104.652 20.54 139.266 ; 
      RECT 20.196 104.652 20.332 139.266 ; 
      RECT 19.988 104.652 20.124 139.266 ; 
      RECT 19.78 104.652 19.916 139.266 ; 
      RECT 0 132.204 19.708 139.266 ; 
      RECT 18.74 121.26 38.448 133.068 ; 
      RECT 18.532 104.652 18.668 139.266 ; 
      RECT 18.324 104.652 18.46 139.266 ; 
      RECT 18.116 104.652 18.252 139.266 ; 
      RECT 17.908 104.652 18.044 139.266 ; 
      RECT 0 110.892 17.836 139.266 ; 
      RECT 0 119.532 19.708 131.34 ; 
      RECT 18.74 108.588 23.292 120.396 ; 
      RECT 23.364 110.508 38.448 139.266 ; 
      RECT 20.772 104.972 24.156 120.012 ; 
      RECT 16.02 106.86 19.116 118.668 ; 
      RECT 15.156 107.436 17.836 139.266 ; 
      RECT 0 109.74 15.084 139.266 ; 
      RECT 13.428 104.652 15.228 110.796 ; 
      RECT 28.548 104.652 29.34 139.266 ; 
      RECT 13.428 108.972 28.476 110.412 ; 
      RECT 9.972 107.436 13.356 139.266 ; 
      RECT 0 108.588 9.9 139.266 ; 
      RECT 27.684 104.652 38.448 109.644 ; 
      RECT 26.82 107.436 38.448 109.644 ; 
      RECT 0 108.588 26.748 109.644 ; 
      RECT 25.956 104.652 27.612 108.876 ; 
      RECT 20.612 107.436 38.448 108.876 ; 
      RECT 0.684 107.436 19.708 109.644 ; 
      RECT 18.74 107.244 19.708 139.266 ; 
      RECT 0 106.86 0.612 139.266 ; 
      RECT 19.188 104.652 20.7 107.724 ; 
      RECT 20.772 107.244 25.884 110.412 ; 
      RECT 12.564 107.244 15.948 109.644 ; 
      RECT 10.836 107.244 12.492 139.266 ; 
      RECT 0 106.86 10.764 107.724 ; 
      RECT 25.092 104.652 38.448 107.34 ; 
      RECT 19.188 104.972 25.02 107.34 ; 
      RECT 15.3 106.86 19.116 107.34 ; 
      RECT 11.7 104.652 15.228 107.34 ; 
      RECT 0 106.86 11.628 107.34 ; 
      RECT 23.364 104.652 38.448 107.148 ; 
      RECT 18.74 104.972 38.448 107.148 ; 
      RECT 0.54 104.652 17.836 107.148 ; 
      RECT 0 104.652 0.468 139.266 ; 
      RECT 0 104.652 23.292 105.996 ; 
      RECT 0 104.652 38.448 104.876 ; 
        RECT 0 141.068 38.448 141.588 ; 
        RECT 37.98 137.214 38.448 141.588 ; 
        RECT 23.364 140.684 37.908 141.588 ; 
        RECT 18.036 140.684 23.292 141.588 ; 
        RECT 15.156 137.214 17.676 141.588 ; 
        RECT 0.54 140.684 15.084 141.588 ; 
        RECT 0 137.214 0.468 141.588 ; 
        RECT 37.836 137.214 38.448 140.876 ; 
        RECT 23.58 137.214 37.764 141.588 ; 
        RECT 20.592 137.214 23.508 140.876 ; 
        RECT 19.944 137.996 20.448 141.588 ; 
        RECT 14.94 137.612 19.836 140.876 ; 
        RECT 0.684 137.214 14.868 141.588 ; 
        RECT 0 137.214 0.612 140.876 ; 
        RECT 20.376 137.214 38.448 140.492 ; 
        RECT 0 137.612 20.304 140.492 ; 
        RECT 19.476 137.214 38.448 137.9 ; 
        RECT 0 137.214 19.404 140.492 ; 
        RECT 0 137.214 38.448 137.516 ; 
        RECT 0 145.388 38.448 145.908 ; 
        RECT 37.98 141.534 38.448 145.908 ; 
        RECT 23.364 145.004 37.908 145.908 ; 
        RECT 18.036 145.004 23.292 145.908 ; 
        RECT 15.156 141.534 17.676 145.908 ; 
        RECT 0.54 145.004 15.084 145.908 ; 
        RECT 0 141.534 0.468 145.908 ; 
        RECT 37.836 141.534 38.448 145.196 ; 
        RECT 23.58 141.534 37.764 145.908 ; 
        RECT 20.592 141.534 23.508 145.196 ; 
        RECT 19.944 142.316 20.448 145.908 ; 
        RECT 14.94 141.932 19.836 145.196 ; 
        RECT 0.684 141.534 14.868 145.908 ; 
        RECT 0 141.534 0.612 145.196 ; 
        RECT 20.376 141.534 38.448 144.812 ; 
        RECT 0 141.932 20.304 144.812 ; 
        RECT 19.476 141.534 38.448 142.22 ; 
        RECT 0 141.534 19.404 144.812 ; 
        RECT 0 141.534 38.448 141.836 ; 
        RECT 0 149.708 38.448 150.228 ; 
        RECT 37.98 145.854 38.448 150.228 ; 
        RECT 23.364 149.324 37.908 150.228 ; 
        RECT 18.036 149.324 23.292 150.228 ; 
        RECT 15.156 145.854 17.676 150.228 ; 
        RECT 0.54 149.324 15.084 150.228 ; 
        RECT 0 145.854 0.468 150.228 ; 
        RECT 37.836 145.854 38.448 149.516 ; 
        RECT 23.58 145.854 37.764 150.228 ; 
        RECT 20.592 145.854 23.508 149.516 ; 
        RECT 19.944 146.636 20.448 150.228 ; 
        RECT 14.94 146.252 19.836 149.516 ; 
        RECT 0.684 145.854 14.868 150.228 ; 
        RECT 0 145.854 0.612 149.516 ; 
        RECT 20.376 145.854 38.448 149.132 ; 
        RECT 0 146.252 20.304 149.132 ; 
        RECT 19.476 145.854 38.448 146.54 ; 
        RECT 0 145.854 19.404 149.132 ; 
        RECT 0 145.854 38.448 146.156 ; 
        RECT 0 154.028 38.448 154.548 ; 
        RECT 37.98 150.174 38.448 154.548 ; 
        RECT 23.364 153.644 37.908 154.548 ; 
        RECT 18.036 153.644 23.292 154.548 ; 
        RECT 15.156 150.174 17.676 154.548 ; 
        RECT 0.54 153.644 15.084 154.548 ; 
        RECT 0 150.174 0.468 154.548 ; 
        RECT 37.836 150.174 38.448 153.836 ; 
        RECT 23.58 150.174 37.764 154.548 ; 
        RECT 20.592 150.174 23.508 153.836 ; 
        RECT 19.944 150.956 20.448 154.548 ; 
        RECT 14.94 150.572 19.836 153.836 ; 
        RECT 0.684 150.174 14.868 154.548 ; 
        RECT 0 150.174 0.612 153.836 ; 
        RECT 20.376 150.174 38.448 153.452 ; 
        RECT 0 150.572 20.304 153.452 ; 
        RECT 19.476 150.174 38.448 150.86 ; 
        RECT 0 150.174 19.404 153.452 ; 
        RECT 0 150.174 38.448 150.476 ; 
        RECT 0 158.348 38.448 158.868 ; 
        RECT 37.98 154.494 38.448 158.868 ; 
        RECT 23.364 157.964 37.908 158.868 ; 
        RECT 18.036 157.964 23.292 158.868 ; 
        RECT 15.156 154.494 17.676 158.868 ; 
        RECT 0.54 157.964 15.084 158.868 ; 
        RECT 0 154.494 0.468 158.868 ; 
        RECT 37.836 154.494 38.448 158.156 ; 
        RECT 23.58 154.494 37.764 158.868 ; 
        RECT 20.592 154.494 23.508 158.156 ; 
        RECT 19.944 155.276 20.448 158.868 ; 
        RECT 14.94 154.892 19.836 158.156 ; 
        RECT 0.684 154.494 14.868 158.868 ; 
        RECT 0 154.494 0.612 158.156 ; 
        RECT 20.376 154.494 38.448 157.772 ; 
        RECT 0 154.892 20.304 157.772 ; 
        RECT 19.476 154.494 38.448 155.18 ; 
        RECT 0 154.494 19.404 157.772 ; 
        RECT 0 154.494 38.448 154.796 ; 
        RECT 0 162.668 38.448 163.188 ; 
        RECT 37.98 158.814 38.448 163.188 ; 
        RECT 23.364 162.284 37.908 163.188 ; 
        RECT 18.036 162.284 23.292 163.188 ; 
        RECT 15.156 158.814 17.676 163.188 ; 
        RECT 0.54 162.284 15.084 163.188 ; 
        RECT 0 158.814 0.468 163.188 ; 
        RECT 37.836 158.814 38.448 162.476 ; 
        RECT 23.58 158.814 37.764 163.188 ; 
        RECT 20.592 158.814 23.508 162.476 ; 
        RECT 19.944 159.596 20.448 163.188 ; 
        RECT 14.94 159.212 19.836 162.476 ; 
        RECT 0.684 158.814 14.868 163.188 ; 
        RECT 0 158.814 0.612 162.476 ; 
        RECT 20.376 158.814 38.448 162.092 ; 
        RECT 0 159.212 20.304 162.092 ; 
        RECT 19.476 158.814 38.448 159.5 ; 
        RECT 0 158.814 19.404 162.092 ; 
        RECT 0 158.814 38.448 159.116 ; 
        RECT 0 166.988 38.448 167.508 ; 
        RECT 37.98 163.134 38.448 167.508 ; 
        RECT 23.364 166.604 37.908 167.508 ; 
        RECT 18.036 166.604 23.292 167.508 ; 
        RECT 15.156 163.134 17.676 167.508 ; 
        RECT 0.54 166.604 15.084 167.508 ; 
        RECT 0 163.134 0.468 167.508 ; 
        RECT 37.836 163.134 38.448 166.796 ; 
        RECT 23.58 163.134 37.764 167.508 ; 
        RECT 20.592 163.134 23.508 166.796 ; 
        RECT 19.944 163.916 20.448 167.508 ; 
        RECT 14.94 163.532 19.836 166.796 ; 
        RECT 0.684 163.134 14.868 167.508 ; 
        RECT 0 163.134 0.612 166.796 ; 
        RECT 20.376 163.134 38.448 166.412 ; 
        RECT 0 163.532 20.304 166.412 ; 
        RECT 19.476 163.134 38.448 163.82 ; 
        RECT 0 163.134 19.404 166.412 ; 
        RECT 0 163.134 38.448 163.436 ; 
        RECT 0 171.308 38.448 171.828 ; 
        RECT 37.98 167.454 38.448 171.828 ; 
        RECT 23.364 170.924 37.908 171.828 ; 
        RECT 18.036 170.924 23.292 171.828 ; 
        RECT 15.156 167.454 17.676 171.828 ; 
        RECT 0.54 170.924 15.084 171.828 ; 
        RECT 0 167.454 0.468 171.828 ; 
        RECT 37.836 167.454 38.448 171.116 ; 
        RECT 23.58 167.454 37.764 171.828 ; 
        RECT 20.592 167.454 23.508 171.116 ; 
        RECT 19.944 168.236 20.448 171.828 ; 
        RECT 14.94 167.852 19.836 171.116 ; 
        RECT 0.684 167.454 14.868 171.828 ; 
        RECT 0 167.454 0.612 171.116 ; 
        RECT 20.376 167.454 38.448 170.732 ; 
        RECT 0 167.852 20.304 170.732 ; 
        RECT 19.476 167.454 38.448 168.14 ; 
        RECT 0 167.454 19.404 170.732 ; 
        RECT 0 167.454 38.448 167.756 ; 
        RECT 0 175.628 38.448 176.148 ; 
        RECT 37.98 171.774 38.448 176.148 ; 
        RECT 23.364 175.244 37.908 176.148 ; 
        RECT 18.036 175.244 23.292 176.148 ; 
        RECT 15.156 171.774 17.676 176.148 ; 
        RECT 0.54 175.244 15.084 176.148 ; 
        RECT 0 171.774 0.468 176.148 ; 
        RECT 37.836 171.774 38.448 175.436 ; 
        RECT 23.58 171.774 37.764 176.148 ; 
        RECT 20.592 171.774 23.508 175.436 ; 
        RECT 19.944 172.556 20.448 176.148 ; 
        RECT 14.94 172.172 19.836 175.436 ; 
        RECT 0.684 171.774 14.868 176.148 ; 
        RECT 0 171.774 0.612 175.436 ; 
        RECT 20.376 171.774 38.448 175.052 ; 
        RECT 0 172.172 20.304 175.052 ; 
        RECT 19.476 171.774 38.448 172.46 ; 
        RECT 0 171.774 19.404 175.052 ; 
        RECT 0 171.774 38.448 172.076 ; 
        RECT 0 179.948 38.448 180.468 ; 
        RECT 37.98 176.094 38.448 180.468 ; 
        RECT 23.364 179.564 37.908 180.468 ; 
        RECT 18.036 179.564 23.292 180.468 ; 
        RECT 15.156 176.094 17.676 180.468 ; 
        RECT 0.54 179.564 15.084 180.468 ; 
        RECT 0 176.094 0.468 180.468 ; 
        RECT 37.836 176.094 38.448 179.756 ; 
        RECT 23.58 176.094 37.764 180.468 ; 
        RECT 20.592 176.094 23.508 179.756 ; 
        RECT 19.944 176.876 20.448 180.468 ; 
        RECT 14.94 176.492 19.836 179.756 ; 
        RECT 0.684 176.094 14.868 180.468 ; 
        RECT 0 176.094 0.612 179.756 ; 
        RECT 20.376 176.094 38.448 179.372 ; 
        RECT 0 176.492 20.304 179.372 ; 
        RECT 19.476 176.094 38.448 176.78 ; 
        RECT 0 176.094 19.404 179.372 ; 
        RECT 0 176.094 38.448 176.396 ; 
        RECT 0 184.268 38.448 184.788 ; 
        RECT 37.98 180.414 38.448 184.788 ; 
        RECT 23.364 183.884 37.908 184.788 ; 
        RECT 18.036 183.884 23.292 184.788 ; 
        RECT 15.156 180.414 17.676 184.788 ; 
        RECT 0.54 183.884 15.084 184.788 ; 
        RECT 0 180.414 0.468 184.788 ; 
        RECT 37.836 180.414 38.448 184.076 ; 
        RECT 23.58 180.414 37.764 184.788 ; 
        RECT 20.592 180.414 23.508 184.076 ; 
        RECT 19.944 181.196 20.448 184.788 ; 
        RECT 14.94 180.812 19.836 184.076 ; 
        RECT 0.684 180.414 14.868 184.788 ; 
        RECT 0 180.414 0.612 184.076 ; 
        RECT 20.376 180.414 38.448 183.692 ; 
        RECT 0 180.812 20.304 183.692 ; 
        RECT 19.476 180.414 38.448 181.1 ; 
        RECT 0 180.414 19.404 183.692 ; 
        RECT 0 180.414 38.448 180.716 ; 
        RECT 0 188.588 38.448 189.108 ; 
        RECT 37.98 184.734 38.448 189.108 ; 
        RECT 23.364 188.204 37.908 189.108 ; 
        RECT 18.036 188.204 23.292 189.108 ; 
        RECT 15.156 184.734 17.676 189.108 ; 
        RECT 0.54 188.204 15.084 189.108 ; 
        RECT 0 184.734 0.468 189.108 ; 
        RECT 37.836 184.734 38.448 188.396 ; 
        RECT 23.58 184.734 37.764 189.108 ; 
        RECT 20.592 184.734 23.508 188.396 ; 
        RECT 19.944 185.516 20.448 189.108 ; 
        RECT 14.94 185.132 19.836 188.396 ; 
        RECT 0.684 184.734 14.868 189.108 ; 
        RECT 0 184.734 0.612 188.396 ; 
        RECT 20.376 184.734 38.448 188.012 ; 
        RECT 0 185.132 20.304 188.012 ; 
        RECT 19.476 184.734 38.448 185.42 ; 
        RECT 0 184.734 19.404 188.012 ; 
        RECT 0 184.734 38.448 185.036 ; 
        RECT 0 192.908 38.448 193.428 ; 
        RECT 37.98 189.054 38.448 193.428 ; 
        RECT 23.364 192.524 37.908 193.428 ; 
        RECT 18.036 192.524 23.292 193.428 ; 
        RECT 15.156 189.054 17.676 193.428 ; 
        RECT 0.54 192.524 15.084 193.428 ; 
        RECT 0 189.054 0.468 193.428 ; 
        RECT 37.836 189.054 38.448 192.716 ; 
        RECT 23.58 189.054 37.764 193.428 ; 
        RECT 20.592 189.054 23.508 192.716 ; 
        RECT 19.944 189.836 20.448 193.428 ; 
        RECT 14.94 189.452 19.836 192.716 ; 
        RECT 0.684 189.054 14.868 193.428 ; 
        RECT 0 189.054 0.612 192.716 ; 
        RECT 20.376 189.054 38.448 192.332 ; 
        RECT 0 189.452 20.304 192.332 ; 
        RECT 19.476 189.054 38.448 189.74 ; 
        RECT 0 189.054 19.404 192.332 ; 
        RECT 0 189.054 38.448 189.356 ; 
        RECT 0 197.228 38.448 197.748 ; 
        RECT 37.98 193.374 38.448 197.748 ; 
        RECT 23.364 196.844 37.908 197.748 ; 
        RECT 18.036 196.844 23.292 197.748 ; 
        RECT 15.156 193.374 17.676 197.748 ; 
        RECT 0.54 196.844 15.084 197.748 ; 
        RECT 0 193.374 0.468 197.748 ; 
        RECT 37.836 193.374 38.448 197.036 ; 
        RECT 23.58 193.374 37.764 197.748 ; 
        RECT 20.592 193.374 23.508 197.036 ; 
        RECT 19.944 194.156 20.448 197.748 ; 
        RECT 14.94 193.772 19.836 197.036 ; 
        RECT 0.684 193.374 14.868 197.748 ; 
        RECT 0 193.374 0.612 197.036 ; 
        RECT 20.376 193.374 38.448 196.652 ; 
        RECT 0 193.772 20.304 196.652 ; 
        RECT 19.476 193.374 38.448 194.06 ; 
        RECT 0 193.374 19.404 196.652 ; 
        RECT 0 193.374 38.448 193.676 ; 
        RECT 0 201.548 38.448 202.068 ; 
        RECT 37.98 197.694 38.448 202.068 ; 
        RECT 23.364 201.164 37.908 202.068 ; 
        RECT 18.036 201.164 23.292 202.068 ; 
        RECT 15.156 197.694 17.676 202.068 ; 
        RECT 0.54 201.164 15.084 202.068 ; 
        RECT 0 197.694 0.468 202.068 ; 
        RECT 37.836 197.694 38.448 201.356 ; 
        RECT 23.58 197.694 37.764 202.068 ; 
        RECT 20.592 197.694 23.508 201.356 ; 
        RECT 19.944 198.476 20.448 202.068 ; 
        RECT 14.94 198.092 19.836 201.356 ; 
        RECT 0.684 197.694 14.868 202.068 ; 
        RECT 0 197.694 0.612 201.356 ; 
        RECT 20.376 197.694 38.448 200.972 ; 
        RECT 0 198.092 20.304 200.972 ; 
        RECT 19.476 197.694 38.448 198.38 ; 
        RECT 0 197.694 19.404 200.972 ; 
        RECT 0 197.694 38.448 197.996 ; 
        RECT 0 205.868 38.448 206.388 ; 
        RECT 37.98 202.014 38.448 206.388 ; 
        RECT 23.364 205.484 37.908 206.388 ; 
        RECT 18.036 205.484 23.292 206.388 ; 
        RECT 15.156 202.014 17.676 206.388 ; 
        RECT 0.54 205.484 15.084 206.388 ; 
        RECT 0 202.014 0.468 206.388 ; 
        RECT 37.836 202.014 38.448 205.676 ; 
        RECT 23.58 202.014 37.764 206.388 ; 
        RECT 20.592 202.014 23.508 205.676 ; 
        RECT 19.944 202.796 20.448 206.388 ; 
        RECT 14.94 202.412 19.836 205.676 ; 
        RECT 0.684 202.014 14.868 206.388 ; 
        RECT 0 202.014 0.612 205.676 ; 
        RECT 20.376 202.014 38.448 205.292 ; 
        RECT 0 202.412 20.304 205.292 ; 
        RECT 19.476 202.014 38.448 202.7 ; 
        RECT 0 202.014 19.404 205.292 ; 
        RECT 0 202.014 38.448 202.316 ; 
        RECT 0 210.188 38.448 210.708 ; 
        RECT 37.98 206.334 38.448 210.708 ; 
        RECT 23.364 209.804 37.908 210.708 ; 
        RECT 18.036 209.804 23.292 210.708 ; 
        RECT 15.156 206.334 17.676 210.708 ; 
        RECT 0.54 209.804 15.084 210.708 ; 
        RECT 0 206.334 0.468 210.708 ; 
        RECT 37.836 206.334 38.448 209.996 ; 
        RECT 23.58 206.334 37.764 210.708 ; 
        RECT 20.592 206.334 23.508 209.996 ; 
        RECT 19.944 207.116 20.448 210.708 ; 
        RECT 14.94 206.732 19.836 209.996 ; 
        RECT 0.684 206.334 14.868 210.708 ; 
        RECT 0 206.334 0.612 209.996 ; 
        RECT 20.376 206.334 38.448 209.612 ; 
        RECT 0 206.732 20.304 209.612 ; 
        RECT 19.476 206.334 38.448 207.02 ; 
        RECT 0 206.334 19.404 209.612 ; 
        RECT 0 206.334 38.448 206.636 ; 
        RECT 0 214.508 38.448 215.028 ; 
        RECT 37.98 210.654 38.448 215.028 ; 
        RECT 23.364 214.124 37.908 215.028 ; 
        RECT 18.036 214.124 23.292 215.028 ; 
        RECT 15.156 210.654 17.676 215.028 ; 
        RECT 0.54 214.124 15.084 215.028 ; 
        RECT 0 210.654 0.468 215.028 ; 
        RECT 37.836 210.654 38.448 214.316 ; 
        RECT 23.58 210.654 37.764 215.028 ; 
        RECT 20.592 210.654 23.508 214.316 ; 
        RECT 19.944 211.436 20.448 215.028 ; 
        RECT 14.94 211.052 19.836 214.316 ; 
        RECT 0.684 210.654 14.868 215.028 ; 
        RECT 0 210.654 0.612 214.316 ; 
        RECT 20.376 210.654 38.448 213.932 ; 
        RECT 0 211.052 20.304 213.932 ; 
        RECT 19.476 210.654 38.448 211.34 ; 
        RECT 0 210.654 19.404 213.932 ; 
        RECT 0 210.654 38.448 210.956 ; 
        RECT 0 218.828 38.448 219.348 ; 
        RECT 37.98 214.974 38.448 219.348 ; 
        RECT 23.364 218.444 37.908 219.348 ; 
        RECT 18.036 218.444 23.292 219.348 ; 
        RECT 15.156 214.974 17.676 219.348 ; 
        RECT 0.54 218.444 15.084 219.348 ; 
        RECT 0 214.974 0.468 219.348 ; 
        RECT 37.836 214.974 38.448 218.636 ; 
        RECT 23.58 214.974 37.764 219.348 ; 
        RECT 20.592 214.974 23.508 218.636 ; 
        RECT 19.944 215.756 20.448 219.348 ; 
        RECT 14.94 215.372 19.836 218.636 ; 
        RECT 0.684 214.974 14.868 219.348 ; 
        RECT 0 214.974 0.612 218.636 ; 
        RECT 20.376 214.974 38.448 218.252 ; 
        RECT 0 215.372 20.304 218.252 ; 
        RECT 19.476 214.974 38.448 215.66 ; 
        RECT 0 214.974 19.404 218.252 ; 
        RECT 0 214.974 38.448 215.276 ; 
        RECT 0 223.148 38.448 223.668 ; 
        RECT 37.98 219.294 38.448 223.668 ; 
        RECT 23.364 222.764 37.908 223.668 ; 
        RECT 18.036 222.764 23.292 223.668 ; 
        RECT 15.156 219.294 17.676 223.668 ; 
        RECT 0.54 222.764 15.084 223.668 ; 
        RECT 0 219.294 0.468 223.668 ; 
        RECT 37.836 219.294 38.448 222.956 ; 
        RECT 23.58 219.294 37.764 223.668 ; 
        RECT 20.592 219.294 23.508 222.956 ; 
        RECT 19.944 220.076 20.448 223.668 ; 
        RECT 14.94 219.692 19.836 222.956 ; 
        RECT 0.684 219.294 14.868 223.668 ; 
        RECT 0 219.294 0.612 222.956 ; 
        RECT 20.376 219.294 38.448 222.572 ; 
        RECT 0 219.692 20.304 222.572 ; 
        RECT 19.476 219.294 38.448 219.98 ; 
        RECT 0 219.294 19.404 222.572 ; 
        RECT 0 219.294 38.448 219.596 ; 
        RECT 0 227.468 38.448 227.988 ; 
        RECT 37.98 223.614 38.448 227.988 ; 
        RECT 23.364 227.084 37.908 227.988 ; 
        RECT 18.036 227.084 23.292 227.988 ; 
        RECT 15.156 223.614 17.676 227.988 ; 
        RECT 0.54 227.084 15.084 227.988 ; 
        RECT 0 223.614 0.468 227.988 ; 
        RECT 37.836 223.614 38.448 227.276 ; 
        RECT 23.58 223.614 37.764 227.988 ; 
        RECT 20.592 223.614 23.508 227.276 ; 
        RECT 19.944 224.396 20.448 227.988 ; 
        RECT 14.94 224.012 19.836 227.276 ; 
        RECT 0.684 223.614 14.868 227.988 ; 
        RECT 0 223.614 0.612 227.276 ; 
        RECT 20.376 223.614 38.448 226.892 ; 
        RECT 0 224.012 20.304 226.892 ; 
        RECT 19.476 223.614 38.448 224.3 ; 
        RECT 0 223.614 19.404 226.892 ; 
        RECT 0 223.614 38.448 223.916 ; 
        RECT 0 231.788 38.448 232.308 ; 
        RECT 37.98 227.934 38.448 232.308 ; 
        RECT 23.364 231.404 37.908 232.308 ; 
        RECT 18.036 231.404 23.292 232.308 ; 
        RECT 15.156 227.934 17.676 232.308 ; 
        RECT 0.54 231.404 15.084 232.308 ; 
        RECT 0 227.934 0.468 232.308 ; 
        RECT 37.836 227.934 38.448 231.596 ; 
        RECT 23.58 227.934 37.764 232.308 ; 
        RECT 20.592 227.934 23.508 231.596 ; 
        RECT 19.944 228.716 20.448 232.308 ; 
        RECT 14.94 228.332 19.836 231.596 ; 
        RECT 0.684 227.934 14.868 232.308 ; 
        RECT 0 227.934 0.612 231.596 ; 
        RECT 20.376 227.934 38.448 231.212 ; 
        RECT 0 228.332 20.304 231.212 ; 
        RECT 19.476 227.934 38.448 228.62 ; 
        RECT 0 227.934 19.404 231.212 ; 
        RECT 0 227.934 38.448 228.236 ; 
        RECT 0 236.108 38.448 236.628 ; 
        RECT 37.98 232.254 38.448 236.628 ; 
        RECT 23.364 235.724 37.908 236.628 ; 
        RECT 18.036 235.724 23.292 236.628 ; 
        RECT 15.156 232.254 17.676 236.628 ; 
        RECT 0.54 235.724 15.084 236.628 ; 
        RECT 0 232.254 0.468 236.628 ; 
        RECT 37.836 232.254 38.448 235.916 ; 
        RECT 23.58 232.254 37.764 236.628 ; 
        RECT 20.592 232.254 23.508 235.916 ; 
        RECT 19.944 233.036 20.448 236.628 ; 
        RECT 14.94 232.652 19.836 235.916 ; 
        RECT 0.684 232.254 14.868 236.628 ; 
        RECT 0 232.254 0.612 235.916 ; 
        RECT 20.376 232.254 38.448 235.532 ; 
        RECT 0 232.652 20.304 235.532 ; 
        RECT 19.476 232.254 38.448 232.94 ; 
        RECT 0 232.254 19.404 235.532 ; 
        RECT 0 232.254 38.448 232.556 ; 
        RECT 0 240.428 38.448 240.948 ; 
        RECT 37.98 236.574 38.448 240.948 ; 
        RECT 23.364 240.044 37.908 240.948 ; 
        RECT 18.036 240.044 23.292 240.948 ; 
        RECT 15.156 236.574 17.676 240.948 ; 
        RECT 0.54 240.044 15.084 240.948 ; 
        RECT 0 236.574 0.468 240.948 ; 
        RECT 37.836 236.574 38.448 240.236 ; 
        RECT 23.58 236.574 37.764 240.948 ; 
        RECT 20.592 236.574 23.508 240.236 ; 
        RECT 19.944 237.356 20.448 240.948 ; 
        RECT 14.94 236.972 19.836 240.236 ; 
        RECT 0.684 236.574 14.868 240.948 ; 
        RECT 0 236.574 0.612 240.236 ; 
        RECT 20.376 236.574 38.448 239.852 ; 
        RECT 0 236.972 20.304 239.852 ; 
        RECT 19.476 236.574 38.448 237.26 ; 
        RECT 0 236.574 19.404 239.852 ; 
        RECT 0 236.574 38.448 236.876 ; 
  LAYER M4 ; 
      RECT 6.428 111.504 32.01 111.6 ; 
      RECT 6.428 112.656 32.01 112.752 ; 
      RECT 6.428 114.192 32.01 114.288 ; 
      RECT 6.428 114.576 32.01 114.672 ; 
      RECT 6.428 115.92 32.01 116.016 ; 
      RECT 29.996 107.34 30.332 107.436 ; 
      RECT 29.276 109.068 29.744 109.164 ; 
      RECT 29.276 111.696 29.744 111.792 ; 
      RECT 29.276 112.848 29.744 112.944 ; 
      RECT 26.714 109.068 28.992 109.164 ; 
      RECT 26.972 112.176 27.404 112.272 ; 
      RECT 21.628 113.676 26 113.772 ; 
      RECT 24.38 111.948 24.716 112.044 ; 
      RECT 21.244 116.748 24.716 116.844 ; 
      RECT 24.38 117.132 24.716 117.228 ; 
      RECT 23.668 110.028 24.004 110.124 ; 
      RECT 23.516 115.404 23.852 115.5 ; 
      RECT 22.804 109.644 23.14 109.74 ; 
      RECT 21.948 104.492 23 104.588 ; 
      RECT 21.948 139.052 23 139.148 ; 
      RECT 22.012 115.596 22.988 115.692 ; 
      RECT 22.652 116.172 22.988 116.268 ; 
      RECT 16.828 117.132 22.988 117.228 ; 
      RECT 22.652 118.284 22.988 118.38 ; 
      RECT 21.716 138.668 22.768 138.764 ; 
      RECT 21.712 104.108 22.764 104.204 ; 
      RECT 21.56 103.724 22.612 103.82 ; 
      RECT 21.56 137.9 22.612 137.996 ; 
      RECT 22.22 120.012 22.556 120.108 ; 
      RECT 19.132 121.548 22.556 121.644 ; 
      RECT 20.668 130.572 22.556 130.668 ; 
      RECT 22.22 130.956 22.556 131.052 ; 
      RECT 21.368 103.34 22.42 103.436 ; 
      RECT 21.368 137.516 22.42 137.612 ; 
      RECT 20.476 126.924 22.256 127.02 ; 
      RECT 21.192 102.956 22.244 103.052 ; 
      RECT 21.192 138.86 22.244 138.956 ; 
      RECT 20.996 104.3 22.048 104.396 ; 
      RECT 20.996 138.476 22.048 138.572 ; 
      RECT 21.52 116.172 22.004 116.268 ; 
      RECT 21.436 124.62 21.968 124.716 ; 
      RECT 20.808 103.916 21.86 104.012 ; 
      RECT 20.808 138.092 21.86 138.188 ; 
      RECT 20.668 102.764 21.72 102.86 ; 
      RECT 20.668 137.708 21.72 137.804 ; 
      RECT 17.404 130.956 21.68 131.052 ; 
      RECT 21.344 135.564 21.68 135.66 ; 
      RECT 20.444 102.188 21.496 102.284 ; 
      RECT 20.444 137.324 21.496 137.42 ; 
      RECT 21.052 120.012 21.392 120.108 ; 
      RECT 16.636 122.316 21.104 122.412 ; 
      RECT 19.216 113.676 21.044 113.772 ; 
      RECT 18.524 105.068 19.592 105.164 ; 
      RECT 18.524 136.748 19.592 136.844 ; 
      RECT 19.072 119.82 19.508 119.916 ; 
      RECT 18.432 104.684 19.4 104.78 ; 
      RECT 18.432 139.244 19.4 139.34 ; 
      RECT 18.208 102.764 19.176 102.86 ; 
      RECT 18.324 139.628 19.176 139.724 ; 
      RECT 18.788 118.284 19.124 118.38 ; 
      RECT 17.992 103.148 18.984 103.244 ; 
      RECT 17.992 139.052 18.984 139.148 ; 
      RECT 17.056 128.652 18.74 128.748 ; 
      RECT 16.928 104.492 17.996 104.588 ; 
      RECT 16.928 139.628 17.996 139.724 ; 
      RECT 17.488 122.892 17.972 122.988 ; 
      RECT 17.456 135.564 17.792 135.66 ; 
      RECT 16.792 104.108 17.78 104.204 ; 
      RECT 16.524 137.9 17.78 137.996 ; 
      RECT 16.688 103.724 17.608 103.82 ; 
      RECT 16.64 139.244 17.608 139.34 ; 
      RECT 16.476 103.34 17.396 103.436 ; 
      RECT 17.06 129.228 17.396 129.324 ; 
      RECT 16.276 137.516 17.396 137.612 ; 
      RECT 16.296 102.956 17.216 103.052 ; 
      RECT 16.296 138.86 17.216 138.956 ; 
      RECT 12.448 118.284 17.204 118.38 ; 
      RECT 16.144 103.916 17.064 104.012 ; 
      RECT 16.144 138.476 17.064 138.572 ; 
      RECT 16.072 103.532 16.844 103.628 ; 
      RECT 16.072 138.092 16.844 138.188 ; 
      RECT 15.876 103.148 16.648 103.244 ; 
      RECT 15.876 137.708 16.648 137.804 ; 
      RECT 15.892 121.932 16.628 122.028 ; 
      RECT 15.668 102.764 16.44 102.86 ; 
      RECT 15.668 137.324 16.44 137.42 ; 
      RECT 13.732 111.18 16.436 111.276 ; 
      RECT 15.892 122.316 16.228 122.412 ; 
      RECT 14.816 104.876 15.868 104.972 ; 
      RECT 15.032 120.012 15.48 120.108 ; 
      RECT 13.58 111.948 13.916 112.044 ; 
  LAYER V4 ; 
      RECT 30.192 107.34 30.288 107.436 ; 
      RECT 30.192 111.504 30.288 111.6 ; 
      RECT 29.52 109.068 29.616 109.164 ; 
      RECT 29.52 111.696 29.616 111.792 ; 
      RECT 29.52 112.848 29.616 112.944 ; 
      RECT 27.024 109.068 27.12 109.164 ; 
      RECT 27.024 112.176 27.12 112.272 ; 
      RECT 24.576 111.948 24.672 112.044 ; 
      RECT 24.576 112.656 24.672 112.752 ; 
      RECT 24.576 116.748 24.672 116.844 ; 
      RECT 24.576 117.132 24.672 117.228 ; 
      RECT 23.712 110.028 23.808 110.124 ; 
      RECT 23.712 114.192 23.808 114.288 ; 
      RECT 23.712 115.404 23.808 115.5 ; 
      RECT 23.712 115.92 23.808 116.016 ; 
      RECT 22.848 109.644 22.944 109.74 ; 
      RECT 22.848 114.576 22.944 114.672 ; 
      RECT 22.848 115.596 22.944 115.692 ; 
      RECT 22.848 116.172 22.944 116.268 ; 
      RECT 22.848 117.132 22.944 117.228 ; 
      RECT 22.848 118.284 22.944 118.38 ; 
      RECT 22.416 120.012 22.512 120.108 ; 
      RECT 22.416 121.548 22.512 121.644 ; 
      RECT 22.416 130.572 22.512 130.668 ; 
      RECT 22.416 130.956 22.512 131.052 ; 
      RECT 22.056 104.492 22.152 104.588 ; 
      RECT 22.056 115.596 22.152 115.692 ; 
      RECT 22.056 139.052 22.152 139.148 ; 
      RECT 21.864 104.108 21.96 104.204 ; 
      RECT 21.864 116.172 21.96 116.268 ; 
      RECT 21.864 138.668 21.96 138.764 ; 
      RECT 21.672 103.724 21.768 103.82 ; 
      RECT 21.672 113.676 21.768 113.772 ; 
      RECT 21.672 137.9 21.768 137.996 ; 
      RECT 21.48 103.34 21.576 103.436 ; 
      RECT 21.48 124.62 21.576 124.716 ; 
      RECT 21.48 135.564 21.576 135.66 ; 
      RECT 21.48 137.516 21.576 137.612 ; 
      RECT 21.288 102.956 21.384 103.052 ; 
      RECT 21.288 116.748 21.384 116.844 ; 
      RECT 21.288 138.86 21.384 138.956 ; 
      RECT 21.096 104.3 21.192 104.396 ; 
      RECT 21.096 120.012 21.192 120.108 ; 
      RECT 21.096 138.476 21.192 138.572 ; 
      RECT 20.904 103.916 21 104.012 ; 
      RECT 20.904 113.676 21 113.772 ; 
      RECT 20.904 138.092 21 138.188 ; 
      RECT 20.712 102.764 20.808 102.86 ; 
      RECT 20.712 130.572 20.808 130.668 ; 
      RECT 20.712 137.708 20.808 137.804 ; 
      RECT 20.52 102.188 20.616 102.284 ; 
      RECT 20.52 126.924 20.616 127.02 ; 
      RECT 20.52 137.324 20.616 137.42 ; 
      RECT 19.368 105.068 19.464 105.164 ; 
      RECT 19.368 119.82 19.464 119.916 ; 
      RECT 19.368 136.748 19.464 136.844 ; 
      RECT 19.176 104.684 19.272 104.78 ; 
      RECT 19.176 121.548 19.272 121.644 ; 
      RECT 19.176 139.244 19.272 139.34 ; 
      RECT 18.984 102.764 19.08 102.86 ; 
      RECT 18.984 118.284 19.08 118.38 ; 
      RECT 18.984 139.628 19.08 139.724 ; 
      RECT 18.6 103.148 18.696 103.244 ; 
      RECT 18.6 128.652 18.696 128.748 ; 
      RECT 18.6 139.052 18.696 139.148 ; 
      RECT 17.832 104.492 17.928 104.588 ; 
      RECT 17.832 122.892 17.928 122.988 ; 
      RECT 17.832 139.628 17.928 139.724 ; 
      RECT 17.64 104.108 17.736 104.204 ; 
      RECT 17.64 135.564 17.736 135.66 ; 
      RECT 17.64 137.9 17.736 137.996 ; 
      RECT 17.448 103.724 17.544 103.82 ; 
      RECT 17.448 130.956 17.544 131.052 ; 
      RECT 17.448 139.244 17.544 139.34 ; 
      RECT 17.256 103.34 17.352 103.436 ; 
      RECT 17.256 129.228 17.352 129.324 ; 
      RECT 17.256 137.516 17.352 137.612 ; 
      RECT 17.064 102.956 17.16 103.052 ; 
      RECT 17.064 118.284 17.16 118.38 ; 
      RECT 17.064 138.86 17.16 138.956 ; 
      RECT 16.872 103.916 16.968 104.012 ; 
      RECT 16.872 117.132 16.968 117.228 ; 
      RECT 16.872 138.476 16.968 138.572 ; 
      RECT 16.68 103.532 16.776 103.628 ; 
      RECT 16.68 122.316 16.776 122.412 ; 
      RECT 16.68 138.092 16.776 138.188 ; 
      RECT 16.488 103.148 16.584 103.244 ; 
      RECT 16.488 121.932 16.584 122.028 ; 
      RECT 16.488 137.708 16.584 137.804 ; 
      RECT 16.296 102.764 16.392 102.86 ; 
      RECT 16.296 111.18 16.392 111.276 ; 
      RECT 16.296 137.324 16.392 137.42 ; 
      RECT 15.936 121.932 16.032 122.028 ; 
      RECT 15.936 122.316 16.032 122.412 ; 
      RECT 15.268 104.876 15.364 104.972 ; 
      RECT 15.268 120.012 15.364 120.108 ; 
      RECT 13.776 111.18 13.872 111.276 ; 
      RECT 13.776 111.948 13.872 112.044 ; 
  LAYER M5 ; 
      RECT 30.192 107.296 30.288 111.644 ; 
      RECT 29.52 109.014 29.616 113.144 ; 
      RECT 27.024 108.99 27.12 112.32 ; 
      RECT 24.576 111.904 24.672 112.796 ; 
      RECT 24.576 116.704 24.672 117.272 ; 
      RECT 23.712 109.984 23.808 114.332 ; 
      RECT 23.712 115.36 23.808 116.06 ; 
      RECT 22.848 109.6 22.944 114.716 ; 
      RECT 22.848 115.552 22.944 116.312 ; 
      RECT 22.848 117.088 22.944 118.424 ; 
      RECT 22.416 119.968 22.512 121.688 ; 
      RECT 22.416 130.528 22.512 131.096 ; 
      RECT 22.056 105.84 22.152 136.172 ; 
      RECT 21.864 105.84 21.96 136.172 ; 
      RECT 21.672 105.84 21.768 136.172 ; 
      RECT 21.48 105.84 21.576 136.172 ; 
      RECT 21.288 105.84 21.384 136.172 ; 
      RECT 21.096 105.84 21.192 136.172 ; 
      RECT 20.904 105.84 21 136.172 ; 
      RECT 20.712 105.84 20.808 136.172 ; 
      RECT 20.52 105.84 20.616 136.172 ; 
      RECT 19.368 104.792 19.464 136.924 ; 
      RECT 19.176 102.708 19.272 140.024 ; 
      RECT 18.984 102.584 19.08 140.02 ; 
      RECT 18.6 102.768 18.696 140.024 ; 
      RECT 17.832 102.764 17.928 139.836 ; 
      RECT 17.64 102.764 17.736 139.836 ; 
      RECT 17.448 102.764 17.544 139.836 ; 
      RECT 17.256 102.764 17.352 139.836 ; 
      RECT 17.064 102.764 17.16 139.836 ; 
      RECT 16.872 102.648 16.968 139.836 ; 
      RECT 16.68 102.472 16.776 139.84 ; 
      RECT 16.488 102.324 16.584 139.844 ; 
      RECT 16.296 102.084 16.392 139.844 ; 
      RECT 15.936 121.888 16.032 122.456 ; 
      RECT 15.268 104.804 15.364 120.18 ; 
      RECT 13.776 111.136 13.872 112.088 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 38.016 241.776 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 38.016 241.776 ; 
  END 
END srambank_64x4x48_6t122 
