VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_128x4x34_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_128x4x34_6t122 0 0 ; 
  SIZE 64 BY 181.44 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.688 65.768 4.88 ; 
        RECT 0.376 9.008 65.768 9.2 ; 
        RECT 0.376 13.328 65.768 13.52 ; 
        RECT 0.376 17.648 65.768 17.84 ; 
        RECT 0.376 21.968 65.768 22.16 ; 
        RECT 0.376 26.288 65.768 26.48 ; 
        RECT 0.376 30.608 65.768 30.8 ; 
        RECT 0.376 34.928 65.768 35.12 ; 
        RECT 0.376 39.248 65.768 39.44 ; 
        RECT 0.376 43.568 65.768 43.76 ; 
        RECT 0.376 47.888 65.768 48.08 ; 
        RECT 0.376 52.208 65.768 52.4 ; 
        RECT 0.376 56.528 65.768 56.72 ; 
        RECT 0.376 60.848 65.768 61.04 ; 
        RECT 0.376 65.168 65.768 65.36 ; 
        RECT 0.376 69.488 65.768 69.68 ; 
        RECT 0.376 73.808 65.768 74 ; 
        RECT 14.256 75.732 51.84 76.596 ; 
        RECT 36.788 89.748 37.352 89.844 ; 
        RECT 36.264 74.612 37.316 74.708 ; 
        RECT 29.592 88.404 36.504 89.268 ; 
        RECT 29.592 101.076 36.504 101.94 ; 
        RECT 0.376 110.636 65.768 110.828 ; 
        RECT 0.376 114.956 65.768 115.148 ; 
        RECT 0.376 119.276 65.768 119.468 ; 
        RECT 0.376 123.596 65.768 123.788 ; 
        RECT 0.376 127.916 65.768 128.108 ; 
        RECT 0.376 132.236 65.768 132.428 ; 
        RECT 0.376 136.556 65.768 136.748 ; 
        RECT 0.376 140.876 65.768 141.068 ; 
        RECT 0.376 145.196 65.768 145.388 ; 
        RECT 0.376 149.516 65.768 149.708 ; 
        RECT 0.376 153.836 65.768 154.028 ; 
        RECT 0.376 158.156 65.768 158.348 ; 
        RECT 0.376 162.476 65.768 162.668 ; 
        RECT 0.376 166.796 65.768 166.988 ; 
        RECT 0.376 171.116 65.768 171.308 ; 
        RECT 0.376 175.436 65.768 175.628 ; 
        RECT 0.376 179.756 65.768 179.948 ; 
      LAYER M3 ; 
        RECT 65.576 0.866 65.648 5.506 ; 
        RECT 37.136 0.868 37.208 5.504 ; 
        RECT 31.52 1.028 31.88 5.484 ; 
        RECT 28.928 0.868 29 5.504 ; 
        RECT 0.488 0.866 0.56 5.506 ; 
        RECT 65.576 5.186 65.648 9.826 ; 
        RECT 37.136 5.188 37.208 9.824 ; 
        RECT 31.52 5.348 31.88 9.804 ; 
        RECT 28.928 5.188 29 9.824 ; 
        RECT 0.488 5.186 0.56 9.826 ; 
        RECT 65.576 9.506 65.648 14.146 ; 
        RECT 37.136 9.508 37.208 14.144 ; 
        RECT 31.52 9.668 31.88 14.124 ; 
        RECT 28.928 9.508 29 14.144 ; 
        RECT 0.488 9.506 0.56 14.146 ; 
        RECT 65.576 13.826 65.648 18.466 ; 
        RECT 37.136 13.828 37.208 18.464 ; 
        RECT 31.52 13.988 31.88 18.444 ; 
        RECT 28.928 13.828 29 18.464 ; 
        RECT 0.488 13.826 0.56 18.466 ; 
        RECT 65.576 18.146 65.648 22.786 ; 
        RECT 37.136 18.148 37.208 22.784 ; 
        RECT 31.52 18.308 31.88 22.764 ; 
        RECT 28.928 18.148 29 22.784 ; 
        RECT 0.488 18.146 0.56 22.786 ; 
        RECT 65.576 22.466 65.648 27.106 ; 
        RECT 37.136 22.468 37.208 27.104 ; 
        RECT 31.52 22.628 31.88 27.084 ; 
        RECT 28.928 22.468 29 27.104 ; 
        RECT 0.488 22.466 0.56 27.106 ; 
        RECT 65.576 26.786 65.648 31.426 ; 
        RECT 37.136 26.788 37.208 31.424 ; 
        RECT 31.52 26.948 31.88 31.404 ; 
        RECT 28.928 26.788 29 31.424 ; 
        RECT 0.488 26.786 0.56 31.426 ; 
        RECT 65.576 31.106 65.648 35.746 ; 
        RECT 37.136 31.108 37.208 35.744 ; 
        RECT 31.52 31.268 31.88 35.724 ; 
        RECT 28.928 31.108 29 35.744 ; 
        RECT 0.488 31.106 0.56 35.746 ; 
        RECT 65.576 35.426 65.648 40.066 ; 
        RECT 37.136 35.428 37.208 40.064 ; 
        RECT 31.52 35.588 31.88 40.044 ; 
        RECT 28.928 35.428 29 40.064 ; 
        RECT 0.488 35.426 0.56 40.066 ; 
        RECT 65.576 39.746 65.648 44.386 ; 
        RECT 37.136 39.748 37.208 44.384 ; 
        RECT 31.52 39.908 31.88 44.364 ; 
        RECT 28.928 39.748 29 44.384 ; 
        RECT 0.488 39.746 0.56 44.386 ; 
        RECT 65.576 44.066 65.648 48.706 ; 
        RECT 37.136 44.068 37.208 48.704 ; 
        RECT 31.52 44.228 31.88 48.684 ; 
        RECT 28.928 44.068 29 48.704 ; 
        RECT 0.488 44.066 0.56 48.706 ; 
        RECT 65.576 48.386 65.648 53.026 ; 
        RECT 37.136 48.388 37.208 53.024 ; 
        RECT 31.52 48.548 31.88 53.004 ; 
        RECT 28.928 48.388 29 53.024 ; 
        RECT 0.488 48.386 0.56 53.026 ; 
        RECT 65.576 52.706 65.648 57.346 ; 
        RECT 37.136 52.708 37.208 57.344 ; 
        RECT 31.52 52.868 31.88 57.324 ; 
        RECT 28.928 52.708 29 57.344 ; 
        RECT 0.488 52.706 0.56 57.346 ; 
        RECT 65.576 57.026 65.648 61.666 ; 
        RECT 37.136 57.028 37.208 61.664 ; 
        RECT 31.52 57.188 31.88 61.644 ; 
        RECT 28.928 57.028 29 61.664 ; 
        RECT 0.488 57.026 0.56 61.666 ; 
        RECT 65.576 61.346 65.648 65.986 ; 
        RECT 37.136 61.348 37.208 65.984 ; 
        RECT 31.52 61.508 31.88 65.964 ; 
        RECT 28.928 61.348 29 65.984 ; 
        RECT 0.488 61.346 0.56 65.986 ; 
        RECT 65.576 65.666 65.648 70.306 ; 
        RECT 37.136 65.668 37.208 70.304 ; 
        RECT 31.52 65.828 31.88 70.284 ; 
        RECT 28.928 65.668 29 70.304 ; 
        RECT 0.488 65.666 0.56 70.306 ; 
        RECT 65.576 69.986 65.648 74.626 ; 
        RECT 37.136 69.988 37.208 74.624 ; 
        RECT 31.52 70.148 31.88 74.604 ; 
        RECT 28.928 69.988 29 74.624 ; 
        RECT 0.488 69.986 0.56 74.626 ; 
        RECT 65.556 74.282 65.628 107.11 ; 
        RECT 37.188 89.56 37.26 106.954 ; 
        RECT 37.116 74.414 37.188 74.966 ; 
        RECT 31.644 75.576 32.58 105.908 ; 
        RECT 31.5 105.576 31.86 107.08 ; 
        RECT 31.5 74.44 31.86 75.944 ; 
        RECT 0.468 74.282 0.54 107.11 ; 
        RECT 65.576 106.814 65.648 111.454 ; 
        RECT 37.136 106.816 37.208 111.452 ; 
        RECT 31.52 106.976 31.88 111.432 ; 
        RECT 28.928 106.816 29 111.452 ; 
        RECT 0.488 106.814 0.56 111.454 ; 
        RECT 65.576 111.134 65.648 115.774 ; 
        RECT 37.136 111.136 37.208 115.772 ; 
        RECT 31.52 111.296 31.88 115.752 ; 
        RECT 28.928 111.136 29 115.772 ; 
        RECT 0.488 111.134 0.56 115.774 ; 
        RECT 65.576 115.454 65.648 120.094 ; 
        RECT 37.136 115.456 37.208 120.092 ; 
        RECT 31.52 115.616 31.88 120.072 ; 
        RECT 28.928 115.456 29 120.092 ; 
        RECT 0.488 115.454 0.56 120.094 ; 
        RECT 65.576 119.774 65.648 124.414 ; 
        RECT 37.136 119.776 37.208 124.412 ; 
        RECT 31.52 119.936 31.88 124.392 ; 
        RECT 28.928 119.776 29 124.412 ; 
        RECT 0.488 119.774 0.56 124.414 ; 
        RECT 65.576 124.094 65.648 128.734 ; 
        RECT 37.136 124.096 37.208 128.732 ; 
        RECT 31.52 124.256 31.88 128.712 ; 
        RECT 28.928 124.096 29 128.732 ; 
        RECT 0.488 124.094 0.56 128.734 ; 
        RECT 65.576 128.414 65.648 133.054 ; 
        RECT 37.136 128.416 37.208 133.052 ; 
        RECT 31.52 128.576 31.88 133.032 ; 
        RECT 28.928 128.416 29 133.052 ; 
        RECT 0.488 128.414 0.56 133.054 ; 
        RECT 65.576 132.734 65.648 137.374 ; 
        RECT 37.136 132.736 37.208 137.372 ; 
        RECT 31.52 132.896 31.88 137.352 ; 
        RECT 28.928 132.736 29 137.372 ; 
        RECT 0.488 132.734 0.56 137.374 ; 
        RECT 65.576 137.054 65.648 141.694 ; 
        RECT 37.136 137.056 37.208 141.692 ; 
        RECT 31.52 137.216 31.88 141.672 ; 
        RECT 28.928 137.056 29 141.692 ; 
        RECT 0.488 137.054 0.56 141.694 ; 
        RECT 65.576 141.374 65.648 146.014 ; 
        RECT 37.136 141.376 37.208 146.012 ; 
        RECT 31.52 141.536 31.88 145.992 ; 
        RECT 28.928 141.376 29 146.012 ; 
        RECT 0.488 141.374 0.56 146.014 ; 
        RECT 65.576 145.694 65.648 150.334 ; 
        RECT 37.136 145.696 37.208 150.332 ; 
        RECT 31.52 145.856 31.88 150.312 ; 
        RECT 28.928 145.696 29 150.332 ; 
        RECT 0.488 145.694 0.56 150.334 ; 
        RECT 65.576 150.014 65.648 154.654 ; 
        RECT 37.136 150.016 37.208 154.652 ; 
        RECT 31.52 150.176 31.88 154.632 ; 
        RECT 28.928 150.016 29 154.652 ; 
        RECT 0.488 150.014 0.56 154.654 ; 
        RECT 65.576 154.334 65.648 158.974 ; 
        RECT 37.136 154.336 37.208 158.972 ; 
        RECT 31.52 154.496 31.88 158.952 ; 
        RECT 28.928 154.336 29 158.972 ; 
        RECT 0.488 154.334 0.56 158.974 ; 
        RECT 65.576 158.654 65.648 163.294 ; 
        RECT 37.136 158.656 37.208 163.292 ; 
        RECT 31.52 158.816 31.88 163.272 ; 
        RECT 28.928 158.656 29 163.292 ; 
        RECT 0.488 158.654 0.56 163.294 ; 
        RECT 65.576 162.974 65.648 167.614 ; 
        RECT 37.136 162.976 37.208 167.612 ; 
        RECT 31.52 163.136 31.88 167.592 ; 
        RECT 28.928 162.976 29 167.612 ; 
        RECT 0.488 162.974 0.56 167.614 ; 
        RECT 65.576 167.294 65.648 171.934 ; 
        RECT 37.136 167.296 37.208 171.932 ; 
        RECT 31.52 167.456 31.88 171.912 ; 
        RECT 28.928 167.296 29 171.932 ; 
        RECT 0.488 167.294 0.56 171.934 ; 
        RECT 65.576 171.614 65.648 176.254 ; 
        RECT 37.136 171.616 37.208 176.252 ; 
        RECT 31.52 171.776 31.88 176.232 ; 
        RECT 28.928 171.616 29 176.252 ; 
        RECT 0.488 171.614 0.56 176.254 ; 
        RECT 65.576 175.934 65.648 180.574 ; 
        RECT 37.136 175.936 37.208 180.572 ; 
        RECT 31.52 176.096 31.88 180.552 ; 
        RECT 28.928 175.936 29 180.572 ; 
        RECT 0.488 175.934 0.56 180.574 ; 
      LAYER V3 ; 
        RECT 0.488 4.688 0.56 4.88 ; 
        RECT 28.928 4.688 29 4.88 ; 
        RECT 31.52 4.688 31.88 4.88 ; 
        RECT 37.136 4.688 37.208 4.88 ; 
        RECT 65.576 4.688 65.648 4.88 ; 
        RECT 0.488 9.008 0.56 9.2 ; 
        RECT 28.928 9.008 29 9.2 ; 
        RECT 31.52 9.008 31.88 9.2 ; 
        RECT 37.136 9.008 37.208 9.2 ; 
        RECT 65.576 9.008 65.648 9.2 ; 
        RECT 0.488 13.328 0.56 13.52 ; 
        RECT 28.928 13.328 29 13.52 ; 
        RECT 31.52 13.328 31.88 13.52 ; 
        RECT 37.136 13.328 37.208 13.52 ; 
        RECT 65.576 13.328 65.648 13.52 ; 
        RECT 0.488 17.648 0.56 17.84 ; 
        RECT 28.928 17.648 29 17.84 ; 
        RECT 31.52 17.648 31.88 17.84 ; 
        RECT 37.136 17.648 37.208 17.84 ; 
        RECT 65.576 17.648 65.648 17.84 ; 
        RECT 0.488 21.968 0.56 22.16 ; 
        RECT 28.928 21.968 29 22.16 ; 
        RECT 31.52 21.968 31.88 22.16 ; 
        RECT 37.136 21.968 37.208 22.16 ; 
        RECT 65.576 21.968 65.648 22.16 ; 
        RECT 0.488 26.288 0.56 26.48 ; 
        RECT 28.928 26.288 29 26.48 ; 
        RECT 31.52 26.288 31.88 26.48 ; 
        RECT 37.136 26.288 37.208 26.48 ; 
        RECT 65.576 26.288 65.648 26.48 ; 
        RECT 0.488 30.608 0.56 30.8 ; 
        RECT 28.928 30.608 29 30.8 ; 
        RECT 31.52 30.608 31.88 30.8 ; 
        RECT 37.136 30.608 37.208 30.8 ; 
        RECT 65.576 30.608 65.648 30.8 ; 
        RECT 0.488 34.928 0.56 35.12 ; 
        RECT 28.928 34.928 29 35.12 ; 
        RECT 31.52 34.928 31.88 35.12 ; 
        RECT 37.136 34.928 37.208 35.12 ; 
        RECT 65.576 34.928 65.648 35.12 ; 
        RECT 0.488 39.248 0.56 39.44 ; 
        RECT 28.928 39.248 29 39.44 ; 
        RECT 31.52 39.248 31.88 39.44 ; 
        RECT 37.136 39.248 37.208 39.44 ; 
        RECT 65.576 39.248 65.648 39.44 ; 
        RECT 0.488 43.568 0.56 43.76 ; 
        RECT 28.928 43.568 29 43.76 ; 
        RECT 31.52 43.568 31.88 43.76 ; 
        RECT 37.136 43.568 37.208 43.76 ; 
        RECT 65.576 43.568 65.648 43.76 ; 
        RECT 0.488 47.888 0.56 48.08 ; 
        RECT 28.928 47.888 29 48.08 ; 
        RECT 31.52 47.888 31.88 48.08 ; 
        RECT 37.136 47.888 37.208 48.08 ; 
        RECT 65.576 47.888 65.648 48.08 ; 
        RECT 0.488 52.208 0.56 52.4 ; 
        RECT 28.928 52.208 29 52.4 ; 
        RECT 31.52 52.208 31.88 52.4 ; 
        RECT 37.136 52.208 37.208 52.4 ; 
        RECT 65.576 52.208 65.648 52.4 ; 
        RECT 0.488 56.528 0.56 56.72 ; 
        RECT 28.928 56.528 29 56.72 ; 
        RECT 31.52 56.528 31.88 56.72 ; 
        RECT 37.136 56.528 37.208 56.72 ; 
        RECT 65.576 56.528 65.648 56.72 ; 
        RECT 0.488 60.848 0.56 61.04 ; 
        RECT 28.928 60.848 29 61.04 ; 
        RECT 31.52 60.848 31.88 61.04 ; 
        RECT 37.136 60.848 37.208 61.04 ; 
        RECT 65.576 60.848 65.648 61.04 ; 
        RECT 0.488 65.168 0.56 65.36 ; 
        RECT 28.928 65.168 29 65.36 ; 
        RECT 31.52 65.168 31.88 65.36 ; 
        RECT 37.136 65.168 37.208 65.36 ; 
        RECT 65.576 65.168 65.648 65.36 ; 
        RECT 0.488 69.488 0.56 69.68 ; 
        RECT 28.928 69.488 29 69.68 ; 
        RECT 31.52 69.488 31.88 69.68 ; 
        RECT 37.136 69.488 37.208 69.68 ; 
        RECT 65.576 69.488 65.648 69.68 ; 
        RECT 0.488 73.808 0.56 74 ; 
        RECT 28.928 73.808 29 74 ; 
        RECT 31.52 73.808 31.88 74 ; 
        RECT 37.136 73.808 37.208 74 ; 
        RECT 65.576 73.808 65.648 74 ; 
        RECT 31.66 101.076 31.732 101.94 ; 
        RECT 31.66 88.404 31.732 89.268 ; 
        RECT 31.66 75.732 31.732 76.596 ; 
        RECT 31.868 101.076 31.94 101.94 ; 
        RECT 31.868 88.404 31.94 89.268 ; 
        RECT 31.868 75.732 31.94 76.596 ; 
        RECT 32.076 101.076 32.148 101.94 ; 
        RECT 32.076 88.404 32.148 89.268 ; 
        RECT 32.076 75.732 32.148 76.596 ; 
        RECT 32.284 101.076 32.356 101.94 ; 
        RECT 32.284 88.404 32.356 89.268 ; 
        RECT 32.284 75.732 32.356 76.596 ; 
        RECT 32.492 101.076 32.564 101.94 ; 
        RECT 32.492 88.404 32.564 89.268 ; 
        RECT 32.492 75.732 32.564 76.596 ; 
        RECT 37.116 74.612 37.188 74.708 ; 
        RECT 37.188 89.748 37.26 89.844 ; 
        RECT 0.488 110.636 0.56 110.828 ; 
        RECT 28.928 110.636 29 110.828 ; 
        RECT 31.52 110.636 31.88 110.828 ; 
        RECT 37.136 110.636 37.208 110.828 ; 
        RECT 65.576 110.636 65.648 110.828 ; 
        RECT 0.488 114.956 0.56 115.148 ; 
        RECT 28.928 114.956 29 115.148 ; 
        RECT 31.52 114.956 31.88 115.148 ; 
        RECT 37.136 114.956 37.208 115.148 ; 
        RECT 65.576 114.956 65.648 115.148 ; 
        RECT 0.488 119.276 0.56 119.468 ; 
        RECT 28.928 119.276 29 119.468 ; 
        RECT 31.52 119.276 31.88 119.468 ; 
        RECT 37.136 119.276 37.208 119.468 ; 
        RECT 65.576 119.276 65.648 119.468 ; 
        RECT 0.488 123.596 0.56 123.788 ; 
        RECT 28.928 123.596 29 123.788 ; 
        RECT 31.52 123.596 31.88 123.788 ; 
        RECT 37.136 123.596 37.208 123.788 ; 
        RECT 65.576 123.596 65.648 123.788 ; 
        RECT 0.488 127.916 0.56 128.108 ; 
        RECT 28.928 127.916 29 128.108 ; 
        RECT 31.52 127.916 31.88 128.108 ; 
        RECT 37.136 127.916 37.208 128.108 ; 
        RECT 65.576 127.916 65.648 128.108 ; 
        RECT 0.488 132.236 0.56 132.428 ; 
        RECT 28.928 132.236 29 132.428 ; 
        RECT 31.52 132.236 31.88 132.428 ; 
        RECT 37.136 132.236 37.208 132.428 ; 
        RECT 65.576 132.236 65.648 132.428 ; 
        RECT 0.488 136.556 0.56 136.748 ; 
        RECT 28.928 136.556 29 136.748 ; 
        RECT 31.52 136.556 31.88 136.748 ; 
        RECT 37.136 136.556 37.208 136.748 ; 
        RECT 65.576 136.556 65.648 136.748 ; 
        RECT 0.488 140.876 0.56 141.068 ; 
        RECT 28.928 140.876 29 141.068 ; 
        RECT 31.52 140.876 31.88 141.068 ; 
        RECT 37.136 140.876 37.208 141.068 ; 
        RECT 65.576 140.876 65.648 141.068 ; 
        RECT 0.488 145.196 0.56 145.388 ; 
        RECT 28.928 145.196 29 145.388 ; 
        RECT 31.52 145.196 31.88 145.388 ; 
        RECT 37.136 145.196 37.208 145.388 ; 
        RECT 65.576 145.196 65.648 145.388 ; 
        RECT 0.488 149.516 0.56 149.708 ; 
        RECT 28.928 149.516 29 149.708 ; 
        RECT 31.52 149.516 31.88 149.708 ; 
        RECT 37.136 149.516 37.208 149.708 ; 
        RECT 65.576 149.516 65.648 149.708 ; 
        RECT 0.488 153.836 0.56 154.028 ; 
        RECT 28.928 153.836 29 154.028 ; 
        RECT 31.52 153.836 31.88 154.028 ; 
        RECT 37.136 153.836 37.208 154.028 ; 
        RECT 65.576 153.836 65.648 154.028 ; 
        RECT 0.488 158.156 0.56 158.348 ; 
        RECT 28.928 158.156 29 158.348 ; 
        RECT 31.52 158.156 31.88 158.348 ; 
        RECT 37.136 158.156 37.208 158.348 ; 
        RECT 65.576 158.156 65.648 158.348 ; 
        RECT 0.488 162.476 0.56 162.668 ; 
        RECT 28.928 162.476 29 162.668 ; 
        RECT 31.52 162.476 31.88 162.668 ; 
        RECT 37.136 162.476 37.208 162.668 ; 
        RECT 65.576 162.476 65.648 162.668 ; 
        RECT 0.488 166.796 0.56 166.988 ; 
        RECT 28.928 166.796 29 166.988 ; 
        RECT 31.52 166.796 31.88 166.988 ; 
        RECT 37.136 166.796 37.208 166.988 ; 
        RECT 65.576 166.796 65.648 166.988 ; 
        RECT 0.488 171.116 0.56 171.308 ; 
        RECT 28.928 171.116 29 171.308 ; 
        RECT 31.52 171.116 31.88 171.308 ; 
        RECT 37.136 171.116 37.208 171.308 ; 
        RECT 65.576 171.116 65.648 171.308 ; 
        RECT 0.488 175.436 0.56 175.628 ; 
        RECT 28.928 175.436 29 175.628 ; 
        RECT 31.52 175.436 31.88 175.628 ; 
        RECT 37.136 175.436 37.208 175.628 ; 
        RECT 65.576 175.436 65.648 175.628 ; 
        RECT 0.488 179.756 0.56 179.948 ; 
        RECT 28.928 179.756 29 179.948 ; 
        RECT 31.52 179.756 31.88 179.948 ; 
        RECT 37.136 179.756 37.208 179.948 ; 
        RECT 65.576 179.756 65.648 179.948 ; 
      LAYER M5 ; 
        RECT 36.864 74.54 36.96 89.916 ; 
      LAYER V4 ; 
        RECT 36.864 89.748 36.96 89.844 ; 
        RECT 36.864 75.732 36.96 76.596 ; 
        RECT 36.864 74.612 36.96 74.708 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.304 65.748 4.496 ; 
        RECT 0.376 8.624 65.748 8.816 ; 
        RECT 0.376 12.944 65.748 13.136 ; 
        RECT 0.376 17.264 65.748 17.456 ; 
        RECT 0.376 21.584 65.748 21.776 ; 
        RECT 0.376 25.904 65.748 26.096 ; 
        RECT 0.376 30.224 65.748 30.416 ; 
        RECT 0.376 34.544 65.748 34.736 ; 
        RECT 0.376 38.864 65.748 39.056 ; 
        RECT 0.376 43.184 65.748 43.376 ; 
        RECT 0.376 47.504 65.748 47.696 ; 
        RECT 0.376 51.824 65.748 52.016 ; 
        RECT 0.376 56.144 65.748 56.336 ; 
        RECT 0.376 60.464 65.748 60.656 ; 
        RECT 0.376 64.784 65.748 64.976 ; 
        RECT 0.376 69.104 65.748 69.296 ; 
        RECT 0.376 73.424 65.748 73.616 ; 
        RECT 14.256 77.46 51.84 78.324 ; 
        RECT 29.592 90.132 36.504 90.996 ; 
        RECT 29.592 102.804 36.504 103.668 ; 
        RECT 0.376 110.252 65.748 110.444 ; 
        RECT 0.376 114.572 65.748 114.764 ; 
        RECT 0.376 118.892 65.748 119.084 ; 
        RECT 0.376 123.212 65.748 123.404 ; 
        RECT 0.376 127.532 65.748 127.724 ; 
        RECT 0.376 131.852 65.748 132.044 ; 
        RECT 0.376 136.172 65.748 136.364 ; 
        RECT 0.376 140.492 65.748 140.684 ; 
        RECT 0.376 144.812 65.748 145.004 ; 
        RECT 0.376 149.132 65.748 149.324 ; 
        RECT 0.376 153.452 65.748 153.644 ; 
        RECT 0.376 157.772 65.748 157.964 ; 
        RECT 0.376 162.092 65.748 162.284 ; 
        RECT 0.376 166.412 65.748 166.604 ; 
        RECT 0.376 170.732 65.748 170.924 ; 
        RECT 0.376 175.052 65.748 175.244 ; 
        RECT 0.376 179.372 65.748 179.564 ; 
      LAYER M3 ; 
        RECT 65.432 0.866 65.504 5.506 ; 
        RECT 37.352 0.866 37.424 5.506 ; 
        RECT 34.292 1.012 34.436 5.468 ; 
        RECT 33.68 1.012 33.788 5.468 ; 
        RECT 28.712 0.866 28.784 5.506 ; 
        RECT 0.632 0.866 0.704 5.506 ; 
        RECT 65.432 5.186 65.504 9.826 ; 
        RECT 37.352 5.186 37.424 9.826 ; 
        RECT 34.292 5.332 34.436 9.788 ; 
        RECT 33.68 5.332 33.788 9.788 ; 
        RECT 28.712 5.186 28.784 9.826 ; 
        RECT 0.632 5.186 0.704 9.826 ; 
        RECT 65.432 9.506 65.504 14.146 ; 
        RECT 37.352 9.506 37.424 14.146 ; 
        RECT 34.292 9.652 34.436 14.108 ; 
        RECT 33.68 9.652 33.788 14.108 ; 
        RECT 28.712 9.506 28.784 14.146 ; 
        RECT 0.632 9.506 0.704 14.146 ; 
        RECT 65.432 13.826 65.504 18.466 ; 
        RECT 37.352 13.826 37.424 18.466 ; 
        RECT 34.292 13.972 34.436 18.428 ; 
        RECT 33.68 13.972 33.788 18.428 ; 
        RECT 28.712 13.826 28.784 18.466 ; 
        RECT 0.632 13.826 0.704 18.466 ; 
        RECT 65.432 18.146 65.504 22.786 ; 
        RECT 37.352 18.146 37.424 22.786 ; 
        RECT 34.292 18.292 34.436 22.748 ; 
        RECT 33.68 18.292 33.788 22.748 ; 
        RECT 28.712 18.146 28.784 22.786 ; 
        RECT 0.632 18.146 0.704 22.786 ; 
        RECT 65.432 22.466 65.504 27.106 ; 
        RECT 37.352 22.466 37.424 27.106 ; 
        RECT 34.292 22.612 34.436 27.068 ; 
        RECT 33.68 22.612 33.788 27.068 ; 
        RECT 28.712 22.466 28.784 27.106 ; 
        RECT 0.632 22.466 0.704 27.106 ; 
        RECT 65.432 26.786 65.504 31.426 ; 
        RECT 37.352 26.786 37.424 31.426 ; 
        RECT 34.292 26.932 34.436 31.388 ; 
        RECT 33.68 26.932 33.788 31.388 ; 
        RECT 28.712 26.786 28.784 31.426 ; 
        RECT 0.632 26.786 0.704 31.426 ; 
        RECT 65.432 31.106 65.504 35.746 ; 
        RECT 37.352 31.106 37.424 35.746 ; 
        RECT 34.292 31.252 34.436 35.708 ; 
        RECT 33.68 31.252 33.788 35.708 ; 
        RECT 28.712 31.106 28.784 35.746 ; 
        RECT 0.632 31.106 0.704 35.746 ; 
        RECT 65.432 35.426 65.504 40.066 ; 
        RECT 37.352 35.426 37.424 40.066 ; 
        RECT 34.292 35.572 34.436 40.028 ; 
        RECT 33.68 35.572 33.788 40.028 ; 
        RECT 28.712 35.426 28.784 40.066 ; 
        RECT 0.632 35.426 0.704 40.066 ; 
        RECT 65.432 39.746 65.504 44.386 ; 
        RECT 37.352 39.746 37.424 44.386 ; 
        RECT 34.292 39.892 34.436 44.348 ; 
        RECT 33.68 39.892 33.788 44.348 ; 
        RECT 28.712 39.746 28.784 44.386 ; 
        RECT 0.632 39.746 0.704 44.386 ; 
        RECT 65.432 44.066 65.504 48.706 ; 
        RECT 37.352 44.066 37.424 48.706 ; 
        RECT 34.292 44.212 34.436 48.668 ; 
        RECT 33.68 44.212 33.788 48.668 ; 
        RECT 28.712 44.066 28.784 48.706 ; 
        RECT 0.632 44.066 0.704 48.706 ; 
        RECT 65.432 48.386 65.504 53.026 ; 
        RECT 37.352 48.386 37.424 53.026 ; 
        RECT 34.292 48.532 34.436 52.988 ; 
        RECT 33.68 48.532 33.788 52.988 ; 
        RECT 28.712 48.386 28.784 53.026 ; 
        RECT 0.632 48.386 0.704 53.026 ; 
        RECT 65.432 52.706 65.504 57.346 ; 
        RECT 37.352 52.706 37.424 57.346 ; 
        RECT 34.292 52.852 34.436 57.308 ; 
        RECT 33.68 52.852 33.788 57.308 ; 
        RECT 28.712 52.706 28.784 57.346 ; 
        RECT 0.632 52.706 0.704 57.346 ; 
        RECT 65.432 57.026 65.504 61.666 ; 
        RECT 37.352 57.026 37.424 61.666 ; 
        RECT 34.292 57.172 34.436 61.628 ; 
        RECT 33.68 57.172 33.788 61.628 ; 
        RECT 28.712 57.026 28.784 61.666 ; 
        RECT 0.632 57.026 0.704 61.666 ; 
        RECT 65.432 61.346 65.504 65.986 ; 
        RECT 37.352 61.346 37.424 65.986 ; 
        RECT 34.292 61.492 34.436 65.948 ; 
        RECT 33.68 61.492 33.788 65.948 ; 
        RECT 28.712 61.346 28.784 65.986 ; 
        RECT 0.632 61.346 0.704 65.986 ; 
        RECT 65.432 65.666 65.504 70.306 ; 
        RECT 37.352 65.666 37.424 70.306 ; 
        RECT 34.292 65.812 34.436 70.268 ; 
        RECT 33.68 65.812 33.788 70.268 ; 
        RECT 28.712 65.666 28.784 70.306 ; 
        RECT 0.632 65.666 0.704 70.306 ; 
        RECT 65.432 69.986 65.504 74.626 ; 
        RECT 37.352 69.986 37.424 74.626 ; 
        RECT 34.292 70.132 34.436 74.588 ; 
        RECT 33.68 70.132 33.788 74.588 ; 
        RECT 28.712 69.986 28.784 74.626 ; 
        RECT 0.632 69.986 0.704 74.626 ; 
        RECT 65.412 74.282 65.484 107.11 ; 
        RECT 37.332 74.282 37.404 107.11 ; 
        RECT 33.516 75.176 34.452 105.908 ; 
        RECT 34.272 74.458 34.416 106.936 ; 
        RECT 33.66 74.456 33.768 106.936 ; 
        RECT 28.692 74.282 28.764 107.11 ; 
        RECT 0.612 74.282 0.684 107.11 ; 
        RECT 65.432 106.814 65.504 111.454 ; 
        RECT 37.352 106.814 37.424 111.454 ; 
        RECT 34.292 106.96 34.436 111.416 ; 
        RECT 33.68 106.96 33.788 111.416 ; 
        RECT 28.712 106.814 28.784 111.454 ; 
        RECT 0.632 106.814 0.704 111.454 ; 
        RECT 65.432 111.134 65.504 115.774 ; 
        RECT 37.352 111.134 37.424 115.774 ; 
        RECT 34.292 111.28 34.436 115.736 ; 
        RECT 33.68 111.28 33.788 115.736 ; 
        RECT 28.712 111.134 28.784 115.774 ; 
        RECT 0.632 111.134 0.704 115.774 ; 
        RECT 65.432 115.454 65.504 120.094 ; 
        RECT 37.352 115.454 37.424 120.094 ; 
        RECT 34.292 115.6 34.436 120.056 ; 
        RECT 33.68 115.6 33.788 120.056 ; 
        RECT 28.712 115.454 28.784 120.094 ; 
        RECT 0.632 115.454 0.704 120.094 ; 
        RECT 65.432 119.774 65.504 124.414 ; 
        RECT 37.352 119.774 37.424 124.414 ; 
        RECT 34.292 119.92 34.436 124.376 ; 
        RECT 33.68 119.92 33.788 124.376 ; 
        RECT 28.712 119.774 28.784 124.414 ; 
        RECT 0.632 119.774 0.704 124.414 ; 
        RECT 65.432 124.094 65.504 128.734 ; 
        RECT 37.352 124.094 37.424 128.734 ; 
        RECT 34.292 124.24 34.436 128.696 ; 
        RECT 33.68 124.24 33.788 128.696 ; 
        RECT 28.712 124.094 28.784 128.734 ; 
        RECT 0.632 124.094 0.704 128.734 ; 
        RECT 65.432 128.414 65.504 133.054 ; 
        RECT 37.352 128.414 37.424 133.054 ; 
        RECT 34.292 128.56 34.436 133.016 ; 
        RECT 33.68 128.56 33.788 133.016 ; 
        RECT 28.712 128.414 28.784 133.054 ; 
        RECT 0.632 128.414 0.704 133.054 ; 
        RECT 65.432 132.734 65.504 137.374 ; 
        RECT 37.352 132.734 37.424 137.374 ; 
        RECT 34.292 132.88 34.436 137.336 ; 
        RECT 33.68 132.88 33.788 137.336 ; 
        RECT 28.712 132.734 28.784 137.374 ; 
        RECT 0.632 132.734 0.704 137.374 ; 
        RECT 65.432 137.054 65.504 141.694 ; 
        RECT 37.352 137.054 37.424 141.694 ; 
        RECT 34.292 137.2 34.436 141.656 ; 
        RECT 33.68 137.2 33.788 141.656 ; 
        RECT 28.712 137.054 28.784 141.694 ; 
        RECT 0.632 137.054 0.704 141.694 ; 
        RECT 65.432 141.374 65.504 146.014 ; 
        RECT 37.352 141.374 37.424 146.014 ; 
        RECT 34.292 141.52 34.436 145.976 ; 
        RECT 33.68 141.52 33.788 145.976 ; 
        RECT 28.712 141.374 28.784 146.014 ; 
        RECT 0.632 141.374 0.704 146.014 ; 
        RECT 65.432 145.694 65.504 150.334 ; 
        RECT 37.352 145.694 37.424 150.334 ; 
        RECT 34.292 145.84 34.436 150.296 ; 
        RECT 33.68 145.84 33.788 150.296 ; 
        RECT 28.712 145.694 28.784 150.334 ; 
        RECT 0.632 145.694 0.704 150.334 ; 
        RECT 65.432 150.014 65.504 154.654 ; 
        RECT 37.352 150.014 37.424 154.654 ; 
        RECT 34.292 150.16 34.436 154.616 ; 
        RECT 33.68 150.16 33.788 154.616 ; 
        RECT 28.712 150.014 28.784 154.654 ; 
        RECT 0.632 150.014 0.704 154.654 ; 
        RECT 65.432 154.334 65.504 158.974 ; 
        RECT 37.352 154.334 37.424 158.974 ; 
        RECT 34.292 154.48 34.436 158.936 ; 
        RECT 33.68 154.48 33.788 158.936 ; 
        RECT 28.712 154.334 28.784 158.974 ; 
        RECT 0.632 154.334 0.704 158.974 ; 
        RECT 65.432 158.654 65.504 163.294 ; 
        RECT 37.352 158.654 37.424 163.294 ; 
        RECT 34.292 158.8 34.436 163.256 ; 
        RECT 33.68 158.8 33.788 163.256 ; 
        RECT 28.712 158.654 28.784 163.294 ; 
        RECT 0.632 158.654 0.704 163.294 ; 
        RECT 65.432 162.974 65.504 167.614 ; 
        RECT 37.352 162.974 37.424 167.614 ; 
        RECT 34.292 163.12 34.436 167.576 ; 
        RECT 33.68 163.12 33.788 167.576 ; 
        RECT 28.712 162.974 28.784 167.614 ; 
        RECT 0.632 162.974 0.704 167.614 ; 
        RECT 65.432 167.294 65.504 171.934 ; 
        RECT 37.352 167.294 37.424 171.934 ; 
        RECT 34.292 167.44 34.436 171.896 ; 
        RECT 33.68 167.44 33.788 171.896 ; 
        RECT 28.712 167.294 28.784 171.934 ; 
        RECT 0.632 167.294 0.704 171.934 ; 
        RECT 65.432 171.614 65.504 176.254 ; 
        RECT 37.352 171.614 37.424 176.254 ; 
        RECT 34.292 171.76 34.436 176.216 ; 
        RECT 33.68 171.76 33.788 176.216 ; 
        RECT 28.712 171.614 28.784 176.254 ; 
        RECT 0.632 171.614 0.704 176.254 ; 
        RECT 65.432 175.934 65.504 180.574 ; 
        RECT 37.352 175.934 37.424 180.574 ; 
        RECT 34.292 176.08 34.436 180.536 ; 
        RECT 33.68 176.08 33.788 180.536 ; 
        RECT 28.712 175.934 28.784 180.574 ; 
        RECT 0.632 175.934 0.704 180.574 ; 
      LAYER V3 ; 
        RECT 0.632 4.304 0.704 4.496 ; 
        RECT 28.712 4.304 28.784 4.496 ; 
        RECT 33.68 4.304 33.788 4.496 ; 
        RECT 34.292 4.304 34.436 4.496 ; 
        RECT 37.352 4.304 37.424 4.496 ; 
        RECT 65.432 4.304 65.504 4.496 ; 
        RECT 0.632 8.624 0.704 8.816 ; 
        RECT 28.712 8.624 28.784 8.816 ; 
        RECT 33.68 8.624 33.788 8.816 ; 
        RECT 34.292 8.624 34.436 8.816 ; 
        RECT 37.352 8.624 37.424 8.816 ; 
        RECT 65.432 8.624 65.504 8.816 ; 
        RECT 0.632 12.944 0.704 13.136 ; 
        RECT 28.712 12.944 28.784 13.136 ; 
        RECT 33.68 12.944 33.788 13.136 ; 
        RECT 34.292 12.944 34.436 13.136 ; 
        RECT 37.352 12.944 37.424 13.136 ; 
        RECT 65.432 12.944 65.504 13.136 ; 
        RECT 0.632 17.264 0.704 17.456 ; 
        RECT 28.712 17.264 28.784 17.456 ; 
        RECT 33.68 17.264 33.788 17.456 ; 
        RECT 34.292 17.264 34.436 17.456 ; 
        RECT 37.352 17.264 37.424 17.456 ; 
        RECT 65.432 17.264 65.504 17.456 ; 
        RECT 0.632 21.584 0.704 21.776 ; 
        RECT 28.712 21.584 28.784 21.776 ; 
        RECT 33.68 21.584 33.788 21.776 ; 
        RECT 34.292 21.584 34.436 21.776 ; 
        RECT 37.352 21.584 37.424 21.776 ; 
        RECT 65.432 21.584 65.504 21.776 ; 
        RECT 0.632 25.904 0.704 26.096 ; 
        RECT 28.712 25.904 28.784 26.096 ; 
        RECT 33.68 25.904 33.788 26.096 ; 
        RECT 34.292 25.904 34.436 26.096 ; 
        RECT 37.352 25.904 37.424 26.096 ; 
        RECT 65.432 25.904 65.504 26.096 ; 
        RECT 0.632 30.224 0.704 30.416 ; 
        RECT 28.712 30.224 28.784 30.416 ; 
        RECT 33.68 30.224 33.788 30.416 ; 
        RECT 34.292 30.224 34.436 30.416 ; 
        RECT 37.352 30.224 37.424 30.416 ; 
        RECT 65.432 30.224 65.504 30.416 ; 
        RECT 0.632 34.544 0.704 34.736 ; 
        RECT 28.712 34.544 28.784 34.736 ; 
        RECT 33.68 34.544 33.788 34.736 ; 
        RECT 34.292 34.544 34.436 34.736 ; 
        RECT 37.352 34.544 37.424 34.736 ; 
        RECT 65.432 34.544 65.504 34.736 ; 
        RECT 0.632 38.864 0.704 39.056 ; 
        RECT 28.712 38.864 28.784 39.056 ; 
        RECT 33.68 38.864 33.788 39.056 ; 
        RECT 34.292 38.864 34.436 39.056 ; 
        RECT 37.352 38.864 37.424 39.056 ; 
        RECT 65.432 38.864 65.504 39.056 ; 
        RECT 0.632 43.184 0.704 43.376 ; 
        RECT 28.712 43.184 28.784 43.376 ; 
        RECT 33.68 43.184 33.788 43.376 ; 
        RECT 34.292 43.184 34.436 43.376 ; 
        RECT 37.352 43.184 37.424 43.376 ; 
        RECT 65.432 43.184 65.504 43.376 ; 
        RECT 0.632 47.504 0.704 47.696 ; 
        RECT 28.712 47.504 28.784 47.696 ; 
        RECT 33.68 47.504 33.788 47.696 ; 
        RECT 34.292 47.504 34.436 47.696 ; 
        RECT 37.352 47.504 37.424 47.696 ; 
        RECT 65.432 47.504 65.504 47.696 ; 
        RECT 0.632 51.824 0.704 52.016 ; 
        RECT 28.712 51.824 28.784 52.016 ; 
        RECT 33.68 51.824 33.788 52.016 ; 
        RECT 34.292 51.824 34.436 52.016 ; 
        RECT 37.352 51.824 37.424 52.016 ; 
        RECT 65.432 51.824 65.504 52.016 ; 
        RECT 0.632 56.144 0.704 56.336 ; 
        RECT 28.712 56.144 28.784 56.336 ; 
        RECT 33.68 56.144 33.788 56.336 ; 
        RECT 34.292 56.144 34.436 56.336 ; 
        RECT 37.352 56.144 37.424 56.336 ; 
        RECT 65.432 56.144 65.504 56.336 ; 
        RECT 0.632 60.464 0.704 60.656 ; 
        RECT 28.712 60.464 28.784 60.656 ; 
        RECT 33.68 60.464 33.788 60.656 ; 
        RECT 34.292 60.464 34.436 60.656 ; 
        RECT 37.352 60.464 37.424 60.656 ; 
        RECT 65.432 60.464 65.504 60.656 ; 
        RECT 0.632 64.784 0.704 64.976 ; 
        RECT 28.712 64.784 28.784 64.976 ; 
        RECT 33.68 64.784 33.788 64.976 ; 
        RECT 34.292 64.784 34.436 64.976 ; 
        RECT 37.352 64.784 37.424 64.976 ; 
        RECT 65.432 64.784 65.504 64.976 ; 
        RECT 0.632 69.104 0.704 69.296 ; 
        RECT 28.712 69.104 28.784 69.296 ; 
        RECT 33.68 69.104 33.788 69.296 ; 
        RECT 34.292 69.104 34.436 69.296 ; 
        RECT 37.352 69.104 37.424 69.296 ; 
        RECT 65.432 69.104 65.504 69.296 ; 
        RECT 0.632 73.424 0.704 73.616 ; 
        RECT 28.712 73.424 28.784 73.616 ; 
        RECT 33.68 73.424 33.788 73.616 ; 
        RECT 34.292 73.424 34.436 73.616 ; 
        RECT 37.352 73.424 37.424 73.616 ; 
        RECT 65.432 73.424 65.504 73.616 ; 
        RECT 33.532 102.804 33.604 103.668 ; 
        RECT 33.532 90.132 33.604 90.996 ; 
        RECT 33.532 77.46 33.604 78.324 ; 
        RECT 33.74 102.804 33.812 103.668 ; 
        RECT 33.74 90.132 33.812 90.996 ; 
        RECT 33.74 77.46 33.812 78.324 ; 
        RECT 33.948 102.804 34.02 103.668 ; 
        RECT 33.948 90.132 34.02 90.996 ; 
        RECT 33.948 77.46 34.02 78.324 ; 
        RECT 34.156 102.804 34.228 103.668 ; 
        RECT 34.156 90.132 34.228 90.996 ; 
        RECT 34.156 77.46 34.228 78.324 ; 
        RECT 34.364 102.804 34.436 103.668 ; 
        RECT 34.364 90.132 34.436 90.996 ; 
        RECT 34.364 77.46 34.436 78.324 ; 
        RECT 37.332 77.462 37.404 78.326 ; 
        RECT 0.632 110.252 0.704 110.444 ; 
        RECT 28.712 110.252 28.784 110.444 ; 
        RECT 33.68 110.252 33.788 110.444 ; 
        RECT 34.292 110.252 34.436 110.444 ; 
        RECT 37.352 110.252 37.424 110.444 ; 
        RECT 65.432 110.252 65.504 110.444 ; 
        RECT 0.632 114.572 0.704 114.764 ; 
        RECT 28.712 114.572 28.784 114.764 ; 
        RECT 33.68 114.572 33.788 114.764 ; 
        RECT 34.292 114.572 34.436 114.764 ; 
        RECT 37.352 114.572 37.424 114.764 ; 
        RECT 65.432 114.572 65.504 114.764 ; 
        RECT 0.632 118.892 0.704 119.084 ; 
        RECT 28.712 118.892 28.784 119.084 ; 
        RECT 33.68 118.892 33.788 119.084 ; 
        RECT 34.292 118.892 34.436 119.084 ; 
        RECT 37.352 118.892 37.424 119.084 ; 
        RECT 65.432 118.892 65.504 119.084 ; 
        RECT 0.632 123.212 0.704 123.404 ; 
        RECT 28.712 123.212 28.784 123.404 ; 
        RECT 33.68 123.212 33.788 123.404 ; 
        RECT 34.292 123.212 34.436 123.404 ; 
        RECT 37.352 123.212 37.424 123.404 ; 
        RECT 65.432 123.212 65.504 123.404 ; 
        RECT 0.632 127.532 0.704 127.724 ; 
        RECT 28.712 127.532 28.784 127.724 ; 
        RECT 33.68 127.532 33.788 127.724 ; 
        RECT 34.292 127.532 34.436 127.724 ; 
        RECT 37.352 127.532 37.424 127.724 ; 
        RECT 65.432 127.532 65.504 127.724 ; 
        RECT 0.632 131.852 0.704 132.044 ; 
        RECT 28.712 131.852 28.784 132.044 ; 
        RECT 33.68 131.852 33.788 132.044 ; 
        RECT 34.292 131.852 34.436 132.044 ; 
        RECT 37.352 131.852 37.424 132.044 ; 
        RECT 65.432 131.852 65.504 132.044 ; 
        RECT 0.632 136.172 0.704 136.364 ; 
        RECT 28.712 136.172 28.784 136.364 ; 
        RECT 33.68 136.172 33.788 136.364 ; 
        RECT 34.292 136.172 34.436 136.364 ; 
        RECT 37.352 136.172 37.424 136.364 ; 
        RECT 65.432 136.172 65.504 136.364 ; 
        RECT 0.632 140.492 0.704 140.684 ; 
        RECT 28.712 140.492 28.784 140.684 ; 
        RECT 33.68 140.492 33.788 140.684 ; 
        RECT 34.292 140.492 34.436 140.684 ; 
        RECT 37.352 140.492 37.424 140.684 ; 
        RECT 65.432 140.492 65.504 140.684 ; 
        RECT 0.632 144.812 0.704 145.004 ; 
        RECT 28.712 144.812 28.784 145.004 ; 
        RECT 33.68 144.812 33.788 145.004 ; 
        RECT 34.292 144.812 34.436 145.004 ; 
        RECT 37.352 144.812 37.424 145.004 ; 
        RECT 65.432 144.812 65.504 145.004 ; 
        RECT 0.632 149.132 0.704 149.324 ; 
        RECT 28.712 149.132 28.784 149.324 ; 
        RECT 33.68 149.132 33.788 149.324 ; 
        RECT 34.292 149.132 34.436 149.324 ; 
        RECT 37.352 149.132 37.424 149.324 ; 
        RECT 65.432 149.132 65.504 149.324 ; 
        RECT 0.632 153.452 0.704 153.644 ; 
        RECT 28.712 153.452 28.784 153.644 ; 
        RECT 33.68 153.452 33.788 153.644 ; 
        RECT 34.292 153.452 34.436 153.644 ; 
        RECT 37.352 153.452 37.424 153.644 ; 
        RECT 65.432 153.452 65.504 153.644 ; 
        RECT 0.632 157.772 0.704 157.964 ; 
        RECT 28.712 157.772 28.784 157.964 ; 
        RECT 33.68 157.772 33.788 157.964 ; 
        RECT 34.292 157.772 34.436 157.964 ; 
        RECT 37.352 157.772 37.424 157.964 ; 
        RECT 65.432 157.772 65.504 157.964 ; 
        RECT 0.632 162.092 0.704 162.284 ; 
        RECT 28.712 162.092 28.784 162.284 ; 
        RECT 33.68 162.092 33.788 162.284 ; 
        RECT 34.292 162.092 34.436 162.284 ; 
        RECT 37.352 162.092 37.424 162.284 ; 
        RECT 65.432 162.092 65.504 162.284 ; 
        RECT 0.632 166.412 0.704 166.604 ; 
        RECT 28.712 166.412 28.784 166.604 ; 
        RECT 33.68 166.412 33.788 166.604 ; 
        RECT 34.292 166.412 34.436 166.604 ; 
        RECT 37.352 166.412 37.424 166.604 ; 
        RECT 65.432 166.412 65.504 166.604 ; 
        RECT 0.632 170.732 0.704 170.924 ; 
        RECT 28.712 170.732 28.784 170.924 ; 
        RECT 33.68 170.732 33.788 170.924 ; 
        RECT 34.292 170.732 34.436 170.924 ; 
        RECT 37.352 170.732 37.424 170.924 ; 
        RECT 65.432 170.732 65.504 170.924 ; 
        RECT 0.632 175.052 0.704 175.244 ; 
        RECT 28.712 175.052 28.784 175.244 ; 
        RECT 33.68 175.052 33.788 175.244 ; 
        RECT 34.292 175.052 34.436 175.244 ; 
        RECT 37.352 175.052 37.424 175.244 ; 
        RECT 65.432 175.052 65.504 175.244 ; 
        RECT 0.632 179.372 0.704 179.564 ; 
        RECT 28.712 179.372 28.784 179.564 ; 
        RECT 33.68 179.372 33.788 179.564 ; 
        RECT 34.292 179.372 34.436 179.564 ; 
        RECT 37.352 179.372 37.424 179.564 ; 
        RECT 65.432 179.372 65.504 179.564 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 43.164 79.348 43.236 79.496 ; 
      LAYER M4 ; 
        RECT 42.956 79.38 43.292 79.476 ; 
      LAYER M5 ; 
        RECT 43.152 75.576 43.248 88.536 ; 
      LAYER V3 ; 
        RECT 43.164 79.38 43.236 79.476 ; 
      LAYER V4 ; 
        RECT 43.152 79.38 43.248 79.476 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 42.3 79.36 42.372 79.508 ; 
      LAYER M4 ; 
        RECT 42.092 79.38 42.428 79.476 ; 
      LAYER M5 ; 
        RECT 42.288 75.576 42.384 88.536 ; 
      LAYER V3 ; 
        RECT 42.3 79.38 42.372 79.476 ; 
      LAYER V4 ; 
        RECT 42.288 79.38 42.384 79.476 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 41.436 77.044 41.508 77.192 ; 
      LAYER M4 ; 
        RECT 41.228 77.076 41.564 77.172 ; 
      LAYER M5 ; 
        RECT 41.424 75.576 41.52 88.536 ; 
      LAYER V3 ; 
        RECT 41.436 77.076 41.508 77.172 ; 
      LAYER V4 ; 
        RECT 41.424 77.076 41.52 77.172 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 40.572 78.004 40.644 78.728 ; 
      LAYER M4 ; 
        RECT 40.364 78.612 40.7 78.708 ; 
      LAYER M5 ; 
        RECT 40.56 75.576 40.656 88.536 ; 
      LAYER V3 ; 
        RECT 40.572 78.612 40.644 78.708 ; 
      LAYER V4 ; 
        RECT 40.56 78.612 40.656 78.708 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 39.708 77.056 39.78 77.324 ; 
      LAYER M4 ; 
        RECT 39.5 77.076 39.836 77.172 ; 
      LAYER M5 ; 
        RECT 39.696 75.576 39.792 88.536 ; 
      LAYER V3 ; 
        RECT 39.708 77.076 39.78 77.172 ; 
      LAYER V4 ; 
        RECT 39.696 77.076 39.792 77.172 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 38.844 75.988 38.916 77 ; 
      LAYER M4 ; 
        RECT 38.636 76.884 38.972 76.98 ; 
      LAYER M5 ; 
        RECT 38.832 75.576 38.928 88.536 ; 
      LAYER V3 ; 
        RECT 38.844 76.884 38.916 76.98 ; 
      LAYER V4 ; 
        RECT 38.832 76.884 38.928 76.98 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.98 80.128 38.052 80.276 ; 
      LAYER M4 ; 
        RECT 37.772 80.148 38.108 80.244 ; 
      LAYER M5 ; 
        RECT 37.968 75.576 38.064 88.536 ; 
      LAYER V3 ; 
        RECT 37.98 80.148 38.052 80.244 ; 
      LAYER V4 ; 
        RECT 37.968 80.148 38.064 80.244 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.116 79.516 37.188 79.88 ; 
      LAYER M4 ; 
        RECT 36.908 79.764 37.244 79.86 ; 
      LAYER M5 ; 
        RECT 37.104 75.576 37.2 88.536 ; 
      LAYER V3 ; 
        RECT 37.116 79.764 37.188 79.86 ; 
      LAYER V4 ; 
        RECT 37.104 79.764 37.2 79.86 ; 
    END 
  END ADDRESS[7] 
  PIN ADDRESS[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 34.524 77.056 34.596 77.324 ; 
      LAYER M4 ; 
        RECT 33.388 77.076 34.64 77.172 ; 
      LAYER M5 ; 
        RECT 33.432 75.576 33.528 88.536 ; 
      LAYER V3 ; 
        RECT 34.524 77.076 34.596 77.172 ; 
      LAYER V4 ; 
        RECT 33.432 77.076 33.528 77.172 ; 
    END 
  END ADDRESS[8] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 32.94 75.988 33.012 77 ; 
      LAYER M4 ; 
        RECT 32.092 76.884 33.056 76.98 ; 
      LAYER M5 ; 
        RECT 32.136 75.576 32.232 88.536 ; 
      LAYER V3 ; 
        RECT 32.94 76.884 33.012 76.98 ; 
      LAYER V4 ; 
        RECT 32.136 76.884 32.232 76.98 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.772 77.056 29.844 77.324 ; 
      LAYER M4 ; 
        RECT 29.564 77.076 29.9 77.172 ; 
      LAYER M5 ; 
        RECT 29.76 75.576 29.856 88.536 ; 
      LAYER V3 ; 
        RECT 29.772 77.076 29.844 77.172 ; 
      LAYER V4 ; 
        RECT 29.76 77.076 29.856 77.172 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.908 80.512 28.98 80.708 ; 
      LAYER M4 ; 
        RECT 28.7 80.532 29.036 80.628 ; 
      LAYER M5 ; 
        RECT 28.896 75.576 28.992 88.536 ; 
      LAYER V3 ; 
        RECT 28.908 80.532 28.98 80.628 ; 
      LAYER V4 ; 
        RECT 28.896 80.532 28.992 80.628 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.052 75.988 29.124 77 ; 
      LAYER M4 ; 
        RECT 27.988 76.884 29.168 76.98 ; 
      LAYER M5 ; 
        RECT 28.032 75.576 28.128 88.536 ; 
      LAYER V3 ; 
        RECT 29.052 76.884 29.124 76.98 ; 
      LAYER V4 ; 
        RECT 28.032 76.884 28.128 76.98 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.18 79.348 27.252 79.496 ; 
      LAYER M4 ; 
        RECT 26.972 79.38 27.308 79.476 ; 
      LAYER M5 ; 
        RECT 27.168 75.576 27.264 88.536 ; 
      LAYER V3 ; 
        RECT 27.18 79.38 27.252 79.476 ; 
      LAYER V4 ; 
        RECT 27.168 79.38 27.264 79.476 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.316 77.056 26.388 77.972 ; 
      LAYER M4 ; 
        RECT 26.108 77.076 26.444 77.172 ; 
      LAYER M5 ; 
        RECT 26.304 75.576 26.4 88.536 ; 
      LAYER V3 ; 
        RECT 26.316 77.076 26.388 77.172 ; 
      LAYER V4 ; 
        RECT 26.304 77.076 26.4 77.172 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.452 75.988 25.524 77 ; 
      LAYER M4 ; 
        RECT 25.244 76.884 25.58 76.98 ; 
      LAYER M5 ; 
        RECT 25.44 75.576 25.536 88.536 ; 
      LAYER V3 ; 
        RECT 25.452 76.884 25.524 76.98 ; 
      LAYER V4 ; 
        RECT 25.44 76.884 25.536 76.98 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.588 77.044 24.66 77.192 ; 
      LAYER M4 ; 
        RECT 24.38 77.076 24.716 77.172 ; 
      LAYER M5 ; 
        RECT 24.576 75.576 24.672 88.536 ; 
      LAYER V3 ; 
        RECT 24.588 77.076 24.66 77.172 ; 
      LAYER V4 ; 
        RECT 24.576 77.076 24.672 77.172 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 23.724 79.348 23.796 79.496 ; 
      LAYER M4 ; 
        RECT 23.516 79.38 23.852 79.476 ; 
      LAYER M5 ; 
        RECT 23.712 75.576 23.808 88.536 ; 
      LAYER V3 ; 
        RECT 23.724 79.38 23.796 79.476 ; 
      LAYER V4 ; 
        RECT 23.712 79.38 23.808 79.476 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.712 34.388 1.808 ; 
      LAYER M3 ; 
        RECT 34.148 1.51 34.22 2.468 ; 
      LAYER V3 ; 
        RECT 34.148 1.712 34.22 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.328 34.66 1.424 ; 
      LAYER M3 ; 
        RECT 33.248 1.08 33.32 2.7 ; 
      LAYER V3 ; 
        RECT 33.248 1.328 33.32 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 6.032 34.388 6.128 ; 
      LAYER M3 ; 
        RECT 34.148 5.83 34.22 6.788 ; 
      LAYER V3 ; 
        RECT 34.148 6.032 34.22 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 5.648 34.66 5.744 ; 
      LAYER M3 ; 
        RECT 33.248 5.4 33.32 7.02 ; 
      LAYER V3 ; 
        RECT 33.248 5.648 33.32 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 10.352 34.388 10.448 ; 
      LAYER M3 ; 
        RECT 34.148 10.15 34.22 11.108 ; 
      LAYER V3 ; 
        RECT 34.148 10.352 34.22 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 9.968 34.66 10.064 ; 
      LAYER M3 ; 
        RECT 33.248 9.72 33.32 11.34 ; 
      LAYER V3 ; 
        RECT 33.248 9.968 33.32 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.672 34.388 14.768 ; 
      LAYER M3 ; 
        RECT 34.148 14.47 34.22 15.428 ; 
      LAYER V3 ; 
        RECT 34.148 14.672 34.22 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.288 34.66 14.384 ; 
      LAYER M3 ; 
        RECT 33.248 14.04 33.32 15.66 ; 
      LAYER V3 ; 
        RECT 33.248 14.288 33.32 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.992 34.388 19.088 ; 
      LAYER M3 ; 
        RECT 34.148 18.79 34.22 19.748 ; 
      LAYER V3 ; 
        RECT 34.148 18.992 34.22 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.608 34.66 18.704 ; 
      LAYER M3 ; 
        RECT 33.248 18.36 33.32 19.98 ; 
      LAYER V3 ; 
        RECT 33.248 18.608 33.32 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 23.312 34.388 23.408 ; 
      LAYER M3 ; 
        RECT 34.148 23.11 34.22 24.068 ; 
      LAYER V3 ; 
        RECT 34.148 23.312 34.22 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 22.928 34.66 23.024 ; 
      LAYER M3 ; 
        RECT 33.248 22.68 33.32 24.3 ; 
      LAYER V3 ; 
        RECT 33.248 22.928 33.32 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.632 34.388 27.728 ; 
      LAYER M3 ; 
        RECT 34.148 27.43 34.22 28.388 ; 
      LAYER V3 ; 
        RECT 34.148 27.632 34.22 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.248 34.66 27.344 ; 
      LAYER M3 ; 
        RECT 33.248 27 33.32 28.62 ; 
      LAYER V3 ; 
        RECT 33.248 27.248 33.32 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.952 34.388 32.048 ; 
      LAYER M3 ; 
        RECT 34.148 31.75 34.22 32.708 ; 
      LAYER V3 ; 
        RECT 34.148 31.952 34.22 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.568 34.66 31.664 ; 
      LAYER M3 ; 
        RECT 33.248 31.32 33.32 32.94 ; 
      LAYER V3 ; 
        RECT 33.248 31.568 33.32 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 36.272 34.388 36.368 ; 
      LAYER M3 ; 
        RECT 34.148 36.07 34.22 37.028 ; 
      LAYER V3 ; 
        RECT 34.148 36.272 34.22 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 35.888 34.66 35.984 ; 
      LAYER M3 ; 
        RECT 33.248 35.64 33.32 37.26 ; 
      LAYER V3 ; 
        RECT 33.248 35.888 33.32 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.592 34.388 40.688 ; 
      LAYER M3 ; 
        RECT 34.148 40.39 34.22 41.348 ; 
      LAYER V3 ; 
        RECT 34.148 40.592 34.22 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.208 34.66 40.304 ; 
      LAYER M3 ; 
        RECT 33.248 39.96 33.32 41.58 ; 
      LAYER V3 ; 
        RECT 33.248 40.208 33.32 40.304 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 44.912 34.388 45.008 ; 
      LAYER M3 ; 
        RECT 34.148 44.71 34.22 45.668 ; 
      LAYER V3 ; 
        RECT 34.148 44.912 34.22 45.008 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 44.528 34.66 44.624 ; 
      LAYER M3 ; 
        RECT 33.248 44.28 33.32 45.9 ; 
      LAYER V3 ; 
        RECT 33.248 44.528 33.32 44.624 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 49.232 34.388 49.328 ; 
      LAYER M3 ; 
        RECT 34.148 49.03 34.22 49.988 ; 
      LAYER V3 ; 
        RECT 34.148 49.232 34.22 49.328 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 48.848 34.66 48.944 ; 
      LAYER M3 ; 
        RECT 33.248 48.6 33.32 50.22 ; 
      LAYER V3 ; 
        RECT 33.248 48.848 33.32 48.944 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 53.552 34.388 53.648 ; 
      LAYER M3 ; 
        RECT 34.148 53.35 34.22 54.308 ; 
      LAYER V3 ; 
        RECT 34.148 53.552 34.22 53.648 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 53.168 34.66 53.264 ; 
      LAYER M3 ; 
        RECT 33.248 52.92 33.32 54.54 ; 
      LAYER V3 ; 
        RECT 33.248 53.168 33.32 53.264 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 57.872 34.388 57.968 ; 
      LAYER M3 ; 
        RECT 34.148 57.67 34.22 58.628 ; 
      LAYER V3 ; 
        RECT 34.148 57.872 34.22 57.968 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 57.488 34.66 57.584 ; 
      LAYER M3 ; 
        RECT 33.248 57.24 33.32 58.86 ; 
      LAYER V3 ; 
        RECT 33.248 57.488 33.32 57.584 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 62.192 34.388 62.288 ; 
      LAYER M3 ; 
        RECT 34.148 61.99 34.22 62.948 ; 
      LAYER V3 ; 
        RECT 34.148 62.192 34.22 62.288 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 61.808 34.66 61.904 ; 
      LAYER M3 ; 
        RECT 33.248 61.56 33.32 63.18 ; 
      LAYER V3 ; 
        RECT 33.248 61.808 33.32 61.904 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 66.512 34.388 66.608 ; 
      LAYER M3 ; 
        RECT 34.148 66.31 34.22 67.268 ; 
      LAYER V3 ; 
        RECT 34.148 66.512 34.22 66.608 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 66.128 34.66 66.224 ; 
      LAYER M3 ; 
        RECT 33.248 65.88 33.32 67.5 ; 
      LAYER V3 ; 
        RECT 33.248 66.128 33.32 66.224 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 70.832 34.388 70.928 ; 
      LAYER M3 ; 
        RECT 34.148 70.63 34.22 71.588 ; 
      LAYER V3 ; 
        RECT 34.148 70.832 34.22 70.928 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 70.448 34.66 70.544 ; 
      LAYER M3 ; 
        RECT 33.248 70.2 33.32 71.82 ; 
      LAYER V3 ; 
        RECT 33.248 70.448 33.32 70.544 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 107.66 34.388 107.756 ; 
      LAYER M3 ; 
        RECT 34.148 107.458 34.22 108.416 ; 
      LAYER V3 ; 
        RECT 34.148 107.66 34.22 107.756 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 107.276 34.66 107.372 ; 
      LAYER M3 ; 
        RECT 33.248 107.028 33.32 108.648 ; 
      LAYER V3 ; 
        RECT 33.248 107.276 33.32 107.372 ; 
    END 
  END wd[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 111.98 34.388 112.076 ; 
      LAYER M3 ; 
        RECT 34.148 111.778 34.22 112.736 ; 
      LAYER V3 ; 
        RECT 34.148 111.98 34.22 112.076 ; 
    END 
  END dataout[18] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 111.596 34.66 111.692 ; 
      LAYER M3 ; 
        RECT 33.248 111.348 33.32 112.968 ; 
      LAYER V3 ; 
        RECT 33.248 111.596 33.32 111.692 ; 
    END 
  END wd[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 116.3 34.388 116.396 ; 
      LAYER M3 ; 
        RECT 34.148 116.098 34.22 117.056 ; 
      LAYER V3 ; 
        RECT 34.148 116.3 34.22 116.396 ; 
    END 
  END dataout[19] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 115.916 34.66 116.012 ; 
      LAYER M3 ; 
        RECT 33.248 115.668 33.32 117.288 ; 
      LAYER V3 ; 
        RECT 33.248 115.916 33.32 116.012 ; 
    END 
  END wd[19] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 120.62 34.388 120.716 ; 
      LAYER M3 ; 
        RECT 34.148 120.418 34.22 121.376 ; 
      LAYER V3 ; 
        RECT 34.148 120.62 34.22 120.716 ; 
    END 
  END dataout[20] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 120.236 34.66 120.332 ; 
      LAYER M3 ; 
        RECT 33.248 119.988 33.32 121.608 ; 
      LAYER V3 ; 
        RECT 33.248 120.236 33.32 120.332 ; 
    END 
  END wd[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 124.94 34.388 125.036 ; 
      LAYER M3 ; 
        RECT 34.148 124.738 34.22 125.696 ; 
      LAYER V3 ; 
        RECT 34.148 124.94 34.22 125.036 ; 
    END 
  END dataout[21] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 124.556 34.66 124.652 ; 
      LAYER M3 ; 
        RECT 33.248 124.308 33.32 125.928 ; 
      LAYER V3 ; 
        RECT 33.248 124.556 33.32 124.652 ; 
    END 
  END wd[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 129.26 34.388 129.356 ; 
      LAYER M3 ; 
        RECT 34.148 129.058 34.22 130.016 ; 
      LAYER V3 ; 
        RECT 34.148 129.26 34.22 129.356 ; 
    END 
  END dataout[22] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 128.876 34.66 128.972 ; 
      LAYER M3 ; 
        RECT 33.248 128.628 33.32 130.248 ; 
      LAYER V3 ; 
        RECT 33.248 128.876 33.32 128.972 ; 
    END 
  END wd[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 133.58 34.388 133.676 ; 
      LAYER M3 ; 
        RECT 34.148 133.378 34.22 134.336 ; 
      LAYER V3 ; 
        RECT 34.148 133.58 34.22 133.676 ; 
    END 
  END dataout[23] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 133.196 34.66 133.292 ; 
      LAYER M3 ; 
        RECT 33.248 132.948 33.32 134.568 ; 
      LAYER V3 ; 
        RECT 33.248 133.196 33.32 133.292 ; 
    END 
  END wd[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 137.9 34.388 137.996 ; 
      LAYER M3 ; 
        RECT 34.148 137.698 34.22 138.656 ; 
      LAYER V3 ; 
        RECT 34.148 137.9 34.22 137.996 ; 
    END 
  END dataout[24] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 137.516 34.66 137.612 ; 
      LAYER M3 ; 
        RECT 33.248 137.268 33.32 138.888 ; 
      LAYER V3 ; 
        RECT 33.248 137.516 33.32 137.612 ; 
    END 
  END wd[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 142.22 34.388 142.316 ; 
      LAYER M3 ; 
        RECT 34.148 142.018 34.22 142.976 ; 
      LAYER V3 ; 
        RECT 34.148 142.22 34.22 142.316 ; 
    END 
  END dataout[25] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 141.836 34.66 141.932 ; 
      LAYER M3 ; 
        RECT 33.248 141.588 33.32 143.208 ; 
      LAYER V3 ; 
        RECT 33.248 141.836 33.32 141.932 ; 
    END 
  END wd[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 146.54 34.388 146.636 ; 
      LAYER M3 ; 
        RECT 34.148 146.338 34.22 147.296 ; 
      LAYER V3 ; 
        RECT 34.148 146.54 34.22 146.636 ; 
    END 
  END dataout[26] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 146.156 34.66 146.252 ; 
      LAYER M3 ; 
        RECT 33.248 145.908 33.32 147.528 ; 
      LAYER V3 ; 
        RECT 33.248 146.156 33.32 146.252 ; 
    END 
  END wd[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 150.86 34.388 150.956 ; 
      LAYER M3 ; 
        RECT 34.148 150.658 34.22 151.616 ; 
      LAYER V3 ; 
        RECT 34.148 150.86 34.22 150.956 ; 
    END 
  END dataout[27] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 150.476 34.66 150.572 ; 
      LAYER M3 ; 
        RECT 33.248 150.228 33.32 151.848 ; 
      LAYER V3 ; 
        RECT 33.248 150.476 33.32 150.572 ; 
    END 
  END wd[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 155.18 34.388 155.276 ; 
      LAYER M3 ; 
        RECT 34.148 154.978 34.22 155.936 ; 
      LAYER V3 ; 
        RECT 34.148 155.18 34.22 155.276 ; 
    END 
  END dataout[28] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 154.796 34.66 154.892 ; 
      LAYER M3 ; 
        RECT 33.248 154.548 33.32 156.168 ; 
      LAYER V3 ; 
        RECT 33.248 154.796 33.32 154.892 ; 
    END 
  END wd[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 159.5 34.388 159.596 ; 
      LAYER M3 ; 
        RECT 34.148 159.298 34.22 160.256 ; 
      LAYER V3 ; 
        RECT 34.148 159.5 34.22 159.596 ; 
    END 
  END dataout[29] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 159.116 34.66 159.212 ; 
      LAYER M3 ; 
        RECT 33.248 158.868 33.32 160.488 ; 
      LAYER V3 ; 
        RECT 33.248 159.116 33.32 159.212 ; 
    END 
  END wd[29] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 163.82 34.388 163.916 ; 
      LAYER M3 ; 
        RECT 34.148 163.618 34.22 164.576 ; 
      LAYER V3 ; 
        RECT 34.148 163.82 34.22 163.916 ; 
    END 
  END dataout[30] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 163.436 34.66 163.532 ; 
      LAYER M3 ; 
        RECT 33.248 163.188 33.32 164.808 ; 
      LAYER V3 ; 
        RECT 33.248 163.436 33.32 163.532 ; 
    END 
  END wd[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 168.14 34.388 168.236 ; 
      LAYER M3 ; 
        RECT 34.148 167.938 34.22 168.896 ; 
      LAYER V3 ; 
        RECT 34.148 168.14 34.22 168.236 ; 
    END 
  END dataout[31] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 167.756 34.66 167.852 ; 
      LAYER M3 ; 
        RECT 33.248 167.508 33.32 169.128 ; 
      LAYER V3 ; 
        RECT 33.248 167.756 33.32 167.852 ; 
    END 
  END wd[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 172.46 34.388 172.556 ; 
      LAYER M3 ; 
        RECT 34.148 172.258 34.22 173.216 ; 
      LAYER V3 ; 
        RECT 34.148 172.46 34.22 172.556 ; 
    END 
  END dataout[32] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 172.076 34.66 172.172 ; 
      LAYER M3 ; 
        RECT 33.248 171.828 33.32 173.448 ; 
      LAYER V3 ; 
        RECT 33.248 172.076 33.32 172.172 ; 
    END 
  END wd[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 176.78 34.388 176.876 ; 
      LAYER M3 ; 
        RECT 34.148 176.578 34.22 177.536 ; 
      LAYER V3 ; 
        RECT 34.148 176.78 34.22 176.876 ; 
    END 
  END dataout[33] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 176.396 34.66 176.492 ; 
      LAYER M3 ; 
        RECT 33.248 176.148 33.32 177.768 ; 
      LAYER V3 ; 
        RECT 33.248 176.396 33.32 176.492 ; 
    END 
  END wd[33] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0 74.388 66.096 109.002 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
        RECT 0.02 119.934 66.116 124.308 ; 
        RECT 0.02 124.254 66.116 128.628 ; 
        RECT 0.02 128.574 66.116 132.948 ; 
        RECT 0.02 132.894 66.116 137.268 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0 74.388 66.096 109.002 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
        RECT 0.02 119.934 66.116 124.308 ; 
        RECT 0.02 124.254 66.116 128.628 ; 
        RECT 0.02 128.574 66.116 132.948 ; 
        RECT 0.02 132.894 66.116 137.268 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
  LAYER V1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0 74.388 66.096 109.002 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
        RECT 0.02 119.934 66.116 124.308 ; 
        RECT 0.02 124.254 66.116 128.628 ; 
        RECT 0.02 128.574 66.116 132.948 ; 
        RECT 0.02 132.894 66.116 137.268 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
  LAYER V2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0 74.388 66.096 109.002 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
        RECT 0.02 119.934 66.116 124.308 ; 
        RECT 0.02 124.254 66.116 128.628 ; 
        RECT 0.02 128.574 66.116 132.948 ; 
        RECT 0.02 132.894 66.116 137.268 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
  LAYER M3 ; 
      RECT 34.796 1.38 34.868 5.122 ; 
      RECT 34.652 1.38 34.724 5.122 ; 
      RECT 34.508 3.688 34.58 4.978 ; 
      RECT 34.04 4.476 34.112 4.914 ; 
      RECT 34.004 1.51 34.076 2.468 ; 
      RECT 33.86 3.834 33.932 4.448 ; 
      RECT 33.536 3.936 33.608 4.968 ; 
      RECT 31.376 1.38 31.448 5.122 ; 
      RECT 31.232 1.38 31.304 5.122 ; 
      RECT 31.088 2.104 31.16 4.376 ; 
      RECT 34.796 5.7 34.868 9.442 ; 
      RECT 34.652 5.7 34.724 9.442 ; 
      RECT 34.508 8.008 34.58 9.298 ; 
      RECT 34.04 8.796 34.112 9.234 ; 
      RECT 34.004 5.83 34.076 6.788 ; 
      RECT 33.86 8.154 33.932 8.768 ; 
      RECT 33.536 8.256 33.608 9.288 ; 
      RECT 31.376 5.7 31.448 9.442 ; 
      RECT 31.232 5.7 31.304 9.442 ; 
      RECT 31.088 6.424 31.16 8.696 ; 
      RECT 34.796 10.02 34.868 13.762 ; 
      RECT 34.652 10.02 34.724 13.762 ; 
      RECT 34.508 12.328 34.58 13.618 ; 
      RECT 34.04 13.116 34.112 13.554 ; 
      RECT 34.004 10.15 34.076 11.108 ; 
      RECT 33.86 12.474 33.932 13.088 ; 
      RECT 33.536 12.576 33.608 13.608 ; 
      RECT 31.376 10.02 31.448 13.762 ; 
      RECT 31.232 10.02 31.304 13.762 ; 
      RECT 31.088 10.744 31.16 13.016 ; 
      RECT 34.796 14.34 34.868 18.082 ; 
      RECT 34.652 14.34 34.724 18.082 ; 
      RECT 34.508 16.648 34.58 17.938 ; 
      RECT 34.04 17.436 34.112 17.874 ; 
      RECT 34.004 14.47 34.076 15.428 ; 
      RECT 33.86 16.794 33.932 17.408 ; 
      RECT 33.536 16.896 33.608 17.928 ; 
      RECT 31.376 14.34 31.448 18.082 ; 
      RECT 31.232 14.34 31.304 18.082 ; 
      RECT 31.088 15.064 31.16 17.336 ; 
      RECT 34.796 18.66 34.868 22.402 ; 
      RECT 34.652 18.66 34.724 22.402 ; 
      RECT 34.508 20.968 34.58 22.258 ; 
      RECT 34.04 21.756 34.112 22.194 ; 
      RECT 34.004 18.79 34.076 19.748 ; 
      RECT 33.86 21.114 33.932 21.728 ; 
      RECT 33.536 21.216 33.608 22.248 ; 
      RECT 31.376 18.66 31.448 22.402 ; 
      RECT 31.232 18.66 31.304 22.402 ; 
      RECT 31.088 19.384 31.16 21.656 ; 
      RECT 34.796 22.98 34.868 26.722 ; 
      RECT 34.652 22.98 34.724 26.722 ; 
      RECT 34.508 25.288 34.58 26.578 ; 
      RECT 34.04 26.076 34.112 26.514 ; 
      RECT 34.004 23.11 34.076 24.068 ; 
      RECT 33.86 25.434 33.932 26.048 ; 
      RECT 33.536 25.536 33.608 26.568 ; 
      RECT 31.376 22.98 31.448 26.722 ; 
      RECT 31.232 22.98 31.304 26.722 ; 
      RECT 31.088 23.704 31.16 25.976 ; 
      RECT 34.796 27.3 34.868 31.042 ; 
      RECT 34.652 27.3 34.724 31.042 ; 
      RECT 34.508 29.608 34.58 30.898 ; 
      RECT 34.04 30.396 34.112 30.834 ; 
      RECT 34.004 27.43 34.076 28.388 ; 
      RECT 33.86 29.754 33.932 30.368 ; 
      RECT 33.536 29.856 33.608 30.888 ; 
      RECT 31.376 27.3 31.448 31.042 ; 
      RECT 31.232 27.3 31.304 31.042 ; 
      RECT 31.088 28.024 31.16 30.296 ; 
      RECT 34.796 31.62 34.868 35.362 ; 
      RECT 34.652 31.62 34.724 35.362 ; 
      RECT 34.508 33.928 34.58 35.218 ; 
      RECT 34.04 34.716 34.112 35.154 ; 
      RECT 34.004 31.75 34.076 32.708 ; 
      RECT 33.86 34.074 33.932 34.688 ; 
      RECT 33.536 34.176 33.608 35.208 ; 
      RECT 31.376 31.62 31.448 35.362 ; 
      RECT 31.232 31.62 31.304 35.362 ; 
      RECT 31.088 32.344 31.16 34.616 ; 
      RECT 34.796 35.94 34.868 39.682 ; 
      RECT 34.652 35.94 34.724 39.682 ; 
      RECT 34.508 38.248 34.58 39.538 ; 
      RECT 34.04 39.036 34.112 39.474 ; 
      RECT 34.004 36.07 34.076 37.028 ; 
      RECT 33.86 38.394 33.932 39.008 ; 
      RECT 33.536 38.496 33.608 39.528 ; 
      RECT 31.376 35.94 31.448 39.682 ; 
      RECT 31.232 35.94 31.304 39.682 ; 
      RECT 31.088 36.664 31.16 38.936 ; 
      RECT 34.796 40.26 34.868 44.002 ; 
      RECT 34.652 40.26 34.724 44.002 ; 
      RECT 34.508 42.568 34.58 43.858 ; 
      RECT 34.04 43.356 34.112 43.794 ; 
      RECT 34.004 40.39 34.076 41.348 ; 
      RECT 33.86 42.714 33.932 43.328 ; 
      RECT 33.536 42.816 33.608 43.848 ; 
      RECT 31.376 40.26 31.448 44.002 ; 
      RECT 31.232 40.26 31.304 44.002 ; 
      RECT 31.088 40.984 31.16 43.256 ; 
      RECT 34.796 44.58 34.868 48.322 ; 
      RECT 34.652 44.58 34.724 48.322 ; 
      RECT 34.508 46.888 34.58 48.178 ; 
      RECT 34.04 47.676 34.112 48.114 ; 
      RECT 34.004 44.71 34.076 45.668 ; 
      RECT 33.86 47.034 33.932 47.648 ; 
      RECT 33.536 47.136 33.608 48.168 ; 
      RECT 31.376 44.58 31.448 48.322 ; 
      RECT 31.232 44.58 31.304 48.322 ; 
      RECT 31.088 45.304 31.16 47.576 ; 
      RECT 34.796 48.9 34.868 52.642 ; 
      RECT 34.652 48.9 34.724 52.642 ; 
      RECT 34.508 51.208 34.58 52.498 ; 
      RECT 34.04 51.996 34.112 52.434 ; 
      RECT 34.004 49.03 34.076 49.988 ; 
      RECT 33.86 51.354 33.932 51.968 ; 
      RECT 33.536 51.456 33.608 52.488 ; 
      RECT 31.376 48.9 31.448 52.642 ; 
      RECT 31.232 48.9 31.304 52.642 ; 
      RECT 31.088 49.624 31.16 51.896 ; 
      RECT 34.796 53.22 34.868 56.962 ; 
      RECT 34.652 53.22 34.724 56.962 ; 
      RECT 34.508 55.528 34.58 56.818 ; 
      RECT 34.04 56.316 34.112 56.754 ; 
      RECT 34.004 53.35 34.076 54.308 ; 
      RECT 33.86 55.674 33.932 56.288 ; 
      RECT 33.536 55.776 33.608 56.808 ; 
      RECT 31.376 53.22 31.448 56.962 ; 
      RECT 31.232 53.22 31.304 56.962 ; 
      RECT 31.088 53.944 31.16 56.216 ; 
      RECT 34.796 57.54 34.868 61.282 ; 
      RECT 34.652 57.54 34.724 61.282 ; 
      RECT 34.508 59.848 34.58 61.138 ; 
      RECT 34.04 60.636 34.112 61.074 ; 
      RECT 34.004 57.67 34.076 58.628 ; 
      RECT 33.86 59.994 33.932 60.608 ; 
      RECT 33.536 60.096 33.608 61.128 ; 
      RECT 31.376 57.54 31.448 61.282 ; 
      RECT 31.232 57.54 31.304 61.282 ; 
      RECT 31.088 58.264 31.16 60.536 ; 
      RECT 34.796 61.86 34.868 65.602 ; 
      RECT 34.652 61.86 34.724 65.602 ; 
      RECT 34.508 64.168 34.58 65.458 ; 
      RECT 34.04 64.956 34.112 65.394 ; 
      RECT 34.004 61.99 34.076 62.948 ; 
      RECT 33.86 64.314 33.932 64.928 ; 
      RECT 33.536 64.416 33.608 65.448 ; 
      RECT 31.376 61.86 31.448 65.602 ; 
      RECT 31.232 61.86 31.304 65.602 ; 
      RECT 31.088 62.584 31.16 64.856 ; 
      RECT 34.796 66.18 34.868 69.922 ; 
      RECT 34.652 66.18 34.724 69.922 ; 
      RECT 34.508 68.488 34.58 69.778 ; 
      RECT 34.04 69.276 34.112 69.714 ; 
      RECT 34.004 66.31 34.076 67.268 ; 
      RECT 33.86 68.634 33.932 69.248 ; 
      RECT 33.536 68.736 33.608 69.768 ; 
      RECT 31.376 66.18 31.448 69.922 ; 
      RECT 31.232 66.18 31.304 69.922 ; 
      RECT 31.088 66.904 31.16 69.176 ; 
      RECT 34.796 70.5 34.868 74.242 ; 
      RECT 34.652 70.5 34.724 74.242 ; 
      RECT 34.508 72.808 34.58 74.098 ; 
      RECT 34.04 73.596 34.112 74.034 ; 
      RECT 34.004 70.63 34.076 71.588 ; 
      RECT 33.86 72.954 33.932 73.568 ; 
      RECT 33.536 73.056 33.608 74.088 ; 
      RECT 31.376 70.5 31.448 74.242 ; 
      RECT 31.232 70.5 31.304 74.242 ; 
      RECT 31.088 71.224 31.16 73.496 ; 
      RECT 65.268 89.56 65.34 106.976 ; 
      RECT 65.124 84.3 65.196 84.576 ; 
      RECT 65.124 90.78 65.196 91.112 ; 
      RECT 64.98 74.282 65.052 107.11 ; 
      RECT 64.836 89.69 64.908 92.45 ; 
      RECT 64.836 92.654 64.908 96.6 ; 
      RECT 64.836 96.76 64.908 99.228 ; 
      RECT 64.692 89.436 64.764 92.2548 ; 
      RECT 64.692 95.268 64.764 99.948 ; 
      RECT 64.548 74.282 64.62 88.668 ; 
      RECT 64.116 74.282 64.188 88.668 ; 
      RECT 63.684 74.282 63.756 88.668 ; 
      RECT 63.252 74.282 63.324 88.668 ; 
      RECT 62.82 74.282 62.892 88.668 ; 
      RECT 62.388 74.282 62.46 88.668 ; 
      RECT 61.956 74.282 62.028 88.668 ; 
      RECT 61.524 74.282 61.596 88.668 ; 
      RECT 61.092 74.282 61.164 88.668 ; 
      RECT 60.66 74.282 60.732 88.668 ; 
      RECT 60.228 74.282 60.3 88.668 ; 
      RECT 59.796 74.282 59.868 88.668 ; 
      RECT 59.364 74.282 59.436 88.668 ; 
      RECT 58.932 74.282 59.004 88.668 ; 
      RECT 58.5 74.282 58.572 88.668 ; 
      RECT 58.068 74.282 58.14 88.668 ; 
      RECT 57.636 74.282 57.708 88.668 ; 
      RECT 57.204 74.282 57.276 88.668 ; 
      RECT 56.772 74.282 56.844 88.668 ; 
      RECT 56.34 74.282 56.412 88.668 ; 
      RECT 55.908 74.282 55.98 88.668 ; 
      RECT 55.476 74.282 55.548 88.668 ; 
      RECT 55.044 74.282 55.116 88.668 ; 
      RECT 54.612 74.282 54.684 88.668 ; 
      RECT 54.18 74.282 54.252 88.668 ; 
      RECT 53.748 74.282 53.82 88.668 ; 
      RECT 53.316 74.282 53.388 88.668 ; 
      RECT 52.884 74.282 52.956 88.668 ; 
      RECT 52.452 74.282 52.524 88.668 ; 
      RECT 52.02 74.282 52.092 88.668 ; 
      RECT 51.588 74.282 51.66 88.668 ; 
      RECT 51.156 74.282 51.228 88.668 ; 
      RECT 50.724 74.282 50.796 88.668 ; 
      RECT 50.292 74.282 50.364 88.668 ; 
      RECT 49.86 74.282 49.932 88.668 ; 
      RECT 49.428 74.282 49.5 88.668 ; 
      RECT 48.996 74.282 49.068 88.668 ; 
      RECT 48.564 74.282 48.636 88.668 ; 
      RECT 48.132 74.282 48.204 88.668 ; 
      RECT 47.7 74.282 47.772 88.668 ; 
      RECT 47.268 74.282 47.34 88.668 ; 
      RECT 46.836 74.282 46.908 88.668 ; 
      RECT 46.404 74.282 46.476 88.668 ; 
      RECT 45.972 74.282 46.044 88.668 ; 
      RECT 45.54 74.282 45.612 88.668 ; 
      RECT 45.108 74.282 45.18 88.668 ; 
      RECT 44.676 74.282 44.748 88.668 ; 
      RECT 44.244 74.282 44.316 88.668 ; 
      RECT 43.812 74.282 43.884 88.668 ; 
      RECT 43.38 74.282 43.452 88.668 ; 
      RECT 42.948 74.282 43.02 88.668 ; 
      RECT 42.516 74.282 42.588 88.668 ; 
      RECT 42.084 74.282 42.156 88.668 ; 
      RECT 41.652 74.282 41.724 88.668 ; 
      RECT 41.22 74.282 41.292 88.668 ; 
      RECT 40.788 74.282 40.86 88.668 ; 
      RECT 40.356 74.282 40.428 88.668 ; 
      RECT 39.924 74.282 39.996 88.668 ; 
      RECT 39.492 74.282 39.564 88.668 ; 
      RECT 39.06 74.282 39.132 88.668 ; 
      RECT 38.628 74.282 38.7 88.668 ; 
      RECT 38.196 74.282 38.268 88.668 ; 
      RECT 38.052 89.702 38.124 92.27 ; 
      RECT 38.052 94.98 38.124 97.108 ; 
      RECT 37.98 76.924 38.052 79.628 ; 
      RECT 37.98 82.612 38.052 83.804 ; 
      RECT 37.98 87.076 38.052 88.124 ; 
      RECT 37.908 89.36 37.98 92.45 ; 
      RECT 37.908 92.6548 37.98 94.62 ; 
      RECT 37.908 94.8 37.98 96.284 ; 
      RECT 37.908 96.588 37.98 99.228 ; 
      RECT 37.764 74.282 37.836 107.11 ; 
      RECT 37.62 91.532 37.692 93.39 ; 
      RECT 37.548 77.356 37.62 79.88 ; 
      RECT 37.548 81.532 37.62 82.292 ; 
      RECT 37.548 85.06 37.62 85.256 ; 
      RECT 37.548 87.988 37.62 88.136 ; 
      RECT 37.476 89.56 37.548 106.958 ; 
      RECT 37.116 75.844 37.188 79.052 ; 
      RECT 37.116 81.244 37.188 83.516 ; 
      RECT 36.972 81.532 37.044 83.012 ; 
      RECT 36.828 78.94 36.9 79.484 ; 
      RECT 36.828 82.9 36.9 83.804 ; 
      RECT 36.828 87.868 36.9 88.124 ; 
      RECT 36.684 79.348 36.756 79.496 ; 
      RECT 36.684 85.852 36.756 86.024 ; 
      RECT 36.684 87.988 36.756 88.136 ; 
      RECT 36.54 80.596 36.612 82.58 ; 
      RECT 36.54 82.756 36.612 83.516 ; 
      RECT 36.54 86.596 36.612 87.836 ; 
      RECT 36.396 80.164 36.468 85.152 ; 
      RECT 36.396 95.716 36.468 98.636 ; 
      RECT 36.396 100.036 36.468 102.956 ; 
      RECT 35.1 79.084 35.172 80.276 ; 
      RECT 35.1 83.836 35.172 84.092 ; 
      RECT 35.1 84.916 35.172 86.756 ; 
      RECT 35.1 89.716 35.172 89.864 ; 
      RECT 35.1 97.876 35.172 99.068 ; 
      RECT 34.956 79.372 35.028 81.392 ; 
      RECT 34.956 82.468 35.028 85.676 ; 
      RECT 34.956 89.848 35.028 90.932 ; 
      RECT 34.956 91.252 35.028 92.156 ; 
      RECT 34.812 79.084 34.884 81.788 ; 
      RECT 34.812 82.18 34.884 83.516 ; 
      RECT 34.812 84.34 34.884 84.884 ; 
      RECT 34.812 87.076 34.884 90.284 ; 
      RECT 34.812 92.02 34.884 92.168 ; 
      RECT 34.812 100.684 34.884 102.02 ; 
      RECT 34.668 80.02 34.74 80.564 ; 
      RECT 34.668 87.58 34.74 91.508 ; 
      RECT 34.668 93.268 34.74 94.46 ; 
      RECT 34.668 100.036 34.74 101.084 ; 
      RECT 34.524 76.276 34.596 76.892 ; 
      RECT 34.524 79.516 34.596 86.66 ; 
      RECT 34.524 90.82 34.596 100.148 ; 
      RECT 34.524 100.972 34.596 105.404 ; 
      RECT 33.372 77.356 33.444 78.404 ; 
      RECT 33.372 78.94 33.444 79.196 ; 
      RECT 33.372 79.516 33.444 80.42 ; 
      RECT 33.372 80.596 33.444 81.356 ; 
      RECT 33.372 81.676 33.444 92.156 ; 
      RECT 33.372 92.332 33.444 97.556 ; 
      RECT 33.372 101.908 33.444 102.956 ; 
      RECT 33.228 81.352 33.3 82.436 ; 
      RECT 33.228 82.756 33.3 86.108 ; 
      RECT 33.228 86.788 33.3 90.14 ; 
      RECT 33.228 90.316 33.3 95.396 ; 
      RECT 33.228 96.22 33.3 96.908 ; 
      RECT 33.228 99.748 33.3 104.036 ; 
      RECT 33.084 81.676 33.156 82.76 ; 
      RECT 33.084 83.38 33.156 83.528 ; 
      RECT 33.084 86.5 33.156 90.428 ; 
      RECT 33.084 91.396 33.156 93.236 ; 
      RECT 33.084 94.636 33.156 97.592 ; 
      RECT 32.94 78.148 33.012 82.436 ; 
      RECT 32.94 88.804 33.012 89.672 ; 
      RECT 32.94 94.348 33.012 95.54 ; 
      RECT 32.796 80.74 32.868 82.58 ; 
      RECT 32.796 87.076 32.868 87.836 ; 
      RECT 32.796 88 32.868 88.148 ; 
      RECT 32.796 89.092 32.868 90.428 ; 
      RECT 32.796 90.964 32.868 96.332 ; 
      RECT 32.796 96.76 32.868 101.228 ; 
      RECT 32.652 78.436 32.724 79.196 ; 
      RECT 32.652 80.02 32.724 80.564 ; 
      RECT 32.652 81.676 32.724 94.316 ; 
      RECT 32.652 94.636 32.724 96.476 ; 
      RECT 32.652 98.956 32.724 100.796 ; 
      RECT 32.652 104.212 32.724 105.116 ; 
      RECT 32.508 74.388 32.58 75.004 ; 
      RECT 32.508 106.368 32.58 107.032 ; 
      RECT 32.364 74.388 32.436 74.588 ; 
      RECT 32.076 74.388 32.148 74.674 ; 
      RECT 32.076 106.646 32.148 107.11 ; 
      RECT 31.5 80.452 31.572 81.212 ; 
      RECT 31.5 83.404 31.572 84.884 ; 
      RECT 31.5 91.252 31.572 92.156 ; 
      RECT 31.5 93.412 31.572 97.988 ; 
      RECT 31.5 101.116 31.572 102.956 ; 
      RECT 31.5 105.268 31.572 105.416 ; 
      RECT 31.356 76.276 31.428 78.26 ; 
      RECT 31.356 92.596 31.428 92.744 ; 
      RECT 31.356 96.904 31.428 100.148 ; 
      RECT 31.212 78.148 31.284 79.196 ; 
      RECT 31.212 80.308 31.284 81.644 ; 
      RECT 31.212 82.468 31.284 82.868 ; 
      RECT 31.212 85.996 31.284 97.052 ; 
      RECT 31.212 97.588 31.284 98.492 ; 
      RECT 31.068 76.78 31.14 81.356 ; 
      RECT 31.068 95.716 31.14 96.476 ; 
      RECT 31.068 98.932 31.14 99.08 ; 
      RECT 31.068 100.036 31.14 103.244 ; 
      RECT 30.924 80.596 30.996 84.596 ; 
      RECT 30.924 98.356 30.996 98.504 ; 
      RECT 29.484 78.94 29.556 80.564 ; 
      RECT 29.196 79.084 29.268 81.5 ; 
      RECT 29.052 78.436 29.124 78.692 ; 
      RECT 28.908 74.6 28.98 74.804 ; 
      RECT 28.908 87.076 28.98 87.836 ; 
      RECT 28.836 89.56 28.908 106.954 ; 
      RECT 28.548 89.56 28.62 106.958 ; 
      RECT 28.476 76.276 28.548 77.036 ; 
      RECT 28.476 79.372 28.548 88.412 ; 
      RECT 28.404 91.532 28.476 93.39 ; 
      RECT 28.26 74.282 28.332 107.11 ; 
      RECT 28.116 89.36 28.188 92.45 ; 
      RECT 28.116 92.6548 28.188 94.62 ; 
      RECT 28.116 94.8 28.188 96.284 ; 
      RECT 28.116 96.588 28.188 99.228 ; 
      RECT 28.044 76.276 28.116 78.26 ; 
      RECT 28.044 81.388 28.116 83.66 ; 
      RECT 28.044 84.916 28.116 87.836 ; 
      RECT 27.972 89.702 28.044 92.27 ; 
      RECT 27.972 94.98 28.044 97.108 ; 
      RECT 27.828 74.282 27.9 88.668 ; 
      RECT 27.396 74.282 27.468 88.668 ; 
      RECT 26.964 74.282 27.036 88.668 ; 
      RECT 26.532 74.282 26.604 88.668 ; 
      RECT 26.1 74.282 26.172 88.668 ; 
      RECT 25.668 74.282 25.74 88.668 ; 
      RECT 25.236 74.282 25.308 88.668 ; 
      RECT 24.804 74.282 24.876 88.668 ; 
      RECT 24.372 74.282 24.444 88.668 ; 
      RECT 23.94 74.282 24.012 88.668 ; 
      RECT 23.508 74.282 23.58 88.668 ; 
      RECT 23.076 74.282 23.148 88.668 ; 
      RECT 22.644 74.282 22.716 88.668 ; 
      RECT 22.212 74.282 22.284 88.668 ; 
      RECT 21.78 74.282 21.852 88.668 ; 
      RECT 21.348 74.282 21.42 88.668 ; 
      RECT 20.916 74.282 20.988 88.668 ; 
      RECT 20.484 74.282 20.556 88.668 ; 
      RECT 20.052 74.282 20.124 88.668 ; 
      RECT 19.62 74.282 19.692 88.668 ; 
      RECT 19.188 74.282 19.26 88.668 ; 
      RECT 18.756 74.282 18.828 88.668 ; 
      RECT 18.324 74.282 18.396 88.668 ; 
      RECT 17.892 74.282 17.964 88.668 ; 
      RECT 17.46 74.282 17.532 88.668 ; 
      RECT 17.028 74.282 17.1 88.668 ; 
      RECT 16.596 74.282 16.668 88.668 ; 
      RECT 16.164 74.282 16.236 88.668 ; 
      RECT 15.732 74.282 15.804 88.668 ; 
      RECT 15.3 74.282 15.372 88.668 ; 
      RECT 14.868 74.282 14.94 88.668 ; 
      RECT 14.436 74.282 14.508 88.668 ; 
      RECT 14.004 74.282 14.076 88.668 ; 
      RECT 13.572 74.282 13.644 88.668 ; 
      RECT 13.14 74.282 13.212 88.668 ; 
      RECT 12.708 74.282 12.78 88.668 ; 
      RECT 12.276 74.282 12.348 88.668 ; 
      RECT 11.844 74.282 11.916 88.668 ; 
      RECT 11.412 74.282 11.484 88.668 ; 
      RECT 10.98 74.282 11.052 88.668 ; 
      RECT 10.548 74.282 10.62 88.668 ; 
      RECT 10.116 74.282 10.188 88.668 ; 
      RECT 9.684 74.282 9.756 88.668 ; 
      RECT 9.252 74.282 9.324 88.668 ; 
      RECT 8.82 74.282 8.892 88.668 ; 
      RECT 8.388 74.282 8.46 88.668 ; 
      RECT 7.956 74.282 8.028 88.668 ; 
      RECT 7.524 74.282 7.596 88.668 ; 
      RECT 7.092 74.282 7.164 88.668 ; 
      RECT 6.66 74.282 6.732 88.668 ; 
      RECT 6.228 74.282 6.3 88.668 ; 
      RECT 5.796 74.282 5.868 88.668 ; 
      RECT 5.364 74.282 5.436 88.668 ; 
      RECT 4.932 74.282 5.004 88.668 ; 
      RECT 4.5 74.282 4.572 88.668 ; 
      RECT 4.068 74.282 4.14 88.668 ; 
      RECT 3.636 74.282 3.708 88.668 ; 
      RECT 3.204 74.282 3.276 88.668 ; 
      RECT 2.772 74.282 2.844 88.668 ; 
      RECT 2.34 74.282 2.412 88.668 ; 
      RECT 1.908 74.282 1.98 88.668 ; 
      RECT 1.476 74.282 1.548 88.668 ; 
      RECT 1.332 89.436 1.404 92.2548 ; 
      RECT 1.332 95.268 1.404 99.948 ; 
      RECT 1.188 89.69 1.26 92.45 ; 
      RECT 1.188 92.654 1.26 96.6 ; 
      RECT 1.188 96.76 1.26 99.228 ; 
      RECT 1.044 74.282 1.116 107.11 ; 
      RECT 0.9 84.3 0.972 84.576 ; 
      RECT 0.9 90.78 0.972 91.112 ; 
      RECT 0.756 89.56 0.828 106.976 ; 
        RECT 34.796 107.328 34.868 111.07 ; 
        RECT 34.652 107.328 34.724 111.07 ; 
        RECT 34.508 109.636 34.58 110.926 ; 
        RECT 34.04 110.424 34.112 110.862 ; 
        RECT 34.004 107.458 34.076 108.416 ; 
        RECT 33.86 109.782 33.932 110.396 ; 
        RECT 33.536 109.884 33.608 110.916 ; 
        RECT 31.376 107.328 31.448 111.07 ; 
        RECT 31.232 107.328 31.304 111.07 ; 
        RECT 31.088 108.052 31.16 110.324 ; 
        RECT 34.796 111.648 34.868 115.39 ; 
        RECT 34.652 111.648 34.724 115.39 ; 
        RECT 34.508 113.956 34.58 115.246 ; 
        RECT 34.04 114.744 34.112 115.182 ; 
        RECT 34.004 111.778 34.076 112.736 ; 
        RECT 33.86 114.102 33.932 114.716 ; 
        RECT 33.536 114.204 33.608 115.236 ; 
        RECT 31.376 111.648 31.448 115.39 ; 
        RECT 31.232 111.648 31.304 115.39 ; 
        RECT 31.088 112.372 31.16 114.644 ; 
        RECT 34.796 115.968 34.868 119.71 ; 
        RECT 34.652 115.968 34.724 119.71 ; 
        RECT 34.508 118.276 34.58 119.566 ; 
        RECT 34.04 119.064 34.112 119.502 ; 
        RECT 34.004 116.098 34.076 117.056 ; 
        RECT 33.86 118.422 33.932 119.036 ; 
        RECT 33.536 118.524 33.608 119.556 ; 
        RECT 31.376 115.968 31.448 119.71 ; 
        RECT 31.232 115.968 31.304 119.71 ; 
        RECT 31.088 116.692 31.16 118.964 ; 
        RECT 34.796 120.288 34.868 124.03 ; 
        RECT 34.652 120.288 34.724 124.03 ; 
        RECT 34.508 122.596 34.58 123.886 ; 
        RECT 34.04 123.384 34.112 123.822 ; 
        RECT 34.004 120.418 34.076 121.376 ; 
        RECT 33.86 122.742 33.932 123.356 ; 
        RECT 33.536 122.844 33.608 123.876 ; 
        RECT 31.376 120.288 31.448 124.03 ; 
        RECT 31.232 120.288 31.304 124.03 ; 
        RECT 31.088 121.012 31.16 123.284 ; 
        RECT 34.796 124.608 34.868 128.35 ; 
        RECT 34.652 124.608 34.724 128.35 ; 
        RECT 34.508 126.916 34.58 128.206 ; 
        RECT 34.04 127.704 34.112 128.142 ; 
        RECT 34.004 124.738 34.076 125.696 ; 
        RECT 33.86 127.062 33.932 127.676 ; 
        RECT 33.536 127.164 33.608 128.196 ; 
        RECT 31.376 124.608 31.448 128.35 ; 
        RECT 31.232 124.608 31.304 128.35 ; 
        RECT 31.088 125.332 31.16 127.604 ; 
        RECT 34.796 128.928 34.868 132.67 ; 
        RECT 34.652 128.928 34.724 132.67 ; 
        RECT 34.508 131.236 34.58 132.526 ; 
        RECT 34.04 132.024 34.112 132.462 ; 
        RECT 34.004 129.058 34.076 130.016 ; 
        RECT 33.86 131.382 33.932 131.996 ; 
        RECT 33.536 131.484 33.608 132.516 ; 
        RECT 31.376 128.928 31.448 132.67 ; 
        RECT 31.232 128.928 31.304 132.67 ; 
        RECT 31.088 129.652 31.16 131.924 ; 
        RECT 34.796 133.248 34.868 136.99 ; 
        RECT 34.652 133.248 34.724 136.99 ; 
        RECT 34.508 135.556 34.58 136.846 ; 
        RECT 34.04 136.344 34.112 136.782 ; 
        RECT 34.004 133.378 34.076 134.336 ; 
        RECT 33.86 135.702 33.932 136.316 ; 
        RECT 33.536 135.804 33.608 136.836 ; 
        RECT 31.376 133.248 31.448 136.99 ; 
        RECT 31.232 133.248 31.304 136.99 ; 
        RECT 31.088 133.972 31.16 136.244 ; 
        RECT 34.796 137.568 34.868 141.31 ; 
        RECT 34.652 137.568 34.724 141.31 ; 
        RECT 34.508 139.876 34.58 141.166 ; 
        RECT 34.04 140.664 34.112 141.102 ; 
        RECT 34.004 137.698 34.076 138.656 ; 
        RECT 33.86 140.022 33.932 140.636 ; 
        RECT 33.536 140.124 33.608 141.156 ; 
        RECT 31.376 137.568 31.448 141.31 ; 
        RECT 31.232 137.568 31.304 141.31 ; 
        RECT 31.088 138.292 31.16 140.564 ; 
        RECT 34.796 141.888 34.868 145.63 ; 
        RECT 34.652 141.888 34.724 145.63 ; 
        RECT 34.508 144.196 34.58 145.486 ; 
        RECT 34.04 144.984 34.112 145.422 ; 
        RECT 34.004 142.018 34.076 142.976 ; 
        RECT 33.86 144.342 33.932 144.956 ; 
        RECT 33.536 144.444 33.608 145.476 ; 
        RECT 31.376 141.888 31.448 145.63 ; 
        RECT 31.232 141.888 31.304 145.63 ; 
        RECT 31.088 142.612 31.16 144.884 ; 
        RECT 34.796 146.208 34.868 149.95 ; 
        RECT 34.652 146.208 34.724 149.95 ; 
        RECT 34.508 148.516 34.58 149.806 ; 
        RECT 34.04 149.304 34.112 149.742 ; 
        RECT 34.004 146.338 34.076 147.296 ; 
        RECT 33.86 148.662 33.932 149.276 ; 
        RECT 33.536 148.764 33.608 149.796 ; 
        RECT 31.376 146.208 31.448 149.95 ; 
        RECT 31.232 146.208 31.304 149.95 ; 
        RECT 31.088 146.932 31.16 149.204 ; 
        RECT 34.796 150.528 34.868 154.27 ; 
        RECT 34.652 150.528 34.724 154.27 ; 
        RECT 34.508 152.836 34.58 154.126 ; 
        RECT 34.04 153.624 34.112 154.062 ; 
        RECT 34.004 150.658 34.076 151.616 ; 
        RECT 33.86 152.982 33.932 153.596 ; 
        RECT 33.536 153.084 33.608 154.116 ; 
        RECT 31.376 150.528 31.448 154.27 ; 
        RECT 31.232 150.528 31.304 154.27 ; 
        RECT 31.088 151.252 31.16 153.524 ; 
        RECT 34.796 154.848 34.868 158.59 ; 
        RECT 34.652 154.848 34.724 158.59 ; 
        RECT 34.508 157.156 34.58 158.446 ; 
        RECT 34.04 157.944 34.112 158.382 ; 
        RECT 34.004 154.978 34.076 155.936 ; 
        RECT 33.86 157.302 33.932 157.916 ; 
        RECT 33.536 157.404 33.608 158.436 ; 
        RECT 31.376 154.848 31.448 158.59 ; 
        RECT 31.232 154.848 31.304 158.59 ; 
        RECT 31.088 155.572 31.16 157.844 ; 
        RECT 34.796 159.168 34.868 162.91 ; 
        RECT 34.652 159.168 34.724 162.91 ; 
        RECT 34.508 161.476 34.58 162.766 ; 
        RECT 34.04 162.264 34.112 162.702 ; 
        RECT 34.004 159.298 34.076 160.256 ; 
        RECT 33.86 161.622 33.932 162.236 ; 
        RECT 33.536 161.724 33.608 162.756 ; 
        RECT 31.376 159.168 31.448 162.91 ; 
        RECT 31.232 159.168 31.304 162.91 ; 
        RECT 31.088 159.892 31.16 162.164 ; 
        RECT 34.796 163.488 34.868 167.23 ; 
        RECT 34.652 163.488 34.724 167.23 ; 
        RECT 34.508 165.796 34.58 167.086 ; 
        RECT 34.04 166.584 34.112 167.022 ; 
        RECT 34.004 163.618 34.076 164.576 ; 
        RECT 33.86 165.942 33.932 166.556 ; 
        RECT 33.536 166.044 33.608 167.076 ; 
        RECT 31.376 163.488 31.448 167.23 ; 
        RECT 31.232 163.488 31.304 167.23 ; 
        RECT 31.088 164.212 31.16 166.484 ; 
        RECT 34.796 167.808 34.868 171.55 ; 
        RECT 34.652 167.808 34.724 171.55 ; 
        RECT 34.508 170.116 34.58 171.406 ; 
        RECT 34.04 170.904 34.112 171.342 ; 
        RECT 34.004 167.938 34.076 168.896 ; 
        RECT 33.86 170.262 33.932 170.876 ; 
        RECT 33.536 170.364 33.608 171.396 ; 
        RECT 31.376 167.808 31.448 171.55 ; 
        RECT 31.232 167.808 31.304 171.55 ; 
        RECT 31.088 168.532 31.16 170.804 ; 
        RECT 34.796 172.128 34.868 175.87 ; 
        RECT 34.652 172.128 34.724 175.87 ; 
        RECT 34.508 174.436 34.58 175.726 ; 
        RECT 34.04 175.224 34.112 175.662 ; 
        RECT 34.004 172.258 34.076 173.216 ; 
        RECT 33.86 174.582 33.932 175.196 ; 
        RECT 33.536 174.684 33.608 175.716 ; 
        RECT 31.376 172.128 31.448 175.87 ; 
        RECT 31.232 172.128 31.304 175.87 ; 
        RECT 31.088 172.852 31.16 175.124 ; 
        RECT 34.796 176.448 34.868 180.19 ; 
        RECT 34.652 176.448 34.724 180.19 ; 
        RECT 34.508 178.756 34.58 180.046 ; 
        RECT 34.04 179.544 34.112 179.982 ; 
        RECT 34.004 176.578 34.076 177.536 ; 
        RECT 33.86 178.902 33.932 179.516 ; 
        RECT 33.536 179.004 33.608 180.036 ; 
        RECT 31.376 176.448 31.448 180.19 ; 
        RECT 31.232 176.448 31.304 180.19 ; 
        RECT 31.088 177.172 31.16 179.444 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 34.564 1.026 35.076 5.4 ; 
      RECT 34.508 3.688 35.076 4.978 ; 
      RECT 33.916 2.596 34.164 5.4 ; 
      RECT 33.86 3.834 34.164 4.448 ; 
      RECT 33.916 1.026 34.02 5.4 ; 
      RECT 33.916 1.51 34.076 2.468 ; 
      RECT 33.916 1.026 34.164 1.382 ; 
      RECT 32.728 2.828 33.552 5.4 ; 
      RECT 33.448 1.026 33.552 5.4 ; 
      RECT 32.728 3.936 33.608 4.968 ; 
      RECT 32.728 1.026 33.12 5.4 ; 
      RECT 31.06 1.026 31.392 5.4 ; 
      RECT 31.06 1.38 31.448 5.122 ; 
      RECT 65.776 1.026 66.116 5.4 ; 
      RECT 65.2 1.026 65.304 5.4 ; 
      RECT 64.768 1.026 64.872 5.4 ; 
      RECT 64.336 1.026 64.44 5.4 ; 
      RECT 63.904 1.026 64.008 5.4 ; 
      RECT 63.472 1.026 63.576 5.4 ; 
      RECT 63.04 1.026 63.144 5.4 ; 
      RECT 62.608 1.026 62.712 5.4 ; 
      RECT 62.176 1.026 62.28 5.4 ; 
      RECT 61.744 1.026 61.848 5.4 ; 
      RECT 61.312 1.026 61.416 5.4 ; 
      RECT 60.88 1.026 60.984 5.4 ; 
      RECT 60.448 1.026 60.552 5.4 ; 
      RECT 60.016 1.026 60.12 5.4 ; 
      RECT 59.584 1.026 59.688 5.4 ; 
      RECT 59.152 1.026 59.256 5.4 ; 
      RECT 58.72 1.026 58.824 5.4 ; 
      RECT 58.288 1.026 58.392 5.4 ; 
      RECT 57.856 1.026 57.96 5.4 ; 
      RECT 57.424 1.026 57.528 5.4 ; 
      RECT 56.992 1.026 57.096 5.4 ; 
      RECT 56.56 1.026 56.664 5.4 ; 
      RECT 56.128 1.026 56.232 5.4 ; 
      RECT 55.696 1.026 55.8 5.4 ; 
      RECT 55.264 1.026 55.368 5.4 ; 
      RECT 54.832 1.026 54.936 5.4 ; 
      RECT 54.4 1.026 54.504 5.4 ; 
      RECT 53.968 1.026 54.072 5.4 ; 
      RECT 53.536 1.026 53.64 5.4 ; 
      RECT 53.104 1.026 53.208 5.4 ; 
      RECT 52.672 1.026 52.776 5.4 ; 
      RECT 52.24 1.026 52.344 5.4 ; 
      RECT 51.808 1.026 51.912 5.4 ; 
      RECT 51.376 1.026 51.48 5.4 ; 
      RECT 50.944 1.026 51.048 5.4 ; 
      RECT 50.512 1.026 50.616 5.4 ; 
      RECT 50.08 1.026 50.184 5.4 ; 
      RECT 49.648 1.026 49.752 5.4 ; 
      RECT 49.216 1.026 49.32 5.4 ; 
      RECT 48.784 1.026 48.888 5.4 ; 
      RECT 48.352 1.026 48.456 5.4 ; 
      RECT 47.92 1.026 48.024 5.4 ; 
      RECT 47.488 1.026 47.592 5.4 ; 
      RECT 47.056 1.026 47.16 5.4 ; 
      RECT 46.624 1.026 46.728 5.4 ; 
      RECT 46.192 1.026 46.296 5.4 ; 
      RECT 45.76 1.026 45.864 5.4 ; 
      RECT 45.328 1.026 45.432 5.4 ; 
      RECT 44.896 1.026 45 5.4 ; 
      RECT 44.464 1.026 44.568 5.4 ; 
      RECT 44.032 1.026 44.136 5.4 ; 
      RECT 43.6 1.026 43.704 5.4 ; 
      RECT 43.168 1.026 43.272 5.4 ; 
      RECT 42.736 1.026 42.84 5.4 ; 
      RECT 42.304 1.026 42.408 5.4 ; 
      RECT 41.872 1.026 41.976 5.4 ; 
      RECT 41.44 1.026 41.544 5.4 ; 
      RECT 41.008 1.026 41.112 5.4 ; 
      RECT 40.576 1.026 40.68 5.4 ; 
      RECT 40.144 1.026 40.248 5.4 ; 
      RECT 39.712 1.026 39.816 5.4 ; 
      RECT 39.28 1.026 39.384 5.4 ; 
      RECT 38.848 1.026 38.952 5.4 ; 
      RECT 38.416 1.026 38.52 5.4 ; 
      RECT 37.984 1.026 38.088 5.4 ; 
      RECT 37.552 1.026 37.656 5.4 ; 
      RECT 36.7 1.026 37.008 5.4 ; 
      RECT 29.128 1.026 29.436 5.4 ; 
      RECT 28.48 1.026 28.584 5.4 ; 
      RECT 28.048 1.026 28.152 5.4 ; 
      RECT 27.616 1.026 27.72 5.4 ; 
      RECT 27.184 1.026 27.288 5.4 ; 
      RECT 26.752 1.026 26.856 5.4 ; 
      RECT 26.32 1.026 26.424 5.4 ; 
      RECT 25.888 1.026 25.992 5.4 ; 
      RECT 25.456 1.026 25.56 5.4 ; 
      RECT 25.024 1.026 25.128 5.4 ; 
      RECT 24.592 1.026 24.696 5.4 ; 
      RECT 24.16 1.026 24.264 5.4 ; 
      RECT 23.728 1.026 23.832 5.4 ; 
      RECT 23.296 1.026 23.4 5.4 ; 
      RECT 22.864 1.026 22.968 5.4 ; 
      RECT 22.432 1.026 22.536 5.4 ; 
      RECT 22 1.026 22.104 5.4 ; 
      RECT 21.568 1.026 21.672 5.4 ; 
      RECT 21.136 1.026 21.24 5.4 ; 
      RECT 20.704 1.026 20.808 5.4 ; 
      RECT 20.272 1.026 20.376 5.4 ; 
      RECT 19.84 1.026 19.944 5.4 ; 
      RECT 19.408 1.026 19.512 5.4 ; 
      RECT 18.976 1.026 19.08 5.4 ; 
      RECT 18.544 1.026 18.648 5.4 ; 
      RECT 18.112 1.026 18.216 5.4 ; 
      RECT 17.68 1.026 17.784 5.4 ; 
      RECT 17.248 1.026 17.352 5.4 ; 
      RECT 16.816 1.026 16.92 5.4 ; 
      RECT 16.384 1.026 16.488 5.4 ; 
      RECT 15.952 1.026 16.056 5.4 ; 
      RECT 15.52 1.026 15.624 5.4 ; 
      RECT 15.088 1.026 15.192 5.4 ; 
      RECT 14.656 1.026 14.76 5.4 ; 
      RECT 14.224 1.026 14.328 5.4 ; 
      RECT 13.792 1.026 13.896 5.4 ; 
      RECT 13.36 1.026 13.464 5.4 ; 
      RECT 12.928 1.026 13.032 5.4 ; 
      RECT 12.496 1.026 12.6 5.4 ; 
      RECT 12.064 1.026 12.168 5.4 ; 
      RECT 11.632 1.026 11.736 5.4 ; 
      RECT 11.2 1.026 11.304 5.4 ; 
      RECT 10.768 1.026 10.872 5.4 ; 
      RECT 10.336 1.026 10.44 5.4 ; 
      RECT 9.904 1.026 10.008 5.4 ; 
      RECT 9.472 1.026 9.576 5.4 ; 
      RECT 9.04 1.026 9.144 5.4 ; 
      RECT 8.608 1.026 8.712 5.4 ; 
      RECT 8.176 1.026 8.28 5.4 ; 
      RECT 7.744 1.026 7.848 5.4 ; 
      RECT 7.312 1.026 7.416 5.4 ; 
      RECT 6.88 1.026 6.984 5.4 ; 
      RECT 6.448 1.026 6.552 5.4 ; 
      RECT 6.016 1.026 6.12 5.4 ; 
      RECT 5.584 1.026 5.688 5.4 ; 
      RECT 5.152 1.026 5.256 5.4 ; 
      RECT 4.72 1.026 4.824 5.4 ; 
      RECT 4.288 1.026 4.392 5.4 ; 
      RECT 3.856 1.026 3.96 5.4 ; 
      RECT 3.424 1.026 3.528 5.4 ; 
      RECT 2.992 1.026 3.096 5.4 ; 
      RECT 2.56 1.026 2.664 5.4 ; 
      RECT 2.128 1.026 2.232 5.4 ; 
      RECT 1.696 1.026 1.8 5.4 ; 
      RECT 1.264 1.026 1.368 5.4 ; 
      RECT 0.832 1.026 0.936 5.4 ; 
      RECT 0.02 1.026 0.36 5.4 ; 
      RECT 34.564 5.346 35.076 9.72 ; 
      RECT 34.508 8.008 35.076 9.298 ; 
      RECT 33.916 6.916 34.164 9.72 ; 
      RECT 33.86 8.154 34.164 8.768 ; 
      RECT 33.916 5.346 34.02 9.72 ; 
      RECT 33.916 5.83 34.076 6.788 ; 
      RECT 33.916 5.346 34.164 5.702 ; 
      RECT 32.728 7.148 33.552 9.72 ; 
      RECT 33.448 5.346 33.552 9.72 ; 
      RECT 32.728 8.256 33.608 9.288 ; 
      RECT 32.728 5.346 33.12 9.72 ; 
      RECT 31.06 5.346 31.392 9.72 ; 
      RECT 31.06 5.7 31.448 9.442 ; 
      RECT 65.776 5.346 66.116 9.72 ; 
      RECT 65.2 5.346 65.304 9.72 ; 
      RECT 64.768 5.346 64.872 9.72 ; 
      RECT 64.336 5.346 64.44 9.72 ; 
      RECT 63.904 5.346 64.008 9.72 ; 
      RECT 63.472 5.346 63.576 9.72 ; 
      RECT 63.04 5.346 63.144 9.72 ; 
      RECT 62.608 5.346 62.712 9.72 ; 
      RECT 62.176 5.346 62.28 9.72 ; 
      RECT 61.744 5.346 61.848 9.72 ; 
      RECT 61.312 5.346 61.416 9.72 ; 
      RECT 60.88 5.346 60.984 9.72 ; 
      RECT 60.448 5.346 60.552 9.72 ; 
      RECT 60.016 5.346 60.12 9.72 ; 
      RECT 59.584 5.346 59.688 9.72 ; 
      RECT 59.152 5.346 59.256 9.72 ; 
      RECT 58.72 5.346 58.824 9.72 ; 
      RECT 58.288 5.346 58.392 9.72 ; 
      RECT 57.856 5.346 57.96 9.72 ; 
      RECT 57.424 5.346 57.528 9.72 ; 
      RECT 56.992 5.346 57.096 9.72 ; 
      RECT 56.56 5.346 56.664 9.72 ; 
      RECT 56.128 5.346 56.232 9.72 ; 
      RECT 55.696 5.346 55.8 9.72 ; 
      RECT 55.264 5.346 55.368 9.72 ; 
      RECT 54.832 5.346 54.936 9.72 ; 
      RECT 54.4 5.346 54.504 9.72 ; 
      RECT 53.968 5.346 54.072 9.72 ; 
      RECT 53.536 5.346 53.64 9.72 ; 
      RECT 53.104 5.346 53.208 9.72 ; 
      RECT 52.672 5.346 52.776 9.72 ; 
      RECT 52.24 5.346 52.344 9.72 ; 
      RECT 51.808 5.346 51.912 9.72 ; 
      RECT 51.376 5.346 51.48 9.72 ; 
      RECT 50.944 5.346 51.048 9.72 ; 
      RECT 50.512 5.346 50.616 9.72 ; 
      RECT 50.08 5.346 50.184 9.72 ; 
      RECT 49.648 5.346 49.752 9.72 ; 
      RECT 49.216 5.346 49.32 9.72 ; 
      RECT 48.784 5.346 48.888 9.72 ; 
      RECT 48.352 5.346 48.456 9.72 ; 
      RECT 47.92 5.346 48.024 9.72 ; 
      RECT 47.488 5.346 47.592 9.72 ; 
      RECT 47.056 5.346 47.16 9.72 ; 
      RECT 46.624 5.346 46.728 9.72 ; 
      RECT 46.192 5.346 46.296 9.72 ; 
      RECT 45.76 5.346 45.864 9.72 ; 
      RECT 45.328 5.346 45.432 9.72 ; 
      RECT 44.896 5.346 45 9.72 ; 
      RECT 44.464 5.346 44.568 9.72 ; 
      RECT 44.032 5.346 44.136 9.72 ; 
      RECT 43.6 5.346 43.704 9.72 ; 
      RECT 43.168 5.346 43.272 9.72 ; 
      RECT 42.736 5.346 42.84 9.72 ; 
      RECT 42.304 5.346 42.408 9.72 ; 
      RECT 41.872 5.346 41.976 9.72 ; 
      RECT 41.44 5.346 41.544 9.72 ; 
      RECT 41.008 5.346 41.112 9.72 ; 
      RECT 40.576 5.346 40.68 9.72 ; 
      RECT 40.144 5.346 40.248 9.72 ; 
      RECT 39.712 5.346 39.816 9.72 ; 
      RECT 39.28 5.346 39.384 9.72 ; 
      RECT 38.848 5.346 38.952 9.72 ; 
      RECT 38.416 5.346 38.52 9.72 ; 
      RECT 37.984 5.346 38.088 9.72 ; 
      RECT 37.552 5.346 37.656 9.72 ; 
      RECT 36.7 5.346 37.008 9.72 ; 
      RECT 29.128 5.346 29.436 9.72 ; 
      RECT 28.48 5.346 28.584 9.72 ; 
      RECT 28.048 5.346 28.152 9.72 ; 
      RECT 27.616 5.346 27.72 9.72 ; 
      RECT 27.184 5.346 27.288 9.72 ; 
      RECT 26.752 5.346 26.856 9.72 ; 
      RECT 26.32 5.346 26.424 9.72 ; 
      RECT 25.888 5.346 25.992 9.72 ; 
      RECT 25.456 5.346 25.56 9.72 ; 
      RECT 25.024 5.346 25.128 9.72 ; 
      RECT 24.592 5.346 24.696 9.72 ; 
      RECT 24.16 5.346 24.264 9.72 ; 
      RECT 23.728 5.346 23.832 9.72 ; 
      RECT 23.296 5.346 23.4 9.72 ; 
      RECT 22.864 5.346 22.968 9.72 ; 
      RECT 22.432 5.346 22.536 9.72 ; 
      RECT 22 5.346 22.104 9.72 ; 
      RECT 21.568 5.346 21.672 9.72 ; 
      RECT 21.136 5.346 21.24 9.72 ; 
      RECT 20.704 5.346 20.808 9.72 ; 
      RECT 20.272 5.346 20.376 9.72 ; 
      RECT 19.84 5.346 19.944 9.72 ; 
      RECT 19.408 5.346 19.512 9.72 ; 
      RECT 18.976 5.346 19.08 9.72 ; 
      RECT 18.544 5.346 18.648 9.72 ; 
      RECT 18.112 5.346 18.216 9.72 ; 
      RECT 17.68 5.346 17.784 9.72 ; 
      RECT 17.248 5.346 17.352 9.72 ; 
      RECT 16.816 5.346 16.92 9.72 ; 
      RECT 16.384 5.346 16.488 9.72 ; 
      RECT 15.952 5.346 16.056 9.72 ; 
      RECT 15.52 5.346 15.624 9.72 ; 
      RECT 15.088 5.346 15.192 9.72 ; 
      RECT 14.656 5.346 14.76 9.72 ; 
      RECT 14.224 5.346 14.328 9.72 ; 
      RECT 13.792 5.346 13.896 9.72 ; 
      RECT 13.36 5.346 13.464 9.72 ; 
      RECT 12.928 5.346 13.032 9.72 ; 
      RECT 12.496 5.346 12.6 9.72 ; 
      RECT 12.064 5.346 12.168 9.72 ; 
      RECT 11.632 5.346 11.736 9.72 ; 
      RECT 11.2 5.346 11.304 9.72 ; 
      RECT 10.768 5.346 10.872 9.72 ; 
      RECT 10.336 5.346 10.44 9.72 ; 
      RECT 9.904 5.346 10.008 9.72 ; 
      RECT 9.472 5.346 9.576 9.72 ; 
      RECT 9.04 5.346 9.144 9.72 ; 
      RECT 8.608 5.346 8.712 9.72 ; 
      RECT 8.176 5.346 8.28 9.72 ; 
      RECT 7.744 5.346 7.848 9.72 ; 
      RECT 7.312 5.346 7.416 9.72 ; 
      RECT 6.88 5.346 6.984 9.72 ; 
      RECT 6.448 5.346 6.552 9.72 ; 
      RECT 6.016 5.346 6.12 9.72 ; 
      RECT 5.584 5.346 5.688 9.72 ; 
      RECT 5.152 5.346 5.256 9.72 ; 
      RECT 4.72 5.346 4.824 9.72 ; 
      RECT 4.288 5.346 4.392 9.72 ; 
      RECT 3.856 5.346 3.96 9.72 ; 
      RECT 3.424 5.346 3.528 9.72 ; 
      RECT 2.992 5.346 3.096 9.72 ; 
      RECT 2.56 5.346 2.664 9.72 ; 
      RECT 2.128 5.346 2.232 9.72 ; 
      RECT 1.696 5.346 1.8 9.72 ; 
      RECT 1.264 5.346 1.368 9.72 ; 
      RECT 0.832 5.346 0.936 9.72 ; 
      RECT 0.02 5.346 0.36 9.72 ; 
      RECT 34.564 9.666 35.076 14.04 ; 
      RECT 34.508 12.328 35.076 13.618 ; 
      RECT 33.916 11.236 34.164 14.04 ; 
      RECT 33.86 12.474 34.164 13.088 ; 
      RECT 33.916 9.666 34.02 14.04 ; 
      RECT 33.916 10.15 34.076 11.108 ; 
      RECT 33.916 9.666 34.164 10.022 ; 
      RECT 32.728 11.468 33.552 14.04 ; 
      RECT 33.448 9.666 33.552 14.04 ; 
      RECT 32.728 12.576 33.608 13.608 ; 
      RECT 32.728 9.666 33.12 14.04 ; 
      RECT 31.06 9.666 31.392 14.04 ; 
      RECT 31.06 10.02 31.448 13.762 ; 
      RECT 65.776 9.666 66.116 14.04 ; 
      RECT 65.2 9.666 65.304 14.04 ; 
      RECT 64.768 9.666 64.872 14.04 ; 
      RECT 64.336 9.666 64.44 14.04 ; 
      RECT 63.904 9.666 64.008 14.04 ; 
      RECT 63.472 9.666 63.576 14.04 ; 
      RECT 63.04 9.666 63.144 14.04 ; 
      RECT 62.608 9.666 62.712 14.04 ; 
      RECT 62.176 9.666 62.28 14.04 ; 
      RECT 61.744 9.666 61.848 14.04 ; 
      RECT 61.312 9.666 61.416 14.04 ; 
      RECT 60.88 9.666 60.984 14.04 ; 
      RECT 60.448 9.666 60.552 14.04 ; 
      RECT 60.016 9.666 60.12 14.04 ; 
      RECT 59.584 9.666 59.688 14.04 ; 
      RECT 59.152 9.666 59.256 14.04 ; 
      RECT 58.72 9.666 58.824 14.04 ; 
      RECT 58.288 9.666 58.392 14.04 ; 
      RECT 57.856 9.666 57.96 14.04 ; 
      RECT 57.424 9.666 57.528 14.04 ; 
      RECT 56.992 9.666 57.096 14.04 ; 
      RECT 56.56 9.666 56.664 14.04 ; 
      RECT 56.128 9.666 56.232 14.04 ; 
      RECT 55.696 9.666 55.8 14.04 ; 
      RECT 55.264 9.666 55.368 14.04 ; 
      RECT 54.832 9.666 54.936 14.04 ; 
      RECT 54.4 9.666 54.504 14.04 ; 
      RECT 53.968 9.666 54.072 14.04 ; 
      RECT 53.536 9.666 53.64 14.04 ; 
      RECT 53.104 9.666 53.208 14.04 ; 
      RECT 52.672 9.666 52.776 14.04 ; 
      RECT 52.24 9.666 52.344 14.04 ; 
      RECT 51.808 9.666 51.912 14.04 ; 
      RECT 51.376 9.666 51.48 14.04 ; 
      RECT 50.944 9.666 51.048 14.04 ; 
      RECT 50.512 9.666 50.616 14.04 ; 
      RECT 50.08 9.666 50.184 14.04 ; 
      RECT 49.648 9.666 49.752 14.04 ; 
      RECT 49.216 9.666 49.32 14.04 ; 
      RECT 48.784 9.666 48.888 14.04 ; 
      RECT 48.352 9.666 48.456 14.04 ; 
      RECT 47.92 9.666 48.024 14.04 ; 
      RECT 47.488 9.666 47.592 14.04 ; 
      RECT 47.056 9.666 47.16 14.04 ; 
      RECT 46.624 9.666 46.728 14.04 ; 
      RECT 46.192 9.666 46.296 14.04 ; 
      RECT 45.76 9.666 45.864 14.04 ; 
      RECT 45.328 9.666 45.432 14.04 ; 
      RECT 44.896 9.666 45 14.04 ; 
      RECT 44.464 9.666 44.568 14.04 ; 
      RECT 44.032 9.666 44.136 14.04 ; 
      RECT 43.6 9.666 43.704 14.04 ; 
      RECT 43.168 9.666 43.272 14.04 ; 
      RECT 42.736 9.666 42.84 14.04 ; 
      RECT 42.304 9.666 42.408 14.04 ; 
      RECT 41.872 9.666 41.976 14.04 ; 
      RECT 41.44 9.666 41.544 14.04 ; 
      RECT 41.008 9.666 41.112 14.04 ; 
      RECT 40.576 9.666 40.68 14.04 ; 
      RECT 40.144 9.666 40.248 14.04 ; 
      RECT 39.712 9.666 39.816 14.04 ; 
      RECT 39.28 9.666 39.384 14.04 ; 
      RECT 38.848 9.666 38.952 14.04 ; 
      RECT 38.416 9.666 38.52 14.04 ; 
      RECT 37.984 9.666 38.088 14.04 ; 
      RECT 37.552 9.666 37.656 14.04 ; 
      RECT 36.7 9.666 37.008 14.04 ; 
      RECT 29.128 9.666 29.436 14.04 ; 
      RECT 28.48 9.666 28.584 14.04 ; 
      RECT 28.048 9.666 28.152 14.04 ; 
      RECT 27.616 9.666 27.72 14.04 ; 
      RECT 27.184 9.666 27.288 14.04 ; 
      RECT 26.752 9.666 26.856 14.04 ; 
      RECT 26.32 9.666 26.424 14.04 ; 
      RECT 25.888 9.666 25.992 14.04 ; 
      RECT 25.456 9.666 25.56 14.04 ; 
      RECT 25.024 9.666 25.128 14.04 ; 
      RECT 24.592 9.666 24.696 14.04 ; 
      RECT 24.16 9.666 24.264 14.04 ; 
      RECT 23.728 9.666 23.832 14.04 ; 
      RECT 23.296 9.666 23.4 14.04 ; 
      RECT 22.864 9.666 22.968 14.04 ; 
      RECT 22.432 9.666 22.536 14.04 ; 
      RECT 22 9.666 22.104 14.04 ; 
      RECT 21.568 9.666 21.672 14.04 ; 
      RECT 21.136 9.666 21.24 14.04 ; 
      RECT 20.704 9.666 20.808 14.04 ; 
      RECT 20.272 9.666 20.376 14.04 ; 
      RECT 19.84 9.666 19.944 14.04 ; 
      RECT 19.408 9.666 19.512 14.04 ; 
      RECT 18.976 9.666 19.08 14.04 ; 
      RECT 18.544 9.666 18.648 14.04 ; 
      RECT 18.112 9.666 18.216 14.04 ; 
      RECT 17.68 9.666 17.784 14.04 ; 
      RECT 17.248 9.666 17.352 14.04 ; 
      RECT 16.816 9.666 16.92 14.04 ; 
      RECT 16.384 9.666 16.488 14.04 ; 
      RECT 15.952 9.666 16.056 14.04 ; 
      RECT 15.52 9.666 15.624 14.04 ; 
      RECT 15.088 9.666 15.192 14.04 ; 
      RECT 14.656 9.666 14.76 14.04 ; 
      RECT 14.224 9.666 14.328 14.04 ; 
      RECT 13.792 9.666 13.896 14.04 ; 
      RECT 13.36 9.666 13.464 14.04 ; 
      RECT 12.928 9.666 13.032 14.04 ; 
      RECT 12.496 9.666 12.6 14.04 ; 
      RECT 12.064 9.666 12.168 14.04 ; 
      RECT 11.632 9.666 11.736 14.04 ; 
      RECT 11.2 9.666 11.304 14.04 ; 
      RECT 10.768 9.666 10.872 14.04 ; 
      RECT 10.336 9.666 10.44 14.04 ; 
      RECT 9.904 9.666 10.008 14.04 ; 
      RECT 9.472 9.666 9.576 14.04 ; 
      RECT 9.04 9.666 9.144 14.04 ; 
      RECT 8.608 9.666 8.712 14.04 ; 
      RECT 8.176 9.666 8.28 14.04 ; 
      RECT 7.744 9.666 7.848 14.04 ; 
      RECT 7.312 9.666 7.416 14.04 ; 
      RECT 6.88 9.666 6.984 14.04 ; 
      RECT 6.448 9.666 6.552 14.04 ; 
      RECT 6.016 9.666 6.12 14.04 ; 
      RECT 5.584 9.666 5.688 14.04 ; 
      RECT 5.152 9.666 5.256 14.04 ; 
      RECT 4.72 9.666 4.824 14.04 ; 
      RECT 4.288 9.666 4.392 14.04 ; 
      RECT 3.856 9.666 3.96 14.04 ; 
      RECT 3.424 9.666 3.528 14.04 ; 
      RECT 2.992 9.666 3.096 14.04 ; 
      RECT 2.56 9.666 2.664 14.04 ; 
      RECT 2.128 9.666 2.232 14.04 ; 
      RECT 1.696 9.666 1.8 14.04 ; 
      RECT 1.264 9.666 1.368 14.04 ; 
      RECT 0.832 9.666 0.936 14.04 ; 
      RECT 0.02 9.666 0.36 14.04 ; 
      RECT 34.564 13.986 35.076 18.36 ; 
      RECT 34.508 16.648 35.076 17.938 ; 
      RECT 33.916 15.556 34.164 18.36 ; 
      RECT 33.86 16.794 34.164 17.408 ; 
      RECT 33.916 13.986 34.02 18.36 ; 
      RECT 33.916 14.47 34.076 15.428 ; 
      RECT 33.916 13.986 34.164 14.342 ; 
      RECT 32.728 15.788 33.552 18.36 ; 
      RECT 33.448 13.986 33.552 18.36 ; 
      RECT 32.728 16.896 33.608 17.928 ; 
      RECT 32.728 13.986 33.12 18.36 ; 
      RECT 31.06 13.986 31.392 18.36 ; 
      RECT 31.06 14.34 31.448 18.082 ; 
      RECT 65.776 13.986 66.116 18.36 ; 
      RECT 65.2 13.986 65.304 18.36 ; 
      RECT 64.768 13.986 64.872 18.36 ; 
      RECT 64.336 13.986 64.44 18.36 ; 
      RECT 63.904 13.986 64.008 18.36 ; 
      RECT 63.472 13.986 63.576 18.36 ; 
      RECT 63.04 13.986 63.144 18.36 ; 
      RECT 62.608 13.986 62.712 18.36 ; 
      RECT 62.176 13.986 62.28 18.36 ; 
      RECT 61.744 13.986 61.848 18.36 ; 
      RECT 61.312 13.986 61.416 18.36 ; 
      RECT 60.88 13.986 60.984 18.36 ; 
      RECT 60.448 13.986 60.552 18.36 ; 
      RECT 60.016 13.986 60.12 18.36 ; 
      RECT 59.584 13.986 59.688 18.36 ; 
      RECT 59.152 13.986 59.256 18.36 ; 
      RECT 58.72 13.986 58.824 18.36 ; 
      RECT 58.288 13.986 58.392 18.36 ; 
      RECT 57.856 13.986 57.96 18.36 ; 
      RECT 57.424 13.986 57.528 18.36 ; 
      RECT 56.992 13.986 57.096 18.36 ; 
      RECT 56.56 13.986 56.664 18.36 ; 
      RECT 56.128 13.986 56.232 18.36 ; 
      RECT 55.696 13.986 55.8 18.36 ; 
      RECT 55.264 13.986 55.368 18.36 ; 
      RECT 54.832 13.986 54.936 18.36 ; 
      RECT 54.4 13.986 54.504 18.36 ; 
      RECT 53.968 13.986 54.072 18.36 ; 
      RECT 53.536 13.986 53.64 18.36 ; 
      RECT 53.104 13.986 53.208 18.36 ; 
      RECT 52.672 13.986 52.776 18.36 ; 
      RECT 52.24 13.986 52.344 18.36 ; 
      RECT 51.808 13.986 51.912 18.36 ; 
      RECT 51.376 13.986 51.48 18.36 ; 
      RECT 50.944 13.986 51.048 18.36 ; 
      RECT 50.512 13.986 50.616 18.36 ; 
      RECT 50.08 13.986 50.184 18.36 ; 
      RECT 49.648 13.986 49.752 18.36 ; 
      RECT 49.216 13.986 49.32 18.36 ; 
      RECT 48.784 13.986 48.888 18.36 ; 
      RECT 48.352 13.986 48.456 18.36 ; 
      RECT 47.92 13.986 48.024 18.36 ; 
      RECT 47.488 13.986 47.592 18.36 ; 
      RECT 47.056 13.986 47.16 18.36 ; 
      RECT 46.624 13.986 46.728 18.36 ; 
      RECT 46.192 13.986 46.296 18.36 ; 
      RECT 45.76 13.986 45.864 18.36 ; 
      RECT 45.328 13.986 45.432 18.36 ; 
      RECT 44.896 13.986 45 18.36 ; 
      RECT 44.464 13.986 44.568 18.36 ; 
      RECT 44.032 13.986 44.136 18.36 ; 
      RECT 43.6 13.986 43.704 18.36 ; 
      RECT 43.168 13.986 43.272 18.36 ; 
      RECT 42.736 13.986 42.84 18.36 ; 
      RECT 42.304 13.986 42.408 18.36 ; 
      RECT 41.872 13.986 41.976 18.36 ; 
      RECT 41.44 13.986 41.544 18.36 ; 
      RECT 41.008 13.986 41.112 18.36 ; 
      RECT 40.576 13.986 40.68 18.36 ; 
      RECT 40.144 13.986 40.248 18.36 ; 
      RECT 39.712 13.986 39.816 18.36 ; 
      RECT 39.28 13.986 39.384 18.36 ; 
      RECT 38.848 13.986 38.952 18.36 ; 
      RECT 38.416 13.986 38.52 18.36 ; 
      RECT 37.984 13.986 38.088 18.36 ; 
      RECT 37.552 13.986 37.656 18.36 ; 
      RECT 36.7 13.986 37.008 18.36 ; 
      RECT 29.128 13.986 29.436 18.36 ; 
      RECT 28.48 13.986 28.584 18.36 ; 
      RECT 28.048 13.986 28.152 18.36 ; 
      RECT 27.616 13.986 27.72 18.36 ; 
      RECT 27.184 13.986 27.288 18.36 ; 
      RECT 26.752 13.986 26.856 18.36 ; 
      RECT 26.32 13.986 26.424 18.36 ; 
      RECT 25.888 13.986 25.992 18.36 ; 
      RECT 25.456 13.986 25.56 18.36 ; 
      RECT 25.024 13.986 25.128 18.36 ; 
      RECT 24.592 13.986 24.696 18.36 ; 
      RECT 24.16 13.986 24.264 18.36 ; 
      RECT 23.728 13.986 23.832 18.36 ; 
      RECT 23.296 13.986 23.4 18.36 ; 
      RECT 22.864 13.986 22.968 18.36 ; 
      RECT 22.432 13.986 22.536 18.36 ; 
      RECT 22 13.986 22.104 18.36 ; 
      RECT 21.568 13.986 21.672 18.36 ; 
      RECT 21.136 13.986 21.24 18.36 ; 
      RECT 20.704 13.986 20.808 18.36 ; 
      RECT 20.272 13.986 20.376 18.36 ; 
      RECT 19.84 13.986 19.944 18.36 ; 
      RECT 19.408 13.986 19.512 18.36 ; 
      RECT 18.976 13.986 19.08 18.36 ; 
      RECT 18.544 13.986 18.648 18.36 ; 
      RECT 18.112 13.986 18.216 18.36 ; 
      RECT 17.68 13.986 17.784 18.36 ; 
      RECT 17.248 13.986 17.352 18.36 ; 
      RECT 16.816 13.986 16.92 18.36 ; 
      RECT 16.384 13.986 16.488 18.36 ; 
      RECT 15.952 13.986 16.056 18.36 ; 
      RECT 15.52 13.986 15.624 18.36 ; 
      RECT 15.088 13.986 15.192 18.36 ; 
      RECT 14.656 13.986 14.76 18.36 ; 
      RECT 14.224 13.986 14.328 18.36 ; 
      RECT 13.792 13.986 13.896 18.36 ; 
      RECT 13.36 13.986 13.464 18.36 ; 
      RECT 12.928 13.986 13.032 18.36 ; 
      RECT 12.496 13.986 12.6 18.36 ; 
      RECT 12.064 13.986 12.168 18.36 ; 
      RECT 11.632 13.986 11.736 18.36 ; 
      RECT 11.2 13.986 11.304 18.36 ; 
      RECT 10.768 13.986 10.872 18.36 ; 
      RECT 10.336 13.986 10.44 18.36 ; 
      RECT 9.904 13.986 10.008 18.36 ; 
      RECT 9.472 13.986 9.576 18.36 ; 
      RECT 9.04 13.986 9.144 18.36 ; 
      RECT 8.608 13.986 8.712 18.36 ; 
      RECT 8.176 13.986 8.28 18.36 ; 
      RECT 7.744 13.986 7.848 18.36 ; 
      RECT 7.312 13.986 7.416 18.36 ; 
      RECT 6.88 13.986 6.984 18.36 ; 
      RECT 6.448 13.986 6.552 18.36 ; 
      RECT 6.016 13.986 6.12 18.36 ; 
      RECT 5.584 13.986 5.688 18.36 ; 
      RECT 5.152 13.986 5.256 18.36 ; 
      RECT 4.72 13.986 4.824 18.36 ; 
      RECT 4.288 13.986 4.392 18.36 ; 
      RECT 3.856 13.986 3.96 18.36 ; 
      RECT 3.424 13.986 3.528 18.36 ; 
      RECT 2.992 13.986 3.096 18.36 ; 
      RECT 2.56 13.986 2.664 18.36 ; 
      RECT 2.128 13.986 2.232 18.36 ; 
      RECT 1.696 13.986 1.8 18.36 ; 
      RECT 1.264 13.986 1.368 18.36 ; 
      RECT 0.832 13.986 0.936 18.36 ; 
      RECT 0.02 13.986 0.36 18.36 ; 
      RECT 34.564 18.306 35.076 22.68 ; 
      RECT 34.508 20.968 35.076 22.258 ; 
      RECT 33.916 19.876 34.164 22.68 ; 
      RECT 33.86 21.114 34.164 21.728 ; 
      RECT 33.916 18.306 34.02 22.68 ; 
      RECT 33.916 18.79 34.076 19.748 ; 
      RECT 33.916 18.306 34.164 18.662 ; 
      RECT 32.728 20.108 33.552 22.68 ; 
      RECT 33.448 18.306 33.552 22.68 ; 
      RECT 32.728 21.216 33.608 22.248 ; 
      RECT 32.728 18.306 33.12 22.68 ; 
      RECT 31.06 18.306 31.392 22.68 ; 
      RECT 31.06 18.66 31.448 22.402 ; 
      RECT 65.776 18.306 66.116 22.68 ; 
      RECT 65.2 18.306 65.304 22.68 ; 
      RECT 64.768 18.306 64.872 22.68 ; 
      RECT 64.336 18.306 64.44 22.68 ; 
      RECT 63.904 18.306 64.008 22.68 ; 
      RECT 63.472 18.306 63.576 22.68 ; 
      RECT 63.04 18.306 63.144 22.68 ; 
      RECT 62.608 18.306 62.712 22.68 ; 
      RECT 62.176 18.306 62.28 22.68 ; 
      RECT 61.744 18.306 61.848 22.68 ; 
      RECT 61.312 18.306 61.416 22.68 ; 
      RECT 60.88 18.306 60.984 22.68 ; 
      RECT 60.448 18.306 60.552 22.68 ; 
      RECT 60.016 18.306 60.12 22.68 ; 
      RECT 59.584 18.306 59.688 22.68 ; 
      RECT 59.152 18.306 59.256 22.68 ; 
      RECT 58.72 18.306 58.824 22.68 ; 
      RECT 58.288 18.306 58.392 22.68 ; 
      RECT 57.856 18.306 57.96 22.68 ; 
      RECT 57.424 18.306 57.528 22.68 ; 
      RECT 56.992 18.306 57.096 22.68 ; 
      RECT 56.56 18.306 56.664 22.68 ; 
      RECT 56.128 18.306 56.232 22.68 ; 
      RECT 55.696 18.306 55.8 22.68 ; 
      RECT 55.264 18.306 55.368 22.68 ; 
      RECT 54.832 18.306 54.936 22.68 ; 
      RECT 54.4 18.306 54.504 22.68 ; 
      RECT 53.968 18.306 54.072 22.68 ; 
      RECT 53.536 18.306 53.64 22.68 ; 
      RECT 53.104 18.306 53.208 22.68 ; 
      RECT 52.672 18.306 52.776 22.68 ; 
      RECT 52.24 18.306 52.344 22.68 ; 
      RECT 51.808 18.306 51.912 22.68 ; 
      RECT 51.376 18.306 51.48 22.68 ; 
      RECT 50.944 18.306 51.048 22.68 ; 
      RECT 50.512 18.306 50.616 22.68 ; 
      RECT 50.08 18.306 50.184 22.68 ; 
      RECT 49.648 18.306 49.752 22.68 ; 
      RECT 49.216 18.306 49.32 22.68 ; 
      RECT 48.784 18.306 48.888 22.68 ; 
      RECT 48.352 18.306 48.456 22.68 ; 
      RECT 47.92 18.306 48.024 22.68 ; 
      RECT 47.488 18.306 47.592 22.68 ; 
      RECT 47.056 18.306 47.16 22.68 ; 
      RECT 46.624 18.306 46.728 22.68 ; 
      RECT 46.192 18.306 46.296 22.68 ; 
      RECT 45.76 18.306 45.864 22.68 ; 
      RECT 45.328 18.306 45.432 22.68 ; 
      RECT 44.896 18.306 45 22.68 ; 
      RECT 44.464 18.306 44.568 22.68 ; 
      RECT 44.032 18.306 44.136 22.68 ; 
      RECT 43.6 18.306 43.704 22.68 ; 
      RECT 43.168 18.306 43.272 22.68 ; 
      RECT 42.736 18.306 42.84 22.68 ; 
      RECT 42.304 18.306 42.408 22.68 ; 
      RECT 41.872 18.306 41.976 22.68 ; 
      RECT 41.44 18.306 41.544 22.68 ; 
      RECT 41.008 18.306 41.112 22.68 ; 
      RECT 40.576 18.306 40.68 22.68 ; 
      RECT 40.144 18.306 40.248 22.68 ; 
      RECT 39.712 18.306 39.816 22.68 ; 
      RECT 39.28 18.306 39.384 22.68 ; 
      RECT 38.848 18.306 38.952 22.68 ; 
      RECT 38.416 18.306 38.52 22.68 ; 
      RECT 37.984 18.306 38.088 22.68 ; 
      RECT 37.552 18.306 37.656 22.68 ; 
      RECT 36.7 18.306 37.008 22.68 ; 
      RECT 29.128 18.306 29.436 22.68 ; 
      RECT 28.48 18.306 28.584 22.68 ; 
      RECT 28.048 18.306 28.152 22.68 ; 
      RECT 27.616 18.306 27.72 22.68 ; 
      RECT 27.184 18.306 27.288 22.68 ; 
      RECT 26.752 18.306 26.856 22.68 ; 
      RECT 26.32 18.306 26.424 22.68 ; 
      RECT 25.888 18.306 25.992 22.68 ; 
      RECT 25.456 18.306 25.56 22.68 ; 
      RECT 25.024 18.306 25.128 22.68 ; 
      RECT 24.592 18.306 24.696 22.68 ; 
      RECT 24.16 18.306 24.264 22.68 ; 
      RECT 23.728 18.306 23.832 22.68 ; 
      RECT 23.296 18.306 23.4 22.68 ; 
      RECT 22.864 18.306 22.968 22.68 ; 
      RECT 22.432 18.306 22.536 22.68 ; 
      RECT 22 18.306 22.104 22.68 ; 
      RECT 21.568 18.306 21.672 22.68 ; 
      RECT 21.136 18.306 21.24 22.68 ; 
      RECT 20.704 18.306 20.808 22.68 ; 
      RECT 20.272 18.306 20.376 22.68 ; 
      RECT 19.84 18.306 19.944 22.68 ; 
      RECT 19.408 18.306 19.512 22.68 ; 
      RECT 18.976 18.306 19.08 22.68 ; 
      RECT 18.544 18.306 18.648 22.68 ; 
      RECT 18.112 18.306 18.216 22.68 ; 
      RECT 17.68 18.306 17.784 22.68 ; 
      RECT 17.248 18.306 17.352 22.68 ; 
      RECT 16.816 18.306 16.92 22.68 ; 
      RECT 16.384 18.306 16.488 22.68 ; 
      RECT 15.952 18.306 16.056 22.68 ; 
      RECT 15.52 18.306 15.624 22.68 ; 
      RECT 15.088 18.306 15.192 22.68 ; 
      RECT 14.656 18.306 14.76 22.68 ; 
      RECT 14.224 18.306 14.328 22.68 ; 
      RECT 13.792 18.306 13.896 22.68 ; 
      RECT 13.36 18.306 13.464 22.68 ; 
      RECT 12.928 18.306 13.032 22.68 ; 
      RECT 12.496 18.306 12.6 22.68 ; 
      RECT 12.064 18.306 12.168 22.68 ; 
      RECT 11.632 18.306 11.736 22.68 ; 
      RECT 11.2 18.306 11.304 22.68 ; 
      RECT 10.768 18.306 10.872 22.68 ; 
      RECT 10.336 18.306 10.44 22.68 ; 
      RECT 9.904 18.306 10.008 22.68 ; 
      RECT 9.472 18.306 9.576 22.68 ; 
      RECT 9.04 18.306 9.144 22.68 ; 
      RECT 8.608 18.306 8.712 22.68 ; 
      RECT 8.176 18.306 8.28 22.68 ; 
      RECT 7.744 18.306 7.848 22.68 ; 
      RECT 7.312 18.306 7.416 22.68 ; 
      RECT 6.88 18.306 6.984 22.68 ; 
      RECT 6.448 18.306 6.552 22.68 ; 
      RECT 6.016 18.306 6.12 22.68 ; 
      RECT 5.584 18.306 5.688 22.68 ; 
      RECT 5.152 18.306 5.256 22.68 ; 
      RECT 4.72 18.306 4.824 22.68 ; 
      RECT 4.288 18.306 4.392 22.68 ; 
      RECT 3.856 18.306 3.96 22.68 ; 
      RECT 3.424 18.306 3.528 22.68 ; 
      RECT 2.992 18.306 3.096 22.68 ; 
      RECT 2.56 18.306 2.664 22.68 ; 
      RECT 2.128 18.306 2.232 22.68 ; 
      RECT 1.696 18.306 1.8 22.68 ; 
      RECT 1.264 18.306 1.368 22.68 ; 
      RECT 0.832 18.306 0.936 22.68 ; 
      RECT 0.02 18.306 0.36 22.68 ; 
      RECT 34.564 22.626 35.076 27 ; 
      RECT 34.508 25.288 35.076 26.578 ; 
      RECT 33.916 24.196 34.164 27 ; 
      RECT 33.86 25.434 34.164 26.048 ; 
      RECT 33.916 22.626 34.02 27 ; 
      RECT 33.916 23.11 34.076 24.068 ; 
      RECT 33.916 22.626 34.164 22.982 ; 
      RECT 32.728 24.428 33.552 27 ; 
      RECT 33.448 22.626 33.552 27 ; 
      RECT 32.728 25.536 33.608 26.568 ; 
      RECT 32.728 22.626 33.12 27 ; 
      RECT 31.06 22.626 31.392 27 ; 
      RECT 31.06 22.98 31.448 26.722 ; 
      RECT 65.776 22.626 66.116 27 ; 
      RECT 65.2 22.626 65.304 27 ; 
      RECT 64.768 22.626 64.872 27 ; 
      RECT 64.336 22.626 64.44 27 ; 
      RECT 63.904 22.626 64.008 27 ; 
      RECT 63.472 22.626 63.576 27 ; 
      RECT 63.04 22.626 63.144 27 ; 
      RECT 62.608 22.626 62.712 27 ; 
      RECT 62.176 22.626 62.28 27 ; 
      RECT 61.744 22.626 61.848 27 ; 
      RECT 61.312 22.626 61.416 27 ; 
      RECT 60.88 22.626 60.984 27 ; 
      RECT 60.448 22.626 60.552 27 ; 
      RECT 60.016 22.626 60.12 27 ; 
      RECT 59.584 22.626 59.688 27 ; 
      RECT 59.152 22.626 59.256 27 ; 
      RECT 58.72 22.626 58.824 27 ; 
      RECT 58.288 22.626 58.392 27 ; 
      RECT 57.856 22.626 57.96 27 ; 
      RECT 57.424 22.626 57.528 27 ; 
      RECT 56.992 22.626 57.096 27 ; 
      RECT 56.56 22.626 56.664 27 ; 
      RECT 56.128 22.626 56.232 27 ; 
      RECT 55.696 22.626 55.8 27 ; 
      RECT 55.264 22.626 55.368 27 ; 
      RECT 54.832 22.626 54.936 27 ; 
      RECT 54.4 22.626 54.504 27 ; 
      RECT 53.968 22.626 54.072 27 ; 
      RECT 53.536 22.626 53.64 27 ; 
      RECT 53.104 22.626 53.208 27 ; 
      RECT 52.672 22.626 52.776 27 ; 
      RECT 52.24 22.626 52.344 27 ; 
      RECT 51.808 22.626 51.912 27 ; 
      RECT 51.376 22.626 51.48 27 ; 
      RECT 50.944 22.626 51.048 27 ; 
      RECT 50.512 22.626 50.616 27 ; 
      RECT 50.08 22.626 50.184 27 ; 
      RECT 49.648 22.626 49.752 27 ; 
      RECT 49.216 22.626 49.32 27 ; 
      RECT 48.784 22.626 48.888 27 ; 
      RECT 48.352 22.626 48.456 27 ; 
      RECT 47.92 22.626 48.024 27 ; 
      RECT 47.488 22.626 47.592 27 ; 
      RECT 47.056 22.626 47.16 27 ; 
      RECT 46.624 22.626 46.728 27 ; 
      RECT 46.192 22.626 46.296 27 ; 
      RECT 45.76 22.626 45.864 27 ; 
      RECT 45.328 22.626 45.432 27 ; 
      RECT 44.896 22.626 45 27 ; 
      RECT 44.464 22.626 44.568 27 ; 
      RECT 44.032 22.626 44.136 27 ; 
      RECT 43.6 22.626 43.704 27 ; 
      RECT 43.168 22.626 43.272 27 ; 
      RECT 42.736 22.626 42.84 27 ; 
      RECT 42.304 22.626 42.408 27 ; 
      RECT 41.872 22.626 41.976 27 ; 
      RECT 41.44 22.626 41.544 27 ; 
      RECT 41.008 22.626 41.112 27 ; 
      RECT 40.576 22.626 40.68 27 ; 
      RECT 40.144 22.626 40.248 27 ; 
      RECT 39.712 22.626 39.816 27 ; 
      RECT 39.28 22.626 39.384 27 ; 
      RECT 38.848 22.626 38.952 27 ; 
      RECT 38.416 22.626 38.52 27 ; 
      RECT 37.984 22.626 38.088 27 ; 
      RECT 37.552 22.626 37.656 27 ; 
      RECT 36.7 22.626 37.008 27 ; 
      RECT 29.128 22.626 29.436 27 ; 
      RECT 28.48 22.626 28.584 27 ; 
      RECT 28.048 22.626 28.152 27 ; 
      RECT 27.616 22.626 27.72 27 ; 
      RECT 27.184 22.626 27.288 27 ; 
      RECT 26.752 22.626 26.856 27 ; 
      RECT 26.32 22.626 26.424 27 ; 
      RECT 25.888 22.626 25.992 27 ; 
      RECT 25.456 22.626 25.56 27 ; 
      RECT 25.024 22.626 25.128 27 ; 
      RECT 24.592 22.626 24.696 27 ; 
      RECT 24.16 22.626 24.264 27 ; 
      RECT 23.728 22.626 23.832 27 ; 
      RECT 23.296 22.626 23.4 27 ; 
      RECT 22.864 22.626 22.968 27 ; 
      RECT 22.432 22.626 22.536 27 ; 
      RECT 22 22.626 22.104 27 ; 
      RECT 21.568 22.626 21.672 27 ; 
      RECT 21.136 22.626 21.24 27 ; 
      RECT 20.704 22.626 20.808 27 ; 
      RECT 20.272 22.626 20.376 27 ; 
      RECT 19.84 22.626 19.944 27 ; 
      RECT 19.408 22.626 19.512 27 ; 
      RECT 18.976 22.626 19.08 27 ; 
      RECT 18.544 22.626 18.648 27 ; 
      RECT 18.112 22.626 18.216 27 ; 
      RECT 17.68 22.626 17.784 27 ; 
      RECT 17.248 22.626 17.352 27 ; 
      RECT 16.816 22.626 16.92 27 ; 
      RECT 16.384 22.626 16.488 27 ; 
      RECT 15.952 22.626 16.056 27 ; 
      RECT 15.52 22.626 15.624 27 ; 
      RECT 15.088 22.626 15.192 27 ; 
      RECT 14.656 22.626 14.76 27 ; 
      RECT 14.224 22.626 14.328 27 ; 
      RECT 13.792 22.626 13.896 27 ; 
      RECT 13.36 22.626 13.464 27 ; 
      RECT 12.928 22.626 13.032 27 ; 
      RECT 12.496 22.626 12.6 27 ; 
      RECT 12.064 22.626 12.168 27 ; 
      RECT 11.632 22.626 11.736 27 ; 
      RECT 11.2 22.626 11.304 27 ; 
      RECT 10.768 22.626 10.872 27 ; 
      RECT 10.336 22.626 10.44 27 ; 
      RECT 9.904 22.626 10.008 27 ; 
      RECT 9.472 22.626 9.576 27 ; 
      RECT 9.04 22.626 9.144 27 ; 
      RECT 8.608 22.626 8.712 27 ; 
      RECT 8.176 22.626 8.28 27 ; 
      RECT 7.744 22.626 7.848 27 ; 
      RECT 7.312 22.626 7.416 27 ; 
      RECT 6.88 22.626 6.984 27 ; 
      RECT 6.448 22.626 6.552 27 ; 
      RECT 6.016 22.626 6.12 27 ; 
      RECT 5.584 22.626 5.688 27 ; 
      RECT 5.152 22.626 5.256 27 ; 
      RECT 4.72 22.626 4.824 27 ; 
      RECT 4.288 22.626 4.392 27 ; 
      RECT 3.856 22.626 3.96 27 ; 
      RECT 3.424 22.626 3.528 27 ; 
      RECT 2.992 22.626 3.096 27 ; 
      RECT 2.56 22.626 2.664 27 ; 
      RECT 2.128 22.626 2.232 27 ; 
      RECT 1.696 22.626 1.8 27 ; 
      RECT 1.264 22.626 1.368 27 ; 
      RECT 0.832 22.626 0.936 27 ; 
      RECT 0.02 22.626 0.36 27 ; 
      RECT 34.564 26.946 35.076 31.32 ; 
      RECT 34.508 29.608 35.076 30.898 ; 
      RECT 33.916 28.516 34.164 31.32 ; 
      RECT 33.86 29.754 34.164 30.368 ; 
      RECT 33.916 26.946 34.02 31.32 ; 
      RECT 33.916 27.43 34.076 28.388 ; 
      RECT 33.916 26.946 34.164 27.302 ; 
      RECT 32.728 28.748 33.552 31.32 ; 
      RECT 33.448 26.946 33.552 31.32 ; 
      RECT 32.728 29.856 33.608 30.888 ; 
      RECT 32.728 26.946 33.12 31.32 ; 
      RECT 31.06 26.946 31.392 31.32 ; 
      RECT 31.06 27.3 31.448 31.042 ; 
      RECT 65.776 26.946 66.116 31.32 ; 
      RECT 65.2 26.946 65.304 31.32 ; 
      RECT 64.768 26.946 64.872 31.32 ; 
      RECT 64.336 26.946 64.44 31.32 ; 
      RECT 63.904 26.946 64.008 31.32 ; 
      RECT 63.472 26.946 63.576 31.32 ; 
      RECT 63.04 26.946 63.144 31.32 ; 
      RECT 62.608 26.946 62.712 31.32 ; 
      RECT 62.176 26.946 62.28 31.32 ; 
      RECT 61.744 26.946 61.848 31.32 ; 
      RECT 61.312 26.946 61.416 31.32 ; 
      RECT 60.88 26.946 60.984 31.32 ; 
      RECT 60.448 26.946 60.552 31.32 ; 
      RECT 60.016 26.946 60.12 31.32 ; 
      RECT 59.584 26.946 59.688 31.32 ; 
      RECT 59.152 26.946 59.256 31.32 ; 
      RECT 58.72 26.946 58.824 31.32 ; 
      RECT 58.288 26.946 58.392 31.32 ; 
      RECT 57.856 26.946 57.96 31.32 ; 
      RECT 57.424 26.946 57.528 31.32 ; 
      RECT 56.992 26.946 57.096 31.32 ; 
      RECT 56.56 26.946 56.664 31.32 ; 
      RECT 56.128 26.946 56.232 31.32 ; 
      RECT 55.696 26.946 55.8 31.32 ; 
      RECT 55.264 26.946 55.368 31.32 ; 
      RECT 54.832 26.946 54.936 31.32 ; 
      RECT 54.4 26.946 54.504 31.32 ; 
      RECT 53.968 26.946 54.072 31.32 ; 
      RECT 53.536 26.946 53.64 31.32 ; 
      RECT 53.104 26.946 53.208 31.32 ; 
      RECT 52.672 26.946 52.776 31.32 ; 
      RECT 52.24 26.946 52.344 31.32 ; 
      RECT 51.808 26.946 51.912 31.32 ; 
      RECT 51.376 26.946 51.48 31.32 ; 
      RECT 50.944 26.946 51.048 31.32 ; 
      RECT 50.512 26.946 50.616 31.32 ; 
      RECT 50.08 26.946 50.184 31.32 ; 
      RECT 49.648 26.946 49.752 31.32 ; 
      RECT 49.216 26.946 49.32 31.32 ; 
      RECT 48.784 26.946 48.888 31.32 ; 
      RECT 48.352 26.946 48.456 31.32 ; 
      RECT 47.92 26.946 48.024 31.32 ; 
      RECT 47.488 26.946 47.592 31.32 ; 
      RECT 47.056 26.946 47.16 31.32 ; 
      RECT 46.624 26.946 46.728 31.32 ; 
      RECT 46.192 26.946 46.296 31.32 ; 
      RECT 45.76 26.946 45.864 31.32 ; 
      RECT 45.328 26.946 45.432 31.32 ; 
      RECT 44.896 26.946 45 31.32 ; 
      RECT 44.464 26.946 44.568 31.32 ; 
      RECT 44.032 26.946 44.136 31.32 ; 
      RECT 43.6 26.946 43.704 31.32 ; 
      RECT 43.168 26.946 43.272 31.32 ; 
      RECT 42.736 26.946 42.84 31.32 ; 
      RECT 42.304 26.946 42.408 31.32 ; 
      RECT 41.872 26.946 41.976 31.32 ; 
      RECT 41.44 26.946 41.544 31.32 ; 
      RECT 41.008 26.946 41.112 31.32 ; 
      RECT 40.576 26.946 40.68 31.32 ; 
      RECT 40.144 26.946 40.248 31.32 ; 
      RECT 39.712 26.946 39.816 31.32 ; 
      RECT 39.28 26.946 39.384 31.32 ; 
      RECT 38.848 26.946 38.952 31.32 ; 
      RECT 38.416 26.946 38.52 31.32 ; 
      RECT 37.984 26.946 38.088 31.32 ; 
      RECT 37.552 26.946 37.656 31.32 ; 
      RECT 36.7 26.946 37.008 31.32 ; 
      RECT 29.128 26.946 29.436 31.32 ; 
      RECT 28.48 26.946 28.584 31.32 ; 
      RECT 28.048 26.946 28.152 31.32 ; 
      RECT 27.616 26.946 27.72 31.32 ; 
      RECT 27.184 26.946 27.288 31.32 ; 
      RECT 26.752 26.946 26.856 31.32 ; 
      RECT 26.32 26.946 26.424 31.32 ; 
      RECT 25.888 26.946 25.992 31.32 ; 
      RECT 25.456 26.946 25.56 31.32 ; 
      RECT 25.024 26.946 25.128 31.32 ; 
      RECT 24.592 26.946 24.696 31.32 ; 
      RECT 24.16 26.946 24.264 31.32 ; 
      RECT 23.728 26.946 23.832 31.32 ; 
      RECT 23.296 26.946 23.4 31.32 ; 
      RECT 22.864 26.946 22.968 31.32 ; 
      RECT 22.432 26.946 22.536 31.32 ; 
      RECT 22 26.946 22.104 31.32 ; 
      RECT 21.568 26.946 21.672 31.32 ; 
      RECT 21.136 26.946 21.24 31.32 ; 
      RECT 20.704 26.946 20.808 31.32 ; 
      RECT 20.272 26.946 20.376 31.32 ; 
      RECT 19.84 26.946 19.944 31.32 ; 
      RECT 19.408 26.946 19.512 31.32 ; 
      RECT 18.976 26.946 19.08 31.32 ; 
      RECT 18.544 26.946 18.648 31.32 ; 
      RECT 18.112 26.946 18.216 31.32 ; 
      RECT 17.68 26.946 17.784 31.32 ; 
      RECT 17.248 26.946 17.352 31.32 ; 
      RECT 16.816 26.946 16.92 31.32 ; 
      RECT 16.384 26.946 16.488 31.32 ; 
      RECT 15.952 26.946 16.056 31.32 ; 
      RECT 15.52 26.946 15.624 31.32 ; 
      RECT 15.088 26.946 15.192 31.32 ; 
      RECT 14.656 26.946 14.76 31.32 ; 
      RECT 14.224 26.946 14.328 31.32 ; 
      RECT 13.792 26.946 13.896 31.32 ; 
      RECT 13.36 26.946 13.464 31.32 ; 
      RECT 12.928 26.946 13.032 31.32 ; 
      RECT 12.496 26.946 12.6 31.32 ; 
      RECT 12.064 26.946 12.168 31.32 ; 
      RECT 11.632 26.946 11.736 31.32 ; 
      RECT 11.2 26.946 11.304 31.32 ; 
      RECT 10.768 26.946 10.872 31.32 ; 
      RECT 10.336 26.946 10.44 31.32 ; 
      RECT 9.904 26.946 10.008 31.32 ; 
      RECT 9.472 26.946 9.576 31.32 ; 
      RECT 9.04 26.946 9.144 31.32 ; 
      RECT 8.608 26.946 8.712 31.32 ; 
      RECT 8.176 26.946 8.28 31.32 ; 
      RECT 7.744 26.946 7.848 31.32 ; 
      RECT 7.312 26.946 7.416 31.32 ; 
      RECT 6.88 26.946 6.984 31.32 ; 
      RECT 6.448 26.946 6.552 31.32 ; 
      RECT 6.016 26.946 6.12 31.32 ; 
      RECT 5.584 26.946 5.688 31.32 ; 
      RECT 5.152 26.946 5.256 31.32 ; 
      RECT 4.72 26.946 4.824 31.32 ; 
      RECT 4.288 26.946 4.392 31.32 ; 
      RECT 3.856 26.946 3.96 31.32 ; 
      RECT 3.424 26.946 3.528 31.32 ; 
      RECT 2.992 26.946 3.096 31.32 ; 
      RECT 2.56 26.946 2.664 31.32 ; 
      RECT 2.128 26.946 2.232 31.32 ; 
      RECT 1.696 26.946 1.8 31.32 ; 
      RECT 1.264 26.946 1.368 31.32 ; 
      RECT 0.832 26.946 0.936 31.32 ; 
      RECT 0.02 26.946 0.36 31.32 ; 
      RECT 34.564 31.266 35.076 35.64 ; 
      RECT 34.508 33.928 35.076 35.218 ; 
      RECT 33.916 32.836 34.164 35.64 ; 
      RECT 33.86 34.074 34.164 34.688 ; 
      RECT 33.916 31.266 34.02 35.64 ; 
      RECT 33.916 31.75 34.076 32.708 ; 
      RECT 33.916 31.266 34.164 31.622 ; 
      RECT 32.728 33.068 33.552 35.64 ; 
      RECT 33.448 31.266 33.552 35.64 ; 
      RECT 32.728 34.176 33.608 35.208 ; 
      RECT 32.728 31.266 33.12 35.64 ; 
      RECT 31.06 31.266 31.392 35.64 ; 
      RECT 31.06 31.62 31.448 35.362 ; 
      RECT 65.776 31.266 66.116 35.64 ; 
      RECT 65.2 31.266 65.304 35.64 ; 
      RECT 64.768 31.266 64.872 35.64 ; 
      RECT 64.336 31.266 64.44 35.64 ; 
      RECT 63.904 31.266 64.008 35.64 ; 
      RECT 63.472 31.266 63.576 35.64 ; 
      RECT 63.04 31.266 63.144 35.64 ; 
      RECT 62.608 31.266 62.712 35.64 ; 
      RECT 62.176 31.266 62.28 35.64 ; 
      RECT 61.744 31.266 61.848 35.64 ; 
      RECT 61.312 31.266 61.416 35.64 ; 
      RECT 60.88 31.266 60.984 35.64 ; 
      RECT 60.448 31.266 60.552 35.64 ; 
      RECT 60.016 31.266 60.12 35.64 ; 
      RECT 59.584 31.266 59.688 35.64 ; 
      RECT 59.152 31.266 59.256 35.64 ; 
      RECT 58.72 31.266 58.824 35.64 ; 
      RECT 58.288 31.266 58.392 35.64 ; 
      RECT 57.856 31.266 57.96 35.64 ; 
      RECT 57.424 31.266 57.528 35.64 ; 
      RECT 56.992 31.266 57.096 35.64 ; 
      RECT 56.56 31.266 56.664 35.64 ; 
      RECT 56.128 31.266 56.232 35.64 ; 
      RECT 55.696 31.266 55.8 35.64 ; 
      RECT 55.264 31.266 55.368 35.64 ; 
      RECT 54.832 31.266 54.936 35.64 ; 
      RECT 54.4 31.266 54.504 35.64 ; 
      RECT 53.968 31.266 54.072 35.64 ; 
      RECT 53.536 31.266 53.64 35.64 ; 
      RECT 53.104 31.266 53.208 35.64 ; 
      RECT 52.672 31.266 52.776 35.64 ; 
      RECT 52.24 31.266 52.344 35.64 ; 
      RECT 51.808 31.266 51.912 35.64 ; 
      RECT 51.376 31.266 51.48 35.64 ; 
      RECT 50.944 31.266 51.048 35.64 ; 
      RECT 50.512 31.266 50.616 35.64 ; 
      RECT 50.08 31.266 50.184 35.64 ; 
      RECT 49.648 31.266 49.752 35.64 ; 
      RECT 49.216 31.266 49.32 35.64 ; 
      RECT 48.784 31.266 48.888 35.64 ; 
      RECT 48.352 31.266 48.456 35.64 ; 
      RECT 47.92 31.266 48.024 35.64 ; 
      RECT 47.488 31.266 47.592 35.64 ; 
      RECT 47.056 31.266 47.16 35.64 ; 
      RECT 46.624 31.266 46.728 35.64 ; 
      RECT 46.192 31.266 46.296 35.64 ; 
      RECT 45.76 31.266 45.864 35.64 ; 
      RECT 45.328 31.266 45.432 35.64 ; 
      RECT 44.896 31.266 45 35.64 ; 
      RECT 44.464 31.266 44.568 35.64 ; 
      RECT 44.032 31.266 44.136 35.64 ; 
      RECT 43.6 31.266 43.704 35.64 ; 
      RECT 43.168 31.266 43.272 35.64 ; 
      RECT 42.736 31.266 42.84 35.64 ; 
      RECT 42.304 31.266 42.408 35.64 ; 
      RECT 41.872 31.266 41.976 35.64 ; 
      RECT 41.44 31.266 41.544 35.64 ; 
      RECT 41.008 31.266 41.112 35.64 ; 
      RECT 40.576 31.266 40.68 35.64 ; 
      RECT 40.144 31.266 40.248 35.64 ; 
      RECT 39.712 31.266 39.816 35.64 ; 
      RECT 39.28 31.266 39.384 35.64 ; 
      RECT 38.848 31.266 38.952 35.64 ; 
      RECT 38.416 31.266 38.52 35.64 ; 
      RECT 37.984 31.266 38.088 35.64 ; 
      RECT 37.552 31.266 37.656 35.64 ; 
      RECT 36.7 31.266 37.008 35.64 ; 
      RECT 29.128 31.266 29.436 35.64 ; 
      RECT 28.48 31.266 28.584 35.64 ; 
      RECT 28.048 31.266 28.152 35.64 ; 
      RECT 27.616 31.266 27.72 35.64 ; 
      RECT 27.184 31.266 27.288 35.64 ; 
      RECT 26.752 31.266 26.856 35.64 ; 
      RECT 26.32 31.266 26.424 35.64 ; 
      RECT 25.888 31.266 25.992 35.64 ; 
      RECT 25.456 31.266 25.56 35.64 ; 
      RECT 25.024 31.266 25.128 35.64 ; 
      RECT 24.592 31.266 24.696 35.64 ; 
      RECT 24.16 31.266 24.264 35.64 ; 
      RECT 23.728 31.266 23.832 35.64 ; 
      RECT 23.296 31.266 23.4 35.64 ; 
      RECT 22.864 31.266 22.968 35.64 ; 
      RECT 22.432 31.266 22.536 35.64 ; 
      RECT 22 31.266 22.104 35.64 ; 
      RECT 21.568 31.266 21.672 35.64 ; 
      RECT 21.136 31.266 21.24 35.64 ; 
      RECT 20.704 31.266 20.808 35.64 ; 
      RECT 20.272 31.266 20.376 35.64 ; 
      RECT 19.84 31.266 19.944 35.64 ; 
      RECT 19.408 31.266 19.512 35.64 ; 
      RECT 18.976 31.266 19.08 35.64 ; 
      RECT 18.544 31.266 18.648 35.64 ; 
      RECT 18.112 31.266 18.216 35.64 ; 
      RECT 17.68 31.266 17.784 35.64 ; 
      RECT 17.248 31.266 17.352 35.64 ; 
      RECT 16.816 31.266 16.92 35.64 ; 
      RECT 16.384 31.266 16.488 35.64 ; 
      RECT 15.952 31.266 16.056 35.64 ; 
      RECT 15.52 31.266 15.624 35.64 ; 
      RECT 15.088 31.266 15.192 35.64 ; 
      RECT 14.656 31.266 14.76 35.64 ; 
      RECT 14.224 31.266 14.328 35.64 ; 
      RECT 13.792 31.266 13.896 35.64 ; 
      RECT 13.36 31.266 13.464 35.64 ; 
      RECT 12.928 31.266 13.032 35.64 ; 
      RECT 12.496 31.266 12.6 35.64 ; 
      RECT 12.064 31.266 12.168 35.64 ; 
      RECT 11.632 31.266 11.736 35.64 ; 
      RECT 11.2 31.266 11.304 35.64 ; 
      RECT 10.768 31.266 10.872 35.64 ; 
      RECT 10.336 31.266 10.44 35.64 ; 
      RECT 9.904 31.266 10.008 35.64 ; 
      RECT 9.472 31.266 9.576 35.64 ; 
      RECT 9.04 31.266 9.144 35.64 ; 
      RECT 8.608 31.266 8.712 35.64 ; 
      RECT 8.176 31.266 8.28 35.64 ; 
      RECT 7.744 31.266 7.848 35.64 ; 
      RECT 7.312 31.266 7.416 35.64 ; 
      RECT 6.88 31.266 6.984 35.64 ; 
      RECT 6.448 31.266 6.552 35.64 ; 
      RECT 6.016 31.266 6.12 35.64 ; 
      RECT 5.584 31.266 5.688 35.64 ; 
      RECT 5.152 31.266 5.256 35.64 ; 
      RECT 4.72 31.266 4.824 35.64 ; 
      RECT 4.288 31.266 4.392 35.64 ; 
      RECT 3.856 31.266 3.96 35.64 ; 
      RECT 3.424 31.266 3.528 35.64 ; 
      RECT 2.992 31.266 3.096 35.64 ; 
      RECT 2.56 31.266 2.664 35.64 ; 
      RECT 2.128 31.266 2.232 35.64 ; 
      RECT 1.696 31.266 1.8 35.64 ; 
      RECT 1.264 31.266 1.368 35.64 ; 
      RECT 0.832 31.266 0.936 35.64 ; 
      RECT 0.02 31.266 0.36 35.64 ; 
      RECT 34.564 35.586 35.076 39.96 ; 
      RECT 34.508 38.248 35.076 39.538 ; 
      RECT 33.916 37.156 34.164 39.96 ; 
      RECT 33.86 38.394 34.164 39.008 ; 
      RECT 33.916 35.586 34.02 39.96 ; 
      RECT 33.916 36.07 34.076 37.028 ; 
      RECT 33.916 35.586 34.164 35.942 ; 
      RECT 32.728 37.388 33.552 39.96 ; 
      RECT 33.448 35.586 33.552 39.96 ; 
      RECT 32.728 38.496 33.608 39.528 ; 
      RECT 32.728 35.586 33.12 39.96 ; 
      RECT 31.06 35.586 31.392 39.96 ; 
      RECT 31.06 35.94 31.448 39.682 ; 
      RECT 65.776 35.586 66.116 39.96 ; 
      RECT 65.2 35.586 65.304 39.96 ; 
      RECT 64.768 35.586 64.872 39.96 ; 
      RECT 64.336 35.586 64.44 39.96 ; 
      RECT 63.904 35.586 64.008 39.96 ; 
      RECT 63.472 35.586 63.576 39.96 ; 
      RECT 63.04 35.586 63.144 39.96 ; 
      RECT 62.608 35.586 62.712 39.96 ; 
      RECT 62.176 35.586 62.28 39.96 ; 
      RECT 61.744 35.586 61.848 39.96 ; 
      RECT 61.312 35.586 61.416 39.96 ; 
      RECT 60.88 35.586 60.984 39.96 ; 
      RECT 60.448 35.586 60.552 39.96 ; 
      RECT 60.016 35.586 60.12 39.96 ; 
      RECT 59.584 35.586 59.688 39.96 ; 
      RECT 59.152 35.586 59.256 39.96 ; 
      RECT 58.72 35.586 58.824 39.96 ; 
      RECT 58.288 35.586 58.392 39.96 ; 
      RECT 57.856 35.586 57.96 39.96 ; 
      RECT 57.424 35.586 57.528 39.96 ; 
      RECT 56.992 35.586 57.096 39.96 ; 
      RECT 56.56 35.586 56.664 39.96 ; 
      RECT 56.128 35.586 56.232 39.96 ; 
      RECT 55.696 35.586 55.8 39.96 ; 
      RECT 55.264 35.586 55.368 39.96 ; 
      RECT 54.832 35.586 54.936 39.96 ; 
      RECT 54.4 35.586 54.504 39.96 ; 
      RECT 53.968 35.586 54.072 39.96 ; 
      RECT 53.536 35.586 53.64 39.96 ; 
      RECT 53.104 35.586 53.208 39.96 ; 
      RECT 52.672 35.586 52.776 39.96 ; 
      RECT 52.24 35.586 52.344 39.96 ; 
      RECT 51.808 35.586 51.912 39.96 ; 
      RECT 51.376 35.586 51.48 39.96 ; 
      RECT 50.944 35.586 51.048 39.96 ; 
      RECT 50.512 35.586 50.616 39.96 ; 
      RECT 50.08 35.586 50.184 39.96 ; 
      RECT 49.648 35.586 49.752 39.96 ; 
      RECT 49.216 35.586 49.32 39.96 ; 
      RECT 48.784 35.586 48.888 39.96 ; 
      RECT 48.352 35.586 48.456 39.96 ; 
      RECT 47.92 35.586 48.024 39.96 ; 
      RECT 47.488 35.586 47.592 39.96 ; 
      RECT 47.056 35.586 47.16 39.96 ; 
      RECT 46.624 35.586 46.728 39.96 ; 
      RECT 46.192 35.586 46.296 39.96 ; 
      RECT 45.76 35.586 45.864 39.96 ; 
      RECT 45.328 35.586 45.432 39.96 ; 
      RECT 44.896 35.586 45 39.96 ; 
      RECT 44.464 35.586 44.568 39.96 ; 
      RECT 44.032 35.586 44.136 39.96 ; 
      RECT 43.6 35.586 43.704 39.96 ; 
      RECT 43.168 35.586 43.272 39.96 ; 
      RECT 42.736 35.586 42.84 39.96 ; 
      RECT 42.304 35.586 42.408 39.96 ; 
      RECT 41.872 35.586 41.976 39.96 ; 
      RECT 41.44 35.586 41.544 39.96 ; 
      RECT 41.008 35.586 41.112 39.96 ; 
      RECT 40.576 35.586 40.68 39.96 ; 
      RECT 40.144 35.586 40.248 39.96 ; 
      RECT 39.712 35.586 39.816 39.96 ; 
      RECT 39.28 35.586 39.384 39.96 ; 
      RECT 38.848 35.586 38.952 39.96 ; 
      RECT 38.416 35.586 38.52 39.96 ; 
      RECT 37.984 35.586 38.088 39.96 ; 
      RECT 37.552 35.586 37.656 39.96 ; 
      RECT 36.7 35.586 37.008 39.96 ; 
      RECT 29.128 35.586 29.436 39.96 ; 
      RECT 28.48 35.586 28.584 39.96 ; 
      RECT 28.048 35.586 28.152 39.96 ; 
      RECT 27.616 35.586 27.72 39.96 ; 
      RECT 27.184 35.586 27.288 39.96 ; 
      RECT 26.752 35.586 26.856 39.96 ; 
      RECT 26.32 35.586 26.424 39.96 ; 
      RECT 25.888 35.586 25.992 39.96 ; 
      RECT 25.456 35.586 25.56 39.96 ; 
      RECT 25.024 35.586 25.128 39.96 ; 
      RECT 24.592 35.586 24.696 39.96 ; 
      RECT 24.16 35.586 24.264 39.96 ; 
      RECT 23.728 35.586 23.832 39.96 ; 
      RECT 23.296 35.586 23.4 39.96 ; 
      RECT 22.864 35.586 22.968 39.96 ; 
      RECT 22.432 35.586 22.536 39.96 ; 
      RECT 22 35.586 22.104 39.96 ; 
      RECT 21.568 35.586 21.672 39.96 ; 
      RECT 21.136 35.586 21.24 39.96 ; 
      RECT 20.704 35.586 20.808 39.96 ; 
      RECT 20.272 35.586 20.376 39.96 ; 
      RECT 19.84 35.586 19.944 39.96 ; 
      RECT 19.408 35.586 19.512 39.96 ; 
      RECT 18.976 35.586 19.08 39.96 ; 
      RECT 18.544 35.586 18.648 39.96 ; 
      RECT 18.112 35.586 18.216 39.96 ; 
      RECT 17.68 35.586 17.784 39.96 ; 
      RECT 17.248 35.586 17.352 39.96 ; 
      RECT 16.816 35.586 16.92 39.96 ; 
      RECT 16.384 35.586 16.488 39.96 ; 
      RECT 15.952 35.586 16.056 39.96 ; 
      RECT 15.52 35.586 15.624 39.96 ; 
      RECT 15.088 35.586 15.192 39.96 ; 
      RECT 14.656 35.586 14.76 39.96 ; 
      RECT 14.224 35.586 14.328 39.96 ; 
      RECT 13.792 35.586 13.896 39.96 ; 
      RECT 13.36 35.586 13.464 39.96 ; 
      RECT 12.928 35.586 13.032 39.96 ; 
      RECT 12.496 35.586 12.6 39.96 ; 
      RECT 12.064 35.586 12.168 39.96 ; 
      RECT 11.632 35.586 11.736 39.96 ; 
      RECT 11.2 35.586 11.304 39.96 ; 
      RECT 10.768 35.586 10.872 39.96 ; 
      RECT 10.336 35.586 10.44 39.96 ; 
      RECT 9.904 35.586 10.008 39.96 ; 
      RECT 9.472 35.586 9.576 39.96 ; 
      RECT 9.04 35.586 9.144 39.96 ; 
      RECT 8.608 35.586 8.712 39.96 ; 
      RECT 8.176 35.586 8.28 39.96 ; 
      RECT 7.744 35.586 7.848 39.96 ; 
      RECT 7.312 35.586 7.416 39.96 ; 
      RECT 6.88 35.586 6.984 39.96 ; 
      RECT 6.448 35.586 6.552 39.96 ; 
      RECT 6.016 35.586 6.12 39.96 ; 
      RECT 5.584 35.586 5.688 39.96 ; 
      RECT 5.152 35.586 5.256 39.96 ; 
      RECT 4.72 35.586 4.824 39.96 ; 
      RECT 4.288 35.586 4.392 39.96 ; 
      RECT 3.856 35.586 3.96 39.96 ; 
      RECT 3.424 35.586 3.528 39.96 ; 
      RECT 2.992 35.586 3.096 39.96 ; 
      RECT 2.56 35.586 2.664 39.96 ; 
      RECT 2.128 35.586 2.232 39.96 ; 
      RECT 1.696 35.586 1.8 39.96 ; 
      RECT 1.264 35.586 1.368 39.96 ; 
      RECT 0.832 35.586 0.936 39.96 ; 
      RECT 0.02 35.586 0.36 39.96 ; 
      RECT 34.564 39.906 35.076 44.28 ; 
      RECT 34.508 42.568 35.076 43.858 ; 
      RECT 33.916 41.476 34.164 44.28 ; 
      RECT 33.86 42.714 34.164 43.328 ; 
      RECT 33.916 39.906 34.02 44.28 ; 
      RECT 33.916 40.39 34.076 41.348 ; 
      RECT 33.916 39.906 34.164 40.262 ; 
      RECT 32.728 41.708 33.552 44.28 ; 
      RECT 33.448 39.906 33.552 44.28 ; 
      RECT 32.728 42.816 33.608 43.848 ; 
      RECT 32.728 39.906 33.12 44.28 ; 
      RECT 31.06 39.906 31.392 44.28 ; 
      RECT 31.06 40.26 31.448 44.002 ; 
      RECT 65.776 39.906 66.116 44.28 ; 
      RECT 65.2 39.906 65.304 44.28 ; 
      RECT 64.768 39.906 64.872 44.28 ; 
      RECT 64.336 39.906 64.44 44.28 ; 
      RECT 63.904 39.906 64.008 44.28 ; 
      RECT 63.472 39.906 63.576 44.28 ; 
      RECT 63.04 39.906 63.144 44.28 ; 
      RECT 62.608 39.906 62.712 44.28 ; 
      RECT 62.176 39.906 62.28 44.28 ; 
      RECT 61.744 39.906 61.848 44.28 ; 
      RECT 61.312 39.906 61.416 44.28 ; 
      RECT 60.88 39.906 60.984 44.28 ; 
      RECT 60.448 39.906 60.552 44.28 ; 
      RECT 60.016 39.906 60.12 44.28 ; 
      RECT 59.584 39.906 59.688 44.28 ; 
      RECT 59.152 39.906 59.256 44.28 ; 
      RECT 58.72 39.906 58.824 44.28 ; 
      RECT 58.288 39.906 58.392 44.28 ; 
      RECT 57.856 39.906 57.96 44.28 ; 
      RECT 57.424 39.906 57.528 44.28 ; 
      RECT 56.992 39.906 57.096 44.28 ; 
      RECT 56.56 39.906 56.664 44.28 ; 
      RECT 56.128 39.906 56.232 44.28 ; 
      RECT 55.696 39.906 55.8 44.28 ; 
      RECT 55.264 39.906 55.368 44.28 ; 
      RECT 54.832 39.906 54.936 44.28 ; 
      RECT 54.4 39.906 54.504 44.28 ; 
      RECT 53.968 39.906 54.072 44.28 ; 
      RECT 53.536 39.906 53.64 44.28 ; 
      RECT 53.104 39.906 53.208 44.28 ; 
      RECT 52.672 39.906 52.776 44.28 ; 
      RECT 52.24 39.906 52.344 44.28 ; 
      RECT 51.808 39.906 51.912 44.28 ; 
      RECT 51.376 39.906 51.48 44.28 ; 
      RECT 50.944 39.906 51.048 44.28 ; 
      RECT 50.512 39.906 50.616 44.28 ; 
      RECT 50.08 39.906 50.184 44.28 ; 
      RECT 49.648 39.906 49.752 44.28 ; 
      RECT 49.216 39.906 49.32 44.28 ; 
      RECT 48.784 39.906 48.888 44.28 ; 
      RECT 48.352 39.906 48.456 44.28 ; 
      RECT 47.92 39.906 48.024 44.28 ; 
      RECT 47.488 39.906 47.592 44.28 ; 
      RECT 47.056 39.906 47.16 44.28 ; 
      RECT 46.624 39.906 46.728 44.28 ; 
      RECT 46.192 39.906 46.296 44.28 ; 
      RECT 45.76 39.906 45.864 44.28 ; 
      RECT 45.328 39.906 45.432 44.28 ; 
      RECT 44.896 39.906 45 44.28 ; 
      RECT 44.464 39.906 44.568 44.28 ; 
      RECT 44.032 39.906 44.136 44.28 ; 
      RECT 43.6 39.906 43.704 44.28 ; 
      RECT 43.168 39.906 43.272 44.28 ; 
      RECT 42.736 39.906 42.84 44.28 ; 
      RECT 42.304 39.906 42.408 44.28 ; 
      RECT 41.872 39.906 41.976 44.28 ; 
      RECT 41.44 39.906 41.544 44.28 ; 
      RECT 41.008 39.906 41.112 44.28 ; 
      RECT 40.576 39.906 40.68 44.28 ; 
      RECT 40.144 39.906 40.248 44.28 ; 
      RECT 39.712 39.906 39.816 44.28 ; 
      RECT 39.28 39.906 39.384 44.28 ; 
      RECT 38.848 39.906 38.952 44.28 ; 
      RECT 38.416 39.906 38.52 44.28 ; 
      RECT 37.984 39.906 38.088 44.28 ; 
      RECT 37.552 39.906 37.656 44.28 ; 
      RECT 36.7 39.906 37.008 44.28 ; 
      RECT 29.128 39.906 29.436 44.28 ; 
      RECT 28.48 39.906 28.584 44.28 ; 
      RECT 28.048 39.906 28.152 44.28 ; 
      RECT 27.616 39.906 27.72 44.28 ; 
      RECT 27.184 39.906 27.288 44.28 ; 
      RECT 26.752 39.906 26.856 44.28 ; 
      RECT 26.32 39.906 26.424 44.28 ; 
      RECT 25.888 39.906 25.992 44.28 ; 
      RECT 25.456 39.906 25.56 44.28 ; 
      RECT 25.024 39.906 25.128 44.28 ; 
      RECT 24.592 39.906 24.696 44.28 ; 
      RECT 24.16 39.906 24.264 44.28 ; 
      RECT 23.728 39.906 23.832 44.28 ; 
      RECT 23.296 39.906 23.4 44.28 ; 
      RECT 22.864 39.906 22.968 44.28 ; 
      RECT 22.432 39.906 22.536 44.28 ; 
      RECT 22 39.906 22.104 44.28 ; 
      RECT 21.568 39.906 21.672 44.28 ; 
      RECT 21.136 39.906 21.24 44.28 ; 
      RECT 20.704 39.906 20.808 44.28 ; 
      RECT 20.272 39.906 20.376 44.28 ; 
      RECT 19.84 39.906 19.944 44.28 ; 
      RECT 19.408 39.906 19.512 44.28 ; 
      RECT 18.976 39.906 19.08 44.28 ; 
      RECT 18.544 39.906 18.648 44.28 ; 
      RECT 18.112 39.906 18.216 44.28 ; 
      RECT 17.68 39.906 17.784 44.28 ; 
      RECT 17.248 39.906 17.352 44.28 ; 
      RECT 16.816 39.906 16.92 44.28 ; 
      RECT 16.384 39.906 16.488 44.28 ; 
      RECT 15.952 39.906 16.056 44.28 ; 
      RECT 15.52 39.906 15.624 44.28 ; 
      RECT 15.088 39.906 15.192 44.28 ; 
      RECT 14.656 39.906 14.76 44.28 ; 
      RECT 14.224 39.906 14.328 44.28 ; 
      RECT 13.792 39.906 13.896 44.28 ; 
      RECT 13.36 39.906 13.464 44.28 ; 
      RECT 12.928 39.906 13.032 44.28 ; 
      RECT 12.496 39.906 12.6 44.28 ; 
      RECT 12.064 39.906 12.168 44.28 ; 
      RECT 11.632 39.906 11.736 44.28 ; 
      RECT 11.2 39.906 11.304 44.28 ; 
      RECT 10.768 39.906 10.872 44.28 ; 
      RECT 10.336 39.906 10.44 44.28 ; 
      RECT 9.904 39.906 10.008 44.28 ; 
      RECT 9.472 39.906 9.576 44.28 ; 
      RECT 9.04 39.906 9.144 44.28 ; 
      RECT 8.608 39.906 8.712 44.28 ; 
      RECT 8.176 39.906 8.28 44.28 ; 
      RECT 7.744 39.906 7.848 44.28 ; 
      RECT 7.312 39.906 7.416 44.28 ; 
      RECT 6.88 39.906 6.984 44.28 ; 
      RECT 6.448 39.906 6.552 44.28 ; 
      RECT 6.016 39.906 6.12 44.28 ; 
      RECT 5.584 39.906 5.688 44.28 ; 
      RECT 5.152 39.906 5.256 44.28 ; 
      RECT 4.72 39.906 4.824 44.28 ; 
      RECT 4.288 39.906 4.392 44.28 ; 
      RECT 3.856 39.906 3.96 44.28 ; 
      RECT 3.424 39.906 3.528 44.28 ; 
      RECT 2.992 39.906 3.096 44.28 ; 
      RECT 2.56 39.906 2.664 44.28 ; 
      RECT 2.128 39.906 2.232 44.28 ; 
      RECT 1.696 39.906 1.8 44.28 ; 
      RECT 1.264 39.906 1.368 44.28 ; 
      RECT 0.832 39.906 0.936 44.28 ; 
      RECT 0.02 39.906 0.36 44.28 ; 
      RECT 34.564 44.226 35.076 48.6 ; 
      RECT 34.508 46.888 35.076 48.178 ; 
      RECT 33.916 45.796 34.164 48.6 ; 
      RECT 33.86 47.034 34.164 47.648 ; 
      RECT 33.916 44.226 34.02 48.6 ; 
      RECT 33.916 44.71 34.076 45.668 ; 
      RECT 33.916 44.226 34.164 44.582 ; 
      RECT 32.728 46.028 33.552 48.6 ; 
      RECT 33.448 44.226 33.552 48.6 ; 
      RECT 32.728 47.136 33.608 48.168 ; 
      RECT 32.728 44.226 33.12 48.6 ; 
      RECT 31.06 44.226 31.392 48.6 ; 
      RECT 31.06 44.58 31.448 48.322 ; 
      RECT 65.776 44.226 66.116 48.6 ; 
      RECT 65.2 44.226 65.304 48.6 ; 
      RECT 64.768 44.226 64.872 48.6 ; 
      RECT 64.336 44.226 64.44 48.6 ; 
      RECT 63.904 44.226 64.008 48.6 ; 
      RECT 63.472 44.226 63.576 48.6 ; 
      RECT 63.04 44.226 63.144 48.6 ; 
      RECT 62.608 44.226 62.712 48.6 ; 
      RECT 62.176 44.226 62.28 48.6 ; 
      RECT 61.744 44.226 61.848 48.6 ; 
      RECT 61.312 44.226 61.416 48.6 ; 
      RECT 60.88 44.226 60.984 48.6 ; 
      RECT 60.448 44.226 60.552 48.6 ; 
      RECT 60.016 44.226 60.12 48.6 ; 
      RECT 59.584 44.226 59.688 48.6 ; 
      RECT 59.152 44.226 59.256 48.6 ; 
      RECT 58.72 44.226 58.824 48.6 ; 
      RECT 58.288 44.226 58.392 48.6 ; 
      RECT 57.856 44.226 57.96 48.6 ; 
      RECT 57.424 44.226 57.528 48.6 ; 
      RECT 56.992 44.226 57.096 48.6 ; 
      RECT 56.56 44.226 56.664 48.6 ; 
      RECT 56.128 44.226 56.232 48.6 ; 
      RECT 55.696 44.226 55.8 48.6 ; 
      RECT 55.264 44.226 55.368 48.6 ; 
      RECT 54.832 44.226 54.936 48.6 ; 
      RECT 54.4 44.226 54.504 48.6 ; 
      RECT 53.968 44.226 54.072 48.6 ; 
      RECT 53.536 44.226 53.64 48.6 ; 
      RECT 53.104 44.226 53.208 48.6 ; 
      RECT 52.672 44.226 52.776 48.6 ; 
      RECT 52.24 44.226 52.344 48.6 ; 
      RECT 51.808 44.226 51.912 48.6 ; 
      RECT 51.376 44.226 51.48 48.6 ; 
      RECT 50.944 44.226 51.048 48.6 ; 
      RECT 50.512 44.226 50.616 48.6 ; 
      RECT 50.08 44.226 50.184 48.6 ; 
      RECT 49.648 44.226 49.752 48.6 ; 
      RECT 49.216 44.226 49.32 48.6 ; 
      RECT 48.784 44.226 48.888 48.6 ; 
      RECT 48.352 44.226 48.456 48.6 ; 
      RECT 47.92 44.226 48.024 48.6 ; 
      RECT 47.488 44.226 47.592 48.6 ; 
      RECT 47.056 44.226 47.16 48.6 ; 
      RECT 46.624 44.226 46.728 48.6 ; 
      RECT 46.192 44.226 46.296 48.6 ; 
      RECT 45.76 44.226 45.864 48.6 ; 
      RECT 45.328 44.226 45.432 48.6 ; 
      RECT 44.896 44.226 45 48.6 ; 
      RECT 44.464 44.226 44.568 48.6 ; 
      RECT 44.032 44.226 44.136 48.6 ; 
      RECT 43.6 44.226 43.704 48.6 ; 
      RECT 43.168 44.226 43.272 48.6 ; 
      RECT 42.736 44.226 42.84 48.6 ; 
      RECT 42.304 44.226 42.408 48.6 ; 
      RECT 41.872 44.226 41.976 48.6 ; 
      RECT 41.44 44.226 41.544 48.6 ; 
      RECT 41.008 44.226 41.112 48.6 ; 
      RECT 40.576 44.226 40.68 48.6 ; 
      RECT 40.144 44.226 40.248 48.6 ; 
      RECT 39.712 44.226 39.816 48.6 ; 
      RECT 39.28 44.226 39.384 48.6 ; 
      RECT 38.848 44.226 38.952 48.6 ; 
      RECT 38.416 44.226 38.52 48.6 ; 
      RECT 37.984 44.226 38.088 48.6 ; 
      RECT 37.552 44.226 37.656 48.6 ; 
      RECT 36.7 44.226 37.008 48.6 ; 
      RECT 29.128 44.226 29.436 48.6 ; 
      RECT 28.48 44.226 28.584 48.6 ; 
      RECT 28.048 44.226 28.152 48.6 ; 
      RECT 27.616 44.226 27.72 48.6 ; 
      RECT 27.184 44.226 27.288 48.6 ; 
      RECT 26.752 44.226 26.856 48.6 ; 
      RECT 26.32 44.226 26.424 48.6 ; 
      RECT 25.888 44.226 25.992 48.6 ; 
      RECT 25.456 44.226 25.56 48.6 ; 
      RECT 25.024 44.226 25.128 48.6 ; 
      RECT 24.592 44.226 24.696 48.6 ; 
      RECT 24.16 44.226 24.264 48.6 ; 
      RECT 23.728 44.226 23.832 48.6 ; 
      RECT 23.296 44.226 23.4 48.6 ; 
      RECT 22.864 44.226 22.968 48.6 ; 
      RECT 22.432 44.226 22.536 48.6 ; 
      RECT 22 44.226 22.104 48.6 ; 
      RECT 21.568 44.226 21.672 48.6 ; 
      RECT 21.136 44.226 21.24 48.6 ; 
      RECT 20.704 44.226 20.808 48.6 ; 
      RECT 20.272 44.226 20.376 48.6 ; 
      RECT 19.84 44.226 19.944 48.6 ; 
      RECT 19.408 44.226 19.512 48.6 ; 
      RECT 18.976 44.226 19.08 48.6 ; 
      RECT 18.544 44.226 18.648 48.6 ; 
      RECT 18.112 44.226 18.216 48.6 ; 
      RECT 17.68 44.226 17.784 48.6 ; 
      RECT 17.248 44.226 17.352 48.6 ; 
      RECT 16.816 44.226 16.92 48.6 ; 
      RECT 16.384 44.226 16.488 48.6 ; 
      RECT 15.952 44.226 16.056 48.6 ; 
      RECT 15.52 44.226 15.624 48.6 ; 
      RECT 15.088 44.226 15.192 48.6 ; 
      RECT 14.656 44.226 14.76 48.6 ; 
      RECT 14.224 44.226 14.328 48.6 ; 
      RECT 13.792 44.226 13.896 48.6 ; 
      RECT 13.36 44.226 13.464 48.6 ; 
      RECT 12.928 44.226 13.032 48.6 ; 
      RECT 12.496 44.226 12.6 48.6 ; 
      RECT 12.064 44.226 12.168 48.6 ; 
      RECT 11.632 44.226 11.736 48.6 ; 
      RECT 11.2 44.226 11.304 48.6 ; 
      RECT 10.768 44.226 10.872 48.6 ; 
      RECT 10.336 44.226 10.44 48.6 ; 
      RECT 9.904 44.226 10.008 48.6 ; 
      RECT 9.472 44.226 9.576 48.6 ; 
      RECT 9.04 44.226 9.144 48.6 ; 
      RECT 8.608 44.226 8.712 48.6 ; 
      RECT 8.176 44.226 8.28 48.6 ; 
      RECT 7.744 44.226 7.848 48.6 ; 
      RECT 7.312 44.226 7.416 48.6 ; 
      RECT 6.88 44.226 6.984 48.6 ; 
      RECT 6.448 44.226 6.552 48.6 ; 
      RECT 6.016 44.226 6.12 48.6 ; 
      RECT 5.584 44.226 5.688 48.6 ; 
      RECT 5.152 44.226 5.256 48.6 ; 
      RECT 4.72 44.226 4.824 48.6 ; 
      RECT 4.288 44.226 4.392 48.6 ; 
      RECT 3.856 44.226 3.96 48.6 ; 
      RECT 3.424 44.226 3.528 48.6 ; 
      RECT 2.992 44.226 3.096 48.6 ; 
      RECT 2.56 44.226 2.664 48.6 ; 
      RECT 2.128 44.226 2.232 48.6 ; 
      RECT 1.696 44.226 1.8 48.6 ; 
      RECT 1.264 44.226 1.368 48.6 ; 
      RECT 0.832 44.226 0.936 48.6 ; 
      RECT 0.02 44.226 0.36 48.6 ; 
      RECT 34.564 48.546 35.076 52.92 ; 
      RECT 34.508 51.208 35.076 52.498 ; 
      RECT 33.916 50.116 34.164 52.92 ; 
      RECT 33.86 51.354 34.164 51.968 ; 
      RECT 33.916 48.546 34.02 52.92 ; 
      RECT 33.916 49.03 34.076 49.988 ; 
      RECT 33.916 48.546 34.164 48.902 ; 
      RECT 32.728 50.348 33.552 52.92 ; 
      RECT 33.448 48.546 33.552 52.92 ; 
      RECT 32.728 51.456 33.608 52.488 ; 
      RECT 32.728 48.546 33.12 52.92 ; 
      RECT 31.06 48.546 31.392 52.92 ; 
      RECT 31.06 48.9 31.448 52.642 ; 
      RECT 65.776 48.546 66.116 52.92 ; 
      RECT 65.2 48.546 65.304 52.92 ; 
      RECT 64.768 48.546 64.872 52.92 ; 
      RECT 64.336 48.546 64.44 52.92 ; 
      RECT 63.904 48.546 64.008 52.92 ; 
      RECT 63.472 48.546 63.576 52.92 ; 
      RECT 63.04 48.546 63.144 52.92 ; 
      RECT 62.608 48.546 62.712 52.92 ; 
      RECT 62.176 48.546 62.28 52.92 ; 
      RECT 61.744 48.546 61.848 52.92 ; 
      RECT 61.312 48.546 61.416 52.92 ; 
      RECT 60.88 48.546 60.984 52.92 ; 
      RECT 60.448 48.546 60.552 52.92 ; 
      RECT 60.016 48.546 60.12 52.92 ; 
      RECT 59.584 48.546 59.688 52.92 ; 
      RECT 59.152 48.546 59.256 52.92 ; 
      RECT 58.72 48.546 58.824 52.92 ; 
      RECT 58.288 48.546 58.392 52.92 ; 
      RECT 57.856 48.546 57.96 52.92 ; 
      RECT 57.424 48.546 57.528 52.92 ; 
      RECT 56.992 48.546 57.096 52.92 ; 
      RECT 56.56 48.546 56.664 52.92 ; 
      RECT 56.128 48.546 56.232 52.92 ; 
      RECT 55.696 48.546 55.8 52.92 ; 
      RECT 55.264 48.546 55.368 52.92 ; 
      RECT 54.832 48.546 54.936 52.92 ; 
      RECT 54.4 48.546 54.504 52.92 ; 
      RECT 53.968 48.546 54.072 52.92 ; 
      RECT 53.536 48.546 53.64 52.92 ; 
      RECT 53.104 48.546 53.208 52.92 ; 
      RECT 52.672 48.546 52.776 52.92 ; 
      RECT 52.24 48.546 52.344 52.92 ; 
      RECT 51.808 48.546 51.912 52.92 ; 
      RECT 51.376 48.546 51.48 52.92 ; 
      RECT 50.944 48.546 51.048 52.92 ; 
      RECT 50.512 48.546 50.616 52.92 ; 
      RECT 50.08 48.546 50.184 52.92 ; 
      RECT 49.648 48.546 49.752 52.92 ; 
      RECT 49.216 48.546 49.32 52.92 ; 
      RECT 48.784 48.546 48.888 52.92 ; 
      RECT 48.352 48.546 48.456 52.92 ; 
      RECT 47.92 48.546 48.024 52.92 ; 
      RECT 47.488 48.546 47.592 52.92 ; 
      RECT 47.056 48.546 47.16 52.92 ; 
      RECT 46.624 48.546 46.728 52.92 ; 
      RECT 46.192 48.546 46.296 52.92 ; 
      RECT 45.76 48.546 45.864 52.92 ; 
      RECT 45.328 48.546 45.432 52.92 ; 
      RECT 44.896 48.546 45 52.92 ; 
      RECT 44.464 48.546 44.568 52.92 ; 
      RECT 44.032 48.546 44.136 52.92 ; 
      RECT 43.6 48.546 43.704 52.92 ; 
      RECT 43.168 48.546 43.272 52.92 ; 
      RECT 42.736 48.546 42.84 52.92 ; 
      RECT 42.304 48.546 42.408 52.92 ; 
      RECT 41.872 48.546 41.976 52.92 ; 
      RECT 41.44 48.546 41.544 52.92 ; 
      RECT 41.008 48.546 41.112 52.92 ; 
      RECT 40.576 48.546 40.68 52.92 ; 
      RECT 40.144 48.546 40.248 52.92 ; 
      RECT 39.712 48.546 39.816 52.92 ; 
      RECT 39.28 48.546 39.384 52.92 ; 
      RECT 38.848 48.546 38.952 52.92 ; 
      RECT 38.416 48.546 38.52 52.92 ; 
      RECT 37.984 48.546 38.088 52.92 ; 
      RECT 37.552 48.546 37.656 52.92 ; 
      RECT 36.7 48.546 37.008 52.92 ; 
      RECT 29.128 48.546 29.436 52.92 ; 
      RECT 28.48 48.546 28.584 52.92 ; 
      RECT 28.048 48.546 28.152 52.92 ; 
      RECT 27.616 48.546 27.72 52.92 ; 
      RECT 27.184 48.546 27.288 52.92 ; 
      RECT 26.752 48.546 26.856 52.92 ; 
      RECT 26.32 48.546 26.424 52.92 ; 
      RECT 25.888 48.546 25.992 52.92 ; 
      RECT 25.456 48.546 25.56 52.92 ; 
      RECT 25.024 48.546 25.128 52.92 ; 
      RECT 24.592 48.546 24.696 52.92 ; 
      RECT 24.16 48.546 24.264 52.92 ; 
      RECT 23.728 48.546 23.832 52.92 ; 
      RECT 23.296 48.546 23.4 52.92 ; 
      RECT 22.864 48.546 22.968 52.92 ; 
      RECT 22.432 48.546 22.536 52.92 ; 
      RECT 22 48.546 22.104 52.92 ; 
      RECT 21.568 48.546 21.672 52.92 ; 
      RECT 21.136 48.546 21.24 52.92 ; 
      RECT 20.704 48.546 20.808 52.92 ; 
      RECT 20.272 48.546 20.376 52.92 ; 
      RECT 19.84 48.546 19.944 52.92 ; 
      RECT 19.408 48.546 19.512 52.92 ; 
      RECT 18.976 48.546 19.08 52.92 ; 
      RECT 18.544 48.546 18.648 52.92 ; 
      RECT 18.112 48.546 18.216 52.92 ; 
      RECT 17.68 48.546 17.784 52.92 ; 
      RECT 17.248 48.546 17.352 52.92 ; 
      RECT 16.816 48.546 16.92 52.92 ; 
      RECT 16.384 48.546 16.488 52.92 ; 
      RECT 15.952 48.546 16.056 52.92 ; 
      RECT 15.52 48.546 15.624 52.92 ; 
      RECT 15.088 48.546 15.192 52.92 ; 
      RECT 14.656 48.546 14.76 52.92 ; 
      RECT 14.224 48.546 14.328 52.92 ; 
      RECT 13.792 48.546 13.896 52.92 ; 
      RECT 13.36 48.546 13.464 52.92 ; 
      RECT 12.928 48.546 13.032 52.92 ; 
      RECT 12.496 48.546 12.6 52.92 ; 
      RECT 12.064 48.546 12.168 52.92 ; 
      RECT 11.632 48.546 11.736 52.92 ; 
      RECT 11.2 48.546 11.304 52.92 ; 
      RECT 10.768 48.546 10.872 52.92 ; 
      RECT 10.336 48.546 10.44 52.92 ; 
      RECT 9.904 48.546 10.008 52.92 ; 
      RECT 9.472 48.546 9.576 52.92 ; 
      RECT 9.04 48.546 9.144 52.92 ; 
      RECT 8.608 48.546 8.712 52.92 ; 
      RECT 8.176 48.546 8.28 52.92 ; 
      RECT 7.744 48.546 7.848 52.92 ; 
      RECT 7.312 48.546 7.416 52.92 ; 
      RECT 6.88 48.546 6.984 52.92 ; 
      RECT 6.448 48.546 6.552 52.92 ; 
      RECT 6.016 48.546 6.12 52.92 ; 
      RECT 5.584 48.546 5.688 52.92 ; 
      RECT 5.152 48.546 5.256 52.92 ; 
      RECT 4.72 48.546 4.824 52.92 ; 
      RECT 4.288 48.546 4.392 52.92 ; 
      RECT 3.856 48.546 3.96 52.92 ; 
      RECT 3.424 48.546 3.528 52.92 ; 
      RECT 2.992 48.546 3.096 52.92 ; 
      RECT 2.56 48.546 2.664 52.92 ; 
      RECT 2.128 48.546 2.232 52.92 ; 
      RECT 1.696 48.546 1.8 52.92 ; 
      RECT 1.264 48.546 1.368 52.92 ; 
      RECT 0.832 48.546 0.936 52.92 ; 
      RECT 0.02 48.546 0.36 52.92 ; 
      RECT 34.564 52.866 35.076 57.24 ; 
      RECT 34.508 55.528 35.076 56.818 ; 
      RECT 33.916 54.436 34.164 57.24 ; 
      RECT 33.86 55.674 34.164 56.288 ; 
      RECT 33.916 52.866 34.02 57.24 ; 
      RECT 33.916 53.35 34.076 54.308 ; 
      RECT 33.916 52.866 34.164 53.222 ; 
      RECT 32.728 54.668 33.552 57.24 ; 
      RECT 33.448 52.866 33.552 57.24 ; 
      RECT 32.728 55.776 33.608 56.808 ; 
      RECT 32.728 52.866 33.12 57.24 ; 
      RECT 31.06 52.866 31.392 57.24 ; 
      RECT 31.06 53.22 31.448 56.962 ; 
      RECT 65.776 52.866 66.116 57.24 ; 
      RECT 65.2 52.866 65.304 57.24 ; 
      RECT 64.768 52.866 64.872 57.24 ; 
      RECT 64.336 52.866 64.44 57.24 ; 
      RECT 63.904 52.866 64.008 57.24 ; 
      RECT 63.472 52.866 63.576 57.24 ; 
      RECT 63.04 52.866 63.144 57.24 ; 
      RECT 62.608 52.866 62.712 57.24 ; 
      RECT 62.176 52.866 62.28 57.24 ; 
      RECT 61.744 52.866 61.848 57.24 ; 
      RECT 61.312 52.866 61.416 57.24 ; 
      RECT 60.88 52.866 60.984 57.24 ; 
      RECT 60.448 52.866 60.552 57.24 ; 
      RECT 60.016 52.866 60.12 57.24 ; 
      RECT 59.584 52.866 59.688 57.24 ; 
      RECT 59.152 52.866 59.256 57.24 ; 
      RECT 58.72 52.866 58.824 57.24 ; 
      RECT 58.288 52.866 58.392 57.24 ; 
      RECT 57.856 52.866 57.96 57.24 ; 
      RECT 57.424 52.866 57.528 57.24 ; 
      RECT 56.992 52.866 57.096 57.24 ; 
      RECT 56.56 52.866 56.664 57.24 ; 
      RECT 56.128 52.866 56.232 57.24 ; 
      RECT 55.696 52.866 55.8 57.24 ; 
      RECT 55.264 52.866 55.368 57.24 ; 
      RECT 54.832 52.866 54.936 57.24 ; 
      RECT 54.4 52.866 54.504 57.24 ; 
      RECT 53.968 52.866 54.072 57.24 ; 
      RECT 53.536 52.866 53.64 57.24 ; 
      RECT 53.104 52.866 53.208 57.24 ; 
      RECT 52.672 52.866 52.776 57.24 ; 
      RECT 52.24 52.866 52.344 57.24 ; 
      RECT 51.808 52.866 51.912 57.24 ; 
      RECT 51.376 52.866 51.48 57.24 ; 
      RECT 50.944 52.866 51.048 57.24 ; 
      RECT 50.512 52.866 50.616 57.24 ; 
      RECT 50.08 52.866 50.184 57.24 ; 
      RECT 49.648 52.866 49.752 57.24 ; 
      RECT 49.216 52.866 49.32 57.24 ; 
      RECT 48.784 52.866 48.888 57.24 ; 
      RECT 48.352 52.866 48.456 57.24 ; 
      RECT 47.92 52.866 48.024 57.24 ; 
      RECT 47.488 52.866 47.592 57.24 ; 
      RECT 47.056 52.866 47.16 57.24 ; 
      RECT 46.624 52.866 46.728 57.24 ; 
      RECT 46.192 52.866 46.296 57.24 ; 
      RECT 45.76 52.866 45.864 57.24 ; 
      RECT 45.328 52.866 45.432 57.24 ; 
      RECT 44.896 52.866 45 57.24 ; 
      RECT 44.464 52.866 44.568 57.24 ; 
      RECT 44.032 52.866 44.136 57.24 ; 
      RECT 43.6 52.866 43.704 57.24 ; 
      RECT 43.168 52.866 43.272 57.24 ; 
      RECT 42.736 52.866 42.84 57.24 ; 
      RECT 42.304 52.866 42.408 57.24 ; 
      RECT 41.872 52.866 41.976 57.24 ; 
      RECT 41.44 52.866 41.544 57.24 ; 
      RECT 41.008 52.866 41.112 57.24 ; 
      RECT 40.576 52.866 40.68 57.24 ; 
      RECT 40.144 52.866 40.248 57.24 ; 
      RECT 39.712 52.866 39.816 57.24 ; 
      RECT 39.28 52.866 39.384 57.24 ; 
      RECT 38.848 52.866 38.952 57.24 ; 
      RECT 38.416 52.866 38.52 57.24 ; 
      RECT 37.984 52.866 38.088 57.24 ; 
      RECT 37.552 52.866 37.656 57.24 ; 
      RECT 36.7 52.866 37.008 57.24 ; 
      RECT 29.128 52.866 29.436 57.24 ; 
      RECT 28.48 52.866 28.584 57.24 ; 
      RECT 28.048 52.866 28.152 57.24 ; 
      RECT 27.616 52.866 27.72 57.24 ; 
      RECT 27.184 52.866 27.288 57.24 ; 
      RECT 26.752 52.866 26.856 57.24 ; 
      RECT 26.32 52.866 26.424 57.24 ; 
      RECT 25.888 52.866 25.992 57.24 ; 
      RECT 25.456 52.866 25.56 57.24 ; 
      RECT 25.024 52.866 25.128 57.24 ; 
      RECT 24.592 52.866 24.696 57.24 ; 
      RECT 24.16 52.866 24.264 57.24 ; 
      RECT 23.728 52.866 23.832 57.24 ; 
      RECT 23.296 52.866 23.4 57.24 ; 
      RECT 22.864 52.866 22.968 57.24 ; 
      RECT 22.432 52.866 22.536 57.24 ; 
      RECT 22 52.866 22.104 57.24 ; 
      RECT 21.568 52.866 21.672 57.24 ; 
      RECT 21.136 52.866 21.24 57.24 ; 
      RECT 20.704 52.866 20.808 57.24 ; 
      RECT 20.272 52.866 20.376 57.24 ; 
      RECT 19.84 52.866 19.944 57.24 ; 
      RECT 19.408 52.866 19.512 57.24 ; 
      RECT 18.976 52.866 19.08 57.24 ; 
      RECT 18.544 52.866 18.648 57.24 ; 
      RECT 18.112 52.866 18.216 57.24 ; 
      RECT 17.68 52.866 17.784 57.24 ; 
      RECT 17.248 52.866 17.352 57.24 ; 
      RECT 16.816 52.866 16.92 57.24 ; 
      RECT 16.384 52.866 16.488 57.24 ; 
      RECT 15.952 52.866 16.056 57.24 ; 
      RECT 15.52 52.866 15.624 57.24 ; 
      RECT 15.088 52.866 15.192 57.24 ; 
      RECT 14.656 52.866 14.76 57.24 ; 
      RECT 14.224 52.866 14.328 57.24 ; 
      RECT 13.792 52.866 13.896 57.24 ; 
      RECT 13.36 52.866 13.464 57.24 ; 
      RECT 12.928 52.866 13.032 57.24 ; 
      RECT 12.496 52.866 12.6 57.24 ; 
      RECT 12.064 52.866 12.168 57.24 ; 
      RECT 11.632 52.866 11.736 57.24 ; 
      RECT 11.2 52.866 11.304 57.24 ; 
      RECT 10.768 52.866 10.872 57.24 ; 
      RECT 10.336 52.866 10.44 57.24 ; 
      RECT 9.904 52.866 10.008 57.24 ; 
      RECT 9.472 52.866 9.576 57.24 ; 
      RECT 9.04 52.866 9.144 57.24 ; 
      RECT 8.608 52.866 8.712 57.24 ; 
      RECT 8.176 52.866 8.28 57.24 ; 
      RECT 7.744 52.866 7.848 57.24 ; 
      RECT 7.312 52.866 7.416 57.24 ; 
      RECT 6.88 52.866 6.984 57.24 ; 
      RECT 6.448 52.866 6.552 57.24 ; 
      RECT 6.016 52.866 6.12 57.24 ; 
      RECT 5.584 52.866 5.688 57.24 ; 
      RECT 5.152 52.866 5.256 57.24 ; 
      RECT 4.72 52.866 4.824 57.24 ; 
      RECT 4.288 52.866 4.392 57.24 ; 
      RECT 3.856 52.866 3.96 57.24 ; 
      RECT 3.424 52.866 3.528 57.24 ; 
      RECT 2.992 52.866 3.096 57.24 ; 
      RECT 2.56 52.866 2.664 57.24 ; 
      RECT 2.128 52.866 2.232 57.24 ; 
      RECT 1.696 52.866 1.8 57.24 ; 
      RECT 1.264 52.866 1.368 57.24 ; 
      RECT 0.832 52.866 0.936 57.24 ; 
      RECT 0.02 52.866 0.36 57.24 ; 
      RECT 34.564 57.186 35.076 61.56 ; 
      RECT 34.508 59.848 35.076 61.138 ; 
      RECT 33.916 58.756 34.164 61.56 ; 
      RECT 33.86 59.994 34.164 60.608 ; 
      RECT 33.916 57.186 34.02 61.56 ; 
      RECT 33.916 57.67 34.076 58.628 ; 
      RECT 33.916 57.186 34.164 57.542 ; 
      RECT 32.728 58.988 33.552 61.56 ; 
      RECT 33.448 57.186 33.552 61.56 ; 
      RECT 32.728 60.096 33.608 61.128 ; 
      RECT 32.728 57.186 33.12 61.56 ; 
      RECT 31.06 57.186 31.392 61.56 ; 
      RECT 31.06 57.54 31.448 61.282 ; 
      RECT 65.776 57.186 66.116 61.56 ; 
      RECT 65.2 57.186 65.304 61.56 ; 
      RECT 64.768 57.186 64.872 61.56 ; 
      RECT 64.336 57.186 64.44 61.56 ; 
      RECT 63.904 57.186 64.008 61.56 ; 
      RECT 63.472 57.186 63.576 61.56 ; 
      RECT 63.04 57.186 63.144 61.56 ; 
      RECT 62.608 57.186 62.712 61.56 ; 
      RECT 62.176 57.186 62.28 61.56 ; 
      RECT 61.744 57.186 61.848 61.56 ; 
      RECT 61.312 57.186 61.416 61.56 ; 
      RECT 60.88 57.186 60.984 61.56 ; 
      RECT 60.448 57.186 60.552 61.56 ; 
      RECT 60.016 57.186 60.12 61.56 ; 
      RECT 59.584 57.186 59.688 61.56 ; 
      RECT 59.152 57.186 59.256 61.56 ; 
      RECT 58.72 57.186 58.824 61.56 ; 
      RECT 58.288 57.186 58.392 61.56 ; 
      RECT 57.856 57.186 57.96 61.56 ; 
      RECT 57.424 57.186 57.528 61.56 ; 
      RECT 56.992 57.186 57.096 61.56 ; 
      RECT 56.56 57.186 56.664 61.56 ; 
      RECT 56.128 57.186 56.232 61.56 ; 
      RECT 55.696 57.186 55.8 61.56 ; 
      RECT 55.264 57.186 55.368 61.56 ; 
      RECT 54.832 57.186 54.936 61.56 ; 
      RECT 54.4 57.186 54.504 61.56 ; 
      RECT 53.968 57.186 54.072 61.56 ; 
      RECT 53.536 57.186 53.64 61.56 ; 
      RECT 53.104 57.186 53.208 61.56 ; 
      RECT 52.672 57.186 52.776 61.56 ; 
      RECT 52.24 57.186 52.344 61.56 ; 
      RECT 51.808 57.186 51.912 61.56 ; 
      RECT 51.376 57.186 51.48 61.56 ; 
      RECT 50.944 57.186 51.048 61.56 ; 
      RECT 50.512 57.186 50.616 61.56 ; 
      RECT 50.08 57.186 50.184 61.56 ; 
      RECT 49.648 57.186 49.752 61.56 ; 
      RECT 49.216 57.186 49.32 61.56 ; 
      RECT 48.784 57.186 48.888 61.56 ; 
      RECT 48.352 57.186 48.456 61.56 ; 
      RECT 47.92 57.186 48.024 61.56 ; 
      RECT 47.488 57.186 47.592 61.56 ; 
      RECT 47.056 57.186 47.16 61.56 ; 
      RECT 46.624 57.186 46.728 61.56 ; 
      RECT 46.192 57.186 46.296 61.56 ; 
      RECT 45.76 57.186 45.864 61.56 ; 
      RECT 45.328 57.186 45.432 61.56 ; 
      RECT 44.896 57.186 45 61.56 ; 
      RECT 44.464 57.186 44.568 61.56 ; 
      RECT 44.032 57.186 44.136 61.56 ; 
      RECT 43.6 57.186 43.704 61.56 ; 
      RECT 43.168 57.186 43.272 61.56 ; 
      RECT 42.736 57.186 42.84 61.56 ; 
      RECT 42.304 57.186 42.408 61.56 ; 
      RECT 41.872 57.186 41.976 61.56 ; 
      RECT 41.44 57.186 41.544 61.56 ; 
      RECT 41.008 57.186 41.112 61.56 ; 
      RECT 40.576 57.186 40.68 61.56 ; 
      RECT 40.144 57.186 40.248 61.56 ; 
      RECT 39.712 57.186 39.816 61.56 ; 
      RECT 39.28 57.186 39.384 61.56 ; 
      RECT 38.848 57.186 38.952 61.56 ; 
      RECT 38.416 57.186 38.52 61.56 ; 
      RECT 37.984 57.186 38.088 61.56 ; 
      RECT 37.552 57.186 37.656 61.56 ; 
      RECT 36.7 57.186 37.008 61.56 ; 
      RECT 29.128 57.186 29.436 61.56 ; 
      RECT 28.48 57.186 28.584 61.56 ; 
      RECT 28.048 57.186 28.152 61.56 ; 
      RECT 27.616 57.186 27.72 61.56 ; 
      RECT 27.184 57.186 27.288 61.56 ; 
      RECT 26.752 57.186 26.856 61.56 ; 
      RECT 26.32 57.186 26.424 61.56 ; 
      RECT 25.888 57.186 25.992 61.56 ; 
      RECT 25.456 57.186 25.56 61.56 ; 
      RECT 25.024 57.186 25.128 61.56 ; 
      RECT 24.592 57.186 24.696 61.56 ; 
      RECT 24.16 57.186 24.264 61.56 ; 
      RECT 23.728 57.186 23.832 61.56 ; 
      RECT 23.296 57.186 23.4 61.56 ; 
      RECT 22.864 57.186 22.968 61.56 ; 
      RECT 22.432 57.186 22.536 61.56 ; 
      RECT 22 57.186 22.104 61.56 ; 
      RECT 21.568 57.186 21.672 61.56 ; 
      RECT 21.136 57.186 21.24 61.56 ; 
      RECT 20.704 57.186 20.808 61.56 ; 
      RECT 20.272 57.186 20.376 61.56 ; 
      RECT 19.84 57.186 19.944 61.56 ; 
      RECT 19.408 57.186 19.512 61.56 ; 
      RECT 18.976 57.186 19.08 61.56 ; 
      RECT 18.544 57.186 18.648 61.56 ; 
      RECT 18.112 57.186 18.216 61.56 ; 
      RECT 17.68 57.186 17.784 61.56 ; 
      RECT 17.248 57.186 17.352 61.56 ; 
      RECT 16.816 57.186 16.92 61.56 ; 
      RECT 16.384 57.186 16.488 61.56 ; 
      RECT 15.952 57.186 16.056 61.56 ; 
      RECT 15.52 57.186 15.624 61.56 ; 
      RECT 15.088 57.186 15.192 61.56 ; 
      RECT 14.656 57.186 14.76 61.56 ; 
      RECT 14.224 57.186 14.328 61.56 ; 
      RECT 13.792 57.186 13.896 61.56 ; 
      RECT 13.36 57.186 13.464 61.56 ; 
      RECT 12.928 57.186 13.032 61.56 ; 
      RECT 12.496 57.186 12.6 61.56 ; 
      RECT 12.064 57.186 12.168 61.56 ; 
      RECT 11.632 57.186 11.736 61.56 ; 
      RECT 11.2 57.186 11.304 61.56 ; 
      RECT 10.768 57.186 10.872 61.56 ; 
      RECT 10.336 57.186 10.44 61.56 ; 
      RECT 9.904 57.186 10.008 61.56 ; 
      RECT 9.472 57.186 9.576 61.56 ; 
      RECT 9.04 57.186 9.144 61.56 ; 
      RECT 8.608 57.186 8.712 61.56 ; 
      RECT 8.176 57.186 8.28 61.56 ; 
      RECT 7.744 57.186 7.848 61.56 ; 
      RECT 7.312 57.186 7.416 61.56 ; 
      RECT 6.88 57.186 6.984 61.56 ; 
      RECT 6.448 57.186 6.552 61.56 ; 
      RECT 6.016 57.186 6.12 61.56 ; 
      RECT 5.584 57.186 5.688 61.56 ; 
      RECT 5.152 57.186 5.256 61.56 ; 
      RECT 4.72 57.186 4.824 61.56 ; 
      RECT 4.288 57.186 4.392 61.56 ; 
      RECT 3.856 57.186 3.96 61.56 ; 
      RECT 3.424 57.186 3.528 61.56 ; 
      RECT 2.992 57.186 3.096 61.56 ; 
      RECT 2.56 57.186 2.664 61.56 ; 
      RECT 2.128 57.186 2.232 61.56 ; 
      RECT 1.696 57.186 1.8 61.56 ; 
      RECT 1.264 57.186 1.368 61.56 ; 
      RECT 0.832 57.186 0.936 61.56 ; 
      RECT 0.02 57.186 0.36 61.56 ; 
      RECT 34.564 61.506 35.076 65.88 ; 
      RECT 34.508 64.168 35.076 65.458 ; 
      RECT 33.916 63.076 34.164 65.88 ; 
      RECT 33.86 64.314 34.164 64.928 ; 
      RECT 33.916 61.506 34.02 65.88 ; 
      RECT 33.916 61.99 34.076 62.948 ; 
      RECT 33.916 61.506 34.164 61.862 ; 
      RECT 32.728 63.308 33.552 65.88 ; 
      RECT 33.448 61.506 33.552 65.88 ; 
      RECT 32.728 64.416 33.608 65.448 ; 
      RECT 32.728 61.506 33.12 65.88 ; 
      RECT 31.06 61.506 31.392 65.88 ; 
      RECT 31.06 61.86 31.448 65.602 ; 
      RECT 65.776 61.506 66.116 65.88 ; 
      RECT 65.2 61.506 65.304 65.88 ; 
      RECT 64.768 61.506 64.872 65.88 ; 
      RECT 64.336 61.506 64.44 65.88 ; 
      RECT 63.904 61.506 64.008 65.88 ; 
      RECT 63.472 61.506 63.576 65.88 ; 
      RECT 63.04 61.506 63.144 65.88 ; 
      RECT 62.608 61.506 62.712 65.88 ; 
      RECT 62.176 61.506 62.28 65.88 ; 
      RECT 61.744 61.506 61.848 65.88 ; 
      RECT 61.312 61.506 61.416 65.88 ; 
      RECT 60.88 61.506 60.984 65.88 ; 
      RECT 60.448 61.506 60.552 65.88 ; 
      RECT 60.016 61.506 60.12 65.88 ; 
      RECT 59.584 61.506 59.688 65.88 ; 
      RECT 59.152 61.506 59.256 65.88 ; 
      RECT 58.72 61.506 58.824 65.88 ; 
      RECT 58.288 61.506 58.392 65.88 ; 
      RECT 57.856 61.506 57.96 65.88 ; 
      RECT 57.424 61.506 57.528 65.88 ; 
      RECT 56.992 61.506 57.096 65.88 ; 
      RECT 56.56 61.506 56.664 65.88 ; 
      RECT 56.128 61.506 56.232 65.88 ; 
      RECT 55.696 61.506 55.8 65.88 ; 
      RECT 55.264 61.506 55.368 65.88 ; 
      RECT 54.832 61.506 54.936 65.88 ; 
      RECT 54.4 61.506 54.504 65.88 ; 
      RECT 53.968 61.506 54.072 65.88 ; 
      RECT 53.536 61.506 53.64 65.88 ; 
      RECT 53.104 61.506 53.208 65.88 ; 
      RECT 52.672 61.506 52.776 65.88 ; 
      RECT 52.24 61.506 52.344 65.88 ; 
      RECT 51.808 61.506 51.912 65.88 ; 
      RECT 51.376 61.506 51.48 65.88 ; 
      RECT 50.944 61.506 51.048 65.88 ; 
      RECT 50.512 61.506 50.616 65.88 ; 
      RECT 50.08 61.506 50.184 65.88 ; 
      RECT 49.648 61.506 49.752 65.88 ; 
      RECT 49.216 61.506 49.32 65.88 ; 
      RECT 48.784 61.506 48.888 65.88 ; 
      RECT 48.352 61.506 48.456 65.88 ; 
      RECT 47.92 61.506 48.024 65.88 ; 
      RECT 47.488 61.506 47.592 65.88 ; 
      RECT 47.056 61.506 47.16 65.88 ; 
      RECT 46.624 61.506 46.728 65.88 ; 
      RECT 46.192 61.506 46.296 65.88 ; 
      RECT 45.76 61.506 45.864 65.88 ; 
      RECT 45.328 61.506 45.432 65.88 ; 
      RECT 44.896 61.506 45 65.88 ; 
      RECT 44.464 61.506 44.568 65.88 ; 
      RECT 44.032 61.506 44.136 65.88 ; 
      RECT 43.6 61.506 43.704 65.88 ; 
      RECT 43.168 61.506 43.272 65.88 ; 
      RECT 42.736 61.506 42.84 65.88 ; 
      RECT 42.304 61.506 42.408 65.88 ; 
      RECT 41.872 61.506 41.976 65.88 ; 
      RECT 41.44 61.506 41.544 65.88 ; 
      RECT 41.008 61.506 41.112 65.88 ; 
      RECT 40.576 61.506 40.68 65.88 ; 
      RECT 40.144 61.506 40.248 65.88 ; 
      RECT 39.712 61.506 39.816 65.88 ; 
      RECT 39.28 61.506 39.384 65.88 ; 
      RECT 38.848 61.506 38.952 65.88 ; 
      RECT 38.416 61.506 38.52 65.88 ; 
      RECT 37.984 61.506 38.088 65.88 ; 
      RECT 37.552 61.506 37.656 65.88 ; 
      RECT 36.7 61.506 37.008 65.88 ; 
      RECT 29.128 61.506 29.436 65.88 ; 
      RECT 28.48 61.506 28.584 65.88 ; 
      RECT 28.048 61.506 28.152 65.88 ; 
      RECT 27.616 61.506 27.72 65.88 ; 
      RECT 27.184 61.506 27.288 65.88 ; 
      RECT 26.752 61.506 26.856 65.88 ; 
      RECT 26.32 61.506 26.424 65.88 ; 
      RECT 25.888 61.506 25.992 65.88 ; 
      RECT 25.456 61.506 25.56 65.88 ; 
      RECT 25.024 61.506 25.128 65.88 ; 
      RECT 24.592 61.506 24.696 65.88 ; 
      RECT 24.16 61.506 24.264 65.88 ; 
      RECT 23.728 61.506 23.832 65.88 ; 
      RECT 23.296 61.506 23.4 65.88 ; 
      RECT 22.864 61.506 22.968 65.88 ; 
      RECT 22.432 61.506 22.536 65.88 ; 
      RECT 22 61.506 22.104 65.88 ; 
      RECT 21.568 61.506 21.672 65.88 ; 
      RECT 21.136 61.506 21.24 65.88 ; 
      RECT 20.704 61.506 20.808 65.88 ; 
      RECT 20.272 61.506 20.376 65.88 ; 
      RECT 19.84 61.506 19.944 65.88 ; 
      RECT 19.408 61.506 19.512 65.88 ; 
      RECT 18.976 61.506 19.08 65.88 ; 
      RECT 18.544 61.506 18.648 65.88 ; 
      RECT 18.112 61.506 18.216 65.88 ; 
      RECT 17.68 61.506 17.784 65.88 ; 
      RECT 17.248 61.506 17.352 65.88 ; 
      RECT 16.816 61.506 16.92 65.88 ; 
      RECT 16.384 61.506 16.488 65.88 ; 
      RECT 15.952 61.506 16.056 65.88 ; 
      RECT 15.52 61.506 15.624 65.88 ; 
      RECT 15.088 61.506 15.192 65.88 ; 
      RECT 14.656 61.506 14.76 65.88 ; 
      RECT 14.224 61.506 14.328 65.88 ; 
      RECT 13.792 61.506 13.896 65.88 ; 
      RECT 13.36 61.506 13.464 65.88 ; 
      RECT 12.928 61.506 13.032 65.88 ; 
      RECT 12.496 61.506 12.6 65.88 ; 
      RECT 12.064 61.506 12.168 65.88 ; 
      RECT 11.632 61.506 11.736 65.88 ; 
      RECT 11.2 61.506 11.304 65.88 ; 
      RECT 10.768 61.506 10.872 65.88 ; 
      RECT 10.336 61.506 10.44 65.88 ; 
      RECT 9.904 61.506 10.008 65.88 ; 
      RECT 9.472 61.506 9.576 65.88 ; 
      RECT 9.04 61.506 9.144 65.88 ; 
      RECT 8.608 61.506 8.712 65.88 ; 
      RECT 8.176 61.506 8.28 65.88 ; 
      RECT 7.744 61.506 7.848 65.88 ; 
      RECT 7.312 61.506 7.416 65.88 ; 
      RECT 6.88 61.506 6.984 65.88 ; 
      RECT 6.448 61.506 6.552 65.88 ; 
      RECT 6.016 61.506 6.12 65.88 ; 
      RECT 5.584 61.506 5.688 65.88 ; 
      RECT 5.152 61.506 5.256 65.88 ; 
      RECT 4.72 61.506 4.824 65.88 ; 
      RECT 4.288 61.506 4.392 65.88 ; 
      RECT 3.856 61.506 3.96 65.88 ; 
      RECT 3.424 61.506 3.528 65.88 ; 
      RECT 2.992 61.506 3.096 65.88 ; 
      RECT 2.56 61.506 2.664 65.88 ; 
      RECT 2.128 61.506 2.232 65.88 ; 
      RECT 1.696 61.506 1.8 65.88 ; 
      RECT 1.264 61.506 1.368 65.88 ; 
      RECT 0.832 61.506 0.936 65.88 ; 
      RECT 0.02 61.506 0.36 65.88 ; 
      RECT 34.564 65.826 35.076 70.2 ; 
      RECT 34.508 68.488 35.076 69.778 ; 
      RECT 33.916 67.396 34.164 70.2 ; 
      RECT 33.86 68.634 34.164 69.248 ; 
      RECT 33.916 65.826 34.02 70.2 ; 
      RECT 33.916 66.31 34.076 67.268 ; 
      RECT 33.916 65.826 34.164 66.182 ; 
      RECT 32.728 67.628 33.552 70.2 ; 
      RECT 33.448 65.826 33.552 70.2 ; 
      RECT 32.728 68.736 33.608 69.768 ; 
      RECT 32.728 65.826 33.12 70.2 ; 
      RECT 31.06 65.826 31.392 70.2 ; 
      RECT 31.06 66.18 31.448 69.922 ; 
      RECT 65.776 65.826 66.116 70.2 ; 
      RECT 65.2 65.826 65.304 70.2 ; 
      RECT 64.768 65.826 64.872 70.2 ; 
      RECT 64.336 65.826 64.44 70.2 ; 
      RECT 63.904 65.826 64.008 70.2 ; 
      RECT 63.472 65.826 63.576 70.2 ; 
      RECT 63.04 65.826 63.144 70.2 ; 
      RECT 62.608 65.826 62.712 70.2 ; 
      RECT 62.176 65.826 62.28 70.2 ; 
      RECT 61.744 65.826 61.848 70.2 ; 
      RECT 61.312 65.826 61.416 70.2 ; 
      RECT 60.88 65.826 60.984 70.2 ; 
      RECT 60.448 65.826 60.552 70.2 ; 
      RECT 60.016 65.826 60.12 70.2 ; 
      RECT 59.584 65.826 59.688 70.2 ; 
      RECT 59.152 65.826 59.256 70.2 ; 
      RECT 58.72 65.826 58.824 70.2 ; 
      RECT 58.288 65.826 58.392 70.2 ; 
      RECT 57.856 65.826 57.96 70.2 ; 
      RECT 57.424 65.826 57.528 70.2 ; 
      RECT 56.992 65.826 57.096 70.2 ; 
      RECT 56.56 65.826 56.664 70.2 ; 
      RECT 56.128 65.826 56.232 70.2 ; 
      RECT 55.696 65.826 55.8 70.2 ; 
      RECT 55.264 65.826 55.368 70.2 ; 
      RECT 54.832 65.826 54.936 70.2 ; 
      RECT 54.4 65.826 54.504 70.2 ; 
      RECT 53.968 65.826 54.072 70.2 ; 
      RECT 53.536 65.826 53.64 70.2 ; 
      RECT 53.104 65.826 53.208 70.2 ; 
      RECT 52.672 65.826 52.776 70.2 ; 
      RECT 52.24 65.826 52.344 70.2 ; 
      RECT 51.808 65.826 51.912 70.2 ; 
      RECT 51.376 65.826 51.48 70.2 ; 
      RECT 50.944 65.826 51.048 70.2 ; 
      RECT 50.512 65.826 50.616 70.2 ; 
      RECT 50.08 65.826 50.184 70.2 ; 
      RECT 49.648 65.826 49.752 70.2 ; 
      RECT 49.216 65.826 49.32 70.2 ; 
      RECT 48.784 65.826 48.888 70.2 ; 
      RECT 48.352 65.826 48.456 70.2 ; 
      RECT 47.92 65.826 48.024 70.2 ; 
      RECT 47.488 65.826 47.592 70.2 ; 
      RECT 47.056 65.826 47.16 70.2 ; 
      RECT 46.624 65.826 46.728 70.2 ; 
      RECT 46.192 65.826 46.296 70.2 ; 
      RECT 45.76 65.826 45.864 70.2 ; 
      RECT 45.328 65.826 45.432 70.2 ; 
      RECT 44.896 65.826 45 70.2 ; 
      RECT 44.464 65.826 44.568 70.2 ; 
      RECT 44.032 65.826 44.136 70.2 ; 
      RECT 43.6 65.826 43.704 70.2 ; 
      RECT 43.168 65.826 43.272 70.2 ; 
      RECT 42.736 65.826 42.84 70.2 ; 
      RECT 42.304 65.826 42.408 70.2 ; 
      RECT 41.872 65.826 41.976 70.2 ; 
      RECT 41.44 65.826 41.544 70.2 ; 
      RECT 41.008 65.826 41.112 70.2 ; 
      RECT 40.576 65.826 40.68 70.2 ; 
      RECT 40.144 65.826 40.248 70.2 ; 
      RECT 39.712 65.826 39.816 70.2 ; 
      RECT 39.28 65.826 39.384 70.2 ; 
      RECT 38.848 65.826 38.952 70.2 ; 
      RECT 38.416 65.826 38.52 70.2 ; 
      RECT 37.984 65.826 38.088 70.2 ; 
      RECT 37.552 65.826 37.656 70.2 ; 
      RECT 36.7 65.826 37.008 70.2 ; 
      RECT 29.128 65.826 29.436 70.2 ; 
      RECT 28.48 65.826 28.584 70.2 ; 
      RECT 28.048 65.826 28.152 70.2 ; 
      RECT 27.616 65.826 27.72 70.2 ; 
      RECT 27.184 65.826 27.288 70.2 ; 
      RECT 26.752 65.826 26.856 70.2 ; 
      RECT 26.32 65.826 26.424 70.2 ; 
      RECT 25.888 65.826 25.992 70.2 ; 
      RECT 25.456 65.826 25.56 70.2 ; 
      RECT 25.024 65.826 25.128 70.2 ; 
      RECT 24.592 65.826 24.696 70.2 ; 
      RECT 24.16 65.826 24.264 70.2 ; 
      RECT 23.728 65.826 23.832 70.2 ; 
      RECT 23.296 65.826 23.4 70.2 ; 
      RECT 22.864 65.826 22.968 70.2 ; 
      RECT 22.432 65.826 22.536 70.2 ; 
      RECT 22 65.826 22.104 70.2 ; 
      RECT 21.568 65.826 21.672 70.2 ; 
      RECT 21.136 65.826 21.24 70.2 ; 
      RECT 20.704 65.826 20.808 70.2 ; 
      RECT 20.272 65.826 20.376 70.2 ; 
      RECT 19.84 65.826 19.944 70.2 ; 
      RECT 19.408 65.826 19.512 70.2 ; 
      RECT 18.976 65.826 19.08 70.2 ; 
      RECT 18.544 65.826 18.648 70.2 ; 
      RECT 18.112 65.826 18.216 70.2 ; 
      RECT 17.68 65.826 17.784 70.2 ; 
      RECT 17.248 65.826 17.352 70.2 ; 
      RECT 16.816 65.826 16.92 70.2 ; 
      RECT 16.384 65.826 16.488 70.2 ; 
      RECT 15.952 65.826 16.056 70.2 ; 
      RECT 15.52 65.826 15.624 70.2 ; 
      RECT 15.088 65.826 15.192 70.2 ; 
      RECT 14.656 65.826 14.76 70.2 ; 
      RECT 14.224 65.826 14.328 70.2 ; 
      RECT 13.792 65.826 13.896 70.2 ; 
      RECT 13.36 65.826 13.464 70.2 ; 
      RECT 12.928 65.826 13.032 70.2 ; 
      RECT 12.496 65.826 12.6 70.2 ; 
      RECT 12.064 65.826 12.168 70.2 ; 
      RECT 11.632 65.826 11.736 70.2 ; 
      RECT 11.2 65.826 11.304 70.2 ; 
      RECT 10.768 65.826 10.872 70.2 ; 
      RECT 10.336 65.826 10.44 70.2 ; 
      RECT 9.904 65.826 10.008 70.2 ; 
      RECT 9.472 65.826 9.576 70.2 ; 
      RECT 9.04 65.826 9.144 70.2 ; 
      RECT 8.608 65.826 8.712 70.2 ; 
      RECT 8.176 65.826 8.28 70.2 ; 
      RECT 7.744 65.826 7.848 70.2 ; 
      RECT 7.312 65.826 7.416 70.2 ; 
      RECT 6.88 65.826 6.984 70.2 ; 
      RECT 6.448 65.826 6.552 70.2 ; 
      RECT 6.016 65.826 6.12 70.2 ; 
      RECT 5.584 65.826 5.688 70.2 ; 
      RECT 5.152 65.826 5.256 70.2 ; 
      RECT 4.72 65.826 4.824 70.2 ; 
      RECT 4.288 65.826 4.392 70.2 ; 
      RECT 3.856 65.826 3.96 70.2 ; 
      RECT 3.424 65.826 3.528 70.2 ; 
      RECT 2.992 65.826 3.096 70.2 ; 
      RECT 2.56 65.826 2.664 70.2 ; 
      RECT 2.128 65.826 2.232 70.2 ; 
      RECT 1.696 65.826 1.8 70.2 ; 
      RECT 1.264 65.826 1.368 70.2 ; 
      RECT 0.832 65.826 0.936 70.2 ; 
      RECT 0.02 65.826 0.36 70.2 ; 
      RECT 34.564 70.146 35.076 74.52 ; 
      RECT 34.508 72.808 35.076 74.098 ; 
      RECT 33.916 71.716 34.164 74.52 ; 
      RECT 33.86 72.954 34.164 73.568 ; 
      RECT 33.916 70.146 34.02 74.52 ; 
      RECT 33.916 70.63 34.076 71.588 ; 
      RECT 33.916 70.146 34.164 70.502 ; 
      RECT 32.728 71.948 33.552 74.52 ; 
      RECT 33.448 70.146 33.552 74.52 ; 
      RECT 32.728 73.056 33.608 74.088 ; 
      RECT 32.728 70.146 33.12 74.52 ; 
      RECT 31.06 70.146 31.392 74.52 ; 
      RECT 31.06 70.5 31.448 74.242 ; 
      RECT 65.776 70.146 66.116 74.52 ; 
      RECT 65.2 70.146 65.304 74.52 ; 
      RECT 64.768 70.146 64.872 74.52 ; 
      RECT 64.336 70.146 64.44 74.52 ; 
      RECT 63.904 70.146 64.008 74.52 ; 
      RECT 63.472 70.146 63.576 74.52 ; 
      RECT 63.04 70.146 63.144 74.52 ; 
      RECT 62.608 70.146 62.712 74.52 ; 
      RECT 62.176 70.146 62.28 74.52 ; 
      RECT 61.744 70.146 61.848 74.52 ; 
      RECT 61.312 70.146 61.416 74.52 ; 
      RECT 60.88 70.146 60.984 74.52 ; 
      RECT 60.448 70.146 60.552 74.52 ; 
      RECT 60.016 70.146 60.12 74.52 ; 
      RECT 59.584 70.146 59.688 74.52 ; 
      RECT 59.152 70.146 59.256 74.52 ; 
      RECT 58.72 70.146 58.824 74.52 ; 
      RECT 58.288 70.146 58.392 74.52 ; 
      RECT 57.856 70.146 57.96 74.52 ; 
      RECT 57.424 70.146 57.528 74.52 ; 
      RECT 56.992 70.146 57.096 74.52 ; 
      RECT 56.56 70.146 56.664 74.52 ; 
      RECT 56.128 70.146 56.232 74.52 ; 
      RECT 55.696 70.146 55.8 74.52 ; 
      RECT 55.264 70.146 55.368 74.52 ; 
      RECT 54.832 70.146 54.936 74.52 ; 
      RECT 54.4 70.146 54.504 74.52 ; 
      RECT 53.968 70.146 54.072 74.52 ; 
      RECT 53.536 70.146 53.64 74.52 ; 
      RECT 53.104 70.146 53.208 74.52 ; 
      RECT 52.672 70.146 52.776 74.52 ; 
      RECT 52.24 70.146 52.344 74.52 ; 
      RECT 51.808 70.146 51.912 74.52 ; 
      RECT 51.376 70.146 51.48 74.52 ; 
      RECT 50.944 70.146 51.048 74.52 ; 
      RECT 50.512 70.146 50.616 74.52 ; 
      RECT 50.08 70.146 50.184 74.52 ; 
      RECT 49.648 70.146 49.752 74.52 ; 
      RECT 49.216 70.146 49.32 74.52 ; 
      RECT 48.784 70.146 48.888 74.52 ; 
      RECT 48.352 70.146 48.456 74.52 ; 
      RECT 47.92 70.146 48.024 74.52 ; 
      RECT 47.488 70.146 47.592 74.52 ; 
      RECT 47.056 70.146 47.16 74.52 ; 
      RECT 46.624 70.146 46.728 74.52 ; 
      RECT 46.192 70.146 46.296 74.52 ; 
      RECT 45.76 70.146 45.864 74.52 ; 
      RECT 45.328 70.146 45.432 74.52 ; 
      RECT 44.896 70.146 45 74.52 ; 
      RECT 44.464 70.146 44.568 74.52 ; 
      RECT 44.032 70.146 44.136 74.52 ; 
      RECT 43.6 70.146 43.704 74.52 ; 
      RECT 43.168 70.146 43.272 74.52 ; 
      RECT 42.736 70.146 42.84 74.52 ; 
      RECT 42.304 70.146 42.408 74.52 ; 
      RECT 41.872 70.146 41.976 74.52 ; 
      RECT 41.44 70.146 41.544 74.52 ; 
      RECT 41.008 70.146 41.112 74.52 ; 
      RECT 40.576 70.146 40.68 74.52 ; 
      RECT 40.144 70.146 40.248 74.52 ; 
      RECT 39.712 70.146 39.816 74.52 ; 
      RECT 39.28 70.146 39.384 74.52 ; 
      RECT 38.848 70.146 38.952 74.52 ; 
      RECT 38.416 70.146 38.52 74.52 ; 
      RECT 37.984 70.146 38.088 74.52 ; 
      RECT 37.552 70.146 37.656 74.52 ; 
      RECT 36.7 70.146 37.008 74.52 ; 
      RECT 29.128 70.146 29.436 74.52 ; 
      RECT 28.48 70.146 28.584 74.52 ; 
      RECT 28.048 70.146 28.152 74.52 ; 
      RECT 27.616 70.146 27.72 74.52 ; 
      RECT 27.184 70.146 27.288 74.52 ; 
      RECT 26.752 70.146 26.856 74.52 ; 
      RECT 26.32 70.146 26.424 74.52 ; 
      RECT 25.888 70.146 25.992 74.52 ; 
      RECT 25.456 70.146 25.56 74.52 ; 
      RECT 25.024 70.146 25.128 74.52 ; 
      RECT 24.592 70.146 24.696 74.52 ; 
      RECT 24.16 70.146 24.264 74.52 ; 
      RECT 23.728 70.146 23.832 74.52 ; 
      RECT 23.296 70.146 23.4 74.52 ; 
      RECT 22.864 70.146 22.968 74.52 ; 
      RECT 22.432 70.146 22.536 74.52 ; 
      RECT 22 70.146 22.104 74.52 ; 
      RECT 21.568 70.146 21.672 74.52 ; 
      RECT 21.136 70.146 21.24 74.52 ; 
      RECT 20.704 70.146 20.808 74.52 ; 
      RECT 20.272 70.146 20.376 74.52 ; 
      RECT 19.84 70.146 19.944 74.52 ; 
      RECT 19.408 70.146 19.512 74.52 ; 
      RECT 18.976 70.146 19.08 74.52 ; 
      RECT 18.544 70.146 18.648 74.52 ; 
      RECT 18.112 70.146 18.216 74.52 ; 
      RECT 17.68 70.146 17.784 74.52 ; 
      RECT 17.248 70.146 17.352 74.52 ; 
      RECT 16.816 70.146 16.92 74.52 ; 
      RECT 16.384 70.146 16.488 74.52 ; 
      RECT 15.952 70.146 16.056 74.52 ; 
      RECT 15.52 70.146 15.624 74.52 ; 
      RECT 15.088 70.146 15.192 74.52 ; 
      RECT 14.656 70.146 14.76 74.52 ; 
      RECT 14.224 70.146 14.328 74.52 ; 
      RECT 13.792 70.146 13.896 74.52 ; 
      RECT 13.36 70.146 13.464 74.52 ; 
      RECT 12.928 70.146 13.032 74.52 ; 
      RECT 12.496 70.146 12.6 74.52 ; 
      RECT 12.064 70.146 12.168 74.52 ; 
      RECT 11.632 70.146 11.736 74.52 ; 
      RECT 11.2 70.146 11.304 74.52 ; 
      RECT 10.768 70.146 10.872 74.52 ; 
      RECT 10.336 70.146 10.44 74.52 ; 
      RECT 9.904 70.146 10.008 74.52 ; 
      RECT 9.472 70.146 9.576 74.52 ; 
      RECT 9.04 70.146 9.144 74.52 ; 
      RECT 8.608 70.146 8.712 74.52 ; 
      RECT 8.176 70.146 8.28 74.52 ; 
      RECT 7.744 70.146 7.848 74.52 ; 
      RECT 7.312 70.146 7.416 74.52 ; 
      RECT 6.88 70.146 6.984 74.52 ; 
      RECT 6.448 70.146 6.552 74.52 ; 
      RECT 6.016 70.146 6.12 74.52 ; 
      RECT 5.584 70.146 5.688 74.52 ; 
      RECT 5.152 70.146 5.256 74.52 ; 
      RECT 4.72 70.146 4.824 74.52 ; 
      RECT 4.288 70.146 4.392 74.52 ; 
      RECT 3.856 70.146 3.96 74.52 ; 
      RECT 3.424 70.146 3.528 74.52 ; 
      RECT 2.992 70.146 3.096 74.52 ; 
      RECT 2.56 70.146 2.664 74.52 ; 
      RECT 2.128 70.146 2.232 74.52 ; 
      RECT 1.696 70.146 1.8 74.52 ; 
      RECT 1.264 70.146 1.368 74.52 ; 
      RECT 0.832 70.146 0.936 74.52 ; 
      RECT 0.02 70.146 0.36 74.52 ; 
      RECT 0 107.238 66.096 109.002 ; 
      RECT 65.756 74.388 66.096 109.002 ; 
      RECT 37.532 80.404 65.284 109.002 ; 
      RECT 43.364 74.388 65.284 109.002 ; 
      RECT 28.892 107.208 37.204 109.002 ; 
      RECT 31.988 107.082 37.204 109.002 ; 
      RECT 0.812 79.624 28.564 109.002 ; 
      RECT 27.38 74.388 28.564 109.002 ; 
      RECT 0 74.388 0.34 109.002 ; 
      RECT 28.892 80.836 31.372 109.002 ; 
      RECT 31.988 107.064 37.06 109.002 ; 
      RECT 34.58 80.008 37.06 109.002 ; 
      RECT 34.544 106.036 37.06 109.002 ; 
      RECT 33.896 106.036 34.144 109.002 ; 
      RECT 31.988 106.036 33.532 109.002 ; 
      RECT 37.532 89.56 65.34 106.976 ; 
      RECT 0.756 89.56 28.564 106.976 ; 
      RECT 37.476 89.56 65.34 106.958 ; 
      RECT 0.756 89.56 28.62 106.958 ; 
      RECT 28.836 89.56 31.372 106.954 ; 
      RECT 32.708 77.128 33.388 109.002 ; 
      RECT 33.14 74.388 33.388 109.002 ; 
      RECT 29.972 76.072 31.516 105.448 ; 
      RECT 28.836 105.268 31.572 105.416 ; 
      RECT 34.524 100.972 37.06 105.404 ; 
      RECT 32.652 104.212 33.388 105.116 ; 
      RECT 32.708 101.908 33.444 102.956 ; 
      RECT 28.836 101.116 31.572 102.956 ; 
      RECT 32.652 98.956 33.388 100.796 ; 
      RECT 34.524 90.82 37.06 100.148 ; 
      RECT 28.836 93.412 31.572 97.988 ; 
      RECT 32.708 92.332 33.444 97.556 ; 
      RECT 32.652 94.636 33.444 96.476 ; 
      RECT 32.652 81.676 33.388 94.316 ; 
      RECT 32.652 81.676 33.444 92.156 ; 
      RECT 28.836 91.252 31.572 92.156 ; 
      RECT 34.58 80.008 37.204 89.432 ; 
      RECT 34.524 79.516 36.988 86.66 ; 
      RECT 28.892 83.404 31.572 84.884 ; 
      RECT 32.708 80.596 33.444 81.356 ; 
      RECT 29.108 80.452 31.572 81.212 ; 
      RECT 32.652 80.02 33.388 80.564 ; 
      RECT 29.108 77.452 31.516 105.448 ; 
      RECT 32.708 79.516 33.444 80.42 ; 
      RECT 38.18 79.636 65.284 109.002 ; 
      RECT 42.5 79.624 65.284 109.002 ; 
      RECT 37.532 74.388 37.852 109.002 ; 
      RECT 28.892 77.128 29.644 80.384 ; 
      RECT 37.532 74.388 38.716 80 ; 
      RECT 37.532 78.856 42.172 80 ; 
      RECT 42.5 74.388 43.036 109.002 ; 
      RECT 23.924 78.1 27.052 109.002 ; 
      RECT 0.812 74.388 23.596 109.002 ; 
      RECT 34.58 77.452 36.988 109.002 ; 
      RECT 34.724 75.094 37.204 79.388 ; 
      RECT 37.532 78.856 43.036 79.232 ; 
      RECT 41.636 74.388 65.284 79.22 ; 
      RECT 26.516 74.388 28.564 79.22 ; 
      RECT 32.652 78.94 33.444 79.196 ; 
      RECT 32.652 78.436 33.388 79.196 ; 
      RECT 40.772 77.32 65.284 79.22 ; 
      RECT 37.532 77.452 40.444 80 ; 
      RECT 32.708 77.356 33.444 78.404 ; 
      RECT 0.812 77.32 26.188 79.22 ; 
      RECT 25.652 74.388 26.188 109.002 ; 
      RECT 39.908 74.388 41.308 77.876 ; 
      RECT 37.532 77.128 39.58 80 ; 
      RECT 39.044 74.388 39.58 109.002 ; 
      RECT 24.788 77.128 26.188 109.002 ; 
      RECT 0.812 74.388 24.46 79.22 ; 
      RECT 32.708 74.388 32.812 109.002 ; 
      RECT 29.252 74.388 29.644 109.002 ; 
      RECT 24.788 74.388 25.324 109.002 ; 
      RECT 39.044 74.388 41.308 76.928 ; 
      RECT 34.58 74.388 36.988 76.928 ; 
      RECT 29.252 74.388 31.372 76.928 ; 
      RECT 25.652 74.388 28.564 76.928 ; 
      RECT 39.044 74.388 65.284 76.916 ; 
      RECT 0.812 74.388 25.324 76.916 ; 
      RECT 34.524 76.276 37.204 76.892 ; 
      RECT 37.532 74.388 65.284 75.86 ; 
      RECT 32.708 74.388 33.388 75.86 ; 
      RECT 28.892 74.388 31.372 75.86 ; 
      RECT 0.812 74.388 28.564 75.86 ; 
      RECT 31.988 74.388 33.388 75.448 ; 
      RECT 34.544 74.388 36.988 75.048 ; 
      RECT 31.988 74.388 33.532 75.048 ; 
      RECT 39.06 74.282 39.132 109.002 ; 
      RECT 38.628 74.282 38.7 109.002 ; 
      RECT 27.396 74.332 27.468 109.002 ; 
      RECT 26.964 74.332 27.036 109.002 ; 
      RECT 26.532 74.332 26.604 109.002 ; 
      RECT 26.1 74.332 26.172 109.002 ; 
      RECT 25.668 74.282 25.74 109.002 ; 
      RECT 25.236 74.282 25.308 109.002 ; 
      RECT 24.804 74.332 24.876 109.002 ; 
      RECT 24.372 74.332 24.444 109.002 ; 
      RECT 23.94 74.332 24.012 109.002 ; 
      RECT 23.508 74.332 23.58 109.002 ; 
      RECT 33.896 74.388 34.144 75.048 ; 
        RECT 34.564 106.974 35.076 111.348 ; 
        RECT 34.508 109.636 35.076 110.926 ; 
        RECT 33.916 108.544 34.164 111.348 ; 
        RECT 33.86 109.782 34.164 110.396 ; 
        RECT 33.916 106.974 34.02 111.348 ; 
        RECT 33.916 107.458 34.076 108.416 ; 
        RECT 33.916 106.974 34.164 107.33 ; 
        RECT 32.728 108.776 33.552 111.348 ; 
        RECT 33.448 106.974 33.552 111.348 ; 
        RECT 32.728 109.884 33.608 110.916 ; 
        RECT 32.728 106.974 33.12 111.348 ; 
        RECT 31.06 106.974 31.392 111.348 ; 
        RECT 31.06 107.328 31.448 111.07 ; 
        RECT 65.776 106.974 66.116 111.348 ; 
        RECT 65.2 106.974 65.304 111.348 ; 
        RECT 64.768 106.974 64.872 111.348 ; 
        RECT 64.336 106.974 64.44 111.348 ; 
        RECT 63.904 106.974 64.008 111.348 ; 
        RECT 63.472 106.974 63.576 111.348 ; 
        RECT 63.04 106.974 63.144 111.348 ; 
        RECT 62.608 106.974 62.712 111.348 ; 
        RECT 62.176 106.974 62.28 111.348 ; 
        RECT 61.744 106.974 61.848 111.348 ; 
        RECT 61.312 106.974 61.416 111.348 ; 
        RECT 60.88 106.974 60.984 111.348 ; 
        RECT 60.448 106.974 60.552 111.348 ; 
        RECT 60.016 106.974 60.12 111.348 ; 
        RECT 59.584 106.974 59.688 111.348 ; 
        RECT 59.152 106.974 59.256 111.348 ; 
        RECT 58.72 106.974 58.824 111.348 ; 
        RECT 58.288 106.974 58.392 111.348 ; 
        RECT 57.856 106.974 57.96 111.348 ; 
        RECT 57.424 106.974 57.528 111.348 ; 
        RECT 56.992 106.974 57.096 111.348 ; 
        RECT 56.56 106.974 56.664 111.348 ; 
        RECT 56.128 106.974 56.232 111.348 ; 
        RECT 55.696 106.974 55.8 111.348 ; 
        RECT 55.264 106.974 55.368 111.348 ; 
        RECT 54.832 106.974 54.936 111.348 ; 
        RECT 54.4 106.974 54.504 111.348 ; 
        RECT 53.968 106.974 54.072 111.348 ; 
        RECT 53.536 106.974 53.64 111.348 ; 
        RECT 53.104 106.974 53.208 111.348 ; 
        RECT 52.672 106.974 52.776 111.348 ; 
        RECT 52.24 106.974 52.344 111.348 ; 
        RECT 51.808 106.974 51.912 111.348 ; 
        RECT 51.376 106.974 51.48 111.348 ; 
        RECT 50.944 106.974 51.048 111.348 ; 
        RECT 50.512 106.974 50.616 111.348 ; 
        RECT 50.08 106.974 50.184 111.348 ; 
        RECT 49.648 106.974 49.752 111.348 ; 
        RECT 49.216 106.974 49.32 111.348 ; 
        RECT 48.784 106.974 48.888 111.348 ; 
        RECT 48.352 106.974 48.456 111.348 ; 
        RECT 47.92 106.974 48.024 111.348 ; 
        RECT 47.488 106.974 47.592 111.348 ; 
        RECT 47.056 106.974 47.16 111.348 ; 
        RECT 46.624 106.974 46.728 111.348 ; 
        RECT 46.192 106.974 46.296 111.348 ; 
        RECT 45.76 106.974 45.864 111.348 ; 
        RECT 45.328 106.974 45.432 111.348 ; 
        RECT 44.896 106.974 45 111.348 ; 
        RECT 44.464 106.974 44.568 111.348 ; 
        RECT 44.032 106.974 44.136 111.348 ; 
        RECT 43.6 106.974 43.704 111.348 ; 
        RECT 43.168 106.974 43.272 111.348 ; 
        RECT 42.736 106.974 42.84 111.348 ; 
        RECT 42.304 106.974 42.408 111.348 ; 
        RECT 41.872 106.974 41.976 111.348 ; 
        RECT 41.44 106.974 41.544 111.348 ; 
        RECT 41.008 106.974 41.112 111.348 ; 
        RECT 40.576 106.974 40.68 111.348 ; 
        RECT 40.144 106.974 40.248 111.348 ; 
        RECT 39.712 106.974 39.816 111.348 ; 
        RECT 39.28 106.974 39.384 111.348 ; 
        RECT 38.848 106.974 38.952 111.348 ; 
        RECT 38.416 106.974 38.52 111.348 ; 
        RECT 37.984 106.974 38.088 111.348 ; 
        RECT 37.552 106.974 37.656 111.348 ; 
        RECT 36.7 106.974 37.008 111.348 ; 
        RECT 29.128 106.974 29.436 111.348 ; 
        RECT 28.48 106.974 28.584 111.348 ; 
        RECT 28.048 106.974 28.152 111.348 ; 
        RECT 27.616 106.974 27.72 111.348 ; 
        RECT 27.184 106.974 27.288 111.348 ; 
        RECT 26.752 106.974 26.856 111.348 ; 
        RECT 26.32 106.974 26.424 111.348 ; 
        RECT 25.888 106.974 25.992 111.348 ; 
        RECT 25.456 106.974 25.56 111.348 ; 
        RECT 25.024 106.974 25.128 111.348 ; 
        RECT 24.592 106.974 24.696 111.348 ; 
        RECT 24.16 106.974 24.264 111.348 ; 
        RECT 23.728 106.974 23.832 111.348 ; 
        RECT 23.296 106.974 23.4 111.348 ; 
        RECT 22.864 106.974 22.968 111.348 ; 
        RECT 22.432 106.974 22.536 111.348 ; 
        RECT 22 106.974 22.104 111.348 ; 
        RECT 21.568 106.974 21.672 111.348 ; 
        RECT 21.136 106.974 21.24 111.348 ; 
        RECT 20.704 106.974 20.808 111.348 ; 
        RECT 20.272 106.974 20.376 111.348 ; 
        RECT 19.84 106.974 19.944 111.348 ; 
        RECT 19.408 106.974 19.512 111.348 ; 
        RECT 18.976 106.974 19.08 111.348 ; 
        RECT 18.544 106.974 18.648 111.348 ; 
        RECT 18.112 106.974 18.216 111.348 ; 
        RECT 17.68 106.974 17.784 111.348 ; 
        RECT 17.248 106.974 17.352 111.348 ; 
        RECT 16.816 106.974 16.92 111.348 ; 
        RECT 16.384 106.974 16.488 111.348 ; 
        RECT 15.952 106.974 16.056 111.348 ; 
        RECT 15.52 106.974 15.624 111.348 ; 
        RECT 15.088 106.974 15.192 111.348 ; 
        RECT 14.656 106.974 14.76 111.348 ; 
        RECT 14.224 106.974 14.328 111.348 ; 
        RECT 13.792 106.974 13.896 111.348 ; 
        RECT 13.36 106.974 13.464 111.348 ; 
        RECT 12.928 106.974 13.032 111.348 ; 
        RECT 12.496 106.974 12.6 111.348 ; 
        RECT 12.064 106.974 12.168 111.348 ; 
        RECT 11.632 106.974 11.736 111.348 ; 
        RECT 11.2 106.974 11.304 111.348 ; 
        RECT 10.768 106.974 10.872 111.348 ; 
        RECT 10.336 106.974 10.44 111.348 ; 
        RECT 9.904 106.974 10.008 111.348 ; 
        RECT 9.472 106.974 9.576 111.348 ; 
        RECT 9.04 106.974 9.144 111.348 ; 
        RECT 8.608 106.974 8.712 111.348 ; 
        RECT 8.176 106.974 8.28 111.348 ; 
        RECT 7.744 106.974 7.848 111.348 ; 
        RECT 7.312 106.974 7.416 111.348 ; 
        RECT 6.88 106.974 6.984 111.348 ; 
        RECT 6.448 106.974 6.552 111.348 ; 
        RECT 6.016 106.974 6.12 111.348 ; 
        RECT 5.584 106.974 5.688 111.348 ; 
        RECT 5.152 106.974 5.256 111.348 ; 
        RECT 4.72 106.974 4.824 111.348 ; 
        RECT 4.288 106.974 4.392 111.348 ; 
        RECT 3.856 106.974 3.96 111.348 ; 
        RECT 3.424 106.974 3.528 111.348 ; 
        RECT 2.992 106.974 3.096 111.348 ; 
        RECT 2.56 106.974 2.664 111.348 ; 
        RECT 2.128 106.974 2.232 111.348 ; 
        RECT 1.696 106.974 1.8 111.348 ; 
        RECT 1.264 106.974 1.368 111.348 ; 
        RECT 0.832 106.974 0.936 111.348 ; 
        RECT 0.02 106.974 0.36 111.348 ; 
        RECT 34.564 111.294 35.076 115.668 ; 
        RECT 34.508 113.956 35.076 115.246 ; 
        RECT 33.916 112.864 34.164 115.668 ; 
        RECT 33.86 114.102 34.164 114.716 ; 
        RECT 33.916 111.294 34.02 115.668 ; 
        RECT 33.916 111.778 34.076 112.736 ; 
        RECT 33.916 111.294 34.164 111.65 ; 
        RECT 32.728 113.096 33.552 115.668 ; 
        RECT 33.448 111.294 33.552 115.668 ; 
        RECT 32.728 114.204 33.608 115.236 ; 
        RECT 32.728 111.294 33.12 115.668 ; 
        RECT 31.06 111.294 31.392 115.668 ; 
        RECT 31.06 111.648 31.448 115.39 ; 
        RECT 65.776 111.294 66.116 115.668 ; 
        RECT 65.2 111.294 65.304 115.668 ; 
        RECT 64.768 111.294 64.872 115.668 ; 
        RECT 64.336 111.294 64.44 115.668 ; 
        RECT 63.904 111.294 64.008 115.668 ; 
        RECT 63.472 111.294 63.576 115.668 ; 
        RECT 63.04 111.294 63.144 115.668 ; 
        RECT 62.608 111.294 62.712 115.668 ; 
        RECT 62.176 111.294 62.28 115.668 ; 
        RECT 61.744 111.294 61.848 115.668 ; 
        RECT 61.312 111.294 61.416 115.668 ; 
        RECT 60.88 111.294 60.984 115.668 ; 
        RECT 60.448 111.294 60.552 115.668 ; 
        RECT 60.016 111.294 60.12 115.668 ; 
        RECT 59.584 111.294 59.688 115.668 ; 
        RECT 59.152 111.294 59.256 115.668 ; 
        RECT 58.72 111.294 58.824 115.668 ; 
        RECT 58.288 111.294 58.392 115.668 ; 
        RECT 57.856 111.294 57.96 115.668 ; 
        RECT 57.424 111.294 57.528 115.668 ; 
        RECT 56.992 111.294 57.096 115.668 ; 
        RECT 56.56 111.294 56.664 115.668 ; 
        RECT 56.128 111.294 56.232 115.668 ; 
        RECT 55.696 111.294 55.8 115.668 ; 
        RECT 55.264 111.294 55.368 115.668 ; 
        RECT 54.832 111.294 54.936 115.668 ; 
        RECT 54.4 111.294 54.504 115.668 ; 
        RECT 53.968 111.294 54.072 115.668 ; 
        RECT 53.536 111.294 53.64 115.668 ; 
        RECT 53.104 111.294 53.208 115.668 ; 
        RECT 52.672 111.294 52.776 115.668 ; 
        RECT 52.24 111.294 52.344 115.668 ; 
        RECT 51.808 111.294 51.912 115.668 ; 
        RECT 51.376 111.294 51.48 115.668 ; 
        RECT 50.944 111.294 51.048 115.668 ; 
        RECT 50.512 111.294 50.616 115.668 ; 
        RECT 50.08 111.294 50.184 115.668 ; 
        RECT 49.648 111.294 49.752 115.668 ; 
        RECT 49.216 111.294 49.32 115.668 ; 
        RECT 48.784 111.294 48.888 115.668 ; 
        RECT 48.352 111.294 48.456 115.668 ; 
        RECT 47.92 111.294 48.024 115.668 ; 
        RECT 47.488 111.294 47.592 115.668 ; 
        RECT 47.056 111.294 47.16 115.668 ; 
        RECT 46.624 111.294 46.728 115.668 ; 
        RECT 46.192 111.294 46.296 115.668 ; 
        RECT 45.76 111.294 45.864 115.668 ; 
        RECT 45.328 111.294 45.432 115.668 ; 
        RECT 44.896 111.294 45 115.668 ; 
        RECT 44.464 111.294 44.568 115.668 ; 
        RECT 44.032 111.294 44.136 115.668 ; 
        RECT 43.6 111.294 43.704 115.668 ; 
        RECT 43.168 111.294 43.272 115.668 ; 
        RECT 42.736 111.294 42.84 115.668 ; 
        RECT 42.304 111.294 42.408 115.668 ; 
        RECT 41.872 111.294 41.976 115.668 ; 
        RECT 41.44 111.294 41.544 115.668 ; 
        RECT 41.008 111.294 41.112 115.668 ; 
        RECT 40.576 111.294 40.68 115.668 ; 
        RECT 40.144 111.294 40.248 115.668 ; 
        RECT 39.712 111.294 39.816 115.668 ; 
        RECT 39.28 111.294 39.384 115.668 ; 
        RECT 38.848 111.294 38.952 115.668 ; 
        RECT 38.416 111.294 38.52 115.668 ; 
        RECT 37.984 111.294 38.088 115.668 ; 
        RECT 37.552 111.294 37.656 115.668 ; 
        RECT 36.7 111.294 37.008 115.668 ; 
        RECT 29.128 111.294 29.436 115.668 ; 
        RECT 28.48 111.294 28.584 115.668 ; 
        RECT 28.048 111.294 28.152 115.668 ; 
        RECT 27.616 111.294 27.72 115.668 ; 
        RECT 27.184 111.294 27.288 115.668 ; 
        RECT 26.752 111.294 26.856 115.668 ; 
        RECT 26.32 111.294 26.424 115.668 ; 
        RECT 25.888 111.294 25.992 115.668 ; 
        RECT 25.456 111.294 25.56 115.668 ; 
        RECT 25.024 111.294 25.128 115.668 ; 
        RECT 24.592 111.294 24.696 115.668 ; 
        RECT 24.16 111.294 24.264 115.668 ; 
        RECT 23.728 111.294 23.832 115.668 ; 
        RECT 23.296 111.294 23.4 115.668 ; 
        RECT 22.864 111.294 22.968 115.668 ; 
        RECT 22.432 111.294 22.536 115.668 ; 
        RECT 22 111.294 22.104 115.668 ; 
        RECT 21.568 111.294 21.672 115.668 ; 
        RECT 21.136 111.294 21.24 115.668 ; 
        RECT 20.704 111.294 20.808 115.668 ; 
        RECT 20.272 111.294 20.376 115.668 ; 
        RECT 19.84 111.294 19.944 115.668 ; 
        RECT 19.408 111.294 19.512 115.668 ; 
        RECT 18.976 111.294 19.08 115.668 ; 
        RECT 18.544 111.294 18.648 115.668 ; 
        RECT 18.112 111.294 18.216 115.668 ; 
        RECT 17.68 111.294 17.784 115.668 ; 
        RECT 17.248 111.294 17.352 115.668 ; 
        RECT 16.816 111.294 16.92 115.668 ; 
        RECT 16.384 111.294 16.488 115.668 ; 
        RECT 15.952 111.294 16.056 115.668 ; 
        RECT 15.52 111.294 15.624 115.668 ; 
        RECT 15.088 111.294 15.192 115.668 ; 
        RECT 14.656 111.294 14.76 115.668 ; 
        RECT 14.224 111.294 14.328 115.668 ; 
        RECT 13.792 111.294 13.896 115.668 ; 
        RECT 13.36 111.294 13.464 115.668 ; 
        RECT 12.928 111.294 13.032 115.668 ; 
        RECT 12.496 111.294 12.6 115.668 ; 
        RECT 12.064 111.294 12.168 115.668 ; 
        RECT 11.632 111.294 11.736 115.668 ; 
        RECT 11.2 111.294 11.304 115.668 ; 
        RECT 10.768 111.294 10.872 115.668 ; 
        RECT 10.336 111.294 10.44 115.668 ; 
        RECT 9.904 111.294 10.008 115.668 ; 
        RECT 9.472 111.294 9.576 115.668 ; 
        RECT 9.04 111.294 9.144 115.668 ; 
        RECT 8.608 111.294 8.712 115.668 ; 
        RECT 8.176 111.294 8.28 115.668 ; 
        RECT 7.744 111.294 7.848 115.668 ; 
        RECT 7.312 111.294 7.416 115.668 ; 
        RECT 6.88 111.294 6.984 115.668 ; 
        RECT 6.448 111.294 6.552 115.668 ; 
        RECT 6.016 111.294 6.12 115.668 ; 
        RECT 5.584 111.294 5.688 115.668 ; 
        RECT 5.152 111.294 5.256 115.668 ; 
        RECT 4.72 111.294 4.824 115.668 ; 
        RECT 4.288 111.294 4.392 115.668 ; 
        RECT 3.856 111.294 3.96 115.668 ; 
        RECT 3.424 111.294 3.528 115.668 ; 
        RECT 2.992 111.294 3.096 115.668 ; 
        RECT 2.56 111.294 2.664 115.668 ; 
        RECT 2.128 111.294 2.232 115.668 ; 
        RECT 1.696 111.294 1.8 115.668 ; 
        RECT 1.264 111.294 1.368 115.668 ; 
        RECT 0.832 111.294 0.936 115.668 ; 
        RECT 0.02 111.294 0.36 115.668 ; 
        RECT 34.564 115.614 35.076 119.988 ; 
        RECT 34.508 118.276 35.076 119.566 ; 
        RECT 33.916 117.184 34.164 119.988 ; 
        RECT 33.86 118.422 34.164 119.036 ; 
        RECT 33.916 115.614 34.02 119.988 ; 
        RECT 33.916 116.098 34.076 117.056 ; 
        RECT 33.916 115.614 34.164 115.97 ; 
        RECT 32.728 117.416 33.552 119.988 ; 
        RECT 33.448 115.614 33.552 119.988 ; 
        RECT 32.728 118.524 33.608 119.556 ; 
        RECT 32.728 115.614 33.12 119.988 ; 
        RECT 31.06 115.614 31.392 119.988 ; 
        RECT 31.06 115.968 31.448 119.71 ; 
        RECT 65.776 115.614 66.116 119.988 ; 
        RECT 65.2 115.614 65.304 119.988 ; 
        RECT 64.768 115.614 64.872 119.988 ; 
        RECT 64.336 115.614 64.44 119.988 ; 
        RECT 63.904 115.614 64.008 119.988 ; 
        RECT 63.472 115.614 63.576 119.988 ; 
        RECT 63.04 115.614 63.144 119.988 ; 
        RECT 62.608 115.614 62.712 119.988 ; 
        RECT 62.176 115.614 62.28 119.988 ; 
        RECT 61.744 115.614 61.848 119.988 ; 
        RECT 61.312 115.614 61.416 119.988 ; 
        RECT 60.88 115.614 60.984 119.988 ; 
        RECT 60.448 115.614 60.552 119.988 ; 
        RECT 60.016 115.614 60.12 119.988 ; 
        RECT 59.584 115.614 59.688 119.988 ; 
        RECT 59.152 115.614 59.256 119.988 ; 
        RECT 58.72 115.614 58.824 119.988 ; 
        RECT 58.288 115.614 58.392 119.988 ; 
        RECT 57.856 115.614 57.96 119.988 ; 
        RECT 57.424 115.614 57.528 119.988 ; 
        RECT 56.992 115.614 57.096 119.988 ; 
        RECT 56.56 115.614 56.664 119.988 ; 
        RECT 56.128 115.614 56.232 119.988 ; 
        RECT 55.696 115.614 55.8 119.988 ; 
        RECT 55.264 115.614 55.368 119.988 ; 
        RECT 54.832 115.614 54.936 119.988 ; 
        RECT 54.4 115.614 54.504 119.988 ; 
        RECT 53.968 115.614 54.072 119.988 ; 
        RECT 53.536 115.614 53.64 119.988 ; 
        RECT 53.104 115.614 53.208 119.988 ; 
        RECT 52.672 115.614 52.776 119.988 ; 
        RECT 52.24 115.614 52.344 119.988 ; 
        RECT 51.808 115.614 51.912 119.988 ; 
        RECT 51.376 115.614 51.48 119.988 ; 
        RECT 50.944 115.614 51.048 119.988 ; 
        RECT 50.512 115.614 50.616 119.988 ; 
        RECT 50.08 115.614 50.184 119.988 ; 
        RECT 49.648 115.614 49.752 119.988 ; 
        RECT 49.216 115.614 49.32 119.988 ; 
        RECT 48.784 115.614 48.888 119.988 ; 
        RECT 48.352 115.614 48.456 119.988 ; 
        RECT 47.92 115.614 48.024 119.988 ; 
        RECT 47.488 115.614 47.592 119.988 ; 
        RECT 47.056 115.614 47.16 119.988 ; 
        RECT 46.624 115.614 46.728 119.988 ; 
        RECT 46.192 115.614 46.296 119.988 ; 
        RECT 45.76 115.614 45.864 119.988 ; 
        RECT 45.328 115.614 45.432 119.988 ; 
        RECT 44.896 115.614 45 119.988 ; 
        RECT 44.464 115.614 44.568 119.988 ; 
        RECT 44.032 115.614 44.136 119.988 ; 
        RECT 43.6 115.614 43.704 119.988 ; 
        RECT 43.168 115.614 43.272 119.988 ; 
        RECT 42.736 115.614 42.84 119.988 ; 
        RECT 42.304 115.614 42.408 119.988 ; 
        RECT 41.872 115.614 41.976 119.988 ; 
        RECT 41.44 115.614 41.544 119.988 ; 
        RECT 41.008 115.614 41.112 119.988 ; 
        RECT 40.576 115.614 40.68 119.988 ; 
        RECT 40.144 115.614 40.248 119.988 ; 
        RECT 39.712 115.614 39.816 119.988 ; 
        RECT 39.28 115.614 39.384 119.988 ; 
        RECT 38.848 115.614 38.952 119.988 ; 
        RECT 38.416 115.614 38.52 119.988 ; 
        RECT 37.984 115.614 38.088 119.988 ; 
        RECT 37.552 115.614 37.656 119.988 ; 
        RECT 36.7 115.614 37.008 119.988 ; 
        RECT 29.128 115.614 29.436 119.988 ; 
        RECT 28.48 115.614 28.584 119.988 ; 
        RECT 28.048 115.614 28.152 119.988 ; 
        RECT 27.616 115.614 27.72 119.988 ; 
        RECT 27.184 115.614 27.288 119.988 ; 
        RECT 26.752 115.614 26.856 119.988 ; 
        RECT 26.32 115.614 26.424 119.988 ; 
        RECT 25.888 115.614 25.992 119.988 ; 
        RECT 25.456 115.614 25.56 119.988 ; 
        RECT 25.024 115.614 25.128 119.988 ; 
        RECT 24.592 115.614 24.696 119.988 ; 
        RECT 24.16 115.614 24.264 119.988 ; 
        RECT 23.728 115.614 23.832 119.988 ; 
        RECT 23.296 115.614 23.4 119.988 ; 
        RECT 22.864 115.614 22.968 119.988 ; 
        RECT 22.432 115.614 22.536 119.988 ; 
        RECT 22 115.614 22.104 119.988 ; 
        RECT 21.568 115.614 21.672 119.988 ; 
        RECT 21.136 115.614 21.24 119.988 ; 
        RECT 20.704 115.614 20.808 119.988 ; 
        RECT 20.272 115.614 20.376 119.988 ; 
        RECT 19.84 115.614 19.944 119.988 ; 
        RECT 19.408 115.614 19.512 119.988 ; 
        RECT 18.976 115.614 19.08 119.988 ; 
        RECT 18.544 115.614 18.648 119.988 ; 
        RECT 18.112 115.614 18.216 119.988 ; 
        RECT 17.68 115.614 17.784 119.988 ; 
        RECT 17.248 115.614 17.352 119.988 ; 
        RECT 16.816 115.614 16.92 119.988 ; 
        RECT 16.384 115.614 16.488 119.988 ; 
        RECT 15.952 115.614 16.056 119.988 ; 
        RECT 15.52 115.614 15.624 119.988 ; 
        RECT 15.088 115.614 15.192 119.988 ; 
        RECT 14.656 115.614 14.76 119.988 ; 
        RECT 14.224 115.614 14.328 119.988 ; 
        RECT 13.792 115.614 13.896 119.988 ; 
        RECT 13.36 115.614 13.464 119.988 ; 
        RECT 12.928 115.614 13.032 119.988 ; 
        RECT 12.496 115.614 12.6 119.988 ; 
        RECT 12.064 115.614 12.168 119.988 ; 
        RECT 11.632 115.614 11.736 119.988 ; 
        RECT 11.2 115.614 11.304 119.988 ; 
        RECT 10.768 115.614 10.872 119.988 ; 
        RECT 10.336 115.614 10.44 119.988 ; 
        RECT 9.904 115.614 10.008 119.988 ; 
        RECT 9.472 115.614 9.576 119.988 ; 
        RECT 9.04 115.614 9.144 119.988 ; 
        RECT 8.608 115.614 8.712 119.988 ; 
        RECT 8.176 115.614 8.28 119.988 ; 
        RECT 7.744 115.614 7.848 119.988 ; 
        RECT 7.312 115.614 7.416 119.988 ; 
        RECT 6.88 115.614 6.984 119.988 ; 
        RECT 6.448 115.614 6.552 119.988 ; 
        RECT 6.016 115.614 6.12 119.988 ; 
        RECT 5.584 115.614 5.688 119.988 ; 
        RECT 5.152 115.614 5.256 119.988 ; 
        RECT 4.72 115.614 4.824 119.988 ; 
        RECT 4.288 115.614 4.392 119.988 ; 
        RECT 3.856 115.614 3.96 119.988 ; 
        RECT 3.424 115.614 3.528 119.988 ; 
        RECT 2.992 115.614 3.096 119.988 ; 
        RECT 2.56 115.614 2.664 119.988 ; 
        RECT 2.128 115.614 2.232 119.988 ; 
        RECT 1.696 115.614 1.8 119.988 ; 
        RECT 1.264 115.614 1.368 119.988 ; 
        RECT 0.832 115.614 0.936 119.988 ; 
        RECT 0.02 115.614 0.36 119.988 ; 
        RECT 34.564 119.934 35.076 124.308 ; 
        RECT 34.508 122.596 35.076 123.886 ; 
        RECT 33.916 121.504 34.164 124.308 ; 
        RECT 33.86 122.742 34.164 123.356 ; 
        RECT 33.916 119.934 34.02 124.308 ; 
        RECT 33.916 120.418 34.076 121.376 ; 
        RECT 33.916 119.934 34.164 120.29 ; 
        RECT 32.728 121.736 33.552 124.308 ; 
        RECT 33.448 119.934 33.552 124.308 ; 
        RECT 32.728 122.844 33.608 123.876 ; 
        RECT 32.728 119.934 33.12 124.308 ; 
        RECT 31.06 119.934 31.392 124.308 ; 
        RECT 31.06 120.288 31.448 124.03 ; 
        RECT 65.776 119.934 66.116 124.308 ; 
        RECT 65.2 119.934 65.304 124.308 ; 
        RECT 64.768 119.934 64.872 124.308 ; 
        RECT 64.336 119.934 64.44 124.308 ; 
        RECT 63.904 119.934 64.008 124.308 ; 
        RECT 63.472 119.934 63.576 124.308 ; 
        RECT 63.04 119.934 63.144 124.308 ; 
        RECT 62.608 119.934 62.712 124.308 ; 
        RECT 62.176 119.934 62.28 124.308 ; 
        RECT 61.744 119.934 61.848 124.308 ; 
        RECT 61.312 119.934 61.416 124.308 ; 
        RECT 60.88 119.934 60.984 124.308 ; 
        RECT 60.448 119.934 60.552 124.308 ; 
        RECT 60.016 119.934 60.12 124.308 ; 
        RECT 59.584 119.934 59.688 124.308 ; 
        RECT 59.152 119.934 59.256 124.308 ; 
        RECT 58.72 119.934 58.824 124.308 ; 
        RECT 58.288 119.934 58.392 124.308 ; 
        RECT 57.856 119.934 57.96 124.308 ; 
        RECT 57.424 119.934 57.528 124.308 ; 
        RECT 56.992 119.934 57.096 124.308 ; 
        RECT 56.56 119.934 56.664 124.308 ; 
        RECT 56.128 119.934 56.232 124.308 ; 
        RECT 55.696 119.934 55.8 124.308 ; 
        RECT 55.264 119.934 55.368 124.308 ; 
        RECT 54.832 119.934 54.936 124.308 ; 
        RECT 54.4 119.934 54.504 124.308 ; 
        RECT 53.968 119.934 54.072 124.308 ; 
        RECT 53.536 119.934 53.64 124.308 ; 
        RECT 53.104 119.934 53.208 124.308 ; 
        RECT 52.672 119.934 52.776 124.308 ; 
        RECT 52.24 119.934 52.344 124.308 ; 
        RECT 51.808 119.934 51.912 124.308 ; 
        RECT 51.376 119.934 51.48 124.308 ; 
        RECT 50.944 119.934 51.048 124.308 ; 
        RECT 50.512 119.934 50.616 124.308 ; 
        RECT 50.08 119.934 50.184 124.308 ; 
        RECT 49.648 119.934 49.752 124.308 ; 
        RECT 49.216 119.934 49.32 124.308 ; 
        RECT 48.784 119.934 48.888 124.308 ; 
        RECT 48.352 119.934 48.456 124.308 ; 
        RECT 47.92 119.934 48.024 124.308 ; 
        RECT 47.488 119.934 47.592 124.308 ; 
        RECT 47.056 119.934 47.16 124.308 ; 
        RECT 46.624 119.934 46.728 124.308 ; 
        RECT 46.192 119.934 46.296 124.308 ; 
        RECT 45.76 119.934 45.864 124.308 ; 
        RECT 45.328 119.934 45.432 124.308 ; 
        RECT 44.896 119.934 45 124.308 ; 
        RECT 44.464 119.934 44.568 124.308 ; 
        RECT 44.032 119.934 44.136 124.308 ; 
        RECT 43.6 119.934 43.704 124.308 ; 
        RECT 43.168 119.934 43.272 124.308 ; 
        RECT 42.736 119.934 42.84 124.308 ; 
        RECT 42.304 119.934 42.408 124.308 ; 
        RECT 41.872 119.934 41.976 124.308 ; 
        RECT 41.44 119.934 41.544 124.308 ; 
        RECT 41.008 119.934 41.112 124.308 ; 
        RECT 40.576 119.934 40.68 124.308 ; 
        RECT 40.144 119.934 40.248 124.308 ; 
        RECT 39.712 119.934 39.816 124.308 ; 
        RECT 39.28 119.934 39.384 124.308 ; 
        RECT 38.848 119.934 38.952 124.308 ; 
        RECT 38.416 119.934 38.52 124.308 ; 
        RECT 37.984 119.934 38.088 124.308 ; 
        RECT 37.552 119.934 37.656 124.308 ; 
        RECT 36.7 119.934 37.008 124.308 ; 
        RECT 29.128 119.934 29.436 124.308 ; 
        RECT 28.48 119.934 28.584 124.308 ; 
        RECT 28.048 119.934 28.152 124.308 ; 
        RECT 27.616 119.934 27.72 124.308 ; 
        RECT 27.184 119.934 27.288 124.308 ; 
        RECT 26.752 119.934 26.856 124.308 ; 
        RECT 26.32 119.934 26.424 124.308 ; 
        RECT 25.888 119.934 25.992 124.308 ; 
        RECT 25.456 119.934 25.56 124.308 ; 
        RECT 25.024 119.934 25.128 124.308 ; 
        RECT 24.592 119.934 24.696 124.308 ; 
        RECT 24.16 119.934 24.264 124.308 ; 
        RECT 23.728 119.934 23.832 124.308 ; 
        RECT 23.296 119.934 23.4 124.308 ; 
        RECT 22.864 119.934 22.968 124.308 ; 
        RECT 22.432 119.934 22.536 124.308 ; 
        RECT 22 119.934 22.104 124.308 ; 
        RECT 21.568 119.934 21.672 124.308 ; 
        RECT 21.136 119.934 21.24 124.308 ; 
        RECT 20.704 119.934 20.808 124.308 ; 
        RECT 20.272 119.934 20.376 124.308 ; 
        RECT 19.84 119.934 19.944 124.308 ; 
        RECT 19.408 119.934 19.512 124.308 ; 
        RECT 18.976 119.934 19.08 124.308 ; 
        RECT 18.544 119.934 18.648 124.308 ; 
        RECT 18.112 119.934 18.216 124.308 ; 
        RECT 17.68 119.934 17.784 124.308 ; 
        RECT 17.248 119.934 17.352 124.308 ; 
        RECT 16.816 119.934 16.92 124.308 ; 
        RECT 16.384 119.934 16.488 124.308 ; 
        RECT 15.952 119.934 16.056 124.308 ; 
        RECT 15.52 119.934 15.624 124.308 ; 
        RECT 15.088 119.934 15.192 124.308 ; 
        RECT 14.656 119.934 14.76 124.308 ; 
        RECT 14.224 119.934 14.328 124.308 ; 
        RECT 13.792 119.934 13.896 124.308 ; 
        RECT 13.36 119.934 13.464 124.308 ; 
        RECT 12.928 119.934 13.032 124.308 ; 
        RECT 12.496 119.934 12.6 124.308 ; 
        RECT 12.064 119.934 12.168 124.308 ; 
        RECT 11.632 119.934 11.736 124.308 ; 
        RECT 11.2 119.934 11.304 124.308 ; 
        RECT 10.768 119.934 10.872 124.308 ; 
        RECT 10.336 119.934 10.44 124.308 ; 
        RECT 9.904 119.934 10.008 124.308 ; 
        RECT 9.472 119.934 9.576 124.308 ; 
        RECT 9.04 119.934 9.144 124.308 ; 
        RECT 8.608 119.934 8.712 124.308 ; 
        RECT 8.176 119.934 8.28 124.308 ; 
        RECT 7.744 119.934 7.848 124.308 ; 
        RECT 7.312 119.934 7.416 124.308 ; 
        RECT 6.88 119.934 6.984 124.308 ; 
        RECT 6.448 119.934 6.552 124.308 ; 
        RECT 6.016 119.934 6.12 124.308 ; 
        RECT 5.584 119.934 5.688 124.308 ; 
        RECT 5.152 119.934 5.256 124.308 ; 
        RECT 4.72 119.934 4.824 124.308 ; 
        RECT 4.288 119.934 4.392 124.308 ; 
        RECT 3.856 119.934 3.96 124.308 ; 
        RECT 3.424 119.934 3.528 124.308 ; 
        RECT 2.992 119.934 3.096 124.308 ; 
        RECT 2.56 119.934 2.664 124.308 ; 
        RECT 2.128 119.934 2.232 124.308 ; 
        RECT 1.696 119.934 1.8 124.308 ; 
        RECT 1.264 119.934 1.368 124.308 ; 
        RECT 0.832 119.934 0.936 124.308 ; 
        RECT 0.02 119.934 0.36 124.308 ; 
        RECT 34.564 124.254 35.076 128.628 ; 
        RECT 34.508 126.916 35.076 128.206 ; 
        RECT 33.916 125.824 34.164 128.628 ; 
        RECT 33.86 127.062 34.164 127.676 ; 
        RECT 33.916 124.254 34.02 128.628 ; 
        RECT 33.916 124.738 34.076 125.696 ; 
        RECT 33.916 124.254 34.164 124.61 ; 
        RECT 32.728 126.056 33.552 128.628 ; 
        RECT 33.448 124.254 33.552 128.628 ; 
        RECT 32.728 127.164 33.608 128.196 ; 
        RECT 32.728 124.254 33.12 128.628 ; 
        RECT 31.06 124.254 31.392 128.628 ; 
        RECT 31.06 124.608 31.448 128.35 ; 
        RECT 65.776 124.254 66.116 128.628 ; 
        RECT 65.2 124.254 65.304 128.628 ; 
        RECT 64.768 124.254 64.872 128.628 ; 
        RECT 64.336 124.254 64.44 128.628 ; 
        RECT 63.904 124.254 64.008 128.628 ; 
        RECT 63.472 124.254 63.576 128.628 ; 
        RECT 63.04 124.254 63.144 128.628 ; 
        RECT 62.608 124.254 62.712 128.628 ; 
        RECT 62.176 124.254 62.28 128.628 ; 
        RECT 61.744 124.254 61.848 128.628 ; 
        RECT 61.312 124.254 61.416 128.628 ; 
        RECT 60.88 124.254 60.984 128.628 ; 
        RECT 60.448 124.254 60.552 128.628 ; 
        RECT 60.016 124.254 60.12 128.628 ; 
        RECT 59.584 124.254 59.688 128.628 ; 
        RECT 59.152 124.254 59.256 128.628 ; 
        RECT 58.72 124.254 58.824 128.628 ; 
        RECT 58.288 124.254 58.392 128.628 ; 
        RECT 57.856 124.254 57.96 128.628 ; 
        RECT 57.424 124.254 57.528 128.628 ; 
        RECT 56.992 124.254 57.096 128.628 ; 
        RECT 56.56 124.254 56.664 128.628 ; 
        RECT 56.128 124.254 56.232 128.628 ; 
        RECT 55.696 124.254 55.8 128.628 ; 
        RECT 55.264 124.254 55.368 128.628 ; 
        RECT 54.832 124.254 54.936 128.628 ; 
        RECT 54.4 124.254 54.504 128.628 ; 
        RECT 53.968 124.254 54.072 128.628 ; 
        RECT 53.536 124.254 53.64 128.628 ; 
        RECT 53.104 124.254 53.208 128.628 ; 
        RECT 52.672 124.254 52.776 128.628 ; 
        RECT 52.24 124.254 52.344 128.628 ; 
        RECT 51.808 124.254 51.912 128.628 ; 
        RECT 51.376 124.254 51.48 128.628 ; 
        RECT 50.944 124.254 51.048 128.628 ; 
        RECT 50.512 124.254 50.616 128.628 ; 
        RECT 50.08 124.254 50.184 128.628 ; 
        RECT 49.648 124.254 49.752 128.628 ; 
        RECT 49.216 124.254 49.32 128.628 ; 
        RECT 48.784 124.254 48.888 128.628 ; 
        RECT 48.352 124.254 48.456 128.628 ; 
        RECT 47.92 124.254 48.024 128.628 ; 
        RECT 47.488 124.254 47.592 128.628 ; 
        RECT 47.056 124.254 47.16 128.628 ; 
        RECT 46.624 124.254 46.728 128.628 ; 
        RECT 46.192 124.254 46.296 128.628 ; 
        RECT 45.76 124.254 45.864 128.628 ; 
        RECT 45.328 124.254 45.432 128.628 ; 
        RECT 44.896 124.254 45 128.628 ; 
        RECT 44.464 124.254 44.568 128.628 ; 
        RECT 44.032 124.254 44.136 128.628 ; 
        RECT 43.6 124.254 43.704 128.628 ; 
        RECT 43.168 124.254 43.272 128.628 ; 
        RECT 42.736 124.254 42.84 128.628 ; 
        RECT 42.304 124.254 42.408 128.628 ; 
        RECT 41.872 124.254 41.976 128.628 ; 
        RECT 41.44 124.254 41.544 128.628 ; 
        RECT 41.008 124.254 41.112 128.628 ; 
        RECT 40.576 124.254 40.68 128.628 ; 
        RECT 40.144 124.254 40.248 128.628 ; 
        RECT 39.712 124.254 39.816 128.628 ; 
        RECT 39.28 124.254 39.384 128.628 ; 
        RECT 38.848 124.254 38.952 128.628 ; 
        RECT 38.416 124.254 38.52 128.628 ; 
        RECT 37.984 124.254 38.088 128.628 ; 
        RECT 37.552 124.254 37.656 128.628 ; 
        RECT 36.7 124.254 37.008 128.628 ; 
        RECT 29.128 124.254 29.436 128.628 ; 
        RECT 28.48 124.254 28.584 128.628 ; 
        RECT 28.048 124.254 28.152 128.628 ; 
        RECT 27.616 124.254 27.72 128.628 ; 
        RECT 27.184 124.254 27.288 128.628 ; 
        RECT 26.752 124.254 26.856 128.628 ; 
        RECT 26.32 124.254 26.424 128.628 ; 
        RECT 25.888 124.254 25.992 128.628 ; 
        RECT 25.456 124.254 25.56 128.628 ; 
        RECT 25.024 124.254 25.128 128.628 ; 
        RECT 24.592 124.254 24.696 128.628 ; 
        RECT 24.16 124.254 24.264 128.628 ; 
        RECT 23.728 124.254 23.832 128.628 ; 
        RECT 23.296 124.254 23.4 128.628 ; 
        RECT 22.864 124.254 22.968 128.628 ; 
        RECT 22.432 124.254 22.536 128.628 ; 
        RECT 22 124.254 22.104 128.628 ; 
        RECT 21.568 124.254 21.672 128.628 ; 
        RECT 21.136 124.254 21.24 128.628 ; 
        RECT 20.704 124.254 20.808 128.628 ; 
        RECT 20.272 124.254 20.376 128.628 ; 
        RECT 19.84 124.254 19.944 128.628 ; 
        RECT 19.408 124.254 19.512 128.628 ; 
        RECT 18.976 124.254 19.08 128.628 ; 
        RECT 18.544 124.254 18.648 128.628 ; 
        RECT 18.112 124.254 18.216 128.628 ; 
        RECT 17.68 124.254 17.784 128.628 ; 
        RECT 17.248 124.254 17.352 128.628 ; 
        RECT 16.816 124.254 16.92 128.628 ; 
        RECT 16.384 124.254 16.488 128.628 ; 
        RECT 15.952 124.254 16.056 128.628 ; 
        RECT 15.52 124.254 15.624 128.628 ; 
        RECT 15.088 124.254 15.192 128.628 ; 
        RECT 14.656 124.254 14.76 128.628 ; 
        RECT 14.224 124.254 14.328 128.628 ; 
        RECT 13.792 124.254 13.896 128.628 ; 
        RECT 13.36 124.254 13.464 128.628 ; 
        RECT 12.928 124.254 13.032 128.628 ; 
        RECT 12.496 124.254 12.6 128.628 ; 
        RECT 12.064 124.254 12.168 128.628 ; 
        RECT 11.632 124.254 11.736 128.628 ; 
        RECT 11.2 124.254 11.304 128.628 ; 
        RECT 10.768 124.254 10.872 128.628 ; 
        RECT 10.336 124.254 10.44 128.628 ; 
        RECT 9.904 124.254 10.008 128.628 ; 
        RECT 9.472 124.254 9.576 128.628 ; 
        RECT 9.04 124.254 9.144 128.628 ; 
        RECT 8.608 124.254 8.712 128.628 ; 
        RECT 8.176 124.254 8.28 128.628 ; 
        RECT 7.744 124.254 7.848 128.628 ; 
        RECT 7.312 124.254 7.416 128.628 ; 
        RECT 6.88 124.254 6.984 128.628 ; 
        RECT 6.448 124.254 6.552 128.628 ; 
        RECT 6.016 124.254 6.12 128.628 ; 
        RECT 5.584 124.254 5.688 128.628 ; 
        RECT 5.152 124.254 5.256 128.628 ; 
        RECT 4.72 124.254 4.824 128.628 ; 
        RECT 4.288 124.254 4.392 128.628 ; 
        RECT 3.856 124.254 3.96 128.628 ; 
        RECT 3.424 124.254 3.528 128.628 ; 
        RECT 2.992 124.254 3.096 128.628 ; 
        RECT 2.56 124.254 2.664 128.628 ; 
        RECT 2.128 124.254 2.232 128.628 ; 
        RECT 1.696 124.254 1.8 128.628 ; 
        RECT 1.264 124.254 1.368 128.628 ; 
        RECT 0.832 124.254 0.936 128.628 ; 
        RECT 0.02 124.254 0.36 128.628 ; 
        RECT 34.564 128.574 35.076 132.948 ; 
        RECT 34.508 131.236 35.076 132.526 ; 
        RECT 33.916 130.144 34.164 132.948 ; 
        RECT 33.86 131.382 34.164 131.996 ; 
        RECT 33.916 128.574 34.02 132.948 ; 
        RECT 33.916 129.058 34.076 130.016 ; 
        RECT 33.916 128.574 34.164 128.93 ; 
        RECT 32.728 130.376 33.552 132.948 ; 
        RECT 33.448 128.574 33.552 132.948 ; 
        RECT 32.728 131.484 33.608 132.516 ; 
        RECT 32.728 128.574 33.12 132.948 ; 
        RECT 31.06 128.574 31.392 132.948 ; 
        RECT 31.06 128.928 31.448 132.67 ; 
        RECT 65.776 128.574 66.116 132.948 ; 
        RECT 65.2 128.574 65.304 132.948 ; 
        RECT 64.768 128.574 64.872 132.948 ; 
        RECT 64.336 128.574 64.44 132.948 ; 
        RECT 63.904 128.574 64.008 132.948 ; 
        RECT 63.472 128.574 63.576 132.948 ; 
        RECT 63.04 128.574 63.144 132.948 ; 
        RECT 62.608 128.574 62.712 132.948 ; 
        RECT 62.176 128.574 62.28 132.948 ; 
        RECT 61.744 128.574 61.848 132.948 ; 
        RECT 61.312 128.574 61.416 132.948 ; 
        RECT 60.88 128.574 60.984 132.948 ; 
        RECT 60.448 128.574 60.552 132.948 ; 
        RECT 60.016 128.574 60.12 132.948 ; 
        RECT 59.584 128.574 59.688 132.948 ; 
        RECT 59.152 128.574 59.256 132.948 ; 
        RECT 58.72 128.574 58.824 132.948 ; 
        RECT 58.288 128.574 58.392 132.948 ; 
        RECT 57.856 128.574 57.96 132.948 ; 
        RECT 57.424 128.574 57.528 132.948 ; 
        RECT 56.992 128.574 57.096 132.948 ; 
        RECT 56.56 128.574 56.664 132.948 ; 
        RECT 56.128 128.574 56.232 132.948 ; 
        RECT 55.696 128.574 55.8 132.948 ; 
        RECT 55.264 128.574 55.368 132.948 ; 
        RECT 54.832 128.574 54.936 132.948 ; 
        RECT 54.4 128.574 54.504 132.948 ; 
        RECT 53.968 128.574 54.072 132.948 ; 
        RECT 53.536 128.574 53.64 132.948 ; 
        RECT 53.104 128.574 53.208 132.948 ; 
        RECT 52.672 128.574 52.776 132.948 ; 
        RECT 52.24 128.574 52.344 132.948 ; 
        RECT 51.808 128.574 51.912 132.948 ; 
        RECT 51.376 128.574 51.48 132.948 ; 
        RECT 50.944 128.574 51.048 132.948 ; 
        RECT 50.512 128.574 50.616 132.948 ; 
        RECT 50.08 128.574 50.184 132.948 ; 
        RECT 49.648 128.574 49.752 132.948 ; 
        RECT 49.216 128.574 49.32 132.948 ; 
        RECT 48.784 128.574 48.888 132.948 ; 
        RECT 48.352 128.574 48.456 132.948 ; 
        RECT 47.92 128.574 48.024 132.948 ; 
        RECT 47.488 128.574 47.592 132.948 ; 
        RECT 47.056 128.574 47.16 132.948 ; 
        RECT 46.624 128.574 46.728 132.948 ; 
        RECT 46.192 128.574 46.296 132.948 ; 
        RECT 45.76 128.574 45.864 132.948 ; 
        RECT 45.328 128.574 45.432 132.948 ; 
        RECT 44.896 128.574 45 132.948 ; 
        RECT 44.464 128.574 44.568 132.948 ; 
        RECT 44.032 128.574 44.136 132.948 ; 
        RECT 43.6 128.574 43.704 132.948 ; 
        RECT 43.168 128.574 43.272 132.948 ; 
        RECT 42.736 128.574 42.84 132.948 ; 
        RECT 42.304 128.574 42.408 132.948 ; 
        RECT 41.872 128.574 41.976 132.948 ; 
        RECT 41.44 128.574 41.544 132.948 ; 
        RECT 41.008 128.574 41.112 132.948 ; 
        RECT 40.576 128.574 40.68 132.948 ; 
        RECT 40.144 128.574 40.248 132.948 ; 
        RECT 39.712 128.574 39.816 132.948 ; 
        RECT 39.28 128.574 39.384 132.948 ; 
        RECT 38.848 128.574 38.952 132.948 ; 
        RECT 38.416 128.574 38.52 132.948 ; 
        RECT 37.984 128.574 38.088 132.948 ; 
        RECT 37.552 128.574 37.656 132.948 ; 
        RECT 36.7 128.574 37.008 132.948 ; 
        RECT 29.128 128.574 29.436 132.948 ; 
        RECT 28.48 128.574 28.584 132.948 ; 
        RECT 28.048 128.574 28.152 132.948 ; 
        RECT 27.616 128.574 27.72 132.948 ; 
        RECT 27.184 128.574 27.288 132.948 ; 
        RECT 26.752 128.574 26.856 132.948 ; 
        RECT 26.32 128.574 26.424 132.948 ; 
        RECT 25.888 128.574 25.992 132.948 ; 
        RECT 25.456 128.574 25.56 132.948 ; 
        RECT 25.024 128.574 25.128 132.948 ; 
        RECT 24.592 128.574 24.696 132.948 ; 
        RECT 24.16 128.574 24.264 132.948 ; 
        RECT 23.728 128.574 23.832 132.948 ; 
        RECT 23.296 128.574 23.4 132.948 ; 
        RECT 22.864 128.574 22.968 132.948 ; 
        RECT 22.432 128.574 22.536 132.948 ; 
        RECT 22 128.574 22.104 132.948 ; 
        RECT 21.568 128.574 21.672 132.948 ; 
        RECT 21.136 128.574 21.24 132.948 ; 
        RECT 20.704 128.574 20.808 132.948 ; 
        RECT 20.272 128.574 20.376 132.948 ; 
        RECT 19.84 128.574 19.944 132.948 ; 
        RECT 19.408 128.574 19.512 132.948 ; 
        RECT 18.976 128.574 19.08 132.948 ; 
        RECT 18.544 128.574 18.648 132.948 ; 
        RECT 18.112 128.574 18.216 132.948 ; 
        RECT 17.68 128.574 17.784 132.948 ; 
        RECT 17.248 128.574 17.352 132.948 ; 
        RECT 16.816 128.574 16.92 132.948 ; 
        RECT 16.384 128.574 16.488 132.948 ; 
        RECT 15.952 128.574 16.056 132.948 ; 
        RECT 15.52 128.574 15.624 132.948 ; 
        RECT 15.088 128.574 15.192 132.948 ; 
        RECT 14.656 128.574 14.76 132.948 ; 
        RECT 14.224 128.574 14.328 132.948 ; 
        RECT 13.792 128.574 13.896 132.948 ; 
        RECT 13.36 128.574 13.464 132.948 ; 
        RECT 12.928 128.574 13.032 132.948 ; 
        RECT 12.496 128.574 12.6 132.948 ; 
        RECT 12.064 128.574 12.168 132.948 ; 
        RECT 11.632 128.574 11.736 132.948 ; 
        RECT 11.2 128.574 11.304 132.948 ; 
        RECT 10.768 128.574 10.872 132.948 ; 
        RECT 10.336 128.574 10.44 132.948 ; 
        RECT 9.904 128.574 10.008 132.948 ; 
        RECT 9.472 128.574 9.576 132.948 ; 
        RECT 9.04 128.574 9.144 132.948 ; 
        RECT 8.608 128.574 8.712 132.948 ; 
        RECT 8.176 128.574 8.28 132.948 ; 
        RECT 7.744 128.574 7.848 132.948 ; 
        RECT 7.312 128.574 7.416 132.948 ; 
        RECT 6.88 128.574 6.984 132.948 ; 
        RECT 6.448 128.574 6.552 132.948 ; 
        RECT 6.016 128.574 6.12 132.948 ; 
        RECT 5.584 128.574 5.688 132.948 ; 
        RECT 5.152 128.574 5.256 132.948 ; 
        RECT 4.72 128.574 4.824 132.948 ; 
        RECT 4.288 128.574 4.392 132.948 ; 
        RECT 3.856 128.574 3.96 132.948 ; 
        RECT 3.424 128.574 3.528 132.948 ; 
        RECT 2.992 128.574 3.096 132.948 ; 
        RECT 2.56 128.574 2.664 132.948 ; 
        RECT 2.128 128.574 2.232 132.948 ; 
        RECT 1.696 128.574 1.8 132.948 ; 
        RECT 1.264 128.574 1.368 132.948 ; 
        RECT 0.832 128.574 0.936 132.948 ; 
        RECT 0.02 128.574 0.36 132.948 ; 
        RECT 34.564 132.894 35.076 137.268 ; 
        RECT 34.508 135.556 35.076 136.846 ; 
        RECT 33.916 134.464 34.164 137.268 ; 
        RECT 33.86 135.702 34.164 136.316 ; 
        RECT 33.916 132.894 34.02 137.268 ; 
        RECT 33.916 133.378 34.076 134.336 ; 
        RECT 33.916 132.894 34.164 133.25 ; 
        RECT 32.728 134.696 33.552 137.268 ; 
        RECT 33.448 132.894 33.552 137.268 ; 
        RECT 32.728 135.804 33.608 136.836 ; 
        RECT 32.728 132.894 33.12 137.268 ; 
        RECT 31.06 132.894 31.392 137.268 ; 
        RECT 31.06 133.248 31.448 136.99 ; 
        RECT 65.776 132.894 66.116 137.268 ; 
        RECT 65.2 132.894 65.304 137.268 ; 
        RECT 64.768 132.894 64.872 137.268 ; 
        RECT 64.336 132.894 64.44 137.268 ; 
        RECT 63.904 132.894 64.008 137.268 ; 
        RECT 63.472 132.894 63.576 137.268 ; 
        RECT 63.04 132.894 63.144 137.268 ; 
        RECT 62.608 132.894 62.712 137.268 ; 
        RECT 62.176 132.894 62.28 137.268 ; 
        RECT 61.744 132.894 61.848 137.268 ; 
        RECT 61.312 132.894 61.416 137.268 ; 
        RECT 60.88 132.894 60.984 137.268 ; 
        RECT 60.448 132.894 60.552 137.268 ; 
        RECT 60.016 132.894 60.12 137.268 ; 
        RECT 59.584 132.894 59.688 137.268 ; 
        RECT 59.152 132.894 59.256 137.268 ; 
        RECT 58.72 132.894 58.824 137.268 ; 
        RECT 58.288 132.894 58.392 137.268 ; 
        RECT 57.856 132.894 57.96 137.268 ; 
        RECT 57.424 132.894 57.528 137.268 ; 
        RECT 56.992 132.894 57.096 137.268 ; 
        RECT 56.56 132.894 56.664 137.268 ; 
        RECT 56.128 132.894 56.232 137.268 ; 
        RECT 55.696 132.894 55.8 137.268 ; 
        RECT 55.264 132.894 55.368 137.268 ; 
        RECT 54.832 132.894 54.936 137.268 ; 
        RECT 54.4 132.894 54.504 137.268 ; 
        RECT 53.968 132.894 54.072 137.268 ; 
        RECT 53.536 132.894 53.64 137.268 ; 
        RECT 53.104 132.894 53.208 137.268 ; 
        RECT 52.672 132.894 52.776 137.268 ; 
        RECT 52.24 132.894 52.344 137.268 ; 
        RECT 51.808 132.894 51.912 137.268 ; 
        RECT 51.376 132.894 51.48 137.268 ; 
        RECT 50.944 132.894 51.048 137.268 ; 
        RECT 50.512 132.894 50.616 137.268 ; 
        RECT 50.08 132.894 50.184 137.268 ; 
        RECT 49.648 132.894 49.752 137.268 ; 
        RECT 49.216 132.894 49.32 137.268 ; 
        RECT 48.784 132.894 48.888 137.268 ; 
        RECT 48.352 132.894 48.456 137.268 ; 
        RECT 47.92 132.894 48.024 137.268 ; 
        RECT 47.488 132.894 47.592 137.268 ; 
        RECT 47.056 132.894 47.16 137.268 ; 
        RECT 46.624 132.894 46.728 137.268 ; 
        RECT 46.192 132.894 46.296 137.268 ; 
        RECT 45.76 132.894 45.864 137.268 ; 
        RECT 45.328 132.894 45.432 137.268 ; 
        RECT 44.896 132.894 45 137.268 ; 
        RECT 44.464 132.894 44.568 137.268 ; 
        RECT 44.032 132.894 44.136 137.268 ; 
        RECT 43.6 132.894 43.704 137.268 ; 
        RECT 43.168 132.894 43.272 137.268 ; 
        RECT 42.736 132.894 42.84 137.268 ; 
        RECT 42.304 132.894 42.408 137.268 ; 
        RECT 41.872 132.894 41.976 137.268 ; 
        RECT 41.44 132.894 41.544 137.268 ; 
        RECT 41.008 132.894 41.112 137.268 ; 
        RECT 40.576 132.894 40.68 137.268 ; 
        RECT 40.144 132.894 40.248 137.268 ; 
        RECT 39.712 132.894 39.816 137.268 ; 
        RECT 39.28 132.894 39.384 137.268 ; 
        RECT 38.848 132.894 38.952 137.268 ; 
        RECT 38.416 132.894 38.52 137.268 ; 
        RECT 37.984 132.894 38.088 137.268 ; 
        RECT 37.552 132.894 37.656 137.268 ; 
        RECT 36.7 132.894 37.008 137.268 ; 
        RECT 29.128 132.894 29.436 137.268 ; 
        RECT 28.48 132.894 28.584 137.268 ; 
        RECT 28.048 132.894 28.152 137.268 ; 
        RECT 27.616 132.894 27.72 137.268 ; 
        RECT 27.184 132.894 27.288 137.268 ; 
        RECT 26.752 132.894 26.856 137.268 ; 
        RECT 26.32 132.894 26.424 137.268 ; 
        RECT 25.888 132.894 25.992 137.268 ; 
        RECT 25.456 132.894 25.56 137.268 ; 
        RECT 25.024 132.894 25.128 137.268 ; 
        RECT 24.592 132.894 24.696 137.268 ; 
        RECT 24.16 132.894 24.264 137.268 ; 
        RECT 23.728 132.894 23.832 137.268 ; 
        RECT 23.296 132.894 23.4 137.268 ; 
        RECT 22.864 132.894 22.968 137.268 ; 
        RECT 22.432 132.894 22.536 137.268 ; 
        RECT 22 132.894 22.104 137.268 ; 
        RECT 21.568 132.894 21.672 137.268 ; 
        RECT 21.136 132.894 21.24 137.268 ; 
        RECT 20.704 132.894 20.808 137.268 ; 
        RECT 20.272 132.894 20.376 137.268 ; 
        RECT 19.84 132.894 19.944 137.268 ; 
        RECT 19.408 132.894 19.512 137.268 ; 
        RECT 18.976 132.894 19.08 137.268 ; 
        RECT 18.544 132.894 18.648 137.268 ; 
        RECT 18.112 132.894 18.216 137.268 ; 
        RECT 17.68 132.894 17.784 137.268 ; 
        RECT 17.248 132.894 17.352 137.268 ; 
        RECT 16.816 132.894 16.92 137.268 ; 
        RECT 16.384 132.894 16.488 137.268 ; 
        RECT 15.952 132.894 16.056 137.268 ; 
        RECT 15.52 132.894 15.624 137.268 ; 
        RECT 15.088 132.894 15.192 137.268 ; 
        RECT 14.656 132.894 14.76 137.268 ; 
        RECT 14.224 132.894 14.328 137.268 ; 
        RECT 13.792 132.894 13.896 137.268 ; 
        RECT 13.36 132.894 13.464 137.268 ; 
        RECT 12.928 132.894 13.032 137.268 ; 
        RECT 12.496 132.894 12.6 137.268 ; 
        RECT 12.064 132.894 12.168 137.268 ; 
        RECT 11.632 132.894 11.736 137.268 ; 
        RECT 11.2 132.894 11.304 137.268 ; 
        RECT 10.768 132.894 10.872 137.268 ; 
        RECT 10.336 132.894 10.44 137.268 ; 
        RECT 9.904 132.894 10.008 137.268 ; 
        RECT 9.472 132.894 9.576 137.268 ; 
        RECT 9.04 132.894 9.144 137.268 ; 
        RECT 8.608 132.894 8.712 137.268 ; 
        RECT 8.176 132.894 8.28 137.268 ; 
        RECT 7.744 132.894 7.848 137.268 ; 
        RECT 7.312 132.894 7.416 137.268 ; 
        RECT 6.88 132.894 6.984 137.268 ; 
        RECT 6.448 132.894 6.552 137.268 ; 
        RECT 6.016 132.894 6.12 137.268 ; 
        RECT 5.584 132.894 5.688 137.268 ; 
        RECT 5.152 132.894 5.256 137.268 ; 
        RECT 4.72 132.894 4.824 137.268 ; 
        RECT 4.288 132.894 4.392 137.268 ; 
        RECT 3.856 132.894 3.96 137.268 ; 
        RECT 3.424 132.894 3.528 137.268 ; 
        RECT 2.992 132.894 3.096 137.268 ; 
        RECT 2.56 132.894 2.664 137.268 ; 
        RECT 2.128 132.894 2.232 137.268 ; 
        RECT 1.696 132.894 1.8 137.268 ; 
        RECT 1.264 132.894 1.368 137.268 ; 
        RECT 0.832 132.894 0.936 137.268 ; 
        RECT 0.02 132.894 0.36 137.268 ; 
        RECT 34.564 137.214 35.076 141.588 ; 
        RECT 34.508 139.876 35.076 141.166 ; 
        RECT 33.916 138.784 34.164 141.588 ; 
        RECT 33.86 140.022 34.164 140.636 ; 
        RECT 33.916 137.214 34.02 141.588 ; 
        RECT 33.916 137.698 34.076 138.656 ; 
        RECT 33.916 137.214 34.164 137.57 ; 
        RECT 32.728 139.016 33.552 141.588 ; 
        RECT 33.448 137.214 33.552 141.588 ; 
        RECT 32.728 140.124 33.608 141.156 ; 
        RECT 32.728 137.214 33.12 141.588 ; 
        RECT 31.06 137.214 31.392 141.588 ; 
        RECT 31.06 137.568 31.448 141.31 ; 
        RECT 65.776 137.214 66.116 141.588 ; 
        RECT 65.2 137.214 65.304 141.588 ; 
        RECT 64.768 137.214 64.872 141.588 ; 
        RECT 64.336 137.214 64.44 141.588 ; 
        RECT 63.904 137.214 64.008 141.588 ; 
        RECT 63.472 137.214 63.576 141.588 ; 
        RECT 63.04 137.214 63.144 141.588 ; 
        RECT 62.608 137.214 62.712 141.588 ; 
        RECT 62.176 137.214 62.28 141.588 ; 
        RECT 61.744 137.214 61.848 141.588 ; 
        RECT 61.312 137.214 61.416 141.588 ; 
        RECT 60.88 137.214 60.984 141.588 ; 
        RECT 60.448 137.214 60.552 141.588 ; 
        RECT 60.016 137.214 60.12 141.588 ; 
        RECT 59.584 137.214 59.688 141.588 ; 
        RECT 59.152 137.214 59.256 141.588 ; 
        RECT 58.72 137.214 58.824 141.588 ; 
        RECT 58.288 137.214 58.392 141.588 ; 
        RECT 57.856 137.214 57.96 141.588 ; 
        RECT 57.424 137.214 57.528 141.588 ; 
        RECT 56.992 137.214 57.096 141.588 ; 
        RECT 56.56 137.214 56.664 141.588 ; 
        RECT 56.128 137.214 56.232 141.588 ; 
        RECT 55.696 137.214 55.8 141.588 ; 
        RECT 55.264 137.214 55.368 141.588 ; 
        RECT 54.832 137.214 54.936 141.588 ; 
        RECT 54.4 137.214 54.504 141.588 ; 
        RECT 53.968 137.214 54.072 141.588 ; 
        RECT 53.536 137.214 53.64 141.588 ; 
        RECT 53.104 137.214 53.208 141.588 ; 
        RECT 52.672 137.214 52.776 141.588 ; 
        RECT 52.24 137.214 52.344 141.588 ; 
        RECT 51.808 137.214 51.912 141.588 ; 
        RECT 51.376 137.214 51.48 141.588 ; 
        RECT 50.944 137.214 51.048 141.588 ; 
        RECT 50.512 137.214 50.616 141.588 ; 
        RECT 50.08 137.214 50.184 141.588 ; 
        RECT 49.648 137.214 49.752 141.588 ; 
        RECT 49.216 137.214 49.32 141.588 ; 
        RECT 48.784 137.214 48.888 141.588 ; 
        RECT 48.352 137.214 48.456 141.588 ; 
        RECT 47.92 137.214 48.024 141.588 ; 
        RECT 47.488 137.214 47.592 141.588 ; 
        RECT 47.056 137.214 47.16 141.588 ; 
        RECT 46.624 137.214 46.728 141.588 ; 
        RECT 46.192 137.214 46.296 141.588 ; 
        RECT 45.76 137.214 45.864 141.588 ; 
        RECT 45.328 137.214 45.432 141.588 ; 
        RECT 44.896 137.214 45 141.588 ; 
        RECT 44.464 137.214 44.568 141.588 ; 
        RECT 44.032 137.214 44.136 141.588 ; 
        RECT 43.6 137.214 43.704 141.588 ; 
        RECT 43.168 137.214 43.272 141.588 ; 
        RECT 42.736 137.214 42.84 141.588 ; 
        RECT 42.304 137.214 42.408 141.588 ; 
        RECT 41.872 137.214 41.976 141.588 ; 
        RECT 41.44 137.214 41.544 141.588 ; 
        RECT 41.008 137.214 41.112 141.588 ; 
        RECT 40.576 137.214 40.68 141.588 ; 
        RECT 40.144 137.214 40.248 141.588 ; 
        RECT 39.712 137.214 39.816 141.588 ; 
        RECT 39.28 137.214 39.384 141.588 ; 
        RECT 38.848 137.214 38.952 141.588 ; 
        RECT 38.416 137.214 38.52 141.588 ; 
        RECT 37.984 137.214 38.088 141.588 ; 
        RECT 37.552 137.214 37.656 141.588 ; 
        RECT 36.7 137.214 37.008 141.588 ; 
        RECT 29.128 137.214 29.436 141.588 ; 
        RECT 28.48 137.214 28.584 141.588 ; 
        RECT 28.048 137.214 28.152 141.588 ; 
        RECT 27.616 137.214 27.72 141.588 ; 
        RECT 27.184 137.214 27.288 141.588 ; 
        RECT 26.752 137.214 26.856 141.588 ; 
        RECT 26.32 137.214 26.424 141.588 ; 
        RECT 25.888 137.214 25.992 141.588 ; 
        RECT 25.456 137.214 25.56 141.588 ; 
        RECT 25.024 137.214 25.128 141.588 ; 
        RECT 24.592 137.214 24.696 141.588 ; 
        RECT 24.16 137.214 24.264 141.588 ; 
        RECT 23.728 137.214 23.832 141.588 ; 
        RECT 23.296 137.214 23.4 141.588 ; 
        RECT 22.864 137.214 22.968 141.588 ; 
        RECT 22.432 137.214 22.536 141.588 ; 
        RECT 22 137.214 22.104 141.588 ; 
        RECT 21.568 137.214 21.672 141.588 ; 
        RECT 21.136 137.214 21.24 141.588 ; 
        RECT 20.704 137.214 20.808 141.588 ; 
        RECT 20.272 137.214 20.376 141.588 ; 
        RECT 19.84 137.214 19.944 141.588 ; 
        RECT 19.408 137.214 19.512 141.588 ; 
        RECT 18.976 137.214 19.08 141.588 ; 
        RECT 18.544 137.214 18.648 141.588 ; 
        RECT 18.112 137.214 18.216 141.588 ; 
        RECT 17.68 137.214 17.784 141.588 ; 
        RECT 17.248 137.214 17.352 141.588 ; 
        RECT 16.816 137.214 16.92 141.588 ; 
        RECT 16.384 137.214 16.488 141.588 ; 
        RECT 15.952 137.214 16.056 141.588 ; 
        RECT 15.52 137.214 15.624 141.588 ; 
        RECT 15.088 137.214 15.192 141.588 ; 
        RECT 14.656 137.214 14.76 141.588 ; 
        RECT 14.224 137.214 14.328 141.588 ; 
        RECT 13.792 137.214 13.896 141.588 ; 
        RECT 13.36 137.214 13.464 141.588 ; 
        RECT 12.928 137.214 13.032 141.588 ; 
        RECT 12.496 137.214 12.6 141.588 ; 
        RECT 12.064 137.214 12.168 141.588 ; 
        RECT 11.632 137.214 11.736 141.588 ; 
        RECT 11.2 137.214 11.304 141.588 ; 
        RECT 10.768 137.214 10.872 141.588 ; 
        RECT 10.336 137.214 10.44 141.588 ; 
        RECT 9.904 137.214 10.008 141.588 ; 
        RECT 9.472 137.214 9.576 141.588 ; 
        RECT 9.04 137.214 9.144 141.588 ; 
        RECT 8.608 137.214 8.712 141.588 ; 
        RECT 8.176 137.214 8.28 141.588 ; 
        RECT 7.744 137.214 7.848 141.588 ; 
        RECT 7.312 137.214 7.416 141.588 ; 
        RECT 6.88 137.214 6.984 141.588 ; 
        RECT 6.448 137.214 6.552 141.588 ; 
        RECT 6.016 137.214 6.12 141.588 ; 
        RECT 5.584 137.214 5.688 141.588 ; 
        RECT 5.152 137.214 5.256 141.588 ; 
        RECT 4.72 137.214 4.824 141.588 ; 
        RECT 4.288 137.214 4.392 141.588 ; 
        RECT 3.856 137.214 3.96 141.588 ; 
        RECT 3.424 137.214 3.528 141.588 ; 
        RECT 2.992 137.214 3.096 141.588 ; 
        RECT 2.56 137.214 2.664 141.588 ; 
        RECT 2.128 137.214 2.232 141.588 ; 
        RECT 1.696 137.214 1.8 141.588 ; 
        RECT 1.264 137.214 1.368 141.588 ; 
        RECT 0.832 137.214 0.936 141.588 ; 
        RECT 0.02 137.214 0.36 141.588 ; 
        RECT 34.564 141.534 35.076 145.908 ; 
        RECT 34.508 144.196 35.076 145.486 ; 
        RECT 33.916 143.104 34.164 145.908 ; 
        RECT 33.86 144.342 34.164 144.956 ; 
        RECT 33.916 141.534 34.02 145.908 ; 
        RECT 33.916 142.018 34.076 142.976 ; 
        RECT 33.916 141.534 34.164 141.89 ; 
        RECT 32.728 143.336 33.552 145.908 ; 
        RECT 33.448 141.534 33.552 145.908 ; 
        RECT 32.728 144.444 33.608 145.476 ; 
        RECT 32.728 141.534 33.12 145.908 ; 
        RECT 31.06 141.534 31.392 145.908 ; 
        RECT 31.06 141.888 31.448 145.63 ; 
        RECT 65.776 141.534 66.116 145.908 ; 
        RECT 65.2 141.534 65.304 145.908 ; 
        RECT 64.768 141.534 64.872 145.908 ; 
        RECT 64.336 141.534 64.44 145.908 ; 
        RECT 63.904 141.534 64.008 145.908 ; 
        RECT 63.472 141.534 63.576 145.908 ; 
        RECT 63.04 141.534 63.144 145.908 ; 
        RECT 62.608 141.534 62.712 145.908 ; 
        RECT 62.176 141.534 62.28 145.908 ; 
        RECT 61.744 141.534 61.848 145.908 ; 
        RECT 61.312 141.534 61.416 145.908 ; 
        RECT 60.88 141.534 60.984 145.908 ; 
        RECT 60.448 141.534 60.552 145.908 ; 
        RECT 60.016 141.534 60.12 145.908 ; 
        RECT 59.584 141.534 59.688 145.908 ; 
        RECT 59.152 141.534 59.256 145.908 ; 
        RECT 58.72 141.534 58.824 145.908 ; 
        RECT 58.288 141.534 58.392 145.908 ; 
        RECT 57.856 141.534 57.96 145.908 ; 
        RECT 57.424 141.534 57.528 145.908 ; 
        RECT 56.992 141.534 57.096 145.908 ; 
        RECT 56.56 141.534 56.664 145.908 ; 
        RECT 56.128 141.534 56.232 145.908 ; 
        RECT 55.696 141.534 55.8 145.908 ; 
        RECT 55.264 141.534 55.368 145.908 ; 
        RECT 54.832 141.534 54.936 145.908 ; 
        RECT 54.4 141.534 54.504 145.908 ; 
        RECT 53.968 141.534 54.072 145.908 ; 
        RECT 53.536 141.534 53.64 145.908 ; 
        RECT 53.104 141.534 53.208 145.908 ; 
        RECT 52.672 141.534 52.776 145.908 ; 
        RECT 52.24 141.534 52.344 145.908 ; 
        RECT 51.808 141.534 51.912 145.908 ; 
        RECT 51.376 141.534 51.48 145.908 ; 
        RECT 50.944 141.534 51.048 145.908 ; 
        RECT 50.512 141.534 50.616 145.908 ; 
        RECT 50.08 141.534 50.184 145.908 ; 
        RECT 49.648 141.534 49.752 145.908 ; 
        RECT 49.216 141.534 49.32 145.908 ; 
        RECT 48.784 141.534 48.888 145.908 ; 
        RECT 48.352 141.534 48.456 145.908 ; 
        RECT 47.92 141.534 48.024 145.908 ; 
        RECT 47.488 141.534 47.592 145.908 ; 
        RECT 47.056 141.534 47.16 145.908 ; 
        RECT 46.624 141.534 46.728 145.908 ; 
        RECT 46.192 141.534 46.296 145.908 ; 
        RECT 45.76 141.534 45.864 145.908 ; 
        RECT 45.328 141.534 45.432 145.908 ; 
        RECT 44.896 141.534 45 145.908 ; 
        RECT 44.464 141.534 44.568 145.908 ; 
        RECT 44.032 141.534 44.136 145.908 ; 
        RECT 43.6 141.534 43.704 145.908 ; 
        RECT 43.168 141.534 43.272 145.908 ; 
        RECT 42.736 141.534 42.84 145.908 ; 
        RECT 42.304 141.534 42.408 145.908 ; 
        RECT 41.872 141.534 41.976 145.908 ; 
        RECT 41.44 141.534 41.544 145.908 ; 
        RECT 41.008 141.534 41.112 145.908 ; 
        RECT 40.576 141.534 40.68 145.908 ; 
        RECT 40.144 141.534 40.248 145.908 ; 
        RECT 39.712 141.534 39.816 145.908 ; 
        RECT 39.28 141.534 39.384 145.908 ; 
        RECT 38.848 141.534 38.952 145.908 ; 
        RECT 38.416 141.534 38.52 145.908 ; 
        RECT 37.984 141.534 38.088 145.908 ; 
        RECT 37.552 141.534 37.656 145.908 ; 
        RECT 36.7 141.534 37.008 145.908 ; 
        RECT 29.128 141.534 29.436 145.908 ; 
        RECT 28.48 141.534 28.584 145.908 ; 
        RECT 28.048 141.534 28.152 145.908 ; 
        RECT 27.616 141.534 27.72 145.908 ; 
        RECT 27.184 141.534 27.288 145.908 ; 
        RECT 26.752 141.534 26.856 145.908 ; 
        RECT 26.32 141.534 26.424 145.908 ; 
        RECT 25.888 141.534 25.992 145.908 ; 
        RECT 25.456 141.534 25.56 145.908 ; 
        RECT 25.024 141.534 25.128 145.908 ; 
        RECT 24.592 141.534 24.696 145.908 ; 
        RECT 24.16 141.534 24.264 145.908 ; 
        RECT 23.728 141.534 23.832 145.908 ; 
        RECT 23.296 141.534 23.4 145.908 ; 
        RECT 22.864 141.534 22.968 145.908 ; 
        RECT 22.432 141.534 22.536 145.908 ; 
        RECT 22 141.534 22.104 145.908 ; 
        RECT 21.568 141.534 21.672 145.908 ; 
        RECT 21.136 141.534 21.24 145.908 ; 
        RECT 20.704 141.534 20.808 145.908 ; 
        RECT 20.272 141.534 20.376 145.908 ; 
        RECT 19.84 141.534 19.944 145.908 ; 
        RECT 19.408 141.534 19.512 145.908 ; 
        RECT 18.976 141.534 19.08 145.908 ; 
        RECT 18.544 141.534 18.648 145.908 ; 
        RECT 18.112 141.534 18.216 145.908 ; 
        RECT 17.68 141.534 17.784 145.908 ; 
        RECT 17.248 141.534 17.352 145.908 ; 
        RECT 16.816 141.534 16.92 145.908 ; 
        RECT 16.384 141.534 16.488 145.908 ; 
        RECT 15.952 141.534 16.056 145.908 ; 
        RECT 15.52 141.534 15.624 145.908 ; 
        RECT 15.088 141.534 15.192 145.908 ; 
        RECT 14.656 141.534 14.76 145.908 ; 
        RECT 14.224 141.534 14.328 145.908 ; 
        RECT 13.792 141.534 13.896 145.908 ; 
        RECT 13.36 141.534 13.464 145.908 ; 
        RECT 12.928 141.534 13.032 145.908 ; 
        RECT 12.496 141.534 12.6 145.908 ; 
        RECT 12.064 141.534 12.168 145.908 ; 
        RECT 11.632 141.534 11.736 145.908 ; 
        RECT 11.2 141.534 11.304 145.908 ; 
        RECT 10.768 141.534 10.872 145.908 ; 
        RECT 10.336 141.534 10.44 145.908 ; 
        RECT 9.904 141.534 10.008 145.908 ; 
        RECT 9.472 141.534 9.576 145.908 ; 
        RECT 9.04 141.534 9.144 145.908 ; 
        RECT 8.608 141.534 8.712 145.908 ; 
        RECT 8.176 141.534 8.28 145.908 ; 
        RECT 7.744 141.534 7.848 145.908 ; 
        RECT 7.312 141.534 7.416 145.908 ; 
        RECT 6.88 141.534 6.984 145.908 ; 
        RECT 6.448 141.534 6.552 145.908 ; 
        RECT 6.016 141.534 6.12 145.908 ; 
        RECT 5.584 141.534 5.688 145.908 ; 
        RECT 5.152 141.534 5.256 145.908 ; 
        RECT 4.72 141.534 4.824 145.908 ; 
        RECT 4.288 141.534 4.392 145.908 ; 
        RECT 3.856 141.534 3.96 145.908 ; 
        RECT 3.424 141.534 3.528 145.908 ; 
        RECT 2.992 141.534 3.096 145.908 ; 
        RECT 2.56 141.534 2.664 145.908 ; 
        RECT 2.128 141.534 2.232 145.908 ; 
        RECT 1.696 141.534 1.8 145.908 ; 
        RECT 1.264 141.534 1.368 145.908 ; 
        RECT 0.832 141.534 0.936 145.908 ; 
        RECT 0.02 141.534 0.36 145.908 ; 
        RECT 34.564 145.854 35.076 150.228 ; 
        RECT 34.508 148.516 35.076 149.806 ; 
        RECT 33.916 147.424 34.164 150.228 ; 
        RECT 33.86 148.662 34.164 149.276 ; 
        RECT 33.916 145.854 34.02 150.228 ; 
        RECT 33.916 146.338 34.076 147.296 ; 
        RECT 33.916 145.854 34.164 146.21 ; 
        RECT 32.728 147.656 33.552 150.228 ; 
        RECT 33.448 145.854 33.552 150.228 ; 
        RECT 32.728 148.764 33.608 149.796 ; 
        RECT 32.728 145.854 33.12 150.228 ; 
        RECT 31.06 145.854 31.392 150.228 ; 
        RECT 31.06 146.208 31.448 149.95 ; 
        RECT 65.776 145.854 66.116 150.228 ; 
        RECT 65.2 145.854 65.304 150.228 ; 
        RECT 64.768 145.854 64.872 150.228 ; 
        RECT 64.336 145.854 64.44 150.228 ; 
        RECT 63.904 145.854 64.008 150.228 ; 
        RECT 63.472 145.854 63.576 150.228 ; 
        RECT 63.04 145.854 63.144 150.228 ; 
        RECT 62.608 145.854 62.712 150.228 ; 
        RECT 62.176 145.854 62.28 150.228 ; 
        RECT 61.744 145.854 61.848 150.228 ; 
        RECT 61.312 145.854 61.416 150.228 ; 
        RECT 60.88 145.854 60.984 150.228 ; 
        RECT 60.448 145.854 60.552 150.228 ; 
        RECT 60.016 145.854 60.12 150.228 ; 
        RECT 59.584 145.854 59.688 150.228 ; 
        RECT 59.152 145.854 59.256 150.228 ; 
        RECT 58.72 145.854 58.824 150.228 ; 
        RECT 58.288 145.854 58.392 150.228 ; 
        RECT 57.856 145.854 57.96 150.228 ; 
        RECT 57.424 145.854 57.528 150.228 ; 
        RECT 56.992 145.854 57.096 150.228 ; 
        RECT 56.56 145.854 56.664 150.228 ; 
        RECT 56.128 145.854 56.232 150.228 ; 
        RECT 55.696 145.854 55.8 150.228 ; 
        RECT 55.264 145.854 55.368 150.228 ; 
        RECT 54.832 145.854 54.936 150.228 ; 
        RECT 54.4 145.854 54.504 150.228 ; 
        RECT 53.968 145.854 54.072 150.228 ; 
        RECT 53.536 145.854 53.64 150.228 ; 
        RECT 53.104 145.854 53.208 150.228 ; 
        RECT 52.672 145.854 52.776 150.228 ; 
        RECT 52.24 145.854 52.344 150.228 ; 
        RECT 51.808 145.854 51.912 150.228 ; 
        RECT 51.376 145.854 51.48 150.228 ; 
        RECT 50.944 145.854 51.048 150.228 ; 
        RECT 50.512 145.854 50.616 150.228 ; 
        RECT 50.08 145.854 50.184 150.228 ; 
        RECT 49.648 145.854 49.752 150.228 ; 
        RECT 49.216 145.854 49.32 150.228 ; 
        RECT 48.784 145.854 48.888 150.228 ; 
        RECT 48.352 145.854 48.456 150.228 ; 
        RECT 47.92 145.854 48.024 150.228 ; 
        RECT 47.488 145.854 47.592 150.228 ; 
        RECT 47.056 145.854 47.16 150.228 ; 
        RECT 46.624 145.854 46.728 150.228 ; 
        RECT 46.192 145.854 46.296 150.228 ; 
        RECT 45.76 145.854 45.864 150.228 ; 
        RECT 45.328 145.854 45.432 150.228 ; 
        RECT 44.896 145.854 45 150.228 ; 
        RECT 44.464 145.854 44.568 150.228 ; 
        RECT 44.032 145.854 44.136 150.228 ; 
        RECT 43.6 145.854 43.704 150.228 ; 
        RECT 43.168 145.854 43.272 150.228 ; 
        RECT 42.736 145.854 42.84 150.228 ; 
        RECT 42.304 145.854 42.408 150.228 ; 
        RECT 41.872 145.854 41.976 150.228 ; 
        RECT 41.44 145.854 41.544 150.228 ; 
        RECT 41.008 145.854 41.112 150.228 ; 
        RECT 40.576 145.854 40.68 150.228 ; 
        RECT 40.144 145.854 40.248 150.228 ; 
        RECT 39.712 145.854 39.816 150.228 ; 
        RECT 39.28 145.854 39.384 150.228 ; 
        RECT 38.848 145.854 38.952 150.228 ; 
        RECT 38.416 145.854 38.52 150.228 ; 
        RECT 37.984 145.854 38.088 150.228 ; 
        RECT 37.552 145.854 37.656 150.228 ; 
        RECT 36.7 145.854 37.008 150.228 ; 
        RECT 29.128 145.854 29.436 150.228 ; 
        RECT 28.48 145.854 28.584 150.228 ; 
        RECT 28.048 145.854 28.152 150.228 ; 
        RECT 27.616 145.854 27.72 150.228 ; 
        RECT 27.184 145.854 27.288 150.228 ; 
        RECT 26.752 145.854 26.856 150.228 ; 
        RECT 26.32 145.854 26.424 150.228 ; 
        RECT 25.888 145.854 25.992 150.228 ; 
        RECT 25.456 145.854 25.56 150.228 ; 
        RECT 25.024 145.854 25.128 150.228 ; 
        RECT 24.592 145.854 24.696 150.228 ; 
        RECT 24.16 145.854 24.264 150.228 ; 
        RECT 23.728 145.854 23.832 150.228 ; 
        RECT 23.296 145.854 23.4 150.228 ; 
        RECT 22.864 145.854 22.968 150.228 ; 
        RECT 22.432 145.854 22.536 150.228 ; 
        RECT 22 145.854 22.104 150.228 ; 
        RECT 21.568 145.854 21.672 150.228 ; 
        RECT 21.136 145.854 21.24 150.228 ; 
        RECT 20.704 145.854 20.808 150.228 ; 
        RECT 20.272 145.854 20.376 150.228 ; 
        RECT 19.84 145.854 19.944 150.228 ; 
        RECT 19.408 145.854 19.512 150.228 ; 
        RECT 18.976 145.854 19.08 150.228 ; 
        RECT 18.544 145.854 18.648 150.228 ; 
        RECT 18.112 145.854 18.216 150.228 ; 
        RECT 17.68 145.854 17.784 150.228 ; 
        RECT 17.248 145.854 17.352 150.228 ; 
        RECT 16.816 145.854 16.92 150.228 ; 
        RECT 16.384 145.854 16.488 150.228 ; 
        RECT 15.952 145.854 16.056 150.228 ; 
        RECT 15.52 145.854 15.624 150.228 ; 
        RECT 15.088 145.854 15.192 150.228 ; 
        RECT 14.656 145.854 14.76 150.228 ; 
        RECT 14.224 145.854 14.328 150.228 ; 
        RECT 13.792 145.854 13.896 150.228 ; 
        RECT 13.36 145.854 13.464 150.228 ; 
        RECT 12.928 145.854 13.032 150.228 ; 
        RECT 12.496 145.854 12.6 150.228 ; 
        RECT 12.064 145.854 12.168 150.228 ; 
        RECT 11.632 145.854 11.736 150.228 ; 
        RECT 11.2 145.854 11.304 150.228 ; 
        RECT 10.768 145.854 10.872 150.228 ; 
        RECT 10.336 145.854 10.44 150.228 ; 
        RECT 9.904 145.854 10.008 150.228 ; 
        RECT 9.472 145.854 9.576 150.228 ; 
        RECT 9.04 145.854 9.144 150.228 ; 
        RECT 8.608 145.854 8.712 150.228 ; 
        RECT 8.176 145.854 8.28 150.228 ; 
        RECT 7.744 145.854 7.848 150.228 ; 
        RECT 7.312 145.854 7.416 150.228 ; 
        RECT 6.88 145.854 6.984 150.228 ; 
        RECT 6.448 145.854 6.552 150.228 ; 
        RECT 6.016 145.854 6.12 150.228 ; 
        RECT 5.584 145.854 5.688 150.228 ; 
        RECT 5.152 145.854 5.256 150.228 ; 
        RECT 4.72 145.854 4.824 150.228 ; 
        RECT 4.288 145.854 4.392 150.228 ; 
        RECT 3.856 145.854 3.96 150.228 ; 
        RECT 3.424 145.854 3.528 150.228 ; 
        RECT 2.992 145.854 3.096 150.228 ; 
        RECT 2.56 145.854 2.664 150.228 ; 
        RECT 2.128 145.854 2.232 150.228 ; 
        RECT 1.696 145.854 1.8 150.228 ; 
        RECT 1.264 145.854 1.368 150.228 ; 
        RECT 0.832 145.854 0.936 150.228 ; 
        RECT 0.02 145.854 0.36 150.228 ; 
        RECT 34.564 150.174 35.076 154.548 ; 
        RECT 34.508 152.836 35.076 154.126 ; 
        RECT 33.916 151.744 34.164 154.548 ; 
        RECT 33.86 152.982 34.164 153.596 ; 
        RECT 33.916 150.174 34.02 154.548 ; 
        RECT 33.916 150.658 34.076 151.616 ; 
        RECT 33.916 150.174 34.164 150.53 ; 
        RECT 32.728 151.976 33.552 154.548 ; 
        RECT 33.448 150.174 33.552 154.548 ; 
        RECT 32.728 153.084 33.608 154.116 ; 
        RECT 32.728 150.174 33.12 154.548 ; 
        RECT 31.06 150.174 31.392 154.548 ; 
        RECT 31.06 150.528 31.448 154.27 ; 
        RECT 65.776 150.174 66.116 154.548 ; 
        RECT 65.2 150.174 65.304 154.548 ; 
        RECT 64.768 150.174 64.872 154.548 ; 
        RECT 64.336 150.174 64.44 154.548 ; 
        RECT 63.904 150.174 64.008 154.548 ; 
        RECT 63.472 150.174 63.576 154.548 ; 
        RECT 63.04 150.174 63.144 154.548 ; 
        RECT 62.608 150.174 62.712 154.548 ; 
        RECT 62.176 150.174 62.28 154.548 ; 
        RECT 61.744 150.174 61.848 154.548 ; 
        RECT 61.312 150.174 61.416 154.548 ; 
        RECT 60.88 150.174 60.984 154.548 ; 
        RECT 60.448 150.174 60.552 154.548 ; 
        RECT 60.016 150.174 60.12 154.548 ; 
        RECT 59.584 150.174 59.688 154.548 ; 
        RECT 59.152 150.174 59.256 154.548 ; 
        RECT 58.72 150.174 58.824 154.548 ; 
        RECT 58.288 150.174 58.392 154.548 ; 
        RECT 57.856 150.174 57.96 154.548 ; 
        RECT 57.424 150.174 57.528 154.548 ; 
        RECT 56.992 150.174 57.096 154.548 ; 
        RECT 56.56 150.174 56.664 154.548 ; 
        RECT 56.128 150.174 56.232 154.548 ; 
        RECT 55.696 150.174 55.8 154.548 ; 
        RECT 55.264 150.174 55.368 154.548 ; 
        RECT 54.832 150.174 54.936 154.548 ; 
        RECT 54.4 150.174 54.504 154.548 ; 
        RECT 53.968 150.174 54.072 154.548 ; 
        RECT 53.536 150.174 53.64 154.548 ; 
        RECT 53.104 150.174 53.208 154.548 ; 
        RECT 52.672 150.174 52.776 154.548 ; 
        RECT 52.24 150.174 52.344 154.548 ; 
        RECT 51.808 150.174 51.912 154.548 ; 
        RECT 51.376 150.174 51.48 154.548 ; 
        RECT 50.944 150.174 51.048 154.548 ; 
        RECT 50.512 150.174 50.616 154.548 ; 
        RECT 50.08 150.174 50.184 154.548 ; 
        RECT 49.648 150.174 49.752 154.548 ; 
        RECT 49.216 150.174 49.32 154.548 ; 
        RECT 48.784 150.174 48.888 154.548 ; 
        RECT 48.352 150.174 48.456 154.548 ; 
        RECT 47.92 150.174 48.024 154.548 ; 
        RECT 47.488 150.174 47.592 154.548 ; 
        RECT 47.056 150.174 47.16 154.548 ; 
        RECT 46.624 150.174 46.728 154.548 ; 
        RECT 46.192 150.174 46.296 154.548 ; 
        RECT 45.76 150.174 45.864 154.548 ; 
        RECT 45.328 150.174 45.432 154.548 ; 
        RECT 44.896 150.174 45 154.548 ; 
        RECT 44.464 150.174 44.568 154.548 ; 
        RECT 44.032 150.174 44.136 154.548 ; 
        RECT 43.6 150.174 43.704 154.548 ; 
        RECT 43.168 150.174 43.272 154.548 ; 
        RECT 42.736 150.174 42.84 154.548 ; 
        RECT 42.304 150.174 42.408 154.548 ; 
        RECT 41.872 150.174 41.976 154.548 ; 
        RECT 41.44 150.174 41.544 154.548 ; 
        RECT 41.008 150.174 41.112 154.548 ; 
        RECT 40.576 150.174 40.68 154.548 ; 
        RECT 40.144 150.174 40.248 154.548 ; 
        RECT 39.712 150.174 39.816 154.548 ; 
        RECT 39.28 150.174 39.384 154.548 ; 
        RECT 38.848 150.174 38.952 154.548 ; 
        RECT 38.416 150.174 38.52 154.548 ; 
        RECT 37.984 150.174 38.088 154.548 ; 
        RECT 37.552 150.174 37.656 154.548 ; 
        RECT 36.7 150.174 37.008 154.548 ; 
        RECT 29.128 150.174 29.436 154.548 ; 
        RECT 28.48 150.174 28.584 154.548 ; 
        RECT 28.048 150.174 28.152 154.548 ; 
        RECT 27.616 150.174 27.72 154.548 ; 
        RECT 27.184 150.174 27.288 154.548 ; 
        RECT 26.752 150.174 26.856 154.548 ; 
        RECT 26.32 150.174 26.424 154.548 ; 
        RECT 25.888 150.174 25.992 154.548 ; 
        RECT 25.456 150.174 25.56 154.548 ; 
        RECT 25.024 150.174 25.128 154.548 ; 
        RECT 24.592 150.174 24.696 154.548 ; 
        RECT 24.16 150.174 24.264 154.548 ; 
        RECT 23.728 150.174 23.832 154.548 ; 
        RECT 23.296 150.174 23.4 154.548 ; 
        RECT 22.864 150.174 22.968 154.548 ; 
        RECT 22.432 150.174 22.536 154.548 ; 
        RECT 22 150.174 22.104 154.548 ; 
        RECT 21.568 150.174 21.672 154.548 ; 
        RECT 21.136 150.174 21.24 154.548 ; 
        RECT 20.704 150.174 20.808 154.548 ; 
        RECT 20.272 150.174 20.376 154.548 ; 
        RECT 19.84 150.174 19.944 154.548 ; 
        RECT 19.408 150.174 19.512 154.548 ; 
        RECT 18.976 150.174 19.08 154.548 ; 
        RECT 18.544 150.174 18.648 154.548 ; 
        RECT 18.112 150.174 18.216 154.548 ; 
        RECT 17.68 150.174 17.784 154.548 ; 
        RECT 17.248 150.174 17.352 154.548 ; 
        RECT 16.816 150.174 16.92 154.548 ; 
        RECT 16.384 150.174 16.488 154.548 ; 
        RECT 15.952 150.174 16.056 154.548 ; 
        RECT 15.52 150.174 15.624 154.548 ; 
        RECT 15.088 150.174 15.192 154.548 ; 
        RECT 14.656 150.174 14.76 154.548 ; 
        RECT 14.224 150.174 14.328 154.548 ; 
        RECT 13.792 150.174 13.896 154.548 ; 
        RECT 13.36 150.174 13.464 154.548 ; 
        RECT 12.928 150.174 13.032 154.548 ; 
        RECT 12.496 150.174 12.6 154.548 ; 
        RECT 12.064 150.174 12.168 154.548 ; 
        RECT 11.632 150.174 11.736 154.548 ; 
        RECT 11.2 150.174 11.304 154.548 ; 
        RECT 10.768 150.174 10.872 154.548 ; 
        RECT 10.336 150.174 10.44 154.548 ; 
        RECT 9.904 150.174 10.008 154.548 ; 
        RECT 9.472 150.174 9.576 154.548 ; 
        RECT 9.04 150.174 9.144 154.548 ; 
        RECT 8.608 150.174 8.712 154.548 ; 
        RECT 8.176 150.174 8.28 154.548 ; 
        RECT 7.744 150.174 7.848 154.548 ; 
        RECT 7.312 150.174 7.416 154.548 ; 
        RECT 6.88 150.174 6.984 154.548 ; 
        RECT 6.448 150.174 6.552 154.548 ; 
        RECT 6.016 150.174 6.12 154.548 ; 
        RECT 5.584 150.174 5.688 154.548 ; 
        RECT 5.152 150.174 5.256 154.548 ; 
        RECT 4.72 150.174 4.824 154.548 ; 
        RECT 4.288 150.174 4.392 154.548 ; 
        RECT 3.856 150.174 3.96 154.548 ; 
        RECT 3.424 150.174 3.528 154.548 ; 
        RECT 2.992 150.174 3.096 154.548 ; 
        RECT 2.56 150.174 2.664 154.548 ; 
        RECT 2.128 150.174 2.232 154.548 ; 
        RECT 1.696 150.174 1.8 154.548 ; 
        RECT 1.264 150.174 1.368 154.548 ; 
        RECT 0.832 150.174 0.936 154.548 ; 
        RECT 0.02 150.174 0.36 154.548 ; 
        RECT 34.564 154.494 35.076 158.868 ; 
        RECT 34.508 157.156 35.076 158.446 ; 
        RECT 33.916 156.064 34.164 158.868 ; 
        RECT 33.86 157.302 34.164 157.916 ; 
        RECT 33.916 154.494 34.02 158.868 ; 
        RECT 33.916 154.978 34.076 155.936 ; 
        RECT 33.916 154.494 34.164 154.85 ; 
        RECT 32.728 156.296 33.552 158.868 ; 
        RECT 33.448 154.494 33.552 158.868 ; 
        RECT 32.728 157.404 33.608 158.436 ; 
        RECT 32.728 154.494 33.12 158.868 ; 
        RECT 31.06 154.494 31.392 158.868 ; 
        RECT 31.06 154.848 31.448 158.59 ; 
        RECT 65.776 154.494 66.116 158.868 ; 
        RECT 65.2 154.494 65.304 158.868 ; 
        RECT 64.768 154.494 64.872 158.868 ; 
        RECT 64.336 154.494 64.44 158.868 ; 
        RECT 63.904 154.494 64.008 158.868 ; 
        RECT 63.472 154.494 63.576 158.868 ; 
        RECT 63.04 154.494 63.144 158.868 ; 
        RECT 62.608 154.494 62.712 158.868 ; 
        RECT 62.176 154.494 62.28 158.868 ; 
        RECT 61.744 154.494 61.848 158.868 ; 
        RECT 61.312 154.494 61.416 158.868 ; 
        RECT 60.88 154.494 60.984 158.868 ; 
        RECT 60.448 154.494 60.552 158.868 ; 
        RECT 60.016 154.494 60.12 158.868 ; 
        RECT 59.584 154.494 59.688 158.868 ; 
        RECT 59.152 154.494 59.256 158.868 ; 
        RECT 58.72 154.494 58.824 158.868 ; 
        RECT 58.288 154.494 58.392 158.868 ; 
        RECT 57.856 154.494 57.96 158.868 ; 
        RECT 57.424 154.494 57.528 158.868 ; 
        RECT 56.992 154.494 57.096 158.868 ; 
        RECT 56.56 154.494 56.664 158.868 ; 
        RECT 56.128 154.494 56.232 158.868 ; 
        RECT 55.696 154.494 55.8 158.868 ; 
        RECT 55.264 154.494 55.368 158.868 ; 
        RECT 54.832 154.494 54.936 158.868 ; 
        RECT 54.4 154.494 54.504 158.868 ; 
        RECT 53.968 154.494 54.072 158.868 ; 
        RECT 53.536 154.494 53.64 158.868 ; 
        RECT 53.104 154.494 53.208 158.868 ; 
        RECT 52.672 154.494 52.776 158.868 ; 
        RECT 52.24 154.494 52.344 158.868 ; 
        RECT 51.808 154.494 51.912 158.868 ; 
        RECT 51.376 154.494 51.48 158.868 ; 
        RECT 50.944 154.494 51.048 158.868 ; 
        RECT 50.512 154.494 50.616 158.868 ; 
        RECT 50.08 154.494 50.184 158.868 ; 
        RECT 49.648 154.494 49.752 158.868 ; 
        RECT 49.216 154.494 49.32 158.868 ; 
        RECT 48.784 154.494 48.888 158.868 ; 
        RECT 48.352 154.494 48.456 158.868 ; 
        RECT 47.92 154.494 48.024 158.868 ; 
        RECT 47.488 154.494 47.592 158.868 ; 
        RECT 47.056 154.494 47.16 158.868 ; 
        RECT 46.624 154.494 46.728 158.868 ; 
        RECT 46.192 154.494 46.296 158.868 ; 
        RECT 45.76 154.494 45.864 158.868 ; 
        RECT 45.328 154.494 45.432 158.868 ; 
        RECT 44.896 154.494 45 158.868 ; 
        RECT 44.464 154.494 44.568 158.868 ; 
        RECT 44.032 154.494 44.136 158.868 ; 
        RECT 43.6 154.494 43.704 158.868 ; 
        RECT 43.168 154.494 43.272 158.868 ; 
        RECT 42.736 154.494 42.84 158.868 ; 
        RECT 42.304 154.494 42.408 158.868 ; 
        RECT 41.872 154.494 41.976 158.868 ; 
        RECT 41.44 154.494 41.544 158.868 ; 
        RECT 41.008 154.494 41.112 158.868 ; 
        RECT 40.576 154.494 40.68 158.868 ; 
        RECT 40.144 154.494 40.248 158.868 ; 
        RECT 39.712 154.494 39.816 158.868 ; 
        RECT 39.28 154.494 39.384 158.868 ; 
        RECT 38.848 154.494 38.952 158.868 ; 
        RECT 38.416 154.494 38.52 158.868 ; 
        RECT 37.984 154.494 38.088 158.868 ; 
        RECT 37.552 154.494 37.656 158.868 ; 
        RECT 36.7 154.494 37.008 158.868 ; 
        RECT 29.128 154.494 29.436 158.868 ; 
        RECT 28.48 154.494 28.584 158.868 ; 
        RECT 28.048 154.494 28.152 158.868 ; 
        RECT 27.616 154.494 27.72 158.868 ; 
        RECT 27.184 154.494 27.288 158.868 ; 
        RECT 26.752 154.494 26.856 158.868 ; 
        RECT 26.32 154.494 26.424 158.868 ; 
        RECT 25.888 154.494 25.992 158.868 ; 
        RECT 25.456 154.494 25.56 158.868 ; 
        RECT 25.024 154.494 25.128 158.868 ; 
        RECT 24.592 154.494 24.696 158.868 ; 
        RECT 24.16 154.494 24.264 158.868 ; 
        RECT 23.728 154.494 23.832 158.868 ; 
        RECT 23.296 154.494 23.4 158.868 ; 
        RECT 22.864 154.494 22.968 158.868 ; 
        RECT 22.432 154.494 22.536 158.868 ; 
        RECT 22 154.494 22.104 158.868 ; 
        RECT 21.568 154.494 21.672 158.868 ; 
        RECT 21.136 154.494 21.24 158.868 ; 
        RECT 20.704 154.494 20.808 158.868 ; 
        RECT 20.272 154.494 20.376 158.868 ; 
        RECT 19.84 154.494 19.944 158.868 ; 
        RECT 19.408 154.494 19.512 158.868 ; 
        RECT 18.976 154.494 19.08 158.868 ; 
        RECT 18.544 154.494 18.648 158.868 ; 
        RECT 18.112 154.494 18.216 158.868 ; 
        RECT 17.68 154.494 17.784 158.868 ; 
        RECT 17.248 154.494 17.352 158.868 ; 
        RECT 16.816 154.494 16.92 158.868 ; 
        RECT 16.384 154.494 16.488 158.868 ; 
        RECT 15.952 154.494 16.056 158.868 ; 
        RECT 15.52 154.494 15.624 158.868 ; 
        RECT 15.088 154.494 15.192 158.868 ; 
        RECT 14.656 154.494 14.76 158.868 ; 
        RECT 14.224 154.494 14.328 158.868 ; 
        RECT 13.792 154.494 13.896 158.868 ; 
        RECT 13.36 154.494 13.464 158.868 ; 
        RECT 12.928 154.494 13.032 158.868 ; 
        RECT 12.496 154.494 12.6 158.868 ; 
        RECT 12.064 154.494 12.168 158.868 ; 
        RECT 11.632 154.494 11.736 158.868 ; 
        RECT 11.2 154.494 11.304 158.868 ; 
        RECT 10.768 154.494 10.872 158.868 ; 
        RECT 10.336 154.494 10.44 158.868 ; 
        RECT 9.904 154.494 10.008 158.868 ; 
        RECT 9.472 154.494 9.576 158.868 ; 
        RECT 9.04 154.494 9.144 158.868 ; 
        RECT 8.608 154.494 8.712 158.868 ; 
        RECT 8.176 154.494 8.28 158.868 ; 
        RECT 7.744 154.494 7.848 158.868 ; 
        RECT 7.312 154.494 7.416 158.868 ; 
        RECT 6.88 154.494 6.984 158.868 ; 
        RECT 6.448 154.494 6.552 158.868 ; 
        RECT 6.016 154.494 6.12 158.868 ; 
        RECT 5.584 154.494 5.688 158.868 ; 
        RECT 5.152 154.494 5.256 158.868 ; 
        RECT 4.72 154.494 4.824 158.868 ; 
        RECT 4.288 154.494 4.392 158.868 ; 
        RECT 3.856 154.494 3.96 158.868 ; 
        RECT 3.424 154.494 3.528 158.868 ; 
        RECT 2.992 154.494 3.096 158.868 ; 
        RECT 2.56 154.494 2.664 158.868 ; 
        RECT 2.128 154.494 2.232 158.868 ; 
        RECT 1.696 154.494 1.8 158.868 ; 
        RECT 1.264 154.494 1.368 158.868 ; 
        RECT 0.832 154.494 0.936 158.868 ; 
        RECT 0.02 154.494 0.36 158.868 ; 
        RECT 34.564 158.814 35.076 163.188 ; 
        RECT 34.508 161.476 35.076 162.766 ; 
        RECT 33.916 160.384 34.164 163.188 ; 
        RECT 33.86 161.622 34.164 162.236 ; 
        RECT 33.916 158.814 34.02 163.188 ; 
        RECT 33.916 159.298 34.076 160.256 ; 
        RECT 33.916 158.814 34.164 159.17 ; 
        RECT 32.728 160.616 33.552 163.188 ; 
        RECT 33.448 158.814 33.552 163.188 ; 
        RECT 32.728 161.724 33.608 162.756 ; 
        RECT 32.728 158.814 33.12 163.188 ; 
        RECT 31.06 158.814 31.392 163.188 ; 
        RECT 31.06 159.168 31.448 162.91 ; 
        RECT 65.776 158.814 66.116 163.188 ; 
        RECT 65.2 158.814 65.304 163.188 ; 
        RECT 64.768 158.814 64.872 163.188 ; 
        RECT 64.336 158.814 64.44 163.188 ; 
        RECT 63.904 158.814 64.008 163.188 ; 
        RECT 63.472 158.814 63.576 163.188 ; 
        RECT 63.04 158.814 63.144 163.188 ; 
        RECT 62.608 158.814 62.712 163.188 ; 
        RECT 62.176 158.814 62.28 163.188 ; 
        RECT 61.744 158.814 61.848 163.188 ; 
        RECT 61.312 158.814 61.416 163.188 ; 
        RECT 60.88 158.814 60.984 163.188 ; 
        RECT 60.448 158.814 60.552 163.188 ; 
        RECT 60.016 158.814 60.12 163.188 ; 
        RECT 59.584 158.814 59.688 163.188 ; 
        RECT 59.152 158.814 59.256 163.188 ; 
        RECT 58.72 158.814 58.824 163.188 ; 
        RECT 58.288 158.814 58.392 163.188 ; 
        RECT 57.856 158.814 57.96 163.188 ; 
        RECT 57.424 158.814 57.528 163.188 ; 
        RECT 56.992 158.814 57.096 163.188 ; 
        RECT 56.56 158.814 56.664 163.188 ; 
        RECT 56.128 158.814 56.232 163.188 ; 
        RECT 55.696 158.814 55.8 163.188 ; 
        RECT 55.264 158.814 55.368 163.188 ; 
        RECT 54.832 158.814 54.936 163.188 ; 
        RECT 54.4 158.814 54.504 163.188 ; 
        RECT 53.968 158.814 54.072 163.188 ; 
        RECT 53.536 158.814 53.64 163.188 ; 
        RECT 53.104 158.814 53.208 163.188 ; 
        RECT 52.672 158.814 52.776 163.188 ; 
        RECT 52.24 158.814 52.344 163.188 ; 
        RECT 51.808 158.814 51.912 163.188 ; 
        RECT 51.376 158.814 51.48 163.188 ; 
        RECT 50.944 158.814 51.048 163.188 ; 
        RECT 50.512 158.814 50.616 163.188 ; 
        RECT 50.08 158.814 50.184 163.188 ; 
        RECT 49.648 158.814 49.752 163.188 ; 
        RECT 49.216 158.814 49.32 163.188 ; 
        RECT 48.784 158.814 48.888 163.188 ; 
        RECT 48.352 158.814 48.456 163.188 ; 
        RECT 47.92 158.814 48.024 163.188 ; 
        RECT 47.488 158.814 47.592 163.188 ; 
        RECT 47.056 158.814 47.16 163.188 ; 
        RECT 46.624 158.814 46.728 163.188 ; 
        RECT 46.192 158.814 46.296 163.188 ; 
        RECT 45.76 158.814 45.864 163.188 ; 
        RECT 45.328 158.814 45.432 163.188 ; 
        RECT 44.896 158.814 45 163.188 ; 
        RECT 44.464 158.814 44.568 163.188 ; 
        RECT 44.032 158.814 44.136 163.188 ; 
        RECT 43.6 158.814 43.704 163.188 ; 
        RECT 43.168 158.814 43.272 163.188 ; 
        RECT 42.736 158.814 42.84 163.188 ; 
        RECT 42.304 158.814 42.408 163.188 ; 
        RECT 41.872 158.814 41.976 163.188 ; 
        RECT 41.44 158.814 41.544 163.188 ; 
        RECT 41.008 158.814 41.112 163.188 ; 
        RECT 40.576 158.814 40.68 163.188 ; 
        RECT 40.144 158.814 40.248 163.188 ; 
        RECT 39.712 158.814 39.816 163.188 ; 
        RECT 39.28 158.814 39.384 163.188 ; 
        RECT 38.848 158.814 38.952 163.188 ; 
        RECT 38.416 158.814 38.52 163.188 ; 
        RECT 37.984 158.814 38.088 163.188 ; 
        RECT 37.552 158.814 37.656 163.188 ; 
        RECT 36.7 158.814 37.008 163.188 ; 
        RECT 29.128 158.814 29.436 163.188 ; 
        RECT 28.48 158.814 28.584 163.188 ; 
        RECT 28.048 158.814 28.152 163.188 ; 
        RECT 27.616 158.814 27.72 163.188 ; 
        RECT 27.184 158.814 27.288 163.188 ; 
        RECT 26.752 158.814 26.856 163.188 ; 
        RECT 26.32 158.814 26.424 163.188 ; 
        RECT 25.888 158.814 25.992 163.188 ; 
        RECT 25.456 158.814 25.56 163.188 ; 
        RECT 25.024 158.814 25.128 163.188 ; 
        RECT 24.592 158.814 24.696 163.188 ; 
        RECT 24.16 158.814 24.264 163.188 ; 
        RECT 23.728 158.814 23.832 163.188 ; 
        RECT 23.296 158.814 23.4 163.188 ; 
        RECT 22.864 158.814 22.968 163.188 ; 
        RECT 22.432 158.814 22.536 163.188 ; 
        RECT 22 158.814 22.104 163.188 ; 
        RECT 21.568 158.814 21.672 163.188 ; 
        RECT 21.136 158.814 21.24 163.188 ; 
        RECT 20.704 158.814 20.808 163.188 ; 
        RECT 20.272 158.814 20.376 163.188 ; 
        RECT 19.84 158.814 19.944 163.188 ; 
        RECT 19.408 158.814 19.512 163.188 ; 
        RECT 18.976 158.814 19.08 163.188 ; 
        RECT 18.544 158.814 18.648 163.188 ; 
        RECT 18.112 158.814 18.216 163.188 ; 
        RECT 17.68 158.814 17.784 163.188 ; 
        RECT 17.248 158.814 17.352 163.188 ; 
        RECT 16.816 158.814 16.92 163.188 ; 
        RECT 16.384 158.814 16.488 163.188 ; 
        RECT 15.952 158.814 16.056 163.188 ; 
        RECT 15.52 158.814 15.624 163.188 ; 
        RECT 15.088 158.814 15.192 163.188 ; 
        RECT 14.656 158.814 14.76 163.188 ; 
        RECT 14.224 158.814 14.328 163.188 ; 
        RECT 13.792 158.814 13.896 163.188 ; 
        RECT 13.36 158.814 13.464 163.188 ; 
        RECT 12.928 158.814 13.032 163.188 ; 
        RECT 12.496 158.814 12.6 163.188 ; 
        RECT 12.064 158.814 12.168 163.188 ; 
        RECT 11.632 158.814 11.736 163.188 ; 
        RECT 11.2 158.814 11.304 163.188 ; 
        RECT 10.768 158.814 10.872 163.188 ; 
        RECT 10.336 158.814 10.44 163.188 ; 
        RECT 9.904 158.814 10.008 163.188 ; 
        RECT 9.472 158.814 9.576 163.188 ; 
        RECT 9.04 158.814 9.144 163.188 ; 
        RECT 8.608 158.814 8.712 163.188 ; 
        RECT 8.176 158.814 8.28 163.188 ; 
        RECT 7.744 158.814 7.848 163.188 ; 
        RECT 7.312 158.814 7.416 163.188 ; 
        RECT 6.88 158.814 6.984 163.188 ; 
        RECT 6.448 158.814 6.552 163.188 ; 
        RECT 6.016 158.814 6.12 163.188 ; 
        RECT 5.584 158.814 5.688 163.188 ; 
        RECT 5.152 158.814 5.256 163.188 ; 
        RECT 4.72 158.814 4.824 163.188 ; 
        RECT 4.288 158.814 4.392 163.188 ; 
        RECT 3.856 158.814 3.96 163.188 ; 
        RECT 3.424 158.814 3.528 163.188 ; 
        RECT 2.992 158.814 3.096 163.188 ; 
        RECT 2.56 158.814 2.664 163.188 ; 
        RECT 2.128 158.814 2.232 163.188 ; 
        RECT 1.696 158.814 1.8 163.188 ; 
        RECT 1.264 158.814 1.368 163.188 ; 
        RECT 0.832 158.814 0.936 163.188 ; 
        RECT 0.02 158.814 0.36 163.188 ; 
        RECT 34.564 163.134 35.076 167.508 ; 
        RECT 34.508 165.796 35.076 167.086 ; 
        RECT 33.916 164.704 34.164 167.508 ; 
        RECT 33.86 165.942 34.164 166.556 ; 
        RECT 33.916 163.134 34.02 167.508 ; 
        RECT 33.916 163.618 34.076 164.576 ; 
        RECT 33.916 163.134 34.164 163.49 ; 
        RECT 32.728 164.936 33.552 167.508 ; 
        RECT 33.448 163.134 33.552 167.508 ; 
        RECT 32.728 166.044 33.608 167.076 ; 
        RECT 32.728 163.134 33.12 167.508 ; 
        RECT 31.06 163.134 31.392 167.508 ; 
        RECT 31.06 163.488 31.448 167.23 ; 
        RECT 65.776 163.134 66.116 167.508 ; 
        RECT 65.2 163.134 65.304 167.508 ; 
        RECT 64.768 163.134 64.872 167.508 ; 
        RECT 64.336 163.134 64.44 167.508 ; 
        RECT 63.904 163.134 64.008 167.508 ; 
        RECT 63.472 163.134 63.576 167.508 ; 
        RECT 63.04 163.134 63.144 167.508 ; 
        RECT 62.608 163.134 62.712 167.508 ; 
        RECT 62.176 163.134 62.28 167.508 ; 
        RECT 61.744 163.134 61.848 167.508 ; 
        RECT 61.312 163.134 61.416 167.508 ; 
        RECT 60.88 163.134 60.984 167.508 ; 
        RECT 60.448 163.134 60.552 167.508 ; 
        RECT 60.016 163.134 60.12 167.508 ; 
        RECT 59.584 163.134 59.688 167.508 ; 
        RECT 59.152 163.134 59.256 167.508 ; 
        RECT 58.72 163.134 58.824 167.508 ; 
        RECT 58.288 163.134 58.392 167.508 ; 
        RECT 57.856 163.134 57.96 167.508 ; 
        RECT 57.424 163.134 57.528 167.508 ; 
        RECT 56.992 163.134 57.096 167.508 ; 
        RECT 56.56 163.134 56.664 167.508 ; 
        RECT 56.128 163.134 56.232 167.508 ; 
        RECT 55.696 163.134 55.8 167.508 ; 
        RECT 55.264 163.134 55.368 167.508 ; 
        RECT 54.832 163.134 54.936 167.508 ; 
        RECT 54.4 163.134 54.504 167.508 ; 
        RECT 53.968 163.134 54.072 167.508 ; 
        RECT 53.536 163.134 53.64 167.508 ; 
        RECT 53.104 163.134 53.208 167.508 ; 
        RECT 52.672 163.134 52.776 167.508 ; 
        RECT 52.24 163.134 52.344 167.508 ; 
        RECT 51.808 163.134 51.912 167.508 ; 
        RECT 51.376 163.134 51.48 167.508 ; 
        RECT 50.944 163.134 51.048 167.508 ; 
        RECT 50.512 163.134 50.616 167.508 ; 
        RECT 50.08 163.134 50.184 167.508 ; 
        RECT 49.648 163.134 49.752 167.508 ; 
        RECT 49.216 163.134 49.32 167.508 ; 
        RECT 48.784 163.134 48.888 167.508 ; 
        RECT 48.352 163.134 48.456 167.508 ; 
        RECT 47.92 163.134 48.024 167.508 ; 
        RECT 47.488 163.134 47.592 167.508 ; 
        RECT 47.056 163.134 47.16 167.508 ; 
        RECT 46.624 163.134 46.728 167.508 ; 
        RECT 46.192 163.134 46.296 167.508 ; 
        RECT 45.76 163.134 45.864 167.508 ; 
        RECT 45.328 163.134 45.432 167.508 ; 
        RECT 44.896 163.134 45 167.508 ; 
        RECT 44.464 163.134 44.568 167.508 ; 
        RECT 44.032 163.134 44.136 167.508 ; 
        RECT 43.6 163.134 43.704 167.508 ; 
        RECT 43.168 163.134 43.272 167.508 ; 
        RECT 42.736 163.134 42.84 167.508 ; 
        RECT 42.304 163.134 42.408 167.508 ; 
        RECT 41.872 163.134 41.976 167.508 ; 
        RECT 41.44 163.134 41.544 167.508 ; 
        RECT 41.008 163.134 41.112 167.508 ; 
        RECT 40.576 163.134 40.68 167.508 ; 
        RECT 40.144 163.134 40.248 167.508 ; 
        RECT 39.712 163.134 39.816 167.508 ; 
        RECT 39.28 163.134 39.384 167.508 ; 
        RECT 38.848 163.134 38.952 167.508 ; 
        RECT 38.416 163.134 38.52 167.508 ; 
        RECT 37.984 163.134 38.088 167.508 ; 
        RECT 37.552 163.134 37.656 167.508 ; 
        RECT 36.7 163.134 37.008 167.508 ; 
        RECT 29.128 163.134 29.436 167.508 ; 
        RECT 28.48 163.134 28.584 167.508 ; 
        RECT 28.048 163.134 28.152 167.508 ; 
        RECT 27.616 163.134 27.72 167.508 ; 
        RECT 27.184 163.134 27.288 167.508 ; 
        RECT 26.752 163.134 26.856 167.508 ; 
        RECT 26.32 163.134 26.424 167.508 ; 
        RECT 25.888 163.134 25.992 167.508 ; 
        RECT 25.456 163.134 25.56 167.508 ; 
        RECT 25.024 163.134 25.128 167.508 ; 
        RECT 24.592 163.134 24.696 167.508 ; 
        RECT 24.16 163.134 24.264 167.508 ; 
        RECT 23.728 163.134 23.832 167.508 ; 
        RECT 23.296 163.134 23.4 167.508 ; 
        RECT 22.864 163.134 22.968 167.508 ; 
        RECT 22.432 163.134 22.536 167.508 ; 
        RECT 22 163.134 22.104 167.508 ; 
        RECT 21.568 163.134 21.672 167.508 ; 
        RECT 21.136 163.134 21.24 167.508 ; 
        RECT 20.704 163.134 20.808 167.508 ; 
        RECT 20.272 163.134 20.376 167.508 ; 
        RECT 19.84 163.134 19.944 167.508 ; 
        RECT 19.408 163.134 19.512 167.508 ; 
        RECT 18.976 163.134 19.08 167.508 ; 
        RECT 18.544 163.134 18.648 167.508 ; 
        RECT 18.112 163.134 18.216 167.508 ; 
        RECT 17.68 163.134 17.784 167.508 ; 
        RECT 17.248 163.134 17.352 167.508 ; 
        RECT 16.816 163.134 16.92 167.508 ; 
        RECT 16.384 163.134 16.488 167.508 ; 
        RECT 15.952 163.134 16.056 167.508 ; 
        RECT 15.52 163.134 15.624 167.508 ; 
        RECT 15.088 163.134 15.192 167.508 ; 
        RECT 14.656 163.134 14.76 167.508 ; 
        RECT 14.224 163.134 14.328 167.508 ; 
        RECT 13.792 163.134 13.896 167.508 ; 
        RECT 13.36 163.134 13.464 167.508 ; 
        RECT 12.928 163.134 13.032 167.508 ; 
        RECT 12.496 163.134 12.6 167.508 ; 
        RECT 12.064 163.134 12.168 167.508 ; 
        RECT 11.632 163.134 11.736 167.508 ; 
        RECT 11.2 163.134 11.304 167.508 ; 
        RECT 10.768 163.134 10.872 167.508 ; 
        RECT 10.336 163.134 10.44 167.508 ; 
        RECT 9.904 163.134 10.008 167.508 ; 
        RECT 9.472 163.134 9.576 167.508 ; 
        RECT 9.04 163.134 9.144 167.508 ; 
        RECT 8.608 163.134 8.712 167.508 ; 
        RECT 8.176 163.134 8.28 167.508 ; 
        RECT 7.744 163.134 7.848 167.508 ; 
        RECT 7.312 163.134 7.416 167.508 ; 
        RECT 6.88 163.134 6.984 167.508 ; 
        RECT 6.448 163.134 6.552 167.508 ; 
        RECT 6.016 163.134 6.12 167.508 ; 
        RECT 5.584 163.134 5.688 167.508 ; 
        RECT 5.152 163.134 5.256 167.508 ; 
        RECT 4.72 163.134 4.824 167.508 ; 
        RECT 4.288 163.134 4.392 167.508 ; 
        RECT 3.856 163.134 3.96 167.508 ; 
        RECT 3.424 163.134 3.528 167.508 ; 
        RECT 2.992 163.134 3.096 167.508 ; 
        RECT 2.56 163.134 2.664 167.508 ; 
        RECT 2.128 163.134 2.232 167.508 ; 
        RECT 1.696 163.134 1.8 167.508 ; 
        RECT 1.264 163.134 1.368 167.508 ; 
        RECT 0.832 163.134 0.936 167.508 ; 
        RECT 0.02 163.134 0.36 167.508 ; 
        RECT 34.564 167.454 35.076 171.828 ; 
        RECT 34.508 170.116 35.076 171.406 ; 
        RECT 33.916 169.024 34.164 171.828 ; 
        RECT 33.86 170.262 34.164 170.876 ; 
        RECT 33.916 167.454 34.02 171.828 ; 
        RECT 33.916 167.938 34.076 168.896 ; 
        RECT 33.916 167.454 34.164 167.81 ; 
        RECT 32.728 169.256 33.552 171.828 ; 
        RECT 33.448 167.454 33.552 171.828 ; 
        RECT 32.728 170.364 33.608 171.396 ; 
        RECT 32.728 167.454 33.12 171.828 ; 
        RECT 31.06 167.454 31.392 171.828 ; 
        RECT 31.06 167.808 31.448 171.55 ; 
        RECT 65.776 167.454 66.116 171.828 ; 
        RECT 65.2 167.454 65.304 171.828 ; 
        RECT 64.768 167.454 64.872 171.828 ; 
        RECT 64.336 167.454 64.44 171.828 ; 
        RECT 63.904 167.454 64.008 171.828 ; 
        RECT 63.472 167.454 63.576 171.828 ; 
        RECT 63.04 167.454 63.144 171.828 ; 
        RECT 62.608 167.454 62.712 171.828 ; 
        RECT 62.176 167.454 62.28 171.828 ; 
        RECT 61.744 167.454 61.848 171.828 ; 
        RECT 61.312 167.454 61.416 171.828 ; 
        RECT 60.88 167.454 60.984 171.828 ; 
        RECT 60.448 167.454 60.552 171.828 ; 
        RECT 60.016 167.454 60.12 171.828 ; 
        RECT 59.584 167.454 59.688 171.828 ; 
        RECT 59.152 167.454 59.256 171.828 ; 
        RECT 58.72 167.454 58.824 171.828 ; 
        RECT 58.288 167.454 58.392 171.828 ; 
        RECT 57.856 167.454 57.96 171.828 ; 
        RECT 57.424 167.454 57.528 171.828 ; 
        RECT 56.992 167.454 57.096 171.828 ; 
        RECT 56.56 167.454 56.664 171.828 ; 
        RECT 56.128 167.454 56.232 171.828 ; 
        RECT 55.696 167.454 55.8 171.828 ; 
        RECT 55.264 167.454 55.368 171.828 ; 
        RECT 54.832 167.454 54.936 171.828 ; 
        RECT 54.4 167.454 54.504 171.828 ; 
        RECT 53.968 167.454 54.072 171.828 ; 
        RECT 53.536 167.454 53.64 171.828 ; 
        RECT 53.104 167.454 53.208 171.828 ; 
        RECT 52.672 167.454 52.776 171.828 ; 
        RECT 52.24 167.454 52.344 171.828 ; 
        RECT 51.808 167.454 51.912 171.828 ; 
        RECT 51.376 167.454 51.48 171.828 ; 
        RECT 50.944 167.454 51.048 171.828 ; 
        RECT 50.512 167.454 50.616 171.828 ; 
        RECT 50.08 167.454 50.184 171.828 ; 
        RECT 49.648 167.454 49.752 171.828 ; 
        RECT 49.216 167.454 49.32 171.828 ; 
        RECT 48.784 167.454 48.888 171.828 ; 
        RECT 48.352 167.454 48.456 171.828 ; 
        RECT 47.92 167.454 48.024 171.828 ; 
        RECT 47.488 167.454 47.592 171.828 ; 
        RECT 47.056 167.454 47.16 171.828 ; 
        RECT 46.624 167.454 46.728 171.828 ; 
        RECT 46.192 167.454 46.296 171.828 ; 
        RECT 45.76 167.454 45.864 171.828 ; 
        RECT 45.328 167.454 45.432 171.828 ; 
        RECT 44.896 167.454 45 171.828 ; 
        RECT 44.464 167.454 44.568 171.828 ; 
        RECT 44.032 167.454 44.136 171.828 ; 
        RECT 43.6 167.454 43.704 171.828 ; 
        RECT 43.168 167.454 43.272 171.828 ; 
        RECT 42.736 167.454 42.84 171.828 ; 
        RECT 42.304 167.454 42.408 171.828 ; 
        RECT 41.872 167.454 41.976 171.828 ; 
        RECT 41.44 167.454 41.544 171.828 ; 
        RECT 41.008 167.454 41.112 171.828 ; 
        RECT 40.576 167.454 40.68 171.828 ; 
        RECT 40.144 167.454 40.248 171.828 ; 
        RECT 39.712 167.454 39.816 171.828 ; 
        RECT 39.28 167.454 39.384 171.828 ; 
        RECT 38.848 167.454 38.952 171.828 ; 
        RECT 38.416 167.454 38.52 171.828 ; 
        RECT 37.984 167.454 38.088 171.828 ; 
        RECT 37.552 167.454 37.656 171.828 ; 
        RECT 36.7 167.454 37.008 171.828 ; 
        RECT 29.128 167.454 29.436 171.828 ; 
        RECT 28.48 167.454 28.584 171.828 ; 
        RECT 28.048 167.454 28.152 171.828 ; 
        RECT 27.616 167.454 27.72 171.828 ; 
        RECT 27.184 167.454 27.288 171.828 ; 
        RECT 26.752 167.454 26.856 171.828 ; 
        RECT 26.32 167.454 26.424 171.828 ; 
        RECT 25.888 167.454 25.992 171.828 ; 
        RECT 25.456 167.454 25.56 171.828 ; 
        RECT 25.024 167.454 25.128 171.828 ; 
        RECT 24.592 167.454 24.696 171.828 ; 
        RECT 24.16 167.454 24.264 171.828 ; 
        RECT 23.728 167.454 23.832 171.828 ; 
        RECT 23.296 167.454 23.4 171.828 ; 
        RECT 22.864 167.454 22.968 171.828 ; 
        RECT 22.432 167.454 22.536 171.828 ; 
        RECT 22 167.454 22.104 171.828 ; 
        RECT 21.568 167.454 21.672 171.828 ; 
        RECT 21.136 167.454 21.24 171.828 ; 
        RECT 20.704 167.454 20.808 171.828 ; 
        RECT 20.272 167.454 20.376 171.828 ; 
        RECT 19.84 167.454 19.944 171.828 ; 
        RECT 19.408 167.454 19.512 171.828 ; 
        RECT 18.976 167.454 19.08 171.828 ; 
        RECT 18.544 167.454 18.648 171.828 ; 
        RECT 18.112 167.454 18.216 171.828 ; 
        RECT 17.68 167.454 17.784 171.828 ; 
        RECT 17.248 167.454 17.352 171.828 ; 
        RECT 16.816 167.454 16.92 171.828 ; 
        RECT 16.384 167.454 16.488 171.828 ; 
        RECT 15.952 167.454 16.056 171.828 ; 
        RECT 15.52 167.454 15.624 171.828 ; 
        RECT 15.088 167.454 15.192 171.828 ; 
        RECT 14.656 167.454 14.76 171.828 ; 
        RECT 14.224 167.454 14.328 171.828 ; 
        RECT 13.792 167.454 13.896 171.828 ; 
        RECT 13.36 167.454 13.464 171.828 ; 
        RECT 12.928 167.454 13.032 171.828 ; 
        RECT 12.496 167.454 12.6 171.828 ; 
        RECT 12.064 167.454 12.168 171.828 ; 
        RECT 11.632 167.454 11.736 171.828 ; 
        RECT 11.2 167.454 11.304 171.828 ; 
        RECT 10.768 167.454 10.872 171.828 ; 
        RECT 10.336 167.454 10.44 171.828 ; 
        RECT 9.904 167.454 10.008 171.828 ; 
        RECT 9.472 167.454 9.576 171.828 ; 
        RECT 9.04 167.454 9.144 171.828 ; 
        RECT 8.608 167.454 8.712 171.828 ; 
        RECT 8.176 167.454 8.28 171.828 ; 
        RECT 7.744 167.454 7.848 171.828 ; 
        RECT 7.312 167.454 7.416 171.828 ; 
        RECT 6.88 167.454 6.984 171.828 ; 
        RECT 6.448 167.454 6.552 171.828 ; 
        RECT 6.016 167.454 6.12 171.828 ; 
        RECT 5.584 167.454 5.688 171.828 ; 
        RECT 5.152 167.454 5.256 171.828 ; 
        RECT 4.72 167.454 4.824 171.828 ; 
        RECT 4.288 167.454 4.392 171.828 ; 
        RECT 3.856 167.454 3.96 171.828 ; 
        RECT 3.424 167.454 3.528 171.828 ; 
        RECT 2.992 167.454 3.096 171.828 ; 
        RECT 2.56 167.454 2.664 171.828 ; 
        RECT 2.128 167.454 2.232 171.828 ; 
        RECT 1.696 167.454 1.8 171.828 ; 
        RECT 1.264 167.454 1.368 171.828 ; 
        RECT 0.832 167.454 0.936 171.828 ; 
        RECT 0.02 167.454 0.36 171.828 ; 
        RECT 34.564 171.774 35.076 176.148 ; 
        RECT 34.508 174.436 35.076 175.726 ; 
        RECT 33.916 173.344 34.164 176.148 ; 
        RECT 33.86 174.582 34.164 175.196 ; 
        RECT 33.916 171.774 34.02 176.148 ; 
        RECT 33.916 172.258 34.076 173.216 ; 
        RECT 33.916 171.774 34.164 172.13 ; 
        RECT 32.728 173.576 33.552 176.148 ; 
        RECT 33.448 171.774 33.552 176.148 ; 
        RECT 32.728 174.684 33.608 175.716 ; 
        RECT 32.728 171.774 33.12 176.148 ; 
        RECT 31.06 171.774 31.392 176.148 ; 
        RECT 31.06 172.128 31.448 175.87 ; 
        RECT 65.776 171.774 66.116 176.148 ; 
        RECT 65.2 171.774 65.304 176.148 ; 
        RECT 64.768 171.774 64.872 176.148 ; 
        RECT 64.336 171.774 64.44 176.148 ; 
        RECT 63.904 171.774 64.008 176.148 ; 
        RECT 63.472 171.774 63.576 176.148 ; 
        RECT 63.04 171.774 63.144 176.148 ; 
        RECT 62.608 171.774 62.712 176.148 ; 
        RECT 62.176 171.774 62.28 176.148 ; 
        RECT 61.744 171.774 61.848 176.148 ; 
        RECT 61.312 171.774 61.416 176.148 ; 
        RECT 60.88 171.774 60.984 176.148 ; 
        RECT 60.448 171.774 60.552 176.148 ; 
        RECT 60.016 171.774 60.12 176.148 ; 
        RECT 59.584 171.774 59.688 176.148 ; 
        RECT 59.152 171.774 59.256 176.148 ; 
        RECT 58.72 171.774 58.824 176.148 ; 
        RECT 58.288 171.774 58.392 176.148 ; 
        RECT 57.856 171.774 57.96 176.148 ; 
        RECT 57.424 171.774 57.528 176.148 ; 
        RECT 56.992 171.774 57.096 176.148 ; 
        RECT 56.56 171.774 56.664 176.148 ; 
        RECT 56.128 171.774 56.232 176.148 ; 
        RECT 55.696 171.774 55.8 176.148 ; 
        RECT 55.264 171.774 55.368 176.148 ; 
        RECT 54.832 171.774 54.936 176.148 ; 
        RECT 54.4 171.774 54.504 176.148 ; 
        RECT 53.968 171.774 54.072 176.148 ; 
        RECT 53.536 171.774 53.64 176.148 ; 
        RECT 53.104 171.774 53.208 176.148 ; 
        RECT 52.672 171.774 52.776 176.148 ; 
        RECT 52.24 171.774 52.344 176.148 ; 
        RECT 51.808 171.774 51.912 176.148 ; 
        RECT 51.376 171.774 51.48 176.148 ; 
        RECT 50.944 171.774 51.048 176.148 ; 
        RECT 50.512 171.774 50.616 176.148 ; 
        RECT 50.08 171.774 50.184 176.148 ; 
        RECT 49.648 171.774 49.752 176.148 ; 
        RECT 49.216 171.774 49.32 176.148 ; 
        RECT 48.784 171.774 48.888 176.148 ; 
        RECT 48.352 171.774 48.456 176.148 ; 
        RECT 47.92 171.774 48.024 176.148 ; 
        RECT 47.488 171.774 47.592 176.148 ; 
        RECT 47.056 171.774 47.16 176.148 ; 
        RECT 46.624 171.774 46.728 176.148 ; 
        RECT 46.192 171.774 46.296 176.148 ; 
        RECT 45.76 171.774 45.864 176.148 ; 
        RECT 45.328 171.774 45.432 176.148 ; 
        RECT 44.896 171.774 45 176.148 ; 
        RECT 44.464 171.774 44.568 176.148 ; 
        RECT 44.032 171.774 44.136 176.148 ; 
        RECT 43.6 171.774 43.704 176.148 ; 
        RECT 43.168 171.774 43.272 176.148 ; 
        RECT 42.736 171.774 42.84 176.148 ; 
        RECT 42.304 171.774 42.408 176.148 ; 
        RECT 41.872 171.774 41.976 176.148 ; 
        RECT 41.44 171.774 41.544 176.148 ; 
        RECT 41.008 171.774 41.112 176.148 ; 
        RECT 40.576 171.774 40.68 176.148 ; 
        RECT 40.144 171.774 40.248 176.148 ; 
        RECT 39.712 171.774 39.816 176.148 ; 
        RECT 39.28 171.774 39.384 176.148 ; 
        RECT 38.848 171.774 38.952 176.148 ; 
        RECT 38.416 171.774 38.52 176.148 ; 
        RECT 37.984 171.774 38.088 176.148 ; 
        RECT 37.552 171.774 37.656 176.148 ; 
        RECT 36.7 171.774 37.008 176.148 ; 
        RECT 29.128 171.774 29.436 176.148 ; 
        RECT 28.48 171.774 28.584 176.148 ; 
        RECT 28.048 171.774 28.152 176.148 ; 
        RECT 27.616 171.774 27.72 176.148 ; 
        RECT 27.184 171.774 27.288 176.148 ; 
        RECT 26.752 171.774 26.856 176.148 ; 
        RECT 26.32 171.774 26.424 176.148 ; 
        RECT 25.888 171.774 25.992 176.148 ; 
        RECT 25.456 171.774 25.56 176.148 ; 
        RECT 25.024 171.774 25.128 176.148 ; 
        RECT 24.592 171.774 24.696 176.148 ; 
        RECT 24.16 171.774 24.264 176.148 ; 
        RECT 23.728 171.774 23.832 176.148 ; 
        RECT 23.296 171.774 23.4 176.148 ; 
        RECT 22.864 171.774 22.968 176.148 ; 
        RECT 22.432 171.774 22.536 176.148 ; 
        RECT 22 171.774 22.104 176.148 ; 
        RECT 21.568 171.774 21.672 176.148 ; 
        RECT 21.136 171.774 21.24 176.148 ; 
        RECT 20.704 171.774 20.808 176.148 ; 
        RECT 20.272 171.774 20.376 176.148 ; 
        RECT 19.84 171.774 19.944 176.148 ; 
        RECT 19.408 171.774 19.512 176.148 ; 
        RECT 18.976 171.774 19.08 176.148 ; 
        RECT 18.544 171.774 18.648 176.148 ; 
        RECT 18.112 171.774 18.216 176.148 ; 
        RECT 17.68 171.774 17.784 176.148 ; 
        RECT 17.248 171.774 17.352 176.148 ; 
        RECT 16.816 171.774 16.92 176.148 ; 
        RECT 16.384 171.774 16.488 176.148 ; 
        RECT 15.952 171.774 16.056 176.148 ; 
        RECT 15.52 171.774 15.624 176.148 ; 
        RECT 15.088 171.774 15.192 176.148 ; 
        RECT 14.656 171.774 14.76 176.148 ; 
        RECT 14.224 171.774 14.328 176.148 ; 
        RECT 13.792 171.774 13.896 176.148 ; 
        RECT 13.36 171.774 13.464 176.148 ; 
        RECT 12.928 171.774 13.032 176.148 ; 
        RECT 12.496 171.774 12.6 176.148 ; 
        RECT 12.064 171.774 12.168 176.148 ; 
        RECT 11.632 171.774 11.736 176.148 ; 
        RECT 11.2 171.774 11.304 176.148 ; 
        RECT 10.768 171.774 10.872 176.148 ; 
        RECT 10.336 171.774 10.44 176.148 ; 
        RECT 9.904 171.774 10.008 176.148 ; 
        RECT 9.472 171.774 9.576 176.148 ; 
        RECT 9.04 171.774 9.144 176.148 ; 
        RECT 8.608 171.774 8.712 176.148 ; 
        RECT 8.176 171.774 8.28 176.148 ; 
        RECT 7.744 171.774 7.848 176.148 ; 
        RECT 7.312 171.774 7.416 176.148 ; 
        RECT 6.88 171.774 6.984 176.148 ; 
        RECT 6.448 171.774 6.552 176.148 ; 
        RECT 6.016 171.774 6.12 176.148 ; 
        RECT 5.584 171.774 5.688 176.148 ; 
        RECT 5.152 171.774 5.256 176.148 ; 
        RECT 4.72 171.774 4.824 176.148 ; 
        RECT 4.288 171.774 4.392 176.148 ; 
        RECT 3.856 171.774 3.96 176.148 ; 
        RECT 3.424 171.774 3.528 176.148 ; 
        RECT 2.992 171.774 3.096 176.148 ; 
        RECT 2.56 171.774 2.664 176.148 ; 
        RECT 2.128 171.774 2.232 176.148 ; 
        RECT 1.696 171.774 1.8 176.148 ; 
        RECT 1.264 171.774 1.368 176.148 ; 
        RECT 0.832 171.774 0.936 176.148 ; 
        RECT 0.02 171.774 0.36 176.148 ; 
        RECT 34.564 176.094 35.076 180.468 ; 
        RECT 34.508 178.756 35.076 180.046 ; 
        RECT 33.916 177.664 34.164 180.468 ; 
        RECT 33.86 178.902 34.164 179.516 ; 
        RECT 33.916 176.094 34.02 180.468 ; 
        RECT 33.916 176.578 34.076 177.536 ; 
        RECT 33.916 176.094 34.164 176.45 ; 
        RECT 32.728 177.896 33.552 180.468 ; 
        RECT 33.448 176.094 33.552 180.468 ; 
        RECT 32.728 179.004 33.608 180.036 ; 
        RECT 32.728 176.094 33.12 180.468 ; 
        RECT 31.06 176.094 31.392 180.468 ; 
        RECT 31.06 176.448 31.448 180.19 ; 
        RECT 65.776 176.094 66.116 180.468 ; 
        RECT 65.2 176.094 65.304 180.468 ; 
        RECT 64.768 176.094 64.872 180.468 ; 
        RECT 64.336 176.094 64.44 180.468 ; 
        RECT 63.904 176.094 64.008 180.468 ; 
        RECT 63.472 176.094 63.576 180.468 ; 
        RECT 63.04 176.094 63.144 180.468 ; 
        RECT 62.608 176.094 62.712 180.468 ; 
        RECT 62.176 176.094 62.28 180.468 ; 
        RECT 61.744 176.094 61.848 180.468 ; 
        RECT 61.312 176.094 61.416 180.468 ; 
        RECT 60.88 176.094 60.984 180.468 ; 
        RECT 60.448 176.094 60.552 180.468 ; 
        RECT 60.016 176.094 60.12 180.468 ; 
        RECT 59.584 176.094 59.688 180.468 ; 
        RECT 59.152 176.094 59.256 180.468 ; 
        RECT 58.72 176.094 58.824 180.468 ; 
        RECT 58.288 176.094 58.392 180.468 ; 
        RECT 57.856 176.094 57.96 180.468 ; 
        RECT 57.424 176.094 57.528 180.468 ; 
        RECT 56.992 176.094 57.096 180.468 ; 
        RECT 56.56 176.094 56.664 180.468 ; 
        RECT 56.128 176.094 56.232 180.468 ; 
        RECT 55.696 176.094 55.8 180.468 ; 
        RECT 55.264 176.094 55.368 180.468 ; 
        RECT 54.832 176.094 54.936 180.468 ; 
        RECT 54.4 176.094 54.504 180.468 ; 
        RECT 53.968 176.094 54.072 180.468 ; 
        RECT 53.536 176.094 53.64 180.468 ; 
        RECT 53.104 176.094 53.208 180.468 ; 
        RECT 52.672 176.094 52.776 180.468 ; 
        RECT 52.24 176.094 52.344 180.468 ; 
        RECT 51.808 176.094 51.912 180.468 ; 
        RECT 51.376 176.094 51.48 180.468 ; 
        RECT 50.944 176.094 51.048 180.468 ; 
        RECT 50.512 176.094 50.616 180.468 ; 
        RECT 50.08 176.094 50.184 180.468 ; 
        RECT 49.648 176.094 49.752 180.468 ; 
        RECT 49.216 176.094 49.32 180.468 ; 
        RECT 48.784 176.094 48.888 180.468 ; 
        RECT 48.352 176.094 48.456 180.468 ; 
        RECT 47.92 176.094 48.024 180.468 ; 
        RECT 47.488 176.094 47.592 180.468 ; 
        RECT 47.056 176.094 47.16 180.468 ; 
        RECT 46.624 176.094 46.728 180.468 ; 
        RECT 46.192 176.094 46.296 180.468 ; 
        RECT 45.76 176.094 45.864 180.468 ; 
        RECT 45.328 176.094 45.432 180.468 ; 
        RECT 44.896 176.094 45 180.468 ; 
        RECT 44.464 176.094 44.568 180.468 ; 
        RECT 44.032 176.094 44.136 180.468 ; 
        RECT 43.6 176.094 43.704 180.468 ; 
        RECT 43.168 176.094 43.272 180.468 ; 
        RECT 42.736 176.094 42.84 180.468 ; 
        RECT 42.304 176.094 42.408 180.468 ; 
        RECT 41.872 176.094 41.976 180.468 ; 
        RECT 41.44 176.094 41.544 180.468 ; 
        RECT 41.008 176.094 41.112 180.468 ; 
        RECT 40.576 176.094 40.68 180.468 ; 
        RECT 40.144 176.094 40.248 180.468 ; 
        RECT 39.712 176.094 39.816 180.468 ; 
        RECT 39.28 176.094 39.384 180.468 ; 
        RECT 38.848 176.094 38.952 180.468 ; 
        RECT 38.416 176.094 38.52 180.468 ; 
        RECT 37.984 176.094 38.088 180.468 ; 
        RECT 37.552 176.094 37.656 180.468 ; 
        RECT 36.7 176.094 37.008 180.468 ; 
        RECT 29.128 176.094 29.436 180.468 ; 
        RECT 28.48 176.094 28.584 180.468 ; 
        RECT 28.048 176.094 28.152 180.468 ; 
        RECT 27.616 176.094 27.72 180.468 ; 
        RECT 27.184 176.094 27.288 180.468 ; 
        RECT 26.752 176.094 26.856 180.468 ; 
        RECT 26.32 176.094 26.424 180.468 ; 
        RECT 25.888 176.094 25.992 180.468 ; 
        RECT 25.456 176.094 25.56 180.468 ; 
        RECT 25.024 176.094 25.128 180.468 ; 
        RECT 24.592 176.094 24.696 180.468 ; 
        RECT 24.16 176.094 24.264 180.468 ; 
        RECT 23.728 176.094 23.832 180.468 ; 
        RECT 23.296 176.094 23.4 180.468 ; 
        RECT 22.864 176.094 22.968 180.468 ; 
        RECT 22.432 176.094 22.536 180.468 ; 
        RECT 22 176.094 22.104 180.468 ; 
        RECT 21.568 176.094 21.672 180.468 ; 
        RECT 21.136 176.094 21.24 180.468 ; 
        RECT 20.704 176.094 20.808 180.468 ; 
        RECT 20.272 176.094 20.376 180.468 ; 
        RECT 19.84 176.094 19.944 180.468 ; 
        RECT 19.408 176.094 19.512 180.468 ; 
        RECT 18.976 176.094 19.08 180.468 ; 
        RECT 18.544 176.094 18.648 180.468 ; 
        RECT 18.112 176.094 18.216 180.468 ; 
        RECT 17.68 176.094 17.784 180.468 ; 
        RECT 17.248 176.094 17.352 180.468 ; 
        RECT 16.816 176.094 16.92 180.468 ; 
        RECT 16.384 176.094 16.488 180.468 ; 
        RECT 15.952 176.094 16.056 180.468 ; 
        RECT 15.52 176.094 15.624 180.468 ; 
        RECT 15.088 176.094 15.192 180.468 ; 
        RECT 14.656 176.094 14.76 180.468 ; 
        RECT 14.224 176.094 14.328 180.468 ; 
        RECT 13.792 176.094 13.896 180.468 ; 
        RECT 13.36 176.094 13.464 180.468 ; 
        RECT 12.928 176.094 13.032 180.468 ; 
        RECT 12.496 176.094 12.6 180.468 ; 
        RECT 12.064 176.094 12.168 180.468 ; 
        RECT 11.632 176.094 11.736 180.468 ; 
        RECT 11.2 176.094 11.304 180.468 ; 
        RECT 10.768 176.094 10.872 180.468 ; 
        RECT 10.336 176.094 10.44 180.468 ; 
        RECT 9.904 176.094 10.008 180.468 ; 
        RECT 9.472 176.094 9.576 180.468 ; 
        RECT 9.04 176.094 9.144 180.468 ; 
        RECT 8.608 176.094 8.712 180.468 ; 
        RECT 8.176 176.094 8.28 180.468 ; 
        RECT 7.744 176.094 7.848 180.468 ; 
        RECT 7.312 176.094 7.416 180.468 ; 
        RECT 6.88 176.094 6.984 180.468 ; 
        RECT 6.448 176.094 6.552 180.468 ; 
        RECT 6.016 176.094 6.12 180.468 ; 
        RECT 5.584 176.094 5.688 180.468 ; 
        RECT 5.152 176.094 5.256 180.468 ; 
        RECT 4.72 176.094 4.824 180.468 ; 
        RECT 4.288 176.094 4.392 180.468 ; 
        RECT 3.856 176.094 3.96 180.468 ; 
        RECT 3.424 176.094 3.528 180.468 ; 
        RECT 2.992 176.094 3.096 180.468 ; 
        RECT 2.56 176.094 2.664 180.468 ; 
        RECT 2.128 176.094 2.232 180.468 ; 
        RECT 1.696 176.094 1.8 180.468 ; 
        RECT 1.264 176.094 1.368 180.468 ; 
        RECT 0.832 176.094 0.936 180.468 ; 
        RECT 0.02 176.094 0.36 180.468 ; 
  LAYER V3 SPACING 0.072 ; 
      RECT 0.02 4.88 66.116 5.4 ; 
      RECT 65.648 1.026 66.116 5.4 ; 
      RECT 37.208 4.496 65.576 5.4 ; 
      RECT 31.88 4.496 37.136 5.4 ; 
      RECT 29 1.026 31.52 5.4 ; 
      RECT 0.56 4.496 28.928 5.4 ; 
      RECT 0.02 1.026 0.488 5.4 ; 
      RECT 65.504 1.026 66.116 4.688 ; 
      RECT 37.424 1.026 65.432 5.4 ; 
      RECT 34.436 1.026 37.352 4.688 ; 
      RECT 33.788 1.808 34.292 5.4 ; 
      RECT 28.784 1.424 33.68 4.688 ; 
      RECT 0.704 1.026 28.712 5.4 ; 
      RECT 0.02 1.026 0.632 4.688 ; 
      RECT 34.22 1.026 66.116 4.304 ; 
      RECT 0.02 1.424 34.148 4.304 ; 
      RECT 33.32 1.026 66.116 1.712 ; 
      RECT 0.02 1.026 33.248 4.304 ; 
      RECT 0.02 1.026 66.116 1.328 ; 
      RECT 0.02 9.2 66.116 9.72 ; 
      RECT 65.648 5.346 66.116 9.72 ; 
      RECT 37.208 8.816 65.576 9.72 ; 
      RECT 31.88 8.816 37.136 9.72 ; 
      RECT 29 5.346 31.52 9.72 ; 
      RECT 0.56 8.816 28.928 9.72 ; 
      RECT 0.02 5.346 0.488 9.72 ; 
      RECT 65.504 5.346 66.116 9.008 ; 
      RECT 37.424 5.346 65.432 9.72 ; 
      RECT 34.436 5.346 37.352 9.008 ; 
      RECT 33.788 6.128 34.292 9.72 ; 
      RECT 28.784 5.744 33.68 9.008 ; 
      RECT 0.704 5.346 28.712 9.72 ; 
      RECT 0.02 5.346 0.632 9.008 ; 
      RECT 34.22 5.346 66.116 8.624 ; 
      RECT 0.02 5.744 34.148 8.624 ; 
      RECT 33.32 5.346 66.116 6.032 ; 
      RECT 0.02 5.346 33.248 8.624 ; 
      RECT 0.02 5.346 66.116 5.648 ; 
      RECT 0.02 13.52 66.116 14.04 ; 
      RECT 65.648 9.666 66.116 14.04 ; 
      RECT 37.208 13.136 65.576 14.04 ; 
      RECT 31.88 13.136 37.136 14.04 ; 
      RECT 29 9.666 31.52 14.04 ; 
      RECT 0.56 13.136 28.928 14.04 ; 
      RECT 0.02 9.666 0.488 14.04 ; 
      RECT 65.504 9.666 66.116 13.328 ; 
      RECT 37.424 9.666 65.432 14.04 ; 
      RECT 34.436 9.666 37.352 13.328 ; 
      RECT 33.788 10.448 34.292 14.04 ; 
      RECT 28.784 10.064 33.68 13.328 ; 
      RECT 0.704 9.666 28.712 14.04 ; 
      RECT 0.02 9.666 0.632 13.328 ; 
      RECT 34.22 9.666 66.116 12.944 ; 
      RECT 0.02 10.064 34.148 12.944 ; 
      RECT 33.32 9.666 66.116 10.352 ; 
      RECT 0.02 9.666 33.248 12.944 ; 
      RECT 0.02 9.666 66.116 9.968 ; 
      RECT 0.02 17.84 66.116 18.36 ; 
      RECT 65.648 13.986 66.116 18.36 ; 
      RECT 37.208 17.456 65.576 18.36 ; 
      RECT 31.88 17.456 37.136 18.36 ; 
      RECT 29 13.986 31.52 18.36 ; 
      RECT 0.56 17.456 28.928 18.36 ; 
      RECT 0.02 13.986 0.488 18.36 ; 
      RECT 65.504 13.986 66.116 17.648 ; 
      RECT 37.424 13.986 65.432 18.36 ; 
      RECT 34.436 13.986 37.352 17.648 ; 
      RECT 33.788 14.768 34.292 18.36 ; 
      RECT 28.784 14.384 33.68 17.648 ; 
      RECT 0.704 13.986 28.712 18.36 ; 
      RECT 0.02 13.986 0.632 17.648 ; 
      RECT 34.22 13.986 66.116 17.264 ; 
      RECT 0.02 14.384 34.148 17.264 ; 
      RECT 33.32 13.986 66.116 14.672 ; 
      RECT 0.02 13.986 33.248 17.264 ; 
      RECT 0.02 13.986 66.116 14.288 ; 
      RECT 0.02 22.16 66.116 22.68 ; 
      RECT 65.648 18.306 66.116 22.68 ; 
      RECT 37.208 21.776 65.576 22.68 ; 
      RECT 31.88 21.776 37.136 22.68 ; 
      RECT 29 18.306 31.52 22.68 ; 
      RECT 0.56 21.776 28.928 22.68 ; 
      RECT 0.02 18.306 0.488 22.68 ; 
      RECT 65.504 18.306 66.116 21.968 ; 
      RECT 37.424 18.306 65.432 22.68 ; 
      RECT 34.436 18.306 37.352 21.968 ; 
      RECT 33.788 19.088 34.292 22.68 ; 
      RECT 28.784 18.704 33.68 21.968 ; 
      RECT 0.704 18.306 28.712 22.68 ; 
      RECT 0.02 18.306 0.632 21.968 ; 
      RECT 34.22 18.306 66.116 21.584 ; 
      RECT 0.02 18.704 34.148 21.584 ; 
      RECT 33.32 18.306 66.116 18.992 ; 
      RECT 0.02 18.306 33.248 21.584 ; 
      RECT 0.02 18.306 66.116 18.608 ; 
      RECT 0.02 26.48 66.116 27 ; 
      RECT 65.648 22.626 66.116 27 ; 
      RECT 37.208 26.096 65.576 27 ; 
      RECT 31.88 26.096 37.136 27 ; 
      RECT 29 22.626 31.52 27 ; 
      RECT 0.56 26.096 28.928 27 ; 
      RECT 0.02 22.626 0.488 27 ; 
      RECT 65.504 22.626 66.116 26.288 ; 
      RECT 37.424 22.626 65.432 27 ; 
      RECT 34.436 22.626 37.352 26.288 ; 
      RECT 33.788 23.408 34.292 27 ; 
      RECT 28.784 23.024 33.68 26.288 ; 
      RECT 0.704 22.626 28.712 27 ; 
      RECT 0.02 22.626 0.632 26.288 ; 
      RECT 34.22 22.626 66.116 25.904 ; 
      RECT 0.02 23.024 34.148 25.904 ; 
      RECT 33.32 22.626 66.116 23.312 ; 
      RECT 0.02 22.626 33.248 25.904 ; 
      RECT 0.02 22.626 66.116 22.928 ; 
      RECT 0.02 30.8 66.116 31.32 ; 
      RECT 65.648 26.946 66.116 31.32 ; 
      RECT 37.208 30.416 65.576 31.32 ; 
      RECT 31.88 30.416 37.136 31.32 ; 
      RECT 29 26.946 31.52 31.32 ; 
      RECT 0.56 30.416 28.928 31.32 ; 
      RECT 0.02 26.946 0.488 31.32 ; 
      RECT 65.504 26.946 66.116 30.608 ; 
      RECT 37.424 26.946 65.432 31.32 ; 
      RECT 34.436 26.946 37.352 30.608 ; 
      RECT 33.788 27.728 34.292 31.32 ; 
      RECT 28.784 27.344 33.68 30.608 ; 
      RECT 0.704 26.946 28.712 31.32 ; 
      RECT 0.02 26.946 0.632 30.608 ; 
      RECT 34.22 26.946 66.116 30.224 ; 
      RECT 0.02 27.344 34.148 30.224 ; 
      RECT 33.32 26.946 66.116 27.632 ; 
      RECT 0.02 26.946 33.248 30.224 ; 
      RECT 0.02 26.946 66.116 27.248 ; 
      RECT 0.02 35.12 66.116 35.64 ; 
      RECT 65.648 31.266 66.116 35.64 ; 
      RECT 37.208 34.736 65.576 35.64 ; 
      RECT 31.88 34.736 37.136 35.64 ; 
      RECT 29 31.266 31.52 35.64 ; 
      RECT 0.56 34.736 28.928 35.64 ; 
      RECT 0.02 31.266 0.488 35.64 ; 
      RECT 65.504 31.266 66.116 34.928 ; 
      RECT 37.424 31.266 65.432 35.64 ; 
      RECT 34.436 31.266 37.352 34.928 ; 
      RECT 33.788 32.048 34.292 35.64 ; 
      RECT 28.784 31.664 33.68 34.928 ; 
      RECT 0.704 31.266 28.712 35.64 ; 
      RECT 0.02 31.266 0.632 34.928 ; 
      RECT 34.22 31.266 66.116 34.544 ; 
      RECT 0.02 31.664 34.148 34.544 ; 
      RECT 33.32 31.266 66.116 31.952 ; 
      RECT 0.02 31.266 33.248 34.544 ; 
      RECT 0.02 31.266 66.116 31.568 ; 
      RECT 0.02 39.44 66.116 39.96 ; 
      RECT 65.648 35.586 66.116 39.96 ; 
      RECT 37.208 39.056 65.576 39.96 ; 
      RECT 31.88 39.056 37.136 39.96 ; 
      RECT 29 35.586 31.52 39.96 ; 
      RECT 0.56 39.056 28.928 39.96 ; 
      RECT 0.02 35.586 0.488 39.96 ; 
      RECT 65.504 35.586 66.116 39.248 ; 
      RECT 37.424 35.586 65.432 39.96 ; 
      RECT 34.436 35.586 37.352 39.248 ; 
      RECT 33.788 36.368 34.292 39.96 ; 
      RECT 28.784 35.984 33.68 39.248 ; 
      RECT 0.704 35.586 28.712 39.96 ; 
      RECT 0.02 35.586 0.632 39.248 ; 
      RECT 34.22 35.586 66.116 38.864 ; 
      RECT 0.02 35.984 34.148 38.864 ; 
      RECT 33.32 35.586 66.116 36.272 ; 
      RECT 0.02 35.586 33.248 38.864 ; 
      RECT 0.02 35.586 66.116 35.888 ; 
      RECT 0.02 43.76 66.116 44.28 ; 
      RECT 65.648 39.906 66.116 44.28 ; 
      RECT 37.208 43.376 65.576 44.28 ; 
      RECT 31.88 43.376 37.136 44.28 ; 
      RECT 29 39.906 31.52 44.28 ; 
      RECT 0.56 43.376 28.928 44.28 ; 
      RECT 0.02 39.906 0.488 44.28 ; 
      RECT 65.504 39.906 66.116 43.568 ; 
      RECT 37.424 39.906 65.432 44.28 ; 
      RECT 34.436 39.906 37.352 43.568 ; 
      RECT 33.788 40.688 34.292 44.28 ; 
      RECT 28.784 40.304 33.68 43.568 ; 
      RECT 0.704 39.906 28.712 44.28 ; 
      RECT 0.02 39.906 0.632 43.568 ; 
      RECT 34.22 39.906 66.116 43.184 ; 
      RECT 0.02 40.304 34.148 43.184 ; 
      RECT 33.32 39.906 66.116 40.592 ; 
      RECT 0.02 39.906 33.248 43.184 ; 
      RECT 0.02 39.906 66.116 40.208 ; 
      RECT 0.02 48.08 66.116 48.6 ; 
      RECT 65.648 44.226 66.116 48.6 ; 
      RECT 37.208 47.696 65.576 48.6 ; 
      RECT 31.88 47.696 37.136 48.6 ; 
      RECT 29 44.226 31.52 48.6 ; 
      RECT 0.56 47.696 28.928 48.6 ; 
      RECT 0.02 44.226 0.488 48.6 ; 
      RECT 65.504 44.226 66.116 47.888 ; 
      RECT 37.424 44.226 65.432 48.6 ; 
      RECT 34.436 44.226 37.352 47.888 ; 
      RECT 33.788 45.008 34.292 48.6 ; 
      RECT 28.784 44.624 33.68 47.888 ; 
      RECT 0.704 44.226 28.712 48.6 ; 
      RECT 0.02 44.226 0.632 47.888 ; 
      RECT 34.22 44.226 66.116 47.504 ; 
      RECT 0.02 44.624 34.148 47.504 ; 
      RECT 33.32 44.226 66.116 44.912 ; 
      RECT 0.02 44.226 33.248 47.504 ; 
      RECT 0.02 44.226 66.116 44.528 ; 
      RECT 0.02 52.4 66.116 52.92 ; 
      RECT 65.648 48.546 66.116 52.92 ; 
      RECT 37.208 52.016 65.576 52.92 ; 
      RECT 31.88 52.016 37.136 52.92 ; 
      RECT 29 48.546 31.52 52.92 ; 
      RECT 0.56 52.016 28.928 52.92 ; 
      RECT 0.02 48.546 0.488 52.92 ; 
      RECT 65.504 48.546 66.116 52.208 ; 
      RECT 37.424 48.546 65.432 52.92 ; 
      RECT 34.436 48.546 37.352 52.208 ; 
      RECT 33.788 49.328 34.292 52.92 ; 
      RECT 28.784 48.944 33.68 52.208 ; 
      RECT 0.704 48.546 28.712 52.92 ; 
      RECT 0.02 48.546 0.632 52.208 ; 
      RECT 34.22 48.546 66.116 51.824 ; 
      RECT 0.02 48.944 34.148 51.824 ; 
      RECT 33.32 48.546 66.116 49.232 ; 
      RECT 0.02 48.546 33.248 51.824 ; 
      RECT 0.02 48.546 66.116 48.848 ; 
      RECT 0.02 56.72 66.116 57.24 ; 
      RECT 65.648 52.866 66.116 57.24 ; 
      RECT 37.208 56.336 65.576 57.24 ; 
      RECT 31.88 56.336 37.136 57.24 ; 
      RECT 29 52.866 31.52 57.24 ; 
      RECT 0.56 56.336 28.928 57.24 ; 
      RECT 0.02 52.866 0.488 57.24 ; 
      RECT 65.504 52.866 66.116 56.528 ; 
      RECT 37.424 52.866 65.432 57.24 ; 
      RECT 34.436 52.866 37.352 56.528 ; 
      RECT 33.788 53.648 34.292 57.24 ; 
      RECT 28.784 53.264 33.68 56.528 ; 
      RECT 0.704 52.866 28.712 57.24 ; 
      RECT 0.02 52.866 0.632 56.528 ; 
      RECT 34.22 52.866 66.116 56.144 ; 
      RECT 0.02 53.264 34.148 56.144 ; 
      RECT 33.32 52.866 66.116 53.552 ; 
      RECT 0.02 52.866 33.248 56.144 ; 
      RECT 0.02 52.866 66.116 53.168 ; 
      RECT 0.02 61.04 66.116 61.56 ; 
      RECT 65.648 57.186 66.116 61.56 ; 
      RECT 37.208 60.656 65.576 61.56 ; 
      RECT 31.88 60.656 37.136 61.56 ; 
      RECT 29 57.186 31.52 61.56 ; 
      RECT 0.56 60.656 28.928 61.56 ; 
      RECT 0.02 57.186 0.488 61.56 ; 
      RECT 65.504 57.186 66.116 60.848 ; 
      RECT 37.424 57.186 65.432 61.56 ; 
      RECT 34.436 57.186 37.352 60.848 ; 
      RECT 33.788 57.968 34.292 61.56 ; 
      RECT 28.784 57.584 33.68 60.848 ; 
      RECT 0.704 57.186 28.712 61.56 ; 
      RECT 0.02 57.186 0.632 60.848 ; 
      RECT 34.22 57.186 66.116 60.464 ; 
      RECT 0.02 57.584 34.148 60.464 ; 
      RECT 33.32 57.186 66.116 57.872 ; 
      RECT 0.02 57.186 33.248 60.464 ; 
      RECT 0.02 57.186 66.116 57.488 ; 
      RECT 0.02 65.36 66.116 65.88 ; 
      RECT 65.648 61.506 66.116 65.88 ; 
      RECT 37.208 64.976 65.576 65.88 ; 
      RECT 31.88 64.976 37.136 65.88 ; 
      RECT 29 61.506 31.52 65.88 ; 
      RECT 0.56 64.976 28.928 65.88 ; 
      RECT 0.02 61.506 0.488 65.88 ; 
      RECT 65.504 61.506 66.116 65.168 ; 
      RECT 37.424 61.506 65.432 65.88 ; 
      RECT 34.436 61.506 37.352 65.168 ; 
      RECT 33.788 62.288 34.292 65.88 ; 
      RECT 28.784 61.904 33.68 65.168 ; 
      RECT 0.704 61.506 28.712 65.88 ; 
      RECT 0.02 61.506 0.632 65.168 ; 
      RECT 34.22 61.506 66.116 64.784 ; 
      RECT 0.02 61.904 34.148 64.784 ; 
      RECT 33.32 61.506 66.116 62.192 ; 
      RECT 0.02 61.506 33.248 64.784 ; 
      RECT 0.02 61.506 66.116 61.808 ; 
      RECT 0.02 69.68 66.116 70.2 ; 
      RECT 65.648 65.826 66.116 70.2 ; 
      RECT 37.208 69.296 65.576 70.2 ; 
      RECT 31.88 69.296 37.136 70.2 ; 
      RECT 29 65.826 31.52 70.2 ; 
      RECT 0.56 69.296 28.928 70.2 ; 
      RECT 0.02 65.826 0.488 70.2 ; 
      RECT 65.504 65.826 66.116 69.488 ; 
      RECT 37.424 65.826 65.432 70.2 ; 
      RECT 34.436 65.826 37.352 69.488 ; 
      RECT 33.788 66.608 34.292 70.2 ; 
      RECT 28.784 66.224 33.68 69.488 ; 
      RECT 0.704 65.826 28.712 70.2 ; 
      RECT 0.02 65.826 0.632 69.488 ; 
      RECT 34.22 65.826 66.116 69.104 ; 
      RECT 0.02 66.224 34.148 69.104 ; 
      RECT 33.32 65.826 66.116 66.512 ; 
      RECT 0.02 65.826 33.248 69.104 ; 
      RECT 0.02 65.826 66.116 66.128 ; 
      RECT 0.02 74 66.116 74.52 ; 
      RECT 65.648 70.146 66.116 74.52 ; 
      RECT 37.208 73.616 65.576 74.52 ; 
      RECT 31.88 73.616 37.136 74.52 ; 
      RECT 29 70.146 31.52 74.52 ; 
      RECT 0.56 73.616 28.928 74.52 ; 
      RECT 0.02 70.146 0.488 74.52 ; 
      RECT 65.504 70.146 66.116 73.808 ; 
      RECT 37.424 70.146 65.432 74.52 ; 
      RECT 34.436 70.146 37.352 73.808 ; 
      RECT 33.788 70.928 34.292 74.52 ; 
      RECT 28.784 70.544 33.68 73.808 ; 
      RECT 0.704 70.146 28.712 74.52 ; 
      RECT 0.02 70.146 0.632 73.808 ; 
      RECT 34.22 70.146 66.116 73.424 ; 
      RECT 0.02 70.544 34.148 73.424 ; 
      RECT 33.32 70.146 66.116 70.832 ; 
      RECT 0.02 70.146 33.248 73.424 ; 
      RECT 0.02 70.146 66.116 70.448 ; 
      RECT 0 103.668 66.096 109.002 ; 
      RECT 43.236 74.388 66.096 109.002 ; 
      RECT 34.436 89.844 66.096 109.002 ; 
      RECT 38.052 79.476 66.096 109.002 ; 
      RECT 34.228 74.388 34.364 109.002 ; 
      RECT 34.02 74.388 34.156 109.002 ; 
      RECT 33.812 74.388 33.948 109.002 ; 
      RECT 33.604 74.388 33.74 109.002 ; 
      RECT 0 101.94 33.532 109.002 ; 
      RECT 32.564 90.996 66.096 102.804 ; 
      RECT 32.356 74.388 32.492 109.002 ; 
      RECT 32.148 74.388 32.284 109.002 ; 
      RECT 31.94 74.388 32.076 109.002 ; 
      RECT 31.732 74.388 31.868 109.002 ; 
      RECT 0 80.628 31.66 109.002 ; 
      RECT 0 89.268 33.532 101.076 ; 
      RECT 32.564 78.324 37.116 90.132 ; 
      RECT 37.26 80.244 66.096 109.002 ; 
      RECT 0 89.268 37.188 90.132 ; 
      RECT 32.564 80.244 66.096 89.748 ; 
      RECT 29.844 76.596 32.94 88.404 ; 
      RECT 28.98 77.172 31.66 109.002 ; 
      RECT 0 79.476 28.908 109.002 ; 
      RECT 27.252 74.388 29.052 80.532 ; 
      RECT 0 79.86 37.98 80.532 ; 
      RECT 37.188 79.476 66.096 80.148 ; 
      RECT 42.372 74.388 43.164 109.002 ; 
      RECT 27.252 78.708 42.3 79.764 ; 
      RECT 23.796 77.172 27.18 109.002 ; 
      RECT 0 74.388 23.724 109.002 ; 
      RECT 41.508 74.388 66.096 79.38 ; 
      RECT 40.644 77.172 66.096 79.38 ; 
      RECT 0 78.326 40.572 79.38 ; 
      RECT 39.78 74.388 41.436 78.612 ; 
      RECT 37.404 77.172 66.096 78.612 ; 
      RECT 34.436 77.172 37.332 79.764 ; 
      RECT 32.564 76.98 33.532 109.002 ; 
      RECT 33.012 74.388 34.524 77.46 ; 
      RECT 34.596 76.98 39.708 77.462 ; 
      RECT 26.388 76.98 29.772 79.38 ; 
      RECT 24.66 76.98 26.316 109.002 ; 
      RECT 0 74.388 24.588 79.38 ; 
      RECT 38.916 74.388 66.096 77.076 ; 
      RECT 33.012 74.708 38.844 77.076 ; 
      RECT 29.124 76.596 32.94 77.076 ; 
      RECT 25.524 74.388 29.052 77.076 ; 
      RECT 0 74.388 25.452 77.076 ; 
      RECT 37.188 74.388 66.096 76.884 ; 
      RECT 32.564 74.708 66.096 76.884 ; 
      RECT 0 74.388 31.66 76.884 ; 
      RECT 0 74.388 37.116 75.732 ; 
      RECT 0 74.388 66.096 74.612 ; 
        RECT 0.02 110.828 66.116 111.348 ; 
        RECT 65.648 106.974 66.116 111.348 ; 
        RECT 37.208 110.444 65.576 111.348 ; 
        RECT 31.88 110.444 37.136 111.348 ; 
        RECT 29 106.974 31.52 111.348 ; 
        RECT 0.56 110.444 28.928 111.348 ; 
        RECT 0.02 106.974 0.488 111.348 ; 
        RECT 65.504 106.974 66.116 110.636 ; 
        RECT 37.424 106.974 65.432 111.348 ; 
        RECT 34.436 106.974 37.352 110.636 ; 
        RECT 33.788 107.756 34.292 111.348 ; 
        RECT 28.784 107.372 33.68 110.636 ; 
        RECT 0.704 106.974 28.712 111.348 ; 
        RECT 0.02 106.974 0.632 110.636 ; 
        RECT 34.22 106.974 66.116 110.252 ; 
        RECT 0.02 107.372 34.148 110.252 ; 
        RECT 33.32 106.974 66.116 107.66 ; 
        RECT 0.02 106.974 33.248 110.252 ; 
        RECT 0.02 106.974 66.116 107.276 ; 
        RECT 0.02 115.148 66.116 115.668 ; 
        RECT 65.648 111.294 66.116 115.668 ; 
        RECT 37.208 114.764 65.576 115.668 ; 
        RECT 31.88 114.764 37.136 115.668 ; 
        RECT 29 111.294 31.52 115.668 ; 
        RECT 0.56 114.764 28.928 115.668 ; 
        RECT 0.02 111.294 0.488 115.668 ; 
        RECT 65.504 111.294 66.116 114.956 ; 
        RECT 37.424 111.294 65.432 115.668 ; 
        RECT 34.436 111.294 37.352 114.956 ; 
        RECT 33.788 112.076 34.292 115.668 ; 
        RECT 28.784 111.692 33.68 114.956 ; 
        RECT 0.704 111.294 28.712 115.668 ; 
        RECT 0.02 111.294 0.632 114.956 ; 
        RECT 34.22 111.294 66.116 114.572 ; 
        RECT 0.02 111.692 34.148 114.572 ; 
        RECT 33.32 111.294 66.116 111.98 ; 
        RECT 0.02 111.294 33.248 114.572 ; 
        RECT 0.02 111.294 66.116 111.596 ; 
        RECT 0.02 119.468 66.116 119.988 ; 
        RECT 65.648 115.614 66.116 119.988 ; 
        RECT 37.208 119.084 65.576 119.988 ; 
        RECT 31.88 119.084 37.136 119.988 ; 
        RECT 29 115.614 31.52 119.988 ; 
        RECT 0.56 119.084 28.928 119.988 ; 
        RECT 0.02 115.614 0.488 119.988 ; 
        RECT 65.504 115.614 66.116 119.276 ; 
        RECT 37.424 115.614 65.432 119.988 ; 
        RECT 34.436 115.614 37.352 119.276 ; 
        RECT 33.788 116.396 34.292 119.988 ; 
        RECT 28.784 116.012 33.68 119.276 ; 
        RECT 0.704 115.614 28.712 119.988 ; 
        RECT 0.02 115.614 0.632 119.276 ; 
        RECT 34.22 115.614 66.116 118.892 ; 
        RECT 0.02 116.012 34.148 118.892 ; 
        RECT 33.32 115.614 66.116 116.3 ; 
        RECT 0.02 115.614 33.248 118.892 ; 
        RECT 0.02 115.614 66.116 115.916 ; 
        RECT 0.02 123.788 66.116 124.308 ; 
        RECT 65.648 119.934 66.116 124.308 ; 
        RECT 37.208 123.404 65.576 124.308 ; 
        RECT 31.88 123.404 37.136 124.308 ; 
        RECT 29 119.934 31.52 124.308 ; 
        RECT 0.56 123.404 28.928 124.308 ; 
        RECT 0.02 119.934 0.488 124.308 ; 
        RECT 65.504 119.934 66.116 123.596 ; 
        RECT 37.424 119.934 65.432 124.308 ; 
        RECT 34.436 119.934 37.352 123.596 ; 
        RECT 33.788 120.716 34.292 124.308 ; 
        RECT 28.784 120.332 33.68 123.596 ; 
        RECT 0.704 119.934 28.712 124.308 ; 
        RECT 0.02 119.934 0.632 123.596 ; 
        RECT 34.22 119.934 66.116 123.212 ; 
        RECT 0.02 120.332 34.148 123.212 ; 
        RECT 33.32 119.934 66.116 120.62 ; 
        RECT 0.02 119.934 33.248 123.212 ; 
        RECT 0.02 119.934 66.116 120.236 ; 
        RECT 0.02 128.108 66.116 128.628 ; 
        RECT 65.648 124.254 66.116 128.628 ; 
        RECT 37.208 127.724 65.576 128.628 ; 
        RECT 31.88 127.724 37.136 128.628 ; 
        RECT 29 124.254 31.52 128.628 ; 
        RECT 0.56 127.724 28.928 128.628 ; 
        RECT 0.02 124.254 0.488 128.628 ; 
        RECT 65.504 124.254 66.116 127.916 ; 
        RECT 37.424 124.254 65.432 128.628 ; 
        RECT 34.436 124.254 37.352 127.916 ; 
        RECT 33.788 125.036 34.292 128.628 ; 
        RECT 28.784 124.652 33.68 127.916 ; 
        RECT 0.704 124.254 28.712 128.628 ; 
        RECT 0.02 124.254 0.632 127.916 ; 
        RECT 34.22 124.254 66.116 127.532 ; 
        RECT 0.02 124.652 34.148 127.532 ; 
        RECT 33.32 124.254 66.116 124.94 ; 
        RECT 0.02 124.254 33.248 127.532 ; 
        RECT 0.02 124.254 66.116 124.556 ; 
        RECT 0.02 132.428 66.116 132.948 ; 
        RECT 65.648 128.574 66.116 132.948 ; 
        RECT 37.208 132.044 65.576 132.948 ; 
        RECT 31.88 132.044 37.136 132.948 ; 
        RECT 29 128.574 31.52 132.948 ; 
        RECT 0.56 132.044 28.928 132.948 ; 
        RECT 0.02 128.574 0.488 132.948 ; 
        RECT 65.504 128.574 66.116 132.236 ; 
        RECT 37.424 128.574 65.432 132.948 ; 
        RECT 34.436 128.574 37.352 132.236 ; 
        RECT 33.788 129.356 34.292 132.948 ; 
        RECT 28.784 128.972 33.68 132.236 ; 
        RECT 0.704 128.574 28.712 132.948 ; 
        RECT 0.02 128.574 0.632 132.236 ; 
        RECT 34.22 128.574 66.116 131.852 ; 
        RECT 0.02 128.972 34.148 131.852 ; 
        RECT 33.32 128.574 66.116 129.26 ; 
        RECT 0.02 128.574 33.248 131.852 ; 
        RECT 0.02 128.574 66.116 128.876 ; 
        RECT 0.02 136.748 66.116 137.268 ; 
        RECT 65.648 132.894 66.116 137.268 ; 
        RECT 37.208 136.364 65.576 137.268 ; 
        RECT 31.88 136.364 37.136 137.268 ; 
        RECT 29 132.894 31.52 137.268 ; 
        RECT 0.56 136.364 28.928 137.268 ; 
        RECT 0.02 132.894 0.488 137.268 ; 
        RECT 65.504 132.894 66.116 136.556 ; 
        RECT 37.424 132.894 65.432 137.268 ; 
        RECT 34.436 132.894 37.352 136.556 ; 
        RECT 33.788 133.676 34.292 137.268 ; 
        RECT 28.784 133.292 33.68 136.556 ; 
        RECT 0.704 132.894 28.712 137.268 ; 
        RECT 0.02 132.894 0.632 136.556 ; 
        RECT 34.22 132.894 66.116 136.172 ; 
        RECT 0.02 133.292 34.148 136.172 ; 
        RECT 33.32 132.894 66.116 133.58 ; 
        RECT 0.02 132.894 33.248 136.172 ; 
        RECT 0.02 132.894 66.116 133.196 ; 
        RECT 0.02 141.068 66.116 141.588 ; 
        RECT 65.648 137.214 66.116 141.588 ; 
        RECT 37.208 140.684 65.576 141.588 ; 
        RECT 31.88 140.684 37.136 141.588 ; 
        RECT 29 137.214 31.52 141.588 ; 
        RECT 0.56 140.684 28.928 141.588 ; 
        RECT 0.02 137.214 0.488 141.588 ; 
        RECT 65.504 137.214 66.116 140.876 ; 
        RECT 37.424 137.214 65.432 141.588 ; 
        RECT 34.436 137.214 37.352 140.876 ; 
        RECT 33.788 137.996 34.292 141.588 ; 
        RECT 28.784 137.612 33.68 140.876 ; 
        RECT 0.704 137.214 28.712 141.588 ; 
        RECT 0.02 137.214 0.632 140.876 ; 
        RECT 34.22 137.214 66.116 140.492 ; 
        RECT 0.02 137.612 34.148 140.492 ; 
        RECT 33.32 137.214 66.116 137.9 ; 
        RECT 0.02 137.214 33.248 140.492 ; 
        RECT 0.02 137.214 66.116 137.516 ; 
        RECT 0.02 145.388 66.116 145.908 ; 
        RECT 65.648 141.534 66.116 145.908 ; 
        RECT 37.208 145.004 65.576 145.908 ; 
        RECT 31.88 145.004 37.136 145.908 ; 
        RECT 29 141.534 31.52 145.908 ; 
        RECT 0.56 145.004 28.928 145.908 ; 
        RECT 0.02 141.534 0.488 145.908 ; 
        RECT 65.504 141.534 66.116 145.196 ; 
        RECT 37.424 141.534 65.432 145.908 ; 
        RECT 34.436 141.534 37.352 145.196 ; 
        RECT 33.788 142.316 34.292 145.908 ; 
        RECT 28.784 141.932 33.68 145.196 ; 
        RECT 0.704 141.534 28.712 145.908 ; 
        RECT 0.02 141.534 0.632 145.196 ; 
        RECT 34.22 141.534 66.116 144.812 ; 
        RECT 0.02 141.932 34.148 144.812 ; 
        RECT 33.32 141.534 66.116 142.22 ; 
        RECT 0.02 141.534 33.248 144.812 ; 
        RECT 0.02 141.534 66.116 141.836 ; 
        RECT 0.02 149.708 66.116 150.228 ; 
        RECT 65.648 145.854 66.116 150.228 ; 
        RECT 37.208 149.324 65.576 150.228 ; 
        RECT 31.88 149.324 37.136 150.228 ; 
        RECT 29 145.854 31.52 150.228 ; 
        RECT 0.56 149.324 28.928 150.228 ; 
        RECT 0.02 145.854 0.488 150.228 ; 
        RECT 65.504 145.854 66.116 149.516 ; 
        RECT 37.424 145.854 65.432 150.228 ; 
        RECT 34.436 145.854 37.352 149.516 ; 
        RECT 33.788 146.636 34.292 150.228 ; 
        RECT 28.784 146.252 33.68 149.516 ; 
        RECT 0.704 145.854 28.712 150.228 ; 
        RECT 0.02 145.854 0.632 149.516 ; 
        RECT 34.22 145.854 66.116 149.132 ; 
        RECT 0.02 146.252 34.148 149.132 ; 
        RECT 33.32 145.854 66.116 146.54 ; 
        RECT 0.02 145.854 33.248 149.132 ; 
        RECT 0.02 145.854 66.116 146.156 ; 
        RECT 0.02 154.028 66.116 154.548 ; 
        RECT 65.648 150.174 66.116 154.548 ; 
        RECT 37.208 153.644 65.576 154.548 ; 
        RECT 31.88 153.644 37.136 154.548 ; 
        RECT 29 150.174 31.52 154.548 ; 
        RECT 0.56 153.644 28.928 154.548 ; 
        RECT 0.02 150.174 0.488 154.548 ; 
        RECT 65.504 150.174 66.116 153.836 ; 
        RECT 37.424 150.174 65.432 154.548 ; 
        RECT 34.436 150.174 37.352 153.836 ; 
        RECT 33.788 150.956 34.292 154.548 ; 
        RECT 28.784 150.572 33.68 153.836 ; 
        RECT 0.704 150.174 28.712 154.548 ; 
        RECT 0.02 150.174 0.632 153.836 ; 
        RECT 34.22 150.174 66.116 153.452 ; 
        RECT 0.02 150.572 34.148 153.452 ; 
        RECT 33.32 150.174 66.116 150.86 ; 
        RECT 0.02 150.174 33.248 153.452 ; 
        RECT 0.02 150.174 66.116 150.476 ; 
        RECT 0.02 158.348 66.116 158.868 ; 
        RECT 65.648 154.494 66.116 158.868 ; 
        RECT 37.208 157.964 65.576 158.868 ; 
        RECT 31.88 157.964 37.136 158.868 ; 
        RECT 29 154.494 31.52 158.868 ; 
        RECT 0.56 157.964 28.928 158.868 ; 
        RECT 0.02 154.494 0.488 158.868 ; 
        RECT 65.504 154.494 66.116 158.156 ; 
        RECT 37.424 154.494 65.432 158.868 ; 
        RECT 34.436 154.494 37.352 158.156 ; 
        RECT 33.788 155.276 34.292 158.868 ; 
        RECT 28.784 154.892 33.68 158.156 ; 
        RECT 0.704 154.494 28.712 158.868 ; 
        RECT 0.02 154.494 0.632 158.156 ; 
        RECT 34.22 154.494 66.116 157.772 ; 
        RECT 0.02 154.892 34.148 157.772 ; 
        RECT 33.32 154.494 66.116 155.18 ; 
        RECT 0.02 154.494 33.248 157.772 ; 
        RECT 0.02 154.494 66.116 154.796 ; 
        RECT 0.02 162.668 66.116 163.188 ; 
        RECT 65.648 158.814 66.116 163.188 ; 
        RECT 37.208 162.284 65.576 163.188 ; 
        RECT 31.88 162.284 37.136 163.188 ; 
        RECT 29 158.814 31.52 163.188 ; 
        RECT 0.56 162.284 28.928 163.188 ; 
        RECT 0.02 158.814 0.488 163.188 ; 
        RECT 65.504 158.814 66.116 162.476 ; 
        RECT 37.424 158.814 65.432 163.188 ; 
        RECT 34.436 158.814 37.352 162.476 ; 
        RECT 33.788 159.596 34.292 163.188 ; 
        RECT 28.784 159.212 33.68 162.476 ; 
        RECT 0.704 158.814 28.712 163.188 ; 
        RECT 0.02 158.814 0.632 162.476 ; 
        RECT 34.22 158.814 66.116 162.092 ; 
        RECT 0.02 159.212 34.148 162.092 ; 
        RECT 33.32 158.814 66.116 159.5 ; 
        RECT 0.02 158.814 33.248 162.092 ; 
        RECT 0.02 158.814 66.116 159.116 ; 
        RECT 0.02 166.988 66.116 167.508 ; 
        RECT 65.648 163.134 66.116 167.508 ; 
        RECT 37.208 166.604 65.576 167.508 ; 
        RECT 31.88 166.604 37.136 167.508 ; 
        RECT 29 163.134 31.52 167.508 ; 
        RECT 0.56 166.604 28.928 167.508 ; 
        RECT 0.02 163.134 0.488 167.508 ; 
        RECT 65.504 163.134 66.116 166.796 ; 
        RECT 37.424 163.134 65.432 167.508 ; 
        RECT 34.436 163.134 37.352 166.796 ; 
        RECT 33.788 163.916 34.292 167.508 ; 
        RECT 28.784 163.532 33.68 166.796 ; 
        RECT 0.704 163.134 28.712 167.508 ; 
        RECT 0.02 163.134 0.632 166.796 ; 
        RECT 34.22 163.134 66.116 166.412 ; 
        RECT 0.02 163.532 34.148 166.412 ; 
        RECT 33.32 163.134 66.116 163.82 ; 
        RECT 0.02 163.134 33.248 166.412 ; 
        RECT 0.02 163.134 66.116 163.436 ; 
        RECT 0.02 171.308 66.116 171.828 ; 
        RECT 65.648 167.454 66.116 171.828 ; 
        RECT 37.208 170.924 65.576 171.828 ; 
        RECT 31.88 170.924 37.136 171.828 ; 
        RECT 29 167.454 31.52 171.828 ; 
        RECT 0.56 170.924 28.928 171.828 ; 
        RECT 0.02 167.454 0.488 171.828 ; 
        RECT 65.504 167.454 66.116 171.116 ; 
        RECT 37.424 167.454 65.432 171.828 ; 
        RECT 34.436 167.454 37.352 171.116 ; 
        RECT 33.788 168.236 34.292 171.828 ; 
        RECT 28.784 167.852 33.68 171.116 ; 
        RECT 0.704 167.454 28.712 171.828 ; 
        RECT 0.02 167.454 0.632 171.116 ; 
        RECT 34.22 167.454 66.116 170.732 ; 
        RECT 0.02 167.852 34.148 170.732 ; 
        RECT 33.32 167.454 66.116 168.14 ; 
        RECT 0.02 167.454 33.248 170.732 ; 
        RECT 0.02 167.454 66.116 167.756 ; 
        RECT 0.02 175.628 66.116 176.148 ; 
        RECT 65.648 171.774 66.116 176.148 ; 
        RECT 37.208 175.244 65.576 176.148 ; 
        RECT 31.88 175.244 37.136 176.148 ; 
        RECT 29 171.774 31.52 176.148 ; 
        RECT 0.56 175.244 28.928 176.148 ; 
        RECT 0.02 171.774 0.488 176.148 ; 
        RECT 65.504 171.774 66.116 175.436 ; 
        RECT 37.424 171.774 65.432 176.148 ; 
        RECT 34.436 171.774 37.352 175.436 ; 
        RECT 33.788 172.556 34.292 176.148 ; 
        RECT 28.784 172.172 33.68 175.436 ; 
        RECT 0.704 171.774 28.712 176.148 ; 
        RECT 0.02 171.774 0.632 175.436 ; 
        RECT 34.22 171.774 66.116 175.052 ; 
        RECT 0.02 172.172 34.148 175.052 ; 
        RECT 33.32 171.774 66.116 172.46 ; 
        RECT 0.02 171.774 33.248 175.052 ; 
        RECT 0.02 171.774 66.116 172.076 ; 
        RECT 0.02 179.948 66.116 180.468 ; 
        RECT 65.648 176.094 66.116 180.468 ; 
        RECT 37.208 179.564 65.576 180.468 ; 
        RECT 31.88 179.564 37.136 180.468 ; 
        RECT 29 176.094 31.52 180.468 ; 
        RECT 0.56 179.564 28.928 180.468 ; 
        RECT 0.02 176.094 0.488 180.468 ; 
        RECT 65.504 176.094 66.116 179.756 ; 
        RECT 37.424 176.094 65.432 180.468 ; 
        RECT 34.436 176.094 37.352 179.756 ; 
        RECT 33.788 176.876 34.292 180.468 ; 
        RECT 28.784 176.492 33.68 179.756 ; 
        RECT 0.704 176.094 28.712 180.468 ; 
        RECT 0.02 176.094 0.632 179.756 ; 
        RECT 34.22 176.094 66.116 179.372 ; 
        RECT 0.02 176.492 34.148 179.372 ; 
        RECT 33.32 176.094 66.116 176.78 ; 
        RECT 0.02 176.094 33.248 179.372 ; 
        RECT 0.02 176.094 66.116 176.396 ; 
  LAYER M4 ; 
      RECT 6.276 81.24 60.038 81.336 ; 
      RECT 6.276 82.392 60.038 82.488 ; 
      RECT 6.276 83.928 60.038 84.024 ; 
      RECT 6.276 84.312 60.038 84.408 ; 
      RECT 6.276 85.656 60.038 85.752 ; 
      RECT 6.276 87.192 60.038 87.288 ; 
      RECT 43.82 77.076 44.156 77.172 ; 
      RECT 43.068 78.804 43.588 78.9 ; 
      RECT 43.1 81.434 43.568 81.53 ; 
      RECT 43.1 82.584 43.568 82.68 ; 
      RECT 40.544 78.804 42.828 78.9 ; 
      RECT 40.784 81.912 41.216 82.008 ; 
      RECT 35.452 83.412 39.824 83.508 ; 
      RECT 38.204 81.684 38.54 81.78 ; 
      RECT 35.068 86.484 38.54 86.58 ; 
      RECT 38.204 86.868 38.54 86.964 ; 
      RECT 37.492 79.764 37.828 79.86 ; 
      RECT 37.34 85.14 37.676 85.236 ; 
      RECT 37.34 88.02 37.676 88.116 ; 
      RECT 36.628 79.38 36.964 79.476 ; 
      RECT 35.772 74.228 36.824 74.324 ; 
      RECT 35.772 108.724 36.824 108.82 ; 
      RECT 35.836 85.332 36.812 85.428 ; 
      RECT 36.476 85.908 36.812 86.004 ; 
      RECT 30.652 86.868 36.812 86.964 ; 
      RECT 36.476 88.02 36.812 88.116 ; 
      RECT 35.54 108.34 36.592 108.436 ; 
      RECT 35.536 73.844 36.588 73.94 ; 
      RECT 35.384 73.46 36.436 73.556 ; 
      RECT 35.384 107.572 36.436 107.668 ; 
      RECT 36.044 89.748 36.38 89.844 ; 
      RECT 32.956 91.284 36.38 91.38 ; 
      RECT 34.492 100.308 36.38 100.404 ; 
      RECT 36.044 100.692 36.38 100.788 ; 
      RECT 35.192 73.076 36.244 73.172 ; 
      RECT 35.192 107.188 36.244 107.284 ; 
      RECT 34.3 96.66 36.08 96.756 ; 
      RECT 35.016 72.692 36.068 72.788 ; 
      RECT 35.016 108.532 36.068 108.628 ; 
      RECT 34.82 74.036 35.872 74.132 ; 
      RECT 34.82 108.148 35.872 108.244 ; 
      RECT 35.344 85.908 35.828 86.004 ; 
      RECT 35.26 94.356 35.792 94.452 ; 
      RECT 34.632 73.652 35.684 73.748 ; 
      RECT 34.632 107.764 35.684 107.86 ; 
      RECT 34.492 72.5 35.544 72.596 ; 
      RECT 34.492 107.38 35.544 107.476 ; 
      RECT 31.228 100.692 35.504 100.788 ; 
      RECT 35.168 105.3 35.504 105.396 ; 
      RECT 34.268 71.924 35.32 72.02 ; 
      RECT 34.268 106.996 35.32 107.092 ; 
      RECT 34.876 89.748 35.216 89.844 ; 
      RECT 30.46 92.052 34.928 92.148 ; 
      RECT 33.04 83.412 34.868 83.508 ; 
      RECT 32.348 74.804 33.416 74.9 ; 
      RECT 32.348 106.42 33.416 106.516 ; 
      RECT 32.896 89.556 33.332 89.652 ; 
      RECT 32.256 74.42 33.224 74.516 ; 
      RECT 32.256 108.916 33.224 109.012 ; 
      RECT 32.032 72.5 33 72.596 ; 
      RECT 32.148 109.3 33 109.396 ; 
      RECT 32.612 88.02 32.948 88.116 ; 
      RECT 31.816 72.884 32.808 72.98 ; 
      RECT 31.816 108.724 32.808 108.82 ; 
      RECT 30.88 98.388 32.564 98.484 ; 
      RECT 30.752 74.228 31.82 74.324 ; 
      RECT 30.752 109.3 31.82 109.396 ; 
      RECT 31.312 92.628 31.796 92.724 ; 
      RECT 31.28 105.3 31.616 105.396 ; 
      RECT 30.616 73.844 31.604 73.94 ; 
      RECT 30.348 107.572 31.604 107.668 ; 
      RECT 30.512 73.46 31.432 73.556 ; 
      RECT 30.464 108.916 31.432 109.012 ; 
      RECT 30.3 73.076 31.22 73.172 ; 
      RECT 30.884 98.964 31.22 99.06 ; 
      RECT 30.1 107.188 31.22 107.284 ; 
      RECT 30.12 72.692 31.04 72.788 ; 
      RECT 30.12 108.532 31.04 108.628 ; 
      RECT 26.272 88.02 31.028 88.116 ; 
      RECT 29.968 73.652 30.888 73.748 ; 
      RECT 29.968 108.148 30.888 108.244 ; 
      RECT 29.896 73.268 30.668 73.364 ; 
      RECT 29.896 107.764 30.668 107.86 ; 
      RECT 29.7 72.884 30.472 72.98 ; 
      RECT 29.7 107.38 30.472 107.476 ; 
      RECT 29.716 91.668 30.452 91.764 ; 
      RECT 29.492 72.5 30.264 72.596 ; 
      RECT 29.492 106.996 30.264 107.092 ; 
      RECT 27.556 80.916 30.26 81.012 ; 
      RECT 29.716 92.052 30.052 92.148 ; 
      RECT 28.64 74.612 29.692 74.708 ; 
      RECT 28.77 89.748 29.304 89.844 ; 
      RECT 27.404 81.684 27.74 81.78 ; 
  LAYER V4 ; 
      RECT 44.016 77.076 44.112 77.172 ; 
      RECT 44.016 81.24 44.112 81.336 ; 
      RECT 43.344 78.804 43.44 78.9 ; 
      RECT 43.344 81.434 43.44 81.53 ; 
      RECT 43.344 82.584 43.44 82.68 ; 
      RECT 40.848 78.804 40.944 78.9 ; 
      RECT 40.848 81.912 40.944 82.008 ; 
      RECT 38.4 81.684 38.496 81.78 ; 
      RECT 38.4 82.392 38.496 82.488 ; 
      RECT 38.4 86.484 38.496 86.58 ; 
      RECT 38.4 86.868 38.496 86.964 ; 
      RECT 37.536 79.764 37.632 79.86 ; 
      RECT 37.536 83.928 37.632 84.024 ; 
      RECT 37.536 85.14 37.632 85.236 ; 
      RECT 37.536 85.656 37.632 85.752 ; 
      RECT 37.536 87.192 37.632 87.288 ; 
      RECT 37.536 88.02 37.632 88.116 ; 
      RECT 36.672 79.38 36.768 79.476 ; 
      RECT 36.672 84.312 36.768 84.408 ; 
      RECT 36.672 85.332 36.768 85.428 ; 
      RECT 36.672 85.908 36.768 86.004 ; 
      RECT 36.672 86.868 36.768 86.964 ; 
      RECT 36.672 88.02 36.768 88.116 ; 
      RECT 36.24 89.748 36.336 89.844 ; 
      RECT 36.24 91.284 36.336 91.38 ; 
      RECT 36.24 100.308 36.336 100.404 ; 
      RECT 36.24 100.692 36.336 100.788 ; 
      RECT 35.88 74.228 35.976 74.324 ; 
      RECT 35.88 85.332 35.976 85.428 ; 
      RECT 35.88 108.724 35.976 108.82 ; 
      RECT 35.688 73.844 35.784 73.94 ; 
      RECT 35.688 85.908 35.784 86.004 ; 
      RECT 35.688 108.34 35.784 108.436 ; 
      RECT 35.496 73.46 35.592 73.556 ; 
      RECT 35.496 83.412 35.592 83.508 ; 
      RECT 35.496 107.572 35.592 107.668 ; 
      RECT 35.304 73.076 35.4 73.172 ; 
      RECT 35.304 94.356 35.4 94.452 ; 
      RECT 35.304 105.3 35.4 105.396 ; 
      RECT 35.304 107.188 35.4 107.284 ; 
      RECT 35.112 72.692 35.208 72.788 ; 
      RECT 35.112 86.484 35.208 86.58 ; 
      RECT 35.112 108.532 35.208 108.628 ; 
      RECT 34.92 74.036 35.016 74.132 ; 
      RECT 34.92 89.748 35.016 89.844 ; 
      RECT 34.92 108.148 35.016 108.244 ; 
      RECT 34.728 73.652 34.824 73.748 ; 
      RECT 34.728 83.412 34.824 83.508 ; 
      RECT 34.728 107.764 34.824 107.86 ; 
      RECT 34.536 72.5 34.632 72.596 ; 
      RECT 34.536 100.308 34.632 100.404 ; 
      RECT 34.536 107.38 34.632 107.476 ; 
      RECT 34.344 71.924 34.44 72.02 ; 
      RECT 34.344 96.66 34.44 96.756 ; 
      RECT 34.344 106.996 34.44 107.092 ; 
      RECT 33.192 74.804 33.288 74.9 ; 
      RECT 33.192 89.556 33.288 89.652 ; 
      RECT 33.192 106.42 33.288 106.516 ; 
      RECT 33 74.42 33.096 74.516 ; 
      RECT 33 91.284 33.096 91.38 ; 
      RECT 33 108.916 33.096 109.012 ; 
      RECT 32.808 72.5 32.904 72.596 ; 
      RECT 32.808 88.02 32.904 88.116 ; 
      RECT 32.808 109.3 32.904 109.396 ; 
      RECT 32.424 72.884 32.52 72.98 ; 
      RECT 32.424 98.388 32.52 98.484 ; 
      RECT 32.424 108.724 32.52 108.82 ; 
      RECT 31.656 74.228 31.752 74.324 ; 
      RECT 31.656 92.628 31.752 92.724 ; 
      RECT 31.656 109.3 31.752 109.396 ; 
      RECT 31.464 73.844 31.56 73.94 ; 
      RECT 31.464 105.3 31.56 105.396 ; 
      RECT 31.464 107.572 31.56 107.668 ; 
      RECT 31.272 73.46 31.368 73.556 ; 
      RECT 31.272 100.692 31.368 100.788 ; 
      RECT 31.272 108.916 31.368 109.012 ; 
      RECT 31.08 73.076 31.176 73.172 ; 
      RECT 31.08 98.964 31.176 99.06 ; 
      RECT 31.08 107.188 31.176 107.284 ; 
      RECT 30.888 72.692 30.984 72.788 ; 
      RECT 30.888 88.02 30.984 88.116 ; 
      RECT 30.888 108.532 30.984 108.628 ; 
      RECT 30.696 73.652 30.792 73.748 ; 
      RECT 30.696 86.868 30.792 86.964 ; 
      RECT 30.696 108.148 30.792 108.244 ; 
      RECT 30.504 73.268 30.6 73.364 ; 
      RECT 30.504 92.052 30.6 92.148 ; 
      RECT 30.504 107.764 30.6 107.86 ; 
      RECT 30.312 72.884 30.408 72.98 ; 
      RECT 30.312 91.668 30.408 91.764 ; 
      RECT 30.312 107.38 30.408 107.476 ; 
      RECT 30.12 72.5 30.216 72.596 ; 
      RECT 30.12 80.916 30.216 81.012 ; 
      RECT 30.12 106.996 30.216 107.092 ; 
      RECT 29.76 91.668 29.856 91.764 ; 
      RECT 29.76 92.052 29.856 92.148 ; 
      RECT 29.088 74.612 29.184 74.708 ; 
      RECT 29.088 89.748 29.184 89.844 ; 
      RECT 27.6 80.916 27.696 81.012 ; 
      RECT 27.6 81.684 27.696 81.78 ; 
  LAYER M5 ; 
      RECT 44.016 77.032 44.112 81.38 ; 
      RECT 43.344 78.692 43.44 82.934 ; 
      RECT 40.848 78.726 40.944 82.056 ; 
      RECT 38.4 81.64 38.496 82.532 ; 
      RECT 38.4 86.44 38.496 87.008 ; 
      RECT 37.536 79.72 37.632 84.068 ; 
      RECT 37.536 85.096 37.632 85.796 ; 
      RECT 37.536 87.148 37.632 88.16 ; 
      RECT 36.672 79.336 36.768 84.452 ; 
      RECT 36.672 85.288 36.768 86.048 ; 
      RECT 36.672 86.824 36.768 88.16 ; 
      RECT 36.24 89.704 36.336 91.424 ; 
      RECT 36.24 100.264 36.336 100.832 ; 
      RECT 35.88 75.576 35.976 105.908 ; 
      RECT 35.688 75.576 35.784 105.908 ; 
      RECT 35.496 75.576 35.592 105.908 ; 
      RECT 35.304 75.576 35.4 105.908 ; 
      RECT 35.112 75.576 35.208 105.908 ; 
      RECT 34.92 75.576 35.016 105.908 ; 
      RECT 34.728 75.576 34.824 105.908 ; 
      RECT 34.536 75.576 34.632 105.908 ; 
      RECT 34.344 75.576 34.44 105.908 ; 
      RECT 33.192 75.576 33.288 105.908 ; 
      RECT 33 75.576 33.096 105.908 ; 
      RECT 32.808 75.576 32.904 105.908 ; 
      RECT 32.424 75.576 32.52 105.908 ; 
      RECT 31.656 75.576 31.752 105.908 ; 
      RECT 31.464 75.576 31.56 105.908 ; 
      RECT 31.272 75.576 31.368 105.908 ; 
      RECT 31.08 75.576 31.176 105.908 ; 
      RECT 30.888 75.576 30.984 105.908 ; 
      RECT 30.696 75.576 30.792 105.908 ; 
      RECT 30.504 72.208 30.6 108.428 ; 
      RECT 30.312 72.06 30.408 108.244 ; 
      RECT 30.12 71.844 30.216 108.028 ; 
      RECT 29.76 91.624 29.856 92.192 ; 
      RECT 29.088 74.54 29.184 89.916 ; 
      RECT 27.6 80.872 27.696 81.824 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 63.568 181.296 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 63.568 181.296 ; 
  END 
END srambank_128x4x34_6t122 
