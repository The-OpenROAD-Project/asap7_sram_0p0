VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_256x4x32_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_256x4x32_6t122 0 0 ;
  SIZE 30.348 BY 43.2 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1040 1.1720 30.2580 1.2200 ;
        RECT 0.1040 2.2520 30.2580 2.3000 ;
        RECT 0.1040 3.3320 30.2580 3.3800 ;
        RECT 0.1040 4.4120 30.2580 4.4600 ;
        RECT 0.1040 5.4920 30.2580 5.5400 ;
        RECT 0.1040 6.5720 30.2580 6.6200 ;
        RECT 0.1040 7.6520 30.2580 7.7000 ;
        RECT 0.1040 8.7320 30.2580 8.7800 ;
        RECT 0.1040 9.8120 30.2580 9.8600 ;
        RECT 0.1040 10.8920 30.2580 10.9400 ;
        RECT 0.1040 11.9720 30.2580 12.0200 ;
        RECT 0.1040 13.0520 30.2580 13.1000 ;
        RECT 0.1040 14.1320 30.2580 14.1800 ;
        RECT 0.1040 15.2120 30.2580 15.2600 ;
        RECT 0.1040 16.2920 30.2580 16.3400 ;
        RECT 0.1040 17.3720 30.2580 17.4200 ;
        RECT 0.1040 26.5790 30.2580 26.6270 ;
        RECT 0.1040 27.6590 30.2580 27.7070 ;
        RECT 0.1040 28.7390 30.2580 28.7870 ;
        RECT 0.1040 29.8190 30.2580 29.8670 ;
        RECT 0.1040 30.8990 30.2580 30.9470 ;
        RECT 0.1040 31.9790 30.2580 32.0270 ;
        RECT 0.1040 33.0590 30.2580 33.1070 ;
        RECT 0.1040 34.1390 30.2580 34.1870 ;
        RECT 0.1040 35.2190 30.2580 35.2670 ;
        RECT 0.1040 36.2990 30.2580 36.3470 ;
        RECT 0.1040 37.3790 30.2580 37.4270 ;
        RECT 0.1040 38.4590 30.2580 38.5070 ;
        RECT 0.1040 39.5390 30.2580 39.5870 ;
        RECT 0.1040 40.6190 30.2580 40.6670 ;
        RECT 0.1040 41.6990 30.2580 41.7470 ;
        RECT 0.1040 42.7790 30.2580 42.8270 ;
      LAYER M3  ;
        RECT 30.2180 0.2165 30.2360 1.3765 ;
        RECT 16.1960 0.2170 16.2140 1.3760 ;
        RECT 14.7920 0.2530 14.8820 1.3685 ;
        RECT 14.1440 0.2170 14.1620 1.3760 ;
        RECT 0.1220 0.2165 0.1400 1.3765 ;
        RECT 30.2180 1.2965 30.2360 2.4565 ;
        RECT 16.1960 1.2970 16.2140 2.4560 ;
        RECT 14.7920 1.3330 14.8820 2.4485 ;
        RECT 14.1440 1.2970 14.1620 2.4560 ;
        RECT 0.1220 1.2965 0.1400 2.4565 ;
        RECT 30.2180 2.3765 30.2360 3.5365 ;
        RECT 16.1960 2.3770 16.2140 3.5360 ;
        RECT 14.7920 2.4130 14.8820 3.5285 ;
        RECT 14.1440 2.3770 14.1620 3.5360 ;
        RECT 0.1220 2.3765 0.1400 3.5365 ;
        RECT 30.2180 3.4565 30.2360 4.6165 ;
        RECT 16.1960 3.4570 16.2140 4.6160 ;
        RECT 14.7920 3.4930 14.8820 4.6085 ;
        RECT 14.1440 3.4570 14.1620 4.6160 ;
        RECT 0.1220 3.4565 0.1400 4.6165 ;
        RECT 30.2180 4.5365 30.2360 5.6965 ;
        RECT 16.1960 4.5370 16.2140 5.6960 ;
        RECT 14.7920 4.5730 14.8820 5.6885 ;
        RECT 14.1440 4.5370 14.1620 5.6960 ;
        RECT 0.1220 4.5365 0.1400 5.6965 ;
        RECT 30.2180 5.6165 30.2360 6.7765 ;
        RECT 16.1960 5.6170 16.2140 6.7760 ;
        RECT 14.7920 5.6530 14.8820 6.7685 ;
        RECT 14.1440 5.6170 14.1620 6.7760 ;
        RECT 0.1220 5.6165 0.1400 6.7765 ;
        RECT 30.2180 6.6965 30.2360 7.8565 ;
        RECT 16.1960 6.6970 16.2140 7.8560 ;
        RECT 14.7920 6.7330 14.8820 7.8485 ;
        RECT 14.1440 6.6970 14.1620 7.8560 ;
        RECT 0.1220 6.6965 0.1400 7.8565 ;
        RECT 30.2180 7.7765 30.2360 8.9365 ;
        RECT 16.1960 7.7770 16.2140 8.9360 ;
        RECT 14.7920 7.8130 14.8820 8.9285 ;
        RECT 14.1440 7.7770 14.1620 8.9360 ;
        RECT 0.1220 7.7765 0.1400 8.9365 ;
        RECT 30.2180 8.8565 30.2360 10.0165 ;
        RECT 16.1960 8.8570 16.2140 10.0160 ;
        RECT 14.7920 8.8930 14.8820 10.0085 ;
        RECT 14.1440 8.8570 14.1620 10.0160 ;
        RECT 0.1220 8.8565 0.1400 10.0165 ;
        RECT 30.2180 9.9365 30.2360 11.0965 ;
        RECT 16.1960 9.9370 16.2140 11.0960 ;
        RECT 14.7920 9.9730 14.8820 11.0885 ;
        RECT 14.1440 9.9370 14.1620 11.0960 ;
        RECT 0.1220 9.9365 0.1400 11.0965 ;
        RECT 30.2180 11.0165 30.2360 12.1765 ;
        RECT 16.1960 11.0170 16.2140 12.1760 ;
        RECT 14.7920 11.0530 14.8820 12.1685 ;
        RECT 14.1440 11.0170 14.1620 12.1760 ;
        RECT 0.1220 11.0165 0.1400 12.1765 ;
        RECT 30.2180 12.0965 30.2360 13.2565 ;
        RECT 16.1960 12.0970 16.2140 13.2560 ;
        RECT 14.7920 12.1330 14.8820 13.2485 ;
        RECT 14.1440 12.0970 14.1620 13.2560 ;
        RECT 0.1220 12.0965 0.1400 13.2565 ;
        RECT 30.2180 13.1765 30.2360 14.3365 ;
        RECT 16.1960 13.1770 16.2140 14.3360 ;
        RECT 14.7920 13.2130 14.8820 14.3285 ;
        RECT 14.1440 13.1770 14.1620 14.3360 ;
        RECT 0.1220 13.1765 0.1400 14.3365 ;
        RECT 30.2180 14.2565 30.2360 15.4165 ;
        RECT 16.1960 14.2570 16.2140 15.4160 ;
        RECT 14.7920 14.2930 14.8820 15.4085 ;
        RECT 14.1440 14.2570 14.1620 15.4160 ;
        RECT 0.1220 14.2565 0.1400 15.4165 ;
        RECT 30.2180 15.3365 30.2360 16.4965 ;
        RECT 16.1960 15.3370 16.2140 16.4960 ;
        RECT 14.7920 15.3730 14.8820 16.4885 ;
        RECT 14.1440 15.3370 14.1620 16.4960 ;
        RECT 0.1220 15.3365 0.1400 16.4965 ;
        RECT 30.2180 16.4165 30.2360 17.5765 ;
        RECT 16.1960 16.4170 16.2140 17.5760 ;
        RECT 14.7920 16.4530 14.8820 17.5685 ;
        RECT 14.1440 16.4170 14.1620 17.5760 ;
        RECT 0.1220 16.4165 0.1400 17.5765 ;
        RECT 14.0490 21.3650 14.0670 27.4285 ;
        RECT 30.2180 25.6235 30.2360 26.7835 ;
        RECT 16.1960 25.6240 16.2140 26.7830 ;
        RECT 14.7920 25.6600 14.8820 26.7755 ;
        RECT 14.1440 25.6240 14.1620 26.7830 ;
        RECT 0.1220 25.6235 0.1400 26.7835 ;
        RECT 30.2180 26.7035 30.2360 27.8635 ;
        RECT 16.1960 26.7040 16.2140 27.8630 ;
        RECT 14.7920 26.7400 14.8820 27.8555 ;
        RECT 14.1440 26.7040 14.1620 27.8630 ;
        RECT 0.1220 26.7035 0.1400 27.8635 ;
        RECT 30.2180 27.7835 30.2360 28.9435 ;
        RECT 16.1960 27.7840 16.2140 28.9430 ;
        RECT 14.7920 27.8200 14.8820 28.9355 ;
        RECT 14.1440 27.7840 14.1620 28.9430 ;
        RECT 0.1220 27.7835 0.1400 28.9435 ;
        RECT 30.2180 28.8635 30.2360 30.0235 ;
        RECT 16.1960 28.8640 16.2140 30.0230 ;
        RECT 14.7920 28.9000 14.8820 30.0155 ;
        RECT 14.1440 28.8640 14.1620 30.0230 ;
        RECT 0.1220 28.8635 0.1400 30.0235 ;
        RECT 30.2180 29.9435 30.2360 31.1035 ;
        RECT 16.1960 29.9440 16.2140 31.1030 ;
        RECT 14.7920 29.9800 14.8820 31.0955 ;
        RECT 14.1440 29.9440 14.1620 31.1030 ;
        RECT 0.1220 29.9435 0.1400 31.1035 ;
        RECT 30.2180 31.0235 30.2360 32.1835 ;
        RECT 16.1960 31.0240 16.2140 32.1830 ;
        RECT 14.7920 31.0600 14.8820 32.1755 ;
        RECT 14.1440 31.0240 14.1620 32.1830 ;
        RECT 0.1220 31.0235 0.1400 32.1835 ;
        RECT 30.2180 32.1035 30.2360 33.2635 ;
        RECT 16.1960 32.1040 16.2140 33.2630 ;
        RECT 14.7920 32.1400 14.8820 33.2555 ;
        RECT 14.1440 32.1040 14.1620 33.2630 ;
        RECT 0.1220 32.1035 0.1400 33.2635 ;
        RECT 30.2180 33.1835 30.2360 34.3435 ;
        RECT 16.1960 33.1840 16.2140 34.3430 ;
        RECT 14.7920 33.2200 14.8820 34.3355 ;
        RECT 14.1440 33.1840 14.1620 34.3430 ;
        RECT 0.1220 33.1835 0.1400 34.3435 ;
        RECT 30.2180 34.2635 30.2360 35.4235 ;
        RECT 16.1960 34.2640 16.2140 35.4230 ;
        RECT 14.7920 34.3000 14.8820 35.4155 ;
        RECT 14.1440 34.2640 14.1620 35.4230 ;
        RECT 0.1220 34.2635 0.1400 35.4235 ;
        RECT 30.2180 35.3435 30.2360 36.5035 ;
        RECT 16.1960 35.3440 16.2140 36.5030 ;
        RECT 14.7920 35.3800 14.8820 36.4955 ;
        RECT 14.1440 35.3440 14.1620 36.5030 ;
        RECT 0.1220 35.3435 0.1400 36.5035 ;
        RECT 30.2180 36.4235 30.2360 37.5835 ;
        RECT 16.1960 36.4240 16.2140 37.5830 ;
        RECT 14.7920 36.4600 14.8820 37.5755 ;
        RECT 14.1440 36.4240 14.1620 37.5830 ;
        RECT 0.1220 36.4235 0.1400 37.5835 ;
        RECT 30.2180 37.5035 30.2360 38.6635 ;
        RECT 16.1960 37.5040 16.2140 38.6630 ;
        RECT 14.7920 37.5400 14.8820 38.6555 ;
        RECT 14.1440 37.5040 14.1620 38.6630 ;
        RECT 0.1220 37.5035 0.1400 38.6635 ;
        RECT 30.2180 38.5835 30.2360 39.7435 ;
        RECT 16.1960 38.5840 16.2140 39.7430 ;
        RECT 14.7920 38.6200 14.8820 39.7355 ;
        RECT 14.1440 38.5840 14.1620 39.7430 ;
        RECT 0.1220 38.5835 0.1400 39.7435 ;
        RECT 30.2180 39.6635 30.2360 40.8235 ;
        RECT 16.1960 39.6640 16.2140 40.8230 ;
        RECT 14.7920 39.7000 14.8820 40.8155 ;
        RECT 14.1440 39.6640 14.1620 40.8230 ;
        RECT 0.1220 39.6635 0.1400 40.8235 ;
        RECT 30.2180 40.7435 30.2360 41.9035 ;
        RECT 16.1960 40.7440 16.2140 41.9030 ;
        RECT 14.7920 40.7800 14.8820 41.8955 ;
        RECT 14.1440 40.7440 14.1620 41.9030 ;
        RECT 0.1220 40.7435 0.1400 41.9035 ;
        RECT 30.2180 41.8235 30.2360 42.9835 ;
        RECT 16.1960 41.8240 16.2140 42.9830 ;
        RECT 14.7920 41.8600 14.8820 42.9755 ;
        RECT 14.1440 41.8240 14.1620 42.9830 ;
        RECT 0.1220 41.8235 0.1400 42.9835 ;
      LAYER V3  ;
        RECT 0.1220 1.1720 0.1400 1.2200 ;
        RECT 14.1440 1.1720 14.1620 1.2200 ;
        RECT 14.7920 1.1720 14.8820 1.2200 ;
        RECT 16.1960 1.1720 16.2140 1.2200 ;
        RECT 30.2180 1.1720 30.2360 1.2200 ;
        RECT 0.1220 2.2520 0.1400 2.3000 ;
        RECT 14.1440 2.2520 14.1620 2.3000 ;
        RECT 14.7920 2.2520 14.8820 2.3000 ;
        RECT 16.1960 2.2520 16.2140 2.3000 ;
        RECT 30.2180 2.2520 30.2360 2.3000 ;
        RECT 0.1220 3.3320 0.1400 3.3800 ;
        RECT 14.1440 3.3320 14.1620 3.3800 ;
        RECT 14.7920 3.3320 14.8820 3.3800 ;
        RECT 16.1960 3.3320 16.2140 3.3800 ;
        RECT 30.2180 3.3320 30.2360 3.3800 ;
        RECT 0.1220 4.4120 0.1400 4.4600 ;
        RECT 14.1440 4.4120 14.1620 4.4600 ;
        RECT 14.7920 4.4120 14.8820 4.4600 ;
        RECT 16.1960 4.4120 16.2140 4.4600 ;
        RECT 30.2180 4.4120 30.2360 4.4600 ;
        RECT 0.1220 5.4920 0.1400 5.5400 ;
        RECT 14.1440 5.4920 14.1620 5.5400 ;
        RECT 14.7920 5.4920 14.8820 5.5400 ;
        RECT 16.1960 5.4920 16.2140 5.5400 ;
        RECT 30.2180 5.4920 30.2360 5.5400 ;
        RECT 0.1220 6.5720 0.1400 6.6200 ;
        RECT 14.1440 6.5720 14.1620 6.6200 ;
        RECT 14.7920 6.5720 14.8820 6.6200 ;
        RECT 16.1960 6.5720 16.2140 6.6200 ;
        RECT 30.2180 6.5720 30.2360 6.6200 ;
        RECT 0.1220 7.6520 0.1400 7.7000 ;
        RECT 14.1440 7.6520 14.1620 7.7000 ;
        RECT 14.7920 7.6520 14.8820 7.7000 ;
        RECT 16.1960 7.6520 16.2140 7.7000 ;
        RECT 30.2180 7.6520 30.2360 7.7000 ;
        RECT 0.1220 8.7320 0.1400 8.7800 ;
        RECT 14.1440 8.7320 14.1620 8.7800 ;
        RECT 14.7920 8.7320 14.8820 8.7800 ;
        RECT 16.1960 8.7320 16.2140 8.7800 ;
        RECT 30.2180 8.7320 30.2360 8.7800 ;
        RECT 0.1220 9.8120 0.1400 9.8600 ;
        RECT 14.1440 9.8120 14.1620 9.8600 ;
        RECT 14.7920 9.8120 14.8820 9.8600 ;
        RECT 16.1960 9.8120 16.2140 9.8600 ;
        RECT 30.2180 9.8120 30.2360 9.8600 ;
        RECT 0.1220 10.8920 0.1400 10.9400 ;
        RECT 14.1440 10.8920 14.1620 10.9400 ;
        RECT 14.7920 10.8920 14.8820 10.9400 ;
        RECT 16.1960 10.8920 16.2140 10.9400 ;
        RECT 30.2180 10.8920 30.2360 10.9400 ;
        RECT 0.1220 11.9720 0.1400 12.0200 ;
        RECT 14.1440 11.9720 14.1620 12.0200 ;
        RECT 14.7920 11.9720 14.8820 12.0200 ;
        RECT 16.1960 11.9720 16.2140 12.0200 ;
        RECT 30.2180 11.9720 30.2360 12.0200 ;
        RECT 0.1220 13.0520 0.1400 13.1000 ;
        RECT 14.1440 13.0520 14.1620 13.1000 ;
        RECT 14.7920 13.0520 14.8820 13.1000 ;
        RECT 16.1960 13.0520 16.2140 13.1000 ;
        RECT 30.2180 13.0520 30.2360 13.1000 ;
        RECT 0.1220 14.1320 0.1400 14.1800 ;
        RECT 14.1440 14.1320 14.1620 14.1800 ;
        RECT 14.7920 14.1320 14.8820 14.1800 ;
        RECT 16.1960 14.1320 16.2140 14.1800 ;
        RECT 30.2180 14.1320 30.2360 14.1800 ;
        RECT 0.1220 15.2120 0.1400 15.2600 ;
        RECT 14.1440 15.2120 14.1620 15.2600 ;
        RECT 14.7920 15.2120 14.8820 15.2600 ;
        RECT 16.1960 15.2120 16.2140 15.2600 ;
        RECT 30.2180 15.2120 30.2360 15.2600 ;
        RECT 0.1220 16.2920 0.1400 16.3400 ;
        RECT 14.1440 16.2920 14.1620 16.3400 ;
        RECT 14.7920 16.2920 14.8820 16.3400 ;
        RECT 16.1960 16.2920 16.2140 16.3400 ;
        RECT 30.2180 16.2920 30.2360 16.3400 ;
        RECT 0.1220 17.3720 0.1400 17.4200 ;
        RECT 14.1440 17.3720 14.1620 17.4200 ;
        RECT 14.7920 17.3720 14.8820 17.4200 ;
        RECT 16.1960 17.3720 16.2140 17.4200 ;
        RECT 30.2180 17.3720 30.2360 17.4200 ;
        RECT 0.1220 26.5790 0.1400 26.6270 ;
        RECT 14.1440 26.5790 14.1620 26.6270 ;
        RECT 14.7920 26.5790 14.8820 26.6270 ;
        RECT 16.1960 26.5790 16.2140 26.6270 ;
        RECT 30.2180 26.5790 30.2360 26.6270 ;
        RECT 0.1220 27.6590 0.1400 27.7070 ;
        RECT 14.1440 27.6590 14.1620 27.7070 ;
        RECT 14.7920 27.6590 14.8820 27.7070 ;
        RECT 16.1960 27.6590 16.2140 27.7070 ;
        RECT 30.2180 27.6590 30.2360 27.7070 ;
        RECT 0.1220 28.7390 0.1400 28.7870 ;
        RECT 14.1440 28.7390 14.1620 28.7870 ;
        RECT 14.7920 28.7390 14.8820 28.7870 ;
        RECT 16.1960 28.7390 16.2140 28.7870 ;
        RECT 30.2180 28.7390 30.2360 28.7870 ;
        RECT 0.1220 29.8190 0.1400 29.8670 ;
        RECT 14.1440 29.8190 14.1620 29.8670 ;
        RECT 14.7920 29.8190 14.8820 29.8670 ;
        RECT 16.1960 29.8190 16.2140 29.8670 ;
        RECT 30.2180 29.8190 30.2360 29.8670 ;
        RECT 0.1220 30.8990 0.1400 30.9470 ;
        RECT 14.1440 30.8990 14.1620 30.9470 ;
        RECT 14.7920 30.8990 14.8820 30.9470 ;
        RECT 16.1960 30.8990 16.2140 30.9470 ;
        RECT 30.2180 30.8990 30.2360 30.9470 ;
        RECT 0.1220 31.9790 0.1400 32.0270 ;
        RECT 14.1440 31.9790 14.1620 32.0270 ;
        RECT 14.7920 31.9790 14.8820 32.0270 ;
        RECT 16.1960 31.9790 16.2140 32.0270 ;
        RECT 30.2180 31.9790 30.2360 32.0270 ;
        RECT 0.1220 33.0590 0.1400 33.1070 ;
        RECT 14.1440 33.0590 14.1620 33.1070 ;
        RECT 14.7920 33.0590 14.8820 33.1070 ;
        RECT 16.1960 33.0590 16.2140 33.1070 ;
        RECT 30.2180 33.0590 30.2360 33.1070 ;
        RECT 0.1220 34.1390 0.1400 34.1870 ;
        RECT 14.1440 34.1390 14.1620 34.1870 ;
        RECT 14.7920 34.1390 14.8820 34.1870 ;
        RECT 16.1960 34.1390 16.2140 34.1870 ;
        RECT 30.2180 34.1390 30.2360 34.1870 ;
        RECT 0.1220 35.2190 0.1400 35.2670 ;
        RECT 14.1440 35.2190 14.1620 35.2670 ;
        RECT 14.7920 35.2190 14.8820 35.2670 ;
        RECT 16.1960 35.2190 16.2140 35.2670 ;
        RECT 30.2180 35.2190 30.2360 35.2670 ;
        RECT 0.1220 36.2990 0.1400 36.3470 ;
        RECT 14.1440 36.2990 14.1620 36.3470 ;
        RECT 14.7920 36.2990 14.8820 36.3470 ;
        RECT 16.1960 36.2990 16.2140 36.3470 ;
        RECT 30.2180 36.2990 30.2360 36.3470 ;
        RECT 0.1220 37.3790 0.1400 37.4270 ;
        RECT 14.1440 37.3790 14.1620 37.4270 ;
        RECT 14.7920 37.3790 14.8820 37.4270 ;
        RECT 16.1960 37.3790 16.2140 37.4270 ;
        RECT 30.2180 37.3790 30.2360 37.4270 ;
        RECT 0.1220 38.4590 0.1400 38.5070 ;
        RECT 14.1440 38.4590 14.1620 38.5070 ;
        RECT 14.7920 38.4590 14.8820 38.5070 ;
        RECT 16.1960 38.4590 16.2140 38.5070 ;
        RECT 30.2180 38.4590 30.2360 38.5070 ;
        RECT 0.1220 39.5390 0.1400 39.5870 ;
        RECT 14.1440 39.5390 14.1620 39.5870 ;
        RECT 14.7920 39.5390 14.8820 39.5870 ;
        RECT 16.1960 39.5390 16.2140 39.5870 ;
        RECT 30.2180 39.5390 30.2360 39.5870 ;
        RECT 0.1220 40.6190 0.1400 40.6670 ;
        RECT 14.1440 40.6190 14.1620 40.6670 ;
        RECT 14.7920 40.6190 14.8820 40.6670 ;
        RECT 16.1960 40.6190 16.2140 40.6670 ;
        RECT 30.2180 40.6190 30.2360 40.6670 ;
        RECT 0.1220 41.6990 0.1400 41.7470 ;
        RECT 14.1440 41.6990 14.1620 41.7470 ;
        RECT 14.7920 41.6990 14.8820 41.7470 ;
        RECT 16.1960 41.6990 16.2140 41.7470 ;
        RECT 30.2180 41.6990 30.2360 41.7470 ;
        RECT 0.1220 42.7790 0.1400 42.8270 ;
        RECT 14.1440 42.7790 14.1620 42.8270 ;
        RECT 14.7920 42.7790 14.8820 42.8270 ;
        RECT 16.1960 42.7790 16.2140 42.8270 ;
        RECT 30.2180 42.7790 30.2360 42.8270 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1040 1.0760 30.2580 1.1240 ;
        RECT 0.1040 2.1560 30.2580 2.2040 ;
        RECT 0.1040 3.2360 30.2580 3.2840 ;
        RECT 0.1040 4.3160 30.2580 4.3640 ;
        RECT 0.1040 5.3960 30.2580 5.4440 ;
        RECT 0.1040 6.4760 30.2580 6.5240 ;
        RECT 0.1040 7.5560 30.2580 7.6040 ;
        RECT 0.1040 8.6360 30.2580 8.6840 ;
        RECT 0.1040 9.7160 30.2580 9.7640 ;
        RECT 0.1040 10.7960 30.2580 10.8440 ;
        RECT 0.1040 11.8760 30.2580 11.9240 ;
        RECT 0.1040 12.9560 30.2580 13.0040 ;
        RECT 0.1040 14.0360 30.2580 14.0840 ;
        RECT 0.1040 15.1160 30.2580 15.1640 ;
        RECT 0.1040 16.1960 30.2580 16.2440 ;
        RECT 0.1040 17.2760 30.2580 17.3240 ;
        RECT 10.4760 18.3415 19.8720 18.5575 ;
        RECT 14.3100 21.5095 16.0380 21.7255 ;
        RECT 14.3100 24.6775 16.0380 24.8935 ;
        RECT 0.1040 26.4830 30.2580 26.5310 ;
        RECT 0.1040 27.5630 30.2580 27.6110 ;
        RECT 0.1040 28.6430 30.2580 28.6910 ;
        RECT 0.1040 29.7230 30.2580 29.7710 ;
        RECT 0.1040 30.8030 30.2580 30.8510 ;
        RECT 0.1040 31.8830 30.2580 31.9310 ;
        RECT 0.1040 32.9630 30.2580 33.0110 ;
        RECT 0.1040 34.0430 30.2580 34.0910 ;
        RECT 0.1040 35.1230 30.2580 35.1710 ;
        RECT 0.1040 36.2030 30.2580 36.2510 ;
        RECT 0.1040 37.2830 30.2580 37.3310 ;
        RECT 0.1040 38.3630 30.2580 38.4110 ;
        RECT 0.1040 39.4430 30.2580 39.4910 ;
        RECT 0.1040 40.5230 30.2580 40.5710 ;
        RECT 0.1040 41.6030 30.2580 41.6510 ;
        RECT 0.1040 42.6830 30.2580 42.7310 ;
      LAYER M3  ;
        RECT 30.1820 0.2165 30.2000 1.3765 ;
        RECT 16.2500 0.2165 16.2680 1.3765 ;
        RECT 15.4850 0.2530 15.5210 1.3675 ;
        RECT 15.2600 0.2530 15.2870 1.3675 ;
        RECT 14.0900 0.2165 14.1080 1.3765 ;
        RECT 0.1580 0.2165 0.1760 1.3765 ;
        RECT 30.1820 1.2965 30.2000 2.4565 ;
        RECT 16.2500 1.2965 16.2680 2.4565 ;
        RECT 15.4850 1.3330 15.5210 2.4475 ;
        RECT 15.2600 1.3330 15.2870 2.4475 ;
        RECT 14.0900 1.2965 14.1080 2.4565 ;
        RECT 0.1580 1.2965 0.1760 2.4565 ;
        RECT 30.1820 2.3765 30.2000 3.5365 ;
        RECT 16.2500 2.3765 16.2680 3.5365 ;
        RECT 15.4850 2.4130 15.5210 3.5275 ;
        RECT 15.2600 2.4130 15.2870 3.5275 ;
        RECT 14.0900 2.3765 14.1080 3.5365 ;
        RECT 0.1580 2.3765 0.1760 3.5365 ;
        RECT 30.1820 3.4565 30.2000 4.6165 ;
        RECT 16.2500 3.4565 16.2680 4.6165 ;
        RECT 15.4850 3.4930 15.5210 4.6075 ;
        RECT 15.2600 3.4930 15.2870 4.6075 ;
        RECT 14.0900 3.4565 14.1080 4.6165 ;
        RECT 0.1580 3.4565 0.1760 4.6165 ;
        RECT 30.1820 4.5365 30.2000 5.6965 ;
        RECT 16.2500 4.5365 16.2680 5.6965 ;
        RECT 15.4850 4.5730 15.5210 5.6875 ;
        RECT 15.2600 4.5730 15.2870 5.6875 ;
        RECT 14.0900 4.5365 14.1080 5.6965 ;
        RECT 0.1580 4.5365 0.1760 5.6965 ;
        RECT 30.1820 5.6165 30.2000 6.7765 ;
        RECT 16.2500 5.6165 16.2680 6.7765 ;
        RECT 15.4850 5.6530 15.5210 6.7675 ;
        RECT 15.2600 5.6530 15.2870 6.7675 ;
        RECT 14.0900 5.6165 14.1080 6.7765 ;
        RECT 0.1580 5.6165 0.1760 6.7765 ;
        RECT 30.1820 6.6965 30.2000 7.8565 ;
        RECT 16.2500 6.6965 16.2680 7.8565 ;
        RECT 15.4850 6.7330 15.5210 7.8475 ;
        RECT 15.2600 6.7330 15.2870 7.8475 ;
        RECT 14.0900 6.6965 14.1080 7.8565 ;
        RECT 0.1580 6.6965 0.1760 7.8565 ;
        RECT 30.1820 7.7765 30.2000 8.9365 ;
        RECT 16.2500 7.7765 16.2680 8.9365 ;
        RECT 15.4850 7.8130 15.5210 8.9275 ;
        RECT 15.2600 7.8130 15.2870 8.9275 ;
        RECT 14.0900 7.7765 14.1080 8.9365 ;
        RECT 0.1580 7.7765 0.1760 8.9365 ;
        RECT 30.1820 8.8565 30.2000 10.0165 ;
        RECT 16.2500 8.8565 16.2680 10.0165 ;
        RECT 15.4850 8.8930 15.5210 10.0075 ;
        RECT 15.2600 8.8930 15.2870 10.0075 ;
        RECT 14.0900 8.8565 14.1080 10.0165 ;
        RECT 0.1580 8.8565 0.1760 10.0165 ;
        RECT 30.1820 9.9365 30.2000 11.0965 ;
        RECT 16.2500 9.9365 16.2680 11.0965 ;
        RECT 15.4850 9.9730 15.5210 11.0875 ;
        RECT 15.2600 9.9730 15.2870 11.0875 ;
        RECT 14.0900 9.9365 14.1080 11.0965 ;
        RECT 0.1580 9.9365 0.1760 11.0965 ;
        RECT 30.1820 11.0165 30.2000 12.1765 ;
        RECT 16.2500 11.0165 16.2680 12.1765 ;
        RECT 15.4850 11.0530 15.5210 12.1675 ;
        RECT 15.2600 11.0530 15.2870 12.1675 ;
        RECT 14.0900 11.0165 14.1080 12.1765 ;
        RECT 0.1580 11.0165 0.1760 12.1765 ;
        RECT 30.1820 12.0965 30.2000 13.2565 ;
        RECT 16.2500 12.0965 16.2680 13.2565 ;
        RECT 15.4850 12.1330 15.5210 13.2475 ;
        RECT 15.2600 12.1330 15.2870 13.2475 ;
        RECT 14.0900 12.0965 14.1080 13.2565 ;
        RECT 0.1580 12.0965 0.1760 13.2565 ;
        RECT 30.1820 13.1765 30.2000 14.3365 ;
        RECT 16.2500 13.1765 16.2680 14.3365 ;
        RECT 15.4850 13.2130 15.5210 14.3275 ;
        RECT 15.2600 13.2130 15.2870 14.3275 ;
        RECT 14.0900 13.1765 14.1080 14.3365 ;
        RECT 0.1580 13.1765 0.1760 14.3365 ;
        RECT 30.1820 14.2565 30.2000 15.4165 ;
        RECT 16.2500 14.2565 16.2680 15.4165 ;
        RECT 15.4850 14.2930 15.5210 15.4075 ;
        RECT 15.2600 14.2930 15.2870 15.4075 ;
        RECT 14.0900 14.2565 14.1080 15.4165 ;
        RECT 0.1580 14.2565 0.1760 15.4165 ;
        RECT 30.1820 15.3365 30.2000 16.4965 ;
        RECT 16.2500 15.3365 16.2680 16.4965 ;
        RECT 15.4850 15.3730 15.5210 16.4875 ;
        RECT 15.2600 15.3730 15.2870 16.4875 ;
        RECT 14.0900 15.3365 14.1080 16.4965 ;
        RECT 0.1580 15.3365 0.1760 16.4965 ;
        RECT 30.1820 16.4165 30.2000 17.5765 ;
        RECT 16.2500 16.4165 16.2680 17.5765 ;
        RECT 15.4850 16.4530 15.5210 17.5675 ;
        RECT 15.2600 16.4530 15.2870 17.5675 ;
        RECT 14.0900 16.4165 14.1080 17.5765 ;
        RECT 0.1580 16.4165 0.1760 17.5765 ;
        RECT 16.2450 17.5470 16.2630 25.7540 ;
        RECT 15.2910 17.7705 15.5250 25.4535 ;
        RECT 14.0850 17.5470 14.1030 27.4285 ;
        RECT 30.1820 25.6235 30.2000 26.7835 ;
        RECT 16.2500 25.6235 16.2680 26.7835 ;
        RECT 15.4850 25.6600 15.5210 26.7745 ;
        RECT 15.2600 25.6600 15.2870 26.7745 ;
        RECT 14.0900 25.6235 14.1080 26.7835 ;
        RECT 0.1580 25.6235 0.1760 26.7835 ;
        RECT 30.1820 26.7035 30.2000 27.8635 ;
        RECT 16.2500 26.7035 16.2680 27.8635 ;
        RECT 15.4850 26.7400 15.5210 27.8545 ;
        RECT 15.2600 26.7400 15.2870 27.8545 ;
        RECT 14.0900 26.7035 14.1080 27.8635 ;
        RECT 0.1580 26.7035 0.1760 27.8635 ;
        RECT 30.1820 27.7835 30.2000 28.9435 ;
        RECT 16.2500 27.7835 16.2680 28.9435 ;
        RECT 15.4850 27.8200 15.5210 28.9345 ;
        RECT 15.2600 27.8200 15.2870 28.9345 ;
        RECT 14.0900 27.7835 14.1080 28.9435 ;
        RECT 0.1580 27.7835 0.1760 28.9435 ;
        RECT 30.1820 28.8635 30.2000 30.0235 ;
        RECT 16.2500 28.8635 16.2680 30.0235 ;
        RECT 15.4850 28.9000 15.5210 30.0145 ;
        RECT 15.2600 28.9000 15.2870 30.0145 ;
        RECT 14.0900 28.8635 14.1080 30.0235 ;
        RECT 0.1580 28.8635 0.1760 30.0235 ;
        RECT 30.1820 29.9435 30.2000 31.1035 ;
        RECT 16.2500 29.9435 16.2680 31.1035 ;
        RECT 15.4850 29.9800 15.5210 31.0945 ;
        RECT 15.2600 29.9800 15.2870 31.0945 ;
        RECT 14.0900 29.9435 14.1080 31.1035 ;
        RECT 0.1580 29.9435 0.1760 31.1035 ;
        RECT 30.1820 31.0235 30.2000 32.1835 ;
        RECT 16.2500 31.0235 16.2680 32.1835 ;
        RECT 15.4850 31.0600 15.5210 32.1745 ;
        RECT 15.2600 31.0600 15.2870 32.1745 ;
        RECT 14.0900 31.0235 14.1080 32.1835 ;
        RECT 0.1580 31.0235 0.1760 32.1835 ;
        RECT 30.1820 32.1035 30.2000 33.2635 ;
        RECT 16.2500 32.1035 16.2680 33.2635 ;
        RECT 15.4850 32.1400 15.5210 33.2545 ;
        RECT 15.2600 32.1400 15.2870 33.2545 ;
        RECT 14.0900 32.1035 14.1080 33.2635 ;
        RECT 0.1580 32.1035 0.1760 33.2635 ;
        RECT 30.1820 33.1835 30.2000 34.3435 ;
        RECT 16.2500 33.1835 16.2680 34.3435 ;
        RECT 15.4850 33.2200 15.5210 34.3345 ;
        RECT 15.2600 33.2200 15.2870 34.3345 ;
        RECT 14.0900 33.1835 14.1080 34.3435 ;
        RECT 0.1580 33.1835 0.1760 34.3435 ;
        RECT 30.1820 34.2635 30.2000 35.4235 ;
        RECT 16.2500 34.2635 16.2680 35.4235 ;
        RECT 15.4850 34.3000 15.5210 35.4145 ;
        RECT 15.2600 34.3000 15.2870 35.4145 ;
        RECT 14.0900 34.2635 14.1080 35.4235 ;
        RECT 0.1580 34.2635 0.1760 35.4235 ;
        RECT 30.1820 35.3435 30.2000 36.5035 ;
        RECT 16.2500 35.3435 16.2680 36.5035 ;
        RECT 15.4850 35.3800 15.5210 36.4945 ;
        RECT 15.2600 35.3800 15.2870 36.4945 ;
        RECT 14.0900 35.3435 14.1080 36.5035 ;
        RECT 0.1580 35.3435 0.1760 36.5035 ;
        RECT 30.1820 36.4235 30.2000 37.5835 ;
        RECT 16.2500 36.4235 16.2680 37.5835 ;
        RECT 15.4850 36.4600 15.5210 37.5745 ;
        RECT 15.2600 36.4600 15.2870 37.5745 ;
        RECT 14.0900 36.4235 14.1080 37.5835 ;
        RECT 0.1580 36.4235 0.1760 37.5835 ;
        RECT 30.1820 37.5035 30.2000 38.6635 ;
        RECT 16.2500 37.5035 16.2680 38.6635 ;
        RECT 15.4850 37.5400 15.5210 38.6545 ;
        RECT 15.2600 37.5400 15.2870 38.6545 ;
        RECT 14.0900 37.5035 14.1080 38.6635 ;
        RECT 0.1580 37.5035 0.1760 38.6635 ;
        RECT 30.1820 38.5835 30.2000 39.7435 ;
        RECT 16.2500 38.5835 16.2680 39.7435 ;
        RECT 15.4850 38.6200 15.5210 39.7345 ;
        RECT 15.2600 38.6200 15.2870 39.7345 ;
        RECT 14.0900 38.5835 14.1080 39.7435 ;
        RECT 0.1580 38.5835 0.1760 39.7435 ;
        RECT 30.1820 39.6635 30.2000 40.8235 ;
        RECT 16.2500 39.6635 16.2680 40.8235 ;
        RECT 15.4850 39.7000 15.5210 40.8145 ;
        RECT 15.2600 39.7000 15.2870 40.8145 ;
        RECT 14.0900 39.6635 14.1080 40.8235 ;
        RECT 0.1580 39.6635 0.1760 40.8235 ;
        RECT 30.1820 40.7435 30.2000 41.9035 ;
        RECT 16.2500 40.7435 16.2680 41.9035 ;
        RECT 15.4850 40.7800 15.5210 41.8945 ;
        RECT 15.2600 40.7800 15.2870 41.8945 ;
        RECT 14.0900 40.7435 14.1080 41.9035 ;
        RECT 0.1580 40.7435 0.1760 41.9035 ;
        RECT 30.1820 41.8235 30.2000 42.9835 ;
        RECT 16.2500 41.8235 16.2680 42.9835 ;
        RECT 15.4850 41.8600 15.5210 42.9745 ;
        RECT 15.2600 41.8600 15.2870 42.9745 ;
        RECT 14.0900 41.8235 14.1080 42.9835 ;
        RECT 0.1580 41.8235 0.1760 42.9835 ;
      LAYER V3  ;
        RECT 0.1580 1.0760 0.1760 1.1240 ;
        RECT 14.0900 1.0760 14.1080 1.1240 ;
        RECT 15.2600 1.0760 15.2870 1.1240 ;
        RECT 15.4850 1.0760 15.5210 1.1240 ;
        RECT 16.2500 1.0760 16.2680 1.1240 ;
        RECT 30.1820 1.0760 30.2000 1.1240 ;
        RECT 0.1580 2.1560 0.1760 2.2040 ;
        RECT 14.0900 2.1560 14.1080 2.2040 ;
        RECT 15.2600 2.1560 15.2870 2.2040 ;
        RECT 15.4850 2.1560 15.5210 2.2040 ;
        RECT 16.2500 2.1560 16.2680 2.2040 ;
        RECT 30.1820 2.1560 30.2000 2.2040 ;
        RECT 0.1580 3.2360 0.1760 3.2840 ;
        RECT 14.0900 3.2360 14.1080 3.2840 ;
        RECT 15.2600 3.2360 15.2870 3.2840 ;
        RECT 15.4850 3.2360 15.5210 3.2840 ;
        RECT 16.2500 3.2360 16.2680 3.2840 ;
        RECT 30.1820 3.2360 30.2000 3.2840 ;
        RECT 0.1580 4.3160 0.1760 4.3640 ;
        RECT 14.0900 4.3160 14.1080 4.3640 ;
        RECT 15.2600 4.3160 15.2870 4.3640 ;
        RECT 15.4850 4.3160 15.5210 4.3640 ;
        RECT 16.2500 4.3160 16.2680 4.3640 ;
        RECT 30.1820 4.3160 30.2000 4.3640 ;
        RECT 0.1580 5.3960 0.1760 5.4440 ;
        RECT 14.0900 5.3960 14.1080 5.4440 ;
        RECT 15.2600 5.3960 15.2870 5.4440 ;
        RECT 15.4850 5.3960 15.5210 5.4440 ;
        RECT 16.2500 5.3960 16.2680 5.4440 ;
        RECT 30.1820 5.3960 30.2000 5.4440 ;
        RECT 0.1580 6.4760 0.1760 6.5240 ;
        RECT 14.0900 6.4760 14.1080 6.5240 ;
        RECT 15.2600 6.4760 15.2870 6.5240 ;
        RECT 15.4850 6.4760 15.5210 6.5240 ;
        RECT 16.2500 6.4760 16.2680 6.5240 ;
        RECT 30.1820 6.4760 30.2000 6.5240 ;
        RECT 0.1580 7.5560 0.1760 7.6040 ;
        RECT 14.0900 7.5560 14.1080 7.6040 ;
        RECT 15.2600 7.5560 15.2870 7.6040 ;
        RECT 15.4850 7.5560 15.5210 7.6040 ;
        RECT 16.2500 7.5560 16.2680 7.6040 ;
        RECT 30.1820 7.5560 30.2000 7.6040 ;
        RECT 0.1580 8.6360 0.1760 8.6840 ;
        RECT 14.0900 8.6360 14.1080 8.6840 ;
        RECT 15.2600 8.6360 15.2870 8.6840 ;
        RECT 15.4850 8.6360 15.5210 8.6840 ;
        RECT 16.2500 8.6360 16.2680 8.6840 ;
        RECT 30.1820 8.6360 30.2000 8.6840 ;
        RECT 0.1580 9.7160 0.1760 9.7640 ;
        RECT 14.0900 9.7160 14.1080 9.7640 ;
        RECT 15.2600 9.7160 15.2870 9.7640 ;
        RECT 15.4850 9.7160 15.5210 9.7640 ;
        RECT 16.2500 9.7160 16.2680 9.7640 ;
        RECT 30.1820 9.7160 30.2000 9.7640 ;
        RECT 0.1580 10.7960 0.1760 10.8440 ;
        RECT 14.0900 10.7960 14.1080 10.8440 ;
        RECT 15.2600 10.7960 15.2870 10.8440 ;
        RECT 15.4850 10.7960 15.5210 10.8440 ;
        RECT 16.2500 10.7960 16.2680 10.8440 ;
        RECT 30.1820 10.7960 30.2000 10.8440 ;
        RECT 0.1580 11.8760 0.1760 11.9240 ;
        RECT 14.0900 11.8760 14.1080 11.9240 ;
        RECT 15.2600 11.8760 15.2870 11.9240 ;
        RECT 15.4850 11.8760 15.5210 11.9240 ;
        RECT 16.2500 11.8760 16.2680 11.9240 ;
        RECT 30.1820 11.8760 30.2000 11.9240 ;
        RECT 0.1580 12.9560 0.1760 13.0040 ;
        RECT 14.0900 12.9560 14.1080 13.0040 ;
        RECT 15.2600 12.9560 15.2870 13.0040 ;
        RECT 15.4850 12.9560 15.5210 13.0040 ;
        RECT 16.2500 12.9560 16.2680 13.0040 ;
        RECT 30.1820 12.9560 30.2000 13.0040 ;
        RECT 0.1580 14.0360 0.1760 14.0840 ;
        RECT 14.0900 14.0360 14.1080 14.0840 ;
        RECT 15.2600 14.0360 15.2870 14.0840 ;
        RECT 15.4850 14.0360 15.5210 14.0840 ;
        RECT 16.2500 14.0360 16.2680 14.0840 ;
        RECT 30.1820 14.0360 30.2000 14.0840 ;
        RECT 0.1580 15.1160 0.1760 15.1640 ;
        RECT 14.0900 15.1160 14.1080 15.1640 ;
        RECT 15.2600 15.1160 15.2870 15.1640 ;
        RECT 15.4850 15.1160 15.5210 15.1640 ;
        RECT 16.2500 15.1160 16.2680 15.1640 ;
        RECT 30.1820 15.1160 30.2000 15.1640 ;
        RECT 0.1580 16.1960 0.1760 16.2440 ;
        RECT 14.0900 16.1960 14.1080 16.2440 ;
        RECT 15.2600 16.1960 15.2870 16.2440 ;
        RECT 15.4850 16.1960 15.5210 16.2440 ;
        RECT 16.2500 16.1960 16.2680 16.2440 ;
        RECT 30.1820 16.1960 30.2000 16.2440 ;
        RECT 0.1580 17.2760 0.1760 17.3240 ;
        RECT 14.0900 17.2760 14.1080 17.3240 ;
        RECT 15.2600 17.2760 15.2870 17.3240 ;
        RECT 15.4850 17.2760 15.5210 17.3240 ;
        RECT 16.2500 17.2760 16.2680 17.3240 ;
        RECT 30.1820 17.2760 30.2000 17.3240 ;
        RECT 14.0850 18.3415 14.1030 18.5575 ;
        RECT 15.2950 24.6775 15.3130 24.8935 ;
        RECT 15.2950 21.5095 15.3130 21.7255 ;
        RECT 15.2950 18.3415 15.3130 18.5575 ;
        RECT 15.3470 24.6775 15.3650 24.8935 ;
        RECT 15.3470 21.5095 15.3650 21.7255 ;
        RECT 15.3470 18.3415 15.3650 18.5575 ;
        RECT 15.3990 24.6775 15.4170 24.8935 ;
        RECT 15.3990 21.5095 15.4170 21.7255 ;
        RECT 15.3990 18.3415 15.4170 18.5575 ;
        RECT 15.4510 24.6775 15.4690 24.8935 ;
        RECT 15.4510 21.5095 15.4690 21.7255 ;
        RECT 15.4510 18.3415 15.4690 18.5575 ;
        RECT 15.5030 24.6775 15.5210 24.8935 ;
        RECT 15.5030 21.5095 15.5210 21.7255 ;
        RECT 15.5030 18.3415 15.5210 18.5575 ;
        RECT 16.2450 18.3415 16.2630 18.5575 ;
        RECT 0.1580 26.4830 0.1760 26.5310 ;
        RECT 14.0900 26.4830 14.1080 26.5310 ;
        RECT 15.2600 26.4830 15.2870 26.5310 ;
        RECT 15.4850 26.4830 15.5210 26.5310 ;
        RECT 16.2500 26.4830 16.2680 26.5310 ;
        RECT 30.1820 26.4830 30.2000 26.5310 ;
        RECT 0.1580 27.5630 0.1760 27.6110 ;
        RECT 14.0900 27.5630 14.1080 27.6110 ;
        RECT 15.2600 27.5630 15.2870 27.6110 ;
        RECT 15.4850 27.5630 15.5210 27.6110 ;
        RECT 16.2500 27.5630 16.2680 27.6110 ;
        RECT 30.1820 27.5630 30.2000 27.6110 ;
        RECT 0.1580 28.6430 0.1760 28.6910 ;
        RECT 14.0900 28.6430 14.1080 28.6910 ;
        RECT 15.2600 28.6430 15.2870 28.6910 ;
        RECT 15.4850 28.6430 15.5210 28.6910 ;
        RECT 16.2500 28.6430 16.2680 28.6910 ;
        RECT 30.1820 28.6430 30.2000 28.6910 ;
        RECT 0.1580 29.7230 0.1760 29.7710 ;
        RECT 14.0900 29.7230 14.1080 29.7710 ;
        RECT 15.2600 29.7230 15.2870 29.7710 ;
        RECT 15.4850 29.7230 15.5210 29.7710 ;
        RECT 16.2500 29.7230 16.2680 29.7710 ;
        RECT 30.1820 29.7230 30.2000 29.7710 ;
        RECT 0.1580 30.8030 0.1760 30.8510 ;
        RECT 14.0900 30.8030 14.1080 30.8510 ;
        RECT 15.2600 30.8030 15.2870 30.8510 ;
        RECT 15.4850 30.8030 15.5210 30.8510 ;
        RECT 16.2500 30.8030 16.2680 30.8510 ;
        RECT 30.1820 30.8030 30.2000 30.8510 ;
        RECT 0.1580 31.8830 0.1760 31.9310 ;
        RECT 14.0900 31.8830 14.1080 31.9310 ;
        RECT 15.2600 31.8830 15.2870 31.9310 ;
        RECT 15.4850 31.8830 15.5210 31.9310 ;
        RECT 16.2500 31.8830 16.2680 31.9310 ;
        RECT 30.1820 31.8830 30.2000 31.9310 ;
        RECT 0.1580 32.9630 0.1760 33.0110 ;
        RECT 14.0900 32.9630 14.1080 33.0110 ;
        RECT 15.2600 32.9630 15.2870 33.0110 ;
        RECT 15.4850 32.9630 15.5210 33.0110 ;
        RECT 16.2500 32.9630 16.2680 33.0110 ;
        RECT 30.1820 32.9630 30.2000 33.0110 ;
        RECT 0.1580 34.0430 0.1760 34.0910 ;
        RECT 14.0900 34.0430 14.1080 34.0910 ;
        RECT 15.2600 34.0430 15.2870 34.0910 ;
        RECT 15.4850 34.0430 15.5210 34.0910 ;
        RECT 16.2500 34.0430 16.2680 34.0910 ;
        RECT 30.1820 34.0430 30.2000 34.0910 ;
        RECT 0.1580 35.1230 0.1760 35.1710 ;
        RECT 14.0900 35.1230 14.1080 35.1710 ;
        RECT 15.2600 35.1230 15.2870 35.1710 ;
        RECT 15.4850 35.1230 15.5210 35.1710 ;
        RECT 16.2500 35.1230 16.2680 35.1710 ;
        RECT 30.1820 35.1230 30.2000 35.1710 ;
        RECT 0.1580 36.2030 0.1760 36.2510 ;
        RECT 14.0900 36.2030 14.1080 36.2510 ;
        RECT 15.2600 36.2030 15.2870 36.2510 ;
        RECT 15.4850 36.2030 15.5210 36.2510 ;
        RECT 16.2500 36.2030 16.2680 36.2510 ;
        RECT 30.1820 36.2030 30.2000 36.2510 ;
        RECT 0.1580 37.2830 0.1760 37.3310 ;
        RECT 14.0900 37.2830 14.1080 37.3310 ;
        RECT 15.2600 37.2830 15.2870 37.3310 ;
        RECT 15.4850 37.2830 15.5210 37.3310 ;
        RECT 16.2500 37.2830 16.2680 37.3310 ;
        RECT 30.1820 37.2830 30.2000 37.3310 ;
        RECT 0.1580 38.3630 0.1760 38.4110 ;
        RECT 14.0900 38.3630 14.1080 38.4110 ;
        RECT 15.2600 38.3630 15.2870 38.4110 ;
        RECT 15.4850 38.3630 15.5210 38.4110 ;
        RECT 16.2500 38.3630 16.2680 38.4110 ;
        RECT 30.1820 38.3630 30.2000 38.4110 ;
        RECT 0.1580 39.4430 0.1760 39.4910 ;
        RECT 14.0900 39.4430 14.1080 39.4910 ;
        RECT 15.2600 39.4430 15.2870 39.4910 ;
        RECT 15.4850 39.4430 15.5210 39.4910 ;
        RECT 16.2500 39.4430 16.2680 39.4910 ;
        RECT 30.1820 39.4430 30.2000 39.4910 ;
        RECT 0.1580 40.5230 0.1760 40.5710 ;
        RECT 14.0900 40.5230 14.1080 40.5710 ;
        RECT 15.2600 40.5230 15.2870 40.5710 ;
        RECT 15.4850 40.5230 15.5210 40.5710 ;
        RECT 16.2500 40.5230 16.2680 40.5710 ;
        RECT 30.1820 40.5230 30.2000 40.5710 ;
        RECT 0.1580 41.6030 0.1760 41.6510 ;
        RECT 14.0900 41.6030 14.1080 41.6510 ;
        RECT 15.2600 41.6030 15.2870 41.6510 ;
        RECT 15.4850 41.6030 15.5210 41.6510 ;
        RECT 16.2500 41.6030 16.2680 41.6510 ;
        RECT 30.1820 41.6030 30.2000 41.6510 ;
        RECT 0.1580 42.6830 0.1760 42.7310 ;
        RECT 14.0900 42.6830 14.1080 42.7310 ;
        RECT 15.2600 42.6830 15.2870 42.7310 ;
        RECT 15.4850 42.6830 15.5210 42.7310 ;
        RECT 16.2500 42.6830 16.2680 42.7310 ;
        RECT 30.1820 42.6830 30.2000 42.7310 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.7030 18.8135 17.7210 18.8505 ;
      LAYER M4  ;
        RECT 17.6510 18.8215 17.7350 18.8455 ;
      LAYER M5  ;
        RECT 17.7000 17.8705 17.7240 21.1105 ;
      LAYER V3  ;
        RECT 17.7030 18.8215 17.7210 18.8455 ;
      LAYER V4  ;
        RECT 17.7000 18.8215 17.7240 18.8455 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.4870 18.8165 17.5050 18.8535 ;
      LAYER M4  ;
        RECT 17.4350 18.8215 17.5190 18.8455 ;
      LAYER M5  ;
        RECT 17.4840 17.8705 17.5080 21.1105 ;
      LAYER V3  ;
        RECT 17.4870 18.8215 17.5050 18.8455 ;
      LAYER V4  ;
        RECT 17.4840 18.8215 17.5080 18.8455 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.2710 18.2375 17.2890 18.2745 ;
      LAYER M4  ;
        RECT 17.2190 18.2455 17.3030 18.2695 ;
      LAYER M5  ;
        RECT 17.2680 17.8705 17.2920 21.1105 ;
      LAYER V3  ;
        RECT 17.2710 18.2455 17.2890 18.2695 ;
      LAYER V4  ;
        RECT 17.2680 18.2455 17.2920 18.2695 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.0550 18.4775 17.0730 18.6585 ;
      LAYER M4  ;
        RECT 17.0030 18.6295 17.0870 18.6535 ;
      LAYER M5  ;
        RECT 17.0520 17.8705 17.0760 21.1105 ;
      LAYER V3  ;
        RECT 17.0550 18.6295 17.0730 18.6535 ;
      LAYER V4  ;
        RECT 17.0520 18.6295 17.0760 18.6535 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.8390 18.2405 16.8570 18.3075 ;
      LAYER M4  ;
        RECT 16.7870 18.2455 16.8710 18.2695 ;
      LAYER M5  ;
        RECT 16.8360 17.8705 16.8600 21.1105 ;
      LAYER V3  ;
        RECT 16.8390 18.2455 16.8570 18.2695 ;
      LAYER V4  ;
        RECT 16.8360 18.2455 16.8600 18.2695 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.6230 17.9735 16.6410 18.2265 ;
      LAYER M4  ;
        RECT 16.5710 18.1975 16.6550 18.2215 ;
      LAYER M5  ;
        RECT 16.6200 17.8705 16.6440 21.1105 ;
      LAYER V3  ;
        RECT 16.6230 18.1975 16.6410 18.2215 ;
      LAYER V4  ;
        RECT 16.6200 18.1975 16.6440 18.2215 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.4070 19.0085 16.4250 19.0455 ;
      LAYER M4  ;
        RECT 16.3550 19.0135 16.4390 19.0375 ;
      LAYER M5  ;
        RECT 16.4040 17.8705 16.4280 21.1105 ;
      LAYER V3  ;
        RECT 16.4070 19.0135 16.4250 19.0375 ;
      LAYER V4  ;
        RECT 16.4040 19.0135 16.4280 19.0375 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.1910 18.8555 16.2090 18.9465 ;
      LAYER M4  ;
        RECT 16.1390 18.9175 16.2230 18.9415 ;
      LAYER M5  ;
        RECT 16.1880 17.8705 16.2120 21.1105 ;
      LAYER V3  ;
        RECT 16.1910 18.9175 16.2090 18.9415 ;
      LAYER V4  ;
        RECT 16.1880 18.9175 16.2120 18.9415 ;
    END
  END ADDRESS[7]
  PIN ADDRESS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.8310 18.5135 15.8490 18.6585 ;
      LAYER M4  ;
        RECT 15.8200 18.6295 16.0070 18.6535 ;
      LAYER M5  ;
        RECT 15.9720 17.6115 15.9960 21.1105 ;
      LAYER V3  ;
        RECT 15.8310 18.6295 15.8490 18.6535 ;
      LAYER V4  ;
        RECT 15.9720 18.6295 15.9960 18.6535 ;
    END
  END ADDRESS[8]
  PIN ADDRESS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.5430 18.2405 15.5610 18.3075 ;
      LAYER M4  ;
        RECT 15.2590 18.2455 15.5720 18.2695 ;
      LAYER M5  ;
        RECT 15.2700 17.8705 15.2940 21.1105 ;
      LAYER V3  ;
        RECT 15.5430 18.2455 15.5610 18.2695 ;
      LAYER V4  ;
        RECT 15.2700 18.2455 15.2940 18.2695 ;
    END
  END ADDRESS[9]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.1470 17.9735 15.1650 18.2265 ;
      LAYER M4  ;
        RECT 14.9350 18.1975 15.1760 18.2215 ;
      LAYER M5  ;
        RECT 14.9460 17.8705 14.9700 21.1105 ;
      LAYER V3  ;
        RECT 15.1470 18.1975 15.1650 18.2215 ;
      LAYER V4  ;
        RECT 14.9460 18.1975 14.9700 18.2215 ;
    END
  END banksel
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.1390 19.1045 14.1570 19.1535 ;
      LAYER M4  ;
        RECT 14.0870 19.1095 14.1710 19.1335 ;
      LAYER M5  ;
        RECT 14.1360 17.8705 14.1600 21.1105 ;
      LAYER V3  ;
        RECT 14.1390 19.1095 14.1570 19.1335 ;
      LAYER V4  ;
        RECT 14.1360 19.1095 14.1600 19.1335 ;
    END
  END clk
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.3550 18.2405 14.3730 18.3075 ;
      LAYER M4  ;
        RECT 14.3030 18.2455 14.3870 18.2695 ;
      LAYER M5  ;
        RECT 14.3520 17.8705 14.3760 21.1105 ;
      LAYER V3  ;
        RECT 14.3550 18.2455 14.3730 18.2695 ;
      LAYER V4  ;
        RECT 14.3520 18.2455 14.3760 18.2695 ;
    END
  END write
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.1750 17.9735 14.1930 18.2265 ;
      LAYER M4  ;
        RECT 13.9090 18.1975 14.2040 18.2215 ;
      LAYER M5  ;
        RECT 13.9200 17.8705 13.9440 21.1105 ;
      LAYER V3  ;
        RECT 14.1750 18.1975 14.1930 18.2215 ;
      LAYER V4  ;
        RECT 13.9200 18.1975 13.9440 18.2215 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.7070 18.8135 13.7250 18.8505 ;
      LAYER M4  ;
        RECT 13.6550 18.8215 13.7390 18.8455 ;
      LAYER M5  ;
        RECT 13.7040 17.8705 13.7280 21.1105 ;
      LAYER V3  ;
        RECT 13.7070 18.8215 13.7250 18.8455 ;
      LAYER V4  ;
        RECT 13.7040 18.8215 13.7280 18.8455 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.4910 18.2405 13.5090 18.4695 ;
      LAYER M4  ;
        RECT 13.4390 18.2455 13.5230 18.2695 ;
      LAYER M5  ;
        RECT 13.4880 17.8705 13.5120 21.1105 ;
      LAYER V3  ;
        RECT 13.4910 18.2455 13.5090 18.2695 ;
      LAYER V4  ;
        RECT 13.4880 18.2455 13.5120 18.2695 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.2750 17.9735 13.2930 18.2265 ;
      LAYER M4  ;
        RECT 13.2230 18.1975 13.3070 18.2215 ;
      LAYER M5  ;
        RECT 13.2720 17.8705 13.2960 21.1105 ;
      LAYER V3  ;
        RECT 13.2750 18.1975 13.2930 18.2215 ;
      LAYER V4  ;
        RECT 13.2720 18.1975 13.2960 18.2215 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.0590 18.2375 13.0770 18.2745 ;
      LAYER M4  ;
        RECT 13.0070 18.2455 13.0910 18.2695 ;
      LAYER M5  ;
        RECT 13.0560 17.8705 13.0800 21.1105 ;
      LAYER V3  ;
        RECT 13.0590 18.2455 13.0770 18.2695 ;
      LAYER V4  ;
        RECT 13.0560 18.2455 13.0800 18.2695 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 12.8430 18.8135 12.8610 18.8505 ;
      LAYER M4  ;
        RECT 12.7910 18.8215 12.8750 18.8455 ;
      LAYER M5  ;
        RECT 12.8400 17.8705 12.8640 21.1105 ;
      LAYER V3  ;
        RECT 12.8430 18.8215 12.8610 18.8455 ;
      LAYER V4  ;
        RECT 12.8400 18.8215 12.8640 18.8455 ;
    END
  END sdel[4]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 15.4975 15.4670 15.7370 ;
      LAYER M4  ;
        RECT 14.8610 15.5480 15.5090 15.5720 ;
      LAYER V3  ;
        RECT 15.4490 15.5480 15.4670 15.5720 ;
    END
  END dataout[14]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 14.4175 15.4670 14.6570 ;
      LAYER M4  ;
        RECT 14.8610 14.4680 15.5090 14.4920 ;
      LAYER V3  ;
        RECT 15.4490 14.4680 15.4670 14.4920 ;
    END
  END dataout[13]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 13.3375 15.4670 13.5770 ;
      LAYER M4  ;
        RECT 14.8610 13.3880 15.5090 13.4120 ;
      LAYER V3  ;
        RECT 15.4490 13.3880 15.4670 13.4120 ;
    END
  END dataout[12]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 12.2575 15.4670 12.4970 ;
      LAYER M4  ;
        RECT 14.8610 12.3080 15.5090 12.3320 ;
      LAYER V3  ;
        RECT 15.4490 12.3080 15.4670 12.3320 ;
    END
  END dataout[11]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 11.1775 15.4670 11.4170 ;
      LAYER M4  ;
        RECT 14.8610 11.2280 15.5090 11.2520 ;
      LAYER V3  ;
        RECT 15.4490 11.2280 15.4670 11.2520 ;
    END
  END dataout[10]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 0.3775 15.4670 0.6170 ;
      LAYER M4  ;
        RECT 14.8610 0.4280 15.5090 0.4520 ;
      LAYER V3  ;
        RECT 15.4490 0.4280 15.4670 0.4520 ;
    END
  END dataout[0]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 16.5775 15.4670 16.8170 ;
      LAYER M4  ;
        RECT 14.8610 16.6280 15.5090 16.6520 ;
      LAYER V3  ;
        RECT 15.4490 16.6280 15.4670 16.6520 ;
    END
  END dataout[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 25.7845 15.4670 26.0240 ;
      LAYER M4  ;
        RECT 14.8610 25.8350 15.5090 25.8590 ;
      LAYER V3  ;
        RECT 15.4490 25.8350 15.4670 25.8590 ;
    END
  END dataout[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 26.8645 15.4670 27.1040 ;
      LAYER M4  ;
        RECT 14.8610 26.9150 15.5090 26.9390 ;
      LAYER V3  ;
        RECT 15.4490 26.9150 15.4670 26.9390 ;
    END
  END dataout[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 27.9445 15.4670 28.1840 ;
      LAYER M4  ;
        RECT 14.8610 27.9950 15.5090 28.0190 ;
      LAYER V3  ;
        RECT 15.4490 27.9950 15.4670 28.0190 ;
    END
  END dataout[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 29.0245 15.4670 29.2640 ;
      LAYER M4  ;
        RECT 14.8610 29.0750 15.5090 29.0990 ;
      LAYER V3  ;
        RECT 15.4490 29.0750 15.4670 29.0990 ;
    END
  END dataout[19]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 1.4575 15.4670 1.6970 ;
      LAYER M4  ;
        RECT 14.8610 1.5080 15.5090 1.5320 ;
      LAYER V3  ;
        RECT 15.4490 1.5080 15.4670 1.5320 ;
    END
  END dataout[1]
  PIN dataout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 30.1045 15.4670 30.3440 ;
      LAYER M4  ;
        RECT 14.8610 30.1550 15.5090 30.1790 ;
      LAYER V3  ;
        RECT 15.4490 30.1550 15.4670 30.1790 ;
    END
  END dataout[20]
  PIN dataout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 31.1845 15.4670 31.4240 ;
      LAYER M4  ;
        RECT 14.8610 31.2350 15.5090 31.2590 ;
      LAYER V3  ;
        RECT 15.4490 31.2350 15.4670 31.2590 ;
    END
  END dataout[21]
  PIN dataout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 32.2645 15.4670 32.5040 ;
      LAYER M4  ;
        RECT 14.8610 32.3150 15.5090 32.3390 ;
      LAYER V3  ;
        RECT 15.4490 32.3150 15.4670 32.3390 ;
    END
  END dataout[22]
  PIN dataout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 33.3445 15.4670 33.5840 ;
      LAYER M4  ;
        RECT 14.8610 33.3950 15.5090 33.4190 ;
      LAYER V3  ;
        RECT 15.4490 33.3950 15.4670 33.4190 ;
    END
  END dataout[23]
  PIN dataout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 34.4245 15.4670 34.6640 ;
      LAYER M4  ;
        RECT 14.8610 34.4750 15.5090 34.4990 ;
      LAYER V3  ;
        RECT 15.4490 34.4750 15.4670 34.4990 ;
    END
  END dataout[24]
  PIN dataout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 35.5045 15.4670 35.7440 ;
      LAYER M4  ;
        RECT 14.8610 35.5550 15.5090 35.5790 ;
      LAYER V3  ;
        RECT 15.4490 35.5550 15.4670 35.5790 ;
    END
  END dataout[25]
  PIN dataout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 36.5845 15.4670 36.8240 ;
      LAYER M4  ;
        RECT 14.8610 36.6350 15.5090 36.6590 ;
      LAYER V3  ;
        RECT 15.4490 36.6350 15.4670 36.6590 ;
    END
  END dataout[26]
  PIN dataout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 37.6645 15.4670 37.9040 ;
      LAYER M4  ;
        RECT 14.8610 37.7150 15.5090 37.7390 ;
      LAYER V3  ;
        RECT 15.4490 37.7150 15.4670 37.7390 ;
    END
  END dataout[27]
  PIN dataout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 38.7445 15.4670 38.9840 ;
      LAYER M4  ;
        RECT 14.8610 38.7950 15.5090 38.8190 ;
      LAYER V3  ;
        RECT 15.4490 38.7950 15.4670 38.8190 ;
    END
  END dataout[28]
  PIN dataout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 39.8245 15.4670 40.0640 ;
      LAYER M4  ;
        RECT 14.8610 39.8750 15.5090 39.8990 ;
      LAYER V3  ;
        RECT 15.4490 39.8750 15.4670 39.8990 ;
    END
  END dataout[29]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 2.5375 15.4670 2.7770 ;
      LAYER M4  ;
        RECT 14.8610 2.5880 15.5090 2.6120 ;
      LAYER V3  ;
        RECT 15.4490 2.5880 15.4670 2.6120 ;
    END
  END dataout[2]
  PIN dataout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 40.9045 15.4670 41.1440 ;
      LAYER M4  ;
        RECT 14.8610 40.9550 15.5090 40.9790 ;
      LAYER V3  ;
        RECT 15.4490 40.9550 15.4670 40.9790 ;
    END
  END dataout[30]
  PIN dataout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 41.9845 15.4670 42.2240 ;
      LAYER M4  ;
        RECT 14.8610 42.0350 15.5090 42.0590 ;
      LAYER V3  ;
        RECT 15.4490 42.0350 15.4670 42.0590 ;
    END
  END dataout[31]
  PIN dataout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[32]
  PIN dataout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[33]
  PIN dataout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[34]
  PIN dataout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[35]
  PIN dataout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[36]
  PIN dataout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[37]
  PIN dataout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[38]
  PIN dataout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[39]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 3.6175 15.4670 3.8570 ;
      LAYER M4  ;
        RECT 14.8610 3.6680 15.5090 3.6920 ;
      LAYER V3  ;
        RECT 15.4490 3.6680 15.4670 3.6920 ;
    END
  END dataout[3]
  PIN dataout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[40]
  PIN dataout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[41]
  PIN dataout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[42]
  PIN dataout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[43]
  PIN dataout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[44]
  PIN dataout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[45]
  PIN dataout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[46]
  PIN dataout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[47]
  PIN dataout[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[48]
  PIN dataout[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[49]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 4.6975 15.4670 4.9370 ;
      LAYER M4  ;
        RECT 14.8610 4.7480 15.5090 4.7720 ;
      LAYER V3  ;
        RECT 15.4490 4.7480 15.4670 4.7720 ;
    END
  END dataout[4]
  PIN dataout[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[50]
  PIN dataout[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[51]
  PIN dataout[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[52]
  PIN dataout[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[53]
  PIN dataout[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[54]
  PIN dataout[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[55]
  PIN dataout[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[56]
  PIN dataout[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[57]
  PIN dataout[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[58]
  PIN dataout[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[59]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 5.7775 15.4670 6.0170 ;
      LAYER M4  ;
        RECT 14.8610 5.8280 15.5090 5.8520 ;
      LAYER V3  ;
        RECT 15.4490 5.8280 15.4670 5.8520 ;
    END
  END dataout[5]
  PIN dataout[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[60]
  PIN dataout[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[61]
  PIN dataout[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[62]
  PIN dataout[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[63]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 6.8575 15.4670 7.0970 ;
      LAYER M4  ;
        RECT 14.8610 6.9080 15.5090 6.9320 ;
      LAYER V3  ;
        RECT 15.4490 6.9080 15.4670 6.9320 ;
    END
  END dataout[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 7.9375 15.4670 8.1770 ;
      LAYER M4  ;
        RECT 14.8610 7.9880 15.5090 8.0120 ;
      LAYER V3  ;
        RECT 15.4490 7.9880 15.4670 8.0120 ;
    END
  END dataout[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 9.0175 15.4670 9.2570 ;
      LAYER M4  ;
        RECT 14.8610 9.0680 15.5090 9.0920 ;
      LAYER V3  ;
        RECT 15.4490 9.0680 15.4670 9.0920 ;
    END
  END dataout[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 10.0975 15.4670 10.3370 ;
      LAYER M4  ;
        RECT 14.8610 10.1480 15.5090 10.1720 ;
      LAYER V3  ;
        RECT 15.4490 10.1480 15.4670 10.1720 ;
    END
  END dataout[9]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 0.2700 15.2420 0.6750 ;
      LAYER M4  ;
        RECT 14.8610 0.3320 15.4970 0.3560 ;
      LAYER V3  ;
        RECT 15.2240 0.3320 15.2420 0.3560 ;
    END
  END wd[0]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 11.0700 15.2420 11.4750 ;
      LAYER M4  ;
        RECT 14.8610 11.1320 15.4970 11.1560 ;
      LAYER V3  ;
        RECT 15.2240 11.1320 15.2420 11.1560 ;
    END
  END wd[10]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 12.1500 15.2420 12.5550 ;
      LAYER M4  ;
        RECT 14.8610 12.2120 15.4970 12.2360 ;
      LAYER V3  ;
        RECT 15.2240 12.2120 15.2420 12.2360 ;
    END
  END wd[11]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 13.2300 15.2420 13.6350 ;
      LAYER M4  ;
        RECT 14.8610 13.2920 15.4970 13.3160 ;
      LAYER V3  ;
        RECT 15.2240 13.2920 15.2420 13.3160 ;
    END
  END wd[12]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 14.3100 15.2420 14.7150 ;
      LAYER M4  ;
        RECT 14.8610 14.3720 15.4970 14.3960 ;
      LAYER V3  ;
        RECT 15.2240 14.3720 15.2420 14.3960 ;
    END
  END wd[13]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 15.3900 15.2420 15.7950 ;
      LAYER M4  ;
        RECT 14.8610 15.4520 15.4970 15.4760 ;
      LAYER V3  ;
        RECT 15.2240 15.4520 15.2420 15.4760 ;
    END
  END wd[14]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 16.4700 15.2420 16.8750 ;
      LAYER M4  ;
        RECT 14.8610 16.5320 15.4970 16.5560 ;
      LAYER V3  ;
        RECT 15.2240 16.5320 15.2420 16.5560 ;
    END
  END wd[15]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 25.6770 15.2420 26.0820 ;
      LAYER M4  ;
        RECT 14.8610 25.7390 15.4970 25.7630 ;
      LAYER V3  ;
        RECT 15.2240 25.7390 15.2420 25.7630 ;
    END
  END wd[16]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 26.7570 15.2420 27.1620 ;
      LAYER M4  ;
        RECT 14.8610 26.8190 15.4970 26.8430 ;
      LAYER V3  ;
        RECT 15.2240 26.8190 15.2420 26.8430 ;
    END
  END wd[17]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 27.8370 15.2420 28.2420 ;
      LAYER M4  ;
        RECT 14.8610 27.8990 15.4970 27.9230 ;
      LAYER V3  ;
        RECT 15.2240 27.8990 15.2420 27.9230 ;
    END
  END wd[18]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 28.9170 15.2420 29.3220 ;
      LAYER M4  ;
        RECT 14.8610 28.9790 15.4970 29.0030 ;
      LAYER V3  ;
        RECT 15.2240 28.9790 15.2420 29.0030 ;
    END
  END wd[19]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 1.3500 15.2420 1.7550 ;
      LAYER M4  ;
        RECT 14.8610 1.4120 15.4970 1.4360 ;
      LAYER V3  ;
        RECT 15.2240 1.4120 15.2420 1.4360 ;
    END
  END wd[1]
  PIN wd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 29.9970 15.2420 30.4020 ;
      LAYER M4  ;
        RECT 14.8610 30.0590 15.4970 30.0830 ;
      LAYER V3  ;
        RECT 15.2240 30.0590 15.2420 30.0830 ;
    END
  END wd[20]
  PIN wd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 31.0770 15.2420 31.4820 ;
      LAYER M4  ;
        RECT 14.8610 31.1390 15.4970 31.1630 ;
      LAYER V3  ;
        RECT 15.2240 31.1390 15.2420 31.1630 ;
    END
  END wd[21]
  PIN wd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 32.1570 15.2420 32.5620 ;
      LAYER M4  ;
        RECT 14.8610 32.2190 15.4970 32.2430 ;
      LAYER V3  ;
        RECT 15.2240 32.2190 15.2420 32.2430 ;
    END
  END wd[22]
  PIN wd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 33.2370 15.2420 33.6420 ;
      LAYER M4  ;
        RECT 14.8610 33.2990 15.4970 33.3230 ;
      LAYER V3  ;
        RECT 15.2240 33.2990 15.2420 33.3230 ;
    END
  END wd[23]
  PIN wd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 34.3170 15.2420 34.7220 ;
      LAYER M4  ;
        RECT 14.8610 34.3790 15.4970 34.4030 ;
      LAYER V3  ;
        RECT 15.2240 34.3790 15.2420 34.4030 ;
    END
  END wd[24]
  PIN wd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 35.3970 15.2420 35.8020 ;
      LAYER M4  ;
        RECT 14.8610 35.4590 15.4970 35.4830 ;
      LAYER V3  ;
        RECT 15.2240 35.4590 15.2420 35.4830 ;
    END
  END wd[25]
  PIN wd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 36.4770 15.2420 36.8820 ;
      LAYER M4  ;
        RECT 14.8610 36.5390 15.4970 36.5630 ;
      LAYER V3  ;
        RECT 15.2240 36.5390 15.2420 36.5630 ;
    END
  END wd[26]
  PIN wd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 37.5570 15.2420 37.9620 ;
      LAYER M4  ;
        RECT 14.8610 37.6190 15.4970 37.6430 ;
      LAYER V3  ;
        RECT 15.2240 37.6190 15.2420 37.6430 ;
    END
  END wd[27]
  PIN wd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 38.6370 15.2420 39.0420 ;
      LAYER M4  ;
        RECT 14.8610 38.6990 15.4970 38.7230 ;
      LAYER V3  ;
        RECT 15.2240 38.6990 15.2420 38.7230 ;
    END
  END wd[28]
  PIN wd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 39.7170 15.2420 40.1220 ;
      LAYER M4  ;
        RECT 14.8610 39.7790 15.4970 39.8030 ;
      LAYER V3  ;
        RECT 15.2240 39.7790 15.2420 39.8030 ;
    END
  END wd[29]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 2.4300 15.2420 2.8350 ;
      LAYER M4  ;
        RECT 14.8610 2.4920 15.4970 2.5160 ;
      LAYER V3  ;
        RECT 15.2240 2.4920 15.2420 2.5160 ;
    END
  END wd[2]
  PIN wd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 40.7970 15.2420 41.2020 ;
      LAYER M4  ;
        RECT 14.8610 40.8590 15.4970 40.8830 ;
      LAYER V3  ;
        RECT 15.2240 40.8590 15.2420 40.8830 ;
    END
  END wd[30]
  PIN wd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 41.8770 15.2420 42.2820 ;
      LAYER M4  ;
        RECT 14.8610 41.9390 15.4970 41.9630 ;
      LAYER V3  ;
        RECT 15.2240 41.9390 15.2420 41.9630 ;
    END
  END wd[31]
  PIN wd[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[32]
  PIN wd[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[33]
  PIN wd[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[34]
  PIN wd[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[35]
  PIN wd[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[36]
  PIN wd[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[37]
  PIN wd[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[38]
  PIN wd[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[39]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 3.5100 15.2420 3.9150 ;
      LAYER M4  ;
        RECT 14.8610 3.5720 15.4970 3.5960 ;
      LAYER V3  ;
        RECT 15.2240 3.5720 15.2420 3.5960 ;
    END
  END wd[3]
  PIN wd[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[40]
  PIN wd[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[41]
  PIN wd[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[42]
  PIN wd[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[43]
  PIN wd[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[44]
  PIN wd[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[45]
  PIN wd[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[46]
  PIN wd[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[47]
  PIN wd[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[48]
  PIN wd[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[49]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 4.5900 15.2420 4.9950 ;
      LAYER M4  ;
        RECT 14.8610 4.6520 15.4970 4.6760 ;
      LAYER V3  ;
        RECT 15.2240 4.6520 15.2420 4.6760 ;
    END
  END wd[4]
  PIN wd[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[50]
  PIN wd[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[51]
  PIN wd[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[52]
  PIN wd[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[53]
  PIN wd[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[54]
  PIN wd[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[55]
  PIN wd[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[56]
  PIN wd[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[57]
  PIN wd[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[58]
  PIN wd[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[59]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 5.6700 15.2420 6.0750 ;
      LAYER M4  ;
        RECT 14.8610 5.7320 15.4970 5.7560 ;
      LAYER V3  ;
        RECT 15.2240 5.7320 15.2420 5.7560 ;
    END
  END wd[5]
  PIN wd[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[60]
  PIN wd[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[61]
  PIN wd[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[62]
  PIN wd[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[63]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 6.7500 15.2420 7.1550 ;
      LAYER M4  ;
        RECT 14.8610 6.8120 15.4970 6.8360 ;
      LAYER V3  ;
        RECT 15.2240 6.8120 15.2420 6.8360 ;
    END
  END wd[6]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 7.8300 15.2420 8.2350 ;
      LAYER M4  ;
        RECT 14.8610 7.8920 15.4970 7.9160 ;
      LAYER V3  ;
        RECT 15.2240 7.8920 15.2420 7.9160 ;
    END
  END wd[7]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 8.9100 15.2420 9.3150 ;
      LAYER M4  ;
        RECT 14.8610 8.9720 15.4970 8.9960 ;
      LAYER V3  ;
        RECT 15.2240 8.9720 15.2420 8.9960 ;
    END
  END wd[8]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 9.9900 15.2420 10.3950 ;
      LAYER M4  ;
        RECT 14.8610 10.0520 15.4970 10.0760 ;
      LAYER V3  ;
        RECT 15.2240 10.0520 15.2420 10.0760 ;
    END
  END wd[9]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0000 17.5735 30.3480 26.2270 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
        RECT 0.0050 29.9835 30.3530 31.0770 ;
        RECT 0.0050 31.0635 30.3530 32.1570 ;
        RECT 0.0050 32.1435 30.3530 33.2370 ;
        RECT 0.0050 33.2235 30.3530 34.3170 ;
        RECT 0.0050 34.3035 30.3530 35.3970 ;
        RECT 0.0050 35.3835 30.3530 36.4770 ;
        RECT 0.0050 36.4635 30.3530 37.5570 ;
        RECT 0.0050 37.5435 30.3530 38.6370 ;
        RECT 0.0050 38.6235 30.3530 39.7170 ;
        RECT 0.0050 39.7035 30.3530 40.7970 ;
        RECT 0.0050 40.7835 30.3530 41.8770 ;
        RECT 0.0050 41.8635 30.3530 42.9570 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0000 17.5735 30.3480 26.2270 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
        RECT 0.0050 29.9835 30.3530 31.0770 ;
        RECT 0.0050 31.0635 30.3530 32.1570 ;
        RECT 0.0050 32.1435 30.3530 33.2370 ;
        RECT 0.0050 33.2235 30.3530 34.3170 ;
        RECT 0.0050 34.3035 30.3530 35.3970 ;
        RECT 0.0050 35.3835 30.3530 36.4770 ;
        RECT 0.0050 36.4635 30.3530 37.5570 ;
        RECT 0.0050 37.5435 30.3530 38.6370 ;
        RECT 0.0050 38.6235 30.3530 39.7170 ;
        RECT 0.0050 39.7035 30.3530 40.7970 ;
        RECT 0.0050 40.7835 30.3530 41.8770 ;
        RECT 0.0050 41.8635 30.3530 42.9570 ;
  LAYER V1 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0000 17.5735 30.3480 26.2270 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
        RECT 0.0050 29.9835 30.3530 31.0770 ;
        RECT 0.0050 31.0635 30.3530 32.1570 ;
        RECT 0.0050 32.1435 30.3530 33.2370 ;
        RECT 0.0050 33.2235 30.3530 34.3170 ;
        RECT 0.0050 34.3035 30.3530 35.3970 ;
        RECT 0.0050 35.3835 30.3530 36.4770 ;
        RECT 0.0050 36.4635 30.3530 37.5570 ;
        RECT 0.0050 37.5435 30.3530 38.6370 ;
        RECT 0.0050 38.6235 30.3530 39.7170 ;
        RECT 0.0050 39.7035 30.3530 40.7970 ;
        RECT 0.0050 40.7835 30.3530 41.8770 ;
        RECT 0.0050 41.8635 30.3530 42.9570 ;
  LAYER V2 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0000 17.5735 30.3480 26.2270 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
        RECT 0.0050 29.9835 30.3530 31.0770 ;
        RECT 0.0050 31.0635 30.3530 32.1570 ;
        RECT 0.0050 32.1435 30.3530 33.2370 ;
        RECT 0.0050 33.2235 30.3530 34.3170 ;
        RECT 0.0050 34.3035 30.3530 35.3970 ;
        RECT 0.0050 35.3835 30.3530 36.4770 ;
        RECT 0.0050 36.4635 30.3530 37.5570 ;
        RECT 0.0050 37.5435 30.3530 38.6370 ;
        RECT 0.0050 38.6235 30.3530 39.7170 ;
        RECT 0.0050 39.7035 30.3530 40.7970 ;
        RECT 0.0050 40.7835 30.3530 41.8770 ;
        RECT 0.0050 41.8635 30.3530 42.9570 ;
  LAYER M3  ;
      RECT 15.6110 0.3450 15.6290 1.2805 ;
      RECT 15.5750 0.3450 15.5930 1.2805 ;
      RECT 15.5390 0.9220 15.5570 1.2445 ;
      RECT 15.4220 1.1190 15.4400 1.2285 ;
      RECT 15.4130 0.3775 15.4310 0.6170 ;
      RECT 15.3770 0.9585 15.3950 1.1120 ;
      RECT 15.2960 0.9840 15.3140 1.2420 ;
      RECT 14.7560 0.3450 14.7740 1.2805 ;
      RECT 14.7200 0.3450 14.7380 1.2805 ;
      RECT 14.6840 0.5260 14.7020 1.0940 ;
      RECT 15.6110 1.4250 15.6290 2.3605 ;
      RECT 15.5750 1.4250 15.5930 2.3605 ;
      RECT 15.5390 2.0020 15.5570 2.3245 ;
      RECT 15.4220 2.1990 15.4400 2.3085 ;
      RECT 15.4130 1.4575 15.4310 1.6970 ;
      RECT 15.3770 2.0385 15.3950 2.1920 ;
      RECT 15.2960 2.0640 15.3140 2.3220 ;
      RECT 14.7560 1.4250 14.7740 2.3605 ;
      RECT 14.7200 1.4250 14.7380 2.3605 ;
      RECT 14.6840 1.6060 14.7020 2.1740 ;
      RECT 15.6110 2.5050 15.6290 3.4405 ;
      RECT 15.5750 2.5050 15.5930 3.4405 ;
      RECT 15.5390 3.0820 15.5570 3.4045 ;
      RECT 15.4220 3.2790 15.4400 3.3885 ;
      RECT 15.4130 2.5375 15.4310 2.7770 ;
      RECT 15.3770 3.1185 15.3950 3.2720 ;
      RECT 15.2960 3.1440 15.3140 3.4020 ;
      RECT 14.7560 2.5050 14.7740 3.4405 ;
      RECT 14.7200 2.5050 14.7380 3.4405 ;
      RECT 14.6840 2.6860 14.7020 3.2540 ;
      RECT 15.6110 3.5850 15.6290 4.5205 ;
      RECT 15.5750 3.5850 15.5930 4.5205 ;
      RECT 15.5390 4.1620 15.5570 4.4845 ;
      RECT 15.4220 4.3590 15.4400 4.4685 ;
      RECT 15.4130 3.6175 15.4310 3.8570 ;
      RECT 15.3770 4.1985 15.3950 4.3520 ;
      RECT 15.2960 4.2240 15.3140 4.4820 ;
      RECT 14.7560 3.5850 14.7740 4.5205 ;
      RECT 14.7200 3.5850 14.7380 4.5205 ;
      RECT 14.6840 3.7660 14.7020 4.3340 ;
      RECT 15.6110 4.6650 15.6290 5.6005 ;
      RECT 15.5750 4.6650 15.5930 5.6005 ;
      RECT 15.5390 5.2420 15.5570 5.5645 ;
      RECT 15.4220 5.4390 15.4400 5.5485 ;
      RECT 15.4130 4.6975 15.4310 4.9370 ;
      RECT 15.3770 5.2785 15.3950 5.4320 ;
      RECT 15.2960 5.3040 15.3140 5.5620 ;
      RECT 14.7560 4.6650 14.7740 5.6005 ;
      RECT 14.7200 4.6650 14.7380 5.6005 ;
      RECT 14.6840 4.8460 14.7020 5.4140 ;
      RECT 15.6110 5.7450 15.6290 6.6805 ;
      RECT 15.5750 5.7450 15.5930 6.6805 ;
      RECT 15.5390 6.3220 15.5570 6.6445 ;
      RECT 15.4220 6.5190 15.4400 6.6285 ;
      RECT 15.4130 5.7775 15.4310 6.0170 ;
      RECT 15.3770 6.3585 15.3950 6.5120 ;
      RECT 15.2960 6.3840 15.3140 6.6420 ;
      RECT 14.7560 5.7450 14.7740 6.6805 ;
      RECT 14.7200 5.7450 14.7380 6.6805 ;
      RECT 14.6840 5.9260 14.7020 6.4940 ;
      RECT 15.6110 6.8250 15.6290 7.7605 ;
      RECT 15.5750 6.8250 15.5930 7.7605 ;
      RECT 15.5390 7.4020 15.5570 7.7245 ;
      RECT 15.4220 7.5990 15.4400 7.7085 ;
      RECT 15.4130 6.8575 15.4310 7.0970 ;
      RECT 15.3770 7.4385 15.3950 7.5920 ;
      RECT 15.2960 7.4640 15.3140 7.7220 ;
      RECT 14.7560 6.8250 14.7740 7.7605 ;
      RECT 14.7200 6.8250 14.7380 7.7605 ;
      RECT 14.6840 7.0060 14.7020 7.5740 ;
      RECT 15.6110 7.9050 15.6290 8.8405 ;
      RECT 15.5750 7.9050 15.5930 8.8405 ;
      RECT 15.5390 8.4820 15.5570 8.8045 ;
      RECT 15.4220 8.6790 15.4400 8.7885 ;
      RECT 15.4130 7.9375 15.4310 8.1770 ;
      RECT 15.3770 8.5185 15.3950 8.6720 ;
      RECT 15.2960 8.5440 15.3140 8.8020 ;
      RECT 14.7560 7.9050 14.7740 8.8405 ;
      RECT 14.7200 7.9050 14.7380 8.8405 ;
      RECT 14.6840 8.0860 14.7020 8.6540 ;
      RECT 15.6110 8.9850 15.6290 9.9205 ;
      RECT 15.5750 8.9850 15.5930 9.9205 ;
      RECT 15.5390 9.5620 15.5570 9.8845 ;
      RECT 15.4220 9.7590 15.4400 9.8685 ;
      RECT 15.4130 9.0175 15.4310 9.2570 ;
      RECT 15.3770 9.5985 15.3950 9.7520 ;
      RECT 15.2960 9.6240 15.3140 9.8820 ;
      RECT 14.7560 8.9850 14.7740 9.9205 ;
      RECT 14.7200 8.9850 14.7380 9.9205 ;
      RECT 14.6840 9.1660 14.7020 9.7340 ;
      RECT 15.6110 10.0650 15.6290 11.0005 ;
      RECT 15.5750 10.0650 15.5930 11.0005 ;
      RECT 15.5390 10.6420 15.5570 10.9645 ;
      RECT 15.4220 10.8390 15.4400 10.9485 ;
      RECT 15.4130 10.0975 15.4310 10.3370 ;
      RECT 15.3770 10.6785 15.3950 10.8320 ;
      RECT 15.2960 10.7040 15.3140 10.9620 ;
      RECT 14.7560 10.0650 14.7740 11.0005 ;
      RECT 14.7200 10.0650 14.7380 11.0005 ;
      RECT 14.6840 10.2460 14.7020 10.8140 ;
      RECT 15.6110 11.1450 15.6290 12.0805 ;
      RECT 15.5750 11.1450 15.5930 12.0805 ;
      RECT 15.5390 11.7220 15.5570 12.0445 ;
      RECT 15.4220 11.9190 15.4400 12.0285 ;
      RECT 15.4130 11.1775 15.4310 11.4170 ;
      RECT 15.3770 11.7585 15.3950 11.9120 ;
      RECT 15.2960 11.7840 15.3140 12.0420 ;
      RECT 14.7560 11.1450 14.7740 12.0805 ;
      RECT 14.7200 11.1450 14.7380 12.0805 ;
      RECT 14.6840 11.3260 14.7020 11.8940 ;
      RECT 15.6110 12.2250 15.6290 13.1605 ;
      RECT 15.5750 12.2250 15.5930 13.1605 ;
      RECT 15.5390 12.8020 15.5570 13.1245 ;
      RECT 15.4220 12.9990 15.4400 13.1085 ;
      RECT 15.4130 12.2575 15.4310 12.4970 ;
      RECT 15.3770 12.8385 15.3950 12.9920 ;
      RECT 15.2960 12.8640 15.3140 13.1220 ;
      RECT 14.7560 12.2250 14.7740 13.1605 ;
      RECT 14.7200 12.2250 14.7380 13.1605 ;
      RECT 14.6840 12.4060 14.7020 12.9740 ;
      RECT 15.6110 13.3050 15.6290 14.2405 ;
      RECT 15.5750 13.3050 15.5930 14.2405 ;
      RECT 15.5390 13.8820 15.5570 14.2045 ;
      RECT 15.4220 14.0790 15.4400 14.1885 ;
      RECT 15.4130 13.3375 15.4310 13.5770 ;
      RECT 15.3770 13.9185 15.3950 14.0720 ;
      RECT 15.2960 13.9440 15.3140 14.2020 ;
      RECT 14.7560 13.3050 14.7740 14.2405 ;
      RECT 14.7200 13.3050 14.7380 14.2405 ;
      RECT 14.6840 13.4860 14.7020 14.0540 ;
      RECT 15.6110 14.3850 15.6290 15.3205 ;
      RECT 15.5750 14.3850 15.5930 15.3205 ;
      RECT 15.5390 14.9620 15.5570 15.2845 ;
      RECT 15.4220 15.1590 15.4400 15.2685 ;
      RECT 15.4130 14.4175 15.4310 14.6570 ;
      RECT 15.3770 14.9985 15.3950 15.1520 ;
      RECT 15.2960 15.0240 15.3140 15.2820 ;
      RECT 14.7560 14.3850 14.7740 15.3205 ;
      RECT 14.7200 14.3850 14.7380 15.3205 ;
      RECT 14.6840 14.5660 14.7020 15.1340 ;
      RECT 15.6110 15.4650 15.6290 16.4005 ;
      RECT 15.5750 15.4650 15.5930 16.4005 ;
      RECT 15.5390 16.0420 15.5570 16.3645 ;
      RECT 15.4220 16.2390 15.4400 16.3485 ;
      RECT 15.4130 15.4975 15.4310 15.7370 ;
      RECT 15.3770 16.0785 15.3950 16.2320 ;
      RECT 15.2960 16.1040 15.3140 16.3620 ;
      RECT 14.7560 15.4650 14.7740 16.4005 ;
      RECT 14.7200 15.4650 14.7380 16.4005 ;
      RECT 14.6840 15.6460 14.7020 16.2140 ;
      RECT 15.6110 16.5450 15.6290 17.4805 ;
      RECT 15.5750 16.5450 15.5930 17.4805 ;
      RECT 15.5390 17.1220 15.5570 17.4445 ;
      RECT 15.4220 17.3190 15.4400 17.4285 ;
      RECT 15.4130 16.5775 15.4310 16.8170 ;
      RECT 15.3770 17.1585 15.3950 17.3120 ;
      RECT 15.2960 17.1840 15.3140 17.4420 ;
      RECT 14.7560 16.5450 14.7740 17.4805 ;
      RECT 14.7200 16.5450 14.7380 17.4805 ;
      RECT 14.6840 16.7260 14.7020 17.2940 ;
      RECT 30.2130 17.3835 30.2310 25.7540 ;
      RECT 30.1770 17.3835 30.1950 25.7540 ;
      RECT 30.0690 17.3835 30.0870 21.1245 ;
      RECT 29.9610 17.3835 29.9790 21.1245 ;
      RECT 29.8530 17.3835 29.8710 21.1245 ;
      RECT 29.7450 17.3835 29.7630 21.1245 ;
      RECT 29.6370 17.3835 29.6550 21.1245 ;
      RECT 29.5290 17.3835 29.5470 21.1245 ;
      RECT 29.4210 17.3835 29.4390 21.1245 ;
      RECT 29.3130 17.3835 29.3310 21.1245 ;
      RECT 29.2050 17.3835 29.2230 21.1245 ;
      RECT 29.0970 17.3835 29.1150 21.1245 ;
      RECT 28.9890 17.3835 29.0070 21.1245 ;
      RECT 28.8810 17.3835 28.8990 21.1245 ;
      RECT 28.7730 17.3835 28.7910 21.1245 ;
      RECT 28.6650 17.3835 28.6830 21.1245 ;
      RECT 28.5570 17.3835 28.5750 21.1245 ;
      RECT 28.4490 17.3835 28.4670 21.1245 ;
      RECT 28.3410 17.3835 28.3590 21.1245 ;
      RECT 28.2330 17.3835 28.2510 21.1245 ;
      RECT 28.1250 17.3835 28.1430 21.1245 ;
      RECT 28.0170 17.3835 28.0350 21.1245 ;
      RECT 27.9090 17.3835 27.9270 21.1245 ;
      RECT 27.8010 17.3835 27.8190 21.1245 ;
      RECT 27.6930 17.3835 27.7110 21.1245 ;
      RECT 27.5850 17.3835 27.6030 21.1245 ;
      RECT 27.4770 17.3835 27.4950 21.1245 ;
      RECT 27.3690 17.3835 27.3870 21.1245 ;
      RECT 27.2610 17.3835 27.2790 21.1245 ;
      RECT 27.1530 17.3835 27.1710 21.1245 ;
      RECT 27.0450 17.3835 27.0630 21.1245 ;
      RECT 26.9370 17.3835 26.9550 21.1245 ;
      RECT 26.8290 17.3835 26.8470 21.1245 ;
      RECT 26.7210 17.3835 26.7390 21.1245 ;
      RECT 26.6130 17.3835 26.6310 21.1245 ;
      RECT 26.5050 17.3835 26.5230 21.1245 ;
      RECT 26.3970 17.3835 26.4150 21.1245 ;
      RECT 26.2890 17.3835 26.3070 21.1245 ;
      RECT 26.1810 17.3835 26.1990 21.1245 ;
      RECT 26.0730 17.3835 26.0910 21.1245 ;
      RECT 25.9650 17.3835 25.9830 21.1245 ;
      RECT 25.8570 17.3835 25.8750 21.1245 ;
      RECT 25.7490 17.3835 25.7670 21.1245 ;
      RECT 25.6410 17.3835 25.6590 21.1245 ;
      RECT 25.5330 17.3835 25.5510 21.1245 ;
      RECT 25.4250 17.3835 25.4430 21.1245 ;
      RECT 25.3170 17.3835 25.3350 21.1245 ;
      RECT 25.2090 17.3835 25.2270 21.1245 ;
      RECT 25.1010 17.3835 25.1190 21.1245 ;
      RECT 24.9930 17.3835 25.0110 21.1245 ;
      RECT 24.8850 17.3835 24.9030 21.1245 ;
      RECT 24.7770 17.3835 24.7950 21.1245 ;
      RECT 24.6690 17.3835 24.6870 21.1245 ;
      RECT 24.5610 17.3835 24.5790 21.1245 ;
      RECT 24.4530 17.3835 24.4710 21.1245 ;
      RECT 24.3450 17.3835 24.3630 21.1245 ;
      RECT 24.2370 17.3835 24.2550 21.1245 ;
      RECT 24.1290 17.3835 24.1470 21.1245 ;
      RECT 24.0210 17.3835 24.0390 21.1245 ;
      RECT 23.9130 17.3835 23.9310 21.1245 ;
      RECT 23.8050 17.3835 23.8230 21.1245 ;
      RECT 23.6970 17.3835 23.7150 21.1245 ;
      RECT 23.5890 17.3835 23.6070 21.1245 ;
      RECT 23.4810 17.3835 23.4990 21.1245 ;
      RECT 23.3730 17.3835 23.3910 21.1245 ;
      RECT 23.2650 17.3835 23.2830 21.1245 ;
      RECT 23.1570 17.3835 23.1750 21.1245 ;
      RECT 23.0490 17.3835 23.0670 21.1245 ;
      RECT 22.9410 17.3835 22.9590 21.1245 ;
      RECT 22.8330 17.3835 22.8510 21.1245 ;
      RECT 22.7250 17.3835 22.7430 21.1245 ;
      RECT 22.6170 17.3835 22.6350 21.1245 ;
      RECT 22.5090 17.3835 22.5270 21.1245 ;
      RECT 22.4010 17.3835 22.4190 21.1245 ;
      RECT 22.2930 17.3835 22.3110 21.1245 ;
      RECT 22.1850 17.3835 22.2030 21.1245 ;
      RECT 22.0770 17.3835 22.0950 21.1245 ;
      RECT 21.9690 17.3835 21.9870 21.1245 ;
      RECT 21.8610 17.3835 21.8790 21.1245 ;
      RECT 21.7530 17.3835 21.7710 21.1245 ;
      RECT 21.6450 17.3835 21.6630 21.1245 ;
      RECT 21.5370 17.3835 21.5550 21.1245 ;
      RECT 21.4290 17.3835 21.4470 21.1245 ;
      RECT 21.3210 17.3835 21.3390 21.1245 ;
      RECT 21.2130 17.3835 21.2310 21.1245 ;
      RECT 21.1050 17.3835 21.1230 21.1245 ;
      RECT 20.9970 17.3835 21.0150 21.1245 ;
      RECT 20.8890 17.3835 20.9070 21.1245 ;
      RECT 20.7810 17.3835 20.7990 21.1245 ;
      RECT 20.6730 17.3835 20.6910 21.1245 ;
      RECT 20.5650 17.3835 20.5830 21.1245 ;
      RECT 20.4570 17.3835 20.4750 21.1245 ;
      RECT 20.3490 17.3835 20.3670 21.1245 ;
      RECT 20.2410 17.3835 20.2590 21.1245 ;
      RECT 20.1330 17.3835 20.1510 21.1245 ;
      RECT 20.0250 17.3835 20.0430 21.1245 ;
      RECT 19.9170 17.3835 19.9350 21.1245 ;
      RECT 19.8090 17.5470 19.8270 17.8970 ;
      RECT 19.7010 17.3835 19.7190 21.1245 ;
      RECT 19.5930 17.3835 19.6110 21.1245 ;
      RECT 19.4850 17.3835 19.5030 21.1245 ;
      RECT 19.3770 17.3835 19.3950 21.1245 ;
      RECT 19.2690 17.3835 19.2870 21.1245 ;
      RECT 19.1610 17.3835 19.1790 21.1245 ;
      RECT 19.0530 17.3835 19.0710 21.1245 ;
      RECT 18.9450 17.3835 18.9630 21.1245 ;
      RECT 18.8370 17.3835 18.8550 21.1245 ;
      RECT 18.7290 17.3835 18.7470 21.1245 ;
      RECT 18.6210 17.3835 18.6390 21.1245 ;
      RECT 18.5130 17.3835 18.5310 21.1245 ;
      RECT 18.4050 17.3835 18.4230 21.1245 ;
      RECT 18.2970 17.3835 18.3150 21.1245 ;
      RECT 18.1890 17.3835 18.2070 21.1245 ;
      RECT 18.0810 17.3835 18.0990 21.1245 ;
      RECT 17.9730 17.3835 17.9910 21.1245 ;
      RECT 17.8650 17.3835 17.8830 21.1245 ;
      RECT 17.7570 17.3835 17.7750 21.1245 ;
      RECT 17.6490 17.3835 17.6670 21.1245 ;
      RECT 17.5410 17.3835 17.5590 21.1245 ;
      RECT 17.4330 17.3835 17.4510 21.1245 ;
      RECT 17.3250 17.3835 17.3430 21.1245 ;
      RECT 17.2170 17.3835 17.2350 21.1245 ;
      RECT 17.1090 17.3835 17.1270 21.1245 ;
      RECT 17.0010 17.3835 17.0190 21.1245 ;
      RECT 16.8930 17.3835 16.9110 21.1245 ;
      RECT 16.7850 17.3835 16.8030 21.1245 ;
      RECT 16.6770 17.3835 16.6950 21.1245 ;
      RECT 16.5690 17.3835 16.5870 21.1245 ;
      RECT 16.4610 17.3835 16.4790 21.1245 ;
      RECT 16.4250 21.3355 16.4430 22.0402 ;
      RECT 16.4250 22.7785 16.4430 23.9395 ;
      RECT 16.4070 18.2075 16.4250 18.8835 ;
      RECT 16.4070 19.6295 16.4250 19.9275 ;
      RECT 16.4070 20.7455 16.4250 21.0075 ;
      RECT 16.3890 21.3990 16.4070 22.0890 ;
      RECT 16.3890 22.1400 16.4070 23.1255 ;
      RECT 16.3890 23.1665 16.4070 23.7835 ;
      RECT 16.3530 17.3835 16.3710 25.7540 ;
      RECT 16.3170 21.6715 16.3350 21.7545 ;
      RECT 16.2990 18.3155 16.3170 18.9465 ;
      RECT 16.2990 19.3595 16.3170 19.5495 ;
      RECT 16.2990 20.2415 16.3170 20.2905 ;
      RECT 16.2990 20.9735 16.3170 21.0105 ;
      RECT 16.2810 21.3665 16.2990 24.9595 ;
      RECT 16.1910 17.5800 16.2090 17.7180 ;
      RECT 16.1910 17.9375 16.2090 18.7395 ;
      RECT 16.1910 19.2875 16.2090 19.8555 ;
      RECT 16.1910 21.3665 16.2090 24.9595 ;
      RECT 16.1550 19.3595 16.1730 19.7295 ;
      RECT 16.1190 18.7115 16.1370 18.8475 ;
      RECT 16.1190 19.7015 16.1370 19.9275 ;
      RECT 16.1190 20.9435 16.1370 21.0075 ;
      RECT 16.0830 18.8135 16.1010 18.8505 ;
      RECT 16.0830 20.4395 16.1010 20.4825 ;
      RECT 16.0830 20.9735 16.1010 21.0105 ;
      RECT 16.0470 19.1255 16.0650 19.6215 ;
      RECT 16.0470 19.6655 16.0650 19.8555 ;
      RECT 16.0470 20.6255 16.0650 20.9355 ;
      RECT 16.0110 19.0175 16.0290 20.2645 ;
      RECT 15.0390 17.5735 15.0570 17.7275 ;
      RECT 15.0030 17.5735 15.0210 17.6235 ;
      RECT 14.9310 17.5735 14.9490 17.6450 ;
      RECT 14.2830 18.7115 14.3010 19.1175 ;
      RECT 14.2470 19.8215 14.2650 19.8585 ;
      RECT 14.2110 18.7475 14.2290 19.3515 ;
      RECT 14.1750 18.5855 14.1930 18.6495 ;
      RECT 14.1390 17.6265 14.1570 17.6775 ;
      RECT 14.1390 20.7455 14.1570 20.9355 ;
      RECT 14.1390 21.3665 14.1570 24.9595 ;
      RECT 14.0310 18.0455 14.0490 18.2355 ;
      RECT 14.0310 18.8195 14.0490 21.0795 ;
      RECT 14.0130 21.6715 14.0310 21.7545 ;
      RECT 13.9770 17.5470 13.9950 25.7540 ;
      RECT 13.9410 21.3990 13.9590 22.0890 ;
      RECT 13.9410 22.1400 13.9590 23.1255 ;
      RECT 13.9410 23.1665 13.9590 23.7835 ;
      RECT 13.9230 18.0455 13.9410 18.5415 ;
      RECT 13.9230 19.3235 13.9410 19.8915 ;
      RECT 13.9230 20.2055 13.9410 20.9355 ;
      RECT 13.9050 21.3355 13.9230 22.0402 ;
      RECT 13.9050 22.7785 13.9230 23.9395 ;
      RECT 13.8690 17.5470 13.8870 17.8970 ;
      RECT 13.8690 21.0910 13.8870 25.7540 ;
      RECT 13.7610 17.5470 13.7790 17.8970 ;
      RECT 13.6530 17.5470 13.6710 17.8970 ;
      RECT 13.5450 17.5470 13.5630 17.8970 ;
      RECT 13.4370 17.5470 13.4550 17.8970 ;
      RECT 13.3290 17.5470 13.3470 17.8970 ;
      RECT 13.2210 17.5470 13.2390 17.8970 ;
      RECT 13.1130 17.5470 13.1310 17.8970 ;
      RECT 13.0050 17.5470 13.0230 17.8970 ;
      RECT 12.8970 17.5470 12.9150 17.8970 ;
      RECT 12.7890 17.5470 12.8070 17.8970 ;
      RECT 12.6810 17.5470 12.6990 17.8970 ;
      RECT 12.5730 17.5470 12.5910 17.8970 ;
      RECT 12.4650 17.5470 12.4830 17.8970 ;
      RECT 12.3570 17.5470 12.3750 17.8970 ;
      RECT 12.2490 17.5470 12.2670 17.8970 ;
      RECT 12.1410 17.5470 12.1590 17.8970 ;
      RECT 12.0330 17.5470 12.0510 17.8970 ;
      RECT 11.9250 17.5470 11.9430 17.8970 ;
      RECT 11.8170 17.5470 11.8350 17.8970 ;
      RECT 11.7090 17.5470 11.7270 17.8970 ;
      RECT 11.6010 17.5470 11.6190 17.8970 ;
      RECT 11.4930 17.5470 11.5110 17.8970 ;
      RECT 11.3850 17.5470 11.4030 17.8970 ;
      RECT 11.2770 17.5470 11.2950 17.8970 ;
      RECT 11.1690 17.5470 11.1870 17.8970 ;
      RECT 11.0610 17.5470 11.0790 17.8970 ;
      RECT 10.9530 17.5470 10.9710 17.8970 ;
      RECT 10.8450 17.5470 10.8630 17.8970 ;
      RECT 10.7370 17.5470 10.7550 17.8970 ;
      RECT 10.6290 17.5470 10.6470 17.8970 ;
      RECT 10.5210 17.5470 10.5390 17.8970 ;
      RECT 10.4130 17.5470 10.4310 17.8970 ;
      RECT 10.3050 17.5470 10.3230 17.8970 ;
      RECT 10.1970 17.5470 10.2150 17.8970 ;
      RECT 10.0890 17.5470 10.1070 17.8970 ;
      RECT 9.9810 17.5470 9.9990 17.8970 ;
      RECT 9.8730 17.5470 9.8910 17.8970 ;
      RECT 9.7650 17.5470 9.7830 17.8970 ;
      RECT 9.6570 17.5470 9.6750 17.8970 ;
      RECT 9.5490 17.5470 9.5670 17.8970 ;
      RECT 9.4410 17.5470 9.4590 17.8970 ;
      RECT 9.3330 17.5470 9.3510 17.8970 ;
      RECT 9.2250 17.5470 9.2430 17.8970 ;
      RECT 9.1170 17.5470 9.1350 17.8970 ;
      RECT 9.0090 17.5470 9.0270 17.8970 ;
      RECT 8.9010 17.5470 8.9190 17.8970 ;
      RECT 8.7930 17.5470 8.8110 17.8970 ;
      RECT 8.6850 17.5470 8.7030 17.8970 ;
      RECT 8.5770 17.5470 8.5950 17.8970 ;
      RECT 8.4690 17.5470 8.4870 17.8970 ;
      RECT 8.3610 17.5470 8.3790 17.8970 ;
      RECT 8.2530 17.5470 8.2710 17.8970 ;
      RECT 8.1450 17.5470 8.1630 17.8970 ;
      RECT 8.0370 17.5470 8.0550 17.8970 ;
      RECT 7.9290 17.5470 7.9470 17.8970 ;
      RECT 7.8210 17.5470 7.8390 17.8970 ;
      RECT 7.7130 17.5470 7.7310 17.8970 ;
      RECT 7.6050 17.5470 7.6230 17.8970 ;
      RECT 7.4970 17.5470 7.5150 17.8970 ;
      RECT 7.3890 17.5470 7.4070 17.8970 ;
      RECT 7.2810 17.5470 7.2990 17.8970 ;
      RECT 7.1730 17.5470 7.1910 17.8970 ;
      RECT 7.0650 17.5470 7.0830 17.8970 ;
      RECT 6.9570 17.5470 6.9750 17.8970 ;
      RECT 6.8490 17.5470 6.8670 17.8970 ;
      RECT 6.7410 17.5470 6.7590 17.8970 ;
      RECT 6.6330 17.5470 6.6510 17.8970 ;
      RECT 6.5250 17.5470 6.5430 17.8970 ;
      RECT 6.4170 17.5470 6.4350 17.8970 ;
      RECT 6.3090 17.5470 6.3270 17.8970 ;
      RECT 6.2010 17.5470 6.2190 17.8970 ;
      RECT 6.0930 17.5470 6.1110 17.8970 ;
      RECT 5.9850 17.5470 6.0030 17.8970 ;
      RECT 5.8770 17.5470 5.8950 17.8970 ;
      RECT 5.7690 17.5470 5.7870 17.8970 ;
      RECT 5.6610 17.5470 5.6790 17.8970 ;
      RECT 5.5530 17.5470 5.5710 17.8970 ;
      RECT 5.4450 17.5470 5.4630 17.8970 ;
      RECT 5.3370 17.5470 5.3550 17.8970 ;
      RECT 5.2290 17.5470 5.2470 17.8970 ;
      RECT 5.1210 17.5470 5.1390 17.8970 ;
      RECT 5.0130 17.5470 5.0310 17.8970 ;
      RECT 4.9050 17.5470 4.9230 17.8970 ;
      RECT 4.7970 17.5470 4.8150 17.8970 ;
      RECT 4.6890 17.5470 4.7070 17.8970 ;
      RECT 4.5810 17.5470 4.5990 17.8970 ;
      RECT 4.4730 17.5470 4.4910 17.8970 ;
      RECT 4.3650 17.5470 4.3830 17.8970 ;
      RECT 4.2570 17.5470 4.2750 17.8970 ;
      RECT 4.1490 17.5470 4.1670 17.8970 ;
      RECT 4.0410 17.5470 4.0590 17.8970 ;
      RECT 3.9330 17.5470 3.9510 17.8970 ;
      RECT 3.8250 17.5470 3.8430 17.8970 ;
      RECT 3.7170 17.5470 3.7350 17.8970 ;
      RECT 3.6090 17.5470 3.6270 17.8970 ;
      RECT 3.5010 17.5470 3.5190 17.8970 ;
      RECT 3.3930 17.5470 3.4110 17.8970 ;
      RECT 3.2850 17.5470 3.3030 17.8970 ;
      RECT 3.1770 17.5470 3.1950 17.8970 ;
      RECT 3.0690 17.5470 3.0870 17.8970 ;
      RECT 2.9610 17.5470 2.9790 17.8970 ;
      RECT 2.8530 17.5470 2.8710 17.8970 ;
      RECT 2.7450 17.5470 2.7630 17.8970 ;
      RECT 2.6370 17.5470 2.6550 17.8970 ;
      RECT 2.5290 17.5470 2.5470 17.8970 ;
      RECT 2.4210 17.5470 2.4390 17.8970 ;
      RECT 2.3130 17.5470 2.3310 17.8970 ;
      RECT 2.2050 17.5470 2.2230 17.8970 ;
      RECT 2.0970 17.5470 2.1150 17.8970 ;
      RECT 1.9890 17.5470 2.0070 17.8970 ;
      RECT 1.8810 17.5470 1.8990 17.8970 ;
      RECT 1.7730 17.5470 1.7910 17.8970 ;
      RECT 1.6650 17.5470 1.6830 17.8970 ;
      RECT 1.5570 17.5470 1.5750 17.8970 ;
      RECT 1.4490 17.5470 1.4670 17.8970 ;
      RECT 1.3410 17.5470 1.3590 17.8970 ;
      RECT 1.2330 17.5470 1.2510 17.8970 ;
      RECT 1.1250 17.5470 1.1430 17.8970 ;
      RECT 1.0170 17.5470 1.0350 17.8970 ;
      RECT 0.9090 17.5470 0.9270 17.8970 ;
      RECT 0.8010 17.5470 0.8190 17.8970 ;
      RECT 0.6930 17.5470 0.7110 17.8970 ;
      RECT 0.5850 17.5470 0.6030 17.8970 ;
      RECT 0.4770 17.5470 0.4950 17.8970 ;
      RECT 0.3690 17.5470 0.3870 17.8970 ;
      RECT 0.2610 17.5470 0.2790 17.8970 ;
      RECT 0.1530 17.5470 0.1710 25.7540 ;
      RECT 0.1170 17.5470 0.1350 25.7540 ;
        RECT 15.6110 25.7520 15.6290 26.6875 ;
        RECT 15.5750 25.7520 15.5930 26.6875 ;
        RECT 15.5390 26.3290 15.5570 26.6515 ;
        RECT 15.4220 26.5260 15.4400 26.6355 ;
        RECT 15.4130 25.7845 15.4310 26.0240 ;
        RECT 15.3770 26.3655 15.3950 26.5190 ;
        RECT 15.2960 26.3910 15.3140 26.6490 ;
        RECT 14.7560 25.7520 14.7740 26.6875 ;
        RECT 14.7200 25.7520 14.7380 26.6875 ;
        RECT 14.6840 25.9330 14.7020 26.5010 ;
        RECT 15.6110 26.8320 15.6290 27.7675 ;
        RECT 15.5750 26.8320 15.5930 27.7675 ;
        RECT 15.5390 27.4090 15.5570 27.7315 ;
        RECT 15.4220 27.6060 15.4400 27.7155 ;
        RECT 15.4130 26.8645 15.4310 27.1040 ;
        RECT 15.3770 27.4455 15.3950 27.5990 ;
        RECT 15.2960 27.4710 15.3140 27.7290 ;
        RECT 14.7560 26.8320 14.7740 27.7675 ;
        RECT 14.7200 26.8320 14.7380 27.7675 ;
        RECT 14.6840 27.0130 14.7020 27.5810 ;
        RECT 15.6110 27.9120 15.6290 28.8475 ;
        RECT 15.5750 27.9120 15.5930 28.8475 ;
        RECT 15.5390 28.4890 15.5570 28.8115 ;
        RECT 15.4220 28.6860 15.4400 28.7955 ;
        RECT 15.4130 27.9445 15.4310 28.1840 ;
        RECT 15.3770 28.5255 15.3950 28.6790 ;
        RECT 15.2960 28.5510 15.3140 28.8090 ;
        RECT 14.7560 27.9120 14.7740 28.8475 ;
        RECT 14.7200 27.9120 14.7380 28.8475 ;
        RECT 14.6840 28.0930 14.7020 28.6610 ;
        RECT 15.6110 28.9920 15.6290 29.9275 ;
        RECT 15.5750 28.9920 15.5930 29.9275 ;
        RECT 15.5390 29.5690 15.5570 29.8915 ;
        RECT 15.4220 29.7660 15.4400 29.8755 ;
        RECT 15.4130 29.0245 15.4310 29.2640 ;
        RECT 15.3770 29.6055 15.3950 29.7590 ;
        RECT 15.2960 29.6310 15.3140 29.8890 ;
        RECT 14.7560 28.9920 14.7740 29.9275 ;
        RECT 14.7200 28.9920 14.7380 29.9275 ;
        RECT 14.6840 29.1730 14.7020 29.7410 ;
        RECT 15.6110 30.0720 15.6290 31.0075 ;
        RECT 15.5750 30.0720 15.5930 31.0075 ;
        RECT 15.5390 30.6490 15.5570 30.9715 ;
        RECT 15.4220 30.8460 15.4400 30.9555 ;
        RECT 15.4130 30.1045 15.4310 30.3440 ;
        RECT 15.3770 30.6855 15.3950 30.8390 ;
        RECT 15.2960 30.7110 15.3140 30.9690 ;
        RECT 14.7560 30.0720 14.7740 31.0075 ;
        RECT 14.7200 30.0720 14.7380 31.0075 ;
        RECT 14.6840 30.2530 14.7020 30.8210 ;
        RECT 15.6110 31.1520 15.6290 32.0875 ;
        RECT 15.5750 31.1520 15.5930 32.0875 ;
        RECT 15.5390 31.7290 15.5570 32.0515 ;
        RECT 15.4220 31.9260 15.4400 32.0355 ;
        RECT 15.4130 31.1845 15.4310 31.4240 ;
        RECT 15.3770 31.7655 15.3950 31.9190 ;
        RECT 15.2960 31.7910 15.3140 32.0490 ;
        RECT 14.7560 31.1520 14.7740 32.0875 ;
        RECT 14.7200 31.1520 14.7380 32.0875 ;
        RECT 14.6840 31.3330 14.7020 31.9010 ;
        RECT 15.6110 32.2320 15.6290 33.1675 ;
        RECT 15.5750 32.2320 15.5930 33.1675 ;
        RECT 15.5390 32.8090 15.5570 33.1315 ;
        RECT 15.4220 33.0060 15.4400 33.1155 ;
        RECT 15.4130 32.2645 15.4310 32.5040 ;
        RECT 15.3770 32.8455 15.3950 32.9990 ;
        RECT 15.2960 32.8710 15.3140 33.1290 ;
        RECT 14.7560 32.2320 14.7740 33.1675 ;
        RECT 14.7200 32.2320 14.7380 33.1675 ;
        RECT 14.6840 32.4130 14.7020 32.9810 ;
        RECT 15.6110 33.3120 15.6290 34.2475 ;
        RECT 15.5750 33.3120 15.5930 34.2475 ;
        RECT 15.5390 33.8890 15.5570 34.2115 ;
        RECT 15.4220 34.0860 15.4400 34.1955 ;
        RECT 15.4130 33.3445 15.4310 33.5840 ;
        RECT 15.3770 33.9255 15.3950 34.0790 ;
        RECT 15.2960 33.9510 15.3140 34.2090 ;
        RECT 14.7560 33.3120 14.7740 34.2475 ;
        RECT 14.7200 33.3120 14.7380 34.2475 ;
        RECT 14.6840 33.4930 14.7020 34.0610 ;
        RECT 15.6110 34.3920 15.6290 35.3275 ;
        RECT 15.5750 34.3920 15.5930 35.3275 ;
        RECT 15.5390 34.9690 15.5570 35.2915 ;
        RECT 15.4220 35.1660 15.4400 35.2755 ;
        RECT 15.4130 34.4245 15.4310 34.6640 ;
        RECT 15.3770 35.0055 15.3950 35.1590 ;
        RECT 15.2960 35.0310 15.3140 35.2890 ;
        RECT 14.7560 34.3920 14.7740 35.3275 ;
        RECT 14.7200 34.3920 14.7380 35.3275 ;
        RECT 14.6840 34.5730 14.7020 35.1410 ;
        RECT 15.6110 35.4720 15.6290 36.4075 ;
        RECT 15.5750 35.4720 15.5930 36.4075 ;
        RECT 15.5390 36.0490 15.5570 36.3715 ;
        RECT 15.4220 36.2460 15.4400 36.3555 ;
        RECT 15.4130 35.5045 15.4310 35.7440 ;
        RECT 15.3770 36.0855 15.3950 36.2390 ;
        RECT 15.2960 36.1110 15.3140 36.3690 ;
        RECT 14.7560 35.4720 14.7740 36.4075 ;
        RECT 14.7200 35.4720 14.7380 36.4075 ;
        RECT 14.6840 35.6530 14.7020 36.2210 ;
        RECT 15.6110 36.5520 15.6290 37.4875 ;
        RECT 15.5750 36.5520 15.5930 37.4875 ;
        RECT 15.5390 37.1290 15.5570 37.4515 ;
        RECT 15.4220 37.3260 15.4400 37.4355 ;
        RECT 15.4130 36.5845 15.4310 36.8240 ;
        RECT 15.3770 37.1655 15.3950 37.3190 ;
        RECT 15.2960 37.1910 15.3140 37.4490 ;
        RECT 14.7560 36.5520 14.7740 37.4875 ;
        RECT 14.7200 36.5520 14.7380 37.4875 ;
        RECT 14.6840 36.7330 14.7020 37.3010 ;
        RECT 15.6110 37.6320 15.6290 38.5675 ;
        RECT 15.5750 37.6320 15.5930 38.5675 ;
        RECT 15.5390 38.2090 15.5570 38.5315 ;
        RECT 15.4220 38.4060 15.4400 38.5155 ;
        RECT 15.4130 37.6645 15.4310 37.9040 ;
        RECT 15.3770 38.2455 15.3950 38.3990 ;
        RECT 15.2960 38.2710 15.3140 38.5290 ;
        RECT 14.7560 37.6320 14.7740 38.5675 ;
        RECT 14.7200 37.6320 14.7380 38.5675 ;
        RECT 14.6840 37.8130 14.7020 38.3810 ;
        RECT 15.6110 38.7120 15.6290 39.6475 ;
        RECT 15.5750 38.7120 15.5930 39.6475 ;
        RECT 15.5390 39.2890 15.5570 39.6115 ;
        RECT 15.4220 39.4860 15.4400 39.5955 ;
        RECT 15.4130 38.7445 15.4310 38.9840 ;
        RECT 15.3770 39.3255 15.3950 39.4790 ;
        RECT 15.2960 39.3510 15.3140 39.6090 ;
        RECT 14.7560 38.7120 14.7740 39.6475 ;
        RECT 14.7200 38.7120 14.7380 39.6475 ;
        RECT 14.6840 38.8930 14.7020 39.4610 ;
        RECT 15.6110 39.7920 15.6290 40.7275 ;
        RECT 15.5750 39.7920 15.5930 40.7275 ;
        RECT 15.5390 40.3690 15.5570 40.6915 ;
        RECT 15.4220 40.5660 15.4400 40.6755 ;
        RECT 15.4130 39.8245 15.4310 40.0640 ;
        RECT 15.3770 40.4055 15.3950 40.5590 ;
        RECT 15.2960 40.4310 15.3140 40.6890 ;
        RECT 14.7560 39.7920 14.7740 40.7275 ;
        RECT 14.7200 39.7920 14.7380 40.7275 ;
        RECT 14.6840 39.9730 14.7020 40.5410 ;
        RECT 15.6110 40.8720 15.6290 41.8075 ;
        RECT 15.5750 40.8720 15.5930 41.8075 ;
        RECT 15.5390 41.4490 15.5570 41.7715 ;
        RECT 15.4220 41.6460 15.4400 41.7555 ;
        RECT 15.4130 40.9045 15.4310 41.1440 ;
        RECT 15.3770 41.4855 15.3950 41.6390 ;
        RECT 15.2960 41.5110 15.3140 41.7690 ;
        RECT 14.7560 40.8720 14.7740 41.8075 ;
        RECT 14.7200 40.8720 14.7380 41.8075 ;
        RECT 14.6840 41.0530 14.7020 41.6210 ;
        RECT 15.6110 41.9520 15.6290 42.8875 ;
        RECT 15.5750 41.9520 15.5930 42.8875 ;
        RECT 15.5390 42.5290 15.5570 42.8515 ;
        RECT 15.4220 42.7260 15.4400 42.8355 ;
        RECT 15.4130 41.9845 15.4310 42.2240 ;
        RECT 15.3770 42.5655 15.3950 42.7190 ;
        RECT 15.2960 42.5910 15.3140 42.8490 ;
        RECT 14.7560 41.9520 14.7740 42.8875 ;
        RECT 14.7200 41.9520 14.7380 42.8875 ;
        RECT 14.6840 42.1330 14.7020 42.7010 ;
  LAYER M3 SPACING 0.018  ;
      RECT 15.5530 0.2565 15.6810 1.3500 ;
      RECT 15.5390 0.9220 15.6810 1.2445 ;
      RECT 15.3190 0.6490 15.4530 1.3500 ;
      RECT 15.2960 0.9840 15.4530 1.2420 ;
      RECT 15.3190 0.2565 15.4170 1.3500 ;
      RECT 15.3190 0.3775 15.4310 0.6170 ;
      RECT 15.3190 0.2565 15.4530 0.3455 ;
      RECT 15.0940 0.7070 15.2280 1.3500 ;
      RECT 15.0940 0.2565 15.1920 1.3500 ;
      RECT 14.6770 0.2565 14.7600 1.3500 ;
      RECT 14.6770 0.3450 14.7740 1.2805 ;
      RECT 30.2680 0.2565 30.3530 1.3500 ;
      RECT 30.1240 0.2565 30.1500 1.3500 ;
      RECT 30.0160 0.2565 30.0420 1.3500 ;
      RECT 29.9080 0.2565 29.9340 1.3500 ;
      RECT 29.8000 0.2565 29.8260 1.3500 ;
      RECT 29.6920 0.2565 29.7180 1.3500 ;
      RECT 29.5840 0.2565 29.6100 1.3500 ;
      RECT 29.4760 0.2565 29.5020 1.3500 ;
      RECT 29.3680 0.2565 29.3940 1.3500 ;
      RECT 29.2600 0.2565 29.2860 1.3500 ;
      RECT 29.1520 0.2565 29.1780 1.3500 ;
      RECT 29.0440 0.2565 29.0700 1.3500 ;
      RECT 28.9360 0.2565 28.9620 1.3500 ;
      RECT 28.8280 0.2565 28.8540 1.3500 ;
      RECT 28.7200 0.2565 28.7460 1.3500 ;
      RECT 28.6120 0.2565 28.6380 1.3500 ;
      RECT 28.5040 0.2565 28.5300 1.3500 ;
      RECT 28.3960 0.2565 28.4220 1.3500 ;
      RECT 28.2880 0.2565 28.3140 1.3500 ;
      RECT 28.1800 0.2565 28.2060 1.3500 ;
      RECT 28.0720 0.2565 28.0980 1.3500 ;
      RECT 27.9640 0.2565 27.9900 1.3500 ;
      RECT 27.8560 0.2565 27.8820 1.3500 ;
      RECT 27.7480 0.2565 27.7740 1.3500 ;
      RECT 27.6400 0.2565 27.6660 1.3500 ;
      RECT 27.5320 0.2565 27.5580 1.3500 ;
      RECT 27.4240 0.2565 27.4500 1.3500 ;
      RECT 27.3160 0.2565 27.3420 1.3500 ;
      RECT 27.2080 0.2565 27.2340 1.3500 ;
      RECT 27.1000 0.2565 27.1260 1.3500 ;
      RECT 26.9920 0.2565 27.0180 1.3500 ;
      RECT 26.8840 0.2565 26.9100 1.3500 ;
      RECT 26.7760 0.2565 26.8020 1.3500 ;
      RECT 26.6680 0.2565 26.6940 1.3500 ;
      RECT 26.5600 0.2565 26.5860 1.3500 ;
      RECT 26.4520 0.2565 26.4780 1.3500 ;
      RECT 26.3440 0.2565 26.3700 1.3500 ;
      RECT 26.2360 0.2565 26.2620 1.3500 ;
      RECT 26.1280 0.2565 26.1540 1.3500 ;
      RECT 26.0200 0.2565 26.0460 1.3500 ;
      RECT 25.9120 0.2565 25.9380 1.3500 ;
      RECT 25.8040 0.2565 25.8300 1.3500 ;
      RECT 25.6960 0.2565 25.7220 1.3500 ;
      RECT 25.5880 0.2565 25.6140 1.3500 ;
      RECT 25.4800 0.2565 25.5060 1.3500 ;
      RECT 25.3720 0.2565 25.3980 1.3500 ;
      RECT 25.2640 0.2565 25.2900 1.3500 ;
      RECT 25.1560 0.2565 25.1820 1.3500 ;
      RECT 25.0480 0.2565 25.0740 1.3500 ;
      RECT 24.9400 0.2565 24.9660 1.3500 ;
      RECT 24.8320 0.2565 24.8580 1.3500 ;
      RECT 24.7240 0.2565 24.7500 1.3500 ;
      RECT 24.6160 0.2565 24.6420 1.3500 ;
      RECT 24.5080 0.2565 24.5340 1.3500 ;
      RECT 24.4000 0.2565 24.4260 1.3500 ;
      RECT 24.2920 0.2565 24.3180 1.3500 ;
      RECT 24.1840 0.2565 24.2100 1.3500 ;
      RECT 24.0760 0.2565 24.1020 1.3500 ;
      RECT 23.9680 0.2565 23.9940 1.3500 ;
      RECT 23.8600 0.2565 23.8860 1.3500 ;
      RECT 23.7520 0.2565 23.7780 1.3500 ;
      RECT 23.6440 0.2565 23.6700 1.3500 ;
      RECT 23.5360 0.2565 23.5620 1.3500 ;
      RECT 23.4280 0.2565 23.4540 1.3500 ;
      RECT 23.3200 0.2565 23.3460 1.3500 ;
      RECT 23.2120 0.2565 23.2380 1.3500 ;
      RECT 23.1040 0.2565 23.1300 1.3500 ;
      RECT 22.9960 0.2565 23.0220 1.3500 ;
      RECT 22.8880 0.2565 22.9140 1.3500 ;
      RECT 22.7800 0.2565 22.8060 1.3500 ;
      RECT 22.6720 0.2565 22.6980 1.3500 ;
      RECT 22.5640 0.2565 22.5900 1.3500 ;
      RECT 22.4560 0.2565 22.4820 1.3500 ;
      RECT 22.3480 0.2565 22.3740 1.3500 ;
      RECT 22.2400 0.2565 22.2660 1.3500 ;
      RECT 22.1320 0.2565 22.1580 1.3500 ;
      RECT 22.0240 0.2565 22.0500 1.3500 ;
      RECT 21.9160 0.2565 21.9420 1.3500 ;
      RECT 21.8080 0.2565 21.8340 1.3500 ;
      RECT 21.7000 0.2565 21.7260 1.3500 ;
      RECT 21.5920 0.2565 21.6180 1.3500 ;
      RECT 21.4840 0.2565 21.5100 1.3500 ;
      RECT 21.3760 0.2565 21.4020 1.3500 ;
      RECT 21.2680 0.2565 21.2940 1.3500 ;
      RECT 21.1600 0.2565 21.1860 1.3500 ;
      RECT 21.0520 0.2565 21.0780 1.3500 ;
      RECT 20.9440 0.2565 20.9700 1.3500 ;
      RECT 20.8360 0.2565 20.8620 1.3500 ;
      RECT 20.7280 0.2565 20.7540 1.3500 ;
      RECT 20.6200 0.2565 20.6460 1.3500 ;
      RECT 20.5120 0.2565 20.5380 1.3500 ;
      RECT 20.4040 0.2565 20.4300 1.3500 ;
      RECT 20.2960 0.2565 20.3220 1.3500 ;
      RECT 20.1880 0.2565 20.2140 1.3500 ;
      RECT 20.0800 0.2565 20.1060 1.3500 ;
      RECT 19.9720 0.2565 19.9980 1.3500 ;
      RECT 19.8640 0.2565 19.8900 1.3500 ;
      RECT 19.7560 0.2565 19.7820 1.3500 ;
      RECT 19.6480 0.2565 19.6740 1.3500 ;
      RECT 19.5400 0.2565 19.5660 1.3500 ;
      RECT 19.4320 0.2565 19.4580 1.3500 ;
      RECT 19.3240 0.2565 19.3500 1.3500 ;
      RECT 19.2160 0.2565 19.2420 1.3500 ;
      RECT 19.1080 0.2565 19.1340 1.3500 ;
      RECT 19.0000 0.2565 19.0260 1.3500 ;
      RECT 18.8920 0.2565 18.9180 1.3500 ;
      RECT 18.7840 0.2565 18.8100 1.3500 ;
      RECT 18.6760 0.2565 18.7020 1.3500 ;
      RECT 18.5680 0.2565 18.5940 1.3500 ;
      RECT 18.4600 0.2565 18.4860 1.3500 ;
      RECT 18.3520 0.2565 18.3780 1.3500 ;
      RECT 18.2440 0.2565 18.2700 1.3500 ;
      RECT 18.1360 0.2565 18.1620 1.3500 ;
      RECT 18.0280 0.2565 18.0540 1.3500 ;
      RECT 17.9200 0.2565 17.9460 1.3500 ;
      RECT 17.8120 0.2565 17.8380 1.3500 ;
      RECT 17.7040 0.2565 17.7300 1.3500 ;
      RECT 17.5960 0.2565 17.6220 1.3500 ;
      RECT 17.4880 0.2565 17.5140 1.3500 ;
      RECT 17.3800 0.2565 17.4060 1.3500 ;
      RECT 17.2720 0.2565 17.2980 1.3500 ;
      RECT 17.1640 0.2565 17.1900 1.3500 ;
      RECT 17.0560 0.2565 17.0820 1.3500 ;
      RECT 16.9480 0.2565 16.9740 1.3500 ;
      RECT 16.8400 0.2565 16.8660 1.3500 ;
      RECT 16.7320 0.2565 16.7580 1.3500 ;
      RECT 16.6240 0.2565 16.6500 1.3500 ;
      RECT 16.5160 0.2565 16.5420 1.3500 ;
      RECT 16.4080 0.2565 16.4340 1.3500 ;
      RECT 16.3000 0.2565 16.3260 1.3500 ;
      RECT 16.0870 0.2565 16.1640 1.3500 ;
      RECT 14.1940 0.2565 14.2710 1.3500 ;
      RECT 14.0320 0.2565 14.0580 1.3500 ;
      RECT 13.9240 0.2565 13.9500 1.3500 ;
      RECT 13.8160 0.2565 13.8420 1.3500 ;
      RECT 13.7080 0.2565 13.7340 1.3500 ;
      RECT 13.6000 0.2565 13.6260 1.3500 ;
      RECT 13.4920 0.2565 13.5180 1.3500 ;
      RECT 13.3840 0.2565 13.4100 1.3500 ;
      RECT 13.2760 0.2565 13.3020 1.3500 ;
      RECT 13.1680 0.2565 13.1940 1.3500 ;
      RECT 13.0600 0.2565 13.0860 1.3500 ;
      RECT 12.9520 0.2565 12.9780 1.3500 ;
      RECT 12.8440 0.2565 12.8700 1.3500 ;
      RECT 12.7360 0.2565 12.7620 1.3500 ;
      RECT 12.6280 0.2565 12.6540 1.3500 ;
      RECT 12.5200 0.2565 12.5460 1.3500 ;
      RECT 12.4120 0.2565 12.4380 1.3500 ;
      RECT 12.3040 0.2565 12.3300 1.3500 ;
      RECT 12.1960 0.2565 12.2220 1.3500 ;
      RECT 12.0880 0.2565 12.1140 1.3500 ;
      RECT 11.9800 0.2565 12.0060 1.3500 ;
      RECT 11.8720 0.2565 11.8980 1.3500 ;
      RECT 11.7640 0.2565 11.7900 1.3500 ;
      RECT 11.6560 0.2565 11.6820 1.3500 ;
      RECT 11.5480 0.2565 11.5740 1.3500 ;
      RECT 11.4400 0.2565 11.4660 1.3500 ;
      RECT 11.3320 0.2565 11.3580 1.3500 ;
      RECT 11.2240 0.2565 11.2500 1.3500 ;
      RECT 11.1160 0.2565 11.1420 1.3500 ;
      RECT 11.0080 0.2565 11.0340 1.3500 ;
      RECT 10.9000 0.2565 10.9260 1.3500 ;
      RECT 10.7920 0.2565 10.8180 1.3500 ;
      RECT 10.6840 0.2565 10.7100 1.3500 ;
      RECT 10.5760 0.2565 10.6020 1.3500 ;
      RECT 10.4680 0.2565 10.4940 1.3500 ;
      RECT 10.3600 0.2565 10.3860 1.3500 ;
      RECT 10.2520 0.2565 10.2780 1.3500 ;
      RECT 10.1440 0.2565 10.1700 1.3500 ;
      RECT 10.0360 0.2565 10.0620 1.3500 ;
      RECT 9.9280 0.2565 9.9540 1.3500 ;
      RECT 9.8200 0.2565 9.8460 1.3500 ;
      RECT 9.7120 0.2565 9.7380 1.3500 ;
      RECT 9.6040 0.2565 9.6300 1.3500 ;
      RECT 9.4960 0.2565 9.5220 1.3500 ;
      RECT 9.3880 0.2565 9.4140 1.3500 ;
      RECT 9.2800 0.2565 9.3060 1.3500 ;
      RECT 9.1720 0.2565 9.1980 1.3500 ;
      RECT 9.0640 0.2565 9.0900 1.3500 ;
      RECT 8.9560 0.2565 8.9820 1.3500 ;
      RECT 8.8480 0.2565 8.8740 1.3500 ;
      RECT 8.7400 0.2565 8.7660 1.3500 ;
      RECT 8.6320 0.2565 8.6580 1.3500 ;
      RECT 8.5240 0.2565 8.5500 1.3500 ;
      RECT 8.4160 0.2565 8.4420 1.3500 ;
      RECT 8.3080 0.2565 8.3340 1.3500 ;
      RECT 8.2000 0.2565 8.2260 1.3500 ;
      RECT 8.0920 0.2565 8.1180 1.3500 ;
      RECT 7.9840 0.2565 8.0100 1.3500 ;
      RECT 7.8760 0.2565 7.9020 1.3500 ;
      RECT 7.7680 0.2565 7.7940 1.3500 ;
      RECT 7.6600 0.2565 7.6860 1.3500 ;
      RECT 7.5520 0.2565 7.5780 1.3500 ;
      RECT 7.4440 0.2565 7.4700 1.3500 ;
      RECT 7.3360 0.2565 7.3620 1.3500 ;
      RECT 7.2280 0.2565 7.2540 1.3500 ;
      RECT 7.1200 0.2565 7.1460 1.3500 ;
      RECT 7.0120 0.2565 7.0380 1.3500 ;
      RECT 6.9040 0.2565 6.9300 1.3500 ;
      RECT 6.7960 0.2565 6.8220 1.3500 ;
      RECT 6.6880 0.2565 6.7140 1.3500 ;
      RECT 6.5800 0.2565 6.6060 1.3500 ;
      RECT 6.4720 0.2565 6.4980 1.3500 ;
      RECT 6.3640 0.2565 6.3900 1.3500 ;
      RECT 6.2560 0.2565 6.2820 1.3500 ;
      RECT 6.1480 0.2565 6.1740 1.3500 ;
      RECT 6.0400 0.2565 6.0660 1.3500 ;
      RECT 5.9320 0.2565 5.9580 1.3500 ;
      RECT 5.8240 0.2565 5.8500 1.3500 ;
      RECT 5.7160 0.2565 5.7420 1.3500 ;
      RECT 5.6080 0.2565 5.6340 1.3500 ;
      RECT 5.5000 0.2565 5.5260 1.3500 ;
      RECT 5.3920 0.2565 5.4180 1.3500 ;
      RECT 5.2840 0.2565 5.3100 1.3500 ;
      RECT 5.1760 0.2565 5.2020 1.3500 ;
      RECT 5.0680 0.2565 5.0940 1.3500 ;
      RECT 4.9600 0.2565 4.9860 1.3500 ;
      RECT 4.8520 0.2565 4.8780 1.3500 ;
      RECT 4.7440 0.2565 4.7700 1.3500 ;
      RECT 4.6360 0.2565 4.6620 1.3500 ;
      RECT 4.5280 0.2565 4.5540 1.3500 ;
      RECT 4.4200 0.2565 4.4460 1.3500 ;
      RECT 4.3120 0.2565 4.3380 1.3500 ;
      RECT 4.2040 0.2565 4.2300 1.3500 ;
      RECT 4.0960 0.2565 4.1220 1.3500 ;
      RECT 3.9880 0.2565 4.0140 1.3500 ;
      RECT 3.8800 0.2565 3.9060 1.3500 ;
      RECT 3.7720 0.2565 3.7980 1.3500 ;
      RECT 3.6640 0.2565 3.6900 1.3500 ;
      RECT 3.5560 0.2565 3.5820 1.3500 ;
      RECT 3.4480 0.2565 3.4740 1.3500 ;
      RECT 3.3400 0.2565 3.3660 1.3500 ;
      RECT 3.2320 0.2565 3.2580 1.3500 ;
      RECT 3.1240 0.2565 3.1500 1.3500 ;
      RECT 3.0160 0.2565 3.0420 1.3500 ;
      RECT 2.9080 0.2565 2.9340 1.3500 ;
      RECT 2.8000 0.2565 2.8260 1.3500 ;
      RECT 2.6920 0.2565 2.7180 1.3500 ;
      RECT 2.5840 0.2565 2.6100 1.3500 ;
      RECT 2.4760 0.2565 2.5020 1.3500 ;
      RECT 2.3680 0.2565 2.3940 1.3500 ;
      RECT 2.2600 0.2565 2.2860 1.3500 ;
      RECT 2.1520 0.2565 2.1780 1.3500 ;
      RECT 2.0440 0.2565 2.0700 1.3500 ;
      RECT 1.9360 0.2565 1.9620 1.3500 ;
      RECT 1.8280 0.2565 1.8540 1.3500 ;
      RECT 1.7200 0.2565 1.7460 1.3500 ;
      RECT 1.6120 0.2565 1.6380 1.3500 ;
      RECT 1.5040 0.2565 1.5300 1.3500 ;
      RECT 1.3960 0.2565 1.4220 1.3500 ;
      RECT 1.2880 0.2565 1.3140 1.3500 ;
      RECT 1.1800 0.2565 1.2060 1.3500 ;
      RECT 1.0720 0.2565 1.0980 1.3500 ;
      RECT 0.9640 0.2565 0.9900 1.3500 ;
      RECT 0.8560 0.2565 0.8820 1.3500 ;
      RECT 0.7480 0.2565 0.7740 1.3500 ;
      RECT 0.6400 0.2565 0.6660 1.3500 ;
      RECT 0.5320 0.2565 0.5580 1.3500 ;
      RECT 0.4240 0.2565 0.4500 1.3500 ;
      RECT 0.3160 0.2565 0.3420 1.3500 ;
      RECT 0.2080 0.2565 0.2340 1.3500 ;
      RECT 0.0050 0.2565 0.0900 1.3500 ;
      RECT 15.5530 1.3365 15.6810 2.4300 ;
      RECT 15.5390 2.0020 15.6810 2.3245 ;
      RECT 15.3190 1.7290 15.4530 2.4300 ;
      RECT 15.2960 2.0640 15.4530 2.3220 ;
      RECT 15.3190 1.3365 15.4170 2.4300 ;
      RECT 15.3190 1.4575 15.4310 1.6970 ;
      RECT 15.3190 1.3365 15.4530 1.4255 ;
      RECT 15.0940 1.7870 15.2280 2.4300 ;
      RECT 15.0940 1.3365 15.1920 2.4300 ;
      RECT 14.6770 1.3365 14.7600 2.4300 ;
      RECT 14.6770 1.4250 14.7740 2.3605 ;
      RECT 30.2680 1.3365 30.3530 2.4300 ;
      RECT 30.1240 1.3365 30.1500 2.4300 ;
      RECT 30.0160 1.3365 30.0420 2.4300 ;
      RECT 29.9080 1.3365 29.9340 2.4300 ;
      RECT 29.8000 1.3365 29.8260 2.4300 ;
      RECT 29.6920 1.3365 29.7180 2.4300 ;
      RECT 29.5840 1.3365 29.6100 2.4300 ;
      RECT 29.4760 1.3365 29.5020 2.4300 ;
      RECT 29.3680 1.3365 29.3940 2.4300 ;
      RECT 29.2600 1.3365 29.2860 2.4300 ;
      RECT 29.1520 1.3365 29.1780 2.4300 ;
      RECT 29.0440 1.3365 29.0700 2.4300 ;
      RECT 28.9360 1.3365 28.9620 2.4300 ;
      RECT 28.8280 1.3365 28.8540 2.4300 ;
      RECT 28.7200 1.3365 28.7460 2.4300 ;
      RECT 28.6120 1.3365 28.6380 2.4300 ;
      RECT 28.5040 1.3365 28.5300 2.4300 ;
      RECT 28.3960 1.3365 28.4220 2.4300 ;
      RECT 28.2880 1.3365 28.3140 2.4300 ;
      RECT 28.1800 1.3365 28.2060 2.4300 ;
      RECT 28.0720 1.3365 28.0980 2.4300 ;
      RECT 27.9640 1.3365 27.9900 2.4300 ;
      RECT 27.8560 1.3365 27.8820 2.4300 ;
      RECT 27.7480 1.3365 27.7740 2.4300 ;
      RECT 27.6400 1.3365 27.6660 2.4300 ;
      RECT 27.5320 1.3365 27.5580 2.4300 ;
      RECT 27.4240 1.3365 27.4500 2.4300 ;
      RECT 27.3160 1.3365 27.3420 2.4300 ;
      RECT 27.2080 1.3365 27.2340 2.4300 ;
      RECT 27.1000 1.3365 27.1260 2.4300 ;
      RECT 26.9920 1.3365 27.0180 2.4300 ;
      RECT 26.8840 1.3365 26.9100 2.4300 ;
      RECT 26.7760 1.3365 26.8020 2.4300 ;
      RECT 26.6680 1.3365 26.6940 2.4300 ;
      RECT 26.5600 1.3365 26.5860 2.4300 ;
      RECT 26.4520 1.3365 26.4780 2.4300 ;
      RECT 26.3440 1.3365 26.3700 2.4300 ;
      RECT 26.2360 1.3365 26.2620 2.4300 ;
      RECT 26.1280 1.3365 26.1540 2.4300 ;
      RECT 26.0200 1.3365 26.0460 2.4300 ;
      RECT 25.9120 1.3365 25.9380 2.4300 ;
      RECT 25.8040 1.3365 25.8300 2.4300 ;
      RECT 25.6960 1.3365 25.7220 2.4300 ;
      RECT 25.5880 1.3365 25.6140 2.4300 ;
      RECT 25.4800 1.3365 25.5060 2.4300 ;
      RECT 25.3720 1.3365 25.3980 2.4300 ;
      RECT 25.2640 1.3365 25.2900 2.4300 ;
      RECT 25.1560 1.3365 25.1820 2.4300 ;
      RECT 25.0480 1.3365 25.0740 2.4300 ;
      RECT 24.9400 1.3365 24.9660 2.4300 ;
      RECT 24.8320 1.3365 24.8580 2.4300 ;
      RECT 24.7240 1.3365 24.7500 2.4300 ;
      RECT 24.6160 1.3365 24.6420 2.4300 ;
      RECT 24.5080 1.3365 24.5340 2.4300 ;
      RECT 24.4000 1.3365 24.4260 2.4300 ;
      RECT 24.2920 1.3365 24.3180 2.4300 ;
      RECT 24.1840 1.3365 24.2100 2.4300 ;
      RECT 24.0760 1.3365 24.1020 2.4300 ;
      RECT 23.9680 1.3365 23.9940 2.4300 ;
      RECT 23.8600 1.3365 23.8860 2.4300 ;
      RECT 23.7520 1.3365 23.7780 2.4300 ;
      RECT 23.6440 1.3365 23.6700 2.4300 ;
      RECT 23.5360 1.3365 23.5620 2.4300 ;
      RECT 23.4280 1.3365 23.4540 2.4300 ;
      RECT 23.3200 1.3365 23.3460 2.4300 ;
      RECT 23.2120 1.3365 23.2380 2.4300 ;
      RECT 23.1040 1.3365 23.1300 2.4300 ;
      RECT 22.9960 1.3365 23.0220 2.4300 ;
      RECT 22.8880 1.3365 22.9140 2.4300 ;
      RECT 22.7800 1.3365 22.8060 2.4300 ;
      RECT 22.6720 1.3365 22.6980 2.4300 ;
      RECT 22.5640 1.3365 22.5900 2.4300 ;
      RECT 22.4560 1.3365 22.4820 2.4300 ;
      RECT 22.3480 1.3365 22.3740 2.4300 ;
      RECT 22.2400 1.3365 22.2660 2.4300 ;
      RECT 22.1320 1.3365 22.1580 2.4300 ;
      RECT 22.0240 1.3365 22.0500 2.4300 ;
      RECT 21.9160 1.3365 21.9420 2.4300 ;
      RECT 21.8080 1.3365 21.8340 2.4300 ;
      RECT 21.7000 1.3365 21.7260 2.4300 ;
      RECT 21.5920 1.3365 21.6180 2.4300 ;
      RECT 21.4840 1.3365 21.5100 2.4300 ;
      RECT 21.3760 1.3365 21.4020 2.4300 ;
      RECT 21.2680 1.3365 21.2940 2.4300 ;
      RECT 21.1600 1.3365 21.1860 2.4300 ;
      RECT 21.0520 1.3365 21.0780 2.4300 ;
      RECT 20.9440 1.3365 20.9700 2.4300 ;
      RECT 20.8360 1.3365 20.8620 2.4300 ;
      RECT 20.7280 1.3365 20.7540 2.4300 ;
      RECT 20.6200 1.3365 20.6460 2.4300 ;
      RECT 20.5120 1.3365 20.5380 2.4300 ;
      RECT 20.4040 1.3365 20.4300 2.4300 ;
      RECT 20.2960 1.3365 20.3220 2.4300 ;
      RECT 20.1880 1.3365 20.2140 2.4300 ;
      RECT 20.0800 1.3365 20.1060 2.4300 ;
      RECT 19.9720 1.3365 19.9980 2.4300 ;
      RECT 19.8640 1.3365 19.8900 2.4300 ;
      RECT 19.7560 1.3365 19.7820 2.4300 ;
      RECT 19.6480 1.3365 19.6740 2.4300 ;
      RECT 19.5400 1.3365 19.5660 2.4300 ;
      RECT 19.4320 1.3365 19.4580 2.4300 ;
      RECT 19.3240 1.3365 19.3500 2.4300 ;
      RECT 19.2160 1.3365 19.2420 2.4300 ;
      RECT 19.1080 1.3365 19.1340 2.4300 ;
      RECT 19.0000 1.3365 19.0260 2.4300 ;
      RECT 18.8920 1.3365 18.9180 2.4300 ;
      RECT 18.7840 1.3365 18.8100 2.4300 ;
      RECT 18.6760 1.3365 18.7020 2.4300 ;
      RECT 18.5680 1.3365 18.5940 2.4300 ;
      RECT 18.4600 1.3365 18.4860 2.4300 ;
      RECT 18.3520 1.3365 18.3780 2.4300 ;
      RECT 18.2440 1.3365 18.2700 2.4300 ;
      RECT 18.1360 1.3365 18.1620 2.4300 ;
      RECT 18.0280 1.3365 18.0540 2.4300 ;
      RECT 17.9200 1.3365 17.9460 2.4300 ;
      RECT 17.8120 1.3365 17.8380 2.4300 ;
      RECT 17.7040 1.3365 17.7300 2.4300 ;
      RECT 17.5960 1.3365 17.6220 2.4300 ;
      RECT 17.4880 1.3365 17.5140 2.4300 ;
      RECT 17.3800 1.3365 17.4060 2.4300 ;
      RECT 17.2720 1.3365 17.2980 2.4300 ;
      RECT 17.1640 1.3365 17.1900 2.4300 ;
      RECT 17.0560 1.3365 17.0820 2.4300 ;
      RECT 16.9480 1.3365 16.9740 2.4300 ;
      RECT 16.8400 1.3365 16.8660 2.4300 ;
      RECT 16.7320 1.3365 16.7580 2.4300 ;
      RECT 16.6240 1.3365 16.6500 2.4300 ;
      RECT 16.5160 1.3365 16.5420 2.4300 ;
      RECT 16.4080 1.3365 16.4340 2.4300 ;
      RECT 16.3000 1.3365 16.3260 2.4300 ;
      RECT 16.0870 1.3365 16.1640 2.4300 ;
      RECT 14.1940 1.3365 14.2710 2.4300 ;
      RECT 14.0320 1.3365 14.0580 2.4300 ;
      RECT 13.9240 1.3365 13.9500 2.4300 ;
      RECT 13.8160 1.3365 13.8420 2.4300 ;
      RECT 13.7080 1.3365 13.7340 2.4300 ;
      RECT 13.6000 1.3365 13.6260 2.4300 ;
      RECT 13.4920 1.3365 13.5180 2.4300 ;
      RECT 13.3840 1.3365 13.4100 2.4300 ;
      RECT 13.2760 1.3365 13.3020 2.4300 ;
      RECT 13.1680 1.3365 13.1940 2.4300 ;
      RECT 13.0600 1.3365 13.0860 2.4300 ;
      RECT 12.9520 1.3365 12.9780 2.4300 ;
      RECT 12.8440 1.3365 12.8700 2.4300 ;
      RECT 12.7360 1.3365 12.7620 2.4300 ;
      RECT 12.6280 1.3365 12.6540 2.4300 ;
      RECT 12.5200 1.3365 12.5460 2.4300 ;
      RECT 12.4120 1.3365 12.4380 2.4300 ;
      RECT 12.3040 1.3365 12.3300 2.4300 ;
      RECT 12.1960 1.3365 12.2220 2.4300 ;
      RECT 12.0880 1.3365 12.1140 2.4300 ;
      RECT 11.9800 1.3365 12.0060 2.4300 ;
      RECT 11.8720 1.3365 11.8980 2.4300 ;
      RECT 11.7640 1.3365 11.7900 2.4300 ;
      RECT 11.6560 1.3365 11.6820 2.4300 ;
      RECT 11.5480 1.3365 11.5740 2.4300 ;
      RECT 11.4400 1.3365 11.4660 2.4300 ;
      RECT 11.3320 1.3365 11.3580 2.4300 ;
      RECT 11.2240 1.3365 11.2500 2.4300 ;
      RECT 11.1160 1.3365 11.1420 2.4300 ;
      RECT 11.0080 1.3365 11.0340 2.4300 ;
      RECT 10.9000 1.3365 10.9260 2.4300 ;
      RECT 10.7920 1.3365 10.8180 2.4300 ;
      RECT 10.6840 1.3365 10.7100 2.4300 ;
      RECT 10.5760 1.3365 10.6020 2.4300 ;
      RECT 10.4680 1.3365 10.4940 2.4300 ;
      RECT 10.3600 1.3365 10.3860 2.4300 ;
      RECT 10.2520 1.3365 10.2780 2.4300 ;
      RECT 10.1440 1.3365 10.1700 2.4300 ;
      RECT 10.0360 1.3365 10.0620 2.4300 ;
      RECT 9.9280 1.3365 9.9540 2.4300 ;
      RECT 9.8200 1.3365 9.8460 2.4300 ;
      RECT 9.7120 1.3365 9.7380 2.4300 ;
      RECT 9.6040 1.3365 9.6300 2.4300 ;
      RECT 9.4960 1.3365 9.5220 2.4300 ;
      RECT 9.3880 1.3365 9.4140 2.4300 ;
      RECT 9.2800 1.3365 9.3060 2.4300 ;
      RECT 9.1720 1.3365 9.1980 2.4300 ;
      RECT 9.0640 1.3365 9.0900 2.4300 ;
      RECT 8.9560 1.3365 8.9820 2.4300 ;
      RECT 8.8480 1.3365 8.8740 2.4300 ;
      RECT 8.7400 1.3365 8.7660 2.4300 ;
      RECT 8.6320 1.3365 8.6580 2.4300 ;
      RECT 8.5240 1.3365 8.5500 2.4300 ;
      RECT 8.4160 1.3365 8.4420 2.4300 ;
      RECT 8.3080 1.3365 8.3340 2.4300 ;
      RECT 8.2000 1.3365 8.2260 2.4300 ;
      RECT 8.0920 1.3365 8.1180 2.4300 ;
      RECT 7.9840 1.3365 8.0100 2.4300 ;
      RECT 7.8760 1.3365 7.9020 2.4300 ;
      RECT 7.7680 1.3365 7.7940 2.4300 ;
      RECT 7.6600 1.3365 7.6860 2.4300 ;
      RECT 7.5520 1.3365 7.5780 2.4300 ;
      RECT 7.4440 1.3365 7.4700 2.4300 ;
      RECT 7.3360 1.3365 7.3620 2.4300 ;
      RECT 7.2280 1.3365 7.2540 2.4300 ;
      RECT 7.1200 1.3365 7.1460 2.4300 ;
      RECT 7.0120 1.3365 7.0380 2.4300 ;
      RECT 6.9040 1.3365 6.9300 2.4300 ;
      RECT 6.7960 1.3365 6.8220 2.4300 ;
      RECT 6.6880 1.3365 6.7140 2.4300 ;
      RECT 6.5800 1.3365 6.6060 2.4300 ;
      RECT 6.4720 1.3365 6.4980 2.4300 ;
      RECT 6.3640 1.3365 6.3900 2.4300 ;
      RECT 6.2560 1.3365 6.2820 2.4300 ;
      RECT 6.1480 1.3365 6.1740 2.4300 ;
      RECT 6.0400 1.3365 6.0660 2.4300 ;
      RECT 5.9320 1.3365 5.9580 2.4300 ;
      RECT 5.8240 1.3365 5.8500 2.4300 ;
      RECT 5.7160 1.3365 5.7420 2.4300 ;
      RECT 5.6080 1.3365 5.6340 2.4300 ;
      RECT 5.5000 1.3365 5.5260 2.4300 ;
      RECT 5.3920 1.3365 5.4180 2.4300 ;
      RECT 5.2840 1.3365 5.3100 2.4300 ;
      RECT 5.1760 1.3365 5.2020 2.4300 ;
      RECT 5.0680 1.3365 5.0940 2.4300 ;
      RECT 4.9600 1.3365 4.9860 2.4300 ;
      RECT 4.8520 1.3365 4.8780 2.4300 ;
      RECT 4.7440 1.3365 4.7700 2.4300 ;
      RECT 4.6360 1.3365 4.6620 2.4300 ;
      RECT 4.5280 1.3365 4.5540 2.4300 ;
      RECT 4.4200 1.3365 4.4460 2.4300 ;
      RECT 4.3120 1.3365 4.3380 2.4300 ;
      RECT 4.2040 1.3365 4.2300 2.4300 ;
      RECT 4.0960 1.3365 4.1220 2.4300 ;
      RECT 3.9880 1.3365 4.0140 2.4300 ;
      RECT 3.8800 1.3365 3.9060 2.4300 ;
      RECT 3.7720 1.3365 3.7980 2.4300 ;
      RECT 3.6640 1.3365 3.6900 2.4300 ;
      RECT 3.5560 1.3365 3.5820 2.4300 ;
      RECT 3.4480 1.3365 3.4740 2.4300 ;
      RECT 3.3400 1.3365 3.3660 2.4300 ;
      RECT 3.2320 1.3365 3.2580 2.4300 ;
      RECT 3.1240 1.3365 3.1500 2.4300 ;
      RECT 3.0160 1.3365 3.0420 2.4300 ;
      RECT 2.9080 1.3365 2.9340 2.4300 ;
      RECT 2.8000 1.3365 2.8260 2.4300 ;
      RECT 2.6920 1.3365 2.7180 2.4300 ;
      RECT 2.5840 1.3365 2.6100 2.4300 ;
      RECT 2.4760 1.3365 2.5020 2.4300 ;
      RECT 2.3680 1.3365 2.3940 2.4300 ;
      RECT 2.2600 1.3365 2.2860 2.4300 ;
      RECT 2.1520 1.3365 2.1780 2.4300 ;
      RECT 2.0440 1.3365 2.0700 2.4300 ;
      RECT 1.9360 1.3365 1.9620 2.4300 ;
      RECT 1.8280 1.3365 1.8540 2.4300 ;
      RECT 1.7200 1.3365 1.7460 2.4300 ;
      RECT 1.6120 1.3365 1.6380 2.4300 ;
      RECT 1.5040 1.3365 1.5300 2.4300 ;
      RECT 1.3960 1.3365 1.4220 2.4300 ;
      RECT 1.2880 1.3365 1.3140 2.4300 ;
      RECT 1.1800 1.3365 1.2060 2.4300 ;
      RECT 1.0720 1.3365 1.0980 2.4300 ;
      RECT 0.9640 1.3365 0.9900 2.4300 ;
      RECT 0.8560 1.3365 0.8820 2.4300 ;
      RECT 0.7480 1.3365 0.7740 2.4300 ;
      RECT 0.6400 1.3365 0.6660 2.4300 ;
      RECT 0.5320 1.3365 0.5580 2.4300 ;
      RECT 0.4240 1.3365 0.4500 2.4300 ;
      RECT 0.3160 1.3365 0.3420 2.4300 ;
      RECT 0.2080 1.3365 0.2340 2.4300 ;
      RECT 0.0050 1.3365 0.0900 2.4300 ;
      RECT 15.5530 2.4165 15.6810 3.5100 ;
      RECT 15.5390 3.0820 15.6810 3.4045 ;
      RECT 15.3190 2.8090 15.4530 3.5100 ;
      RECT 15.2960 3.1440 15.4530 3.4020 ;
      RECT 15.3190 2.4165 15.4170 3.5100 ;
      RECT 15.3190 2.5375 15.4310 2.7770 ;
      RECT 15.3190 2.4165 15.4530 2.5055 ;
      RECT 15.0940 2.8670 15.2280 3.5100 ;
      RECT 15.0940 2.4165 15.1920 3.5100 ;
      RECT 14.6770 2.4165 14.7600 3.5100 ;
      RECT 14.6770 2.5050 14.7740 3.4405 ;
      RECT 30.2680 2.4165 30.3530 3.5100 ;
      RECT 30.1240 2.4165 30.1500 3.5100 ;
      RECT 30.0160 2.4165 30.0420 3.5100 ;
      RECT 29.9080 2.4165 29.9340 3.5100 ;
      RECT 29.8000 2.4165 29.8260 3.5100 ;
      RECT 29.6920 2.4165 29.7180 3.5100 ;
      RECT 29.5840 2.4165 29.6100 3.5100 ;
      RECT 29.4760 2.4165 29.5020 3.5100 ;
      RECT 29.3680 2.4165 29.3940 3.5100 ;
      RECT 29.2600 2.4165 29.2860 3.5100 ;
      RECT 29.1520 2.4165 29.1780 3.5100 ;
      RECT 29.0440 2.4165 29.0700 3.5100 ;
      RECT 28.9360 2.4165 28.9620 3.5100 ;
      RECT 28.8280 2.4165 28.8540 3.5100 ;
      RECT 28.7200 2.4165 28.7460 3.5100 ;
      RECT 28.6120 2.4165 28.6380 3.5100 ;
      RECT 28.5040 2.4165 28.5300 3.5100 ;
      RECT 28.3960 2.4165 28.4220 3.5100 ;
      RECT 28.2880 2.4165 28.3140 3.5100 ;
      RECT 28.1800 2.4165 28.2060 3.5100 ;
      RECT 28.0720 2.4165 28.0980 3.5100 ;
      RECT 27.9640 2.4165 27.9900 3.5100 ;
      RECT 27.8560 2.4165 27.8820 3.5100 ;
      RECT 27.7480 2.4165 27.7740 3.5100 ;
      RECT 27.6400 2.4165 27.6660 3.5100 ;
      RECT 27.5320 2.4165 27.5580 3.5100 ;
      RECT 27.4240 2.4165 27.4500 3.5100 ;
      RECT 27.3160 2.4165 27.3420 3.5100 ;
      RECT 27.2080 2.4165 27.2340 3.5100 ;
      RECT 27.1000 2.4165 27.1260 3.5100 ;
      RECT 26.9920 2.4165 27.0180 3.5100 ;
      RECT 26.8840 2.4165 26.9100 3.5100 ;
      RECT 26.7760 2.4165 26.8020 3.5100 ;
      RECT 26.6680 2.4165 26.6940 3.5100 ;
      RECT 26.5600 2.4165 26.5860 3.5100 ;
      RECT 26.4520 2.4165 26.4780 3.5100 ;
      RECT 26.3440 2.4165 26.3700 3.5100 ;
      RECT 26.2360 2.4165 26.2620 3.5100 ;
      RECT 26.1280 2.4165 26.1540 3.5100 ;
      RECT 26.0200 2.4165 26.0460 3.5100 ;
      RECT 25.9120 2.4165 25.9380 3.5100 ;
      RECT 25.8040 2.4165 25.8300 3.5100 ;
      RECT 25.6960 2.4165 25.7220 3.5100 ;
      RECT 25.5880 2.4165 25.6140 3.5100 ;
      RECT 25.4800 2.4165 25.5060 3.5100 ;
      RECT 25.3720 2.4165 25.3980 3.5100 ;
      RECT 25.2640 2.4165 25.2900 3.5100 ;
      RECT 25.1560 2.4165 25.1820 3.5100 ;
      RECT 25.0480 2.4165 25.0740 3.5100 ;
      RECT 24.9400 2.4165 24.9660 3.5100 ;
      RECT 24.8320 2.4165 24.8580 3.5100 ;
      RECT 24.7240 2.4165 24.7500 3.5100 ;
      RECT 24.6160 2.4165 24.6420 3.5100 ;
      RECT 24.5080 2.4165 24.5340 3.5100 ;
      RECT 24.4000 2.4165 24.4260 3.5100 ;
      RECT 24.2920 2.4165 24.3180 3.5100 ;
      RECT 24.1840 2.4165 24.2100 3.5100 ;
      RECT 24.0760 2.4165 24.1020 3.5100 ;
      RECT 23.9680 2.4165 23.9940 3.5100 ;
      RECT 23.8600 2.4165 23.8860 3.5100 ;
      RECT 23.7520 2.4165 23.7780 3.5100 ;
      RECT 23.6440 2.4165 23.6700 3.5100 ;
      RECT 23.5360 2.4165 23.5620 3.5100 ;
      RECT 23.4280 2.4165 23.4540 3.5100 ;
      RECT 23.3200 2.4165 23.3460 3.5100 ;
      RECT 23.2120 2.4165 23.2380 3.5100 ;
      RECT 23.1040 2.4165 23.1300 3.5100 ;
      RECT 22.9960 2.4165 23.0220 3.5100 ;
      RECT 22.8880 2.4165 22.9140 3.5100 ;
      RECT 22.7800 2.4165 22.8060 3.5100 ;
      RECT 22.6720 2.4165 22.6980 3.5100 ;
      RECT 22.5640 2.4165 22.5900 3.5100 ;
      RECT 22.4560 2.4165 22.4820 3.5100 ;
      RECT 22.3480 2.4165 22.3740 3.5100 ;
      RECT 22.2400 2.4165 22.2660 3.5100 ;
      RECT 22.1320 2.4165 22.1580 3.5100 ;
      RECT 22.0240 2.4165 22.0500 3.5100 ;
      RECT 21.9160 2.4165 21.9420 3.5100 ;
      RECT 21.8080 2.4165 21.8340 3.5100 ;
      RECT 21.7000 2.4165 21.7260 3.5100 ;
      RECT 21.5920 2.4165 21.6180 3.5100 ;
      RECT 21.4840 2.4165 21.5100 3.5100 ;
      RECT 21.3760 2.4165 21.4020 3.5100 ;
      RECT 21.2680 2.4165 21.2940 3.5100 ;
      RECT 21.1600 2.4165 21.1860 3.5100 ;
      RECT 21.0520 2.4165 21.0780 3.5100 ;
      RECT 20.9440 2.4165 20.9700 3.5100 ;
      RECT 20.8360 2.4165 20.8620 3.5100 ;
      RECT 20.7280 2.4165 20.7540 3.5100 ;
      RECT 20.6200 2.4165 20.6460 3.5100 ;
      RECT 20.5120 2.4165 20.5380 3.5100 ;
      RECT 20.4040 2.4165 20.4300 3.5100 ;
      RECT 20.2960 2.4165 20.3220 3.5100 ;
      RECT 20.1880 2.4165 20.2140 3.5100 ;
      RECT 20.0800 2.4165 20.1060 3.5100 ;
      RECT 19.9720 2.4165 19.9980 3.5100 ;
      RECT 19.8640 2.4165 19.8900 3.5100 ;
      RECT 19.7560 2.4165 19.7820 3.5100 ;
      RECT 19.6480 2.4165 19.6740 3.5100 ;
      RECT 19.5400 2.4165 19.5660 3.5100 ;
      RECT 19.4320 2.4165 19.4580 3.5100 ;
      RECT 19.3240 2.4165 19.3500 3.5100 ;
      RECT 19.2160 2.4165 19.2420 3.5100 ;
      RECT 19.1080 2.4165 19.1340 3.5100 ;
      RECT 19.0000 2.4165 19.0260 3.5100 ;
      RECT 18.8920 2.4165 18.9180 3.5100 ;
      RECT 18.7840 2.4165 18.8100 3.5100 ;
      RECT 18.6760 2.4165 18.7020 3.5100 ;
      RECT 18.5680 2.4165 18.5940 3.5100 ;
      RECT 18.4600 2.4165 18.4860 3.5100 ;
      RECT 18.3520 2.4165 18.3780 3.5100 ;
      RECT 18.2440 2.4165 18.2700 3.5100 ;
      RECT 18.1360 2.4165 18.1620 3.5100 ;
      RECT 18.0280 2.4165 18.0540 3.5100 ;
      RECT 17.9200 2.4165 17.9460 3.5100 ;
      RECT 17.8120 2.4165 17.8380 3.5100 ;
      RECT 17.7040 2.4165 17.7300 3.5100 ;
      RECT 17.5960 2.4165 17.6220 3.5100 ;
      RECT 17.4880 2.4165 17.5140 3.5100 ;
      RECT 17.3800 2.4165 17.4060 3.5100 ;
      RECT 17.2720 2.4165 17.2980 3.5100 ;
      RECT 17.1640 2.4165 17.1900 3.5100 ;
      RECT 17.0560 2.4165 17.0820 3.5100 ;
      RECT 16.9480 2.4165 16.9740 3.5100 ;
      RECT 16.8400 2.4165 16.8660 3.5100 ;
      RECT 16.7320 2.4165 16.7580 3.5100 ;
      RECT 16.6240 2.4165 16.6500 3.5100 ;
      RECT 16.5160 2.4165 16.5420 3.5100 ;
      RECT 16.4080 2.4165 16.4340 3.5100 ;
      RECT 16.3000 2.4165 16.3260 3.5100 ;
      RECT 16.0870 2.4165 16.1640 3.5100 ;
      RECT 14.1940 2.4165 14.2710 3.5100 ;
      RECT 14.0320 2.4165 14.0580 3.5100 ;
      RECT 13.9240 2.4165 13.9500 3.5100 ;
      RECT 13.8160 2.4165 13.8420 3.5100 ;
      RECT 13.7080 2.4165 13.7340 3.5100 ;
      RECT 13.6000 2.4165 13.6260 3.5100 ;
      RECT 13.4920 2.4165 13.5180 3.5100 ;
      RECT 13.3840 2.4165 13.4100 3.5100 ;
      RECT 13.2760 2.4165 13.3020 3.5100 ;
      RECT 13.1680 2.4165 13.1940 3.5100 ;
      RECT 13.0600 2.4165 13.0860 3.5100 ;
      RECT 12.9520 2.4165 12.9780 3.5100 ;
      RECT 12.8440 2.4165 12.8700 3.5100 ;
      RECT 12.7360 2.4165 12.7620 3.5100 ;
      RECT 12.6280 2.4165 12.6540 3.5100 ;
      RECT 12.5200 2.4165 12.5460 3.5100 ;
      RECT 12.4120 2.4165 12.4380 3.5100 ;
      RECT 12.3040 2.4165 12.3300 3.5100 ;
      RECT 12.1960 2.4165 12.2220 3.5100 ;
      RECT 12.0880 2.4165 12.1140 3.5100 ;
      RECT 11.9800 2.4165 12.0060 3.5100 ;
      RECT 11.8720 2.4165 11.8980 3.5100 ;
      RECT 11.7640 2.4165 11.7900 3.5100 ;
      RECT 11.6560 2.4165 11.6820 3.5100 ;
      RECT 11.5480 2.4165 11.5740 3.5100 ;
      RECT 11.4400 2.4165 11.4660 3.5100 ;
      RECT 11.3320 2.4165 11.3580 3.5100 ;
      RECT 11.2240 2.4165 11.2500 3.5100 ;
      RECT 11.1160 2.4165 11.1420 3.5100 ;
      RECT 11.0080 2.4165 11.0340 3.5100 ;
      RECT 10.9000 2.4165 10.9260 3.5100 ;
      RECT 10.7920 2.4165 10.8180 3.5100 ;
      RECT 10.6840 2.4165 10.7100 3.5100 ;
      RECT 10.5760 2.4165 10.6020 3.5100 ;
      RECT 10.4680 2.4165 10.4940 3.5100 ;
      RECT 10.3600 2.4165 10.3860 3.5100 ;
      RECT 10.2520 2.4165 10.2780 3.5100 ;
      RECT 10.1440 2.4165 10.1700 3.5100 ;
      RECT 10.0360 2.4165 10.0620 3.5100 ;
      RECT 9.9280 2.4165 9.9540 3.5100 ;
      RECT 9.8200 2.4165 9.8460 3.5100 ;
      RECT 9.7120 2.4165 9.7380 3.5100 ;
      RECT 9.6040 2.4165 9.6300 3.5100 ;
      RECT 9.4960 2.4165 9.5220 3.5100 ;
      RECT 9.3880 2.4165 9.4140 3.5100 ;
      RECT 9.2800 2.4165 9.3060 3.5100 ;
      RECT 9.1720 2.4165 9.1980 3.5100 ;
      RECT 9.0640 2.4165 9.0900 3.5100 ;
      RECT 8.9560 2.4165 8.9820 3.5100 ;
      RECT 8.8480 2.4165 8.8740 3.5100 ;
      RECT 8.7400 2.4165 8.7660 3.5100 ;
      RECT 8.6320 2.4165 8.6580 3.5100 ;
      RECT 8.5240 2.4165 8.5500 3.5100 ;
      RECT 8.4160 2.4165 8.4420 3.5100 ;
      RECT 8.3080 2.4165 8.3340 3.5100 ;
      RECT 8.2000 2.4165 8.2260 3.5100 ;
      RECT 8.0920 2.4165 8.1180 3.5100 ;
      RECT 7.9840 2.4165 8.0100 3.5100 ;
      RECT 7.8760 2.4165 7.9020 3.5100 ;
      RECT 7.7680 2.4165 7.7940 3.5100 ;
      RECT 7.6600 2.4165 7.6860 3.5100 ;
      RECT 7.5520 2.4165 7.5780 3.5100 ;
      RECT 7.4440 2.4165 7.4700 3.5100 ;
      RECT 7.3360 2.4165 7.3620 3.5100 ;
      RECT 7.2280 2.4165 7.2540 3.5100 ;
      RECT 7.1200 2.4165 7.1460 3.5100 ;
      RECT 7.0120 2.4165 7.0380 3.5100 ;
      RECT 6.9040 2.4165 6.9300 3.5100 ;
      RECT 6.7960 2.4165 6.8220 3.5100 ;
      RECT 6.6880 2.4165 6.7140 3.5100 ;
      RECT 6.5800 2.4165 6.6060 3.5100 ;
      RECT 6.4720 2.4165 6.4980 3.5100 ;
      RECT 6.3640 2.4165 6.3900 3.5100 ;
      RECT 6.2560 2.4165 6.2820 3.5100 ;
      RECT 6.1480 2.4165 6.1740 3.5100 ;
      RECT 6.0400 2.4165 6.0660 3.5100 ;
      RECT 5.9320 2.4165 5.9580 3.5100 ;
      RECT 5.8240 2.4165 5.8500 3.5100 ;
      RECT 5.7160 2.4165 5.7420 3.5100 ;
      RECT 5.6080 2.4165 5.6340 3.5100 ;
      RECT 5.5000 2.4165 5.5260 3.5100 ;
      RECT 5.3920 2.4165 5.4180 3.5100 ;
      RECT 5.2840 2.4165 5.3100 3.5100 ;
      RECT 5.1760 2.4165 5.2020 3.5100 ;
      RECT 5.0680 2.4165 5.0940 3.5100 ;
      RECT 4.9600 2.4165 4.9860 3.5100 ;
      RECT 4.8520 2.4165 4.8780 3.5100 ;
      RECT 4.7440 2.4165 4.7700 3.5100 ;
      RECT 4.6360 2.4165 4.6620 3.5100 ;
      RECT 4.5280 2.4165 4.5540 3.5100 ;
      RECT 4.4200 2.4165 4.4460 3.5100 ;
      RECT 4.3120 2.4165 4.3380 3.5100 ;
      RECT 4.2040 2.4165 4.2300 3.5100 ;
      RECT 4.0960 2.4165 4.1220 3.5100 ;
      RECT 3.9880 2.4165 4.0140 3.5100 ;
      RECT 3.8800 2.4165 3.9060 3.5100 ;
      RECT 3.7720 2.4165 3.7980 3.5100 ;
      RECT 3.6640 2.4165 3.6900 3.5100 ;
      RECT 3.5560 2.4165 3.5820 3.5100 ;
      RECT 3.4480 2.4165 3.4740 3.5100 ;
      RECT 3.3400 2.4165 3.3660 3.5100 ;
      RECT 3.2320 2.4165 3.2580 3.5100 ;
      RECT 3.1240 2.4165 3.1500 3.5100 ;
      RECT 3.0160 2.4165 3.0420 3.5100 ;
      RECT 2.9080 2.4165 2.9340 3.5100 ;
      RECT 2.8000 2.4165 2.8260 3.5100 ;
      RECT 2.6920 2.4165 2.7180 3.5100 ;
      RECT 2.5840 2.4165 2.6100 3.5100 ;
      RECT 2.4760 2.4165 2.5020 3.5100 ;
      RECT 2.3680 2.4165 2.3940 3.5100 ;
      RECT 2.2600 2.4165 2.2860 3.5100 ;
      RECT 2.1520 2.4165 2.1780 3.5100 ;
      RECT 2.0440 2.4165 2.0700 3.5100 ;
      RECT 1.9360 2.4165 1.9620 3.5100 ;
      RECT 1.8280 2.4165 1.8540 3.5100 ;
      RECT 1.7200 2.4165 1.7460 3.5100 ;
      RECT 1.6120 2.4165 1.6380 3.5100 ;
      RECT 1.5040 2.4165 1.5300 3.5100 ;
      RECT 1.3960 2.4165 1.4220 3.5100 ;
      RECT 1.2880 2.4165 1.3140 3.5100 ;
      RECT 1.1800 2.4165 1.2060 3.5100 ;
      RECT 1.0720 2.4165 1.0980 3.5100 ;
      RECT 0.9640 2.4165 0.9900 3.5100 ;
      RECT 0.8560 2.4165 0.8820 3.5100 ;
      RECT 0.7480 2.4165 0.7740 3.5100 ;
      RECT 0.6400 2.4165 0.6660 3.5100 ;
      RECT 0.5320 2.4165 0.5580 3.5100 ;
      RECT 0.4240 2.4165 0.4500 3.5100 ;
      RECT 0.3160 2.4165 0.3420 3.5100 ;
      RECT 0.2080 2.4165 0.2340 3.5100 ;
      RECT 0.0050 2.4165 0.0900 3.5100 ;
      RECT 15.5530 3.4965 15.6810 4.5900 ;
      RECT 15.5390 4.1620 15.6810 4.4845 ;
      RECT 15.3190 3.8890 15.4530 4.5900 ;
      RECT 15.2960 4.2240 15.4530 4.4820 ;
      RECT 15.3190 3.4965 15.4170 4.5900 ;
      RECT 15.3190 3.6175 15.4310 3.8570 ;
      RECT 15.3190 3.4965 15.4530 3.5855 ;
      RECT 15.0940 3.9470 15.2280 4.5900 ;
      RECT 15.0940 3.4965 15.1920 4.5900 ;
      RECT 14.6770 3.4965 14.7600 4.5900 ;
      RECT 14.6770 3.5850 14.7740 4.5205 ;
      RECT 30.2680 3.4965 30.3530 4.5900 ;
      RECT 30.1240 3.4965 30.1500 4.5900 ;
      RECT 30.0160 3.4965 30.0420 4.5900 ;
      RECT 29.9080 3.4965 29.9340 4.5900 ;
      RECT 29.8000 3.4965 29.8260 4.5900 ;
      RECT 29.6920 3.4965 29.7180 4.5900 ;
      RECT 29.5840 3.4965 29.6100 4.5900 ;
      RECT 29.4760 3.4965 29.5020 4.5900 ;
      RECT 29.3680 3.4965 29.3940 4.5900 ;
      RECT 29.2600 3.4965 29.2860 4.5900 ;
      RECT 29.1520 3.4965 29.1780 4.5900 ;
      RECT 29.0440 3.4965 29.0700 4.5900 ;
      RECT 28.9360 3.4965 28.9620 4.5900 ;
      RECT 28.8280 3.4965 28.8540 4.5900 ;
      RECT 28.7200 3.4965 28.7460 4.5900 ;
      RECT 28.6120 3.4965 28.6380 4.5900 ;
      RECT 28.5040 3.4965 28.5300 4.5900 ;
      RECT 28.3960 3.4965 28.4220 4.5900 ;
      RECT 28.2880 3.4965 28.3140 4.5900 ;
      RECT 28.1800 3.4965 28.2060 4.5900 ;
      RECT 28.0720 3.4965 28.0980 4.5900 ;
      RECT 27.9640 3.4965 27.9900 4.5900 ;
      RECT 27.8560 3.4965 27.8820 4.5900 ;
      RECT 27.7480 3.4965 27.7740 4.5900 ;
      RECT 27.6400 3.4965 27.6660 4.5900 ;
      RECT 27.5320 3.4965 27.5580 4.5900 ;
      RECT 27.4240 3.4965 27.4500 4.5900 ;
      RECT 27.3160 3.4965 27.3420 4.5900 ;
      RECT 27.2080 3.4965 27.2340 4.5900 ;
      RECT 27.1000 3.4965 27.1260 4.5900 ;
      RECT 26.9920 3.4965 27.0180 4.5900 ;
      RECT 26.8840 3.4965 26.9100 4.5900 ;
      RECT 26.7760 3.4965 26.8020 4.5900 ;
      RECT 26.6680 3.4965 26.6940 4.5900 ;
      RECT 26.5600 3.4965 26.5860 4.5900 ;
      RECT 26.4520 3.4965 26.4780 4.5900 ;
      RECT 26.3440 3.4965 26.3700 4.5900 ;
      RECT 26.2360 3.4965 26.2620 4.5900 ;
      RECT 26.1280 3.4965 26.1540 4.5900 ;
      RECT 26.0200 3.4965 26.0460 4.5900 ;
      RECT 25.9120 3.4965 25.9380 4.5900 ;
      RECT 25.8040 3.4965 25.8300 4.5900 ;
      RECT 25.6960 3.4965 25.7220 4.5900 ;
      RECT 25.5880 3.4965 25.6140 4.5900 ;
      RECT 25.4800 3.4965 25.5060 4.5900 ;
      RECT 25.3720 3.4965 25.3980 4.5900 ;
      RECT 25.2640 3.4965 25.2900 4.5900 ;
      RECT 25.1560 3.4965 25.1820 4.5900 ;
      RECT 25.0480 3.4965 25.0740 4.5900 ;
      RECT 24.9400 3.4965 24.9660 4.5900 ;
      RECT 24.8320 3.4965 24.8580 4.5900 ;
      RECT 24.7240 3.4965 24.7500 4.5900 ;
      RECT 24.6160 3.4965 24.6420 4.5900 ;
      RECT 24.5080 3.4965 24.5340 4.5900 ;
      RECT 24.4000 3.4965 24.4260 4.5900 ;
      RECT 24.2920 3.4965 24.3180 4.5900 ;
      RECT 24.1840 3.4965 24.2100 4.5900 ;
      RECT 24.0760 3.4965 24.1020 4.5900 ;
      RECT 23.9680 3.4965 23.9940 4.5900 ;
      RECT 23.8600 3.4965 23.8860 4.5900 ;
      RECT 23.7520 3.4965 23.7780 4.5900 ;
      RECT 23.6440 3.4965 23.6700 4.5900 ;
      RECT 23.5360 3.4965 23.5620 4.5900 ;
      RECT 23.4280 3.4965 23.4540 4.5900 ;
      RECT 23.3200 3.4965 23.3460 4.5900 ;
      RECT 23.2120 3.4965 23.2380 4.5900 ;
      RECT 23.1040 3.4965 23.1300 4.5900 ;
      RECT 22.9960 3.4965 23.0220 4.5900 ;
      RECT 22.8880 3.4965 22.9140 4.5900 ;
      RECT 22.7800 3.4965 22.8060 4.5900 ;
      RECT 22.6720 3.4965 22.6980 4.5900 ;
      RECT 22.5640 3.4965 22.5900 4.5900 ;
      RECT 22.4560 3.4965 22.4820 4.5900 ;
      RECT 22.3480 3.4965 22.3740 4.5900 ;
      RECT 22.2400 3.4965 22.2660 4.5900 ;
      RECT 22.1320 3.4965 22.1580 4.5900 ;
      RECT 22.0240 3.4965 22.0500 4.5900 ;
      RECT 21.9160 3.4965 21.9420 4.5900 ;
      RECT 21.8080 3.4965 21.8340 4.5900 ;
      RECT 21.7000 3.4965 21.7260 4.5900 ;
      RECT 21.5920 3.4965 21.6180 4.5900 ;
      RECT 21.4840 3.4965 21.5100 4.5900 ;
      RECT 21.3760 3.4965 21.4020 4.5900 ;
      RECT 21.2680 3.4965 21.2940 4.5900 ;
      RECT 21.1600 3.4965 21.1860 4.5900 ;
      RECT 21.0520 3.4965 21.0780 4.5900 ;
      RECT 20.9440 3.4965 20.9700 4.5900 ;
      RECT 20.8360 3.4965 20.8620 4.5900 ;
      RECT 20.7280 3.4965 20.7540 4.5900 ;
      RECT 20.6200 3.4965 20.6460 4.5900 ;
      RECT 20.5120 3.4965 20.5380 4.5900 ;
      RECT 20.4040 3.4965 20.4300 4.5900 ;
      RECT 20.2960 3.4965 20.3220 4.5900 ;
      RECT 20.1880 3.4965 20.2140 4.5900 ;
      RECT 20.0800 3.4965 20.1060 4.5900 ;
      RECT 19.9720 3.4965 19.9980 4.5900 ;
      RECT 19.8640 3.4965 19.8900 4.5900 ;
      RECT 19.7560 3.4965 19.7820 4.5900 ;
      RECT 19.6480 3.4965 19.6740 4.5900 ;
      RECT 19.5400 3.4965 19.5660 4.5900 ;
      RECT 19.4320 3.4965 19.4580 4.5900 ;
      RECT 19.3240 3.4965 19.3500 4.5900 ;
      RECT 19.2160 3.4965 19.2420 4.5900 ;
      RECT 19.1080 3.4965 19.1340 4.5900 ;
      RECT 19.0000 3.4965 19.0260 4.5900 ;
      RECT 18.8920 3.4965 18.9180 4.5900 ;
      RECT 18.7840 3.4965 18.8100 4.5900 ;
      RECT 18.6760 3.4965 18.7020 4.5900 ;
      RECT 18.5680 3.4965 18.5940 4.5900 ;
      RECT 18.4600 3.4965 18.4860 4.5900 ;
      RECT 18.3520 3.4965 18.3780 4.5900 ;
      RECT 18.2440 3.4965 18.2700 4.5900 ;
      RECT 18.1360 3.4965 18.1620 4.5900 ;
      RECT 18.0280 3.4965 18.0540 4.5900 ;
      RECT 17.9200 3.4965 17.9460 4.5900 ;
      RECT 17.8120 3.4965 17.8380 4.5900 ;
      RECT 17.7040 3.4965 17.7300 4.5900 ;
      RECT 17.5960 3.4965 17.6220 4.5900 ;
      RECT 17.4880 3.4965 17.5140 4.5900 ;
      RECT 17.3800 3.4965 17.4060 4.5900 ;
      RECT 17.2720 3.4965 17.2980 4.5900 ;
      RECT 17.1640 3.4965 17.1900 4.5900 ;
      RECT 17.0560 3.4965 17.0820 4.5900 ;
      RECT 16.9480 3.4965 16.9740 4.5900 ;
      RECT 16.8400 3.4965 16.8660 4.5900 ;
      RECT 16.7320 3.4965 16.7580 4.5900 ;
      RECT 16.6240 3.4965 16.6500 4.5900 ;
      RECT 16.5160 3.4965 16.5420 4.5900 ;
      RECT 16.4080 3.4965 16.4340 4.5900 ;
      RECT 16.3000 3.4965 16.3260 4.5900 ;
      RECT 16.0870 3.4965 16.1640 4.5900 ;
      RECT 14.1940 3.4965 14.2710 4.5900 ;
      RECT 14.0320 3.4965 14.0580 4.5900 ;
      RECT 13.9240 3.4965 13.9500 4.5900 ;
      RECT 13.8160 3.4965 13.8420 4.5900 ;
      RECT 13.7080 3.4965 13.7340 4.5900 ;
      RECT 13.6000 3.4965 13.6260 4.5900 ;
      RECT 13.4920 3.4965 13.5180 4.5900 ;
      RECT 13.3840 3.4965 13.4100 4.5900 ;
      RECT 13.2760 3.4965 13.3020 4.5900 ;
      RECT 13.1680 3.4965 13.1940 4.5900 ;
      RECT 13.0600 3.4965 13.0860 4.5900 ;
      RECT 12.9520 3.4965 12.9780 4.5900 ;
      RECT 12.8440 3.4965 12.8700 4.5900 ;
      RECT 12.7360 3.4965 12.7620 4.5900 ;
      RECT 12.6280 3.4965 12.6540 4.5900 ;
      RECT 12.5200 3.4965 12.5460 4.5900 ;
      RECT 12.4120 3.4965 12.4380 4.5900 ;
      RECT 12.3040 3.4965 12.3300 4.5900 ;
      RECT 12.1960 3.4965 12.2220 4.5900 ;
      RECT 12.0880 3.4965 12.1140 4.5900 ;
      RECT 11.9800 3.4965 12.0060 4.5900 ;
      RECT 11.8720 3.4965 11.8980 4.5900 ;
      RECT 11.7640 3.4965 11.7900 4.5900 ;
      RECT 11.6560 3.4965 11.6820 4.5900 ;
      RECT 11.5480 3.4965 11.5740 4.5900 ;
      RECT 11.4400 3.4965 11.4660 4.5900 ;
      RECT 11.3320 3.4965 11.3580 4.5900 ;
      RECT 11.2240 3.4965 11.2500 4.5900 ;
      RECT 11.1160 3.4965 11.1420 4.5900 ;
      RECT 11.0080 3.4965 11.0340 4.5900 ;
      RECT 10.9000 3.4965 10.9260 4.5900 ;
      RECT 10.7920 3.4965 10.8180 4.5900 ;
      RECT 10.6840 3.4965 10.7100 4.5900 ;
      RECT 10.5760 3.4965 10.6020 4.5900 ;
      RECT 10.4680 3.4965 10.4940 4.5900 ;
      RECT 10.3600 3.4965 10.3860 4.5900 ;
      RECT 10.2520 3.4965 10.2780 4.5900 ;
      RECT 10.1440 3.4965 10.1700 4.5900 ;
      RECT 10.0360 3.4965 10.0620 4.5900 ;
      RECT 9.9280 3.4965 9.9540 4.5900 ;
      RECT 9.8200 3.4965 9.8460 4.5900 ;
      RECT 9.7120 3.4965 9.7380 4.5900 ;
      RECT 9.6040 3.4965 9.6300 4.5900 ;
      RECT 9.4960 3.4965 9.5220 4.5900 ;
      RECT 9.3880 3.4965 9.4140 4.5900 ;
      RECT 9.2800 3.4965 9.3060 4.5900 ;
      RECT 9.1720 3.4965 9.1980 4.5900 ;
      RECT 9.0640 3.4965 9.0900 4.5900 ;
      RECT 8.9560 3.4965 8.9820 4.5900 ;
      RECT 8.8480 3.4965 8.8740 4.5900 ;
      RECT 8.7400 3.4965 8.7660 4.5900 ;
      RECT 8.6320 3.4965 8.6580 4.5900 ;
      RECT 8.5240 3.4965 8.5500 4.5900 ;
      RECT 8.4160 3.4965 8.4420 4.5900 ;
      RECT 8.3080 3.4965 8.3340 4.5900 ;
      RECT 8.2000 3.4965 8.2260 4.5900 ;
      RECT 8.0920 3.4965 8.1180 4.5900 ;
      RECT 7.9840 3.4965 8.0100 4.5900 ;
      RECT 7.8760 3.4965 7.9020 4.5900 ;
      RECT 7.7680 3.4965 7.7940 4.5900 ;
      RECT 7.6600 3.4965 7.6860 4.5900 ;
      RECT 7.5520 3.4965 7.5780 4.5900 ;
      RECT 7.4440 3.4965 7.4700 4.5900 ;
      RECT 7.3360 3.4965 7.3620 4.5900 ;
      RECT 7.2280 3.4965 7.2540 4.5900 ;
      RECT 7.1200 3.4965 7.1460 4.5900 ;
      RECT 7.0120 3.4965 7.0380 4.5900 ;
      RECT 6.9040 3.4965 6.9300 4.5900 ;
      RECT 6.7960 3.4965 6.8220 4.5900 ;
      RECT 6.6880 3.4965 6.7140 4.5900 ;
      RECT 6.5800 3.4965 6.6060 4.5900 ;
      RECT 6.4720 3.4965 6.4980 4.5900 ;
      RECT 6.3640 3.4965 6.3900 4.5900 ;
      RECT 6.2560 3.4965 6.2820 4.5900 ;
      RECT 6.1480 3.4965 6.1740 4.5900 ;
      RECT 6.0400 3.4965 6.0660 4.5900 ;
      RECT 5.9320 3.4965 5.9580 4.5900 ;
      RECT 5.8240 3.4965 5.8500 4.5900 ;
      RECT 5.7160 3.4965 5.7420 4.5900 ;
      RECT 5.6080 3.4965 5.6340 4.5900 ;
      RECT 5.5000 3.4965 5.5260 4.5900 ;
      RECT 5.3920 3.4965 5.4180 4.5900 ;
      RECT 5.2840 3.4965 5.3100 4.5900 ;
      RECT 5.1760 3.4965 5.2020 4.5900 ;
      RECT 5.0680 3.4965 5.0940 4.5900 ;
      RECT 4.9600 3.4965 4.9860 4.5900 ;
      RECT 4.8520 3.4965 4.8780 4.5900 ;
      RECT 4.7440 3.4965 4.7700 4.5900 ;
      RECT 4.6360 3.4965 4.6620 4.5900 ;
      RECT 4.5280 3.4965 4.5540 4.5900 ;
      RECT 4.4200 3.4965 4.4460 4.5900 ;
      RECT 4.3120 3.4965 4.3380 4.5900 ;
      RECT 4.2040 3.4965 4.2300 4.5900 ;
      RECT 4.0960 3.4965 4.1220 4.5900 ;
      RECT 3.9880 3.4965 4.0140 4.5900 ;
      RECT 3.8800 3.4965 3.9060 4.5900 ;
      RECT 3.7720 3.4965 3.7980 4.5900 ;
      RECT 3.6640 3.4965 3.6900 4.5900 ;
      RECT 3.5560 3.4965 3.5820 4.5900 ;
      RECT 3.4480 3.4965 3.4740 4.5900 ;
      RECT 3.3400 3.4965 3.3660 4.5900 ;
      RECT 3.2320 3.4965 3.2580 4.5900 ;
      RECT 3.1240 3.4965 3.1500 4.5900 ;
      RECT 3.0160 3.4965 3.0420 4.5900 ;
      RECT 2.9080 3.4965 2.9340 4.5900 ;
      RECT 2.8000 3.4965 2.8260 4.5900 ;
      RECT 2.6920 3.4965 2.7180 4.5900 ;
      RECT 2.5840 3.4965 2.6100 4.5900 ;
      RECT 2.4760 3.4965 2.5020 4.5900 ;
      RECT 2.3680 3.4965 2.3940 4.5900 ;
      RECT 2.2600 3.4965 2.2860 4.5900 ;
      RECT 2.1520 3.4965 2.1780 4.5900 ;
      RECT 2.0440 3.4965 2.0700 4.5900 ;
      RECT 1.9360 3.4965 1.9620 4.5900 ;
      RECT 1.8280 3.4965 1.8540 4.5900 ;
      RECT 1.7200 3.4965 1.7460 4.5900 ;
      RECT 1.6120 3.4965 1.6380 4.5900 ;
      RECT 1.5040 3.4965 1.5300 4.5900 ;
      RECT 1.3960 3.4965 1.4220 4.5900 ;
      RECT 1.2880 3.4965 1.3140 4.5900 ;
      RECT 1.1800 3.4965 1.2060 4.5900 ;
      RECT 1.0720 3.4965 1.0980 4.5900 ;
      RECT 0.9640 3.4965 0.9900 4.5900 ;
      RECT 0.8560 3.4965 0.8820 4.5900 ;
      RECT 0.7480 3.4965 0.7740 4.5900 ;
      RECT 0.6400 3.4965 0.6660 4.5900 ;
      RECT 0.5320 3.4965 0.5580 4.5900 ;
      RECT 0.4240 3.4965 0.4500 4.5900 ;
      RECT 0.3160 3.4965 0.3420 4.5900 ;
      RECT 0.2080 3.4965 0.2340 4.5900 ;
      RECT 0.0050 3.4965 0.0900 4.5900 ;
      RECT 15.5530 4.5765 15.6810 5.6700 ;
      RECT 15.5390 5.2420 15.6810 5.5645 ;
      RECT 15.3190 4.9690 15.4530 5.6700 ;
      RECT 15.2960 5.3040 15.4530 5.5620 ;
      RECT 15.3190 4.5765 15.4170 5.6700 ;
      RECT 15.3190 4.6975 15.4310 4.9370 ;
      RECT 15.3190 4.5765 15.4530 4.6655 ;
      RECT 15.0940 5.0270 15.2280 5.6700 ;
      RECT 15.0940 4.5765 15.1920 5.6700 ;
      RECT 14.6770 4.5765 14.7600 5.6700 ;
      RECT 14.6770 4.6650 14.7740 5.6005 ;
      RECT 30.2680 4.5765 30.3530 5.6700 ;
      RECT 30.1240 4.5765 30.1500 5.6700 ;
      RECT 30.0160 4.5765 30.0420 5.6700 ;
      RECT 29.9080 4.5765 29.9340 5.6700 ;
      RECT 29.8000 4.5765 29.8260 5.6700 ;
      RECT 29.6920 4.5765 29.7180 5.6700 ;
      RECT 29.5840 4.5765 29.6100 5.6700 ;
      RECT 29.4760 4.5765 29.5020 5.6700 ;
      RECT 29.3680 4.5765 29.3940 5.6700 ;
      RECT 29.2600 4.5765 29.2860 5.6700 ;
      RECT 29.1520 4.5765 29.1780 5.6700 ;
      RECT 29.0440 4.5765 29.0700 5.6700 ;
      RECT 28.9360 4.5765 28.9620 5.6700 ;
      RECT 28.8280 4.5765 28.8540 5.6700 ;
      RECT 28.7200 4.5765 28.7460 5.6700 ;
      RECT 28.6120 4.5765 28.6380 5.6700 ;
      RECT 28.5040 4.5765 28.5300 5.6700 ;
      RECT 28.3960 4.5765 28.4220 5.6700 ;
      RECT 28.2880 4.5765 28.3140 5.6700 ;
      RECT 28.1800 4.5765 28.2060 5.6700 ;
      RECT 28.0720 4.5765 28.0980 5.6700 ;
      RECT 27.9640 4.5765 27.9900 5.6700 ;
      RECT 27.8560 4.5765 27.8820 5.6700 ;
      RECT 27.7480 4.5765 27.7740 5.6700 ;
      RECT 27.6400 4.5765 27.6660 5.6700 ;
      RECT 27.5320 4.5765 27.5580 5.6700 ;
      RECT 27.4240 4.5765 27.4500 5.6700 ;
      RECT 27.3160 4.5765 27.3420 5.6700 ;
      RECT 27.2080 4.5765 27.2340 5.6700 ;
      RECT 27.1000 4.5765 27.1260 5.6700 ;
      RECT 26.9920 4.5765 27.0180 5.6700 ;
      RECT 26.8840 4.5765 26.9100 5.6700 ;
      RECT 26.7760 4.5765 26.8020 5.6700 ;
      RECT 26.6680 4.5765 26.6940 5.6700 ;
      RECT 26.5600 4.5765 26.5860 5.6700 ;
      RECT 26.4520 4.5765 26.4780 5.6700 ;
      RECT 26.3440 4.5765 26.3700 5.6700 ;
      RECT 26.2360 4.5765 26.2620 5.6700 ;
      RECT 26.1280 4.5765 26.1540 5.6700 ;
      RECT 26.0200 4.5765 26.0460 5.6700 ;
      RECT 25.9120 4.5765 25.9380 5.6700 ;
      RECT 25.8040 4.5765 25.8300 5.6700 ;
      RECT 25.6960 4.5765 25.7220 5.6700 ;
      RECT 25.5880 4.5765 25.6140 5.6700 ;
      RECT 25.4800 4.5765 25.5060 5.6700 ;
      RECT 25.3720 4.5765 25.3980 5.6700 ;
      RECT 25.2640 4.5765 25.2900 5.6700 ;
      RECT 25.1560 4.5765 25.1820 5.6700 ;
      RECT 25.0480 4.5765 25.0740 5.6700 ;
      RECT 24.9400 4.5765 24.9660 5.6700 ;
      RECT 24.8320 4.5765 24.8580 5.6700 ;
      RECT 24.7240 4.5765 24.7500 5.6700 ;
      RECT 24.6160 4.5765 24.6420 5.6700 ;
      RECT 24.5080 4.5765 24.5340 5.6700 ;
      RECT 24.4000 4.5765 24.4260 5.6700 ;
      RECT 24.2920 4.5765 24.3180 5.6700 ;
      RECT 24.1840 4.5765 24.2100 5.6700 ;
      RECT 24.0760 4.5765 24.1020 5.6700 ;
      RECT 23.9680 4.5765 23.9940 5.6700 ;
      RECT 23.8600 4.5765 23.8860 5.6700 ;
      RECT 23.7520 4.5765 23.7780 5.6700 ;
      RECT 23.6440 4.5765 23.6700 5.6700 ;
      RECT 23.5360 4.5765 23.5620 5.6700 ;
      RECT 23.4280 4.5765 23.4540 5.6700 ;
      RECT 23.3200 4.5765 23.3460 5.6700 ;
      RECT 23.2120 4.5765 23.2380 5.6700 ;
      RECT 23.1040 4.5765 23.1300 5.6700 ;
      RECT 22.9960 4.5765 23.0220 5.6700 ;
      RECT 22.8880 4.5765 22.9140 5.6700 ;
      RECT 22.7800 4.5765 22.8060 5.6700 ;
      RECT 22.6720 4.5765 22.6980 5.6700 ;
      RECT 22.5640 4.5765 22.5900 5.6700 ;
      RECT 22.4560 4.5765 22.4820 5.6700 ;
      RECT 22.3480 4.5765 22.3740 5.6700 ;
      RECT 22.2400 4.5765 22.2660 5.6700 ;
      RECT 22.1320 4.5765 22.1580 5.6700 ;
      RECT 22.0240 4.5765 22.0500 5.6700 ;
      RECT 21.9160 4.5765 21.9420 5.6700 ;
      RECT 21.8080 4.5765 21.8340 5.6700 ;
      RECT 21.7000 4.5765 21.7260 5.6700 ;
      RECT 21.5920 4.5765 21.6180 5.6700 ;
      RECT 21.4840 4.5765 21.5100 5.6700 ;
      RECT 21.3760 4.5765 21.4020 5.6700 ;
      RECT 21.2680 4.5765 21.2940 5.6700 ;
      RECT 21.1600 4.5765 21.1860 5.6700 ;
      RECT 21.0520 4.5765 21.0780 5.6700 ;
      RECT 20.9440 4.5765 20.9700 5.6700 ;
      RECT 20.8360 4.5765 20.8620 5.6700 ;
      RECT 20.7280 4.5765 20.7540 5.6700 ;
      RECT 20.6200 4.5765 20.6460 5.6700 ;
      RECT 20.5120 4.5765 20.5380 5.6700 ;
      RECT 20.4040 4.5765 20.4300 5.6700 ;
      RECT 20.2960 4.5765 20.3220 5.6700 ;
      RECT 20.1880 4.5765 20.2140 5.6700 ;
      RECT 20.0800 4.5765 20.1060 5.6700 ;
      RECT 19.9720 4.5765 19.9980 5.6700 ;
      RECT 19.8640 4.5765 19.8900 5.6700 ;
      RECT 19.7560 4.5765 19.7820 5.6700 ;
      RECT 19.6480 4.5765 19.6740 5.6700 ;
      RECT 19.5400 4.5765 19.5660 5.6700 ;
      RECT 19.4320 4.5765 19.4580 5.6700 ;
      RECT 19.3240 4.5765 19.3500 5.6700 ;
      RECT 19.2160 4.5765 19.2420 5.6700 ;
      RECT 19.1080 4.5765 19.1340 5.6700 ;
      RECT 19.0000 4.5765 19.0260 5.6700 ;
      RECT 18.8920 4.5765 18.9180 5.6700 ;
      RECT 18.7840 4.5765 18.8100 5.6700 ;
      RECT 18.6760 4.5765 18.7020 5.6700 ;
      RECT 18.5680 4.5765 18.5940 5.6700 ;
      RECT 18.4600 4.5765 18.4860 5.6700 ;
      RECT 18.3520 4.5765 18.3780 5.6700 ;
      RECT 18.2440 4.5765 18.2700 5.6700 ;
      RECT 18.1360 4.5765 18.1620 5.6700 ;
      RECT 18.0280 4.5765 18.0540 5.6700 ;
      RECT 17.9200 4.5765 17.9460 5.6700 ;
      RECT 17.8120 4.5765 17.8380 5.6700 ;
      RECT 17.7040 4.5765 17.7300 5.6700 ;
      RECT 17.5960 4.5765 17.6220 5.6700 ;
      RECT 17.4880 4.5765 17.5140 5.6700 ;
      RECT 17.3800 4.5765 17.4060 5.6700 ;
      RECT 17.2720 4.5765 17.2980 5.6700 ;
      RECT 17.1640 4.5765 17.1900 5.6700 ;
      RECT 17.0560 4.5765 17.0820 5.6700 ;
      RECT 16.9480 4.5765 16.9740 5.6700 ;
      RECT 16.8400 4.5765 16.8660 5.6700 ;
      RECT 16.7320 4.5765 16.7580 5.6700 ;
      RECT 16.6240 4.5765 16.6500 5.6700 ;
      RECT 16.5160 4.5765 16.5420 5.6700 ;
      RECT 16.4080 4.5765 16.4340 5.6700 ;
      RECT 16.3000 4.5765 16.3260 5.6700 ;
      RECT 16.0870 4.5765 16.1640 5.6700 ;
      RECT 14.1940 4.5765 14.2710 5.6700 ;
      RECT 14.0320 4.5765 14.0580 5.6700 ;
      RECT 13.9240 4.5765 13.9500 5.6700 ;
      RECT 13.8160 4.5765 13.8420 5.6700 ;
      RECT 13.7080 4.5765 13.7340 5.6700 ;
      RECT 13.6000 4.5765 13.6260 5.6700 ;
      RECT 13.4920 4.5765 13.5180 5.6700 ;
      RECT 13.3840 4.5765 13.4100 5.6700 ;
      RECT 13.2760 4.5765 13.3020 5.6700 ;
      RECT 13.1680 4.5765 13.1940 5.6700 ;
      RECT 13.0600 4.5765 13.0860 5.6700 ;
      RECT 12.9520 4.5765 12.9780 5.6700 ;
      RECT 12.8440 4.5765 12.8700 5.6700 ;
      RECT 12.7360 4.5765 12.7620 5.6700 ;
      RECT 12.6280 4.5765 12.6540 5.6700 ;
      RECT 12.5200 4.5765 12.5460 5.6700 ;
      RECT 12.4120 4.5765 12.4380 5.6700 ;
      RECT 12.3040 4.5765 12.3300 5.6700 ;
      RECT 12.1960 4.5765 12.2220 5.6700 ;
      RECT 12.0880 4.5765 12.1140 5.6700 ;
      RECT 11.9800 4.5765 12.0060 5.6700 ;
      RECT 11.8720 4.5765 11.8980 5.6700 ;
      RECT 11.7640 4.5765 11.7900 5.6700 ;
      RECT 11.6560 4.5765 11.6820 5.6700 ;
      RECT 11.5480 4.5765 11.5740 5.6700 ;
      RECT 11.4400 4.5765 11.4660 5.6700 ;
      RECT 11.3320 4.5765 11.3580 5.6700 ;
      RECT 11.2240 4.5765 11.2500 5.6700 ;
      RECT 11.1160 4.5765 11.1420 5.6700 ;
      RECT 11.0080 4.5765 11.0340 5.6700 ;
      RECT 10.9000 4.5765 10.9260 5.6700 ;
      RECT 10.7920 4.5765 10.8180 5.6700 ;
      RECT 10.6840 4.5765 10.7100 5.6700 ;
      RECT 10.5760 4.5765 10.6020 5.6700 ;
      RECT 10.4680 4.5765 10.4940 5.6700 ;
      RECT 10.3600 4.5765 10.3860 5.6700 ;
      RECT 10.2520 4.5765 10.2780 5.6700 ;
      RECT 10.1440 4.5765 10.1700 5.6700 ;
      RECT 10.0360 4.5765 10.0620 5.6700 ;
      RECT 9.9280 4.5765 9.9540 5.6700 ;
      RECT 9.8200 4.5765 9.8460 5.6700 ;
      RECT 9.7120 4.5765 9.7380 5.6700 ;
      RECT 9.6040 4.5765 9.6300 5.6700 ;
      RECT 9.4960 4.5765 9.5220 5.6700 ;
      RECT 9.3880 4.5765 9.4140 5.6700 ;
      RECT 9.2800 4.5765 9.3060 5.6700 ;
      RECT 9.1720 4.5765 9.1980 5.6700 ;
      RECT 9.0640 4.5765 9.0900 5.6700 ;
      RECT 8.9560 4.5765 8.9820 5.6700 ;
      RECT 8.8480 4.5765 8.8740 5.6700 ;
      RECT 8.7400 4.5765 8.7660 5.6700 ;
      RECT 8.6320 4.5765 8.6580 5.6700 ;
      RECT 8.5240 4.5765 8.5500 5.6700 ;
      RECT 8.4160 4.5765 8.4420 5.6700 ;
      RECT 8.3080 4.5765 8.3340 5.6700 ;
      RECT 8.2000 4.5765 8.2260 5.6700 ;
      RECT 8.0920 4.5765 8.1180 5.6700 ;
      RECT 7.9840 4.5765 8.0100 5.6700 ;
      RECT 7.8760 4.5765 7.9020 5.6700 ;
      RECT 7.7680 4.5765 7.7940 5.6700 ;
      RECT 7.6600 4.5765 7.6860 5.6700 ;
      RECT 7.5520 4.5765 7.5780 5.6700 ;
      RECT 7.4440 4.5765 7.4700 5.6700 ;
      RECT 7.3360 4.5765 7.3620 5.6700 ;
      RECT 7.2280 4.5765 7.2540 5.6700 ;
      RECT 7.1200 4.5765 7.1460 5.6700 ;
      RECT 7.0120 4.5765 7.0380 5.6700 ;
      RECT 6.9040 4.5765 6.9300 5.6700 ;
      RECT 6.7960 4.5765 6.8220 5.6700 ;
      RECT 6.6880 4.5765 6.7140 5.6700 ;
      RECT 6.5800 4.5765 6.6060 5.6700 ;
      RECT 6.4720 4.5765 6.4980 5.6700 ;
      RECT 6.3640 4.5765 6.3900 5.6700 ;
      RECT 6.2560 4.5765 6.2820 5.6700 ;
      RECT 6.1480 4.5765 6.1740 5.6700 ;
      RECT 6.0400 4.5765 6.0660 5.6700 ;
      RECT 5.9320 4.5765 5.9580 5.6700 ;
      RECT 5.8240 4.5765 5.8500 5.6700 ;
      RECT 5.7160 4.5765 5.7420 5.6700 ;
      RECT 5.6080 4.5765 5.6340 5.6700 ;
      RECT 5.5000 4.5765 5.5260 5.6700 ;
      RECT 5.3920 4.5765 5.4180 5.6700 ;
      RECT 5.2840 4.5765 5.3100 5.6700 ;
      RECT 5.1760 4.5765 5.2020 5.6700 ;
      RECT 5.0680 4.5765 5.0940 5.6700 ;
      RECT 4.9600 4.5765 4.9860 5.6700 ;
      RECT 4.8520 4.5765 4.8780 5.6700 ;
      RECT 4.7440 4.5765 4.7700 5.6700 ;
      RECT 4.6360 4.5765 4.6620 5.6700 ;
      RECT 4.5280 4.5765 4.5540 5.6700 ;
      RECT 4.4200 4.5765 4.4460 5.6700 ;
      RECT 4.3120 4.5765 4.3380 5.6700 ;
      RECT 4.2040 4.5765 4.2300 5.6700 ;
      RECT 4.0960 4.5765 4.1220 5.6700 ;
      RECT 3.9880 4.5765 4.0140 5.6700 ;
      RECT 3.8800 4.5765 3.9060 5.6700 ;
      RECT 3.7720 4.5765 3.7980 5.6700 ;
      RECT 3.6640 4.5765 3.6900 5.6700 ;
      RECT 3.5560 4.5765 3.5820 5.6700 ;
      RECT 3.4480 4.5765 3.4740 5.6700 ;
      RECT 3.3400 4.5765 3.3660 5.6700 ;
      RECT 3.2320 4.5765 3.2580 5.6700 ;
      RECT 3.1240 4.5765 3.1500 5.6700 ;
      RECT 3.0160 4.5765 3.0420 5.6700 ;
      RECT 2.9080 4.5765 2.9340 5.6700 ;
      RECT 2.8000 4.5765 2.8260 5.6700 ;
      RECT 2.6920 4.5765 2.7180 5.6700 ;
      RECT 2.5840 4.5765 2.6100 5.6700 ;
      RECT 2.4760 4.5765 2.5020 5.6700 ;
      RECT 2.3680 4.5765 2.3940 5.6700 ;
      RECT 2.2600 4.5765 2.2860 5.6700 ;
      RECT 2.1520 4.5765 2.1780 5.6700 ;
      RECT 2.0440 4.5765 2.0700 5.6700 ;
      RECT 1.9360 4.5765 1.9620 5.6700 ;
      RECT 1.8280 4.5765 1.8540 5.6700 ;
      RECT 1.7200 4.5765 1.7460 5.6700 ;
      RECT 1.6120 4.5765 1.6380 5.6700 ;
      RECT 1.5040 4.5765 1.5300 5.6700 ;
      RECT 1.3960 4.5765 1.4220 5.6700 ;
      RECT 1.2880 4.5765 1.3140 5.6700 ;
      RECT 1.1800 4.5765 1.2060 5.6700 ;
      RECT 1.0720 4.5765 1.0980 5.6700 ;
      RECT 0.9640 4.5765 0.9900 5.6700 ;
      RECT 0.8560 4.5765 0.8820 5.6700 ;
      RECT 0.7480 4.5765 0.7740 5.6700 ;
      RECT 0.6400 4.5765 0.6660 5.6700 ;
      RECT 0.5320 4.5765 0.5580 5.6700 ;
      RECT 0.4240 4.5765 0.4500 5.6700 ;
      RECT 0.3160 4.5765 0.3420 5.6700 ;
      RECT 0.2080 4.5765 0.2340 5.6700 ;
      RECT 0.0050 4.5765 0.0900 5.6700 ;
      RECT 15.5530 5.6565 15.6810 6.7500 ;
      RECT 15.5390 6.3220 15.6810 6.6445 ;
      RECT 15.3190 6.0490 15.4530 6.7500 ;
      RECT 15.2960 6.3840 15.4530 6.6420 ;
      RECT 15.3190 5.6565 15.4170 6.7500 ;
      RECT 15.3190 5.7775 15.4310 6.0170 ;
      RECT 15.3190 5.6565 15.4530 5.7455 ;
      RECT 15.0940 6.1070 15.2280 6.7500 ;
      RECT 15.0940 5.6565 15.1920 6.7500 ;
      RECT 14.6770 5.6565 14.7600 6.7500 ;
      RECT 14.6770 5.7450 14.7740 6.6805 ;
      RECT 30.2680 5.6565 30.3530 6.7500 ;
      RECT 30.1240 5.6565 30.1500 6.7500 ;
      RECT 30.0160 5.6565 30.0420 6.7500 ;
      RECT 29.9080 5.6565 29.9340 6.7500 ;
      RECT 29.8000 5.6565 29.8260 6.7500 ;
      RECT 29.6920 5.6565 29.7180 6.7500 ;
      RECT 29.5840 5.6565 29.6100 6.7500 ;
      RECT 29.4760 5.6565 29.5020 6.7500 ;
      RECT 29.3680 5.6565 29.3940 6.7500 ;
      RECT 29.2600 5.6565 29.2860 6.7500 ;
      RECT 29.1520 5.6565 29.1780 6.7500 ;
      RECT 29.0440 5.6565 29.0700 6.7500 ;
      RECT 28.9360 5.6565 28.9620 6.7500 ;
      RECT 28.8280 5.6565 28.8540 6.7500 ;
      RECT 28.7200 5.6565 28.7460 6.7500 ;
      RECT 28.6120 5.6565 28.6380 6.7500 ;
      RECT 28.5040 5.6565 28.5300 6.7500 ;
      RECT 28.3960 5.6565 28.4220 6.7500 ;
      RECT 28.2880 5.6565 28.3140 6.7500 ;
      RECT 28.1800 5.6565 28.2060 6.7500 ;
      RECT 28.0720 5.6565 28.0980 6.7500 ;
      RECT 27.9640 5.6565 27.9900 6.7500 ;
      RECT 27.8560 5.6565 27.8820 6.7500 ;
      RECT 27.7480 5.6565 27.7740 6.7500 ;
      RECT 27.6400 5.6565 27.6660 6.7500 ;
      RECT 27.5320 5.6565 27.5580 6.7500 ;
      RECT 27.4240 5.6565 27.4500 6.7500 ;
      RECT 27.3160 5.6565 27.3420 6.7500 ;
      RECT 27.2080 5.6565 27.2340 6.7500 ;
      RECT 27.1000 5.6565 27.1260 6.7500 ;
      RECT 26.9920 5.6565 27.0180 6.7500 ;
      RECT 26.8840 5.6565 26.9100 6.7500 ;
      RECT 26.7760 5.6565 26.8020 6.7500 ;
      RECT 26.6680 5.6565 26.6940 6.7500 ;
      RECT 26.5600 5.6565 26.5860 6.7500 ;
      RECT 26.4520 5.6565 26.4780 6.7500 ;
      RECT 26.3440 5.6565 26.3700 6.7500 ;
      RECT 26.2360 5.6565 26.2620 6.7500 ;
      RECT 26.1280 5.6565 26.1540 6.7500 ;
      RECT 26.0200 5.6565 26.0460 6.7500 ;
      RECT 25.9120 5.6565 25.9380 6.7500 ;
      RECT 25.8040 5.6565 25.8300 6.7500 ;
      RECT 25.6960 5.6565 25.7220 6.7500 ;
      RECT 25.5880 5.6565 25.6140 6.7500 ;
      RECT 25.4800 5.6565 25.5060 6.7500 ;
      RECT 25.3720 5.6565 25.3980 6.7500 ;
      RECT 25.2640 5.6565 25.2900 6.7500 ;
      RECT 25.1560 5.6565 25.1820 6.7500 ;
      RECT 25.0480 5.6565 25.0740 6.7500 ;
      RECT 24.9400 5.6565 24.9660 6.7500 ;
      RECT 24.8320 5.6565 24.8580 6.7500 ;
      RECT 24.7240 5.6565 24.7500 6.7500 ;
      RECT 24.6160 5.6565 24.6420 6.7500 ;
      RECT 24.5080 5.6565 24.5340 6.7500 ;
      RECT 24.4000 5.6565 24.4260 6.7500 ;
      RECT 24.2920 5.6565 24.3180 6.7500 ;
      RECT 24.1840 5.6565 24.2100 6.7500 ;
      RECT 24.0760 5.6565 24.1020 6.7500 ;
      RECT 23.9680 5.6565 23.9940 6.7500 ;
      RECT 23.8600 5.6565 23.8860 6.7500 ;
      RECT 23.7520 5.6565 23.7780 6.7500 ;
      RECT 23.6440 5.6565 23.6700 6.7500 ;
      RECT 23.5360 5.6565 23.5620 6.7500 ;
      RECT 23.4280 5.6565 23.4540 6.7500 ;
      RECT 23.3200 5.6565 23.3460 6.7500 ;
      RECT 23.2120 5.6565 23.2380 6.7500 ;
      RECT 23.1040 5.6565 23.1300 6.7500 ;
      RECT 22.9960 5.6565 23.0220 6.7500 ;
      RECT 22.8880 5.6565 22.9140 6.7500 ;
      RECT 22.7800 5.6565 22.8060 6.7500 ;
      RECT 22.6720 5.6565 22.6980 6.7500 ;
      RECT 22.5640 5.6565 22.5900 6.7500 ;
      RECT 22.4560 5.6565 22.4820 6.7500 ;
      RECT 22.3480 5.6565 22.3740 6.7500 ;
      RECT 22.2400 5.6565 22.2660 6.7500 ;
      RECT 22.1320 5.6565 22.1580 6.7500 ;
      RECT 22.0240 5.6565 22.0500 6.7500 ;
      RECT 21.9160 5.6565 21.9420 6.7500 ;
      RECT 21.8080 5.6565 21.8340 6.7500 ;
      RECT 21.7000 5.6565 21.7260 6.7500 ;
      RECT 21.5920 5.6565 21.6180 6.7500 ;
      RECT 21.4840 5.6565 21.5100 6.7500 ;
      RECT 21.3760 5.6565 21.4020 6.7500 ;
      RECT 21.2680 5.6565 21.2940 6.7500 ;
      RECT 21.1600 5.6565 21.1860 6.7500 ;
      RECT 21.0520 5.6565 21.0780 6.7500 ;
      RECT 20.9440 5.6565 20.9700 6.7500 ;
      RECT 20.8360 5.6565 20.8620 6.7500 ;
      RECT 20.7280 5.6565 20.7540 6.7500 ;
      RECT 20.6200 5.6565 20.6460 6.7500 ;
      RECT 20.5120 5.6565 20.5380 6.7500 ;
      RECT 20.4040 5.6565 20.4300 6.7500 ;
      RECT 20.2960 5.6565 20.3220 6.7500 ;
      RECT 20.1880 5.6565 20.2140 6.7500 ;
      RECT 20.0800 5.6565 20.1060 6.7500 ;
      RECT 19.9720 5.6565 19.9980 6.7500 ;
      RECT 19.8640 5.6565 19.8900 6.7500 ;
      RECT 19.7560 5.6565 19.7820 6.7500 ;
      RECT 19.6480 5.6565 19.6740 6.7500 ;
      RECT 19.5400 5.6565 19.5660 6.7500 ;
      RECT 19.4320 5.6565 19.4580 6.7500 ;
      RECT 19.3240 5.6565 19.3500 6.7500 ;
      RECT 19.2160 5.6565 19.2420 6.7500 ;
      RECT 19.1080 5.6565 19.1340 6.7500 ;
      RECT 19.0000 5.6565 19.0260 6.7500 ;
      RECT 18.8920 5.6565 18.9180 6.7500 ;
      RECT 18.7840 5.6565 18.8100 6.7500 ;
      RECT 18.6760 5.6565 18.7020 6.7500 ;
      RECT 18.5680 5.6565 18.5940 6.7500 ;
      RECT 18.4600 5.6565 18.4860 6.7500 ;
      RECT 18.3520 5.6565 18.3780 6.7500 ;
      RECT 18.2440 5.6565 18.2700 6.7500 ;
      RECT 18.1360 5.6565 18.1620 6.7500 ;
      RECT 18.0280 5.6565 18.0540 6.7500 ;
      RECT 17.9200 5.6565 17.9460 6.7500 ;
      RECT 17.8120 5.6565 17.8380 6.7500 ;
      RECT 17.7040 5.6565 17.7300 6.7500 ;
      RECT 17.5960 5.6565 17.6220 6.7500 ;
      RECT 17.4880 5.6565 17.5140 6.7500 ;
      RECT 17.3800 5.6565 17.4060 6.7500 ;
      RECT 17.2720 5.6565 17.2980 6.7500 ;
      RECT 17.1640 5.6565 17.1900 6.7500 ;
      RECT 17.0560 5.6565 17.0820 6.7500 ;
      RECT 16.9480 5.6565 16.9740 6.7500 ;
      RECT 16.8400 5.6565 16.8660 6.7500 ;
      RECT 16.7320 5.6565 16.7580 6.7500 ;
      RECT 16.6240 5.6565 16.6500 6.7500 ;
      RECT 16.5160 5.6565 16.5420 6.7500 ;
      RECT 16.4080 5.6565 16.4340 6.7500 ;
      RECT 16.3000 5.6565 16.3260 6.7500 ;
      RECT 16.0870 5.6565 16.1640 6.7500 ;
      RECT 14.1940 5.6565 14.2710 6.7500 ;
      RECT 14.0320 5.6565 14.0580 6.7500 ;
      RECT 13.9240 5.6565 13.9500 6.7500 ;
      RECT 13.8160 5.6565 13.8420 6.7500 ;
      RECT 13.7080 5.6565 13.7340 6.7500 ;
      RECT 13.6000 5.6565 13.6260 6.7500 ;
      RECT 13.4920 5.6565 13.5180 6.7500 ;
      RECT 13.3840 5.6565 13.4100 6.7500 ;
      RECT 13.2760 5.6565 13.3020 6.7500 ;
      RECT 13.1680 5.6565 13.1940 6.7500 ;
      RECT 13.0600 5.6565 13.0860 6.7500 ;
      RECT 12.9520 5.6565 12.9780 6.7500 ;
      RECT 12.8440 5.6565 12.8700 6.7500 ;
      RECT 12.7360 5.6565 12.7620 6.7500 ;
      RECT 12.6280 5.6565 12.6540 6.7500 ;
      RECT 12.5200 5.6565 12.5460 6.7500 ;
      RECT 12.4120 5.6565 12.4380 6.7500 ;
      RECT 12.3040 5.6565 12.3300 6.7500 ;
      RECT 12.1960 5.6565 12.2220 6.7500 ;
      RECT 12.0880 5.6565 12.1140 6.7500 ;
      RECT 11.9800 5.6565 12.0060 6.7500 ;
      RECT 11.8720 5.6565 11.8980 6.7500 ;
      RECT 11.7640 5.6565 11.7900 6.7500 ;
      RECT 11.6560 5.6565 11.6820 6.7500 ;
      RECT 11.5480 5.6565 11.5740 6.7500 ;
      RECT 11.4400 5.6565 11.4660 6.7500 ;
      RECT 11.3320 5.6565 11.3580 6.7500 ;
      RECT 11.2240 5.6565 11.2500 6.7500 ;
      RECT 11.1160 5.6565 11.1420 6.7500 ;
      RECT 11.0080 5.6565 11.0340 6.7500 ;
      RECT 10.9000 5.6565 10.9260 6.7500 ;
      RECT 10.7920 5.6565 10.8180 6.7500 ;
      RECT 10.6840 5.6565 10.7100 6.7500 ;
      RECT 10.5760 5.6565 10.6020 6.7500 ;
      RECT 10.4680 5.6565 10.4940 6.7500 ;
      RECT 10.3600 5.6565 10.3860 6.7500 ;
      RECT 10.2520 5.6565 10.2780 6.7500 ;
      RECT 10.1440 5.6565 10.1700 6.7500 ;
      RECT 10.0360 5.6565 10.0620 6.7500 ;
      RECT 9.9280 5.6565 9.9540 6.7500 ;
      RECT 9.8200 5.6565 9.8460 6.7500 ;
      RECT 9.7120 5.6565 9.7380 6.7500 ;
      RECT 9.6040 5.6565 9.6300 6.7500 ;
      RECT 9.4960 5.6565 9.5220 6.7500 ;
      RECT 9.3880 5.6565 9.4140 6.7500 ;
      RECT 9.2800 5.6565 9.3060 6.7500 ;
      RECT 9.1720 5.6565 9.1980 6.7500 ;
      RECT 9.0640 5.6565 9.0900 6.7500 ;
      RECT 8.9560 5.6565 8.9820 6.7500 ;
      RECT 8.8480 5.6565 8.8740 6.7500 ;
      RECT 8.7400 5.6565 8.7660 6.7500 ;
      RECT 8.6320 5.6565 8.6580 6.7500 ;
      RECT 8.5240 5.6565 8.5500 6.7500 ;
      RECT 8.4160 5.6565 8.4420 6.7500 ;
      RECT 8.3080 5.6565 8.3340 6.7500 ;
      RECT 8.2000 5.6565 8.2260 6.7500 ;
      RECT 8.0920 5.6565 8.1180 6.7500 ;
      RECT 7.9840 5.6565 8.0100 6.7500 ;
      RECT 7.8760 5.6565 7.9020 6.7500 ;
      RECT 7.7680 5.6565 7.7940 6.7500 ;
      RECT 7.6600 5.6565 7.6860 6.7500 ;
      RECT 7.5520 5.6565 7.5780 6.7500 ;
      RECT 7.4440 5.6565 7.4700 6.7500 ;
      RECT 7.3360 5.6565 7.3620 6.7500 ;
      RECT 7.2280 5.6565 7.2540 6.7500 ;
      RECT 7.1200 5.6565 7.1460 6.7500 ;
      RECT 7.0120 5.6565 7.0380 6.7500 ;
      RECT 6.9040 5.6565 6.9300 6.7500 ;
      RECT 6.7960 5.6565 6.8220 6.7500 ;
      RECT 6.6880 5.6565 6.7140 6.7500 ;
      RECT 6.5800 5.6565 6.6060 6.7500 ;
      RECT 6.4720 5.6565 6.4980 6.7500 ;
      RECT 6.3640 5.6565 6.3900 6.7500 ;
      RECT 6.2560 5.6565 6.2820 6.7500 ;
      RECT 6.1480 5.6565 6.1740 6.7500 ;
      RECT 6.0400 5.6565 6.0660 6.7500 ;
      RECT 5.9320 5.6565 5.9580 6.7500 ;
      RECT 5.8240 5.6565 5.8500 6.7500 ;
      RECT 5.7160 5.6565 5.7420 6.7500 ;
      RECT 5.6080 5.6565 5.6340 6.7500 ;
      RECT 5.5000 5.6565 5.5260 6.7500 ;
      RECT 5.3920 5.6565 5.4180 6.7500 ;
      RECT 5.2840 5.6565 5.3100 6.7500 ;
      RECT 5.1760 5.6565 5.2020 6.7500 ;
      RECT 5.0680 5.6565 5.0940 6.7500 ;
      RECT 4.9600 5.6565 4.9860 6.7500 ;
      RECT 4.8520 5.6565 4.8780 6.7500 ;
      RECT 4.7440 5.6565 4.7700 6.7500 ;
      RECT 4.6360 5.6565 4.6620 6.7500 ;
      RECT 4.5280 5.6565 4.5540 6.7500 ;
      RECT 4.4200 5.6565 4.4460 6.7500 ;
      RECT 4.3120 5.6565 4.3380 6.7500 ;
      RECT 4.2040 5.6565 4.2300 6.7500 ;
      RECT 4.0960 5.6565 4.1220 6.7500 ;
      RECT 3.9880 5.6565 4.0140 6.7500 ;
      RECT 3.8800 5.6565 3.9060 6.7500 ;
      RECT 3.7720 5.6565 3.7980 6.7500 ;
      RECT 3.6640 5.6565 3.6900 6.7500 ;
      RECT 3.5560 5.6565 3.5820 6.7500 ;
      RECT 3.4480 5.6565 3.4740 6.7500 ;
      RECT 3.3400 5.6565 3.3660 6.7500 ;
      RECT 3.2320 5.6565 3.2580 6.7500 ;
      RECT 3.1240 5.6565 3.1500 6.7500 ;
      RECT 3.0160 5.6565 3.0420 6.7500 ;
      RECT 2.9080 5.6565 2.9340 6.7500 ;
      RECT 2.8000 5.6565 2.8260 6.7500 ;
      RECT 2.6920 5.6565 2.7180 6.7500 ;
      RECT 2.5840 5.6565 2.6100 6.7500 ;
      RECT 2.4760 5.6565 2.5020 6.7500 ;
      RECT 2.3680 5.6565 2.3940 6.7500 ;
      RECT 2.2600 5.6565 2.2860 6.7500 ;
      RECT 2.1520 5.6565 2.1780 6.7500 ;
      RECT 2.0440 5.6565 2.0700 6.7500 ;
      RECT 1.9360 5.6565 1.9620 6.7500 ;
      RECT 1.8280 5.6565 1.8540 6.7500 ;
      RECT 1.7200 5.6565 1.7460 6.7500 ;
      RECT 1.6120 5.6565 1.6380 6.7500 ;
      RECT 1.5040 5.6565 1.5300 6.7500 ;
      RECT 1.3960 5.6565 1.4220 6.7500 ;
      RECT 1.2880 5.6565 1.3140 6.7500 ;
      RECT 1.1800 5.6565 1.2060 6.7500 ;
      RECT 1.0720 5.6565 1.0980 6.7500 ;
      RECT 0.9640 5.6565 0.9900 6.7500 ;
      RECT 0.8560 5.6565 0.8820 6.7500 ;
      RECT 0.7480 5.6565 0.7740 6.7500 ;
      RECT 0.6400 5.6565 0.6660 6.7500 ;
      RECT 0.5320 5.6565 0.5580 6.7500 ;
      RECT 0.4240 5.6565 0.4500 6.7500 ;
      RECT 0.3160 5.6565 0.3420 6.7500 ;
      RECT 0.2080 5.6565 0.2340 6.7500 ;
      RECT 0.0050 5.6565 0.0900 6.7500 ;
      RECT 15.5530 6.7365 15.6810 7.8300 ;
      RECT 15.5390 7.4020 15.6810 7.7245 ;
      RECT 15.3190 7.1290 15.4530 7.8300 ;
      RECT 15.2960 7.4640 15.4530 7.7220 ;
      RECT 15.3190 6.7365 15.4170 7.8300 ;
      RECT 15.3190 6.8575 15.4310 7.0970 ;
      RECT 15.3190 6.7365 15.4530 6.8255 ;
      RECT 15.0940 7.1870 15.2280 7.8300 ;
      RECT 15.0940 6.7365 15.1920 7.8300 ;
      RECT 14.6770 6.7365 14.7600 7.8300 ;
      RECT 14.6770 6.8250 14.7740 7.7605 ;
      RECT 30.2680 6.7365 30.3530 7.8300 ;
      RECT 30.1240 6.7365 30.1500 7.8300 ;
      RECT 30.0160 6.7365 30.0420 7.8300 ;
      RECT 29.9080 6.7365 29.9340 7.8300 ;
      RECT 29.8000 6.7365 29.8260 7.8300 ;
      RECT 29.6920 6.7365 29.7180 7.8300 ;
      RECT 29.5840 6.7365 29.6100 7.8300 ;
      RECT 29.4760 6.7365 29.5020 7.8300 ;
      RECT 29.3680 6.7365 29.3940 7.8300 ;
      RECT 29.2600 6.7365 29.2860 7.8300 ;
      RECT 29.1520 6.7365 29.1780 7.8300 ;
      RECT 29.0440 6.7365 29.0700 7.8300 ;
      RECT 28.9360 6.7365 28.9620 7.8300 ;
      RECT 28.8280 6.7365 28.8540 7.8300 ;
      RECT 28.7200 6.7365 28.7460 7.8300 ;
      RECT 28.6120 6.7365 28.6380 7.8300 ;
      RECT 28.5040 6.7365 28.5300 7.8300 ;
      RECT 28.3960 6.7365 28.4220 7.8300 ;
      RECT 28.2880 6.7365 28.3140 7.8300 ;
      RECT 28.1800 6.7365 28.2060 7.8300 ;
      RECT 28.0720 6.7365 28.0980 7.8300 ;
      RECT 27.9640 6.7365 27.9900 7.8300 ;
      RECT 27.8560 6.7365 27.8820 7.8300 ;
      RECT 27.7480 6.7365 27.7740 7.8300 ;
      RECT 27.6400 6.7365 27.6660 7.8300 ;
      RECT 27.5320 6.7365 27.5580 7.8300 ;
      RECT 27.4240 6.7365 27.4500 7.8300 ;
      RECT 27.3160 6.7365 27.3420 7.8300 ;
      RECT 27.2080 6.7365 27.2340 7.8300 ;
      RECT 27.1000 6.7365 27.1260 7.8300 ;
      RECT 26.9920 6.7365 27.0180 7.8300 ;
      RECT 26.8840 6.7365 26.9100 7.8300 ;
      RECT 26.7760 6.7365 26.8020 7.8300 ;
      RECT 26.6680 6.7365 26.6940 7.8300 ;
      RECT 26.5600 6.7365 26.5860 7.8300 ;
      RECT 26.4520 6.7365 26.4780 7.8300 ;
      RECT 26.3440 6.7365 26.3700 7.8300 ;
      RECT 26.2360 6.7365 26.2620 7.8300 ;
      RECT 26.1280 6.7365 26.1540 7.8300 ;
      RECT 26.0200 6.7365 26.0460 7.8300 ;
      RECT 25.9120 6.7365 25.9380 7.8300 ;
      RECT 25.8040 6.7365 25.8300 7.8300 ;
      RECT 25.6960 6.7365 25.7220 7.8300 ;
      RECT 25.5880 6.7365 25.6140 7.8300 ;
      RECT 25.4800 6.7365 25.5060 7.8300 ;
      RECT 25.3720 6.7365 25.3980 7.8300 ;
      RECT 25.2640 6.7365 25.2900 7.8300 ;
      RECT 25.1560 6.7365 25.1820 7.8300 ;
      RECT 25.0480 6.7365 25.0740 7.8300 ;
      RECT 24.9400 6.7365 24.9660 7.8300 ;
      RECT 24.8320 6.7365 24.8580 7.8300 ;
      RECT 24.7240 6.7365 24.7500 7.8300 ;
      RECT 24.6160 6.7365 24.6420 7.8300 ;
      RECT 24.5080 6.7365 24.5340 7.8300 ;
      RECT 24.4000 6.7365 24.4260 7.8300 ;
      RECT 24.2920 6.7365 24.3180 7.8300 ;
      RECT 24.1840 6.7365 24.2100 7.8300 ;
      RECT 24.0760 6.7365 24.1020 7.8300 ;
      RECT 23.9680 6.7365 23.9940 7.8300 ;
      RECT 23.8600 6.7365 23.8860 7.8300 ;
      RECT 23.7520 6.7365 23.7780 7.8300 ;
      RECT 23.6440 6.7365 23.6700 7.8300 ;
      RECT 23.5360 6.7365 23.5620 7.8300 ;
      RECT 23.4280 6.7365 23.4540 7.8300 ;
      RECT 23.3200 6.7365 23.3460 7.8300 ;
      RECT 23.2120 6.7365 23.2380 7.8300 ;
      RECT 23.1040 6.7365 23.1300 7.8300 ;
      RECT 22.9960 6.7365 23.0220 7.8300 ;
      RECT 22.8880 6.7365 22.9140 7.8300 ;
      RECT 22.7800 6.7365 22.8060 7.8300 ;
      RECT 22.6720 6.7365 22.6980 7.8300 ;
      RECT 22.5640 6.7365 22.5900 7.8300 ;
      RECT 22.4560 6.7365 22.4820 7.8300 ;
      RECT 22.3480 6.7365 22.3740 7.8300 ;
      RECT 22.2400 6.7365 22.2660 7.8300 ;
      RECT 22.1320 6.7365 22.1580 7.8300 ;
      RECT 22.0240 6.7365 22.0500 7.8300 ;
      RECT 21.9160 6.7365 21.9420 7.8300 ;
      RECT 21.8080 6.7365 21.8340 7.8300 ;
      RECT 21.7000 6.7365 21.7260 7.8300 ;
      RECT 21.5920 6.7365 21.6180 7.8300 ;
      RECT 21.4840 6.7365 21.5100 7.8300 ;
      RECT 21.3760 6.7365 21.4020 7.8300 ;
      RECT 21.2680 6.7365 21.2940 7.8300 ;
      RECT 21.1600 6.7365 21.1860 7.8300 ;
      RECT 21.0520 6.7365 21.0780 7.8300 ;
      RECT 20.9440 6.7365 20.9700 7.8300 ;
      RECT 20.8360 6.7365 20.8620 7.8300 ;
      RECT 20.7280 6.7365 20.7540 7.8300 ;
      RECT 20.6200 6.7365 20.6460 7.8300 ;
      RECT 20.5120 6.7365 20.5380 7.8300 ;
      RECT 20.4040 6.7365 20.4300 7.8300 ;
      RECT 20.2960 6.7365 20.3220 7.8300 ;
      RECT 20.1880 6.7365 20.2140 7.8300 ;
      RECT 20.0800 6.7365 20.1060 7.8300 ;
      RECT 19.9720 6.7365 19.9980 7.8300 ;
      RECT 19.8640 6.7365 19.8900 7.8300 ;
      RECT 19.7560 6.7365 19.7820 7.8300 ;
      RECT 19.6480 6.7365 19.6740 7.8300 ;
      RECT 19.5400 6.7365 19.5660 7.8300 ;
      RECT 19.4320 6.7365 19.4580 7.8300 ;
      RECT 19.3240 6.7365 19.3500 7.8300 ;
      RECT 19.2160 6.7365 19.2420 7.8300 ;
      RECT 19.1080 6.7365 19.1340 7.8300 ;
      RECT 19.0000 6.7365 19.0260 7.8300 ;
      RECT 18.8920 6.7365 18.9180 7.8300 ;
      RECT 18.7840 6.7365 18.8100 7.8300 ;
      RECT 18.6760 6.7365 18.7020 7.8300 ;
      RECT 18.5680 6.7365 18.5940 7.8300 ;
      RECT 18.4600 6.7365 18.4860 7.8300 ;
      RECT 18.3520 6.7365 18.3780 7.8300 ;
      RECT 18.2440 6.7365 18.2700 7.8300 ;
      RECT 18.1360 6.7365 18.1620 7.8300 ;
      RECT 18.0280 6.7365 18.0540 7.8300 ;
      RECT 17.9200 6.7365 17.9460 7.8300 ;
      RECT 17.8120 6.7365 17.8380 7.8300 ;
      RECT 17.7040 6.7365 17.7300 7.8300 ;
      RECT 17.5960 6.7365 17.6220 7.8300 ;
      RECT 17.4880 6.7365 17.5140 7.8300 ;
      RECT 17.3800 6.7365 17.4060 7.8300 ;
      RECT 17.2720 6.7365 17.2980 7.8300 ;
      RECT 17.1640 6.7365 17.1900 7.8300 ;
      RECT 17.0560 6.7365 17.0820 7.8300 ;
      RECT 16.9480 6.7365 16.9740 7.8300 ;
      RECT 16.8400 6.7365 16.8660 7.8300 ;
      RECT 16.7320 6.7365 16.7580 7.8300 ;
      RECT 16.6240 6.7365 16.6500 7.8300 ;
      RECT 16.5160 6.7365 16.5420 7.8300 ;
      RECT 16.4080 6.7365 16.4340 7.8300 ;
      RECT 16.3000 6.7365 16.3260 7.8300 ;
      RECT 16.0870 6.7365 16.1640 7.8300 ;
      RECT 14.1940 6.7365 14.2710 7.8300 ;
      RECT 14.0320 6.7365 14.0580 7.8300 ;
      RECT 13.9240 6.7365 13.9500 7.8300 ;
      RECT 13.8160 6.7365 13.8420 7.8300 ;
      RECT 13.7080 6.7365 13.7340 7.8300 ;
      RECT 13.6000 6.7365 13.6260 7.8300 ;
      RECT 13.4920 6.7365 13.5180 7.8300 ;
      RECT 13.3840 6.7365 13.4100 7.8300 ;
      RECT 13.2760 6.7365 13.3020 7.8300 ;
      RECT 13.1680 6.7365 13.1940 7.8300 ;
      RECT 13.0600 6.7365 13.0860 7.8300 ;
      RECT 12.9520 6.7365 12.9780 7.8300 ;
      RECT 12.8440 6.7365 12.8700 7.8300 ;
      RECT 12.7360 6.7365 12.7620 7.8300 ;
      RECT 12.6280 6.7365 12.6540 7.8300 ;
      RECT 12.5200 6.7365 12.5460 7.8300 ;
      RECT 12.4120 6.7365 12.4380 7.8300 ;
      RECT 12.3040 6.7365 12.3300 7.8300 ;
      RECT 12.1960 6.7365 12.2220 7.8300 ;
      RECT 12.0880 6.7365 12.1140 7.8300 ;
      RECT 11.9800 6.7365 12.0060 7.8300 ;
      RECT 11.8720 6.7365 11.8980 7.8300 ;
      RECT 11.7640 6.7365 11.7900 7.8300 ;
      RECT 11.6560 6.7365 11.6820 7.8300 ;
      RECT 11.5480 6.7365 11.5740 7.8300 ;
      RECT 11.4400 6.7365 11.4660 7.8300 ;
      RECT 11.3320 6.7365 11.3580 7.8300 ;
      RECT 11.2240 6.7365 11.2500 7.8300 ;
      RECT 11.1160 6.7365 11.1420 7.8300 ;
      RECT 11.0080 6.7365 11.0340 7.8300 ;
      RECT 10.9000 6.7365 10.9260 7.8300 ;
      RECT 10.7920 6.7365 10.8180 7.8300 ;
      RECT 10.6840 6.7365 10.7100 7.8300 ;
      RECT 10.5760 6.7365 10.6020 7.8300 ;
      RECT 10.4680 6.7365 10.4940 7.8300 ;
      RECT 10.3600 6.7365 10.3860 7.8300 ;
      RECT 10.2520 6.7365 10.2780 7.8300 ;
      RECT 10.1440 6.7365 10.1700 7.8300 ;
      RECT 10.0360 6.7365 10.0620 7.8300 ;
      RECT 9.9280 6.7365 9.9540 7.8300 ;
      RECT 9.8200 6.7365 9.8460 7.8300 ;
      RECT 9.7120 6.7365 9.7380 7.8300 ;
      RECT 9.6040 6.7365 9.6300 7.8300 ;
      RECT 9.4960 6.7365 9.5220 7.8300 ;
      RECT 9.3880 6.7365 9.4140 7.8300 ;
      RECT 9.2800 6.7365 9.3060 7.8300 ;
      RECT 9.1720 6.7365 9.1980 7.8300 ;
      RECT 9.0640 6.7365 9.0900 7.8300 ;
      RECT 8.9560 6.7365 8.9820 7.8300 ;
      RECT 8.8480 6.7365 8.8740 7.8300 ;
      RECT 8.7400 6.7365 8.7660 7.8300 ;
      RECT 8.6320 6.7365 8.6580 7.8300 ;
      RECT 8.5240 6.7365 8.5500 7.8300 ;
      RECT 8.4160 6.7365 8.4420 7.8300 ;
      RECT 8.3080 6.7365 8.3340 7.8300 ;
      RECT 8.2000 6.7365 8.2260 7.8300 ;
      RECT 8.0920 6.7365 8.1180 7.8300 ;
      RECT 7.9840 6.7365 8.0100 7.8300 ;
      RECT 7.8760 6.7365 7.9020 7.8300 ;
      RECT 7.7680 6.7365 7.7940 7.8300 ;
      RECT 7.6600 6.7365 7.6860 7.8300 ;
      RECT 7.5520 6.7365 7.5780 7.8300 ;
      RECT 7.4440 6.7365 7.4700 7.8300 ;
      RECT 7.3360 6.7365 7.3620 7.8300 ;
      RECT 7.2280 6.7365 7.2540 7.8300 ;
      RECT 7.1200 6.7365 7.1460 7.8300 ;
      RECT 7.0120 6.7365 7.0380 7.8300 ;
      RECT 6.9040 6.7365 6.9300 7.8300 ;
      RECT 6.7960 6.7365 6.8220 7.8300 ;
      RECT 6.6880 6.7365 6.7140 7.8300 ;
      RECT 6.5800 6.7365 6.6060 7.8300 ;
      RECT 6.4720 6.7365 6.4980 7.8300 ;
      RECT 6.3640 6.7365 6.3900 7.8300 ;
      RECT 6.2560 6.7365 6.2820 7.8300 ;
      RECT 6.1480 6.7365 6.1740 7.8300 ;
      RECT 6.0400 6.7365 6.0660 7.8300 ;
      RECT 5.9320 6.7365 5.9580 7.8300 ;
      RECT 5.8240 6.7365 5.8500 7.8300 ;
      RECT 5.7160 6.7365 5.7420 7.8300 ;
      RECT 5.6080 6.7365 5.6340 7.8300 ;
      RECT 5.5000 6.7365 5.5260 7.8300 ;
      RECT 5.3920 6.7365 5.4180 7.8300 ;
      RECT 5.2840 6.7365 5.3100 7.8300 ;
      RECT 5.1760 6.7365 5.2020 7.8300 ;
      RECT 5.0680 6.7365 5.0940 7.8300 ;
      RECT 4.9600 6.7365 4.9860 7.8300 ;
      RECT 4.8520 6.7365 4.8780 7.8300 ;
      RECT 4.7440 6.7365 4.7700 7.8300 ;
      RECT 4.6360 6.7365 4.6620 7.8300 ;
      RECT 4.5280 6.7365 4.5540 7.8300 ;
      RECT 4.4200 6.7365 4.4460 7.8300 ;
      RECT 4.3120 6.7365 4.3380 7.8300 ;
      RECT 4.2040 6.7365 4.2300 7.8300 ;
      RECT 4.0960 6.7365 4.1220 7.8300 ;
      RECT 3.9880 6.7365 4.0140 7.8300 ;
      RECT 3.8800 6.7365 3.9060 7.8300 ;
      RECT 3.7720 6.7365 3.7980 7.8300 ;
      RECT 3.6640 6.7365 3.6900 7.8300 ;
      RECT 3.5560 6.7365 3.5820 7.8300 ;
      RECT 3.4480 6.7365 3.4740 7.8300 ;
      RECT 3.3400 6.7365 3.3660 7.8300 ;
      RECT 3.2320 6.7365 3.2580 7.8300 ;
      RECT 3.1240 6.7365 3.1500 7.8300 ;
      RECT 3.0160 6.7365 3.0420 7.8300 ;
      RECT 2.9080 6.7365 2.9340 7.8300 ;
      RECT 2.8000 6.7365 2.8260 7.8300 ;
      RECT 2.6920 6.7365 2.7180 7.8300 ;
      RECT 2.5840 6.7365 2.6100 7.8300 ;
      RECT 2.4760 6.7365 2.5020 7.8300 ;
      RECT 2.3680 6.7365 2.3940 7.8300 ;
      RECT 2.2600 6.7365 2.2860 7.8300 ;
      RECT 2.1520 6.7365 2.1780 7.8300 ;
      RECT 2.0440 6.7365 2.0700 7.8300 ;
      RECT 1.9360 6.7365 1.9620 7.8300 ;
      RECT 1.8280 6.7365 1.8540 7.8300 ;
      RECT 1.7200 6.7365 1.7460 7.8300 ;
      RECT 1.6120 6.7365 1.6380 7.8300 ;
      RECT 1.5040 6.7365 1.5300 7.8300 ;
      RECT 1.3960 6.7365 1.4220 7.8300 ;
      RECT 1.2880 6.7365 1.3140 7.8300 ;
      RECT 1.1800 6.7365 1.2060 7.8300 ;
      RECT 1.0720 6.7365 1.0980 7.8300 ;
      RECT 0.9640 6.7365 0.9900 7.8300 ;
      RECT 0.8560 6.7365 0.8820 7.8300 ;
      RECT 0.7480 6.7365 0.7740 7.8300 ;
      RECT 0.6400 6.7365 0.6660 7.8300 ;
      RECT 0.5320 6.7365 0.5580 7.8300 ;
      RECT 0.4240 6.7365 0.4500 7.8300 ;
      RECT 0.3160 6.7365 0.3420 7.8300 ;
      RECT 0.2080 6.7365 0.2340 7.8300 ;
      RECT 0.0050 6.7365 0.0900 7.8300 ;
      RECT 15.5530 7.8165 15.6810 8.9100 ;
      RECT 15.5390 8.4820 15.6810 8.8045 ;
      RECT 15.3190 8.2090 15.4530 8.9100 ;
      RECT 15.2960 8.5440 15.4530 8.8020 ;
      RECT 15.3190 7.8165 15.4170 8.9100 ;
      RECT 15.3190 7.9375 15.4310 8.1770 ;
      RECT 15.3190 7.8165 15.4530 7.9055 ;
      RECT 15.0940 8.2670 15.2280 8.9100 ;
      RECT 15.0940 7.8165 15.1920 8.9100 ;
      RECT 14.6770 7.8165 14.7600 8.9100 ;
      RECT 14.6770 7.9050 14.7740 8.8405 ;
      RECT 30.2680 7.8165 30.3530 8.9100 ;
      RECT 30.1240 7.8165 30.1500 8.9100 ;
      RECT 30.0160 7.8165 30.0420 8.9100 ;
      RECT 29.9080 7.8165 29.9340 8.9100 ;
      RECT 29.8000 7.8165 29.8260 8.9100 ;
      RECT 29.6920 7.8165 29.7180 8.9100 ;
      RECT 29.5840 7.8165 29.6100 8.9100 ;
      RECT 29.4760 7.8165 29.5020 8.9100 ;
      RECT 29.3680 7.8165 29.3940 8.9100 ;
      RECT 29.2600 7.8165 29.2860 8.9100 ;
      RECT 29.1520 7.8165 29.1780 8.9100 ;
      RECT 29.0440 7.8165 29.0700 8.9100 ;
      RECT 28.9360 7.8165 28.9620 8.9100 ;
      RECT 28.8280 7.8165 28.8540 8.9100 ;
      RECT 28.7200 7.8165 28.7460 8.9100 ;
      RECT 28.6120 7.8165 28.6380 8.9100 ;
      RECT 28.5040 7.8165 28.5300 8.9100 ;
      RECT 28.3960 7.8165 28.4220 8.9100 ;
      RECT 28.2880 7.8165 28.3140 8.9100 ;
      RECT 28.1800 7.8165 28.2060 8.9100 ;
      RECT 28.0720 7.8165 28.0980 8.9100 ;
      RECT 27.9640 7.8165 27.9900 8.9100 ;
      RECT 27.8560 7.8165 27.8820 8.9100 ;
      RECT 27.7480 7.8165 27.7740 8.9100 ;
      RECT 27.6400 7.8165 27.6660 8.9100 ;
      RECT 27.5320 7.8165 27.5580 8.9100 ;
      RECT 27.4240 7.8165 27.4500 8.9100 ;
      RECT 27.3160 7.8165 27.3420 8.9100 ;
      RECT 27.2080 7.8165 27.2340 8.9100 ;
      RECT 27.1000 7.8165 27.1260 8.9100 ;
      RECT 26.9920 7.8165 27.0180 8.9100 ;
      RECT 26.8840 7.8165 26.9100 8.9100 ;
      RECT 26.7760 7.8165 26.8020 8.9100 ;
      RECT 26.6680 7.8165 26.6940 8.9100 ;
      RECT 26.5600 7.8165 26.5860 8.9100 ;
      RECT 26.4520 7.8165 26.4780 8.9100 ;
      RECT 26.3440 7.8165 26.3700 8.9100 ;
      RECT 26.2360 7.8165 26.2620 8.9100 ;
      RECT 26.1280 7.8165 26.1540 8.9100 ;
      RECT 26.0200 7.8165 26.0460 8.9100 ;
      RECT 25.9120 7.8165 25.9380 8.9100 ;
      RECT 25.8040 7.8165 25.8300 8.9100 ;
      RECT 25.6960 7.8165 25.7220 8.9100 ;
      RECT 25.5880 7.8165 25.6140 8.9100 ;
      RECT 25.4800 7.8165 25.5060 8.9100 ;
      RECT 25.3720 7.8165 25.3980 8.9100 ;
      RECT 25.2640 7.8165 25.2900 8.9100 ;
      RECT 25.1560 7.8165 25.1820 8.9100 ;
      RECT 25.0480 7.8165 25.0740 8.9100 ;
      RECT 24.9400 7.8165 24.9660 8.9100 ;
      RECT 24.8320 7.8165 24.8580 8.9100 ;
      RECT 24.7240 7.8165 24.7500 8.9100 ;
      RECT 24.6160 7.8165 24.6420 8.9100 ;
      RECT 24.5080 7.8165 24.5340 8.9100 ;
      RECT 24.4000 7.8165 24.4260 8.9100 ;
      RECT 24.2920 7.8165 24.3180 8.9100 ;
      RECT 24.1840 7.8165 24.2100 8.9100 ;
      RECT 24.0760 7.8165 24.1020 8.9100 ;
      RECT 23.9680 7.8165 23.9940 8.9100 ;
      RECT 23.8600 7.8165 23.8860 8.9100 ;
      RECT 23.7520 7.8165 23.7780 8.9100 ;
      RECT 23.6440 7.8165 23.6700 8.9100 ;
      RECT 23.5360 7.8165 23.5620 8.9100 ;
      RECT 23.4280 7.8165 23.4540 8.9100 ;
      RECT 23.3200 7.8165 23.3460 8.9100 ;
      RECT 23.2120 7.8165 23.2380 8.9100 ;
      RECT 23.1040 7.8165 23.1300 8.9100 ;
      RECT 22.9960 7.8165 23.0220 8.9100 ;
      RECT 22.8880 7.8165 22.9140 8.9100 ;
      RECT 22.7800 7.8165 22.8060 8.9100 ;
      RECT 22.6720 7.8165 22.6980 8.9100 ;
      RECT 22.5640 7.8165 22.5900 8.9100 ;
      RECT 22.4560 7.8165 22.4820 8.9100 ;
      RECT 22.3480 7.8165 22.3740 8.9100 ;
      RECT 22.2400 7.8165 22.2660 8.9100 ;
      RECT 22.1320 7.8165 22.1580 8.9100 ;
      RECT 22.0240 7.8165 22.0500 8.9100 ;
      RECT 21.9160 7.8165 21.9420 8.9100 ;
      RECT 21.8080 7.8165 21.8340 8.9100 ;
      RECT 21.7000 7.8165 21.7260 8.9100 ;
      RECT 21.5920 7.8165 21.6180 8.9100 ;
      RECT 21.4840 7.8165 21.5100 8.9100 ;
      RECT 21.3760 7.8165 21.4020 8.9100 ;
      RECT 21.2680 7.8165 21.2940 8.9100 ;
      RECT 21.1600 7.8165 21.1860 8.9100 ;
      RECT 21.0520 7.8165 21.0780 8.9100 ;
      RECT 20.9440 7.8165 20.9700 8.9100 ;
      RECT 20.8360 7.8165 20.8620 8.9100 ;
      RECT 20.7280 7.8165 20.7540 8.9100 ;
      RECT 20.6200 7.8165 20.6460 8.9100 ;
      RECT 20.5120 7.8165 20.5380 8.9100 ;
      RECT 20.4040 7.8165 20.4300 8.9100 ;
      RECT 20.2960 7.8165 20.3220 8.9100 ;
      RECT 20.1880 7.8165 20.2140 8.9100 ;
      RECT 20.0800 7.8165 20.1060 8.9100 ;
      RECT 19.9720 7.8165 19.9980 8.9100 ;
      RECT 19.8640 7.8165 19.8900 8.9100 ;
      RECT 19.7560 7.8165 19.7820 8.9100 ;
      RECT 19.6480 7.8165 19.6740 8.9100 ;
      RECT 19.5400 7.8165 19.5660 8.9100 ;
      RECT 19.4320 7.8165 19.4580 8.9100 ;
      RECT 19.3240 7.8165 19.3500 8.9100 ;
      RECT 19.2160 7.8165 19.2420 8.9100 ;
      RECT 19.1080 7.8165 19.1340 8.9100 ;
      RECT 19.0000 7.8165 19.0260 8.9100 ;
      RECT 18.8920 7.8165 18.9180 8.9100 ;
      RECT 18.7840 7.8165 18.8100 8.9100 ;
      RECT 18.6760 7.8165 18.7020 8.9100 ;
      RECT 18.5680 7.8165 18.5940 8.9100 ;
      RECT 18.4600 7.8165 18.4860 8.9100 ;
      RECT 18.3520 7.8165 18.3780 8.9100 ;
      RECT 18.2440 7.8165 18.2700 8.9100 ;
      RECT 18.1360 7.8165 18.1620 8.9100 ;
      RECT 18.0280 7.8165 18.0540 8.9100 ;
      RECT 17.9200 7.8165 17.9460 8.9100 ;
      RECT 17.8120 7.8165 17.8380 8.9100 ;
      RECT 17.7040 7.8165 17.7300 8.9100 ;
      RECT 17.5960 7.8165 17.6220 8.9100 ;
      RECT 17.4880 7.8165 17.5140 8.9100 ;
      RECT 17.3800 7.8165 17.4060 8.9100 ;
      RECT 17.2720 7.8165 17.2980 8.9100 ;
      RECT 17.1640 7.8165 17.1900 8.9100 ;
      RECT 17.0560 7.8165 17.0820 8.9100 ;
      RECT 16.9480 7.8165 16.9740 8.9100 ;
      RECT 16.8400 7.8165 16.8660 8.9100 ;
      RECT 16.7320 7.8165 16.7580 8.9100 ;
      RECT 16.6240 7.8165 16.6500 8.9100 ;
      RECT 16.5160 7.8165 16.5420 8.9100 ;
      RECT 16.4080 7.8165 16.4340 8.9100 ;
      RECT 16.3000 7.8165 16.3260 8.9100 ;
      RECT 16.0870 7.8165 16.1640 8.9100 ;
      RECT 14.1940 7.8165 14.2710 8.9100 ;
      RECT 14.0320 7.8165 14.0580 8.9100 ;
      RECT 13.9240 7.8165 13.9500 8.9100 ;
      RECT 13.8160 7.8165 13.8420 8.9100 ;
      RECT 13.7080 7.8165 13.7340 8.9100 ;
      RECT 13.6000 7.8165 13.6260 8.9100 ;
      RECT 13.4920 7.8165 13.5180 8.9100 ;
      RECT 13.3840 7.8165 13.4100 8.9100 ;
      RECT 13.2760 7.8165 13.3020 8.9100 ;
      RECT 13.1680 7.8165 13.1940 8.9100 ;
      RECT 13.0600 7.8165 13.0860 8.9100 ;
      RECT 12.9520 7.8165 12.9780 8.9100 ;
      RECT 12.8440 7.8165 12.8700 8.9100 ;
      RECT 12.7360 7.8165 12.7620 8.9100 ;
      RECT 12.6280 7.8165 12.6540 8.9100 ;
      RECT 12.5200 7.8165 12.5460 8.9100 ;
      RECT 12.4120 7.8165 12.4380 8.9100 ;
      RECT 12.3040 7.8165 12.3300 8.9100 ;
      RECT 12.1960 7.8165 12.2220 8.9100 ;
      RECT 12.0880 7.8165 12.1140 8.9100 ;
      RECT 11.9800 7.8165 12.0060 8.9100 ;
      RECT 11.8720 7.8165 11.8980 8.9100 ;
      RECT 11.7640 7.8165 11.7900 8.9100 ;
      RECT 11.6560 7.8165 11.6820 8.9100 ;
      RECT 11.5480 7.8165 11.5740 8.9100 ;
      RECT 11.4400 7.8165 11.4660 8.9100 ;
      RECT 11.3320 7.8165 11.3580 8.9100 ;
      RECT 11.2240 7.8165 11.2500 8.9100 ;
      RECT 11.1160 7.8165 11.1420 8.9100 ;
      RECT 11.0080 7.8165 11.0340 8.9100 ;
      RECT 10.9000 7.8165 10.9260 8.9100 ;
      RECT 10.7920 7.8165 10.8180 8.9100 ;
      RECT 10.6840 7.8165 10.7100 8.9100 ;
      RECT 10.5760 7.8165 10.6020 8.9100 ;
      RECT 10.4680 7.8165 10.4940 8.9100 ;
      RECT 10.3600 7.8165 10.3860 8.9100 ;
      RECT 10.2520 7.8165 10.2780 8.9100 ;
      RECT 10.1440 7.8165 10.1700 8.9100 ;
      RECT 10.0360 7.8165 10.0620 8.9100 ;
      RECT 9.9280 7.8165 9.9540 8.9100 ;
      RECT 9.8200 7.8165 9.8460 8.9100 ;
      RECT 9.7120 7.8165 9.7380 8.9100 ;
      RECT 9.6040 7.8165 9.6300 8.9100 ;
      RECT 9.4960 7.8165 9.5220 8.9100 ;
      RECT 9.3880 7.8165 9.4140 8.9100 ;
      RECT 9.2800 7.8165 9.3060 8.9100 ;
      RECT 9.1720 7.8165 9.1980 8.9100 ;
      RECT 9.0640 7.8165 9.0900 8.9100 ;
      RECT 8.9560 7.8165 8.9820 8.9100 ;
      RECT 8.8480 7.8165 8.8740 8.9100 ;
      RECT 8.7400 7.8165 8.7660 8.9100 ;
      RECT 8.6320 7.8165 8.6580 8.9100 ;
      RECT 8.5240 7.8165 8.5500 8.9100 ;
      RECT 8.4160 7.8165 8.4420 8.9100 ;
      RECT 8.3080 7.8165 8.3340 8.9100 ;
      RECT 8.2000 7.8165 8.2260 8.9100 ;
      RECT 8.0920 7.8165 8.1180 8.9100 ;
      RECT 7.9840 7.8165 8.0100 8.9100 ;
      RECT 7.8760 7.8165 7.9020 8.9100 ;
      RECT 7.7680 7.8165 7.7940 8.9100 ;
      RECT 7.6600 7.8165 7.6860 8.9100 ;
      RECT 7.5520 7.8165 7.5780 8.9100 ;
      RECT 7.4440 7.8165 7.4700 8.9100 ;
      RECT 7.3360 7.8165 7.3620 8.9100 ;
      RECT 7.2280 7.8165 7.2540 8.9100 ;
      RECT 7.1200 7.8165 7.1460 8.9100 ;
      RECT 7.0120 7.8165 7.0380 8.9100 ;
      RECT 6.9040 7.8165 6.9300 8.9100 ;
      RECT 6.7960 7.8165 6.8220 8.9100 ;
      RECT 6.6880 7.8165 6.7140 8.9100 ;
      RECT 6.5800 7.8165 6.6060 8.9100 ;
      RECT 6.4720 7.8165 6.4980 8.9100 ;
      RECT 6.3640 7.8165 6.3900 8.9100 ;
      RECT 6.2560 7.8165 6.2820 8.9100 ;
      RECT 6.1480 7.8165 6.1740 8.9100 ;
      RECT 6.0400 7.8165 6.0660 8.9100 ;
      RECT 5.9320 7.8165 5.9580 8.9100 ;
      RECT 5.8240 7.8165 5.8500 8.9100 ;
      RECT 5.7160 7.8165 5.7420 8.9100 ;
      RECT 5.6080 7.8165 5.6340 8.9100 ;
      RECT 5.5000 7.8165 5.5260 8.9100 ;
      RECT 5.3920 7.8165 5.4180 8.9100 ;
      RECT 5.2840 7.8165 5.3100 8.9100 ;
      RECT 5.1760 7.8165 5.2020 8.9100 ;
      RECT 5.0680 7.8165 5.0940 8.9100 ;
      RECT 4.9600 7.8165 4.9860 8.9100 ;
      RECT 4.8520 7.8165 4.8780 8.9100 ;
      RECT 4.7440 7.8165 4.7700 8.9100 ;
      RECT 4.6360 7.8165 4.6620 8.9100 ;
      RECT 4.5280 7.8165 4.5540 8.9100 ;
      RECT 4.4200 7.8165 4.4460 8.9100 ;
      RECT 4.3120 7.8165 4.3380 8.9100 ;
      RECT 4.2040 7.8165 4.2300 8.9100 ;
      RECT 4.0960 7.8165 4.1220 8.9100 ;
      RECT 3.9880 7.8165 4.0140 8.9100 ;
      RECT 3.8800 7.8165 3.9060 8.9100 ;
      RECT 3.7720 7.8165 3.7980 8.9100 ;
      RECT 3.6640 7.8165 3.6900 8.9100 ;
      RECT 3.5560 7.8165 3.5820 8.9100 ;
      RECT 3.4480 7.8165 3.4740 8.9100 ;
      RECT 3.3400 7.8165 3.3660 8.9100 ;
      RECT 3.2320 7.8165 3.2580 8.9100 ;
      RECT 3.1240 7.8165 3.1500 8.9100 ;
      RECT 3.0160 7.8165 3.0420 8.9100 ;
      RECT 2.9080 7.8165 2.9340 8.9100 ;
      RECT 2.8000 7.8165 2.8260 8.9100 ;
      RECT 2.6920 7.8165 2.7180 8.9100 ;
      RECT 2.5840 7.8165 2.6100 8.9100 ;
      RECT 2.4760 7.8165 2.5020 8.9100 ;
      RECT 2.3680 7.8165 2.3940 8.9100 ;
      RECT 2.2600 7.8165 2.2860 8.9100 ;
      RECT 2.1520 7.8165 2.1780 8.9100 ;
      RECT 2.0440 7.8165 2.0700 8.9100 ;
      RECT 1.9360 7.8165 1.9620 8.9100 ;
      RECT 1.8280 7.8165 1.8540 8.9100 ;
      RECT 1.7200 7.8165 1.7460 8.9100 ;
      RECT 1.6120 7.8165 1.6380 8.9100 ;
      RECT 1.5040 7.8165 1.5300 8.9100 ;
      RECT 1.3960 7.8165 1.4220 8.9100 ;
      RECT 1.2880 7.8165 1.3140 8.9100 ;
      RECT 1.1800 7.8165 1.2060 8.9100 ;
      RECT 1.0720 7.8165 1.0980 8.9100 ;
      RECT 0.9640 7.8165 0.9900 8.9100 ;
      RECT 0.8560 7.8165 0.8820 8.9100 ;
      RECT 0.7480 7.8165 0.7740 8.9100 ;
      RECT 0.6400 7.8165 0.6660 8.9100 ;
      RECT 0.5320 7.8165 0.5580 8.9100 ;
      RECT 0.4240 7.8165 0.4500 8.9100 ;
      RECT 0.3160 7.8165 0.3420 8.9100 ;
      RECT 0.2080 7.8165 0.2340 8.9100 ;
      RECT 0.0050 7.8165 0.0900 8.9100 ;
      RECT 15.5530 8.8965 15.6810 9.9900 ;
      RECT 15.5390 9.5620 15.6810 9.8845 ;
      RECT 15.3190 9.2890 15.4530 9.9900 ;
      RECT 15.2960 9.6240 15.4530 9.8820 ;
      RECT 15.3190 8.8965 15.4170 9.9900 ;
      RECT 15.3190 9.0175 15.4310 9.2570 ;
      RECT 15.3190 8.8965 15.4530 8.9855 ;
      RECT 15.0940 9.3470 15.2280 9.9900 ;
      RECT 15.0940 8.8965 15.1920 9.9900 ;
      RECT 14.6770 8.8965 14.7600 9.9900 ;
      RECT 14.6770 8.9850 14.7740 9.9205 ;
      RECT 30.2680 8.8965 30.3530 9.9900 ;
      RECT 30.1240 8.8965 30.1500 9.9900 ;
      RECT 30.0160 8.8965 30.0420 9.9900 ;
      RECT 29.9080 8.8965 29.9340 9.9900 ;
      RECT 29.8000 8.8965 29.8260 9.9900 ;
      RECT 29.6920 8.8965 29.7180 9.9900 ;
      RECT 29.5840 8.8965 29.6100 9.9900 ;
      RECT 29.4760 8.8965 29.5020 9.9900 ;
      RECT 29.3680 8.8965 29.3940 9.9900 ;
      RECT 29.2600 8.8965 29.2860 9.9900 ;
      RECT 29.1520 8.8965 29.1780 9.9900 ;
      RECT 29.0440 8.8965 29.0700 9.9900 ;
      RECT 28.9360 8.8965 28.9620 9.9900 ;
      RECT 28.8280 8.8965 28.8540 9.9900 ;
      RECT 28.7200 8.8965 28.7460 9.9900 ;
      RECT 28.6120 8.8965 28.6380 9.9900 ;
      RECT 28.5040 8.8965 28.5300 9.9900 ;
      RECT 28.3960 8.8965 28.4220 9.9900 ;
      RECT 28.2880 8.8965 28.3140 9.9900 ;
      RECT 28.1800 8.8965 28.2060 9.9900 ;
      RECT 28.0720 8.8965 28.0980 9.9900 ;
      RECT 27.9640 8.8965 27.9900 9.9900 ;
      RECT 27.8560 8.8965 27.8820 9.9900 ;
      RECT 27.7480 8.8965 27.7740 9.9900 ;
      RECT 27.6400 8.8965 27.6660 9.9900 ;
      RECT 27.5320 8.8965 27.5580 9.9900 ;
      RECT 27.4240 8.8965 27.4500 9.9900 ;
      RECT 27.3160 8.8965 27.3420 9.9900 ;
      RECT 27.2080 8.8965 27.2340 9.9900 ;
      RECT 27.1000 8.8965 27.1260 9.9900 ;
      RECT 26.9920 8.8965 27.0180 9.9900 ;
      RECT 26.8840 8.8965 26.9100 9.9900 ;
      RECT 26.7760 8.8965 26.8020 9.9900 ;
      RECT 26.6680 8.8965 26.6940 9.9900 ;
      RECT 26.5600 8.8965 26.5860 9.9900 ;
      RECT 26.4520 8.8965 26.4780 9.9900 ;
      RECT 26.3440 8.8965 26.3700 9.9900 ;
      RECT 26.2360 8.8965 26.2620 9.9900 ;
      RECT 26.1280 8.8965 26.1540 9.9900 ;
      RECT 26.0200 8.8965 26.0460 9.9900 ;
      RECT 25.9120 8.8965 25.9380 9.9900 ;
      RECT 25.8040 8.8965 25.8300 9.9900 ;
      RECT 25.6960 8.8965 25.7220 9.9900 ;
      RECT 25.5880 8.8965 25.6140 9.9900 ;
      RECT 25.4800 8.8965 25.5060 9.9900 ;
      RECT 25.3720 8.8965 25.3980 9.9900 ;
      RECT 25.2640 8.8965 25.2900 9.9900 ;
      RECT 25.1560 8.8965 25.1820 9.9900 ;
      RECT 25.0480 8.8965 25.0740 9.9900 ;
      RECT 24.9400 8.8965 24.9660 9.9900 ;
      RECT 24.8320 8.8965 24.8580 9.9900 ;
      RECT 24.7240 8.8965 24.7500 9.9900 ;
      RECT 24.6160 8.8965 24.6420 9.9900 ;
      RECT 24.5080 8.8965 24.5340 9.9900 ;
      RECT 24.4000 8.8965 24.4260 9.9900 ;
      RECT 24.2920 8.8965 24.3180 9.9900 ;
      RECT 24.1840 8.8965 24.2100 9.9900 ;
      RECT 24.0760 8.8965 24.1020 9.9900 ;
      RECT 23.9680 8.8965 23.9940 9.9900 ;
      RECT 23.8600 8.8965 23.8860 9.9900 ;
      RECT 23.7520 8.8965 23.7780 9.9900 ;
      RECT 23.6440 8.8965 23.6700 9.9900 ;
      RECT 23.5360 8.8965 23.5620 9.9900 ;
      RECT 23.4280 8.8965 23.4540 9.9900 ;
      RECT 23.3200 8.8965 23.3460 9.9900 ;
      RECT 23.2120 8.8965 23.2380 9.9900 ;
      RECT 23.1040 8.8965 23.1300 9.9900 ;
      RECT 22.9960 8.8965 23.0220 9.9900 ;
      RECT 22.8880 8.8965 22.9140 9.9900 ;
      RECT 22.7800 8.8965 22.8060 9.9900 ;
      RECT 22.6720 8.8965 22.6980 9.9900 ;
      RECT 22.5640 8.8965 22.5900 9.9900 ;
      RECT 22.4560 8.8965 22.4820 9.9900 ;
      RECT 22.3480 8.8965 22.3740 9.9900 ;
      RECT 22.2400 8.8965 22.2660 9.9900 ;
      RECT 22.1320 8.8965 22.1580 9.9900 ;
      RECT 22.0240 8.8965 22.0500 9.9900 ;
      RECT 21.9160 8.8965 21.9420 9.9900 ;
      RECT 21.8080 8.8965 21.8340 9.9900 ;
      RECT 21.7000 8.8965 21.7260 9.9900 ;
      RECT 21.5920 8.8965 21.6180 9.9900 ;
      RECT 21.4840 8.8965 21.5100 9.9900 ;
      RECT 21.3760 8.8965 21.4020 9.9900 ;
      RECT 21.2680 8.8965 21.2940 9.9900 ;
      RECT 21.1600 8.8965 21.1860 9.9900 ;
      RECT 21.0520 8.8965 21.0780 9.9900 ;
      RECT 20.9440 8.8965 20.9700 9.9900 ;
      RECT 20.8360 8.8965 20.8620 9.9900 ;
      RECT 20.7280 8.8965 20.7540 9.9900 ;
      RECT 20.6200 8.8965 20.6460 9.9900 ;
      RECT 20.5120 8.8965 20.5380 9.9900 ;
      RECT 20.4040 8.8965 20.4300 9.9900 ;
      RECT 20.2960 8.8965 20.3220 9.9900 ;
      RECT 20.1880 8.8965 20.2140 9.9900 ;
      RECT 20.0800 8.8965 20.1060 9.9900 ;
      RECT 19.9720 8.8965 19.9980 9.9900 ;
      RECT 19.8640 8.8965 19.8900 9.9900 ;
      RECT 19.7560 8.8965 19.7820 9.9900 ;
      RECT 19.6480 8.8965 19.6740 9.9900 ;
      RECT 19.5400 8.8965 19.5660 9.9900 ;
      RECT 19.4320 8.8965 19.4580 9.9900 ;
      RECT 19.3240 8.8965 19.3500 9.9900 ;
      RECT 19.2160 8.8965 19.2420 9.9900 ;
      RECT 19.1080 8.8965 19.1340 9.9900 ;
      RECT 19.0000 8.8965 19.0260 9.9900 ;
      RECT 18.8920 8.8965 18.9180 9.9900 ;
      RECT 18.7840 8.8965 18.8100 9.9900 ;
      RECT 18.6760 8.8965 18.7020 9.9900 ;
      RECT 18.5680 8.8965 18.5940 9.9900 ;
      RECT 18.4600 8.8965 18.4860 9.9900 ;
      RECT 18.3520 8.8965 18.3780 9.9900 ;
      RECT 18.2440 8.8965 18.2700 9.9900 ;
      RECT 18.1360 8.8965 18.1620 9.9900 ;
      RECT 18.0280 8.8965 18.0540 9.9900 ;
      RECT 17.9200 8.8965 17.9460 9.9900 ;
      RECT 17.8120 8.8965 17.8380 9.9900 ;
      RECT 17.7040 8.8965 17.7300 9.9900 ;
      RECT 17.5960 8.8965 17.6220 9.9900 ;
      RECT 17.4880 8.8965 17.5140 9.9900 ;
      RECT 17.3800 8.8965 17.4060 9.9900 ;
      RECT 17.2720 8.8965 17.2980 9.9900 ;
      RECT 17.1640 8.8965 17.1900 9.9900 ;
      RECT 17.0560 8.8965 17.0820 9.9900 ;
      RECT 16.9480 8.8965 16.9740 9.9900 ;
      RECT 16.8400 8.8965 16.8660 9.9900 ;
      RECT 16.7320 8.8965 16.7580 9.9900 ;
      RECT 16.6240 8.8965 16.6500 9.9900 ;
      RECT 16.5160 8.8965 16.5420 9.9900 ;
      RECT 16.4080 8.8965 16.4340 9.9900 ;
      RECT 16.3000 8.8965 16.3260 9.9900 ;
      RECT 16.0870 8.8965 16.1640 9.9900 ;
      RECT 14.1940 8.8965 14.2710 9.9900 ;
      RECT 14.0320 8.8965 14.0580 9.9900 ;
      RECT 13.9240 8.8965 13.9500 9.9900 ;
      RECT 13.8160 8.8965 13.8420 9.9900 ;
      RECT 13.7080 8.8965 13.7340 9.9900 ;
      RECT 13.6000 8.8965 13.6260 9.9900 ;
      RECT 13.4920 8.8965 13.5180 9.9900 ;
      RECT 13.3840 8.8965 13.4100 9.9900 ;
      RECT 13.2760 8.8965 13.3020 9.9900 ;
      RECT 13.1680 8.8965 13.1940 9.9900 ;
      RECT 13.0600 8.8965 13.0860 9.9900 ;
      RECT 12.9520 8.8965 12.9780 9.9900 ;
      RECT 12.8440 8.8965 12.8700 9.9900 ;
      RECT 12.7360 8.8965 12.7620 9.9900 ;
      RECT 12.6280 8.8965 12.6540 9.9900 ;
      RECT 12.5200 8.8965 12.5460 9.9900 ;
      RECT 12.4120 8.8965 12.4380 9.9900 ;
      RECT 12.3040 8.8965 12.3300 9.9900 ;
      RECT 12.1960 8.8965 12.2220 9.9900 ;
      RECT 12.0880 8.8965 12.1140 9.9900 ;
      RECT 11.9800 8.8965 12.0060 9.9900 ;
      RECT 11.8720 8.8965 11.8980 9.9900 ;
      RECT 11.7640 8.8965 11.7900 9.9900 ;
      RECT 11.6560 8.8965 11.6820 9.9900 ;
      RECT 11.5480 8.8965 11.5740 9.9900 ;
      RECT 11.4400 8.8965 11.4660 9.9900 ;
      RECT 11.3320 8.8965 11.3580 9.9900 ;
      RECT 11.2240 8.8965 11.2500 9.9900 ;
      RECT 11.1160 8.8965 11.1420 9.9900 ;
      RECT 11.0080 8.8965 11.0340 9.9900 ;
      RECT 10.9000 8.8965 10.9260 9.9900 ;
      RECT 10.7920 8.8965 10.8180 9.9900 ;
      RECT 10.6840 8.8965 10.7100 9.9900 ;
      RECT 10.5760 8.8965 10.6020 9.9900 ;
      RECT 10.4680 8.8965 10.4940 9.9900 ;
      RECT 10.3600 8.8965 10.3860 9.9900 ;
      RECT 10.2520 8.8965 10.2780 9.9900 ;
      RECT 10.1440 8.8965 10.1700 9.9900 ;
      RECT 10.0360 8.8965 10.0620 9.9900 ;
      RECT 9.9280 8.8965 9.9540 9.9900 ;
      RECT 9.8200 8.8965 9.8460 9.9900 ;
      RECT 9.7120 8.8965 9.7380 9.9900 ;
      RECT 9.6040 8.8965 9.6300 9.9900 ;
      RECT 9.4960 8.8965 9.5220 9.9900 ;
      RECT 9.3880 8.8965 9.4140 9.9900 ;
      RECT 9.2800 8.8965 9.3060 9.9900 ;
      RECT 9.1720 8.8965 9.1980 9.9900 ;
      RECT 9.0640 8.8965 9.0900 9.9900 ;
      RECT 8.9560 8.8965 8.9820 9.9900 ;
      RECT 8.8480 8.8965 8.8740 9.9900 ;
      RECT 8.7400 8.8965 8.7660 9.9900 ;
      RECT 8.6320 8.8965 8.6580 9.9900 ;
      RECT 8.5240 8.8965 8.5500 9.9900 ;
      RECT 8.4160 8.8965 8.4420 9.9900 ;
      RECT 8.3080 8.8965 8.3340 9.9900 ;
      RECT 8.2000 8.8965 8.2260 9.9900 ;
      RECT 8.0920 8.8965 8.1180 9.9900 ;
      RECT 7.9840 8.8965 8.0100 9.9900 ;
      RECT 7.8760 8.8965 7.9020 9.9900 ;
      RECT 7.7680 8.8965 7.7940 9.9900 ;
      RECT 7.6600 8.8965 7.6860 9.9900 ;
      RECT 7.5520 8.8965 7.5780 9.9900 ;
      RECT 7.4440 8.8965 7.4700 9.9900 ;
      RECT 7.3360 8.8965 7.3620 9.9900 ;
      RECT 7.2280 8.8965 7.2540 9.9900 ;
      RECT 7.1200 8.8965 7.1460 9.9900 ;
      RECT 7.0120 8.8965 7.0380 9.9900 ;
      RECT 6.9040 8.8965 6.9300 9.9900 ;
      RECT 6.7960 8.8965 6.8220 9.9900 ;
      RECT 6.6880 8.8965 6.7140 9.9900 ;
      RECT 6.5800 8.8965 6.6060 9.9900 ;
      RECT 6.4720 8.8965 6.4980 9.9900 ;
      RECT 6.3640 8.8965 6.3900 9.9900 ;
      RECT 6.2560 8.8965 6.2820 9.9900 ;
      RECT 6.1480 8.8965 6.1740 9.9900 ;
      RECT 6.0400 8.8965 6.0660 9.9900 ;
      RECT 5.9320 8.8965 5.9580 9.9900 ;
      RECT 5.8240 8.8965 5.8500 9.9900 ;
      RECT 5.7160 8.8965 5.7420 9.9900 ;
      RECT 5.6080 8.8965 5.6340 9.9900 ;
      RECT 5.5000 8.8965 5.5260 9.9900 ;
      RECT 5.3920 8.8965 5.4180 9.9900 ;
      RECT 5.2840 8.8965 5.3100 9.9900 ;
      RECT 5.1760 8.8965 5.2020 9.9900 ;
      RECT 5.0680 8.8965 5.0940 9.9900 ;
      RECT 4.9600 8.8965 4.9860 9.9900 ;
      RECT 4.8520 8.8965 4.8780 9.9900 ;
      RECT 4.7440 8.8965 4.7700 9.9900 ;
      RECT 4.6360 8.8965 4.6620 9.9900 ;
      RECT 4.5280 8.8965 4.5540 9.9900 ;
      RECT 4.4200 8.8965 4.4460 9.9900 ;
      RECT 4.3120 8.8965 4.3380 9.9900 ;
      RECT 4.2040 8.8965 4.2300 9.9900 ;
      RECT 4.0960 8.8965 4.1220 9.9900 ;
      RECT 3.9880 8.8965 4.0140 9.9900 ;
      RECT 3.8800 8.8965 3.9060 9.9900 ;
      RECT 3.7720 8.8965 3.7980 9.9900 ;
      RECT 3.6640 8.8965 3.6900 9.9900 ;
      RECT 3.5560 8.8965 3.5820 9.9900 ;
      RECT 3.4480 8.8965 3.4740 9.9900 ;
      RECT 3.3400 8.8965 3.3660 9.9900 ;
      RECT 3.2320 8.8965 3.2580 9.9900 ;
      RECT 3.1240 8.8965 3.1500 9.9900 ;
      RECT 3.0160 8.8965 3.0420 9.9900 ;
      RECT 2.9080 8.8965 2.9340 9.9900 ;
      RECT 2.8000 8.8965 2.8260 9.9900 ;
      RECT 2.6920 8.8965 2.7180 9.9900 ;
      RECT 2.5840 8.8965 2.6100 9.9900 ;
      RECT 2.4760 8.8965 2.5020 9.9900 ;
      RECT 2.3680 8.8965 2.3940 9.9900 ;
      RECT 2.2600 8.8965 2.2860 9.9900 ;
      RECT 2.1520 8.8965 2.1780 9.9900 ;
      RECT 2.0440 8.8965 2.0700 9.9900 ;
      RECT 1.9360 8.8965 1.9620 9.9900 ;
      RECT 1.8280 8.8965 1.8540 9.9900 ;
      RECT 1.7200 8.8965 1.7460 9.9900 ;
      RECT 1.6120 8.8965 1.6380 9.9900 ;
      RECT 1.5040 8.8965 1.5300 9.9900 ;
      RECT 1.3960 8.8965 1.4220 9.9900 ;
      RECT 1.2880 8.8965 1.3140 9.9900 ;
      RECT 1.1800 8.8965 1.2060 9.9900 ;
      RECT 1.0720 8.8965 1.0980 9.9900 ;
      RECT 0.9640 8.8965 0.9900 9.9900 ;
      RECT 0.8560 8.8965 0.8820 9.9900 ;
      RECT 0.7480 8.8965 0.7740 9.9900 ;
      RECT 0.6400 8.8965 0.6660 9.9900 ;
      RECT 0.5320 8.8965 0.5580 9.9900 ;
      RECT 0.4240 8.8965 0.4500 9.9900 ;
      RECT 0.3160 8.8965 0.3420 9.9900 ;
      RECT 0.2080 8.8965 0.2340 9.9900 ;
      RECT 0.0050 8.8965 0.0900 9.9900 ;
      RECT 15.5530 9.9765 15.6810 11.0700 ;
      RECT 15.5390 10.6420 15.6810 10.9645 ;
      RECT 15.3190 10.3690 15.4530 11.0700 ;
      RECT 15.2960 10.7040 15.4530 10.9620 ;
      RECT 15.3190 9.9765 15.4170 11.0700 ;
      RECT 15.3190 10.0975 15.4310 10.3370 ;
      RECT 15.3190 9.9765 15.4530 10.0655 ;
      RECT 15.0940 10.4270 15.2280 11.0700 ;
      RECT 15.0940 9.9765 15.1920 11.0700 ;
      RECT 14.6770 9.9765 14.7600 11.0700 ;
      RECT 14.6770 10.0650 14.7740 11.0005 ;
      RECT 30.2680 9.9765 30.3530 11.0700 ;
      RECT 30.1240 9.9765 30.1500 11.0700 ;
      RECT 30.0160 9.9765 30.0420 11.0700 ;
      RECT 29.9080 9.9765 29.9340 11.0700 ;
      RECT 29.8000 9.9765 29.8260 11.0700 ;
      RECT 29.6920 9.9765 29.7180 11.0700 ;
      RECT 29.5840 9.9765 29.6100 11.0700 ;
      RECT 29.4760 9.9765 29.5020 11.0700 ;
      RECT 29.3680 9.9765 29.3940 11.0700 ;
      RECT 29.2600 9.9765 29.2860 11.0700 ;
      RECT 29.1520 9.9765 29.1780 11.0700 ;
      RECT 29.0440 9.9765 29.0700 11.0700 ;
      RECT 28.9360 9.9765 28.9620 11.0700 ;
      RECT 28.8280 9.9765 28.8540 11.0700 ;
      RECT 28.7200 9.9765 28.7460 11.0700 ;
      RECT 28.6120 9.9765 28.6380 11.0700 ;
      RECT 28.5040 9.9765 28.5300 11.0700 ;
      RECT 28.3960 9.9765 28.4220 11.0700 ;
      RECT 28.2880 9.9765 28.3140 11.0700 ;
      RECT 28.1800 9.9765 28.2060 11.0700 ;
      RECT 28.0720 9.9765 28.0980 11.0700 ;
      RECT 27.9640 9.9765 27.9900 11.0700 ;
      RECT 27.8560 9.9765 27.8820 11.0700 ;
      RECT 27.7480 9.9765 27.7740 11.0700 ;
      RECT 27.6400 9.9765 27.6660 11.0700 ;
      RECT 27.5320 9.9765 27.5580 11.0700 ;
      RECT 27.4240 9.9765 27.4500 11.0700 ;
      RECT 27.3160 9.9765 27.3420 11.0700 ;
      RECT 27.2080 9.9765 27.2340 11.0700 ;
      RECT 27.1000 9.9765 27.1260 11.0700 ;
      RECT 26.9920 9.9765 27.0180 11.0700 ;
      RECT 26.8840 9.9765 26.9100 11.0700 ;
      RECT 26.7760 9.9765 26.8020 11.0700 ;
      RECT 26.6680 9.9765 26.6940 11.0700 ;
      RECT 26.5600 9.9765 26.5860 11.0700 ;
      RECT 26.4520 9.9765 26.4780 11.0700 ;
      RECT 26.3440 9.9765 26.3700 11.0700 ;
      RECT 26.2360 9.9765 26.2620 11.0700 ;
      RECT 26.1280 9.9765 26.1540 11.0700 ;
      RECT 26.0200 9.9765 26.0460 11.0700 ;
      RECT 25.9120 9.9765 25.9380 11.0700 ;
      RECT 25.8040 9.9765 25.8300 11.0700 ;
      RECT 25.6960 9.9765 25.7220 11.0700 ;
      RECT 25.5880 9.9765 25.6140 11.0700 ;
      RECT 25.4800 9.9765 25.5060 11.0700 ;
      RECT 25.3720 9.9765 25.3980 11.0700 ;
      RECT 25.2640 9.9765 25.2900 11.0700 ;
      RECT 25.1560 9.9765 25.1820 11.0700 ;
      RECT 25.0480 9.9765 25.0740 11.0700 ;
      RECT 24.9400 9.9765 24.9660 11.0700 ;
      RECT 24.8320 9.9765 24.8580 11.0700 ;
      RECT 24.7240 9.9765 24.7500 11.0700 ;
      RECT 24.6160 9.9765 24.6420 11.0700 ;
      RECT 24.5080 9.9765 24.5340 11.0700 ;
      RECT 24.4000 9.9765 24.4260 11.0700 ;
      RECT 24.2920 9.9765 24.3180 11.0700 ;
      RECT 24.1840 9.9765 24.2100 11.0700 ;
      RECT 24.0760 9.9765 24.1020 11.0700 ;
      RECT 23.9680 9.9765 23.9940 11.0700 ;
      RECT 23.8600 9.9765 23.8860 11.0700 ;
      RECT 23.7520 9.9765 23.7780 11.0700 ;
      RECT 23.6440 9.9765 23.6700 11.0700 ;
      RECT 23.5360 9.9765 23.5620 11.0700 ;
      RECT 23.4280 9.9765 23.4540 11.0700 ;
      RECT 23.3200 9.9765 23.3460 11.0700 ;
      RECT 23.2120 9.9765 23.2380 11.0700 ;
      RECT 23.1040 9.9765 23.1300 11.0700 ;
      RECT 22.9960 9.9765 23.0220 11.0700 ;
      RECT 22.8880 9.9765 22.9140 11.0700 ;
      RECT 22.7800 9.9765 22.8060 11.0700 ;
      RECT 22.6720 9.9765 22.6980 11.0700 ;
      RECT 22.5640 9.9765 22.5900 11.0700 ;
      RECT 22.4560 9.9765 22.4820 11.0700 ;
      RECT 22.3480 9.9765 22.3740 11.0700 ;
      RECT 22.2400 9.9765 22.2660 11.0700 ;
      RECT 22.1320 9.9765 22.1580 11.0700 ;
      RECT 22.0240 9.9765 22.0500 11.0700 ;
      RECT 21.9160 9.9765 21.9420 11.0700 ;
      RECT 21.8080 9.9765 21.8340 11.0700 ;
      RECT 21.7000 9.9765 21.7260 11.0700 ;
      RECT 21.5920 9.9765 21.6180 11.0700 ;
      RECT 21.4840 9.9765 21.5100 11.0700 ;
      RECT 21.3760 9.9765 21.4020 11.0700 ;
      RECT 21.2680 9.9765 21.2940 11.0700 ;
      RECT 21.1600 9.9765 21.1860 11.0700 ;
      RECT 21.0520 9.9765 21.0780 11.0700 ;
      RECT 20.9440 9.9765 20.9700 11.0700 ;
      RECT 20.8360 9.9765 20.8620 11.0700 ;
      RECT 20.7280 9.9765 20.7540 11.0700 ;
      RECT 20.6200 9.9765 20.6460 11.0700 ;
      RECT 20.5120 9.9765 20.5380 11.0700 ;
      RECT 20.4040 9.9765 20.4300 11.0700 ;
      RECT 20.2960 9.9765 20.3220 11.0700 ;
      RECT 20.1880 9.9765 20.2140 11.0700 ;
      RECT 20.0800 9.9765 20.1060 11.0700 ;
      RECT 19.9720 9.9765 19.9980 11.0700 ;
      RECT 19.8640 9.9765 19.8900 11.0700 ;
      RECT 19.7560 9.9765 19.7820 11.0700 ;
      RECT 19.6480 9.9765 19.6740 11.0700 ;
      RECT 19.5400 9.9765 19.5660 11.0700 ;
      RECT 19.4320 9.9765 19.4580 11.0700 ;
      RECT 19.3240 9.9765 19.3500 11.0700 ;
      RECT 19.2160 9.9765 19.2420 11.0700 ;
      RECT 19.1080 9.9765 19.1340 11.0700 ;
      RECT 19.0000 9.9765 19.0260 11.0700 ;
      RECT 18.8920 9.9765 18.9180 11.0700 ;
      RECT 18.7840 9.9765 18.8100 11.0700 ;
      RECT 18.6760 9.9765 18.7020 11.0700 ;
      RECT 18.5680 9.9765 18.5940 11.0700 ;
      RECT 18.4600 9.9765 18.4860 11.0700 ;
      RECT 18.3520 9.9765 18.3780 11.0700 ;
      RECT 18.2440 9.9765 18.2700 11.0700 ;
      RECT 18.1360 9.9765 18.1620 11.0700 ;
      RECT 18.0280 9.9765 18.0540 11.0700 ;
      RECT 17.9200 9.9765 17.9460 11.0700 ;
      RECT 17.8120 9.9765 17.8380 11.0700 ;
      RECT 17.7040 9.9765 17.7300 11.0700 ;
      RECT 17.5960 9.9765 17.6220 11.0700 ;
      RECT 17.4880 9.9765 17.5140 11.0700 ;
      RECT 17.3800 9.9765 17.4060 11.0700 ;
      RECT 17.2720 9.9765 17.2980 11.0700 ;
      RECT 17.1640 9.9765 17.1900 11.0700 ;
      RECT 17.0560 9.9765 17.0820 11.0700 ;
      RECT 16.9480 9.9765 16.9740 11.0700 ;
      RECT 16.8400 9.9765 16.8660 11.0700 ;
      RECT 16.7320 9.9765 16.7580 11.0700 ;
      RECT 16.6240 9.9765 16.6500 11.0700 ;
      RECT 16.5160 9.9765 16.5420 11.0700 ;
      RECT 16.4080 9.9765 16.4340 11.0700 ;
      RECT 16.3000 9.9765 16.3260 11.0700 ;
      RECT 16.0870 9.9765 16.1640 11.0700 ;
      RECT 14.1940 9.9765 14.2710 11.0700 ;
      RECT 14.0320 9.9765 14.0580 11.0700 ;
      RECT 13.9240 9.9765 13.9500 11.0700 ;
      RECT 13.8160 9.9765 13.8420 11.0700 ;
      RECT 13.7080 9.9765 13.7340 11.0700 ;
      RECT 13.6000 9.9765 13.6260 11.0700 ;
      RECT 13.4920 9.9765 13.5180 11.0700 ;
      RECT 13.3840 9.9765 13.4100 11.0700 ;
      RECT 13.2760 9.9765 13.3020 11.0700 ;
      RECT 13.1680 9.9765 13.1940 11.0700 ;
      RECT 13.0600 9.9765 13.0860 11.0700 ;
      RECT 12.9520 9.9765 12.9780 11.0700 ;
      RECT 12.8440 9.9765 12.8700 11.0700 ;
      RECT 12.7360 9.9765 12.7620 11.0700 ;
      RECT 12.6280 9.9765 12.6540 11.0700 ;
      RECT 12.5200 9.9765 12.5460 11.0700 ;
      RECT 12.4120 9.9765 12.4380 11.0700 ;
      RECT 12.3040 9.9765 12.3300 11.0700 ;
      RECT 12.1960 9.9765 12.2220 11.0700 ;
      RECT 12.0880 9.9765 12.1140 11.0700 ;
      RECT 11.9800 9.9765 12.0060 11.0700 ;
      RECT 11.8720 9.9765 11.8980 11.0700 ;
      RECT 11.7640 9.9765 11.7900 11.0700 ;
      RECT 11.6560 9.9765 11.6820 11.0700 ;
      RECT 11.5480 9.9765 11.5740 11.0700 ;
      RECT 11.4400 9.9765 11.4660 11.0700 ;
      RECT 11.3320 9.9765 11.3580 11.0700 ;
      RECT 11.2240 9.9765 11.2500 11.0700 ;
      RECT 11.1160 9.9765 11.1420 11.0700 ;
      RECT 11.0080 9.9765 11.0340 11.0700 ;
      RECT 10.9000 9.9765 10.9260 11.0700 ;
      RECT 10.7920 9.9765 10.8180 11.0700 ;
      RECT 10.6840 9.9765 10.7100 11.0700 ;
      RECT 10.5760 9.9765 10.6020 11.0700 ;
      RECT 10.4680 9.9765 10.4940 11.0700 ;
      RECT 10.3600 9.9765 10.3860 11.0700 ;
      RECT 10.2520 9.9765 10.2780 11.0700 ;
      RECT 10.1440 9.9765 10.1700 11.0700 ;
      RECT 10.0360 9.9765 10.0620 11.0700 ;
      RECT 9.9280 9.9765 9.9540 11.0700 ;
      RECT 9.8200 9.9765 9.8460 11.0700 ;
      RECT 9.7120 9.9765 9.7380 11.0700 ;
      RECT 9.6040 9.9765 9.6300 11.0700 ;
      RECT 9.4960 9.9765 9.5220 11.0700 ;
      RECT 9.3880 9.9765 9.4140 11.0700 ;
      RECT 9.2800 9.9765 9.3060 11.0700 ;
      RECT 9.1720 9.9765 9.1980 11.0700 ;
      RECT 9.0640 9.9765 9.0900 11.0700 ;
      RECT 8.9560 9.9765 8.9820 11.0700 ;
      RECT 8.8480 9.9765 8.8740 11.0700 ;
      RECT 8.7400 9.9765 8.7660 11.0700 ;
      RECT 8.6320 9.9765 8.6580 11.0700 ;
      RECT 8.5240 9.9765 8.5500 11.0700 ;
      RECT 8.4160 9.9765 8.4420 11.0700 ;
      RECT 8.3080 9.9765 8.3340 11.0700 ;
      RECT 8.2000 9.9765 8.2260 11.0700 ;
      RECT 8.0920 9.9765 8.1180 11.0700 ;
      RECT 7.9840 9.9765 8.0100 11.0700 ;
      RECT 7.8760 9.9765 7.9020 11.0700 ;
      RECT 7.7680 9.9765 7.7940 11.0700 ;
      RECT 7.6600 9.9765 7.6860 11.0700 ;
      RECT 7.5520 9.9765 7.5780 11.0700 ;
      RECT 7.4440 9.9765 7.4700 11.0700 ;
      RECT 7.3360 9.9765 7.3620 11.0700 ;
      RECT 7.2280 9.9765 7.2540 11.0700 ;
      RECT 7.1200 9.9765 7.1460 11.0700 ;
      RECT 7.0120 9.9765 7.0380 11.0700 ;
      RECT 6.9040 9.9765 6.9300 11.0700 ;
      RECT 6.7960 9.9765 6.8220 11.0700 ;
      RECT 6.6880 9.9765 6.7140 11.0700 ;
      RECT 6.5800 9.9765 6.6060 11.0700 ;
      RECT 6.4720 9.9765 6.4980 11.0700 ;
      RECT 6.3640 9.9765 6.3900 11.0700 ;
      RECT 6.2560 9.9765 6.2820 11.0700 ;
      RECT 6.1480 9.9765 6.1740 11.0700 ;
      RECT 6.0400 9.9765 6.0660 11.0700 ;
      RECT 5.9320 9.9765 5.9580 11.0700 ;
      RECT 5.8240 9.9765 5.8500 11.0700 ;
      RECT 5.7160 9.9765 5.7420 11.0700 ;
      RECT 5.6080 9.9765 5.6340 11.0700 ;
      RECT 5.5000 9.9765 5.5260 11.0700 ;
      RECT 5.3920 9.9765 5.4180 11.0700 ;
      RECT 5.2840 9.9765 5.3100 11.0700 ;
      RECT 5.1760 9.9765 5.2020 11.0700 ;
      RECT 5.0680 9.9765 5.0940 11.0700 ;
      RECT 4.9600 9.9765 4.9860 11.0700 ;
      RECT 4.8520 9.9765 4.8780 11.0700 ;
      RECT 4.7440 9.9765 4.7700 11.0700 ;
      RECT 4.6360 9.9765 4.6620 11.0700 ;
      RECT 4.5280 9.9765 4.5540 11.0700 ;
      RECT 4.4200 9.9765 4.4460 11.0700 ;
      RECT 4.3120 9.9765 4.3380 11.0700 ;
      RECT 4.2040 9.9765 4.2300 11.0700 ;
      RECT 4.0960 9.9765 4.1220 11.0700 ;
      RECT 3.9880 9.9765 4.0140 11.0700 ;
      RECT 3.8800 9.9765 3.9060 11.0700 ;
      RECT 3.7720 9.9765 3.7980 11.0700 ;
      RECT 3.6640 9.9765 3.6900 11.0700 ;
      RECT 3.5560 9.9765 3.5820 11.0700 ;
      RECT 3.4480 9.9765 3.4740 11.0700 ;
      RECT 3.3400 9.9765 3.3660 11.0700 ;
      RECT 3.2320 9.9765 3.2580 11.0700 ;
      RECT 3.1240 9.9765 3.1500 11.0700 ;
      RECT 3.0160 9.9765 3.0420 11.0700 ;
      RECT 2.9080 9.9765 2.9340 11.0700 ;
      RECT 2.8000 9.9765 2.8260 11.0700 ;
      RECT 2.6920 9.9765 2.7180 11.0700 ;
      RECT 2.5840 9.9765 2.6100 11.0700 ;
      RECT 2.4760 9.9765 2.5020 11.0700 ;
      RECT 2.3680 9.9765 2.3940 11.0700 ;
      RECT 2.2600 9.9765 2.2860 11.0700 ;
      RECT 2.1520 9.9765 2.1780 11.0700 ;
      RECT 2.0440 9.9765 2.0700 11.0700 ;
      RECT 1.9360 9.9765 1.9620 11.0700 ;
      RECT 1.8280 9.9765 1.8540 11.0700 ;
      RECT 1.7200 9.9765 1.7460 11.0700 ;
      RECT 1.6120 9.9765 1.6380 11.0700 ;
      RECT 1.5040 9.9765 1.5300 11.0700 ;
      RECT 1.3960 9.9765 1.4220 11.0700 ;
      RECT 1.2880 9.9765 1.3140 11.0700 ;
      RECT 1.1800 9.9765 1.2060 11.0700 ;
      RECT 1.0720 9.9765 1.0980 11.0700 ;
      RECT 0.9640 9.9765 0.9900 11.0700 ;
      RECT 0.8560 9.9765 0.8820 11.0700 ;
      RECT 0.7480 9.9765 0.7740 11.0700 ;
      RECT 0.6400 9.9765 0.6660 11.0700 ;
      RECT 0.5320 9.9765 0.5580 11.0700 ;
      RECT 0.4240 9.9765 0.4500 11.0700 ;
      RECT 0.3160 9.9765 0.3420 11.0700 ;
      RECT 0.2080 9.9765 0.2340 11.0700 ;
      RECT 0.0050 9.9765 0.0900 11.0700 ;
      RECT 15.5530 11.0565 15.6810 12.1500 ;
      RECT 15.5390 11.7220 15.6810 12.0445 ;
      RECT 15.3190 11.4490 15.4530 12.1500 ;
      RECT 15.2960 11.7840 15.4530 12.0420 ;
      RECT 15.3190 11.0565 15.4170 12.1500 ;
      RECT 15.3190 11.1775 15.4310 11.4170 ;
      RECT 15.3190 11.0565 15.4530 11.1455 ;
      RECT 15.0940 11.5070 15.2280 12.1500 ;
      RECT 15.0940 11.0565 15.1920 12.1500 ;
      RECT 14.6770 11.0565 14.7600 12.1500 ;
      RECT 14.6770 11.1450 14.7740 12.0805 ;
      RECT 30.2680 11.0565 30.3530 12.1500 ;
      RECT 30.1240 11.0565 30.1500 12.1500 ;
      RECT 30.0160 11.0565 30.0420 12.1500 ;
      RECT 29.9080 11.0565 29.9340 12.1500 ;
      RECT 29.8000 11.0565 29.8260 12.1500 ;
      RECT 29.6920 11.0565 29.7180 12.1500 ;
      RECT 29.5840 11.0565 29.6100 12.1500 ;
      RECT 29.4760 11.0565 29.5020 12.1500 ;
      RECT 29.3680 11.0565 29.3940 12.1500 ;
      RECT 29.2600 11.0565 29.2860 12.1500 ;
      RECT 29.1520 11.0565 29.1780 12.1500 ;
      RECT 29.0440 11.0565 29.0700 12.1500 ;
      RECT 28.9360 11.0565 28.9620 12.1500 ;
      RECT 28.8280 11.0565 28.8540 12.1500 ;
      RECT 28.7200 11.0565 28.7460 12.1500 ;
      RECT 28.6120 11.0565 28.6380 12.1500 ;
      RECT 28.5040 11.0565 28.5300 12.1500 ;
      RECT 28.3960 11.0565 28.4220 12.1500 ;
      RECT 28.2880 11.0565 28.3140 12.1500 ;
      RECT 28.1800 11.0565 28.2060 12.1500 ;
      RECT 28.0720 11.0565 28.0980 12.1500 ;
      RECT 27.9640 11.0565 27.9900 12.1500 ;
      RECT 27.8560 11.0565 27.8820 12.1500 ;
      RECT 27.7480 11.0565 27.7740 12.1500 ;
      RECT 27.6400 11.0565 27.6660 12.1500 ;
      RECT 27.5320 11.0565 27.5580 12.1500 ;
      RECT 27.4240 11.0565 27.4500 12.1500 ;
      RECT 27.3160 11.0565 27.3420 12.1500 ;
      RECT 27.2080 11.0565 27.2340 12.1500 ;
      RECT 27.1000 11.0565 27.1260 12.1500 ;
      RECT 26.9920 11.0565 27.0180 12.1500 ;
      RECT 26.8840 11.0565 26.9100 12.1500 ;
      RECT 26.7760 11.0565 26.8020 12.1500 ;
      RECT 26.6680 11.0565 26.6940 12.1500 ;
      RECT 26.5600 11.0565 26.5860 12.1500 ;
      RECT 26.4520 11.0565 26.4780 12.1500 ;
      RECT 26.3440 11.0565 26.3700 12.1500 ;
      RECT 26.2360 11.0565 26.2620 12.1500 ;
      RECT 26.1280 11.0565 26.1540 12.1500 ;
      RECT 26.0200 11.0565 26.0460 12.1500 ;
      RECT 25.9120 11.0565 25.9380 12.1500 ;
      RECT 25.8040 11.0565 25.8300 12.1500 ;
      RECT 25.6960 11.0565 25.7220 12.1500 ;
      RECT 25.5880 11.0565 25.6140 12.1500 ;
      RECT 25.4800 11.0565 25.5060 12.1500 ;
      RECT 25.3720 11.0565 25.3980 12.1500 ;
      RECT 25.2640 11.0565 25.2900 12.1500 ;
      RECT 25.1560 11.0565 25.1820 12.1500 ;
      RECT 25.0480 11.0565 25.0740 12.1500 ;
      RECT 24.9400 11.0565 24.9660 12.1500 ;
      RECT 24.8320 11.0565 24.8580 12.1500 ;
      RECT 24.7240 11.0565 24.7500 12.1500 ;
      RECT 24.6160 11.0565 24.6420 12.1500 ;
      RECT 24.5080 11.0565 24.5340 12.1500 ;
      RECT 24.4000 11.0565 24.4260 12.1500 ;
      RECT 24.2920 11.0565 24.3180 12.1500 ;
      RECT 24.1840 11.0565 24.2100 12.1500 ;
      RECT 24.0760 11.0565 24.1020 12.1500 ;
      RECT 23.9680 11.0565 23.9940 12.1500 ;
      RECT 23.8600 11.0565 23.8860 12.1500 ;
      RECT 23.7520 11.0565 23.7780 12.1500 ;
      RECT 23.6440 11.0565 23.6700 12.1500 ;
      RECT 23.5360 11.0565 23.5620 12.1500 ;
      RECT 23.4280 11.0565 23.4540 12.1500 ;
      RECT 23.3200 11.0565 23.3460 12.1500 ;
      RECT 23.2120 11.0565 23.2380 12.1500 ;
      RECT 23.1040 11.0565 23.1300 12.1500 ;
      RECT 22.9960 11.0565 23.0220 12.1500 ;
      RECT 22.8880 11.0565 22.9140 12.1500 ;
      RECT 22.7800 11.0565 22.8060 12.1500 ;
      RECT 22.6720 11.0565 22.6980 12.1500 ;
      RECT 22.5640 11.0565 22.5900 12.1500 ;
      RECT 22.4560 11.0565 22.4820 12.1500 ;
      RECT 22.3480 11.0565 22.3740 12.1500 ;
      RECT 22.2400 11.0565 22.2660 12.1500 ;
      RECT 22.1320 11.0565 22.1580 12.1500 ;
      RECT 22.0240 11.0565 22.0500 12.1500 ;
      RECT 21.9160 11.0565 21.9420 12.1500 ;
      RECT 21.8080 11.0565 21.8340 12.1500 ;
      RECT 21.7000 11.0565 21.7260 12.1500 ;
      RECT 21.5920 11.0565 21.6180 12.1500 ;
      RECT 21.4840 11.0565 21.5100 12.1500 ;
      RECT 21.3760 11.0565 21.4020 12.1500 ;
      RECT 21.2680 11.0565 21.2940 12.1500 ;
      RECT 21.1600 11.0565 21.1860 12.1500 ;
      RECT 21.0520 11.0565 21.0780 12.1500 ;
      RECT 20.9440 11.0565 20.9700 12.1500 ;
      RECT 20.8360 11.0565 20.8620 12.1500 ;
      RECT 20.7280 11.0565 20.7540 12.1500 ;
      RECT 20.6200 11.0565 20.6460 12.1500 ;
      RECT 20.5120 11.0565 20.5380 12.1500 ;
      RECT 20.4040 11.0565 20.4300 12.1500 ;
      RECT 20.2960 11.0565 20.3220 12.1500 ;
      RECT 20.1880 11.0565 20.2140 12.1500 ;
      RECT 20.0800 11.0565 20.1060 12.1500 ;
      RECT 19.9720 11.0565 19.9980 12.1500 ;
      RECT 19.8640 11.0565 19.8900 12.1500 ;
      RECT 19.7560 11.0565 19.7820 12.1500 ;
      RECT 19.6480 11.0565 19.6740 12.1500 ;
      RECT 19.5400 11.0565 19.5660 12.1500 ;
      RECT 19.4320 11.0565 19.4580 12.1500 ;
      RECT 19.3240 11.0565 19.3500 12.1500 ;
      RECT 19.2160 11.0565 19.2420 12.1500 ;
      RECT 19.1080 11.0565 19.1340 12.1500 ;
      RECT 19.0000 11.0565 19.0260 12.1500 ;
      RECT 18.8920 11.0565 18.9180 12.1500 ;
      RECT 18.7840 11.0565 18.8100 12.1500 ;
      RECT 18.6760 11.0565 18.7020 12.1500 ;
      RECT 18.5680 11.0565 18.5940 12.1500 ;
      RECT 18.4600 11.0565 18.4860 12.1500 ;
      RECT 18.3520 11.0565 18.3780 12.1500 ;
      RECT 18.2440 11.0565 18.2700 12.1500 ;
      RECT 18.1360 11.0565 18.1620 12.1500 ;
      RECT 18.0280 11.0565 18.0540 12.1500 ;
      RECT 17.9200 11.0565 17.9460 12.1500 ;
      RECT 17.8120 11.0565 17.8380 12.1500 ;
      RECT 17.7040 11.0565 17.7300 12.1500 ;
      RECT 17.5960 11.0565 17.6220 12.1500 ;
      RECT 17.4880 11.0565 17.5140 12.1500 ;
      RECT 17.3800 11.0565 17.4060 12.1500 ;
      RECT 17.2720 11.0565 17.2980 12.1500 ;
      RECT 17.1640 11.0565 17.1900 12.1500 ;
      RECT 17.0560 11.0565 17.0820 12.1500 ;
      RECT 16.9480 11.0565 16.9740 12.1500 ;
      RECT 16.8400 11.0565 16.8660 12.1500 ;
      RECT 16.7320 11.0565 16.7580 12.1500 ;
      RECT 16.6240 11.0565 16.6500 12.1500 ;
      RECT 16.5160 11.0565 16.5420 12.1500 ;
      RECT 16.4080 11.0565 16.4340 12.1500 ;
      RECT 16.3000 11.0565 16.3260 12.1500 ;
      RECT 16.0870 11.0565 16.1640 12.1500 ;
      RECT 14.1940 11.0565 14.2710 12.1500 ;
      RECT 14.0320 11.0565 14.0580 12.1500 ;
      RECT 13.9240 11.0565 13.9500 12.1500 ;
      RECT 13.8160 11.0565 13.8420 12.1500 ;
      RECT 13.7080 11.0565 13.7340 12.1500 ;
      RECT 13.6000 11.0565 13.6260 12.1500 ;
      RECT 13.4920 11.0565 13.5180 12.1500 ;
      RECT 13.3840 11.0565 13.4100 12.1500 ;
      RECT 13.2760 11.0565 13.3020 12.1500 ;
      RECT 13.1680 11.0565 13.1940 12.1500 ;
      RECT 13.0600 11.0565 13.0860 12.1500 ;
      RECT 12.9520 11.0565 12.9780 12.1500 ;
      RECT 12.8440 11.0565 12.8700 12.1500 ;
      RECT 12.7360 11.0565 12.7620 12.1500 ;
      RECT 12.6280 11.0565 12.6540 12.1500 ;
      RECT 12.5200 11.0565 12.5460 12.1500 ;
      RECT 12.4120 11.0565 12.4380 12.1500 ;
      RECT 12.3040 11.0565 12.3300 12.1500 ;
      RECT 12.1960 11.0565 12.2220 12.1500 ;
      RECT 12.0880 11.0565 12.1140 12.1500 ;
      RECT 11.9800 11.0565 12.0060 12.1500 ;
      RECT 11.8720 11.0565 11.8980 12.1500 ;
      RECT 11.7640 11.0565 11.7900 12.1500 ;
      RECT 11.6560 11.0565 11.6820 12.1500 ;
      RECT 11.5480 11.0565 11.5740 12.1500 ;
      RECT 11.4400 11.0565 11.4660 12.1500 ;
      RECT 11.3320 11.0565 11.3580 12.1500 ;
      RECT 11.2240 11.0565 11.2500 12.1500 ;
      RECT 11.1160 11.0565 11.1420 12.1500 ;
      RECT 11.0080 11.0565 11.0340 12.1500 ;
      RECT 10.9000 11.0565 10.9260 12.1500 ;
      RECT 10.7920 11.0565 10.8180 12.1500 ;
      RECT 10.6840 11.0565 10.7100 12.1500 ;
      RECT 10.5760 11.0565 10.6020 12.1500 ;
      RECT 10.4680 11.0565 10.4940 12.1500 ;
      RECT 10.3600 11.0565 10.3860 12.1500 ;
      RECT 10.2520 11.0565 10.2780 12.1500 ;
      RECT 10.1440 11.0565 10.1700 12.1500 ;
      RECT 10.0360 11.0565 10.0620 12.1500 ;
      RECT 9.9280 11.0565 9.9540 12.1500 ;
      RECT 9.8200 11.0565 9.8460 12.1500 ;
      RECT 9.7120 11.0565 9.7380 12.1500 ;
      RECT 9.6040 11.0565 9.6300 12.1500 ;
      RECT 9.4960 11.0565 9.5220 12.1500 ;
      RECT 9.3880 11.0565 9.4140 12.1500 ;
      RECT 9.2800 11.0565 9.3060 12.1500 ;
      RECT 9.1720 11.0565 9.1980 12.1500 ;
      RECT 9.0640 11.0565 9.0900 12.1500 ;
      RECT 8.9560 11.0565 8.9820 12.1500 ;
      RECT 8.8480 11.0565 8.8740 12.1500 ;
      RECT 8.7400 11.0565 8.7660 12.1500 ;
      RECT 8.6320 11.0565 8.6580 12.1500 ;
      RECT 8.5240 11.0565 8.5500 12.1500 ;
      RECT 8.4160 11.0565 8.4420 12.1500 ;
      RECT 8.3080 11.0565 8.3340 12.1500 ;
      RECT 8.2000 11.0565 8.2260 12.1500 ;
      RECT 8.0920 11.0565 8.1180 12.1500 ;
      RECT 7.9840 11.0565 8.0100 12.1500 ;
      RECT 7.8760 11.0565 7.9020 12.1500 ;
      RECT 7.7680 11.0565 7.7940 12.1500 ;
      RECT 7.6600 11.0565 7.6860 12.1500 ;
      RECT 7.5520 11.0565 7.5780 12.1500 ;
      RECT 7.4440 11.0565 7.4700 12.1500 ;
      RECT 7.3360 11.0565 7.3620 12.1500 ;
      RECT 7.2280 11.0565 7.2540 12.1500 ;
      RECT 7.1200 11.0565 7.1460 12.1500 ;
      RECT 7.0120 11.0565 7.0380 12.1500 ;
      RECT 6.9040 11.0565 6.9300 12.1500 ;
      RECT 6.7960 11.0565 6.8220 12.1500 ;
      RECT 6.6880 11.0565 6.7140 12.1500 ;
      RECT 6.5800 11.0565 6.6060 12.1500 ;
      RECT 6.4720 11.0565 6.4980 12.1500 ;
      RECT 6.3640 11.0565 6.3900 12.1500 ;
      RECT 6.2560 11.0565 6.2820 12.1500 ;
      RECT 6.1480 11.0565 6.1740 12.1500 ;
      RECT 6.0400 11.0565 6.0660 12.1500 ;
      RECT 5.9320 11.0565 5.9580 12.1500 ;
      RECT 5.8240 11.0565 5.8500 12.1500 ;
      RECT 5.7160 11.0565 5.7420 12.1500 ;
      RECT 5.6080 11.0565 5.6340 12.1500 ;
      RECT 5.5000 11.0565 5.5260 12.1500 ;
      RECT 5.3920 11.0565 5.4180 12.1500 ;
      RECT 5.2840 11.0565 5.3100 12.1500 ;
      RECT 5.1760 11.0565 5.2020 12.1500 ;
      RECT 5.0680 11.0565 5.0940 12.1500 ;
      RECT 4.9600 11.0565 4.9860 12.1500 ;
      RECT 4.8520 11.0565 4.8780 12.1500 ;
      RECT 4.7440 11.0565 4.7700 12.1500 ;
      RECT 4.6360 11.0565 4.6620 12.1500 ;
      RECT 4.5280 11.0565 4.5540 12.1500 ;
      RECT 4.4200 11.0565 4.4460 12.1500 ;
      RECT 4.3120 11.0565 4.3380 12.1500 ;
      RECT 4.2040 11.0565 4.2300 12.1500 ;
      RECT 4.0960 11.0565 4.1220 12.1500 ;
      RECT 3.9880 11.0565 4.0140 12.1500 ;
      RECT 3.8800 11.0565 3.9060 12.1500 ;
      RECT 3.7720 11.0565 3.7980 12.1500 ;
      RECT 3.6640 11.0565 3.6900 12.1500 ;
      RECT 3.5560 11.0565 3.5820 12.1500 ;
      RECT 3.4480 11.0565 3.4740 12.1500 ;
      RECT 3.3400 11.0565 3.3660 12.1500 ;
      RECT 3.2320 11.0565 3.2580 12.1500 ;
      RECT 3.1240 11.0565 3.1500 12.1500 ;
      RECT 3.0160 11.0565 3.0420 12.1500 ;
      RECT 2.9080 11.0565 2.9340 12.1500 ;
      RECT 2.8000 11.0565 2.8260 12.1500 ;
      RECT 2.6920 11.0565 2.7180 12.1500 ;
      RECT 2.5840 11.0565 2.6100 12.1500 ;
      RECT 2.4760 11.0565 2.5020 12.1500 ;
      RECT 2.3680 11.0565 2.3940 12.1500 ;
      RECT 2.2600 11.0565 2.2860 12.1500 ;
      RECT 2.1520 11.0565 2.1780 12.1500 ;
      RECT 2.0440 11.0565 2.0700 12.1500 ;
      RECT 1.9360 11.0565 1.9620 12.1500 ;
      RECT 1.8280 11.0565 1.8540 12.1500 ;
      RECT 1.7200 11.0565 1.7460 12.1500 ;
      RECT 1.6120 11.0565 1.6380 12.1500 ;
      RECT 1.5040 11.0565 1.5300 12.1500 ;
      RECT 1.3960 11.0565 1.4220 12.1500 ;
      RECT 1.2880 11.0565 1.3140 12.1500 ;
      RECT 1.1800 11.0565 1.2060 12.1500 ;
      RECT 1.0720 11.0565 1.0980 12.1500 ;
      RECT 0.9640 11.0565 0.9900 12.1500 ;
      RECT 0.8560 11.0565 0.8820 12.1500 ;
      RECT 0.7480 11.0565 0.7740 12.1500 ;
      RECT 0.6400 11.0565 0.6660 12.1500 ;
      RECT 0.5320 11.0565 0.5580 12.1500 ;
      RECT 0.4240 11.0565 0.4500 12.1500 ;
      RECT 0.3160 11.0565 0.3420 12.1500 ;
      RECT 0.2080 11.0565 0.2340 12.1500 ;
      RECT 0.0050 11.0565 0.0900 12.1500 ;
      RECT 15.5530 12.1365 15.6810 13.2300 ;
      RECT 15.5390 12.8020 15.6810 13.1245 ;
      RECT 15.3190 12.5290 15.4530 13.2300 ;
      RECT 15.2960 12.8640 15.4530 13.1220 ;
      RECT 15.3190 12.1365 15.4170 13.2300 ;
      RECT 15.3190 12.2575 15.4310 12.4970 ;
      RECT 15.3190 12.1365 15.4530 12.2255 ;
      RECT 15.0940 12.5870 15.2280 13.2300 ;
      RECT 15.0940 12.1365 15.1920 13.2300 ;
      RECT 14.6770 12.1365 14.7600 13.2300 ;
      RECT 14.6770 12.2250 14.7740 13.1605 ;
      RECT 30.2680 12.1365 30.3530 13.2300 ;
      RECT 30.1240 12.1365 30.1500 13.2300 ;
      RECT 30.0160 12.1365 30.0420 13.2300 ;
      RECT 29.9080 12.1365 29.9340 13.2300 ;
      RECT 29.8000 12.1365 29.8260 13.2300 ;
      RECT 29.6920 12.1365 29.7180 13.2300 ;
      RECT 29.5840 12.1365 29.6100 13.2300 ;
      RECT 29.4760 12.1365 29.5020 13.2300 ;
      RECT 29.3680 12.1365 29.3940 13.2300 ;
      RECT 29.2600 12.1365 29.2860 13.2300 ;
      RECT 29.1520 12.1365 29.1780 13.2300 ;
      RECT 29.0440 12.1365 29.0700 13.2300 ;
      RECT 28.9360 12.1365 28.9620 13.2300 ;
      RECT 28.8280 12.1365 28.8540 13.2300 ;
      RECT 28.7200 12.1365 28.7460 13.2300 ;
      RECT 28.6120 12.1365 28.6380 13.2300 ;
      RECT 28.5040 12.1365 28.5300 13.2300 ;
      RECT 28.3960 12.1365 28.4220 13.2300 ;
      RECT 28.2880 12.1365 28.3140 13.2300 ;
      RECT 28.1800 12.1365 28.2060 13.2300 ;
      RECT 28.0720 12.1365 28.0980 13.2300 ;
      RECT 27.9640 12.1365 27.9900 13.2300 ;
      RECT 27.8560 12.1365 27.8820 13.2300 ;
      RECT 27.7480 12.1365 27.7740 13.2300 ;
      RECT 27.6400 12.1365 27.6660 13.2300 ;
      RECT 27.5320 12.1365 27.5580 13.2300 ;
      RECT 27.4240 12.1365 27.4500 13.2300 ;
      RECT 27.3160 12.1365 27.3420 13.2300 ;
      RECT 27.2080 12.1365 27.2340 13.2300 ;
      RECT 27.1000 12.1365 27.1260 13.2300 ;
      RECT 26.9920 12.1365 27.0180 13.2300 ;
      RECT 26.8840 12.1365 26.9100 13.2300 ;
      RECT 26.7760 12.1365 26.8020 13.2300 ;
      RECT 26.6680 12.1365 26.6940 13.2300 ;
      RECT 26.5600 12.1365 26.5860 13.2300 ;
      RECT 26.4520 12.1365 26.4780 13.2300 ;
      RECT 26.3440 12.1365 26.3700 13.2300 ;
      RECT 26.2360 12.1365 26.2620 13.2300 ;
      RECT 26.1280 12.1365 26.1540 13.2300 ;
      RECT 26.0200 12.1365 26.0460 13.2300 ;
      RECT 25.9120 12.1365 25.9380 13.2300 ;
      RECT 25.8040 12.1365 25.8300 13.2300 ;
      RECT 25.6960 12.1365 25.7220 13.2300 ;
      RECT 25.5880 12.1365 25.6140 13.2300 ;
      RECT 25.4800 12.1365 25.5060 13.2300 ;
      RECT 25.3720 12.1365 25.3980 13.2300 ;
      RECT 25.2640 12.1365 25.2900 13.2300 ;
      RECT 25.1560 12.1365 25.1820 13.2300 ;
      RECT 25.0480 12.1365 25.0740 13.2300 ;
      RECT 24.9400 12.1365 24.9660 13.2300 ;
      RECT 24.8320 12.1365 24.8580 13.2300 ;
      RECT 24.7240 12.1365 24.7500 13.2300 ;
      RECT 24.6160 12.1365 24.6420 13.2300 ;
      RECT 24.5080 12.1365 24.5340 13.2300 ;
      RECT 24.4000 12.1365 24.4260 13.2300 ;
      RECT 24.2920 12.1365 24.3180 13.2300 ;
      RECT 24.1840 12.1365 24.2100 13.2300 ;
      RECT 24.0760 12.1365 24.1020 13.2300 ;
      RECT 23.9680 12.1365 23.9940 13.2300 ;
      RECT 23.8600 12.1365 23.8860 13.2300 ;
      RECT 23.7520 12.1365 23.7780 13.2300 ;
      RECT 23.6440 12.1365 23.6700 13.2300 ;
      RECT 23.5360 12.1365 23.5620 13.2300 ;
      RECT 23.4280 12.1365 23.4540 13.2300 ;
      RECT 23.3200 12.1365 23.3460 13.2300 ;
      RECT 23.2120 12.1365 23.2380 13.2300 ;
      RECT 23.1040 12.1365 23.1300 13.2300 ;
      RECT 22.9960 12.1365 23.0220 13.2300 ;
      RECT 22.8880 12.1365 22.9140 13.2300 ;
      RECT 22.7800 12.1365 22.8060 13.2300 ;
      RECT 22.6720 12.1365 22.6980 13.2300 ;
      RECT 22.5640 12.1365 22.5900 13.2300 ;
      RECT 22.4560 12.1365 22.4820 13.2300 ;
      RECT 22.3480 12.1365 22.3740 13.2300 ;
      RECT 22.2400 12.1365 22.2660 13.2300 ;
      RECT 22.1320 12.1365 22.1580 13.2300 ;
      RECT 22.0240 12.1365 22.0500 13.2300 ;
      RECT 21.9160 12.1365 21.9420 13.2300 ;
      RECT 21.8080 12.1365 21.8340 13.2300 ;
      RECT 21.7000 12.1365 21.7260 13.2300 ;
      RECT 21.5920 12.1365 21.6180 13.2300 ;
      RECT 21.4840 12.1365 21.5100 13.2300 ;
      RECT 21.3760 12.1365 21.4020 13.2300 ;
      RECT 21.2680 12.1365 21.2940 13.2300 ;
      RECT 21.1600 12.1365 21.1860 13.2300 ;
      RECT 21.0520 12.1365 21.0780 13.2300 ;
      RECT 20.9440 12.1365 20.9700 13.2300 ;
      RECT 20.8360 12.1365 20.8620 13.2300 ;
      RECT 20.7280 12.1365 20.7540 13.2300 ;
      RECT 20.6200 12.1365 20.6460 13.2300 ;
      RECT 20.5120 12.1365 20.5380 13.2300 ;
      RECT 20.4040 12.1365 20.4300 13.2300 ;
      RECT 20.2960 12.1365 20.3220 13.2300 ;
      RECT 20.1880 12.1365 20.2140 13.2300 ;
      RECT 20.0800 12.1365 20.1060 13.2300 ;
      RECT 19.9720 12.1365 19.9980 13.2300 ;
      RECT 19.8640 12.1365 19.8900 13.2300 ;
      RECT 19.7560 12.1365 19.7820 13.2300 ;
      RECT 19.6480 12.1365 19.6740 13.2300 ;
      RECT 19.5400 12.1365 19.5660 13.2300 ;
      RECT 19.4320 12.1365 19.4580 13.2300 ;
      RECT 19.3240 12.1365 19.3500 13.2300 ;
      RECT 19.2160 12.1365 19.2420 13.2300 ;
      RECT 19.1080 12.1365 19.1340 13.2300 ;
      RECT 19.0000 12.1365 19.0260 13.2300 ;
      RECT 18.8920 12.1365 18.9180 13.2300 ;
      RECT 18.7840 12.1365 18.8100 13.2300 ;
      RECT 18.6760 12.1365 18.7020 13.2300 ;
      RECT 18.5680 12.1365 18.5940 13.2300 ;
      RECT 18.4600 12.1365 18.4860 13.2300 ;
      RECT 18.3520 12.1365 18.3780 13.2300 ;
      RECT 18.2440 12.1365 18.2700 13.2300 ;
      RECT 18.1360 12.1365 18.1620 13.2300 ;
      RECT 18.0280 12.1365 18.0540 13.2300 ;
      RECT 17.9200 12.1365 17.9460 13.2300 ;
      RECT 17.8120 12.1365 17.8380 13.2300 ;
      RECT 17.7040 12.1365 17.7300 13.2300 ;
      RECT 17.5960 12.1365 17.6220 13.2300 ;
      RECT 17.4880 12.1365 17.5140 13.2300 ;
      RECT 17.3800 12.1365 17.4060 13.2300 ;
      RECT 17.2720 12.1365 17.2980 13.2300 ;
      RECT 17.1640 12.1365 17.1900 13.2300 ;
      RECT 17.0560 12.1365 17.0820 13.2300 ;
      RECT 16.9480 12.1365 16.9740 13.2300 ;
      RECT 16.8400 12.1365 16.8660 13.2300 ;
      RECT 16.7320 12.1365 16.7580 13.2300 ;
      RECT 16.6240 12.1365 16.6500 13.2300 ;
      RECT 16.5160 12.1365 16.5420 13.2300 ;
      RECT 16.4080 12.1365 16.4340 13.2300 ;
      RECT 16.3000 12.1365 16.3260 13.2300 ;
      RECT 16.0870 12.1365 16.1640 13.2300 ;
      RECT 14.1940 12.1365 14.2710 13.2300 ;
      RECT 14.0320 12.1365 14.0580 13.2300 ;
      RECT 13.9240 12.1365 13.9500 13.2300 ;
      RECT 13.8160 12.1365 13.8420 13.2300 ;
      RECT 13.7080 12.1365 13.7340 13.2300 ;
      RECT 13.6000 12.1365 13.6260 13.2300 ;
      RECT 13.4920 12.1365 13.5180 13.2300 ;
      RECT 13.3840 12.1365 13.4100 13.2300 ;
      RECT 13.2760 12.1365 13.3020 13.2300 ;
      RECT 13.1680 12.1365 13.1940 13.2300 ;
      RECT 13.0600 12.1365 13.0860 13.2300 ;
      RECT 12.9520 12.1365 12.9780 13.2300 ;
      RECT 12.8440 12.1365 12.8700 13.2300 ;
      RECT 12.7360 12.1365 12.7620 13.2300 ;
      RECT 12.6280 12.1365 12.6540 13.2300 ;
      RECT 12.5200 12.1365 12.5460 13.2300 ;
      RECT 12.4120 12.1365 12.4380 13.2300 ;
      RECT 12.3040 12.1365 12.3300 13.2300 ;
      RECT 12.1960 12.1365 12.2220 13.2300 ;
      RECT 12.0880 12.1365 12.1140 13.2300 ;
      RECT 11.9800 12.1365 12.0060 13.2300 ;
      RECT 11.8720 12.1365 11.8980 13.2300 ;
      RECT 11.7640 12.1365 11.7900 13.2300 ;
      RECT 11.6560 12.1365 11.6820 13.2300 ;
      RECT 11.5480 12.1365 11.5740 13.2300 ;
      RECT 11.4400 12.1365 11.4660 13.2300 ;
      RECT 11.3320 12.1365 11.3580 13.2300 ;
      RECT 11.2240 12.1365 11.2500 13.2300 ;
      RECT 11.1160 12.1365 11.1420 13.2300 ;
      RECT 11.0080 12.1365 11.0340 13.2300 ;
      RECT 10.9000 12.1365 10.9260 13.2300 ;
      RECT 10.7920 12.1365 10.8180 13.2300 ;
      RECT 10.6840 12.1365 10.7100 13.2300 ;
      RECT 10.5760 12.1365 10.6020 13.2300 ;
      RECT 10.4680 12.1365 10.4940 13.2300 ;
      RECT 10.3600 12.1365 10.3860 13.2300 ;
      RECT 10.2520 12.1365 10.2780 13.2300 ;
      RECT 10.1440 12.1365 10.1700 13.2300 ;
      RECT 10.0360 12.1365 10.0620 13.2300 ;
      RECT 9.9280 12.1365 9.9540 13.2300 ;
      RECT 9.8200 12.1365 9.8460 13.2300 ;
      RECT 9.7120 12.1365 9.7380 13.2300 ;
      RECT 9.6040 12.1365 9.6300 13.2300 ;
      RECT 9.4960 12.1365 9.5220 13.2300 ;
      RECT 9.3880 12.1365 9.4140 13.2300 ;
      RECT 9.2800 12.1365 9.3060 13.2300 ;
      RECT 9.1720 12.1365 9.1980 13.2300 ;
      RECT 9.0640 12.1365 9.0900 13.2300 ;
      RECT 8.9560 12.1365 8.9820 13.2300 ;
      RECT 8.8480 12.1365 8.8740 13.2300 ;
      RECT 8.7400 12.1365 8.7660 13.2300 ;
      RECT 8.6320 12.1365 8.6580 13.2300 ;
      RECT 8.5240 12.1365 8.5500 13.2300 ;
      RECT 8.4160 12.1365 8.4420 13.2300 ;
      RECT 8.3080 12.1365 8.3340 13.2300 ;
      RECT 8.2000 12.1365 8.2260 13.2300 ;
      RECT 8.0920 12.1365 8.1180 13.2300 ;
      RECT 7.9840 12.1365 8.0100 13.2300 ;
      RECT 7.8760 12.1365 7.9020 13.2300 ;
      RECT 7.7680 12.1365 7.7940 13.2300 ;
      RECT 7.6600 12.1365 7.6860 13.2300 ;
      RECT 7.5520 12.1365 7.5780 13.2300 ;
      RECT 7.4440 12.1365 7.4700 13.2300 ;
      RECT 7.3360 12.1365 7.3620 13.2300 ;
      RECT 7.2280 12.1365 7.2540 13.2300 ;
      RECT 7.1200 12.1365 7.1460 13.2300 ;
      RECT 7.0120 12.1365 7.0380 13.2300 ;
      RECT 6.9040 12.1365 6.9300 13.2300 ;
      RECT 6.7960 12.1365 6.8220 13.2300 ;
      RECT 6.6880 12.1365 6.7140 13.2300 ;
      RECT 6.5800 12.1365 6.6060 13.2300 ;
      RECT 6.4720 12.1365 6.4980 13.2300 ;
      RECT 6.3640 12.1365 6.3900 13.2300 ;
      RECT 6.2560 12.1365 6.2820 13.2300 ;
      RECT 6.1480 12.1365 6.1740 13.2300 ;
      RECT 6.0400 12.1365 6.0660 13.2300 ;
      RECT 5.9320 12.1365 5.9580 13.2300 ;
      RECT 5.8240 12.1365 5.8500 13.2300 ;
      RECT 5.7160 12.1365 5.7420 13.2300 ;
      RECT 5.6080 12.1365 5.6340 13.2300 ;
      RECT 5.5000 12.1365 5.5260 13.2300 ;
      RECT 5.3920 12.1365 5.4180 13.2300 ;
      RECT 5.2840 12.1365 5.3100 13.2300 ;
      RECT 5.1760 12.1365 5.2020 13.2300 ;
      RECT 5.0680 12.1365 5.0940 13.2300 ;
      RECT 4.9600 12.1365 4.9860 13.2300 ;
      RECT 4.8520 12.1365 4.8780 13.2300 ;
      RECT 4.7440 12.1365 4.7700 13.2300 ;
      RECT 4.6360 12.1365 4.6620 13.2300 ;
      RECT 4.5280 12.1365 4.5540 13.2300 ;
      RECT 4.4200 12.1365 4.4460 13.2300 ;
      RECT 4.3120 12.1365 4.3380 13.2300 ;
      RECT 4.2040 12.1365 4.2300 13.2300 ;
      RECT 4.0960 12.1365 4.1220 13.2300 ;
      RECT 3.9880 12.1365 4.0140 13.2300 ;
      RECT 3.8800 12.1365 3.9060 13.2300 ;
      RECT 3.7720 12.1365 3.7980 13.2300 ;
      RECT 3.6640 12.1365 3.6900 13.2300 ;
      RECT 3.5560 12.1365 3.5820 13.2300 ;
      RECT 3.4480 12.1365 3.4740 13.2300 ;
      RECT 3.3400 12.1365 3.3660 13.2300 ;
      RECT 3.2320 12.1365 3.2580 13.2300 ;
      RECT 3.1240 12.1365 3.1500 13.2300 ;
      RECT 3.0160 12.1365 3.0420 13.2300 ;
      RECT 2.9080 12.1365 2.9340 13.2300 ;
      RECT 2.8000 12.1365 2.8260 13.2300 ;
      RECT 2.6920 12.1365 2.7180 13.2300 ;
      RECT 2.5840 12.1365 2.6100 13.2300 ;
      RECT 2.4760 12.1365 2.5020 13.2300 ;
      RECT 2.3680 12.1365 2.3940 13.2300 ;
      RECT 2.2600 12.1365 2.2860 13.2300 ;
      RECT 2.1520 12.1365 2.1780 13.2300 ;
      RECT 2.0440 12.1365 2.0700 13.2300 ;
      RECT 1.9360 12.1365 1.9620 13.2300 ;
      RECT 1.8280 12.1365 1.8540 13.2300 ;
      RECT 1.7200 12.1365 1.7460 13.2300 ;
      RECT 1.6120 12.1365 1.6380 13.2300 ;
      RECT 1.5040 12.1365 1.5300 13.2300 ;
      RECT 1.3960 12.1365 1.4220 13.2300 ;
      RECT 1.2880 12.1365 1.3140 13.2300 ;
      RECT 1.1800 12.1365 1.2060 13.2300 ;
      RECT 1.0720 12.1365 1.0980 13.2300 ;
      RECT 0.9640 12.1365 0.9900 13.2300 ;
      RECT 0.8560 12.1365 0.8820 13.2300 ;
      RECT 0.7480 12.1365 0.7740 13.2300 ;
      RECT 0.6400 12.1365 0.6660 13.2300 ;
      RECT 0.5320 12.1365 0.5580 13.2300 ;
      RECT 0.4240 12.1365 0.4500 13.2300 ;
      RECT 0.3160 12.1365 0.3420 13.2300 ;
      RECT 0.2080 12.1365 0.2340 13.2300 ;
      RECT 0.0050 12.1365 0.0900 13.2300 ;
      RECT 15.5530 13.2165 15.6810 14.3100 ;
      RECT 15.5390 13.8820 15.6810 14.2045 ;
      RECT 15.3190 13.6090 15.4530 14.3100 ;
      RECT 15.2960 13.9440 15.4530 14.2020 ;
      RECT 15.3190 13.2165 15.4170 14.3100 ;
      RECT 15.3190 13.3375 15.4310 13.5770 ;
      RECT 15.3190 13.2165 15.4530 13.3055 ;
      RECT 15.0940 13.6670 15.2280 14.3100 ;
      RECT 15.0940 13.2165 15.1920 14.3100 ;
      RECT 14.6770 13.2165 14.7600 14.3100 ;
      RECT 14.6770 13.3050 14.7740 14.2405 ;
      RECT 30.2680 13.2165 30.3530 14.3100 ;
      RECT 30.1240 13.2165 30.1500 14.3100 ;
      RECT 30.0160 13.2165 30.0420 14.3100 ;
      RECT 29.9080 13.2165 29.9340 14.3100 ;
      RECT 29.8000 13.2165 29.8260 14.3100 ;
      RECT 29.6920 13.2165 29.7180 14.3100 ;
      RECT 29.5840 13.2165 29.6100 14.3100 ;
      RECT 29.4760 13.2165 29.5020 14.3100 ;
      RECT 29.3680 13.2165 29.3940 14.3100 ;
      RECT 29.2600 13.2165 29.2860 14.3100 ;
      RECT 29.1520 13.2165 29.1780 14.3100 ;
      RECT 29.0440 13.2165 29.0700 14.3100 ;
      RECT 28.9360 13.2165 28.9620 14.3100 ;
      RECT 28.8280 13.2165 28.8540 14.3100 ;
      RECT 28.7200 13.2165 28.7460 14.3100 ;
      RECT 28.6120 13.2165 28.6380 14.3100 ;
      RECT 28.5040 13.2165 28.5300 14.3100 ;
      RECT 28.3960 13.2165 28.4220 14.3100 ;
      RECT 28.2880 13.2165 28.3140 14.3100 ;
      RECT 28.1800 13.2165 28.2060 14.3100 ;
      RECT 28.0720 13.2165 28.0980 14.3100 ;
      RECT 27.9640 13.2165 27.9900 14.3100 ;
      RECT 27.8560 13.2165 27.8820 14.3100 ;
      RECT 27.7480 13.2165 27.7740 14.3100 ;
      RECT 27.6400 13.2165 27.6660 14.3100 ;
      RECT 27.5320 13.2165 27.5580 14.3100 ;
      RECT 27.4240 13.2165 27.4500 14.3100 ;
      RECT 27.3160 13.2165 27.3420 14.3100 ;
      RECT 27.2080 13.2165 27.2340 14.3100 ;
      RECT 27.1000 13.2165 27.1260 14.3100 ;
      RECT 26.9920 13.2165 27.0180 14.3100 ;
      RECT 26.8840 13.2165 26.9100 14.3100 ;
      RECT 26.7760 13.2165 26.8020 14.3100 ;
      RECT 26.6680 13.2165 26.6940 14.3100 ;
      RECT 26.5600 13.2165 26.5860 14.3100 ;
      RECT 26.4520 13.2165 26.4780 14.3100 ;
      RECT 26.3440 13.2165 26.3700 14.3100 ;
      RECT 26.2360 13.2165 26.2620 14.3100 ;
      RECT 26.1280 13.2165 26.1540 14.3100 ;
      RECT 26.0200 13.2165 26.0460 14.3100 ;
      RECT 25.9120 13.2165 25.9380 14.3100 ;
      RECT 25.8040 13.2165 25.8300 14.3100 ;
      RECT 25.6960 13.2165 25.7220 14.3100 ;
      RECT 25.5880 13.2165 25.6140 14.3100 ;
      RECT 25.4800 13.2165 25.5060 14.3100 ;
      RECT 25.3720 13.2165 25.3980 14.3100 ;
      RECT 25.2640 13.2165 25.2900 14.3100 ;
      RECT 25.1560 13.2165 25.1820 14.3100 ;
      RECT 25.0480 13.2165 25.0740 14.3100 ;
      RECT 24.9400 13.2165 24.9660 14.3100 ;
      RECT 24.8320 13.2165 24.8580 14.3100 ;
      RECT 24.7240 13.2165 24.7500 14.3100 ;
      RECT 24.6160 13.2165 24.6420 14.3100 ;
      RECT 24.5080 13.2165 24.5340 14.3100 ;
      RECT 24.4000 13.2165 24.4260 14.3100 ;
      RECT 24.2920 13.2165 24.3180 14.3100 ;
      RECT 24.1840 13.2165 24.2100 14.3100 ;
      RECT 24.0760 13.2165 24.1020 14.3100 ;
      RECT 23.9680 13.2165 23.9940 14.3100 ;
      RECT 23.8600 13.2165 23.8860 14.3100 ;
      RECT 23.7520 13.2165 23.7780 14.3100 ;
      RECT 23.6440 13.2165 23.6700 14.3100 ;
      RECT 23.5360 13.2165 23.5620 14.3100 ;
      RECT 23.4280 13.2165 23.4540 14.3100 ;
      RECT 23.3200 13.2165 23.3460 14.3100 ;
      RECT 23.2120 13.2165 23.2380 14.3100 ;
      RECT 23.1040 13.2165 23.1300 14.3100 ;
      RECT 22.9960 13.2165 23.0220 14.3100 ;
      RECT 22.8880 13.2165 22.9140 14.3100 ;
      RECT 22.7800 13.2165 22.8060 14.3100 ;
      RECT 22.6720 13.2165 22.6980 14.3100 ;
      RECT 22.5640 13.2165 22.5900 14.3100 ;
      RECT 22.4560 13.2165 22.4820 14.3100 ;
      RECT 22.3480 13.2165 22.3740 14.3100 ;
      RECT 22.2400 13.2165 22.2660 14.3100 ;
      RECT 22.1320 13.2165 22.1580 14.3100 ;
      RECT 22.0240 13.2165 22.0500 14.3100 ;
      RECT 21.9160 13.2165 21.9420 14.3100 ;
      RECT 21.8080 13.2165 21.8340 14.3100 ;
      RECT 21.7000 13.2165 21.7260 14.3100 ;
      RECT 21.5920 13.2165 21.6180 14.3100 ;
      RECT 21.4840 13.2165 21.5100 14.3100 ;
      RECT 21.3760 13.2165 21.4020 14.3100 ;
      RECT 21.2680 13.2165 21.2940 14.3100 ;
      RECT 21.1600 13.2165 21.1860 14.3100 ;
      RECT 21.0520 13.2165 21.0780 14.3100 ;
      RECT 20.9440 13.2165 20.9700 14.3100 ;
      RECT 20.8360 13.2165 20.8620 14.3100 ;
      RECT 20.7280 13.2165 20.7540 14.3100 ;
      RECT 20.6200 13.2165 20.6460 14.3100 ;
      RECT 20.5120 13.2165 20.5380 14.3100 ;
      RECT 20.4040 13.2165 20.4300 14.3100 ;
      RECT 20.2960 13.2165 20.3220 14.3100 ;
      RECT 20.1880 13.2165 20.2140 14.3100 ;
      RECT 20.0800 13.2165 20.1060 14.3100 ;
      RECT 19.9720 13.2165 19.9980 14.3100 ;
      RECT 19.8640 13.2165 19.8900 14.3100 ;
      RECT 19.7560 13.2165 19.7820 14.3100 ;
      RECT 19.6480 13.2165 19.6740 14.3100 ;
      RECT 19.5400 13.2165 19.5660 14.3100 ;
      RECT 19.4320 13.2165 19.4580 14.3100 ;
      RECT 19.3240 13.2165 19.3500 14.3100 ;
      RECT 19.2160 13.2165 19.2420 14.3100 ;
      RECT 19.1080 13.2165 19.1340 14.3100 ;
      RECT 19.0000 13.2165 19.0260 14.3100 ;
      RECT 18.8920 13.2165 18.9180 14.3100 ;
      RECT 18.7840 13.2165 18.8100 14.3100 ;
      RECT 18.6760 13.2165 18.7020 14.3100 ;
      RECT 18.5680 13.2165 18.5940 14.3100 ;
      RECT 18.4600 13.2165 18.4860 14.3100 ;
      RECT 18.3520 13.2165 18.3780 14.3100 ;
      RECT 18.2440 13.2165 18.2700 14.3100 ;
      RECT 18.1360 13.2165 18.1620 14.3100 ;
      RECT 18.0280 13.2165 18.0540 14.3100 ;
      RECT 17.9200 13.2165 17.9460 14.3100 ;
      RECT 17.8120 13.2165 17.8380 14.3100 ;
      RECT 17.7040 13.2165 17.7300 14.3100 ;
      RECT 17.5960 13.2165 17.6220 14.3100 ;
      RECT 17.4880 13.2165 17.5140 14.3100 ;
      RECT 17.3800 13.2165 17.4060 14.3100 ;
      RECT 17.2720 13.2165 17.2980 14.3100 ;
      RECT 17.1640 13.2165 17.1900 14.3100 ;
      RECT 17.0560 13.2165 17.0820 14.3100 ;
      RECT 16.9480 13.2165 16.9740 14.3100 ;
      RECT 16.8400 13.2165 16.8660 14.3100 ;
      RECT 16.7320 13.2165 16.7580 14.3100 ;
      RECT 16.6240 13.2165 16.6500 14.3100 ;
      RECT 16.5160 13.2165 16.5420 14.3100 ;
      RECT 16.4080 13.2165 16.4340 14.3100 ;
      RECT 16.3000 13.2165 16.3260 14.3100 ;
      RECT 16.0870 13.2165 16.1640 14.3100 ;
      RECT 14.1940 13.2165 14.2710 14.3100 ;
      RECT 14.0320 13.2165 14.0580 14.3100 ;
      RECT 13.9240 13.2165 13.9500 14.3100 ;
      RECT 13.8160 13.2165 13.8420 14.3100 ;
      RECT 13.7080 13.2165 13.7340 14.3100 ;
      RECT 13.6000 13.2165 13.6260 14.3100 ;
      RECT 13.4920 13.2165 13.5180 14.3100 ;
      RECT 13.3840 13.2165 13.4100 14.3100 ;
      RECT 13.2760 13.2165 13.3020 14.3100 ;
      RECT 13.1680 13.2165 13.1940 14.3100 ;
      RECT 13.0600 13.2165 13.0860 14.3100 ;
      RECT 12.9520 13.2165 12.9780 14.3100 ;
      RECT 12.8440 13.2165 12.8700 14.3100 ;
      RECT 12.7360 13.2165 12.7620 14.3100 ;
      RECT 12.6280 13.2165 12.6540 14.3100 ;
      RECT 12.5200 13.2165 12.5460 14.3100 ;
      RECT 12.4120 13.2165 12.4380 14.3100 ;
      RECT 12.3040 13.2165 12.3300 14.3100 ;
      RECT 12.1960 13.2165 12.2220 14.3100 ;
      RECT 12.0880 13.2165 12.1140 14.3100 ;
      RECT 11.9800 13.2165 12.0060 14.3100 ;
      RECT 11.8720 13.2165 11.8980 14.3100 ;
      RECT 11.7640 13.2165 11.7900 14.3100 ;
      RECT 11.6560 13.2165 11.6820 14.3100 ;
      RECT 11.5480 13.2165 11.5740 14.3100 ;
      RECT 11.4400 13.2165 11.4660 14.3100 ;
      RECT 11.3320 13.2165 11.3580 14.3100 ;
      RECT 11.2240 13.2165 11.2500 14.3100 ;
      RECT 11.1160 13.2165 11.1420 14.3100 ;
      RECT 11.0080 13.2165 11.0340 14.3100 ;
      RECT 10.9000 13.2165 10.9260 14.3100 ;
      RECT 10.7920 13.2165 10.8180 14.3100 ;
      RECT 10.6840 13.2165 10.7100 14.3100 ;
      RECT 10.5760 13.2165 10.6020 14.3100 ;
      RECT 10.4680 13.2165 10.4940 14.3100 ;
      RECT 10.3600 13.2165 10.3860 14.3100 ;
      RECT 10.2520 13.2165 10.2780 14.3100 ;
      RECT 10.1440 13.2165 10.1700 14.3100 ;
      RECT 10.0360 13.2165 10.0620 14.3100 ;
      RECT 9.9280 13.2165 9.9540 14.3100 ;
      RECT 9.8200 13.2165 9.8460 14.3100 ;
      RECT 9.7120 13.2165 9.7380 14.3100 ;
      RECT 9.6040 13.2165 9.6300 14.3100 ;
      RECT 9.4960 13.2165 9.5220 14.3100 ;
      RECT 9.3880 13.2165 9.4140 14.3100 ;
      RECT 9.2800 13.2165 9.3060 14.3100 ;
      RECT 9.1720 13.2165 9.1980 14.3100 ;
      RECT 9.0640 13.2165 9.0900 14.3100 ;
      RECT 8.9560 13.2165 8.9820 14.3100 ;
      RECT 8.8480 13.2165 8.8740 14.3100 ;
      RECT 8.7400 13.2165 8.7660 14.3100 ;
      RECT 8.6320 13.2165 8.6580 14.3100 ;
      RECT 8.5240 13.2165 8.5500 14.3100 ;
      RECT 8.4160 13.2165 8.4420 14.3100 ;
      RECT 8.3080 13.2165 8.3340 14.3100 ;
      RECT 8.2000 13.2165 8.2260 14.3100 ;
      RECT 8.0920 13.2165 8.1180 14.3100 ;
      RECT 7.9840 13.2165 8.0100 14.3100 ;
      RECT 7.8760 13.2165 7.9020 14.3100 ;
      RECT 7.7680 13.2165 7.7940 14.3100 ;
      RECT 7.6600 13.2165 7.6860 14.3100 ;
      RECT 7.5520 13.2165 7.5780 14.3100 ;
      RECT 7.4440 13.2165 7.4700 14.3100 ;
      RECT 7.3360 13.2165 7.3620 14.3100 ;
      RECT 7.2280 13.2165 7.2540 14.3100 ;
      RECT 7.1200 13.2165 7.1460 14.3100 ;
      RECT 7.0120 13.2165 7.0380 14.3100 ;
      RECT 6.9040 13.2165 6.9300 14.3100 ;
      RECT 6.7960 13.2165 6.8220 14.3100 ;
      RECT 6.6880 13.2165 6.7140 14.3100 ;
      RECT 6.5800 13.2165 6.6060 14.3100 ;
      RECT 6.4720 13.2165 6.4980 14.3100 ;
      RECT 6.3640 13.2165 6.3900 14.3100 ;
      RECT 6.2560 13.2165 6.2820 14.3100 ;
      RECT 6.1480 13.2165 6.1740 14.3100 ;
      RECT 6.0400 13.2165 6.0660 14.3100 ;
      RECT 5.9320 13.2165 5.9580 14.3100 ;
      RECT 5.8240 13.2165 5.8500 14.3100 ;
      RECT 5.7160 13.2165 5.7420 14.3100 ;
      RECT 5.6080 13.2165 5.6340 14.3100 ;
      RECT 5.5000 13.2165 5.5260 14.3100 ;
      RECT 5.3920 13.2165 5.4180 14.3100 ;
      RECT 5.2840 13.2165 5.3100 14.3100 ;
      RECT 5.1760 13.2165 5.2020 14.3100 ;
      RECT 5.0680 13.2165 5.0940 14.3100 ;
      RECT 4.9600 13.2165 4.9860 14.3100 ;
      RECT 4.8520 13.2165 4.8780 14.3100 ;
      RECT 4.7440 13.2165 4.7700 14.3100 ;
      RECT 4.6360 13.2165 4.6620 14.3100 ;
      RECT 4.5280 13.2165 4.5540 14.3100 ;
      RECT 4.4200 13.2165 4.4460 14.3100 ;
      RECT 4.3120 13.2165 4.3380 14.3100 ;
      RECT 4.2040 13.2165 4.2300 14.3100 ;
      RECT 4.0960 13.2165 4.1220 14.3100 ;
      RECT 3.9880 13.2165 4.0140 14.3100 ;
      RECT 3.8800 13.2165 3.9060 14.3100 ;
      RECT 3.7720 13.2165 3.7980 14.3100 ;
      RECT 3.6640 13.2165 3.6900 14.3100 ;
      RECT 3.5560 13.2165 3.5820 14.3100 ;
      RECT 3.4480 13.2165 3.4740 14.3100 ;
      RECT 3.3400 13.2165 3.3660 14.3100 ;
      RECT 3.2320 13.2165 3.2580 14.3100 ;
      RECT 3.1240 13.2165 3.1500 14.3100 ;
      RECT 3.0160 13.2165 3.0420 14.3100 ;
      RECT 2.9080 13.2165 2.9340 14.3100 ;
      RECT 2.8000 13.2165 2.8260 14.3100 ;
      RECT 2.6920 13.2165 2.7180 14.3100 ;
      RECT 2.5840 13.2165 2.6100 14.3100 ;
      RECT 2.4760 13.2165 2.5020 14.3100 ;
      RECT 2.3680 13.2165 2.3940 14.3100 ;
      RECT 2.2600 13.2165 2.2860 14.3100 ;
      RECT 2.1520 13.2165 2.1780 14.3100 ;
      RECT 2.0440 13.2165 2.0700 14.3100 ;
      RECT 1.9360 13.2165 1.9620 14.3100 ;
      RECT 1.8280 13.2165 1.8540 14.3100 ;
      RECT 1.7200 13.2165 1.7460 14.3100 ;
      RECT 1.6120 13.2165 1.6380 14.3100 ;
      RECT 1.5040 13.2165 1.5300 14.3100 ;
      RECT 1.3960 13.2165 1.4220 14.3100 ;
      RECT 1.2880 13.2165 1.3140 14.3100 ;
      RECT 1.1800 13.2165 1.2060 14.3100 ;
      RECT 1.0720 13.2165 1.0980 14.3100 ;
      RECT 0.9640 13.2165 0.9900 14.3100 ;
      RECT 0.8560 13.2165 0.8820 14.3100 ;
      RECT 0.7480 13.2165 0.7740 14.3100 ;
      RECT 0.6400 13.2165 0.6660 14.3100 ;
      RECT 0.5320 13.2165 0.5580 14.3100 ;
      RECT 0.4240 13.2165 0.4500 14.3100 ;
      RECT 0.3160 13.2165 0.3420 14.3100 ;
      RECT 0.2080 13.2165 0.2340 14.3100 ;
      RECT 0.0050 13.2165 0.0900 14.3100 ;
      RECT 15.5530 14.2965 15.6810 15.3900 ;
      RECT 15.5390 14.9620 15.6810 15.2845 ;
      RECT 15.3190 14.6890 15.4530 15.3900 ;
      RECT 15.2960 15.0240 15.4530 15.2820 ;
      RECT 15.3190 14.2965 15.4170 15.3900 ;
      RECT 15.3190 14.4175 15.4310 14.6570 ;
      RECT 15.3190 14.2965 15.4530 14.3855 ;
      RECT 15.0940 14.7470 15.2280 15.3900 ;
      RECT 15.0940 14.2965 15.1920 15.3900 ;
      RECT 14.6770 14.2965 14.7600 15.3900 ;
      RECT 14.6770 14.3850 14.7740 15.3205 ;
      RECT 30.2680 14.2965 30.3530 15.3900 ;
      RECT 30.1240 14.2965 30.1500 15.3900 ;
      RECT 30.0160 14.2965 30.0420 15.3900 ;
      RECT 29.9080 14.2965 29.9340 15.3900 ;
      RECT 29.8000 14.2965 29.8260 15.3900 ;
      RECT 29.6920 14.2965 29.7180 15.3900 ;
      RECT 29.5840 14.2965 29.6100 15.3900 ;
      RECT 29.4760 14.2965 29.5020 15.3900 ;
      RECT 29.3680 14.2965 29.3940 15.3900 ;
      RECT 29.2600 14.2965 29.2860 15.3900 ;
      RECT 29.1520 14.2965 29.1780 15.3900 ;
      RECT 29.0440 14.2965 29.0700 15.3900 ;
      RECT 28.9360 14.2965 28.9620 15.3900 ;
      RECT 28.8280 14.2965 28.8540 15.3900 ;
      RECT 28.7200 14.2965 28.7460 15.3900 ;
      RECT 28.6120 14.2965 28.6380 15.3900 ;
      RECT 28.5040 14.2965 28.5300 15.3900 ;
      RECT 28.3960 14.2965 28.4220 15.3900 ;
      RECT 28.2880 14.2965 28.3140 15.3900 ;
      RECT 28.1800 14.2965 28.2060 15.3900 ;
      RECT 28.0720 14.2965 28.0980 15.3900 ;
      RECT 27.9640 14.2965 27.9900 15.3900 ;
      RECT 27.8560 14.2965 27.8820 15.3900 ;
      RECT 27.7480 14.2965 27.7740 15.3900 ;
      RECT 27.6400 14.2965 27.6660 15.3900 ;
      RECT 27.5320 14.2965 27.5580 15.3900 ;
      RECT 27.4240 14.2965 27.4500 15.3900 ;
      RECT 27.3160 14.2965 27.3420 15.3900 ;
      RECT 27.2080 14.2965 27.2340 15.3900 ;
      RECT 27.1000 14.2965 27.1260 15.3900 ;
      RECT 26.9920 14.2965 27.0180 15.3900 ;
      RECT 26.8840 14.2965 26.9100 15.3900 ;
      RECT 26.7760 14.2965 26.8020 15.3900 ;
      RECT 26.6680 14.2965 26.6940 15.3900 ;
      RECT 26.5600 14.2965 26.5860 15.3900 ;
      RECT 26.4520 14.2965 26.4780 15.3900 ;
      RECT 26.3440 14.2965 26.3700 15.3900 ;
      RECT 26.2360 14.2965 26.2620 15.3900 ;
      RECT 26.1280 14.2965 26.1540 15.3900 ;
      RECT 26.0200 14.2965 26.0460 15.3900 ;
      RECT 25.9120 14.2965 25.9380 15.3900 ;
      RECT 25.8040 14.2965 25.8300 15.3900 ;
      RECT 25.6960 14.2965 25.7220 15.3900 ;
      RECT 25.5880 14.2965 25.6140 15.3900 ;
      RECT 25.4800 14.2965 25.5060 15.3900 ;
      RECT 25.3720 14.2965 25.3980 15.3900 ;
      RECT 25.2640 14.2965 25.2900 15.3900 ;
      RECT 25.1560 14.2965 25.1820 15.3900 ;
      RECT 25.0480 14.2965 25.0740 15.3900 ;
      RECT 24.9400 14.2965 24.9660 15.3900 ;
      RECT 24.8320 14.2965 24.8580 15.3900 ;
      RECT 24.7240 14.2965 24.7500 15.3900 ;
      RECT 24.6160 14.2965 24.6420 15.3900 ;
      RECT 24.5080 14.2965 24.5340 15.3900 ;
      RECT 24.4000 14.2965 24.4260 15.3900 ;
      RECT 24.2920 14.2965 24.3180 15.3900 ;
      RECT 24.1840 14.2965 24.2100 15.3900 ;
      RECT 24.0760 14.2965 24.1020 15.3900 ;
      RECT 23.9680 14.2965 23.9940 15.3900 ;
      RECT 23.8600 14.2965 23.8860 15.3900 ;
      RECT 23.7520 14.2965 23.7780 15.3900 ;
      RECT 23.6440 14.2965 23.6700 15.3900 ;
      RECT 23.5360 14.2965 23.5620 15.3900 ;
      RECT 23.4280 14.2965 23.4540 15.3900 ;
      RECT 23.3200 14.2965 23.3460 15.3900 ;
      RECT 23.2120 14.2965 23.2380 15.3900 ;
      RECT 23.1040 14.2965 23.1300 15.3900 ;
      RECT 22.9960 14.2965 23.0220 15.3900 ;
      RECT 22.8880 14.2965 22.9140 15.3900 ;
      RECT 22.7800 14.2965 22.8060 15.3900 ;
      RECT 22.6720 14.2965 22.6980 15.3900 ;
      RECT 22.5640 14.2965 22.5900 15.3900 ;
      RECT 22.4560 14.2965 22.4820 15.3900 ;
      RECT 22.3480 14.2965 22.3740 15.3900 ;
      RECT 22.2400 14.2965 22.2660 15.3900 ;
      RECT 22.1320 14.2965 22.1580 15.3900 ;
      RECT 22.0240 14.2965 22.0500 15.3900 ;
      RECT 21.9160 14.2965 21.9420 15.3900 ;
      RECT 21.8080 14.2965 21.8340 15.3900 ;
      RECT 21.7000 14.2965 21.7260 15.3900 ;
      RECT 21.5920 14.2965 21.6180 15.3900 ;
      RECT 21.4840 14.2965 21.5100 15.3900 ;
      RECT 21.3760 14.2965 21.4020 15.3900 ;
      RECT 21.2680 14.2965 21.2940 15.3900 ;
      RECT 21.1600 14.2965 21.1860 15.3900 ;
      RECT 21.0520 14.2965 21.0780 15.3900 ;
      RECT 20.9440 14.2965 20.9700 15.3900 ;
      RECT 20.8360 14.2965 20.8620 15.3900 ;
      RECT 20.7280 14.2965 20.7540 15.3900 ;
      RECT 20.6200 14.2965 20.6460 15.3900 ;
      RECT 20.5120 14.2965 20.5380 15.3900 ;
      RECT 20.4040 14.2965 20.4300 15.3900 ;
      RECT 20.2960 14.2965 20.3220 15.3900 ;
      RECT 20.1880 14.2965 20.2140 15.3900 ;
      RECT 20.0800 14.2965 20.1060 15.3900 ;
      RECT 19.9720 14.2965 19.9980 15.3900 ;
      RECT 19.8640 14.2965 19.8900 15.3900 ;
      RECT 19.7560 14.2965 19.7820 15.3900 ;
      RECT 19.6480 14.2965 19.6740 15.3900 ;
      RECT 19.5400 14.2965 19.5660 15.3900 ;
      RECT 19.4320 14.2965 19.4580 15.3900 ;
      RECT 19.3240 14.2965 19.3500 15.3900 ;
      RECT 19.2160 14.2965 19.2420 15.3900 ;
      RECT 19.1080 14.2965 19.1340 15.3900 ;
      RECT 19.0000 14.2965 19.0260 15.3900 ;
      RECT 18.8920 14.2965 18.9180 15.3900 ;
      RECT 18.7840 14.2965 18.8100 15.3900 ;
      RECT 18.6760 14.2965 18.7020 15.3900 ;
      RECT 18.5680 14.2965 18.5940 15.3900 ;
      RECT 18.4600 14.2965 18.4860 15.3900 ;
      RECT 18.3520 14.2965 18.3780 15.3900 ;
      RECT 18.2440 14.2965 18.2700 15.3900 ;
      RECT 18.1360 14.2965 18.1620 15.3900 ;
      RECT 18.0280 14.2965 18.0540 15.3900 ;
      RECT 17.9200 14.2965 17.9460 15.3900 ;
      RECT 17.8120 14.2965 17.8380 15.3900 ;
      RECT 17.7040 14.2965 17.7300 15.3900 ;
      RECT 17.5960 14.2965 17.6220 15.3900 ;
      RECT 17.4880 14.2965 17.5140 15.3900 ;
      RECT 17.3800 14.2965 17.4060 15.3900 ;
      RECT 17.2720 14.2965 17.2980 15.3900 ;
      RECT 17.1640 14.2965 17.1900 15.3900 ;
      RECT 17.0560 14.2965 17.0820 15.3900 ;
      RECT 16.9480 14.2965 16.9740 15.3900 ;
      RECT 16.8400 14.2965 16.8660 15.3900 ;
      RECT 16.7320 14.2965 16.7580 15.3900 ;
      RECT 16.6240 14.2965 16.6500 15.3900 ;
      RECT 16.5160 14.2965 16.5420 15.3900 ;
      RECT 16.4080 14.2965 16.4340 15.3900 ;
      RECT 16.3000 14.2965 16.3260 15.3900 ;
      RECT 16.0870 14.2965 16.1640 15.3900 ;
      RECT 14.1940 14.2965 14.2710 15.3900 ;
      RECT 14.0320 14.2965 14.0580 15.3900 ;
      RECT 13.9240 14.2965 13.9500 15.3900 ;
      RECT 13.8160 14.2965 13.8420 15.3900 ;
      RECT 13.7080 14.2965 13.7340 15.3900 ;
      RECT 13.6000 14.2965 13.6260 15.3900 ;
      RECT 13.4920 14.2965 13.5180 15.3900 ;
      RECT 13.3840 14.2965 13.4100 15.3900 ;
      RECT 13.2760 14.2965 13.3020 15.3900 ;
      RECT 13.1680 14.2965 13.1940 15.3900 ;
      RECT 13.0600 14.2965 13.0860 15.3900 ;
      RECT 12.9520 14.2965 12.9780 15.3900 ;
      RECT 12.8440 14.2965 12.8700 15.3900 ;
      RECT 12.7360 14.2965 12.7620 15.3900 ;
      RECT 12.6280 14.2965 12.6540 15.3900 ;
      RECT 12.5200 14.2965 12.5460 15.3900 ;
      RECT 12.4120 14.2965 12.4380 15.3900 ;
      RECT 12.3040 14.2965 12.3300 15.3900 ;
      RECT 12.1960 14.2965 12.2220 15.3900 ;
      RECT 12.0880 14.2965 12.1140 15.3900 ;
      RECT 11.9800 14.2965 12.0060 15.3900 ;
      RECT 11.8720 14.2965 11.8980 15.3900 ;
      RECT 11.7640 14.2965 11.7900 15.3900 ;
      RECT 11.6560 14.2965 11.6820 15.3900 ;
      RECT 11.5480 14.2965 11.5740 15.3900 ;
      RECT 11.4400 14.2965 11.4660 15.3900 ;
      RECT 11.3320 14.2965 11.3580 15.3900 ;
      RECT 11.2240 14.2965 11.2500 15.3900 ;
      RECT 11.1160 14.2965 11.1420 15.3900 ;
      RECT 11.0080 14.2965 11.0340 15.3900 ;
      RECT 10.9000 14.2965 10.9260 15.3900 ;
      RECT 10.7920 14.2965 10.8180 15.3900 ;
      RECT 10.6840 14.2965 10.7100 15.3900 ;
      RECT 10.5760 14.2965 10.6020 15.3900 ;
      RECT 10.4680 14.2965 10.4940 15.3900 ;
      RECT 10.3600 14.2965 10.3860 15.3900 ;
      RECT 10.2520 14.2965 10.2780 15.3900 ;
      RECT 10.1440 14.2965 10.1700 15.3900 ;
      RECT 10.0360 14.2965 10.0620 15.3900 ;
      RECT 9.9280 14.2965 9.9540 15.3900 ;
      RECT 9.8200 14.2965 9.8460 15.3900 ;
      RECT 9.7120 14.2965 9.7380 15.3900 ;
      RECT 9.6040 14.2965 9.6300 15.3900 ;
      RECT 9.4960 14.2965 9.5220 15.3900 ;
      RECT 9.3880 14.2965 9.4140 15.3900 ;
      RECT 9.2800 14.2965 9.3060 15.3900 ;
      RECT 9.1720 14.2965 9.1980 15.3900 ;
      RECT 9.0640 14.2965 9.0900 15.3900 ;
      RECT 8.9560 14.2965 8.9820 15.3900 ;
      RECT 8.8480 14.2965 8.8740 15.3900 ;
      RECT 8.7400 14.2965 8.7660 15.3900 ;
      RECT 8.6320 14.2965 8.6580 15.3900 ;
      RECT 8.5240 14.2965 8.5500 15.3900 ;
      RECT 8.4160 14.2965 8.4420 15.3900 ;
      RECT 8.3080 14.2965 8.3340 15.3900 ;
      RECT 8.2000 14.2965 8.2260 15.3900 ;
      RECT 8.0920 14.2965 8.1180 15.3900 ;
      RECT 7.9840 14.2965 8.0100 15.3900 ;
      RECT 7.8760 14.2965 7.9020 15.3900 ;
      RECT 7.7680 14.2965 7.7940 15.3900 ;
      RECT 7.6600 14.2965 7.6860 15.3900 ;
      RECT 7.5520 14.2965 7.5780 15.3900 ;
      RECT 7.4440 14.2965 7.4700 15.3900 ;
      RECT 7.3360 14.2965 7.3620 15.3900 ;
      RECT 7.2280 14.2965 7.2540 15.3900 ;
      RECT 7.1200 14.2965 7.1460 15.3900 ;
      RECT 7.0120 14.2965 7.0380 15.3900 ;
      RECT 6.9040 14.2965 6.9300 15.3900 ;
      RECT 6.7960 14.2965 6.8220 15.3900 ;
      RECT 6.6880 14.2965 6.7140 15.3900 ;
      RECT 6.5800 14.2965 6.6060 15.3900 ;
      RECT 6.4720 14.2965 6.4980 15.3900 ;
      RECT 6.3640 14.2965 6.3900 15.3900 ;
      RECT 6.2560 14.2965 6.2820 15.3900 ;
      RECT 6.1480 14.2965 6.1740 15.3900 ;
      RECT 6.0400 14.2965 6.0660 15.3900 ;
      RECT 5.9320 14.2965 5.9580 15.3900 ;
      RECT 5.8240 14.2965 5.8500 15.3900 ;
      RECT 5.7160 14.2965 5.7420 15.3900 ;
      RECT 5.6080 14.2965 5.6340 15.3900 ;
      RECT 5.5000 14.2965 5.5260 15.3900 ;
      RECT 5.3920 14.2965 5.4180 15.3900 ;
      RECT 5.2840 14.2965 5.3100 15.3900 ;
      RECT 5.1760 14.2965 5.2020 15.3900 ;
      RECT 5.0680 14.2965 5.0940 15.3900 ;
      RECT 4.9600 14.2965 4.9860 15.3900 ;
      RECT 4.8520 14.2965 4.8780 15.3900 ;
      RECT 4.7440 14.2965 4.7700 15.3900 ;
      RECT 4.6360 14.2965 4.6620 15.3900 ;
      RECT 4.5280 14.2965 4.5540 15.3900 ;
      RECT 4.4200 14.2965 4.4460 15.3900 ;
      RECT 4.3120 14.2965 4.3380 15.3900 ;
      RECT 4.2040 14.2965 4.2300 15.3900 ;
      RECT 4.0960 14.2965 4.1220 15.3900 ;
      RECT 3.9880 14.2965 4.0140 15.3900 ;
      RECT 3.8800 14.2965 3.9060 15.3900 ;
      RECT 3.7720 14.2965 3.7980 15.3900 ;
      RECT 3.6640 14.2965 3.6900 15.3900 ;
      RECT 3.5560 14.2965 3.5820 15.3900 ;
      RECT 3.4480 14.2965 3.4740 15.3900 ;
      RECT 3.3400 14.2965 3.3660 15.3900 ;
      RECT 3.2320 14.2965 3.2580 15.3900 ;
      RECT 3.1240 14.2965 3.1500 15.3900 ;
      RECT 3.0160 14.2965 3.0420 15.3900 ;
      RECT 2.9080 14.2965 2.9340 15.3900 ;
      RECT 2.8000 14.2965 2.8260 15.3900 ;
      RECT 2.6920 14.2965 2.7180 15.3900 ;
      RECT 2.5840 14.2965 2.6100 15.3900 ;
      RECT 2.4760 14.2965 2.5020 15.3900 ;
      RECT 2.3680 14.2965 2.3940 15.3900 ;
      RECT 2.2600 14.2965 2.2860 15.3900 ;
      RECT 2.1520 14.2965 2.1780 15.3900 ;
      RECT 2.0440 14.2965 2.0700 15.3900 ;
      RECT 1.9360 14.2965 1.9620 15.3900 ;
      RECT 1.8280 14.2965 1.8540 15.3900 ;
      RECT 1.7200 14.2965 1.7460 15.3900 ;
      RECT 1.6120 14.2965 1.6380 15.3900 ;
      RECT 1.5040 14.2965 1.5300 15.3900 ;
      RECT 1.3960 14.2965 1.4220 15.3900 ;
      RECT 1.2880 14.2965 1.3140 15.3900 ;
      RECT 1.1800 14.2965 1.2060 15.3900 ;
      RECT 1.0720 14.2965 1.0980 15.3900 ;
      RECT 0.9640 14.2965 0.9900 15.3900 ;
      RECT 0.8560 14.2965 0.8820 15.3900 ;
      RECT 0.7480 14.2965 0.7740 15.3900 ;
      RECT 0.6400 14.2965 0.6660 15.3900 ;
      RECT 0.5320 14.2965 0.5580 15.3900 ;
      RECT 0.4240 14.2965 0.4500 15.3900 ;
      RECT 0.3160 14.2965 0.3420 15.3900 ;
      RECT 0.2080 14.2965 0.2340 15.3900 ;
      RECT 0.0050 14.2965 0.0900 15.3900 ;
      RECT 15.5530 15.3765 15.6810 16.4700 ;
      RECT 15.5390 16.0420 15.6810 16.3645 ;
      RECT 15.3190 15.7690 15.4530 16.4700 ;
      RECT 15.2960 16.1040 15.4530 16.3620 ;
      RECT 15.3190 15.3765 15.4170 16.4700 ;
      RECT 15.3190 15.4975 15.4310 15.7370 ;
      RECT 15.3190 15.3765 15.4530 15.4655 ;
      RECT 15.0940 15.8270 15.2280 16.4700 ;
      RECT 15.0940 15.3765 15.1920 16.4700 ;
      RECT 14.6770 15.3765 14.7600 16.4700 ;
      RECT 14.6770 15.4650 14.7740 16.4005 ;
      RECT 30.2680 15.3765 30.3530 16.4700 ;
      RECT 30.1240 15.3765 30.1500 16.4700 ;
      RECT 30.0160 15.3765 30.0420 16.4700 ;
      RECT 29.9080 15.3765 29.9340 16.4700 ;
      RECT 29.8000 15.3765 29.8260 16.4700 ;
      RECT 29.6920 15.3765 29.7180 16.4700 ;
      RECT 29.5840 15.3765 29.6100 16.4700 ;
      RECT 29.4760 15.3765 29.5020 16.4700 ;
      RECT 29.3680 15.3765 29.3940 16.4700 ;
      RECT 29.2600 15.3765 29.2860 16.4700 ;
      RECT 29.1520 15.3765 29.1780 16.4700 ;
      RECT 29.0440 15.3765 29.0700 16.4700 ;
      RECT 28.9360 15.3765 28.9620 16.4700 ;
      RECT 28.8280 15.3765 28.8540 16.4700 ;
      RECT 28.7200 15.3765 28.7460 16.4700 ;
      RECT 28.6120 15.3765 28.6380 16.4700 ;
      RECT 28.5040 15.3765 28.5300 16.4700 ;
      RECT 28.3960 15.3765 28.4220 16.4700 ;
      RECT 28.2880 15.3765 28.3140 16.4700 ;
      RECT 28.1800 15.3765 28.2060 16.4700 ;
      RECT 28.0720 15.3765 28.0980 16.4700 ;
      RECT 27.9640 15.3765 27.9900 16.4700 ;
      RECT 27.8560 15.3765 27.8820 16.4700 ;
      RECT 27.7480 15.3765 27.7740 16.4700 ;
      RECT 27.6400 15.3765 27.6660 16.4700 ;
      RECT 27.5320 15.3765 27.5580 16.4700 ;
      RECT 27.4240 15.3765 27.4500 16.4700 ;
      RECT 27.3160 15.3765 27.3420 16.4700 ;
      RECT 27.2080 15.3765 27.2340 16.4700 ;
      RECT 27.1000 15.3765 27.1260 16.4700 ;
      RECT 26.9920 15.3765 27.0180 16.4700 ;
      RECT 26.8840 15.3765 26.9100 16.4700 ;
      RECT 26.7760 15.3765 26.8020 16.4700 ;
      RECT 26.6680 15.3765 26.6940 16.4700 ;
      RECT 26.5600 15.3765 26.5860 16.4700 ;
      RECT 26.4520 15.3765 26.4780 16.4700 ;
      RECT 26.3440 15.3765 26.3700 16.4700 ;
      RECT 26.2360 15.3765 26.2620 16.4700 ;
      RECT 26.1280 15.3765 26.1540 16.4700 ;
      RECT 26.0200 15.3765 26.0460 16.4700 ;
      RECT 25.9120 15.3765 25.9380 16.4700 ;
      RECT 25.8040 15.3765 25.8300 16.4700 ;
      RECT 25.6960 15.3765 25.7220 16.4700 ;
      RECT 25.5880 15.3765 25.6140 16.4700 ;
      RECT 25.4800 15.3765 25.5060 16.4700 ;
      RECT 25.3720 15.3765 25.3980 16.4700 ;
      RECT 25.2640 15.3765 25.2900 16.4700 ;
      RECT 25.1560 15.3765 25.1820 16.4700 ;
      RECT 25.0480 15.3765 25.0740 16.4700 ;
      RECT 24.9400 15.3765 24.9660 16.4700 ;
      RECT 24.8320 15.3765 24.8580 16.4700 ;
      RECT 24.7240 15.3765 24.7500 16.4700 ;
      RECT 24.6160 15.3765 24.6420 16.4700 ;
      RECT 24.5080 15.3765 24.5340 16.4700 ;
      RECT 24.4000 15.3765 24.4260 16.4700 ;
      RECT 24.2920 15.3765 24.3180 16.4700 ;
      RECT 24.1840 15.3765 24.2100 16.4700 ;
      RECT 24.0760 15.3765 24.1020 16.4700 ;
      RECT 23.9680 15.3765 23.9940 16.4700 ;
      RECT 23.8600 15.3765 23.8860 16.4700 ;
      RECT 23.7520 15.3765 23.7780 16.4700 ;
      RECT 23.6440 15.3765 23.6700 16.4700 ;
      RECT 23.5360 15.3765 23.5620 16.4700 ;
      RECT 23.4280 15.3765 23.4540 16.4700 ;
      RECT 23.3200 15.3765 23.3460 16.4700 ;
      RECT 23.2120 15.3765 23.2380 16.4700 ;
      RECT 23.1040 15.3765 23.1300 16.4700 ;
      RECT 22.9960 15.3765 23.0220 16.4700 ;
      RECT 22.8880 15.3765 22.9140 16.4700 ;
      RECT 22.7800 15.3765 22.8060 16.4700 ;
      RECT 22.6720 15.3765 22.6980 16.4700 ;
      RECT 22.5640 15.3765 22.5900 16.4700 ;
      RECT 22.4560 15.3765 22.4820 16.4700 ;
      RECT 22.3480 15.3765 22.3740 16.4700 ;
      RECT 22.2400 15.3765 22.2660 16.4700 ;
      RECT 22.1320 15.3765 22.1580 16.4700 ;
      RECT 22.0240 15.3765 22.0500 16.4700 ;
      RECT 21.9160 15.3765 21.9420 16.4700 ;
      RECT 21.8080 15.3765 21.8340 16.4700 ;
      RECT 21.7000 15.3765 21.7260 16.4700 ;
      RECT 21.5920 15.3765 21.6180 16.4700 ;
      RECT 21.4840 15.3765 21.5100 16.4700 ;
      RECT 21.3760 15.3765 21.4020 16.4700 ;
      RECT 21.2680 15.3765 21.2940 16.4700 ;
      RECT 21.1600 15.3765 21.1860 16.4700 ;
      RECT 21.0520 15.3765 21.0780 16.4700 ;
      RECT 20.9440 15.3765 20.9700 16.4700 ;
      RECT 20.8360 15.3765 20.8620 16.4700 ;
      RECT 20.7280 15.3765 20.7540 16.4700 ;
      RECT 20.6200 15.3765 20.6460 16.4700 ;
      RECT 20.5120 15.3765 20.5380 16.4700 ;
      RECT 20.4040 15.3765 20.4300 16.4700 ;
      RECT 20.2960 15.3765 20.3220 16.4700 ;
      RECT 20.1880 15.3765 20.2140 16.4700 ;
      RECT 20.0800 15.3765 20.1060 16.4700 ;
      RECT 19.9720 15.3765 19.9980 16.4700 ;
      RECT 19.8640 15.3765 19.8900 16.4700 ;
      RECT 19.7560 15.3765 19.7820 16.4700 ;
      RECT 19.6480 15.3765 19.6740 16.4700 ;
      RECT 19.5400 15.3765 19.5660 16.4700 ;
      RECT 19.4320 15.3765 19.4580 16.4700 ;
      RECT 19.3240 15.3765 19.3500 16.4700 ;
      RECT 19.2160 15.3765 19.2420 16.4700 ;
      RECT 19.1080 15.3765 19.1340 16.4700 ;
      RECT 19.0000 15.3765 19.0260 16.4700 ;
      RECT 18.8920 15.3765 18.9180 16.4700 ;
      RECT 18.7840 15.3765 18.8100 16.4700 ;
      RECT 18.6760 15.3765 18.7020 16.4700 ;
      RECT 18.5680 15.3765 18.5940 16.4700 ;
      RECT 18.4600 15.3765 18.4860 16.4700 ;
      RECT 18.3520 15.3765 18.3780 16.4700 ;
      RECT 18.2440 15.3765 18.2700 16.4700 ;
      RECT 18.1360 15.3765 18.1620 16.4700 ;
      RECT 18.0280 15.3765 18.0540 16.4700 ;
      RECT 17.9200 15.3765 17.9460 16.4700 ;
      RECT 17.8120 15.3765 17.8380 16.4700 ;
      RECT 17.7040 15.3765 17.7300 16.4700 ;
      RECT 17.5960 15.3765 17.6220 16.4700 ;
      RECT 17.4880 15.3765 17.5140 16.4700 ;
      RECT 17.3800 15.3765 17.4060 16.4700 ;
      RECT 17.2720 15.3765 17.2980 16.4700 ;
      RECT 17.1640 15.3765 17.1900 16.4700 ;
      RECT 17.0560 15.3765 17.0820 16.4700 ;
      RECT 16.9480 15.3765 16.9740 16.4700 ;
      RECT 16.8400 15.3765 16.8660 16.4700 ;
      RECT 16.7320 15.3765 16.7580 16.4700 ;
      RECT 16.6240 15.3765 16.6500 16.4700 ;
      RECT 16.5160 15.3765 16.5420 16.4700 ;
      RECT 16.4080 15.3765 16.4340 16.4700 ;
      RECT 16.3000 15.3765 16.3260 16.4700 ;
      RECT 16.0870 15.3765 16.1640 16.4700 ;
      RECT 14.1940 15.3765 14.2710 16.4700 ;
      RECT 14.0320 15.3765 14.0580 16.4700 ;
      RECT 13.9240 15.3765 13.9500 16.4700 ;
      RECT 13.8160 15.3765 13.8420 16.4700 ;
      RECT 13.7080 15.3765 13.7340 16.4700 ;
      RECT 13.6000 15.3765 13.6260 16.4700 ;
      RECT 13.4920 15.3765 13.5180 16.4700 ;
      RECT 13.3840 15.3765 13.4100 16.4700 ;
      RECT 13.2760 15.3765 13.3020 16.4700 ;
      RECT 13.1680 15.3765 13.1940 16.4700 ;
      RECT 13.0600 15.3765 13.0860 16.4700 ;
      RECT 12.9520 15.3765 12.9780 16.4700 ;
      RECT 12.8440 15.3765 12.8700 16.4700 ;
      RECT 12.7360 15.3765 12.7620 16.4700 ;
      RECT 12.6280 15.3765 12.6540 16.4700 ;
      RECT 12.5200 15.3765 12.5460 16.4700 ;
      RECT 12.4120 15.3765 12.4380 16.4700 ;
      RECT 12.3040 15.3765 12.3300 16.4700 ;
      RECT 12.1960 15.3765 12.2220 16.4700 ;
      RECT 12.0880 15.3765 12.1140 16.4700 ;
      RECT 11.9800 15.3765 12.0060 16.4700 ;
      RECT 11.8720 15.3765 11.8980 16.4700 ;
      RECT 11.7640 15.3765 11.7900 16.4700 ;
      RECT 11.6560 15.3765 11.6820 16.4700 ;
      RECT 11.5480 15.3765 11.5740 16.4700 ;
      RECT 11.4400 15.3765 11.4660 16.4700 ;
      RECT 11.3320 15.3765 11.3580 16.4700 ;
      RECT 11.2240 15.3765 11.2500 16.4700 ;
      RECT 11.1160 15.3765 11.1420 16.4700 ;
      RECT 11.0080 15.3765 11.0340 16.4700 ;
      RECT 10.9000 15.3765 10.9260 16.4700 ;
      RECT 10.7920 15.3765 10.8180 16.4700 ;
      RECT 10.6840 15.3765 10.7100 16.4700 ;
      RECT 10.5760 15.3765 10.6020 16.4700 ;
      RECT 10.4680 15.3765 10.4940 16.4700 ;
      RECT 10.3600 15.3765 10.3860 16.4700 ;
      RECT 10.2520 15.3765 10.2780 16.4700 ;
      RECT 10.1440 15.3765 10.1700 16.4700 ;
      RECT 10.0360 15.3765 10.0620 16.4700 ;
      RECT 9.9280 15.3765 9.9540 16.4700 ;
      RECT 9.8200 15.3765 9.8460 16.4700 ;
      RECT 9.7120 15.3765 9.7380 16.4700 ;
      RECT 9.6040 15.3765 9.6300 16.4700 ;
      RECT 9.4960 15.3765 9.5220 16.4700 ;
      RECT 9.3880 15.3765 9.4140 16.4700 ;
      RECT 9.2800 15.3765 9.3060 16.4700 ;
      RECT 9.1720 15.3765 9.1980 16.4700 ;
      RECT 9.0640 15.3765 9.0900 16.4700 ;
      RECT 8.9560 15.3765 8.9820 16.4700 ;
      RECT 8.8480 15.3765 8.8740 16.4700 ;
      RECT 8.7400 15.3765 8.7660 16.4700 ;
      RECT 8.6320 15.3765 8.6580 16.4700 ;
      RECT 8.5240 15.3765 8.5500 16.4700 ;
      RECT 8.4160 15.3765 8.4420 16.4700 ;
      RECT 8.3080 15.3765 8.3340 16.4700 ;
      RECT 8.2000 15.3765 8.2260 16.4700 ;
      RECT 8.0920 15.3765 8.1180 16.4700 ;
      RECT 7.9840 15.3765 8.0100 16.4700 ;
      RECT 7.8760 15.3765 7.9020 16.4700 ;
      RECT 7.7680 15.3765 7.7940 16.4700 ;
      RECT 7.6600 15.3765 7.6860 16.4700 ;
      RECT 7.5520 15.3765 7.5780 16.4700 ;
      RECT 7.4440 15.3765 7.4700 16.4700 ;
      RECT 7.3360 15.3765 7.3620 16.4700 ;
      RECT 7.2280 15.3765 7.2540 16.4700 ;
      RECT 7.1200 15.3765 7.1460 16.4700 ;
      RECT 7.0120 15.3765 7.0380 16.4700 ;
      RECT 6.9040 15.3765 6.9300 16.4700 ;
      RECT 6.7960 15.3765 6.8220 16.4700 ;
      RECT 6.6880 15.3765 6.7140 16.4700 ;
      RECT 6.5800 15.3765 6.6060 16.4700 ;
      RECT 6.4720 15.3765 6.4980 16.4700 ;
      RECT 6.3640 15.3765 6.3900 16.4700 ;
      RECT 6.2560 15.3765 6.2820 16.4700 ;
      RECT 6.1480 15.3765 6.1740 16.4700 ;
      RECT 6.0400 15.3765 6.0660 16.4700 ;
      RECT 5.9320 15.3765 5.9580 16.4700 ;
      RECT 5.8240 15.3765 5.8500 16.4700 ;
      RECT 5.7160 15.3765 5.7420 16.4700 ;
      RECT 5.6080 15.3765 5.6340 16.4700 ;
      RECT 5.5000 15.3765 5.5260 16.4700 ;
      RECT 5.3920 15.3765 5.4180 16.4700 ;
      RECT 5.2840 15.3765 5.3100 16.4700 ;
      RECT 5.1760 15.3765 5.2020 16.4700 ;
      RECT 5.0680 15.3765 5.0940 16.4700 ;
      RECT 4.9600 15.3765 4.9860 16.4700 ;
      RECT 4.8520 15.3765 4.8780 16.4700 ;
      RECT 4.7440 15.3765 4.7700 16.4700 ;
      RECT 4.6360 15.3765 4.6620 16.4700 ;
      RECT 4.5280 15.3765 4.5540 16.4700 ;
      RECT 4.4200 15.3765 4.4460 16.4700 ;
      RECT 4.3120 15.3765 4.3380 16.4700 ;
      RECT 4.2040 15.3765 4.2300 16.4700 ;
      RECT 4.0960 15.3765 4.1220 16.4700 ;
      RECT 3.9880 15.3765 4.0140 16.4700 ;
      RECT 3.8800 15.3765 3.9060 16.4700 ;
      RECT 3.7720 15.3765 3.7980 16.4700 ;
      RECT 3.6640 15.3765 3.6900 16.4700 ;
      RECT 3.5560 15.3765 3.5820 16.4700 ;
      RECT 3.4480 15.3765 3.4740 16.4700 ;
      RECT 3.3400 15.3765 3.3660 16.4700 ;
      RECT 3.2320 15.3765 3.2580 16.4700 ;
      RECT 3.1240 15.3765 3.1500 16.4700 ;
      RECT 3.0160 15.3765 3.0420 16.4700 ;
      RECT 2.9080 15.3765 2.9340 16.4700 ;
      RECT 2.8000 15.3765 2.8260 16.4700 ;
      RECT 2.6920 15.3765 2.7180 16.4700 ;
      RECT 2.5840 15.3765 2.6100 16.4700 ;
      RECT 2.4760 15.3765 2.5020 16.4700 ;
      RECT 2.3680 15.3765 2.3940 16.4700 ;
      RECT 2.2600 15.3765 2.2860 16.4700 ;
      RECT 2.1520 15.3765 2.1780 16.4700 ;
      RECT 2.0440 15.3765 2.0700 16.4700 ;
      RECT 1.9360 15.3765 1.9620 16.4700 ;
      RECT 1.8280 15.3765 1.8540 16.4700 ;
      RECT 1.7200 15.3765 1.7460 16.4700 ;
      RECT 1.6120 15.3765 1.6380 16.4700 ;
      RECT 1.5040 15.3765 1.5300 16.4700 ;
      RECT 1.3960 15.3765 1.4220 16.4700 ;
      RECT 1.2880 15.3765 1.3140 16.4700 ;
      RECT 1.1800 15.3765 1.2060 16.4700 ;
      RECT 1.0720 15.3765 1.0980 16.4700 ;
      RECT 0.9640 15.3765 0.9900 16.4700 ;
      RECT 0.8560 15.3765 0.8820 16.4700 ;
      RECT 0.7480 15.3765 0.7740 16.4700 ;
      RECT 0.6400 15.3765 0.6660 16.4700 ;
      RECT 0.5320 15.3765 0.5580 16.4700 ;
      RECT 0.4240 15.3765 0.4500 16.4700 ;
      RECT 0.3160 15.3765 0.3420 16.4700 ;
      RECT 0.2080 15.3765 0.2340 16.4700 ;
      RECT 0.0050 15.3765 0.0900 16.4700 ;
      RECT 15.5530 16.4565 15.6810 17.5500 ;
      RECT 15.5390 17.1220 15.6810 17.4445 ;
      RECT 15.3190 16.8490 15.4530 17.5500 ;
      RECT 15.2960 17.1840 15.4530 17.4420 ;
      RECT 15.3190 16.4565 15.4170 17.5500 ;
      RECT 15.3190 16.5775 15.4310 16.8170 ;
      RECT 15.3190 16.4565 15.4530 16.5455 ;
      RECT 15.0940 16.9070 15.2280 17.5500 ;
      RECT 15.0940 16.4565 15.1920 17.5500 ;
      RECT 14.6770 16.4565 14.7600 17.5500 ;
      RECT 14.6770 16.5450 14.7740 17.4805 ;
      RECT 30.2680 16.4565 30.3530 17.5500 ;
      RECT 30.1240 16.4565 30.1500 17.5500 ;
      RECT 30.0160 16.4565 30.0420 17.5500 ;
      RECT 29.9080 16.4565 29.9340 17.5500 ;
      RECT 29.8000 16.4565 29.8260 17.5500 ;
      RECT 29.6920 16.4565 29.7180 17.5500 ;
      RECT 29.5840 16.4565 29.6100 17.5500 ;
      RECT 29.4760 16.4565 29.5020 17.5500 ;
      RECT 29.3680 16.4565 29.3940 17.5500 ;
      RECT 29.2600 16.4565 29.2860 17.5500 ;
      RECT 29.1520 16.4565 29.1780 17.5500 ;
      RECT 29.0440 16.4565 29.0700 17.5500 ;
      RECT 28.9360 16.4565 28.9620 17.5500 ;
      RECT 28.8280 16.4565 28.8540 17.5500 ;
      RECT 28.7200 16.4565 28.7460 17.5500 ;
      RECT 28.6120 16.4565 28.6380 17.5500 ;
      RECT 28.5040 16.4565 28.5300 17.5500 ;
      RECT 28.3960 16.4565 28.4220 17.5500 ;
      RECT 28.2880 16.4565 28.3140 17.5500 ;
      RECT 28.1800 16.4565 28.2060 17.5500 ;
      RECT 28.0720 16.4565 28.0980 17.5500 ;
      RECT 27.9640 16.4565 27.9900 17.5500 ;
      RECT 27.8560 16.4565 27.8820 17.5500 ;
      RECT 27.7480 16.4565 27.7740 17.5500 ;
      RECT 27.6400 16.4565 27.6660 17.5500 ;
      RECT 27.5320 16.4565 27.5580 17.5500 ;
      RECT 27.4240 16.4565 27.4500 17.5500 ;
      RECT 27.3160 16.4565 27.3420 17.5500 ;
      RECT 27.2080 16.4565 27.2340 17.5500 ;
      RECT 27.1000 16.4565 27.1260 17.5500 ;
      RECT 26.9920 16.4565 27.0180 17.5500 ;
      RECT 26.8840 16.4565 26.9100 17.5500 ;
      RECT 26.7760 16.4565 26.8020 17.5500 ;
      RECT 26.6680 16.4565 26.6940 17.5500 ;
      RECT 26.5600 16.4565 26.5860 17.5500 ;
      RECT 26.4520 16.4565 26.4780 17.5500 ;
      RECT 26.3440 16.4565 26.3700 17.5500 ;
      RECT 26.2360 16.4565 26.2620 17.5500 ;
      RECT 26.1280 16.4565 26.1540 17.5500 ;
      RECT 26.0200 16.4565 26.0460 17.5500 ;
      RECT 25.9120 16.4565 25.9380 17.5500 ;
      RECT 25.8040 16.4565 25.8300 17.5500 ;
      RECT 25.6960 16.4565 25.7220 17.5500 ;
      RECT 25.5880 16.4565 25.6140 17.5500 ;
      RECT 25.4800 16.4565 25.5060 17.5500 ;
      RECT 25.3720 16.4565 25.3980 17.5500 ;
      RECT 25.2640 16.4565 25.2900 17.5500 ;
      RECT 25.1560 16.4565 25.1820 17.5500 ;
      RECT 25.0480 16.4565 25.0740 17.5500 ;
      RECT 24.9400 16.4565 24.9660 17.5500 ;
      RECT 24.8320 16.4565 24.8580 17.5500 ;
      RECT 24.7240 16.4565 24.7500 17.5500 ;
      RECT 24.6160 16.4565 24.6420 17.5500 ;
      RECT 24.5080 16.4565 24.5340 17.5500 ;
      RECT 24.4000 16.4565 24.4260 17.5500 ;
      RECT 24.2920 16.4565 24.3180 17.5500 ;
      RECT 24.1840 16.4565 24.2100 17.5500 ;
      RECT 24.0760 16.4565 24.1020 17.5500 ;
      RECT 23.9680 16.4565 23.9940 17.5500 ;
      RECT 23.8600 16.4565 23.8860 17.5500 ;
      RECT 23.7520 16.4565 23.7780 17.5500 ;
      RECT 23.6440 16.4565 23.6700 17.5500 ;
      RECT 23.5360 16.4565 23.5620 17.5500 ;
      RECT 23.4280 16.4565 23.4540 17.5500 ;
      RECT 23.3200 16.4565 23.3460 17.5500 ;
      RECT 23.2120 16.4565 23.2380 17.5500 ;
      RECT 23.1040 16.4565 23.1300 17.5500 ;
      RECT 22.9960 16.4565 23.0220 17.5500 ;
      RECT 22.8880 16.4565 22.9140 17.5500 ;
      RECT 22.7800 16.4565 22.8060 17.5500 ;
      RECT 22.6720 16.4565 22.6980 17.5500 ;
      RECT 22.5640 16.4565 22.5900 17.5500 ;
      RECT 22.4560 16.4565 22.4820 17.5500 ;
      RECT 22.3480 16.4565 22.3740 17.5500 ;
      RECT 22.2400 16.4565 22.2660 17.5500 ;
      RECT 22.1320 16.4565 22.1580 17.5500 ;
      RECT 22.0240 16.4565 22.0500 17.5500 ;
      RECT 21.9160 16.4565 21.9420 17.5500 ;
      RECT 21.8080 16.4565 21.8340 17.5500 ;
      RECT 21.7000 16.4565 21.7260 17.5500 ;
      RECT 21.5920 16.4565 21.6180 17.5500 ;
      RECT 21.4840 16.4565 21.5100 17.5500 ;
      RECT 21.3760 16.4565 21.4020 17.5500 ;
      RECT 21.2680 16.4565 21.2940 17.5500 ;
      RECT 21.1600 16.4565 21.1860 17.5500 ;
      RECT 21.0520 16.4565 21.0780 17.5500 ;
      RECT 20.9440 16.4565 20.9700 17.5500 ;
      RECT 20.8360 16.4565 20.8620 17.5500 ;
      RECT 20.7280 16.4565 20.7540 17.5500 ;
      RECT 20.6200 16.4565 20.6460 17.5500 ;
      RECT 20.5120 16.4565 20.5380 17.5500 ;
      RECT 20.4040 16.4565 20.4300 17.5500 ;
      RECT 20.2960 16.4565 20.3220 17.5500 ;
      RECT 20.1880 16.4565 20.2140 17.5500 ;
      RECT 20.0800 16.4565 20.1060 17.5500 ;
      RECT 19.9720 16.4565 19.9980 17.5500 ;
      RECT 19.8640 16.4565 19.8900 17.5500 ;
      RECT 19.7560 16.4565 19.7820 17.5500 ;
      RECT 19.6480 16.4565 19.6740 17.5500 ;
      RECT 19.5400 16.4565 19.5660 17.5500 ;
      RECT 19.4320 16.4565 19.4580 17.5500 ;
      RECT 19.3240 16.4565 19.3500 17.5500 ;
      RECT 19.2160 16.4565 19.2420 17.5500 ;
      RECT 19.1080 16.4565 19.1340 17.5500 ;
      RECT 19.0000 16.4565 19.0260 17.5500 ;
      RECT 18.8920 16.4565 18.9180 17.5500 ;
      RECT 18.7840 16.4565 18.8100 17.5500 ;
      RECT 18.6760 16.4565 18.7020 17.5500 ;
      RECT 18.5680 16.4565 18.5940 17.5500 ;
      RECT 18.4600 16.4565 18.4860 17.5500 ;
      RECT 18.3520 16.4565 18.3780 17.5500 ;
      RECT 18.2440 16.4565 18.2700 17.5500 ;
      RECT 18.1360 16.4565 18.1620 17.5500 ;
      RECT 18.0280 16.4565 18.0540 17.5500 ;
      RECT 17.9200 16.4565 17.9460 17.5500 ;
      RECT 17.8120 16.4565 17.8380 17.5500 ;
      RECT 17.7040 16.4565 17.7300 17.5500 ;
      RECT 17.5960 16.4565 17.6220 17.5500 ;
      RECT 17.4880 16.4565 17.5140 17.5500 ;
      RECT 17.3800 16.4565 17.4060 17.5500 ;
      RECT 17.2720 16.4565 17.2980 17.5500 ;
      RECT 17.1640 16.4565 17.1900 17.5500 ;
      RECT 17.0560 16.4565 17.0820 17.5500 ;
      RECT 16.9480 16.4565 16.9740 17.5500 ;
      RECT 16.8400 16.4565 16.8660 17.5500 ;
      RECT 16.7320 16.4565 16.7580 17.5500 ;
      RECT 16.6240 16.4565 16.6500 17.5500 ;
      RECT 16.5160 16.4565 16.5420 17.5500 ;
      RECT 16.4080 16.4565 16.4340 17.5500 ;
      RECT 16.3000 16.4565 16.3260 17.5500 ;
      RECT 16.0870 16.4565 16.1640 17.5500 ;
      RECT 14.1940 16.4565 14.2710 17.5500 ;
      RECT 14.0320 16.4565 14.0580 17.5500 ;
      RECT 13.9240 16.4565 13.9500 17.5500 ;
      RECT 13.8160 16.4565 13.8420 17.5500 ;
      RECT 13.7080 16.4565 13.7340 17.5500 ;
      RECT 13.6000 16.4565 13.6260 17.5500 ;
      RECT 13.4920 16.4565 13.5180 17.5500 ;
      RECT 13.3840 16.4565 13.4100 17.5500 ;
      RECT 13.2760 16.4565 13.3020 17.5500 ;
      RECT 13.1680 16.4565 13.1940 17.5500 ;
      RECT 13.0600 16.4565 13.0860 17.5500 ;
      RECT 12.9520 16.4565 12.9780 17.5500 ;
      RECT 12.8440 16.4565 12.8700 17.5500 ;
      RECT 12.7360 16.4565 12.7620 17.5500 ;
      RECT 12.6280 16.4565 12.6540 17.5500 ;
      RECT 12.5200 16.4565 12.5460 17.5500 ;
      RECT 12.4120 16.4565 12.4380 17.5500 ;
      RECT 12.3040 16.4565 12.3300 17.5500 ;
      RECT 12.1960 16.4565 12.2220 17.5500 ;
      RECT 12.0880 16.4565 12.1140 17.5500 ;
      RECT 11.9800 16.4565 12.0060 17.5500 ;
      RECT 11.8720 16.4565 11.8980 17.5500 ;
      RECT 11.7640 16.4565 11.7900 17.5500 ;
      RECT 11.6560 16.4565 11.6820 17.5500 ;
      RECT 11.5480 16.4565 11.5740 17.5500 ;
      RECT 11.4400 16.4565 11.4660 17.5500 ;
      RECT 11.3320 16.4565 11.3580 17.5500 ;
      RECT 11.2240 16.4565 11.2500 17.5500 ;
      RECT 11.1160 16.4565 11.1420 17.5500 ;
      RECT 11.0080 16.4565 11.0340 17.5500 ;
      RECT 10.9000 16.4565 10.9260 17.5500 ;
      RECT 10.7920 16.4565 10.8180 17.5500 ;
      RECT 10.6840 16.4565 10.7100 17.5500 ;
      RECT 10.5760 16.4565 10.6020 17.5500 ;
      RECT 10.4680 16.4565 10.4940 17.5500 ;
      RECT 10.3600 16.4565 10.3860 17.5500 ;
      RECT 10.2520 16.4565 10.2780 17.5500 ;
      RECT 10.1440 16.4565 10.1700 17.5500 ;
      RECT 10.0360 16.4565 10.0620 17.5500 ;
      RECT 9.9280 16.4565 9.9540 17.5500 ;
      RECT 9.8200 16.4565 9.8460 17.5500 ;
      RECT 9.7120 16.4565 9.7380 17.5500 ;
      RECT 9.6040 16.4565 9.6300 17.5500 ;
      RECT 9.4960 16.4565 9.5220 17.5500 ;
      RECT 9.3880 16.4565 9.4140 17.5500 ;
      RECT 9.2800 16.4565 9.3060 17.5500 ;
      RECT 9.1720 16.4565 9.1980 17.5500 ;
      RECT 9.0640 16.4565 9.0900 17.5500 ;
      RECT 8.9560 16.4565 8.9820 17.5500 ;
      RECT 8.8480 16.4565 8.8740 17.5500 ;
      RECT 8.7400 16.4565 8.7660 17.5500 ;
      RECT 8.6320 16.4565 8.6580 17.5500 ;
      RECT 8.5240 16.4565 8.5500 17.5500 ;
      RECT 8.4160 16.4565 8.4420 17.5500 ;
      RECT 8.3080 16.4565 8.3340 17.5500 ;
      RECT 8.2000 16.4565 8.2260 17.5500 ;
      RECT 8.0920 16.4565 8.1180 17.5500 ;
      RECT 7.9840 16.4565 8.0100 17.5500 ;
      RECT 7.8760 16.4565 7.9020 17.5500 ;
      RECT 7.7680 16.4565 7.7940 17.5500 ;
      RECT 7.6600 16.4565 7.6860 17.5500 ;
      RECT 7.5520 16.4565 7.5780 17.5500 ;
      RECT 7.4440 16.4565 7.4700 17.5500 ;
      RECT 7.3360 16.4565 7.3620 17.5500 ;
      RECT 7.2280 16.4565 7.2540 17.5500 ;
      RECT 7.1200 16.4565 7.1460 17.5500 ;
      RECT 7.0120 16.4565 7.0380 17.5500 ;
      RECT 6.9040 16.4565 6.9300 17.5500 ;
      RECT 6.7960 16.4565 6.8220 17.5500 ;
      RECT 6.6880 16.4565 6.7140 17.5500 ;
      RECT 6.5800 16.4565 6.6060 17.5500 ;
      RECT 6.4720 16.4565 6.4980 17.5500 ;
      RECT 6.3640 16.4565 6.3900 17.5500 ;
      RECT 6.2560 16.4565 6.2820 17.5500 ;
      RECT 6.1480 16.4565 6.1740 17.5500 ;
      RECT 6.0400 16.4565 6.0660 17.5500 ;
      RECT 5.9320 16.4565 5.9580 17.5500 ;
      RECT 5.8240 16.4565 5.8500 17.5500 ;
      RECT 5.7160 16.4565 5.7420 17.5500 ;
      RECT 5.6080 16.4565 5.6340 17.5500 ;
      RECT 5.5000 16.4565 5.5260 17.5500 ;
      RECT 5.3920 16.4565 5.4180 17.5500 ;
      RECT 5.2840 16.4565 5.3100 17.5500 ;
      RECT 5.1760 16.4565 5.2020 17.5500 ;
      RECT 5.0680 16.4565 5.0940 17.5500 ;
      RECT 4.9600 16.4565 4.9860 17.5500 ;
      RECT 4.8520 16.4565 4.8780 17.5500 ;
      RECT 4.7440 16.4565 4.7700 17.5500 ;
      RECT 4.6360 16.4565 4.6620 17.5500 ;
      RECT 4.5280 16.4565 4.5540 17.5500 ;
      RECT 4.4200 16.4565 4.4460 17.5500 ;
      RECT 4.3120 16.4565 4.3380 17.5500 ;
      RECT 4.2040 16.4565 4.2300 17.5500 ;
      RECT 4.0960 16.4565 4.1220 17.5500 ;
      RECT 3.9880 16.4565 4.0140 17.5500 ;
      RECT 3.8800 16.4565 3.9060 17.5500 ;
      RECT 3.7720 16.4565 3.7980 17.5500 ;
      RECT 3.6640 16.4565 3.6900 17.5500 ;
      RECT 3.5560 16.4565 3.5820 17.5500 ;
      RECT 3.4480 16.4565 3.4740 17.5500 ;
      RECT 3.3400 16.4565 3.3660 17.5500 ;
      RECT 3.2320 16.4565 3.2580 17.5500 ;
      RECT 3.1240 16.4565 3.1500 17.5500 ;
      RECT 3.0160 16.4565 3.0420 17.5500 ;
      RECT 2.9080 16.4565 2.9340 17.5500 ;
      RECT 2.8000 16.4565 2.8260 17.5500 ;
      RECT 2.6920 16.4565 2.7180 17.5500 ;
      RECT 2.5840 16.4565 2.6100 17.5500 ;
      RECT 2.4760 16.4565 2.5020 17.5500 ;
      RECT 2.3680 16.4565 2.3940 17.5500 ;
      RECT 2.2600 16.4565 2.2860 17.5500 ;
      RECT 2.1520 16.4565 2.1780 17.5500 ;
      RECT 2.0440 16.4565 2.0700 17.5500 ;
      RECT 1.9360 16.4565 1.9620 17.5500 ;
      RECT 1.8280 16.4565 1.8540 17.5500 ;
      RECT 1.7200 16.4565 1.7460 17.5500 ;
      RECT 1.6120 16.4565 1.6380 17.5500 ;
      RECT 1.5040 16.4565 1.5300 17.5500 ;
      RECT 1.3960 16.4565 1.4220 17.5500 ;
      RECT 1.2880 16.4565 1.3140 17.5500 ;
      RECT 1.1800 16.4565 1.2060 17.5500 ;
      RECT 1.0720 16.4565 1.0980 17.5500 ;
      RECT 0.9640 16.4565 0.9900 17.5500 ;
      RECT 0.8560 16.4565 0.8820 17.5500 ;
      RECT 0.7480 16.4565 0.7740 17.5500 ;
      RECT 0.6400 16.4565 0.6660 17.5500 ;
      RECT 0.5320 16.4565 0.5580 17.5500 ;
      RECT 0.4240 16.4565 0.4500 17.5500 ;
      RECT 0.3160 16.4565 0.3420 17.5500 ;
      RECT 0.2080 16.4565 0.2340 17.5500 ;
      RECT 0.0050 16.4565 0.0900 17.5500 ;
      RECT 14.1350 25.7860 30.3480 26.2270 ;
      RECT 17.7530 17.5735 30.3480 26.2270 ;
      RECT 16.2950 19.0775 30.3480 26.2270 ;
      RECT 17.5370 18.8825 30.3480 26.2270 ;
      RECT 14.1350 25.4855 16.2130 26.2270 ;
      RECT 15.5570 18.9785 16.2130 26.2270 ;
      RECT 14.1350 19.1855 15.2590 26.2270 ;
      RECT 15.1970 17.5735 15.2590 26.2270 ;
      RECT 15.5430 24.2195 16.2130 25.3275 ;
      RECT 16.2810 21.3665 30.3480 24.9595 ;
      RECT 14.1350 24.4535 15.2730 24.7155 ;
      RECT 15.5430 21.6815 16.2130 24.0135 ;
      RECT 14.1350 22.0595 15.2730 23.3655 ;
      RECT 14.1350 19.3955 15.2730 22.0155 ;
      RECT 15.5430 18.8555 16.1590 20.6415 ;
      RECT 14.1890 19.1255 15.2730 19.3155 ;
      RECT 14.1890 18.3395 15.2590 26.2270 ;
      RECT 14.4050 18.2585 15.2590 26.2270 ;
      RECT 14.1890 18.8555 15.2730 19.0815 ;
      RECT 16.4570 18.8855 30.3480 26.2270 ;
      RECT 16.2950 17.5735 16.3750 26.2270 ;
      RECT 14.1350 18.2585 14.3230 19.0725 ;
      RECT 16.2950 17.5735 16.5910 18.9765 ;
      RECT 16.2950 18.6905 17.4550 18.9765 ;
      RECT 17.5370 17.5735 17.6710 26.2270 ;
      RECT 15.5570 18.6905 16.1590 26.2270 ;
      RECT 15.8810 17.5735 16.2130 18.8235 ;
      RECT 16.2950 18.6905 17.6710 18.7845 ;
      RECT 17.3210 17.5735 30.3480 18.7815 ;
      RECT 14.1350 18.7115 15.2730 18.7755 ;
      RECT 17.1050 18.3065 30.3480 18.7815 ;
      RECT 16.2950 18.3395 17.0230 18.9765 ;
      RECT 15.5570 18.3395 15.7990 26.2270 ;
      RECT 14.4050 18.3155 15.2730 18.5775 ;
      RECT 15.5930 17.5735 16.2130 18.4815 ;
      RECT 16.8890 17.5735 17.2390 18.4455 ;
      RECT 16.2950 18.2585 16.8070 18.9765 ;
      RECT 16.6730 17.5735 16.8070 26.2270 ;
      RECT 14.4050 17.5735 15.1150 26.2270 ;
      RECT 14.2250 17.5735 14.3230 26.2270 ;
      RECT 16.6730 17.5735 17.2390 18.2085 ;
      RECT 15.5570 17.5735 16.2130 18.2085 ;
      RECT 14.2250 17.5735 15.1150 18.2085 ;
      RECT 16.6730 17.5735 30.3480 18.2055 ;
      RECT 15.5430 18.0455 16.2130 18.1995 ;
      RECT 16.2950 17.5735 30.3480 17.9415 ;
      RECT 14.1350 17.5735 15.2590 17.9415 ;
      RECT 14.1350 17.5735 16.2130 17.7385 ;
      RECT 17.7570 17.3835 17.7750 26.2270 ;
      RECT 17.6490 17.3835 17.6670 26.2270 ;
      RECT 17.5410 17.3835 17.5590 26.2270 ;
      RECT 17.4330 17.3835 17.4510 26.2270 ;
      RECT 17.3250 17.3835 17.3430 26.2270 ;
      RECT 17.2170 17.3835 17.2350 26.2270 ;
      RECT 17.1090 17.3835 17.1270 26.2270 ;
      RECT 17.0010 17.3835 17.0190 26.2270 ;
      RECT 16.8930 17.3835 16.9110 26.2270 ;
      RECT 16.7850 17.3835 16.8030 26.2270 ;
      RECT 16.6770 17.3835 16.6950 26.2270 ;
      RECT 16.5690 17.3835 16.5870 26.2270 ;
      RECT 16.4610 17.3835 16.4790 26.2270 ;
      RECT 16.3530 17.3835 16.3710 26.2270 ;
      RECT 0.0000 18.8825 14.0170 26.2270 ;
      RECT 0.0000 21.6715 14.0310 21.7545 ;
      RECT 13.7570 17.5735 14.0530 21.3330 ;
      RECT 12.8930 18.5015 13.6750 26.2270 ;
      RECT 0.0000 17.5735 12.8110 26.2270 ;
      RECT 13.5410 17.5735 14.0530 18.7815 ;
      RECT 0.0000 18.3065 13.4590 18.7815 ;
      RECT 13.3250 17.5735 13.4590 26.2270 ;
      RECT 13.1090 18.2585 13.4590 26.2270 ;
      RECT 0.0000 17.5735 13.0270 18.7815 ;
      RECT 13.1090 17.5735 13.2430 26.2270 ;
      RECT 13.3250 17.5735 14.0530 18.2085 ;
      RECT 0.0000 17.5735 13.2430 18.2055 ;
      RECT 0.0000 17.5735 14.0530 17.9415 ;
      RECT 13.3290 17.5470 13.3470 26.2270 ;
      RECT 13.2210 17.5470 13.2390 26.2270 ;
        RECT 15.5530 25.6635 15.6810 26.7570 ;
        RECT 15.5390 26.3290 15.6810 26.6515 ;
        RECT 15.3190 26.0560 15.4530 26.7570 ;
        RECT 15.2960 26.3910 15.4530 26.6490 ;
        RECT 15.3190 25.6635 15.4170 26.7570 ;
        RECT 15.3190 25.7845 15.4310 26.0240 ;
        RECT 15.3190 25.6635 15.4530 25.7525 ;
        RECT 15.0940 26.1140 15.2280 26.7570 ;
        RECT 15.0940 25.6635 15.1920 26.7570 ;
        RECT 14.6770 25.6635 14.7600 26.7570 ;
        RECT 14.6770 25.7520 14.7740 26.6875 ;
        RECT 30.2680 25.6635 30.3530 26.7570 ;
        RECT 30.1240 25.6635 30.1500 26.7570 ;
        RECT 30.0160 25.6635 30.0420 26.7570 ;
        RECT 29.9080 25.6635 29.9340 26.7570 ;
        RECT 29.8000 25.6635 29.8260 26.7570 ;
        RECT 29.6920 25.6635 29.7180 26.7570 ;
        RECT 29.5840 25.6635 29.6100 26.7570 ;
        RECT 29.4760 25.6635 29.5020 26.7570 ;
        RECT 29.3680 25.6635 29.3940 26.7570 ;
        RECT 29.2600 25.6635 29.2860 26.7570 ;
        RECT 29.1520 25.6635 29.1780 26.7570 ;
        RECT 29.0440 25.6635 29.0700 26.7570 ;
        RECT 28.9360 25.6635 28.9620 26.7570 ;
        RECT 28.8280 25.6635 28.8540 26.7570 ;
        RECT 28.7200 25.6635 28.7460 26.7570 ;
        RECT 28.6120 25.6635 28.6380 26.7570 ;
        RECT 28.5040 25.6635 28.5300 26.7570 ;
        RECT 28.3960 25.6635 28.4220 26.7570 ;
        RECT 28.2880 25.6635 28.3140 26.7570 ;
        RECT 28.1800 25.6635 28.2060 26.7570 ;
        RECT 28.0720 25.6635 28.0980 26.7570 ;
        RECT 27.9640 25.6635 27.9900 26.7570 ;
        RECT 27.8560 25.6635 27.8820 26.7570 ;
        RECT 27.7480 25.6635 27.7740 26.7570 ;
        RECT 27.6400 25.6635 27.6660 26.7570 ;
        RECT 27.5320 25.6635 27.5580 26.7570 ;
        RECT 27.4240 25.6635 27.4500 26.7570 ;
        RECT 27.3160 25.6635 27.3420 26.7570 ;
        RECT 27.2080 25.6635 27.2340 26.7570 ;
        RECT 27.1000 25.6635 27.1260 26.7570 ;
        RECT 26.9920 25.6635 27.0180 26.7570 ;
        RECT 26.8840 25.6635 26.9100 26.7570 ;
        RECT 26.7760 25.6635 26.8020 26.7570 ;
        RECT 26.6680 25.6635 26.6940 26.7570 ;
        RECT 26.5600 25.6635 26.5860 26.7570 ;
        RECT 26.4520 25.6635 26.4780 26.7570 ;
        RECT 26.3440 25.6635 26.3700 26.7570 ;
        RECT 26.2360 25.6635 26.2620 26.7570 ;
        RECT 26.1280 25.6635 26.1540 26.7570 ;
        RECT 26.0200 25.6635 26.0460 26.7570 ;
        RECT 25.9120 25.6635 25.9380 26.7570 ;
        RECT 25.8040 25.6635 25.8300 26.7570 ;
        RECT 25.6960 25.6635 25.7220 26.7570 ;
        RECT 25.5880 25.6635 25.6140 26.7570 ;
        RECT 25.4800 25.6635 25.5060 26.7570 ;
        RECT 25.3720 25.6635 25.3980 26.7570 ;
        RECT 25.2640 25.6635 25.2900 26.7570 ;
        RECT 25.1560 25.6635 25.1820 26.7570 ;
        RECT 25.0480 25.6635 25.0740 26.7570 ;
        RECT 24.9400 25.6635 24.9660 26.7570 ;
        RECT 24.8320 25.6635 24.8580 26.7570 ;
        RECT 24.7240 25.6635 24.7500 26.7570 ;
        RECT 24.6160 25.6635 24.6420 26.7570 ;
        RECT 24.5080 25.6635 24.5340 26.7570 ;
        RECT 24.4000 25.6635 24.4260 26.7570 ;
        RECT 24.2920 25.6635 24.3180 26.7570 ;
        RECT 24.1840 25.6635 24.2100 26.7570 ;
        RECT 24.0760 25.6635 24.1020 26.7570 ;
        RECT 23.9680 25.6635 23.9940 26.7570 ;
        RECT 23.8600 25.6635 23.8860 26.7570 ;
        RECT 23.7520 25.6635 23.7780 26.7570 ;
        RECT 23.6440 25.6635 23.6700 26.7570 ;
        RECT 23.5360 25.6635 23.5620 26.7570 ;
        RECT 23.4280 25.6635 23.4540 26.7570 ;
        RECT 23.3200 25.6635 23.3460 26.7570 ;
        RECT 23.2120 25.6635 23.2380 26.7570 ;
        RECT 23.1040 25.6635 23.1300 26.7570 ;
        RECT 22.9960 25.6635 23.0220 26.7570 ;
        RECT 22.8880 25.6635 22.9140 26.7570 ;
        RECT 22.7800 25.6635 22.8060 26.7570 ;
        RECT 22.6720 25.6635 22.6980 26.7570 ;
        RECT 22.5640 25.6635 22.5900 26.7570 ;
        RECT 22.4560 25.6635 22.4820 26.7570 ;
        RECT 22.3480 25.6635 22.3740 26.7570 ;
        RECT 22.2400 25.6635 22.2660 26.7570 ;
        RECT 22.1320 25.6635 22.1580 26.7570 ;
        RECT 22.0240 25.6635 22.0500 26.7570 ;
        RECT 21.9160 25.6635 21.9420 26.7570 ;
        RECT 21.8080 25.6635 21.8340 26.7570 ;
        RECT 21.7000 25.6635 21.7260 26.7570 ;
        RECT 21.5920 25.6635 21.6180 26.7570 ;
        RECT 21.4840 25.6635 21.5100 26.7570 ;
        RECT 21.3760 25.6635 21.4020 26.7570 ;
        RECT 21.2680 25.6635 21.2940 26.7570 ;
        RECT 21.1600 25.6635 21.1860 26.7570 ;
        RECT 21.0520 25.6635 21.0780 26.7570 ;
        RECT 20.9440 25.6635 20.9700 26.7570 ;
        RECT 20.8360 25.6635 20.8620 26.7570 ;
        RECT 20.7280 25.6635 20.7540 26.7570 ;
        RECT 20.6200 25.6635 20.6460 26.7570 ;
        RECT 20.5120 25.6635 20.5380 26.7570 ;
        RECT 20.4040 25.6635 20.4300 26.7570 ;
        RECT 20.2960 25.6635 20.3220 26.7570 ;
        RECT 20.1880 25.6635 20.2140 26.7570 ;
        RECT 20.0800 25.6635 20.1060 26.7570 ;
        RECT 19.9720 25.6635 19.9980 26.7570 ;
        RECT 19.8640 25.6635 19.8900 26.7570 ;
        RECT 19.7560 25.6635 19.7820 26.7570 ;
        RECT 19.6480 25.6635 19.6740 26.7570 ;
        RECT 19.5400 25.6635 19.5660 26.7570 ;
        RECT 19.4320 25.6635 19.4580 26.7570 ;
        RECT 19.3240 25.6635 19.3500 26.7570 ;
        RECT 19.2160 25.6635 19.2420 26.7570 ;
        RECT 19.1080 25.6635 19.1340 26.7570 ;
        RECT 19.0000 25.6635 19.0260 26.7570 ;
        RECT 18.8920 25.6635 18.9180 26.7570 ;
        RECT 18.7840 25.6635 18.8100 26.7570 ;
        RECT 18.6760 25.6635 18.7020 26.7570 ;
        RECT 18.5680 25.6635 18.5940 26.7570 ;
        RECT 18.4600 25.6635 18.4860 26.7570 ;
        RECT 18.3520 25.6635 18.3780 26.7570 ;
        RECT 18.2440 25.6635 18.2700 26.7570 ;
        RECT 18.1360 25.6635 18.1620 26.7570 ;
        RECT 18.0280 25.6635 18.0540 26.7570 ;
        RECT 17.9200 25.6635 17.9460 26.7570 ;
        RECT 17.8120 25.6635 17.8380 26.7570 ;
        RECT 17.7040 25.6635 17.7300 26.7570 ;
        RECT 17.5960 25.6635 17.6220 26.7570 ;
        RECT 17.4880 25.6635 17.5140 26.7570 ;
        RECT 17.3800 25.6635 17.4060 26.7570 ;
        RECT 17.2720 25.6635 17.2980 26.7570 ;
        RECT 17.1640 25.6635 17.1900 26.7570 ;
        RECT 17.0560 25.6635 17.0820 26.7570 ;
        RECT 16.9480 25.6635 16.9740 26.7570 ;
        RECT 16.8400 25.6635 16.8660 26.7570 ;
        RECT 16.7320 25.6635 16.7580 26.7570 ;
        RECT 16.6240 25.6635 16.6500 26.7570 ;
        RECT 16.5160 25.6635 16.5420 26.7570 ;
        RECT 16.4080 25.6635 16.4340 26.7570 ;
        RECT 16.3000 25.6635 16.3260 26.7570 ;
        RECT 16.0870 25.6635 16.1640 26.7570 ;
        RECT 14.1940 25.6635 14.2710 26.7570 ;
        RECT 14.0320 25.6635 14.0580 26.7570 ;
        RECT 13.9240 25.6635 13.9500 26.7570 ;
        RECT 13.8160 25.6635 13.8420 26.7570 ;
        RECT 13.7080 25.6635 13.7340 26.7570 ;
        RECT 13.6000 25.6635 13.6260 26.7570 ;
        RECT 13.4920 25.6635 13.5180 26.7570 ;
        RECT 13.3840 25.6635 13.4100 26.7570 ;
        RECT 13.2760 25.6635 13.3020 26.7570 ;
        RECT 13.1680 25.6635 13.1940 26.7570 ;
        RECT 13.0600 25.6635 13.0860 26.7570 ;
        RECT 12.9520 25.6635 12.9780 26.7570 ;
        RECT 12.8440 25.6635 12.8700 26.7570 ;
        RECT 12.7360 25.6635 12.7620 26.7570 ;
        RECT 12.6280 25.6635 12.6540 26.7570 ;
        RECT 12.5200 25.6635 12.5460 26.7570 ;
        RECT 12.4120 25.6635 12.4380 26.7570 ;
        RECT 12.3040 25.6635 12.3300 26.7570 ;
        RECT 12.1960 25.6635 12.2220 26.7570 ;
        RECT 12.0880 25.6635 12.1140 26.7570 ;
        RECT 11.9800 25.6635 12.0060 26.7570 ;
        RECT 11.8720 25.6635 11.8980 26.7570 ;
        RECT 11.7640 25.6635 11.7900 26.7570 ;
        RECT 11.6560 25.6635 11.6820 26.7570 ;
        RECT 11.5480 25.6635 11.5740 26.7570 ;
        RECT 11.4400 25.6635 11.4660 26.7570 ;
        RECT 11.3320 25.6635 11.3580 26.7570 ;
        RECT 11.2240 25.6635 11.2500 26.7570 ;
        RECT 11.1160 25.6635 11.1420 26.7570 ;
        RECT 11.0080 25.6635 11.0340 26.7570 ;
        RECT 10.9000 25.6635 10.9260 26.7570 ;
        RECT 10.7920 25.6635 10.8180 26.7570 ;
        RECT 10.6840 25.6635 10.7100 26.7570 ;
        RECT 10.5760 25.6635 10.6020 26.7570 ;
        RECT 10.4680 25.6635 10.4940 26.7570 ;
        RECT 10.3600 25.6635 10.3860 26.7570 ;
        RECT 10.2520 25.6635 10.2780 26.7570 ;
        RECT 10.1440 25.6635 10.1700 26.7570 ;
        RECT 10.0360 25.6635 10.0620 26.7570 ;
        RECT 9.9280 25.6635 9.9540 26.7570 ;
        RECT 9.8200 25.6635 9.8460 26.7570 ;
        RECT 9.7120 25.6635 9.7380 26.7570 ;
        RECT 9.6040 25.6635 9.6300 26.7570 ;
        RECT 9.4960 25.6635 9.5220 26.7570 ;
        RECT 9.3880 25.6635 9.4140 26.7570 ;
        RECT 9.2800 25.6635 9.3060 26.7570 ;
        RECT 9.1720 25.6635 9.1980 26.7570 ;
        RECT 9.0640 25.6635 9.0900 26.7570 ;
        RECT 8.9560 25.6635 8.9820 26.7570 ;
        RECT 8.8480 25.6635 8.8740 26.7570 ;
        RECT 8.7400 25.6635 8.7660 26.7570 ;
        RECT 8.6320 25.6635 8.6580 26.7570 ;
        RECT 8.5240 25.6635 8.5500 26.7570 ;
        RECT 8.4160 25.6635 8.4420 26.7570 ;
        RECT 8.3080 25.6635 8.3340 26.7570 ;
        RECT 8.2000 25.6635 8.2260 26.7570 ;
        RECT 8.0920 25.6635 8.1180 26.7570 ;
        RECT 7.9840 25.6635 8.0100 26.7570 ;
        RECT 7.8760 25.6635 7.9020 26.7570 ;
        RECT 7.7680 25.6635 7.7940 26.7570 ;
        RECT 7.6600 25.6635 7.6860 26.7570 ;
        RECT 7.5520 25.6635 7.5780 26.7570 ;
        RECT 7.4440 25.6635 7.4700 26.7570 ;
        RECT 7.3360 25.6635 7.3620 26.7570 ;
        RECT 7.2280 25.6635 7.2540 26.7570 ;
        RECT 7.1200 25.6635 7.1460 26.7570 ;
        RECT 7.0120 25.6635 7.0380 26.7570 ;
        RECT 6.9040 25.6635 6.9300 26.7570 ;
        RECT 6.7960 25.6635 6.8220 26.7570 ;
        RECT 6.6880 25.6635 6.7140 26.7570 ;
        RECT 6.5800 25.6635 6.6060 26.7570 ;
        RECT 6.4720 25.6635 6.4980 26.7570 ;
        RECT 6.3640 25.6635 6.3900 26.7570 ;
        RECT 6.2560 25.6635 6.2820 26.7570 ;
        RECT 6.1480 25.6635 6.1740 26.7570 ;
        RECT 6.0400 25.6635 6.0660 26.7570 ;
        RECT 5.9320 25.6635 5.9580 26.7570 ;
        RECT 5.8240 25.6635 5.8500 26.7570 ;
        RECT 5.7160 25.6635 5.7420 26.7570 ;
        RECT 5.6080 25.6635 5.6340 26.7570 ;
        RECT 5.5000 25.6635 5.5260 26.7570 ;
        RECT 5.3920 25.6635 5.4180 26.7570 ;
        RECT 5.2840 25.6635 5.3100 26.7570 ;
        RECT 5.1760 25.6635 5.2020 26.7570 ;
        RECT 5.0680 25.6635 5.0940 26.7570 ;
        RECT 4.9600 25.6635 4.9860 26.7570 ;
        RECT 4.8520 25.6635 4.8780 26.7570 ;
        RECT 4.7440 25.6635 4.7700 26.7570 ;
        RECT 4.6360 25.6635 4.6620 26.7570 ;
        RECT 4.5280 25.6635 4.5540 26.7570 ;
        RECT 4.4200 25.6635 4.4460 26.7570 ;
        RECT 4.3120 25.6635 4.3380 26.7570 ;
        RECT 4.2040 25.6635 4.2300 26.7570 ;
        RECT 4.0960 25.6635 4.1220 26.7570 ;
        RECT 3.9880 25.6635 4.0140 26.7570 ;
        RECT 3.8800 25.6635 3.9060 26.7570 ;
        RECT 3.7720 25.6635 3.7980 26.7570 ;
        RECT 3.6640 25.6635 3.6900 26.7570 ;
        RECT 3.5560 25.6635 3.5820 26.7570 ;
        RECT 3.4480 25.6635 3.4740 26.7570 ;
        RECT 3.3400 25.6635 3.3660 26.7570 ;
        RECT 3.2320 25.6635 3.2580 26.7570 ;
        RECT 3.1240 25.6635 3.1500 26.7570 ;
        RECT 3.0160 25.6635 3.0420 26.7570 ;
        RECT 2.9080 25.6635 2.9340 26.7570 ;
        RECT 2.8000 25.6635 2.8260 26.7570 ;
        RECT 2.6920 25.6635 2.7180 26.7570 ;
        RECT 2.5840 25.6635 2.6100 26.7570 ;
        RECT 2.4760 25.6635 2.5020 26.7570 ;
        RECT 2.3680 25.6635 2.3940 26.7570 ;
        RECT 2.2600 25.6635 2.2860 26.7570 ;
        RECT 2.1520 25.6635 2.1780 26.7570 ;
        RECT 2.0440 25.6635 2.0700 26.7570 ;
        RECT 1.9360 25.6635 1.9620 26.7570 ;
        RECT 1.8280 25.6635 1.8540 26.7570 ;
        RECT 1.7200 25.6635 1.7460 26.7570 ;
        RECT 1.6120 25.6635 1.6380 26.7570 ;
        RECT 1.5040 25.6635 1.5300 26.7570 ;
        RECT 1.3960 25.6635 1.4220 26.7570 ;
        RECT 1.2880 25.6635 1.3140 26.7570 ;
        RECT 1.1800 25.6635 1.2060 26.7570 ;
        RECT 1.0720 25.6635 1.0980 26.7570 ;
        RECT 0.9640 25.6635 0.9900 26.7570 ;
        RECT 0.8560 25.6635 0.8820 26.7570 ;
        RECT 0.7480 25.6635 0.7740 26.7570 ;
        RECT 0.6400 25.6635 0.6660 26.7570 ;
        RECT 0.5320 25.6635 0.5580 26.7570 ;
        RECT 0.4240 25.6635 0.4500 26.7570 ;
        RECT 0.3160 25.6635 0.3420 26.7570 ;
        RECT 0.2080 25.6635 0.2340 26.7570 ;
        RECT 0.0050 25.6635 0.0900 26.7570 ;
        RECT 15.5530 26.7435 15.6810 27.8370 ;
        RECT 15.5390 27.4090 15.6810 27.7315 ;
        RECT 15.3190 27.1360 15.4530 27.8370 ;
        RECT 15.2960 27.4710 15.4530 27.7290 ;
        RECT 15.3190 26.7435 15.4170 27.8370 ;
        RECT 15.3190 26.8645 15.4310 27.1040 ;
        RECT 15.3190 26.7435 15.4530 26.8325 ;
        RECT 15.0940 27.1940 15.2280 27.8370 ;
        RECT 15.0940 26.7435 15.1920 27.8370 ;
        RECT 14.6770 26.7435 14.7600 27.8370 ;
        RECT 14.6770 26.8320 14.7740 27.7675 ;
        RECT 30.2680 26.7435 30.3530 27.8370 ;
        RECT 30.1240 26.7435 30.1500 27.8370 ;
        RECT 30.0160 26.7435 30.0420 27.8370 ;
        RECT 29.9080 26.7435 29.9340 27.8370 ;
        RECT 29.8000 26.7435 29.8260 27.8370 ;
        RECT 29.6920 26.7435 29.7180 27.8370 ;
        RECT 29.5840 26.7435 29.6100 27.8370 ;
        RECT 29.4760 26.7435 29.5020 27.8370 ;
        RECT 29.3680 26.7435 29.3940 27.8370 ;
        RECT 29.2600 26.7435 29.2860 27.8370 ;
        RECT 29.1520 26.7435 29.1780 27.8370 ;
        RECT 29.0440 26.7435 29.0700 27.8370 ;
        RECT 28.9360 26.7435 28.9620 27.8370 ;
        RECT 28.8280 26.7435 28.8540 27.8370 ;
        RECT 28.7200 26.7435 28.7460 27.8370 ;
        RECT 28.6120 26.7435 28.6380 27.8370 ;
        RECT 28.5040 26.7435 28.5300 27.8370 ;
        RECT 28.3960 26.7435 28.4220 27.8370 ;
        RECT 28.2880 26.7435 28.3140 27.8370 ;
        RECT 28.1800 26.7435 28.2060 27.8370 ;
        RECT 28.0720 26.7435 28.0980 27.8370 ;
        RECT 27.9640 26.7435 27.9900 27.8370 ;
        RECT 27.8560 26.7435 27.8820 27.8370 ;
        RECT 27.7480 26.7435 27.7740 27.8370 ;
        RECT 27.6400 26.7435 27.6660 27.8370 ;
        RECT 27.5320 26.7435 27.5580 27.8370 ;
        RECT 27.4240 26.7435 27.4500 27.8370 ;
        RECT 27.3160 26.7435 27.3420 27.8370 ;
        RECT 27.2080 26.7435 27.2340 27.8370 ;
        RECT 27.1000 26.7435 27.1260 27.8370 ;
        RECT 26.9920 26.7435 27.0180 27.8370 ;
        RECT 26.8840 26.7435 26.9100 27.8370 ;
        RECT 26.7760 26.7435 26.8020 27.8370 ;
        RECT 26.6680 26.7435 26.6940 27.8370 ;
        RECT 26.5600 26.7435 26.5860 27.8370 ;
        RECT 26.4520 26.7435 26.4780 27.8370 ;
        RECT 26.3440 26.7435 26.3700 27.8370 ;
        RECT 26.2360 26.7435 26.2620 27.8370 ;
        RECT 26.1280 26.7435 26.1540 27.8370 ;
        RECT 26.0200 26.7435 26.0460 27.8370 ;
        RECT 25.9120 26.7435 25.9380 27.8370 ;
        RECT 25.8040 26.7435 25.8300 27.8370 ;
        RECT 25.6960 26.7435 25.7220 27.8370 ;
        RECT 25.5880 26.7435 25.6140 27.8370 ;
        RECT 25.4800 26.7435 25.5060 27.8370 ;
        RECT 25.3720 26.7435 25.3980 27.8370 ;
        RECT 25.2640 26.7435 25.2900 27.8370 ;
        RECT 25.1560 26.7435 25.1820 27.8370 ;
        RECT 25.0480 26.7435 25.0740 27.8370 ;
        RECT 24.9400 26.7435 24.9660 27.8370 ;
        RECT 24.8320 26.7435 24.8580 27.8370 ;
        RECT 24.7240 26.7435 24.7500 27.8370 ;
        RECT 24.6160 26.7435 24.6420 27.8370 ;
        RECT 24.5080 26.7435 24.5340 27.8370 ;
        RECT 24.4000 26.7435 24.4260 27.8370 ;
        RECT 24.2920 26.7435 24.3180 27.8370 ;
        RECT 24.1840 26.7435 24.2100 27.8370 ;
        RECT 24.0760 26.7435 24.1020 27.8370 ;
        RECT 23.9680 26.7435 23.9940 27.8370 ;
        RECT 23.8600 26.7435 23.8860 27.8370 ;
        RECT 23.7520 26.7435 23.7780 27.8370 ;
        RECT 23.6440 26.7435 23.6700 27.8370 ;
        RECT 23.5360 26.7435 23.5620 27.8370 ;
        RECT 23.4280 26.7435 23.4540 27.8370 ;
        RECT 23.3200 26.7435 23.3460 27.8370 ;
        RECT 23.2120 26.7435 23.2380 27.8370 ;
        RECT 23.1040 26.7435 23.1300 27.8370 ;
        RECT 22.9960 26.7435 23.0220 27.8370 ;
        RECT 22.8880 26.7435 22.9140 27.8370 ;
        RECT 22.7800 26.7435 22.8060 27.8370 ;
        RECT 22.6720 26.7435 22.6980 27.8370 ;
        RECT 22.5640 26.7435 22.5900 27.8370 ;
        RECT 22.4560 26.7435 22.4820 27.8370 ;
        RECT 22.3480 26.7435 22.3740 27.8370 ;
        RECT 22.2400 26.7435 22.2660 27.8370 ;
        RECT 22.1320 26.7435 22.1580 27.8370 ;
        RECT 22.0240 26.7435 22.0500 27.8370 ;
        RECT 21.9160 26.7435 21.9420 27.8370 ;
        RECT 21.8080 26.7435 21.8340 27.8370 ;
        RECT 21.7000 26.7435 21.7260 27.8370 ;
        RECT 21.5920 26.7435 21.6180 27.8370 ;
        RECT 21.4840 26.7435 21.5100 27.8370 ;
        RECT 21.3760 26.7435 21.4020 27.8370 ;
        RECT 21.2680 26.7435 21.2940 27.8370 ;
        RECT 21.1600 26.7435 21.1860 27.8370 ;
        RECT 21.0520 26.7435 21.0780 27.8370 ;
        RECT 20.9440 26.7435 20.9700 27.8370 ;
        RECT 20.8360 26.7435 20.8620 27.8370 ;
        RECT 20.7280 26.7435 20.7540 27.8370 ;
        RECT 20.6200 26.7435 20.6460 27.8370 ;
        RECT 20.5120 26.7435 20.5380 27.8370 ;
        RECT 20.4040 26.7435 20.4300 27.8370 ;
        RECT 20.2960 26.7435 20.3220 27.8370 ;
        RECT 20.1880 26.7435 20.2140 27.8370 ;
        RECT 20.0800 26.7435 20.1060 27.8370 ;
        RECT 19.9720 26.7435 19.9980 27.8370 ;
        RECT 19.8640 26.7435 19.8900 27.8370 ;
        RECT 19.7560 26.7435 19.7820 27.8370 ;
        RECT 19.6480 26.7435 19.6740 27.8370 ;
        RECT 19.5400 26.7435 19.5660 27.8370 ;
        RECT 19.4320 26.7435 19.4580 27.8370 ;
        RECT 19.3240 26.7435 19.3500 27.8370 ;
        RECT 19.2160 26.7435 19.2420 27.8370 ;
        RECT 19.1080 26.7435 19.1340 27.8370 ;
        RECT 19.0000 26.7435 19.0260 27.8370 ;
        RECT 18.8920 26.7435 18.9180 27.8370 ;
        RECT 18.7840 26.7435 18.8100 27.8370 ;
        RECT 18.6760 26.7435 18.7020 27.8370 ;
        RECT 18.5680 26.7435 18.5940 27.8370 ;
        RECT 18.4600 26.7435 18.4860 27.8370 ;
        RECT 18.3520 26.7435 18.3780 27.8370 ;
        RECT 18.2440 26.7435 18.2700 27.8370 ;
        RECT 18.1360 26.7435 18.1620 27.8370 ;
        RECT 18.0280 26.7435 18.0540 27.8370 ;
        RECT 17.9200 26.7435 17.9460 27.8370 ;
        RECT 17.8120 26.7435 17.8380 27.8370 ;
        RECT 17.7040 26.7435 17.7300 27.8370 ;
        RECT 17.5960 26.7435 17.6220 27.8370 ;
        RECT 17.4880 26.7435 17.5140 27.8370 ;
        RECT 17.3800 26.7435 17.4060 27.8370 ;
        RECT 17.2720 26.7435 17.2980 27.8370 ;
        RECT 17.1640 26.7435 17.1900 27.8370 ;
        RECT 17.0560 26.7435 17.0820 27.8370 ;
        RECT 16.9480 26.7435 16.9740 27.8370 ;
        RECT 16.8400 26.7435 16.8660 27.8370 ;
        RECT 16.7320 26.7435 16.7580 27.8370 ;
        RECT 16.6240 26.7435 16.6500 27.8370 ;
        RECT 16.5160 26.7435 16.5420 27.8370 ;
        RECT 16.4080 26.7435 16.4340 27.8370 ;
        RECT 16.3000 26.7435 16.3260 27.8370 ;
        RECT 16.0870 26.7435 16.1640 27.8370 ;
        RECT 14.1940 26.7435 14.2710 27.8370 ;
        RECT 14.0320 26.7435 14.0580 27.8370 ;
        RECT 13.9240 26.7435 13.9500 27.8370 ;
        RECT 13.8160 26.7435 13.8420 27.8370 ;
        RECT 13.7080 26.7435 13.7340 27.8370 ;
        RECT 13.6000 26.7435 13.6260 27.8370 ;
        RECT 13.4920 26.7435 13.5180 27.8370 ;
        RECT 13.3840 26.7435 13.4100 27.8370 ;
        RECT 13.2760 26.7435 13.3020 27.8370 ;
        RECT 13.1680 26.7435 13.1940 27.8370 ;
        RECT 13.0600 26.7435 13.0860 27.8370 ;
        RECT 12.9520 26.7435 12.9780 27.8370 ;
        RECT 12.8440 26.7435 12.8700 27.8370 ;
        RECT 12.7360 26.7435 12.7620 27.8370 ;
        RECT 12.6280 26.7435 12.6540 27.8370 ;
        RECT 12.5200 26.7435 12.5460 27.8370 ;
        RECT 12.4120 26.7435 12.4380 27.8370 ;
        RECT 12.3040 26.7435 12.3300 27.8370 ;
        RECT 12.1960 26.7435 12.2220 27.8370 ;
        RECT 12.0880 26.7435 12.1140 27.8370 ;
        RECT 11.9800 26.7435 12.0060 27.8370 ;
        RECT 11.8720 26.7435 11.8980 27.8370 ;
        RECT 11.7640 26.7435 11.7900 27.8370 ;
        RECT 11.6560 26.7435 11.6820 27.8370 ;
        RECT 11.5480 26.7435 11.5740 27.8370 ;
        RECT 11.4400 26.7435 11.4660 27.8370 ;
        RECT 11.3320 26.7435 11.3580 27.8370 ;
        RECT 11.2240 26.7435 11.2500 27.8370 ;
        RECT 11.1160 26.7435 11.1420 27.8370 ;
        RECT 11.0080 26.7435 11.0340 27.8370 ;
        RECT 10.9000 26.7435 10.9260 27.8370 ;
        RECT 10.7920 26.7435 10.8180 27.8370 ;
        RECT 10.6840 26.7435 10.7100 27.8370 ;
        RECT 10.5760 26.7435 10.6020 27.8370 ;
        RECT 10.4680 26.7435 10.4940 27.8370 ;
        RECT 10.3600 26.7435 10.3860 27.8370 ;
        RECT 10.2520 26.7435 10.2780 27.8370 ;
        RECT 10.1440 26.7435 10.1700 27.8370 ;
        RECT 10.0360 26.7435 10.0620 27.8370 ;
        RECT 9.9280 26.7435 9.9540 27.8370 ;
        RECT 9.8200 26.7435 9.8460 27.8370 ;
        RECT 9.7120 26.7435 9.7380 27.8370 ;
        RECT 9.6040 26.7435 9.6300 27.8370 ;
        RECT 9.4960 26.7435 9.5220 27.8370 ;
        RECT 9.3880 26.7435 9.4140 27.8370 ;
        RECT 9.2800 26.7435 9.3060 27.8370 ;
        RECT 9.1720 26.7435 9.1980 27.8370 ;
        RECT 9.0640 26.7435 9.0900 27.8370 ;
        RECT 8.9560 26.7435 8.9820 27.8370 ;
        RECT 8.8480 26.7435 8.8740 27.8370 ;
        RECT 8.7400 26.7435 8.7660 27.8370 ;
        RECT 8.6320 26.7435 8.6580 27.8370 ;
        RECT 8.5240 26.7435 8.5500 27.8370 ;
        RECT 8.4160 26.7435 8.4420 27.8370 ;
        RECT 8.3080 26.7435 8.3340 27.8370 ;
        RECT 8.2000 26.7435 8.2260 27.8370 ;
        RECT 8.0920 26.7435 8.1180 27.8370 ;
        RECT 7.9840 26.7435 8.0100 27.8370 ;
        RECT 7.8760 26.7435 7.9020 27.8370 ;
        RECT 7.7680 26.7435 7.7940 27.8370 ;
        RECT 7.6600 26.7435 7.6860 27.8370 ;
        RECT 7.5520 26.7435 7.5780 27.8370 ;
        RECT 7.4440 26.7435 7.4700 27.8370 ;
        RECT 7.3360 26.7435 7.3620 27.8370 ;
        RECT 7.2280 26.7435 7.2540 27.8370 ;
        RECT 7.1200 26.7435 7.1460 27.8370 ;
        RECT 7.0120 26.7435 7.0380 27.8370 ;
        RECT 6.9040 26.7435 6.9300 27.8370 ;
        RECT 6.7960 26.7435 6.8220 27.8370 ;
        RECT 6.6880 26.7435 6.7140 27.8370 ;
        RECT 6.5800 26.7435 6.6060 27.8370 ;
        RECT 6.4720 26.7435 6.4980 27.8370 ;
        RECT 6.3640 26.7435 6.3900 27.8370 ;
        RECT 6.2560 26.7435 6.2820 27.8370 ;
        RECT 6.1480 26.7435 6.1740 27.8370 ;
        RECT 6.0400 26.7435 6.0660 27.8370 ;
        RECT 5.9320 26.7435 5.9580 27.8370 ;
        RECT 5.8240 26.7435 5.8500 27.8370 ;
        RECT 5.7160 26.7435 5.7420 27.8370 ;
        RECT 5.6080 26.7435 5.6340 27.8370 ;
        RECT 5.5000 26.7435 5.5260 27.8370 ;
        RECT 5.3920 26.7435 5.4180 27.8370 ;
        RECT 5.2840 26.7435 5.3100 27.8370 ;
        RECT 5.1760 26.7435 5.2020 27.8370 ;
        RECT 5.0680 26.7435 5.0940 27.8370 ;
        RECT 4.9600 26.7435 4.9860 27.8370 ;
        RECT 4.8520 26.7435 4.8780 27.8370 ;
        RECT 4.7440 26.7435 4.7700 27.8370 ;
        RECT 4.6360 26.7435 4.6620 27.8370 ;
        RECT 4.5280 26.7435 4.5540 27.8370 ;
        RECT 4.4200 26.7435 4.4460 27.8370 ;
        RECT 4.3120 26.7435 4.3380 27.8370 ;
        RECT 4.2040 26.7435 4.2300 27.8370 ;
        RECT 4.0960 26.7435 4.1220 27.8370 ;
        RECT 3.9880 26.7435 4.0140 27.8370 ;
        RECT 3.8800 26.7435 3.9060 27.8370 ;
        RECT 3.7720 26.7435 3.7980 27.8370 ;
        RECT 3.6640 26.7435 3.6900 27.8370 ;
        RECT 3.5560 26.7435 3.5820 27.8370 ;
        RECT 3.4480 26.7435 3.4740 27.8370 ;
        RECT 3.3400 26.7435 3.3660 27.8370 ;
        RECT 3.2320 26.7435 3.2580 27.8370 ;
        RECT 3.1240 26.7435 3.1500 27.8370 ;
        RECT 3.0160 26.7435 3.0420 27.8370 ;
        RECT 2.9080 26.7435 2.9340 27.8370 ;
        RECT 2.8000 26.7435 2.8260 27.8370 ;
        RECT 2.6920 26.7435 2.7180 27.8370 ;
        RECT 2.5840 26.7435 2.6100 27.8370 ;
        RECT 2.4760 26.7435 2.5020 27.8370 ;
        RECT 2.3680 26.7435 2.3940 27.8370 ;
        RECT 2.2600 26.7435 2.2860 27.8370 ;
        RECT 2.1520 26.7435 2.1780 27.8370 ;
        RECT 2.0440 26.7435 2.0700 27.8370 ;
        RECT 1.9360 26.7435 1.9620 27.8370 ;
        RECT 1.8280 26.7435 1.8540 27.8370 ;
        RECT 1.7200 26.7435 1.7460 27.8370 ;
        RECT 1.6120 26.7435 1.6380 27.8370 ;
        RECT 1.5040 26.7435 1.5300 27.8370 ;
        RECT 1.3960 26.7435 1.4220 27.8370 ;
        RECT 1.2880 26.7435 1.3140 27.8370 ;
        RECT 1.1800 26.7435 1.2060 27.8370 ;
        RECT 1.0720 26.7435 1.0980 27.8370 ;
        RECT 0.9640 26.7435 0.9900 27.8370 ;
        RECT 0.8560 26.7435 0.8820 27.8370 ;
        RECT 0.7480 26.7435 0.7740 27.8370 ;
        RECT 0.6400 26.7435 0.6660 27.8370 ;
        RECT 0.5320 26.7435 0.5580 27.8370 ;
        RECT 0.4240 26.7435 0.4500 27.8370 ;
        RECT 0.3160 26.7435 0.3420 27.8370 ;
        RECT 0.2080 26.7435 0.2340 27.8370 ;
        RECT 0.0050 26.7435 0.0900 27.8370 ;
        RECT 15.5530 27.8235 15.6810 28.9170 ;
        RECT 15.5390 28.4890 15.6810 28.8115 ;
        RECT 15.3190 28.2160 15.4530 28.9170 ;
        RECT 15.2960 28.5510 15.4530 28.8090 ;
        RECT 15.3190 27.8235 15.4170 28.9170 ;
        RECT 15.3190 27.9445 15.4310 28.1840 ;
        RECT 15.3190 27.8235 15.4530 27.9125 ;
        RECT 15.0940 28.2740 15.2280 28.9170 ;
        RECT 15.0940 27.8235 15.1920 28.9170 ;
        RECT 14.6770 27.8235 14.7600 28.9170 ;
        RECT 14.6770 27.9120 14.7740 28.8475 ;
        RECT 30.2680 27.8235 30.3530 28.9170 ;
        RECT 30.1240 27.8235 30.1500 28.9170 ;
        RECT 30.0160 27.8235 30.0420 28.9170 ;
        RECT 29.9080 27.8235 29.9340 28.9170 ;
        RECT 29.8000 27.8235 29.8260 28.9170 ;
        RECT 29.6920 27.8235 29.7180 28.9170 ;
        RECT 29.5840 27.8235 29.6100 28.9170 ;
        RECT 29.4760 27.8235 29.5020 28.9170 ;
        RECT 29.3680 27.8235 29.3940 28.9170 ;
        RECT 29.2600 27.8235 29.2860 28.9170 ;
        RECT 29.1520 27.8235 29.1780 28.9170 ;
        RECT 29.0440 27.8235 29.0700 28.9170 ;
        RECT 28.9360 27.8235 28.9620 28.9170 ;
        RECT 28.8280 27.8235 28.8540 28.9170 ;
        RECT 28.7200 27.8235 28.7460 28.9170 ;
        RECT 28.6120 27.8235 28.6380 28.9170 ;
        RECT 28.5040 27.8235 28.5300 28.9170 ;
        RECT 28.3960 27.8235 28.4220 28.9170 ;
        RECT 28.2880 27.8235 28.3140 28.9170 ;
        RECT 28.1800 27.8235 28.2060 28.9170 ;
        RECT 28.0720 27.8235 28.0980 28.9170 ;
        RECT 27.9640 27.8235 27.9900 28.9170 ;
        RECT 27.8560 27.8235 27.8820 28.9170 ;
        RECT 27.7480 27.8235 27.7740 28.9170 ;
        RECT 27.6400 27.8235 27.6660 28.9170 ;
        RECT 27.5320 27.8235 27.5580 28.9170 ;
        RECT 27.4240 27.8235 27.4500 28.9170 ;
        RECT 27.3160 27.8235 27.3420 28.9170 ;
        RECT 27.2080 27.8235 27.2340 28.9170 ;
        RECT 27.1000 27.8235 27.1260 28.9170 ;
        RECT 26.9920 27.8235 27.0180 28.9170 ;
        RECT 26.8840 27.8235 26.9100 28.9170 ;
        RECT 26.7760 27.8235 26.8020 28.9170 ;
        RECT 26.6680 27.8235 26.6940 28.9170 ;
        RECT 26.5600 27.8235 26.5860 28.9170 ;
        RECT 26.4520 27.8235 26.4780 28.9170 ;
        RECT 26.3440 27.8235 26.3700 28.9170 ;
        RECT 26.2360 27.8235 26.2620 28.9170 ;
        RECT 26.1280 27.8235 26.1540 28.9170 ;
        RECT 26.0200 27.8235 26.0460 28.9170 ;
        RECT 25.9120 27.8235 25.9380 28.9170 ;
        RECT 25.8040 27.8235 25.8300 28.9170 ;
        RECT 25.6960 27.8235 25.7220 28.9170 ;
        RECT 25.5880 27.8235 25.6140 28.9170 ;
        RECT 25.4800 27.8235 25.5060 28.9170 ;
        RECT 25.3720 27.8235 25.3980 28.9170 ;
        RECT 25.2640 27.8235 25.2900 28.9170 ;
        RECT 25.1560 27.8235 25.1820 28.9170 ;
        RECT 25.0480 27.8235 25.0740 28.9170 ;
        RECT 24.9400 27.8235 24.9660 28.9170 ;
        RECT 24.8320 27.8235 24.8580 28.9170 ;
        RECT 24.7240 27.8235 24.7500 28.9170 ;
        RECT 24.6160 27.8235 24.6420 28.9170 ;
        RECT 24.5080 27.8235 24.5340 28.9170 ;
        RECT 24.4000 27.8235 24.4260 28.9170 ;
        RECT 24.2920 27.8235 24.3180 28.9170 ;
        RECT 24.1840 27.8235 24.2100 28.9170 ;
        RECT 24.0760 27.8235 24.1020 28.9170 ;
        RECT 23.9680 27.8235 23.9940 28.9170 ;
        RECT 23.8600 27.8235 23.8860 28.9170 ;
        RECT 23.7520 27.8235 23.7780 28.9170 ;
        RECT 23.6440 27.8235 23.6700 28.9170 ;
        RECT 23.5360 27.8235 23.5620 28.9170 ;
        RECT 23.4280 27.8235 23.4540 28.9170 ;
        RECT 23.3200 27.8235 23.3460 28.9170 ;
        RECT 23.2120 27.8235 23.2380 28.9170 ;
        RECT 23.1040 27.8235 23.1300 28.9170 ;
        RECT 22.9960 27.8235 23.0220 28.9170 ;
        RECT 22.8880 27.8235 22.9140 28.9170 ;
        RECT 22.7800 27.8235 22.8060 28.9170 ;
        RECT 22.6720 27.8235 22.6980 28.9170 ;
        RECT 22.5640 27.8235 22.5900 28.9170 ;
        RECT 22.4560 27.8235 22.4820 28.9170 ;
        RECT 22.3480 27.8235 22.3740 28.9170 ;
        RECT 22.2400 27.8235 22.2660 28.9170 ;
        RECT 22.1320 27.8235 22.1580 28.9170 ;
        RECT 22.0240 27.8235 22.0500 28.9170 ;
        RECT 21.9160 27.8235 21.9420 28.9170 ;
        RECT 21.8080 27.8235 21.8340 28.9170 ;
        RECT 21.7000 27.8235 21.7260 28.9170 ;
        RECT 21.5920 27.8235 21.6180 28.9170 ;
        RECT 21.4840 27.8235 21.5100 28.9170 ;
        RECT 21.3760 27.8235 21.4020 28.9170 ;
        RECT 21.2680 27.8235 21.2940 28.9170 ;
        RECT 21.1600 27.8235 21.1860 28.9170 ;
        RECT 21.0520 27.8235 21.0780 28.9170 ;
        RECT 20.9440 27.8235 20.9700 28.9170 ;
        RECT 20.8360 27.8235 20.8620 28.9170 ;
        RECT 20.7280 27.8235 20.7540 28.9170 ;
        RECT 20.6200 27.8235 20.6460 28.9170 ;
        RECT 20.5120 27.8235 20.5380 28.9170 ;
        RECT 20.4040 27.8235 20.4300 28.9170 ;
        RECT 20.2960 27.8235 20.3220 28.9170 ;
        RECT 20.1880 27.8235 20.2140 28.9170 ;
        RECT 20.0800 27.8235 20.1060 28.9170 ;
        RECT 19.9720 27.8235 19.9980 28.9170 ;
        RECT 19.8640 27.8235 19.8900 28.9170 ;
        RECT 19.7560 27.8235 19.7820 28.9170 ;
        RECT 19.6480 27.8235 19.6740 28.9170 ;
        RECT 19.5400 27.8235 19.5660 28.9170 ;
        RECT 19.4320 27.8235 19.4580 28.9170 ;
        RECT 19.3240 27.8235 19.3500 28.9170 ;
        RECT 19.2160 27.8235 19.2420 28.9170 ;
        RECT 19.1080 27.8235 19.1340 28.9170 ;
        RECT 19.0000 27.8235 19.0260 28.9170 ;
        RECT 18.8920 27.8235 18.9180 28.9170 ;
        RECT 18.7840 27.8235 18.8100 28.9170 ;
        RECT 18.6760 27.8235 18.7020 28.9170 ;
        RECT 18.5680 27.8235 18.5940 28.9170 ;
        RECT 18.4600 27.8235 18.4860 28.9170 ;
        RECT 18.3520 27.8235 18.3780 28.9170 ;
        RECT 18.2440 27.8235 18.2700 28.9170 ;
        RECT 18.1360 27.8235 18.1620 28.9170 ;
        RECT 18.0280 27.8235 18.0540 28.9170 ;
        RECT 17.9200 27.8235 17.9460 28.9170 ;
        RECT 17.8120 27.8235 17.8380 28.9170 ;
        RECT 17.7040 27.8235 17.7300 28.9170 ;
        RECT 17.5960 27.8235 17.6220 28.9170 ;
        RECT 17.4880 27.8235 17.5140 28.9170 ;
        RECT 17.3800 27.8235 17.4060 28.9170 ;
        RECT 17.2720 27.8235 17.2980 28.9170 ;
        RECT 17.1640 27.8235 17.1900 28.9170 ;
        RECT 17.0560 27.8235 17.0820 28.9170 ;
        RECT 16.9480 27.8235 16.9740 28.9170 ;
        RECT 16.8400 27.8235 16.8660 28.9170 ;
        RECT 16.7320 27.8235 16.7580 28.9170 ;
        RECT 16.6240 27.8235 16.6500 28.9170 ;
        RECT 16.5160 27.8235 16.5420 28.9170 ;
        RECT 16.4080 27.8235 16.4340 28.9170 ;
        RECT 16.3000 27.8235 16.3260 28.9170 ;
        RECT 16.0870 27.8235 16.1640 28.9170 ;
        RECT 14.1940 27.8235 14.2710 28.9170 ;
        RECT 14.0320 27.8235 14.0580 28.9170 ;
        RECT 13.9240 27.8235 13.9500 28.9170 ;
        RECT 13.8160 27.8235 13.8420 28.9170 ;
        RECT 13.7080 27.8235 13.7340 28.9170 ;
        RECT 13.6000 27.8235 13.6260 28.9170 ;
        RECT 13.4920 27.8235 13.5180 28.9170 ;
        RECT 13.3840 27.8235 13.4100 28.9170 ;
        RECT 13.2760 27.8235 13.3020 28.9170 ;
        RECT 13.1680 27.8235 13.1940 28.9170 ;
        RECT 13.0600 27.8235 13.0860 28.9170 ;
        RECT 12.9520 27.8235 12.9780 28.9170 ;
        RECT 12.8440 27.8235 12.8700 28.9170 ;
        RECT 12.7360 27.8235 12.7620 28.9170 ;
        RECT 12.6280 27.8235 12.6540 28.9170 ;
        RECT 12.5200 27.8235 12.5460 28.9170 ;
        RECT 12.4120 27.8235 12.4380 28.9170 ;
        RECT 12.3040 27.8235 12.3300 28.9170 ;
        RECT 12.1960 27.8235 12.2220 28.9170 ;
        RECT 12.0880 27.8235 12.1140 28.9170 ;
        RECT 11.9800 27.8235 12.0060 28.9170 ;
        RECT 11.8720 27.8235 11.8980 28.9170 ;
        RECT 11.7640 27.8235 11.7900 28.9170 ;
        RECT 11.6560 27.8235 11.6820 28.9170 ;
        RECT 11.5480 27.8235 11.5740 28.9170 ;
        RECT 11.4400 27.8235 11.4660 28.9170 ;
        RECT 11.3320 27.8235 11.3580 28.9170 ;
        RECT 11.2240 27.8235 11.2500 28.9170 ;
        RECT 11.1160 27.8235 11.1420 28.9170 ;
        RECT 11.0080 27.8235 11.0340 28.9170 ;
        RECT 10.9000 27.8235 10.9260 28.9170 ;
        RECT 10.7920 27.8235 10.8180 28.9170 ;
        RECT 10.6840 27.8235 10.7100 28.9170 ;
        RECT 10.5760 27.8235 10.6020 28.9170 ;
        RECT 10.4680 27.8235 10.4940 28.9170 ;
        RECT 10.3600 27.8235 10.3860 28.9170 ;
        RECT 10.2520 27.8235 10.2780 28.9170 ;
        RECT 10.1440 27.8235 10.1700 28.9170 ;
        RECT 10.0360 27.8235 10.0620 28.9170 ;
        RECT 9.9280 27.8235 9.9540 28.9170 ;
        RECT 9.8200 27.8235 9.8460 28.9170 ;
        RECT 9.7120 27.8235 9.7380 28.9170 ;
        RECT 9.6040 27.8235 9.6300 28.9170 ;
        RECT 9.4960 27.8235 9.5220 28.9170 ;
        RECT 9.3880 27.8235 9.4140 28.9170 ;
        RECT 9.2800 27.8235 9.3060 28.9170 ;
        RECT 9.1720 27.8235 9.1980 28.9170 ;
        RECT 9.0640 27.8235 9.0900 28.9170 ;
        RECT 8.9560 27.8235 8.9820 28.9170 ;
        RECT 8.8480 27.8235 8.8740 28.9170 ;
        RECT 8.7400 27.8235 8.7660 28.9170 ;
        RECT 8.6320 27.8235 8.6580 28.9170 ;
        RECT 8.5240 27.8235 8.5500 28.9170 ;
        RECT 8.4160 27.8235 8.4420 28.9170 ;
        RECT 8.3080 27.8235 8.3340 28.9170 ;
        RECT 8.2000 27.8235 8.2260 28.9170 ;
        RECT 8.0920 27.8235 8.1180 28.9170 ;
        RECT 7.9840 27.8235 8.0100 28.9170 ;
        RECT 7.8760 27.8235 7.9020 28.9170 ;
        RECT 7.7680 27.8235 7.7940 28.9170 ;
        RECT 7.6600 27.8235 7.6860 28.9170 ;
        RECT 7.5520 27.8235 7.5780 28.9170 ;
        RECT 7.4440 27.8235 7.4700 28.9170 ;
        RECT 7.3360 27.8235 7.3620 28.9170 ;
        RECT 7.2280 27.8235 7.2540 28.9170 ;
        RECT 7.1200 27.8235 7.1460 28.9170 ;
        RECT 7.0120 27.8235 7.0380 28.9170 ;
        RECT 6.9040 27.8235 6.9300 28.9170 ;
        RECT 6.7960 27.8235 6.8220 28.9170 ;
        RECT 6.6880 27.8235 6.7140 28.9170 ;
        RECT 6.5800 27.8235 6.6060 28.9170 ;
        RECT 6.4720 27.8235 6.4980 28.9170 ;
        RECT 6.3640 27.8235 6.3900 28.9170 ;
        RECT 6.2560 27.8235 6.2820 28.9170 ;
        RECT 6.1480 27.8235 6.1740 28.9170 ;
        RECT 6.0400 27.8235 6.0660 28.9170 ;
        RECT 5.9320 27.8235 5.9580 28.9170 ;
        RECT 5.8240 27.8235 5.8500 28.9170 ;
        RECT 5.7160 27.8235 5.7420 28.9170 ;
        RECT 5.6080 27.8235 5.6340 28.9170 ;
        RECT 5.5000 27.8235 5.5260 28.9170 ;
        RECT 5.3920 27.8235 5.4180 28.9170 ;
        RECT 5.2840 27.8235 5.3100 28.9170 ;
        RECT 5.1760 27.8235 5.2020 28.9170 ;
        RECT 5.0680 27.8235 5.0940 28.9170 ;
        RECT 4.9600 27.8235 4.9860 28.9170 ;
        RECT 4.8520 27.8235 4.8780 28.9170 ;
        RECT 4.7440 27.8235 4.7700 28.9170 ;
        RECT 4.6360 27.8235 4.6620 28.9170 ;
        RECT 4.5280 27.8235 4.5540 28.9170 ;
        RECT 4.4200 27.8235 4.4460 28.9170 ;
        RECT 4.3120 27.8235 4.3380 28.9170 ;
        RECT 4.2040 27.8235 4.2300 28.9170 ;
        RECT 4.0960 27.8235 4.1220 28.9170 ;
        RECT 3.9880 27.8235 4.0140 28.9170 ;
        RECT 3.8800 27.8235 3.9060 28.9170 ;
        RECT 3.7720 27.8235 3.7980 28.9170 ;
        RECT 3.6640 27.8235 3.6900 28.9170 ;
        RECT 3.5560 27.8235 3.5820 28.9170 ;
        RECT 3.4480 27.8235 3.4740 28.9170 ;
        RECT 3.3400 27.8235 3.3660 28.9170 ;
        RECT 3.2320 27.8235 3.2580 28.9170 ;
        RECT 3.1240 27.8235 3.1500 28.9170 ;
        RECT 3.0160 27.8235 3.0420 28.9170 ;
        RECT 2.9080 27.8235 2.9340 28.9170 ;
        RECT 2.8000 27.8235 2.8260 28.9170 ;
        RECT 2.6920 27.8235 2.7180 28.9170 ;
        RECT 2.5840 27.8235 2.6100 28.9170 ;
        RECT 2.4760 27.8235 2.5020 28.9170 ;
        RECT 2.3680 27.8235 2.3940 28.9170 ;
        RECT 2.2600 27.8235 2.2860 28.9170 ;
        RECT 2.1520 27.8235 2.1780 28.9170 ;
        RECT 2.0440 27.8235 2.0700 28.9170 ;
        RECT 1.9360 27.8235 1.9620 28.9170 ;
        RECT 1.8280 27.8235 1.8540 28.9170 ;
        RECT 1.7200 27.8235 1.7460 28.9170 ;
        RECT 1.6120 27.8235 1.6380 28.9170 ;
        RECT 1.5040 27.8235 1.5300 28.9170 ;
        RECT 1.3960 27.8235 1.4220 28.9170 ;
        RECT 1.2880 27.8235 1.3140 28.9170 ;
        RECT 1.1800 27.8235 1.2060 28.9170 ;
        RECT 1.0720 27.8235 1.0980 28.9170 ;
        RECT 0.9640 27.8235 0.9900 28.9170 ;
        RECT 0.8560 27.8235 0.8820 28.9170 ;
        RECT 0.7480 27.8235 0.7740 28.9170 ;
        RECT 0.6400 27.8235 0.6660 28.9170 ;
        RECT 0.5320 27.8235 0.5580 28.9170 ;
        RECT 0.4240 27.8235 0.4500 28.9170 ;
        RECT 0.3160 27.8235 0.3420 28.9170 ;
        RECT 0.2080 27.8235 0.2340 28.9170 ;
        RECT 0.0050 27.8235 0.0900 28.9170 ;
        RECT 15.5530 28.9035 15.6810 29.9970 ;
        RECT 15.5390 29.5690 15.6810 29.8915 ;
        RECT 15.3190 29.2960 15.4530 29.9970 ;
        RECT 15.2960 29.6310 15.4530 29.8890 ;
        RECT 15.3190 28.9035 15.4170 29.9970 ;
        RECT 15.3190 29.0245 15.4310 29.2640 ;
        RECT 15.3190 28.9035 15.4530 28.9925 ;
        RECT 15.0940 29.3540 15.2280 29.9970 ;
        RECT 15.0940 28.9035 15.1920 29.9970 ;
        RECT 14.6770 28.9035 14.7600 29.9970 ;
        RECT 14.6770 28.9920 14.7740 29.9275 ;
        RECT 30.2680 28.9035 30.3530 29.9970 ;
        RECT 30.1240 28.9035 30.1500 29.9970 ;
        RECT 30.0160 28.9035 30.0420 29.9970 ;
        RECT 29.9080 28.9035 29.9340 29.9970 ;
        RECT 29.8000 28.9035 29.8260 29.9970 ;
        RECT 29.6920 28.9035 29.7180 29.9970 ;
        RECT 29.5840 28.9035 29.6100 29.9970 ;
        RECT 29.4760 28.9035 29.5020 29.9970 ;
        RECT 29.3680 28.9035 29.3940 29.9970 ;
        RECT 29.2600 28.9035 29.2860 29.9970 ;
        RECT 29.1520 28.9035 29.1780 29.9970 ;
        RECT 29.0440 28.9035 29.0700 29.9970 ;
        RECT 28.9360 28.9035 28.9620 29.9970 ;
        RECT 28.8280 28.9035 28.8540 29.9970 ;
        RECT 28.7200 28.9035 28.7460 29.9970 ;
        RECT 28.6120 28.9035 28.6380 29.9970 ;
        RECT 28.5040 28.9035 28.5300 29.9970 ;
        RECT 28.3960 28.9035 28.4220 29.9970 ;
        RECT 28.2880 28.9035 28.3140 29.9970 ;
        RECT 28.1800 28.9035 28.2060 29.9970 ;
        RECT 28.0720 28.9035 28.0980 29.9970 ;
        RECT 27.9640 28.9035 27.9900 29.9970 ;
        RECT 27.8560 28.9035 27.8820 29.9970 ;
        RECT 27.7480 28.9035 27.7740 29.9970 ;
        RECT 27.6400 28.9035 27.6660 29.9970 ;
        RECT 27.5320 28.9035 27.5580 29.9970 ;
        RECT 27.4240 28.9035 27.4500 29.9970 ;
        RECT 27.3160 28.9035 27.3420 29.9970 ;
        RECT 27.2080 28.9035 27.2340 29.9970 ;
        RECT 27.1000 28.9035 27.1260 29.9970 ;
        RECT 26.9920 28.9035 27.0180 29.9970 ;
        RECT 26.8840 28.9035 26.9100 29.9970 ;
        RECT 26.7760 28.9035 26.8020 29.9970 ;
        RECT 26.6680 28.9035 26.6940 29.9970 ;
        RECT 26.5600 28.9035 26.5860 29.9970 ;
        RECT 26.4520 28.9035 26.4780 29.9970 ;
        RECT 26.3440 28.9035 26.3700 29.9970 ;
        RECT 26.2360 28.9035 26.2620 29.9970 ;
        RECT 26.1280 28.9035 26.1540 29.9970 ;
        RECT 26.0200 28.9035 26.0460 29.9970 ;
        RECT 25.9120 28.9035 25.9380 29.9970 ;
        RECT 25.8040 28.9035 25.8300 29.9970 ;
        RECT 25.6960 28.9035 25.7220 29.9970 ;
        RECT 25.5880 28.9035 25.6140 29.9970 ;
        RECT 25.4800 28.9035 25.5060 29.9970 ;
        RECT 25.3720 28.9035 25.3980 29.9970 ;
        RECT 25.2640 28.9035 25.2900 29.9970 ;
        RECT 25.1560 28.9035 25.1820 29.9970 ;
        RECT 25.0480 28.9035 25.0740 29.9970 ;
        RECT 24.9400 28.9035 24.9660 29.9970 ;
        RECT 24.8320 28.9035 24.8580 29.9970 ;
        RECT 24.7240 28.9035 24.7500 29.9970 ;
        RECT 24.6160 28.9035 24.6420 29.9970 ;
        RECT 24.5080 28.9035 24.5340 29.9970 ;
        RECT 24.4000 28.9035 24.4260 29.9970 ;
        RECT 24.2920 28.9035 24.3180 29.9970 ;
        RECT 24.1840 28.9035 24.2100 29.9970 ;
        RECT 24.0760 28.9035 24.1020 29.9970 ;
        RECT 23.9680 28.9035 23.9940 29.9970 ;
        RECT 23.8600 28.9035 23.8860 29.9970 ;
        RECT 23.7520 28.9035 23.7780 29.9970 ;
        RECT 23.6440 28.9035 23.6700 29.9970 ;
        RECT 23.5360 28.9035 23.5620 29.9970 ;
        RECT 23.4280 28.9035 23.4540 29.9970 ;
        RECT 23.3200 28.9035 23.3460 29.9970 ;
        RECT 23.2120 28.9035 23.2380 29.9970 ;
        RECT 23.1040 28.9035 23.1300 29.9970 ;
        RECT 22.9960 28.9035 23.0220 29.9970 ;
        RECT 22.8880 28.9035 22.9140 29.9970 ;
        RECT 22.7800 28.9035 22.8060 29.9970 ;
        RECT 22.6720 28.9035 22.6980 29.9970 ;
        RECT 22.5640 28.9035 22.5900 29.9970 ;
        RECT 22.4560 28.9035 22.4820 29.9970 ;
        RECT 22.3480 28.9035 22.3740 29.9970 ;
        RECT 22.2400 28.9035 22.2660 29.9970 ;
        RECT 22.1320 28.9035 22.1580 29.9970 ;
        RECT 22.0240 28.9035 22.0500 29.9970 ;
        RECT 21.9160 28.9035 21.9420 29.9970 ;
        RECT 21.8080 28.9035 21.8340 29.9970 ;
        RECT 21.7000 28.9035 21.7260 29.9970 ;
        RECT 21.5920 28.9035 21.6180 29.9970 ;
        RECT 21.4840 28.9035 21.5100 29.9970 ;
        RECT 21.3760 28.9035 21.4020 29.9970 ;
        RECT 21.2680 28.9035 21.2940 29.9970 ;
        RECT 21.1600 28.9035 21.1860 29.9970 ;
        RECT 21.0520 28.9035 21.0780 29.9970 ;
        RECT 20.9440 28.9035 20.9700 29.9970 ;
        RECT 20.8360 28.9035 20.8620 29.9970 ;
        RECT 20.7280 28.9035 20.7540 29.9970 ;
        RECT 20.6200 28.9035 20.6460 29.9970 ;
        RECT 20.5120 28.9035 20.5380 29.9970 ;
        RECT 20.4040 28.9035 20.4300 29.9970 ;
        RECT 20.2960 28.9035 20.3220 29.9970 ;
        RECT 20.1880 28.9035 20.2140 29.9970 ;
        RECT 20.0800 28.9035 20.1060 29.9970 ;
        RECT 19.9720 28.9035 19.9980 29.9970 ;
        RECT 19.8640 28.9035 19.8900 29.9970 ;
        RECT 19.7560 28.9035 19.7820 29.9970 ;
        RECT 19.6480 28.9035 19.6740 29.9970 ;
        RECT 19.5400 28.9035 19.5660 29.9970 ;
        RECT 19.4320 28.9035 19.4580 29.9970 ;
        RECT 19.3240 28.9035 19.3500 29.9970 ;
        RECT 19.2160 28.9035 19.2420 29.9970 ;
        RECT 19.1080 28.9035 19.1340 29.9970 ;
        RECT 19.0000 28.9035 19.0260 29.9970 ;
        RECT 18.8920 28.9035 18.9180 29.9970 ;
        RECT 18.7840 28.9035 18.8100 29.9970 ;
        RECT 18.6760 28.9035 18.7020 29.9970 ;
        RECT 18.5680 28.9035 18.5940 29.9970 ;
        RECT 18.4600 28.9035 18.4860 29.9970 ;
        RECT 18.3520 28.9035 18.3780 29.9970 ;
        RECT 18.2440 28.9035 18.2700 29.9970 ;
        RECT 18.1360 28.9035 18.1620 29.9970 ;
        RECT 18.0280 28.9035 18.0540 29.9970 ;
        RECT 17.9200 28.9035 17.9460 29.9970 ;
        RECT 17.8120 28.9035 17.8380 29.9970 ;
        RECT 17.7040 28.9035 17.7300 29.9970 ;
        RECT 17.5960 28.9035 17.6220 29.9970 ;
        RECT 17.4880 28.9035 17.5140 29.9970 ;
        RECT 17.3800 28.9035 17.4060 29.9970 ;
        RECT 17.2720 28.9035 17.2980 29.9970 ;
        RECT 17.1640 28.9035 17.1900 29.9970 ;
        RECT 17.0560 28.9035 17.0820 29.9970 ;
        RECT 16.9480 28.9035 16.9740 29.9970 ;
        RECT 16.8400 28.9035 16.8660 29.9970 ;
        RECT 16.7320 28.9035 16.7580 29.9970 ;
        RECT 16.6240 28.9035 16.6500 29.9970 ;
        RECT 16.5160 28.9035 16.5420 29.9970 ;
        RECT 16.4080 28.9035 16.4340 29.9970 ;
        RECT 16.3000 28.9035 16.3260 29.9970 ;
        RECT 16.0870 28.9035 16.1640 29.9970 ;
        RECT 14.1940 28.9035 14.2710 29.9970 ;
        RECT 14.0320 28.9035 14.0580 29.9970 ;
        RECT 13.9240 28.9035 13.9500 29.9970 ;
        RECT 13.8160 28.9035 13.8420 29.9970 ;
        RECT 13.7080 28.9035 13.7340 29.9970 ;
        RECT 13.6000 28.9035 13.6260 29.9970 ;
        RECT 13.4920 28.9035 13.5180 29.9970 ;
        RECT 13.3840 28.9035 13.4100 29.9970 ;
        RECT 13.2760 28.9035 13.3020 29.9970 ;
        RECT 13.1680 28.9035 13.1940 29.9970 ;
        RECT 13.0600 28.9035 13.0860 29.9970 ;
        RECT 12.9520 28.9035 12.9780 29.9970 ;
        RECT 12.8440 28.9035 12.8700 29.9970 ;
        RECT 12.7360 28.9035 12.7620 29.9970 ;
        RECT 12.6280 28.9035 12.6540 29.9970 ;
        RECT 12.5200 28.9035 12.5460 29.9970 ;
        RECT 12.4120 28.9035 12.4380 29.9970 ;
        RECT 12.3040 28.9035 12.3300 29.9970 ;
        RECT 12.1960 28.9035 12.2220 29.9970 ;
        RECT 12.0880 28.9035 12.1140 29.9970 ;
        RECT 11.9800 28.9035 12.0060 29.9970 ;
        RECT 11.8720 28.9035 11.8980 29.9970 ;
        RECT 11.7640 28.9035 11.7900 29.9970 ;
        RECT 11.6560 28.9035 11.6820 29.9970 ;
        RECT 11.5480 28.9035 11.5740 29.9970 ;
        RECT 11.4400 28.9035 11.4660 29.9970 ;
        RECT 11.3320 28.9035 11.3580 29.9970 ;
        RECT 11.2240 28.9035 11.2500 29.9970 ;
        RECT 11.1160 28.9035 11.1420 29.9970 ;
        RECT 11.0080 28.9035 11.0340 29.9970 ;
        RECT 10.9000 28.9035 10.9260 29.9970 ;
        RECT 10.7920 28.9035 10.8180 29.9970 ;
        RECT 10.6840 28.9035 10.7100 29.9970 ;
        RECT 10.5760 28.9035 10.6020 29.9970 ;
        RECT 10.4680 28.9035 10.4940 29.9970 ;
        RECT 10.3600 28.9035 10.3860 29.9970 ;
        RECT 10.2520 28.9035 10.2780 29.9970 ;
        RECT 10.1440 28.9035 10.1700 29.9970 ;
        RECT 10.0360 28.9035 10.0620 29.9970 ;
        RECT 9.9280 28.9035 9.9540 29.9970 ;
        RECT 9.8200 28.9035 9.8460 29.9970 ;
        RECT 9.7120 28.9035 9.7380 29.9970 ;
        RECT 9.6040 28.9035 9.6300 29.9970 ;
        RECT 9.4960 28.9035 9.5220 29.9970 ;
        RECT 9.3880 28.9035 9.4140 29.9970 ;
        RECT 9.2800 28.9035 9.3060 29.9970 ;
        RECT 9.1720 28.9035 9.1980 29.9970 ;
        RECT 9.0640 28.9035 9.0900 29.9970 ;
        RECT 8.9560 28.9035 8.9820 29.9970 ;
        RECT 8.8480 28.9035 8.8740 29.9970 ;
        RECT 8.7400 28.9035 8.7660 29.9970 ;
        RECT 8.6320 28.9035 8.6580 29.9970 ;
        RECT 8.5240 28.9035 8.5500 29.9970 ;
        RECT 8.4160 28.9035 8.4420 29.9970 ;
        RECT 8.3080 28.9035 8.3340 29.9970 ;
        RECT 8.2000 28.9035 8.2260 29.9970 ;
        RECT 8.0920 28.9035 8.1180 29.9970 ;
        RECT 7.9840 28.9035 8.0100 29.9970 ;
        RECT 7.8760 28.9035 7.9020 29.9970 ;
        RECT 7.7680 28.9035 7.7940 29.9970 ;
        RECT 7.6600 28.9035 7.6860 29.9970 ;
        RECT 7.5520 28.9035 7.5780 29.9970 ;
        RECT 7.4440 28.9035 7.4700 29.9970 ;
        RECT 7.3360 28.9035 7.3620 29.9970 ;
        RECT 7.2280 28.9035 7.2540 29.9970 ;
        RECT 7.1200 28.9035 7.1460 29.9970 ;
        RECT 7.0120 28.9035 7.0380 29.9970 ;
        RECT 6.9040 28.9035 6.9300 29.9970 ;
        RECT 6.7960 28.9035 6.8220 29.9970 ;
        RECT 6.6880 28.9035 6.7140 29.9970 ;
        RECT 6.5800 28.9035 6.6060 29.9970 ;
        RECT 6.4720 28.9035 6.4980 29.9970 ;
        RECT 6.3640 28.9035 6.3900 29.9970 ;
        RECT 6.2560 28.9035 6.2820 29.9970 ;
        RECT 6.1480 28.9035 6.1740 29.9970 ;
        RECT 6.0400 28.9035 6.0660 29.9970 ;
        RECT 5.9320 28.9035 5.9580 29.9970 ;
        RECT 5.8240 28.9035 5.8500 29.9970 ;
        RECT 5.7160 28.9035 5.7420 29.9970 ;
        RECT 5.6080 28.9035 5.6340 29.9970 ;
        RECT 5.5000 28.9035 5.5260 29.9970 ;
        RECT 5.3920 28.9035 5.4180 29.9970 ;
        RECT 5.2840 28.9035 5.3100 29.9970 ;
        RECT 5.1760 28.9035 5.2020 29.9970 ;
        RECT 5.0680 28.9035 5.0940 29.9970 ;
        RECT 4.9600 28.9035 4.9860 29.9970 ;
        RECT 4.8520 28.9035 4.8780 29.9970 ;
        RECT 4.7440 28.9035 4.7700 29.9970 ;
        RECT 4.6360 28.9035 4.6620 29.9970 ;
        RECT 4.5280 28.9035 4.5540 29.9970 ;
        RECT 4.4200 28.9035 4.4460 29.9970 ;
        RECT 4.3120 28.9035 4.3380 29.9970 ;
        RECT 4.2040 28.9035 4.2300 29.9970 ;
        RECT 4.0960 28.9035 4.1220 29.9970 ;
        RECT 3.9880 28.9035 4.0140 29.9970 ;
        RECT 3.8800 28.9035 3.9060 29.9970 ;
        RECT 3.7720 28.9035 3.7980 29.9970 ;
        RECT 3.6640 28.9035 3.6900 29.9970 ;
        RECT 3.5560 28.9035 3.5820 29.9970 ;
        RECT 3.4480 28.9035 3.4740 29.9970 ;
        RECT 3.3400 28.9035 3.3660 29.9970 ;
        RECT 3.2320 28.9035 3.2580 29.9970 ;
        RECT 3.1240 28.9035 3.1500 29.9970 ;
        RECT 3.0160 28.9035 3.0420 29.9970 ;
        RECT 2.9080 28.9035 2.9340 29.9970 ;
        RECT 2.8000 28.9035 2.8260 29.9970 ;
        RECT 2.6920 28.9035 2.7180 29.9970 ;
        RECT 2.5840 28.9035 2.6100 29.9970 ;
        RECT 2.4760 28.9035 2.5020 29.9970 ;
        RECT 2.3680 28.9035 2.3940 29.9970 ;
        RECT 2.2600 28.9035 2.2860 29.9970 ;
        RECT 2.1520 28.9035 2.1780 29.9970 ;
        RECT 2.0440 28.9035 2.0700 29.9970 ;
        RECT 1.9360 28.9035 1.9620 29.9970 ;
        RECT 1.8280 28.9035 1.8540 29.9970 ;
        RECT 1.7200 28.9035 1.7460 29.9970 ;
        RECT 1.6120 28.9035 1.6380 29.9970 ;
        RECT 1.5040 28.9035 1.5300 29.9970 ;
        RECT 1.3960 28.9035 1.4220 29.9970 ;
        RECT 1.2880 28.9035 1.3140 29.9970 ;
        RECT 1.1800 28.9035 1.2060 29.9970 ;
        RECT 1.0720 28.9035 1.0980 29.9970 ;
        RECT 0.9640 28.9035 0.9900 29.9970 ;
        RECT 0.8560 28.9035 0.8820 29.9970 ;
        RECT 0.7480 28.9035 0.7740 29.9970 ;
        RECT 0.6400 28.9035 0.6660 29.9970 ;
        RECT 0.5320 28.9035 0.5580 29.9970 ;
        RECT 0.4240 28.9035 0.4500 29.9970 ;
        RECT 0.3160 28.9035 0.3420 29.9970 ;
        RECT 0.2080 28.9035 0.2340 29.9970 ;
        RECT 0.0050 28.9035 0.0900 29.9970 ;
        RECT 15.5530 29.9835 15.6810 31.0770 ;
        RECT 15.5390 30.6490 15.6810 30.9715 ;
        RECT 15.3190 30.3760 15.4530 31.0770 ;
        RECT 15.2960 30.7110 15.4530 30.9690 ;
        RECT 15.3190 29.9835 15.4170 31.0770 ;
        RECT 15.3190 30.1045 15.4310 30.3440 ;
        RECT 15.3190 29.9835 15.4530 30.0725 ;
        RECT 15.0940 30.4340 15.2280 31.0770 ;
        RECT 15.0940 29.9835 15.1920 31.0770 ;
        RECT 14.6770 29.9835 14.7600 31.0770 ;
        RECT 14.6770 30.0720 14.7740 31.0075 ;
        RECT 30.2680 29.9835 30.3530 31.0770 ;
        RECT 30.1240 29.9835 30.1500 31.0770 ;
        RECT 30.0160 29.9835 30.0420 31.0770 ;
        RECT 29.9080 29.9835 29.9340 31.0770 ;
        RECT 29.8000 29.9835 29.8260 31.0770 ;
        RECT 29.6920 29.9835 29.7180 31.0770 ;
        RECT 29.5840 29.9835 29.6100 31.0770 ;
        RECT 29.4760 29.9835 29.5020 31.0770 ;
        RECT 29.3680 29.9835 29.3940 31.0770 ;
        RECT 29.2600 29.9835 29.2860 31.0770 ;
        RECT 29.1520 29.9835 29.1780 31.0770 ;
        RECT 29.0440 29.9835 29.0700 31.0770 ;
        RECT 28.9360 29.9835 28.9620 31.0770 ;
        RECT 28.8280 29.9835 28.8540 31.0770 ;
        RECT 28.7200 29.9835 28.7460 31.0770 ;
        RECT 28.6120 29.9835 28.6380 31.0770 ;
        RECT 28.5040 29.9835 28.5300 31.0770 ;
        RECT 28.3960 29.9835 28.4220 31.0770 ;
        RECT 28.2880 29.9835 28.3140 31.0770 ;
        RECT 28.1800 29.9835 28.2060 31.0770 ;
        RECT 28.0720 29.9835 28.0980 31.0770 ;
        RECT 27.9640 29.9835 27.9900 31.0770 ;
        RECT 27.8560 29.9835 27.8820 31.0770 ;
        RECT 27.7480 29.9835 27.7740 31.0770 ;
        RECT 27.6400 29.9835 27.6660 31.0770 ;
        RECT 27.5320 29.9835 27.5580 31.0770 ;
        RECT 27.4240 29.9835 27.4500 31.0770 ;
        RECT 27.3160 29.9835 27.3420 31.0770 ;
        RECT 27.2080 29.9835 27.2340 31.0770 ;
        RECT 27.1000 29.9835 27.1260 31.0770 ;
        RECT 26.9920 29.9835 27.0180 31.0770 ;
        RECT 26.8840 29.9835 26.9100 31.0770 ;
        RECT 26.7760 29.9835 26.8020 31.0770 ;
        RECT 26.6680 29.9835 26.6940 31.0770 ;
        RECT 26.5600 29.9835 26.5860 31.0770 ;
        RECT 26.4520 29.9835 26.4780 31.0770 ;
        RECT 26.3440 29.9835 26.3700 31.0770 ;
        RECT 26.2360 29.9835 26.2620 31.0770 ;
        RECT 26.1280 29.9835 26.1540 31.0770 ;
        RECT 26.0200 29.9835 26.0460 31.0770 ;
        RECT 25.9120 29.9835 25.9380 31.0770 ;
        RECT 25.8040 29.9835 25.8300 31.0770 ;
        RECT 25.6960 29.9835 25.7220 31.0770 ;
        RECT 25.5880 29.9835 25.6140 31.0770 ;
        RECT 25.4800 29.9835 25.5060 31.0770 ;
        RECT 25.3720 29.9835 25.3980 31.0770 ;
        RECT 25.2640 29.9835 25.2900 31.0770 ;
        RECT 25.1560 29.9835 25.1820 31.0770 ;
        RECT 25.0480 29.9835 25.0740 31.0770 ;
        RECT 24.9400 29.9835 24.9660 31.0770 ;
        RECT 24.8320 29.9835 24.8580 31.0770 ;
        RECT 24.7240 29.9835 24.7500 31.0770 ;
        RECT 24.6160 29.9835 24.6420 31.0770 ;
        RECT 24.5080 29.9835 24.5340 31.0770 ;
        RECT 24.4000 29.9835 24.4260 31.0770 ;
        RECT 24.2920 29.9835 24.3180 31.0770 ;
        RECT 24.1840 29.9835 24.2100 31.0770 ;
        RECT 24.0760 29.9835 24.1020 31.0770 ;
        RECT 23.9680 29.9835 23.9940 31.0770 ;
        RECT 23.8600 29.9835 23.8860 31.0770 ;
        RECT 23.7520 29.9835 23.7780 31.0770 ;
        RECT 23.6440 29.9835 23.6700 31.0770 ;
        RECT 23.5360 29.9835 23.5620 31.0770 ;
        RECT 23.4280 29.9835 23.4540 31.0770 ;
        RECT 23.3200 29.9835 23.3460 31.0770 ;
        RECT 23.2120 29.9835 23.2380 31.0770 ;
        RECT 23.1040 29.9835 23.1300 31.0770 ;
        RECT 22.9960 29.9835 23.0220 31.0770 ;
        RECT 22.8880 29.9835 22.9140 31.0770 ;
        RECT 22.7800 29.9835 22.8060 31.0770 ;
        RECT 22.6720 29.9835 22.6980 31.0770 ;
        RECT 22.5640 29.9835 22.5900 31.0770 ;
        RECT 22.4560 29.9835 22.4820 31.0770 ;
        RECT 22.3480 29.9835 22.3740 31.0770 ;
        RECT 22.2400 29.9835 22.2660 31.0770 ;
        RECT 22.1320 29.9835 22.1580 31.0770 ;
        RECT 22.0240 29.9835 22.0500 31.0770 ;
        RECT 21.9160 29.9835 21.9420 31.0770 ;
        RECT 21.8080 29.9835 21.8340 31.0770 ;
        RECT 21.7000 29.9835 21.7260 31.0770 ;
        RECT 21.5920 29.9835 21.6180 31.0770 ;
        RECT 21.4840 29.9835 21.5100 31.0770 ;
        RECT 21.3760 29.9835 21.4020 31.0770 ;
        RECT 21.2680 29.9835 21.2940 31.0770 ;
        RECT 21.1600 29.9835 21.1860 31.0770 ;
        RECT 21.0520 29.9835 21.0780 31.0770 ;
        RECT 20.9440 29.9835 20.9700 31.0770 ;
        RECT 20.8360 29.9835 20.8620 31.0770 ;
        RECT 20.7280 29.9835 20.7540 31.0770 ;
        RECT 20.6200 29.9835 20.6460 31.0770 ;
        RECT 20.5120 29.9835 20.5380 31.0770 ;
        RECT 20.4040 29.9835 20.4300 31.0770 ;
        RECT 20.2960 29.9835 20.3220 31.0770 ;
        RECT 20.1880 29.9835 20.2140 31.0770 ;
        RECT 20.0800 29.9835 20.1060 31.0770 ;
        RECT 19.9720 29.9835 19.9980 31.0770 ;
        RECT 19.8640 29.9835 19.8900 31.0770 ;
        RECT 19.7560 29.9835 19.7820 31.0770 ;
        RECT 19.6480 29.9835 19.6740 31.0770 ;
        RECT 19.5400 29.9835 19.5660 31.0770 ;
        RECT 19.4320 29.9835 19.4580 31.0770 ;
        RECT 19.3240 29.9835 19.3500 31.0770 ;
        RECT 19.2160 29.9835 19.2420 31.0770 ;
        RECT 19.1080 29.9835 19.1340 31.0770 ;
        RECT 19.0000 29.9835 19.0260 31.0770 ;
        RECT 18.8920 29.9835 18.9180 31.0770 ;
        RECT 18.7840 29.9835 18.8100 31.0770 ;
        RECT 18.6760 29.9835 18.7020 31.0770 ;
        RECT 18.5680 29.9835 18.5940 31.0770 ;
        RECT 18.4600 29.9835 18.4860 31.0770 ;
        RECT 18.3520 29.9835 18.3780 31.0770 ;
        RECT 18.2440 29.9835 18.2700 31.0770 ;
        RECT 18.1360 29.9835 18.1620 31.0770 ;
        RECT 18.0280 29.9835 18.0540 31.0770 ;
        RECT 17.9200 29.9835 17.9460 31.0770 ;
        RECT 17.8120 29.9835 17.8380 31.0770 ;
        RECT 17.7040 29.9835 17.7300 31.0770 ;
        RECT 17.5960 29.9835 17.6220 31.0770 ;
        RECT 17.4880 29.9835 17.5140 31.0770 ;
        RECT 17.3800 29.9835 17.4060 31.0770 ;
        RECT 17.2720 29.9835 17.2980 31.0770 ;
        RECT 17.1640 29.9835 17.1900 31.0770 ;
        RECT 17.0560 29.9835 17.0820 31.0770 ;
        RECT 16.9480 29.9835 16.9740 31.0770 ;
        RECT 16.8400 29.9835 16.8660 31.0770 ;
        RECT 16.7320 29.9835 16.7580 31.0770 ;
        RECT 16.6240 29.9835 16.6500 31.0770 ;
        RECT 16.5160 29.9835 16.5420 31.0770 ;
        RECT 16.4080 29.9835 16.4340 31.0770 ;
        RECT 16.3000 29.9835 16.3260 31.0770 ;
        RECT 16.0870 29.9835 16.1640 31.0770 ;
        RECT 14.1940 29.9835 14.2710 31.0770 ;
        RECT 14.0320 29.9835 14.0580 31.0770 ;
        RECT 13.9240 29.9835 13.9500 31.0770 ;
        RECT 13.8160 29.9835 13.8420 31.0770 ;
        RECT 13.7080 29.9835 13.7340 31.0770 ;
        RECT 13.6000 29.9835 13.6260 31.0770 ;
        RECT 13.4920 29.9835 13.5180 31.0770 ;
        RECT 13.3840 29.9835 13.4100 31.0770 ;
        RECT 13.2760 29.9835 13.3020 31.0770 ;
        RECT 13.1680 29.9835 13.1940 31.0770 ;
        RECT 13.0600 29.9835 13.0860 31.0770 ;
        RECT 12.9520 29.9835 12.9780 31.0770 ;
        RECT 12.8440 29.9835 12.8700 31.0770 ;
        RECT 12.7360 29.9835 12.7620 31.0770 ;
        RECT 12.6280 29.9835 12.6540 31.0770 ;
        RECT 12.5200 29.9835 12.5460 31.0770 ;
        RECT 12.4120 29.9835 12.4380 31.0770 ;
        RECT 12.3040 29.9835 12.3300 31.0770 ;
        RECT 12.1960 29.9835 12.2220 31.0770 ;
        RECT 12.0880 29.9835 12.1140 31.0770 ;
        RECT 11.9800 29.9835 12.0060 31.0770 ;
        RECT 11.8720 29.9835 11.8980 31.0770 ;
        RECT 11.7640 29.9835 11.7900 31.0770 ;
        RECT 11.6560 29.9835 11.6820 31.0770 ;
        RECT 11.5480 29.9835 11.5740 31.0770 ;
        RECT 11.4400 29.9835 11.4660 31.0770 ;
        RECT 11.3320 29.9835 11.3580 31.0770 ;
        RECT 11.2240 29.9835 11.2500 31.0770 ;
        RECT 11.1160 29.9835 11.1420 31.0770 ;
        RECT 11.0080 29.9835 11.0340 31.0770 ;
        RECT 10.9000 29.9835 10.9260 31.0770 ;
        RECT 10.7920 29.9835 10.8180 31.0770 ;
        RECT 10.6840 29.9835 10.7100 31.0770 ;
        RECT 10.5760 29.9835 10.6020 31.0770 ;
        RECT 10.4680 29.9835 10.4940 31.0770 ;
        RECT 10.3600 29.9835 10.3860 31.0770 ;
        RECT 10.2520 29.9835 10.2780 31.0770 ;
        RECT 10.1440 29.9835 10.1700 31.0770 ;
        RECT 10.0360 29.9835 10.0620 31.0770 ;
        RECT 9.9280 29.9835 9.9540 31.0770 ;
        RECT 9.8200 29.9835 9.8460 31.0770 ;
        RECT 9.7120 29.9835 9.7380 31.0770 ;
        RECT 9.6040 29.9835 9.6300 31.0770 ;
        RECT 9.4960 29.9835 9.5220 31.0770 ;
        RECT 9.3880 29.9835 9.4140 31.0770 ;
        RECT 9.2800 29.9835 9.3060 31.0770 ;
        RECT 9.1720 29.9835 9.1980 31.0770 ;
        RECT 9.0640 29.9835 9.0900 31.0770 ;
        RECT 8.9560 29.9835 8.9820 31.0770 ;
        RECT 8.8480 29.9835 8.8740 31.0770 ;
        RECT 8.7400 29.9835 8.7660 31.0770 ;
        RECT 8.6320 29.9835 8.6580 31.0770 ;
        RECT 8.5240 29.9835 8.5500 31.0770 ;
        RECT 8.4160 29.9835 8.4420 31.0770 ;
        RECT 8.3080 29.9835 8.3340 31.0770 ;
        RECT 8.2000 29.9835 8.2260 31.0770 ;
        RECT 8.0920 29.9835 8.1180 31.0770 ;
        RECT 7.9840 29.9835 8.0100 31.0770 ;
        RECT 7.8760 29.9835 7.9020 31.0770 ;
        RECT 7.7680 29.9835 7.7940 31.0770 ;
        RECT 7.6600 29.9835 7.6860 31.0770 ;
        RECT 7.5520 29.9835 7.5780 31.0770 ;
        RECT 7.4440 29.9835 7.4700 31.0770 ;
        RECT 7.3360 29.9835 7.3620 31.0770 ;
        RECT 7.2280 29.9835 7.2540 31.0770 ;
        RECT 7.1200 29.9835 7.1460 31.0770 ;
        RECT 7.0120 29.9835 7.0380 31.0770 ;
        RECT 6.9040 29.9835 6.9300 31.0770 ;
        RECT 6.7960 29.9835 6.8220 31.0770 ;
        RECT 6.6880 29.9835 6.7140 31.0770 ;
        RECT 6.5800 29.9835 6.6060 31.0770 ;
        RECT 6.4720 29.9835 6.4980 31.0770 ;
        RECT 6.3640 29.9835 6.3900 31.0770 ;
        RECT 6.2560 29.9835 6.2820 31.0770 ;
        RECT 6.1480 29.9835 6.1740 31.0770 ;
        RECT 6.0400 29.9835 6.0660 31.0770 ;
        RECT 5.9320 29.9835 5.9580 31.0770 ;
        RECT 5.8240 29.9835 5.8500 31.0770 ;
        RECT 5.7160 29.9835 5.7420 31.0770 ;
        RECT 5.6080 29.9835 5.6340 31.0770 ;
        RECT 5.5000 29.9835 5.5260 31.0770 ;
        RECT 5.3920 29.9835 5.4180 31.0770 ;
        RECT 5.2840 29.9835 5.3100 31.0770 ;
        RECT 5.1760 29.9835 5.2020 31.0770 ;
        RECT 5.0680 29.9835 5.0940 31.0770 ;
        RECT 4.9600 29.9835 4.9860 31.0770 ;
        RECT 4.8520 29.9835 4.8780 31.0770 ;
        RECT 4.7440 29.9835 4.7700 31.0770 ;
        RECT 4.6360 29.9835 4.6620 31.0770 ;
        RECT 4.5280 29.9835 4.5540 31.0770 ;
        RECT 4.4200 29.9835 4.4460 31.0770 ;
        RECT 4.3120 29.9835 4.3380 31.0770 ;
        RECT 4.2040 29.9835 4.2300 31.0770 ;
        RECT 4.0960 29.9835 4.1220 31.0770 ;
        RECT 3.9880 29.9835 4.0140 31.0770 ;
        RECT 3.8800 29.9835 3.9060 31.0770 ;
        RECT 3.7720 29.9835 3.7980 31.0770 ;
        RECT 3.6640 29.9835 3.6900 31.0770 ;
        RECT 3.5560 29.9835 3.5820 31.0770 ;
        RECT 3.4480 29.9835 3.4740 31.0770 ;
        RECT 3.3400 29.9835 3.3660 31.0770 ;
        RECT 3.2320 29.9835 3.2580 31.0770 ;
        RECT 3.1240 29.9835 3.1500 31.0770 ;
        RECT 3.0160 29.9835 3.0420 31.0770 ;
        RECT 2.9080 29.9835 2.9340 31.0770 ;
        RECT 2.8000 29.9835 2.8260 31.0770 ;
        RECT 2.6920 29.9835 2.7180 31.0770 ;
        RECT 2.5840 29.9835 2.6100 31.0770 ;
        RECT 2.4760 29.9835 2.5020 31.0770 ;
        RECT 2.3680 29.9835 2.3940 31.0770 ;
        RECT 2.2600 29.9835 2.2860 31.0770 ;
        RECT 2.1520 29.9835 2.1780 31.0770 ;
        RECT 2.0440 29.9835 2.0700 31.0770 ;
        RECT 1.9360 29.9835 1.9620 31.0770 ;
        RECT 1.8280 29.9835 1.8540 31.0770 ;
        RECT 1.7200 29.9835 1.7460 31.0770 ;
        RECT 1.6120 29.9835 1.6380 31.0770 ;
        RECT 1.5040 29.9835 1.5300 31.0770 ;
        RECT 1.3960 29.9835 1.4220 31.0770 ;
        RECT 1.2880 29.9835 1.3140 31.0770 ;
        RECT 1.1800 29.9835 1.2060 31.0770 ;
        RECT 1.0720 29.9835 1.0980 31.0770 ;
        RECT 0.9640 29.9835 0.9900 31.0770 ;
        RECT 0.8560 29.9835 0.8820 31.0770 ;
        RECT 0.7480 29.9835 0.7740 31.0770 ;
        RECT 0.6400 29.9835 0.6660 31.0770 ;
        RECT 0.5320 29.9835 0.5580 31.0770 ;
        RECT 0.4240 29.9835 0.4500 31.0770 ;
        RECT 0.3160 29.9835 0.3420 31.0770 ;
        RECT 0.2080 29.9835 0.2340 31.0770 ;
        RECT 0.0050 29.9835 0.0900 31.0770 ;
        RECT 15.5530 31.0635 15.6810 32.1570 ;
        RECT 15.5390 31.7290 15.6810 32.0515 ;
        RECT 15.3190 31.4560 15.4530 32.1570 ;
        RECT 15.2960 31.7910 15.4530 32.0490 ;
        RECT 15.3190 31.0635 15.4170 32.1570 ;
        RECT 15.3190 31.1845 15.4310 31.4240 ;
        RECT 15.3190 31.0635 15.4530 31.1525 ;
        RECT 15.0940 31.5140 15.2280 32.1570 ;
        RECT 15.0940 31.0635 15.1920 32.1570 ;
        RECT 14.6770 31.0635 14.7600 32.1570 ;
        RECT 14.6770 31.1520 14.7740 32.0875 ;
        RECT 30.2680 31.0635 30.3530 32.1570 ;
        RECT 30.1240 31.0635 30.1500 32.1570 ;
        RECT 30.0160 31.0635 30.0420 32.1570 ;
        RECT 29.9080 31.0635 29.9340 32.1570 ;
        RECT 29.8000 31.0635 29.8260 32.1570 ;
        RECT 29.6920 31.0635 29.7180 32.1570 ;
        RECT 29.5840 31.0635 29.6100 32.1570 ;
        RECT 29.4760 31.0635 29.5020 32.1570 ;
        RECT 29.3680 31.0635 29.3940 32.1570 ;
        RECT 29.2600 31.0635 29.2860 32.1570 ;
        RECT 29.1520 31.0635 29.1780 32.1570 ;
        RECT 29.0440 31.0635 29.0700 32.1570 ;
        RECT 28.9360 31.0635 28.9620 32.1570 ;
        RECT 28.8280 31.0635 28.8540 32.1570 ;
        RECT 28.7200 31.0635 28.7460 32.1570 ;
        RECT 28.6120 31.0635 28.6380 32.1570 ;
        RECT 28.5040 31.0635 28.5300 32.1570 ;
        RECT 28.3960 31.0635 28.4220 32.1570 ;
        RECT 28.2880 31.0635 28.3140 32.1570 ;
        RECT 28.1800 31.0635 28.2060 32.1570 ;
        RECT 28.0720 31.0635 28.0980 32.1570 ;
        RECT 27.9640 31.0635 27.9900 32.1570 ;
        RECT 27.8560 31.0635 27.8820 32.1570 ;
        RECT 27.7480 31.0635 27.7740 32.1570 ;
        RECT 27.6400 31.0635 27.6660 32.1570 ;
        RECT 27.5320 31.0635 27.5580 32.1570 ;
        RECT 27.4240 31.0635 27.4500 32.1570 ;
        RECT 27.3160 31.0635 27.3420 32.1570 ;
        RECT 27.2080 31.0635 27.2340 32.1570 ;
        RECT 27.1000 31.0635 27.1260 32.1570 ;
        RECT 26.9920 31.0635 27.0180 32.1570 ;
        RECT 26.8840 31.0635 26.9100 32.1570 ;
        RECT 26.7760 31.0635 26.8020 32.1570 ;
        RECT 26.6680 31.0635 26.6940 32.1570 ;
        RECT 26.5600 31.0635 26.5860 32.1570 ;
        RECT 26.4520 31.0635 26.4780 32.1570 ;
        RECT 26.3440 31.0635 26.3700 32.1570 ;
        RECT 26.2360 31.0635 26.2620 32.1570 ;
        RECT 26.1280 31.0635 26.1540 32.1570 ;
        RECT 26.0200 31.0635 26.0460 32.1570 ;
        RECT 25.9120 31.0635 25.9380 32.1570 ;
        RECT 25.8040 31.0635 25.8300 32.1570 ;
        RECT 25.6960 31.0635 25.7220 32.1570 ;
        RECT 25.5880 31.0635 25.6140 32.1570 ;
        RECT 25.4800 31.0635 25.5060 32.1570 ;
        RECT 25.3720 31.0635 25.3980 32.1570 ;
        RECT 25.2640 31.0635 25.2900 32.1570 ;
        RECT 25.1560 31.0635 25.1820 32.1570 ;
        RECT 25.0480 31.0635 25.0740 32.1570 ;
        RECT 24.9400 31.0635 24.9660 32.1570 ;
        RECT 24.8320 31.0635 24.8580 32.1570 ;
        RECT 24.7240 31.0635 24.7500 32.1570 ;
        RECT 24.6160 31.0635 24.6420 32.1570 ;
        RECT 24.5080 31.0635 24.5340 32.1570 ;
        RECT 24.4000 31.0635 24.4260 32.1570 ;
        RECT 24.2920 31.0635 24.3180 32.1570 ;
        RECT 24.1840 31.0635 24.2100 32.1570 ;
        RECT 24.0760 31.0635 24.1020 32.1570 ;
        RECT 23.9680 31.0635 23.9940 32.1570 ;
        RECT 23.8600 31.0635 23.8860 32.1570 ;
        RECT 23.7520 31.0635 23.7780 32.1570 ;
        RECT 23.6440 31.0635 23.6700 32.1570 ;
        RECT 23.5360 31.0635 23.5620 32.1570 ;
        RECT 23.4280 31.0635 23.4540 32.1570 ;
        RECT 23.3200 31.0635 23.3460 32.1570 ;
        RECT 23.2120 31.0635 23.2380 32.1570 ;
        RECT 23.1040 31.0635 23.1300 32.1570 ;
        RECT 22.9960 31.0635 23.0220 32.1570 ;
        RECT 22.8880 31.0635 22.9140 32.1570 ;
        RECT 22.7800 31.0635 22.8060 32.1570 ;
        RECT 22.6720 31.0635 22.6980 32.1570 ;
        RECT 22.5640 31.0635 22.5900 32.1570 ;
        RECT 22.4560 31.0635 22.4820 32.1570 ;
        RECT 22.3480 31.0635 22.3740 32.1570 ;
        RECT 22.2400 31.0635 22.2660 32.1570 ;
        RECT 22.1320 31.0635 22.1580 32.1570 ;
        RECT 22.0240 31.0635 22.0500 32.1570 ;
        RECT 21.9160 31.0635 21.9420 32.1570 ;
        RECT 21.8080 31.0635 21.8340 32.1570 ;
        RECT 21.7000 31.0635 21.7260 32.1570 ;
        RECT 21.5920 31.0635 21.6180 32.1570 ;
        RECT 21.4840 31.0635 21.5100 32.1570 ;
        RECT 21.3760 31.0635 21.4020 32.1570 ;
        RECT 21.2680 31.0635 21.2940 32.1570 ;
        RECT 21.1600 31.0635 21.1860 32.1570 ;
        RECT 21.0520 31.0635 21.0780 32.1570 ;
        RECT 20.9440 31.0635 20.9700 32.1570 ;
        RECT 20.8360 31.0635 20.8620 32.1570 ;
        RECT 20.7280 31.0635 20.7540 32.1570 ;
        RECT 20.6200 31.0635 20.6460 32.1570 ;
        RECT 20.5120 31.0635 20.5380 32.1570 ;
        RECT 20.4040 31.0635 20.4300 32.1570 ;
        RECT 20.2960 31.0635 20.3220 32.1570 ;
        RECT 20.1880 31.0635 20.2140 32.1570 ;
        RECT 20.0800 31.0635 20.1060 32.1570 ;
        RECT 19.9720 31.0635 19.9980 32.1570 ;
        RECT 19.8640 31.0635 19.8900 32.1570 ;
        RECT 19.7560 31.0635 19.7820 32.1570 ;
        RECT 19.6480 31.0635 19.6740 32.1570 ;
        RECT 19.5400 31.0635 19.5660 32.1570 ;
        RECT 19.4320 31.0635 19.4580 32.1570 ;
        RECT 19.3240 31.0635 19.3500 32.1570 ;
        RECT 19.2160 31.0635 19.2420 32.1570 ;
        RECT 19.1080 31.0635 19.1340 32.1570 ;
        RECT 19.0000 31.0635 19.0260 32.1570 ;
        RECT 18.8920 31.0635 18.9180 32.1570 ;
        RECT 18.7840 31.0635 18.8100 32.1570 ;
        RECT 18.6760 31.0635 18.7020 32.1570 ;
        RECT 18.5680 31.0635 18.5940 32.1570 ;
        RECT 18.4600 31.0635 18.4860 32.1570 ;
        RECT 18.3520 31.0635 18.3780 32.1570 ;
        RECT 18.2440 31.0635 18.2700 32.1570 ;
        RECT 18.1360 31.0635 18.1620 32.1570 ;
        RECT 18.0280 31.0635 18.0540 32.1570 ;
        RECT 17.9200 31.0635 17.9460 32.1570 ;
        RECT 17.8120 31.0635 17.8380 32.1570 ;
        RECT 17.7040 31.0635 17.7300 32.1570 ;
        RECT 17.5960 31.0635 17.6220 32.1570 ;
        RECT 17.4880 31.0635 17.5140 32.1570 ;
        RECT 17.3800 31.0635 17.4060 32.1570 ;
        RECT 17.2720 31.0635 17.2980 32.1570 ;
        RECT 17.1640 31.0635 17.1900 32.1570 ;
        RECT 17.0560 31.0635 17.0820 32.1570 ;
        RECT 16.9480 31.0635 16.9740 32.1570 ;
        RECT 16.8400 31.0635 16.8660 32.1570 ;
        RECT 16.7320 31.0635 16.7580 32.1570 ;
        RECT 16.6240 31.0635 16.6500 32.1570 ;
        RECT 16.5160 31.0635 16.5420 32.1570 ;
        RECT 16.4080 31.0635 16.4340 32.1570 ;
        RECT 16.3000 31.0635 16.3260 32.1570 ;
        RECT 16.0870 31.0635 16.1640 32.1570 ;
        RECT 14.1940 31.0635 14.2710 32.1570 ;
        RECT 14.0320 31.0635 14.0580 32.1570 ;
        RECT 13.9240 31.0635 13.9500 32.1570 ;
        RECT 13.8160 31.0635 13.8420 32.1570 ;
        RECT 13.7080 31.0635 13.7340 32.1570 ;
        RECT 13.6000 31.0635 13.6260 32.1570 ;
        RECT 13.4920 31.0635 13.5180 32.1570 ;
        RECT 13.3840 31.0635 13.4100 32.1570 ;
        RECT 13.2760 31.0635 13.3020 32.1570 ;
        RECT 13.1680 31.0635 13.1940 32.1570 ;
        RECT 13.0600 31.0635 13.0860 32.1570 ;
        RECT 12.9520 31.0635 12.9780 32.1570 ;
        RECT 12.8440 31.0635 12.8700 32.1570 ;
        RECT 12.7360 31.0635 12.7620 32.1570 ;
        RECT 12.6280 31.0635 12.6540 32.1570 ;
        RECT 12.5200 31.0635 12.5460 32.1570 ;
        RECT 12.4120 31.0635 12.4380 32.1570 ;
        RECT 12.3040 31.0635 12.3300 32.1570 ;
        RECT 12.1960 31.0635 12.2220 32.1570 ;
        RECT 12.0880 31.0635 12.1140 32.1570 ;
        RECT 11.9800 31.0635 12.0060 32.1570 ;
        RECT 11.8720 31.0635 11.8980 32.1570 ;
        RECT 11.7640 31.0635 11.7900 32.1570 ;
        RECT 11.6560 31.0635 11.6820 32.1570 ;
        RECT 11.5480 31.0635 11.5740 32.1570 ;
        RECT 11.4400 31.0635 11.4660 32.1570 ;
        RECT 11.3320 31.0635 11.3580 32.1570 ;
        RECT 11.2240 31.0635 11.2500 32.1570 ;
        RECT 11.1160 31.0635 11.1420 32.1570 ;
        RECT 11.0080 31.0635 11.0340 32.1570 ;
        RECT 10.9000 31.0635 10.9260 32.1570 ;
        RECT 10.7920 31.0635 10.8180 32.1570 ;
        RECT 10.6840 31.0635 10.7100 32.1570 ;
        RECT 10.5760 31.0635 10.6020 32.1570 ;
        RECT 10.4680 31.0635 10.4940 32.1570 ;
        RECT 10.3600 31.0635 10.3860 32.1570 ;
        RECT 10.2520 31.0635 10.2780 32.1570 ;
        RECT 10.1440 31.0635 10.1700 32.1570 ;
        RECT 10.0360 31.0635 10.0620 32.1570 ;
        RECT 9.9280 31.0635 9.9540 32.1570 ;
        RECT 9.8200 31.0635 9.8460 32.1570 ;
        RECT 9.7120 31.0635 9.7380 32.1570 ;
        RECT 9.6040 31.0635 9.6300 32.1570 ;
        RECT 9.4960 31.0635 9.5220 32.1570 ;
        RECT 9.3880 31.0635 9.4140 32.1570 ;
        RECT 9.2800 31.0635 9.3060 32.1570 ;
        RECT 9.1720 31.0635 9.1980 32.1570 ;
        RECT 9.0640 31.0635 9.0900 32.1570 ;
        RECT 8.9560 31.0635 8.9820 32.1570 ;
        RECT 8.8480 31.0635 8.8740 32.1570 ;
        RECT 8.7400 31.0635 8.7660 32.1570 ;
        RECT 8.6320 31.0635 8.6580 32.1570 ;
        RECT 8.5240 31.0635 8.5500 32.1570 ;
        RECT 8.4160 31.0635 8.4420 32.1570 ;
        RECT 8.3080 31.0635 8.3340 32.1570 ;
        RECT 8.2000 31.0635 8.2260 32.1570 ;
        RECT 8.0920 31.0635 8.1180 32.1570 ;
        RECT 7.9840 31.0635 8.0100 32.1570 ;
        RECT 7.8760 31.0635 7.9020 32.1570 ;
        RECT 7.7680 31.0635 7.7940 32.1570 ;
        RECT 7.6600 31.0635 7.6860 32.1570 ;
        RECT 7.5520 31.0635 7.5780 32.1570 ;
        RECT 7.4440 31.0635 7.4700 32.1570 ;
        RECT 7.3360 31.0635 7.3620 32.1570 ;
        RECT 7.2280 31.0635 7.2540 32.1570 ;
        RECT 7.1200 31.0635 7.1460 32.1570 ;
        RECT 7.0120 31.0635 7.0380 32.1570 ;
        RECT 6.9040 31.0635 6.9300 32.1570 ;
        RECT 6.7960 31.0635 6.8220 32.1570 ;
        RECT 6.6880 31.0635 6.7140 32.1570 ;
        RECT 6.5800 31.0635 6.6060 32.1570 ;
        RECT 6.4720 31.0635 6.4980 32.1570 ;
        RECT 6.3640 31.0635 6.3900 32.1570 ;
        RECT 6.2560 31.0635 6.2820 32.1570 ;
        RECT 6.1480 31.0635 6.1740 32.1570 ;
        RECT 6.0400 31.0635 6.0660 32.1570 ;
        RECT 5.9320 31.0635 5.9580 32.1570 ;
        RECT 5.8240 31.0635 5.8500 32.1570 ;
        RECT 5.7160 31.0635 5.7420 32.1570 ;
        RECT 5.6080 31.0635 5.6340 32.1570 ;
        RECT 5.5000 31.0635 5.5260 32.1570 ;
        RECT 5.3920 31.0635 5.4180 32.1570 ;
        RECT 5.2840 31.0635 5.3100 32.1570 ;
        RECT 5.1760 31.0635 5.2020 32.1570 ;
        RECT 5.0680 31.0635 5.0940 32.1570 ;
        RECT 4.9600 31.0635 4.9860 32.1570 ;
        RECT 4.8520 31.0635 4.8780 32.1570 ;
        RECT 4.7440 31.0635 4.7700 32.1570 ;
        RECT 4.6360 31.0635 4.6620 32.1570 ;
        RECT 4.5280 31.0635 4.5540 32.1570 ;
        RECT 4.4200 31.0635 4.4460 32.1570 ;
        RECT 4.3120 31.0635 4.3380 32.1570 ;
        RECT 4.2040 31.0635 4.2300 32.1570 ;
        RECT 4.0960 31.0635 4.1220 32.1570 ;
        RECT 3.9880 31.0635 4.0140 32.1570 ;
        RECT 3.8800 31.0635 3.9060 32.1570 ;
        RECT 3.7720 31.0635 3.7980 32.1570 ;
        RECT 3.6640 31.0635 3.6900 32.1570 ;
        RECT 3.5560 31.0635 3.5820 32.1570 ;
        RECT 3.4480 31.0635 3.4740 32.1570 ;
        RECT 3.3400 31.0635 3.3660 32.1570 ;
        RECT 3.2320 31.0635 3.2580 32.1570 ;
        RECT 3.1240 31.0635 3.1500 32.1570 ;
        RECT 3.0160 31.0635 3.0420 32.1570 ;
        RECT 2.9080 31.0635 2.9340 32.1570 ;
        RECT 2.8000 31.0635 2.8260 32.1570 ;
        RECT 2.6920 31.0635 2.7180 32.1570 ;
        RECT 2.5840 31.0635 2.6100 32.1570 ;
        RECT 2.4760 31.0635 2.5020 32.1570 ;
        RECT 2.3680 31.0635 2.3940 32.1570 ;
        RECT 2.2600 31.0635 2.2860 32.1570 ;
        RECT 2.1520 31.0635 2.1780 32.1570 ;
        RECT 2.0440 31.0635 2.0700 32.1570 ;
        RECT 1.9360 31.0635 1.9620 32.1570 ;
        RECT 1.8280 31.0635 1.8540 32.1570 ;
        RECT 1.7200 31.0635 1.7460 32.1570 ;
        RECT 1.6120 31.0635 1.6380 32.1570 ;
        RECT 1.5040 31.0635 1.5300 32.1570 ;
        RECT 1.3960 31.0635 1.4220 32.1570 ;
        RECT 1.2880 31.0635 1.3140 32.1570 ;
        RECT 1.1800 31.0635 1.2060 32.1570 ;
        RECT 1.0720 31.0635 1.0980 32.1570 ;
        RECT 0.9640 31.0635 0.9900 32.1570 ;
        RECT 0.8560 31.0635 0.8820 32.1570 ;
        RECT 0.7480 31.0635 0.7740 32.1570 ;
        RECT 0.6400 31.0635 0.6660 32.1570 ;
        RECT 0.5320 31.0635 0.5580 32.1570 ;
        RECT 0.4240 31.0635 0.4500 32.1570 ;
        RECT 0.3160 31.0635 0.3420 32.1570 ;
        RECT 0.2080 31.0635 0.2340 32.1570 ;
        RECT 0.0050 31.0635 0.0900 32.1570 ;
        RECT 15.5530 32.1435 15.6810 33.2370 ;
        RECT 15.5390 32.8090 15.6810 33.1315 ;
        RECT 15.3190 32.5360 15.4530 33.2370 ;
        RECT 15.2960 32.8710 15.4530 33.1290 ;
        RECT 15.3190 32.1435 15.4170 33.2370 ;
        RECT 15.3190 32.2645 15.4310 32.5040 ;
        RECT 15.3190 32.1435 15.4530 32.2325 ;
        RECT 15.0940 32.5940 15.2280 33.2370 ;
        RECT 15.0940 32.1435 15.1920 33.2370 ;
        RECT 14.6770 32.1435 14.7600 33.2370 ;
        RECT 14.6770 32.2320 14.7740 33.1675 ;
        RECT 30.2680 32.1435 30.3530 33.2370 ;
        RECT 30.1240 32.1435 30.1500 33.2370 ;
        RECT 30.0160 32.1435 30.0420 33.2370 ;
        RECT 29.9080 32.1435 29.9340 33.2370 ;
        RECT 29.8000 32.1435 29.8260 33.2370 ;
        RECT 29.6920 32.1435 29.7180 33.2370 ;
        RECT 29.5840 32.1435 29.6100 33.2370 ;
        RECT 29.4760 32.1435 29.5020 33.2370 ;
        RECT 29.3680 32.1435 29.3940 33.2370 ;
        RECT 29.2600 32.1435 29.2860 33.2370 ;
        RECT 29.1520 32.1435 29.1780 33.2370 ;
        RECT 29.0440 32.1435 29.0700 33.2370 ;
        RECT 28.9360 32.1435 28.9620 33.2370 ;
        RECT 28.8280 32.1435 28.8540 33.2370 ;
        RECT 28.7200 32.1435 28.7460 33.2370 ;
        RECT 28.6120 32.1435 28.6380 33.2370 ;
        RECT 28.5040 32.1435 28.5300 33.2370 ;
        RECT 28.3960 32.1435 28.4220 33.2370 ;
        RECT 28.2880 32.1435 28.3140 33.2370 ;
        RECT 28.1800 32.1435 28.2060 33.2370 ;
        RECT 28.0720 32.1435 28.0980 33.2370 ;
        RECT 27.9640 32.1435 27.9900 33.2370 ;
        RECT 27.8560 32.1435 27.8820 33.2370 ;
        RECT 27.7480 32.1435 27.7740 33.2370 ;
        RECT 27.6400 32.1435 27.6660 33.2370 ;
        RECT 27.5320 32.1435 27.5580 33.2370 ;
        RECT 27.4240 32.1435 27.4500 33.2370 ;
        RECT 27.3160 32.1435 27.3420 33.2370 ;
        RECT 27.2080 32.1435 27.2340 33.2370 ;
        RECT 27.1000 32.1435 27.1260 33.2370 ;
        RECT 26.9920 32.1435 27.0180 33.2370 ;
        RECT 26.8840 32.1435 26.9100 33.2370 ;
        RECT 26.7760 32.1435 26.8020 33.2370 ;
        RECT 26.6680 32.1435 26.6940 33.2370 ;
        RECT 26.5600 32.1435 26.5860 33.2370 ;
        RECT 26.4520 32.1435 26.4780 33.2370 ;
        RECT 26.3440 32.1435 26.3700 33.2370 ;
        RECT 26.2360 32.1435 26.2620 33.2370 ;
        RECT 26.1280 32.1435 26.1540 33.2370 ;
        RECT 26.0200 32.1435 26.0460 33.2370 ;
        RECT 25.9120 32.1435 25.9380 33.2370 ;
        RECT 25.8040 32.1435 25.8300 33.2370 ;
        RECT 25.6960 32.1435 25.7220 33.2370 ;
        RECT 25.5880 32.1435 25.6140 33.2370 ;
        RECT 25.4800 32.1435 25.5060 33.2370 ;
        RECT 25.3720 32.1435 25.3980 33.2370 ;
        RECT 25.2640 32.1435 25.2900 33.2370 ;
        RECT 25.1560 32.1435 25.1820 33.2370 ;
        RECT 25.0480 32.1435 25.0740 33.2370 ;
        RECT 24.9400 32.1435 24.9660 33.2370 ;
        RECT 24.8320 32.1435 24.8580 33.2370 ;
        RECT 24.7240 32.1435 24.7500 33.2370 ;
        RECT 24.6160 32.1435 24.6420 33.2370 ;
        RECT 24.5080 32.1435 24.5340 33.2370 ;
        RECT 24.4000 32.1435 24.4260 33.2370 ;
        RECT 24.2920 32.1435 24.3180 33.2370 ;
        RECT 24.1840 32.1435 24.2100 33.2370 ;
        RECT 24.0760 32.1435 24.1020 33.2370 ;
        RECT 23.9680 32.1435 23.9940 33.2370 ;
        RECT 23.8600 32.1435 23.8860 33.2370 ;
        RECT 23.7520 32.1435 23.7780 33.2370 ;
        RECT 23.6440 32.1435 23.6700 33.2370 ;
        RECT 23.5360 32.1435 23.5620 33.2370 ;
        RECT 23.4280 32.1435 23.4540 33.2370 ;
        RECT 23.3200 32.1435 23.3460 33.2370 ;
        RECT 23.2120 32.1435 23.2380 33.2370 ;
        RECT 23.1040 32.1435 23.1300 33.2370 ;
        RECT 22.9960 32.1435 23.0220 33.2370 ;
        RECT 22.8880 32.1435 22.9140 33.2370 ;
        RECT 22.7800 32.1435 22.8060 33.2370 ;
        RECT 22.6720 32.1435 22.6980 33.2370 ;
        RECT 22.5640 32.1435 22.5900 33.2370 ;
        RECT 22.4560 32.1435 22.4820 33.2370 ;
        RECT 22.3480 32.1435 22.3740 33.2370 ;
        RECT 22.2400 32.1435 22.2660 33.2370 ;
        RECT 22.1320 32.1435 22.1580 33.2370 ;
        RECT 22.0240 32.1435 22.0500 33.2370 ;
        RECT 21.9160 32.1435 21.9420 33.2370 ;
        RECT 21.8080 32.1435 21.8340 33.2370 ;
        RECT 21.7000 32.1435 21.7260 33.2370 ;
        RECT 21.5920 32.1435 21.6180 33.2370 ;
        RECT 21.4840 32.1435 21.5100 33.2370 ;
        RECT 21.3760 32.1435 21.4020 33.2370 ;
        RECT 21.2680 32.1435 21.2940 33.2370 ;
        RECT 21.1600 32.1435 21.1860 33.2370 ;
        RECT 21.0520 32.1435 21.0780 33.2370 ;
        RECT 20.9440 32.1435 20.9700 33.2370 ;
        RECT 20.8360 32.1435 20.8620 33.2370 ;
        RECT 20.7280 32.1435 20.7540 33.2370 ;
        RECT 20.6200 32.1435 20.6460 33.2370 ;
        RECT 20.5120 32.1435 20.5380 33.2370 ;
        RECT 20.4040 32.1435 20.4300 33.2370 ;
        RECT 20.2960 32.1435 20.3220 33.2370 ;
        RECT 20.1880 32.1435 20.2140 33.2370 ;
        RECT 20.0800 32.1435 20.1060 33.2370 ;
        RECT 19.9720 32.1435 19.9980 33.2370 ;
        RECT 19.8640 32.1435 19.8900 33.2370 ;
        RECT 19.7560 32.1435 19.7820 33.2370 ;
        RECT 19.6480 32.1435 19.6740 33.2370 ;
        RECT 19.5400 32.1435 19.5660 33.2370 ;
        RECT 19.4320 32.1435 19.4580 33.2370 ;
        RECT 19.3240 32.1435 19.3500 33.2370 ;
        RECT 19.2160 32.1435 19.2420 33.2370 ;
        RECT 19.1080 32.1435 19.1340 33.2370 ;
        RECT 19.0000 32.1435 19.0260 33.2370 ;
        RECT 18.8920 32.1435 18.9180 33.2370 ;
        RECT 18.7840 32.1435 18.8100 33.2370 ;
        RECT 18.6760 32.1435 18.7020 33.2370 ;
        RECT 18.5680 32.1435 18.5940 33.2370 ;
        RECT 18.4600 32.1435 18.4860 33.2370 ;
        RECT 18.3520 32.1435 18.3780 33.2370 ;
        RECT 18.2440 32.1435 18.2700 33.2370 ;
        RECT 18.1360 32.1435 18.1620 33.2370 ;
        RECT 18.0280 32.1435 18.0540 33.2370 ;
        RECT 17.9200 32.1435 17.9460 33.2370 ;
        RECT 17.8120 32.1435 17.8380 33.2370 ;
        RECT 17.7040 32.1435 17.7300 33.2370 ;
        RECT 17.5960 32.1435 17.6220 33.2370 ;
        RECT 17.4880 32.1435 17.5140 33.2370 ;
        RECT 17.3800 32.1435 17.4060 33.2370 ;
        RECT 17.2720 32.1435 17.2980 33.2370 ;
        RECT 17.1640 32.1435 17.1900 33.2370 ;
        RECT 17.0560 32.1435 17.0820 33.2370 ;
        RECT 16.9480 32.1435 16.9740 33.2370 ;
        RECT 16.8400 32.1435 16.8660 33.2370 ;
        RECT 16.7320 32.1435 16.7580 33.2370 ;
        RECT 16.6240 32.1435 16.6500 33.2370 ;
        RECT 16.5160 32.1435 16.5420 33.2370 ;
        RECT 16.4080 32.1435 16.4340 33.2370 ;
        RECT 16.3000 32.1435 16.3260 33.2370 ;
        RECT 16.0870 32.1435 16.1640 33.2370 ;
        RECT 14.1940 32.1435 14.2710 33.2370 ;
        RECT 14.0320 32.1435 14.0580 33.2370 ;
        RECT 13.9240 32.1435 13.9500 33.2370 ;
        RECT 13.8160 32.1435 13.8420 33.2370 ;
        RECT 13.7080 32.1435 13.7340 33.2370 ;
        RECT 13.6000 32.1435 13.6260 33.2370 ;
        RECT 13.4920 32.1435 13.5180 33.2370 ;
        RECT 13.3840 32.1435 13.4100 33.2370 ;
        RECT 13.2760 32.1435 13.3020 33.2370 ;
        RECT 13.1680 32.1435 13.1940 33.2370 ;
        RECT 13.0600 32.1435 13.0860 33.2370 ;
        RECT 12.9520 32.1435 12.9780 33.2370 ;
        RECT 12.8440 32.1435 12.8700 33.2370 ;
        RECT 12.7360 32.1435 12.7620 33.2370 ;
        RECT 12.6280 32.1435 12.6540 33.2370 ;
        RECT 12.5200 32.1435 12.5460 33.2370 ;
        RECT 12.4120 32.1435 12.4380 33.2370 ;
        RECT 12.3040 32.1435 12.3300 33.2370 ;
        RECT 12.1960 32.1435 12.2220 33.2370 ;
        RECT 12.0880 32.1435 12.1140 33.2370 ;
        RECT 11.9800 32.1435 12.0060 33.2370 ;
        RECT 11.8720 32.1435 11.8980 33.2370 ;
        RECT 11.7640 32.1435 11.7900 33.2370 ;
        RECT 11.6560 32.1435 11.6820 33.2370 ;
        RECT 11.5480 32.1435 11.5740 33.2370 ;
        RECT 11.4400 32.1435 11.4660 33.2370 ;
        RECT 11.3320 32.1435 11.3580 33.2370 ;
        RECT 11.2240 32.1435 11.2500 33.2370 ;
        RECT 11.1160 32.1435 11.1420 33.2370 ;
        RECT 11.0080 32.1435 11.0340 33.2370 ;
        RECT 10.9000 32.1435 10.9260 33.2370 ;
        RECT 10.7920 32.1435 10.8180 33.2370 ;
        RECT 10.6840 32.1435 10.7100 33.2370 ;
        RECT 10.5760 32.1435 10.6020 33.2370 ;
        RECT 10.4680 32.1435 10.4940 33.2370 ;
        RECT 10.3600 32.1435 10.3860 33.2370 ;
        RECT 10.2520 32.1435 10.2780 33.2370 ;
        RECT 10.1440 32.1435 10.1700 33.2370 ;
        RECT 10.0360 32.1435 10.0620 33.2370 ;
        RECT 9.9280 32.1435 9.9540 33.2370 ;
        RECT 9.8200 32.1435 9.8460 33.2370 ;
        RECT 9.7120 32.1435 9.7380 33.2370 ;
        RECT 9.6040 32.1435 9.6300 33.2370 ;
        RECT 9.4960 32.1435 9.5220 33.2370 ;
        RECT 9.3880 32.1435 9.4140 33.2370 ;
        RECT 9.2800 32.1435 9.3060 33.2370 ;
        RECT 9.1720 32.1435 9.1980 33.2370 ;
        RECT 9.0640 32.1435 9.0900 33.2370 ;
        RECT 8.9560 32.1435 8.9820 33.2370 ;
        RECT 8.8480 32.1435 8.8740 33.2370 ;
        RECT 8.7400 32.1435 8.7660 33.2370 ;
        RECT 8.6320 32.1435 8.6580 33.2370 ;
        RECT 8.5240 32.1435 8.5500 33.2370 ;
        RECT 8.4160 32.1435 8.4420 33.2370 ;
        RECT 8.3080 32.1435 8.3340 33.2370 ;
        RECT 8.2000 32.1435 8.2260 33.2370 ;
        RECT 8.0920 32.1435 8.1180 33.2370 ;
        RECT 7.9840 32.1435 8.0100 33.2370 ;
        RECT 7.8760 32.1435 7.9020 33.2370 ;
        RECT 7.7680 32.1435 7.7940 33.2370 ;
        RECT 7.6600 32.1435 7.6860 33.2370 ;
        RECT 7.5520 32.1435 7.5780 33.2370 ;
        RECT 7.4440 32.1435 7.4700 33.2370 ;
        RECT 7.3360 32.1435 7.3620 33.2370 ;
        RECT 7.2280 32.1435 7.2540 33.2370 ;
        RECT 7.1200 32.1435 7.1460 33.2370 ;
        RECT 7.0120 32.1435 7.0380 33.2370 ;
        RECT 6.9040 32.1435 6.9300 33.2370 ;
        RECT 6.7960 32.1435 6.8220 33.2370 ;
        RECT 6.6880 32.1435 6.7140 33.2370 ;
        RECT 6.5800 32.1435 6.6060 33.2370 ;
        RECT 6.4720 32.1435 6.4980 33.2370 ;
        RECT 6.3640 32.1435 6.3900 33.2370 ;
        RECT 6.2560 32.1435 6.2820 33.2370 ;
        RECT 6.1480 32.1435 6.1740 33.2370 ;
        RECT 6.0400 32.1435 6.0660 33.2370 ;
        RECT 5.9320 32.1435 5.9580 33.2370 ;
        RECT 5.8240 32.1435 5.8500 33.2370 ;
        RECT 5.7160 32.1435 5.7420 33.2370 ;
        RECT 5.6080 32.1435 5.6340 33.2370 ;
        RECT 5.5000 32.1435 5.5260 33.2370 ;
        RECT 5.3920 32.1435 5.4180 33.2370 ;
        RECT 5.2840 32.1435 5.3100 33.2370 ;
        RECT 5.1760 32.1435 5.2020 33.2370 ;
        RECT 5.0680 32.1435 5.0940 33.2370 ;
        RECT 4.9600 32.1435 4.9860 33.2370 ;
        RECT 4.8520 32.1435 4.8780 33.2370 ;
        RECT 4.7440 32.1435 4.7700 33.2370 ;
        RECT 4.6360 32.1435 4.6620 33.2370 ;
        RECT 4.5280 32.1435 4.5540 33.2370 ;
        RECT 4.4200 32.1435 4.4460 33.2370 ;
        RECT 4.3120 32.1435 4.3380 33.2370 ;
        RECT 4.2040 32.1435 4.2300 33.2370 ;
        RECT 4.0960 32.1435 4.1220 33.2370 ;
        RECT 3.9880 32.1435 4.0140 33.2370 ;
        RECT 3.8800 32.1435 3.9060 33.2370 ;
        RECT 3.7720 32.1435 3.7980 33.2370 ;
        RECT 3.6640 32.1435 3.6900 33.2370 ;
        RECT 3.5560 32.1435 3.5820 33.2370 ;
        RECT 3.4480 32.1435 3.4740 33.2370 ;
        RECT 3.3400 32.1435 3.3660 33.2370 ;
        RECT 3.2320 32.1435 3.2580 33.2370 ;
        RECT 3.1240 32.1435 3.1500 33.2370 ;
        RECT 3.0160 32.1435 3.0420 33.2370 ;
        RECT 2.9080 32.1435 2.9340 33.2370 ;
        RECT 2.8000 32.1435 2.8260 33.2370 ;
        RECT 2.6920 32.1435 2.7180 33.2370 ;
        RECT 2.5840 32.1435 2.6100 33.2370 ;
        RECT 2.4760 32.1435 2.5020 33.2370 ;
        RECT 2.3680 32.1435 2.3940 33.2370 ;
        RECT 2.2600 32.1435 2.2860 33.2370 ;
        RECT 2.1520 32.1435 2.1780 33.2370 ;
        RECT 2.0440 32.1435 2.0700 33.2370 ;
        RECT 1.9360 32.1435 1.9620 33.2370 ;
        RECT 1.8280 32.1435 1.8540 33.2370 ;
        RECT 1.7200 32.1435 1.7460 33.2370 ;
        RECT 1.6120 32.1435 1.6380 33.2370 ;
        RECT 1.5040 32.1435 1.5300 33.2370 ;
        RECT 1.3960 32.1435 1.4220 33.2370 ;
        RECT 1.2880 32.1435 1.3140 33.2370 ;
        RECT 1.1800 32.1435 1.2060 33.2370 ;
        RECT 1.0720 32.1435 1.0980 33.2370 ;
        RECT 0.9640 32.1435 0.9900 33.2370 ;
        RECT 0.8560 32.1435 0.8820 33.2370 ;
        RECT 0.7480 32.1435 0.7740 33.2370 ;
        RECT 0.6400 32.1435 0.6660 33.2370 ;
        RECT 0.5320 32.1435 0.5580 33.2370 ;
        RECT 0.4240 32.1435 0.4500 33.2370 ;
        RECT 0.3160 32.1435 0.3420 33.2370 ;
        RECT 0.2080 32.1435 0.2340 33.2370 ;
        RECT 0.0050 32.1435 0.0900 33.2370 ;
        RECT 15.5530 33.2235 15.6810 34.3170 ;
        RECT 15.5390 33.8890 15.6810 34.2115 ;
        RECT 15.3190 33.6160 15.4530 34.3170 ;
        RECT 15.2960 33.9510 15.4530 34.2090 ;
        RECT 15.3190 33.2235 15.4170 34.3170 ;
        RECT 15.3190 33.3445 15.4310 33.5840 ;
        RECT 15.3190 33.2235 15.4530 33.3125 ;
        RECT 15.0940 33.6740 15.2280 34.3170 ;
        RECT 15.0940 33.2235 15.1920 34.3170 ;
        RECT 14.6770 33.2235 14.7600 34.3170 ;
        RECT 14.6770 33.3120 14.7740 34.2475 ;
        RECT 30.2680 33.2235 30.3530 34.3170 ;
        RECT 30.1240 33.2235 30.1500 34.3170 ;
        RECT 30.0160 33.2235 30.0420 34.3170 ;
        RECT 29.9080 33.2235 29.9340 34.3170 ;
        RECT 29.8000 33.2235 29.8260 34.3170 ;
        RECT 29.6920 33.2235 29.7180 34.3170 ;
        RECT 29.5840 33.2235 29.6100 34.3170 ;
        RECT 29.4760 33.2235 29.5020 34.3170 ;
        RECT 29.3680 33.2235 29.3940 34.3170 ;
        RECT 29.2600 33.2235 29.2860 34.3170 ;
        RECT 29.1520 33.2235 29.1780 34.3170 ;
        RECT 29.0440 33.2235 29.0700 34.3170 ;
        RECT 28.9360 33.2235 28.9620 34.3170 ;
        RECT 28.8280 33.2235 28.8540 34.3170 ;
        RECT 28.7200 33.2235 28.7460 34.3170 ;
        RECT 28.6120 33.2235 28.6380 34.3170 ;
        RECT 28.5040 33.2235 28.5300 34.3170 ;
        RECT 28.3960 33.2235 28.4220 34.3170 ;
        RECT 28.2880 33.2235 28.3140 34.3170 ;
        RECT 28.1800 33.2235 28.2060 34.3170 ;
        RECT 28.0720 33.2235 28.0980 34.3170 ;
        RECT 27.9640 33.2235 27.9900 34.3170 ;
        RECT 27.8560 33.2235 27.8820 34.3170 ;
        RECT 27.7480 33.2235 27.7740 34.3170 ;
        RECT 27.6400 33.2235 27.6660 34.3170 ;
        RECT 27.5320 33.2235 27.5580 34.3170 ;
        RECT 27.4240 33.2235 27.4500 34.3170 ;
        RECT 27.3160 33.2235 27.3420 34.3170 ;
        RECT 27.2080 33.2235 27.2340 34.3170 ;
        RECT 27.1000 33.2235 27.1260 34.3170 ;
        RECT 26.9920 33.2235 27.0180 34.3170 ;
        RECT 26.8840 33.2235 26.9100 34.3170 ;
        RECT 26.7760 33.2235 26.8020 34.3170 ;
        RECT 26.6680 33.2235 26.6940 34.3170 ;
        RECT 26.5600 33.2235 26.5860 34.3170 ;
        RECT 26.4520 33.2235 26.4780 34.3170 ;
        RECT 26.3440 33.2235 26.3700 34.3170 ;
        RECT 26.2360 33.2235 26.2620 34.3170 ;
        RECT 26.1280 33.2235 26.1540 34.3170 ;
        RECT 26.0200 33.2235 26.0460 34.3170 ;
        RECT 25.9120 33.2235 25.9380 34.3170 ;
        RECT 25.8040 33.2235 25.8300 34.3170 ;
        RECT 25.6960 33.2235 25.7220 34.3170 ;
        RECT 25.5880 33.2235 25.6140 34.3170 ;
        RECT 25.4800 33.2235 25.5060 34.3170 ;
        RECT 25.3720 33.2235 25.3980 34.3170 ;
        RECT 25.2640 33.2235 25.2900 34.3170 ;
        RECT 25.1560 33.2235 25.1820 34.3170 ;
        RECT 25.0480 33.2235 25.0740 34.3170 ;
        RECT 24.9400 33.2235 24.9660 34.3170 ;
        RECT 24.8320 33.2235 24.8580 34.3170 ;
        RECT 24.7240 33.2235 24.7500 34.3170 ;
        RECT 24.6160 33.2235 24.6420 34.3170 ;
        RECT 24.5080 33.2235 24.5340 34.3170 ;
        RECT 24.4000 33.2235 24.4260 34.3170 ;
        RECT 24.2920 33.2235 24.3180 34.3170 ;
        RECT 24.1840 33.2235 24.2100 34.3170 ;
        RECT 24.0760 33.2235 24.1020 34.3170 ;
        RECT 23.9680 33.2235 23.9940 34.3170 ;
        RECT 23.8600 33.2235 23.8860 34.3170 ;
        RECT 23.7520 33.2235 23.7780 34.3170 ;
        RECT 23.6440 33.2235 23.6700 34.3170 ;
        RECT 23.5360 33.2235 23.5620 34.3170 ;
        RECT 23.4280 33.2235 23.4540 34.3170 ;
        RECT 23.3200 33.2235 23.3460 34.3170 ;
        RECT 23.2120 33.2235 23.2380 34.3170 ;
        RECT 23.1040 33.2235 23.1300 34.3170 ;
        RECT 22.9960 33.2235 23.0220 34.3170 ;
        RECT 22.8880 33.2235 22.9140 34.3170 ;
        RECT 22.7800 33.2235 22.8060 34.3170 ;
        RECT 22.6720 33.2235 22.6980 34.3170 ;
        RECT 22.5640 33.2235 22.5900 34.3170 ;
        RECT 22.4560 33.2235 22.4820 34.3170 ;
        RECT 22.3480 33.2235 22.3740 34.3170 ;
        RECT 22.2400 33.2235 22.2660 34.3170 ;
        RECT 22.1320 33.2235 22.1580 34.3170 ;
        RECT 22.0240 33.2235 22.0500 34.3170 ;
        RECT 21.9160 33.2235 21.9420 34.3170 ;
        RECT 21.8080 33.2235 21.8340 34.3170 ;
        RECT 21.7000 33.2235 21.7260 34.3170 ;
        RECT 21.5920 33.2235 21.6180 34.3170 ;
        RECT 21.4840 33.2235 21.5100 34.3170 ;
        RECT 21.3760 33.2235 21.4020 34.3170 ;
        RECT 21.2680 33.2235 21.2940 34.3170 ;
        RECT 21.1600 33.2235 21.1860 34.3170 ;
        RECT 21.0520 33.2235 21.0780 34.3170 ;
        RECT 20.9440 33.2235 20.9700 34.3170 ;
        RECT 20.8360 33.2235 20.8620 34.3170 ;
        RECT 20.7280 33.2235 20.7540 34.3170 ;
        RECT 20.6200 33.2235 20.6460 34.3170 ;
        RECT 20.5120 33.2235 20.5380 34.3170 ;
        RECT 20.4040 33.2235 20.4300 34.3170 ;
        RECT 20.2960 33.2235 20.3220 34.3170 ;
        RECT 20.1880 33.2235 20.2140 34.3170 ;
        RECT 20.0800 33.2235 20.1060 34.3170 ;
        RECT 19.9720 33.2235 19.9980 34.3170 ;
        RECT 19.8640 33.2235 19.8900 34.3170 ;
        RECT 19.7560 33.2235 19.7820 34.3170 ;
        RECT 19.6480 33.2235 19.6740 34.3170 ;
        RECT 19.5400 33.2235 19.5660 34.3170 ;
        RECT 19.4320 33.2235 19.4580 34.3170 ;
        RECT 19.3240 33.2235 19.3500 34.3170 ;
        RECT 19.2160 33.2235 19.2420 34.3170 ;
        RECT 19.1080 33.2235 19.1340 34.3170 ;
        RECT 19.0000 33.2235 19.0260 34.3170 ;
        RECT 18.8920 33.2235 18.9180 34.3170 ;
        RECT 18.7840 33.2235 18.8100 34.3170 ;
        RECT 18.6760 33.2235 18.7020 34.3170 ;
        RECT 18.5680 33.2235 18.5940 34.3170 ;
        RECT 18.4600 33.2235 18.4860 34.3170 ;
        RECT 18.3520 33.2235 18.3780 34.3170 ;
        RECT 18.2440 33.2235 18.2700 34.3170 ;
        RECT 18.1360 33.2235 18.1620 34.3170 ;
        RECT 18.0280 33.2235 18.0540 34.3170 ;
        RECT 17.9200 33.2235 17.9460 34.3170 ;
        RECT 17.8120 33.2235 17.8380 34.3170 ;
        RECT 17.7040 33.2235 17.7300 34.3170 ;
        RECT 17.5960 33.2235 17.6220 34.3170 ;
        RECT 17.4880 33.2235 17.5140 34.3170 ;
        RECT 17.3800 33.2235 17.4060 34.3170 ;
        RECT 17.2720 33.2235 17.2980 34.3170 ;
        RECT 17.1640 33.2235 17.1900 34.3170 ;
        RECT 17.0560 33.2235 17.0820 34.3170 ;
        RECT 16.9480 33.2235 16.9740 34.3170 ;
        RECT 16.8400 33.2235 16.8660 34.3170 ;
        RECT 16.7320 33.2235 16.7580 34.3170 ;
        RECT 16.6240 33.2235 16.6500 34.3170 ;
        RECT 16.5160 33.2235 16.5420 34.3170 ;
        RECT 16.4080 33.2235 16.4340 34.3170 ;
        RECT 16.3000 33.2235 16.3260 34.3170 ;
        RECT 16.0870 33.2235 16.1640 34.3170 ;
        RECT 14.1940 33.2235 14.2710 34.3170 ;
        RECT 14.0320 33.2235 14.0580 34.3170 ;
        RECT 13.9240 33.2235 13.9500 34.3170 ;
        RECT 13.8160 33.2235 13.8420 34.3170 ;
        RECT 13.7080 33.2235 13.7340 34.3170 ;
        RECT 13.6000 33.2235 13.6260 34.3170 ;
        RECT 13.4920 33.2235 13.5180 34.3170 ;
        RECT 13.3840 33.2235 13.4100 34.3170 ;
        RECT 13.2760 33.2235 13.3020 34.3170 ;
        RECT 13.1680 33.2235 13.1940 34.3170 ;
        RECT 13.0600 33.2235 13.0860 34.3170 ;
        RECT 12.9520 33.2235 12.9780 34.3170 ;
        RECT 12.8440 33.2235 12.8700 34.3170 ;
        RECT 12.7360 33.2235 12.7620 34.3170 ;
        RECT 12.6280 33.2235 12.6540 34.3170 ;
        RECT 12.5200 33.2235 12.5460 34.3170 ;
        RECT 12.4120 33.2235 12.4380 34.3170 ;
        RECT 12.3040 33.2235 12.3300 34.3170 ;
        RECT 12.1960 33.2235 12.2220 34.3170 ;
        RECT 12.0880 33.2235 12.1140 34.3170 ;
        RECT 11.9800 33.2235 12.0060 34.3170 ;
        RECT 11.8720 33.2235 11.8980 34.3170 ;
        RECT 11.7640 33.2235 11.7900 34.3170 ;
        RECT 11.6560 33.2235 11.6820 34.3170 ;
        RECT 11.5480 33.2235 11.5740 34.3170 ;
        RECT 11.4400 33.2235 11.4660 34.3170 ;
        RECT 11.3320 33.2235 11.3580 34.3170 ;
        RECT 11.2240 33.2235 11.2500 34.3170 ;
        RECT 11.1160 33.2235 11.1420 34.3170 ;
        RECT 11.0080 33.2235 11.0340 34.3170 ;
        RECT 10.9000 33.2235 10.9260 34.3170 ;
        RECT 10.7920 33.2235 10.8180 34.3170 ;
        RECT 10.6840 33.2235 10.7100 34.3170 ;
        RECT 10.5760 33.2235 10.6020 34.3170 ;
        RECT 10.4680 33.2235 10.4940 34.3170 ;
        RECT 10.3600 33.2235 10.3860 34.3170 ;
        RECT 10.2520 33.2235 10.2780 34.3170 ;
        RECT 10.1440 33.2235 10.1700 34.3170 ;
        RECT 10.0360 33.2235 10.0620 34.3170 ;
        RECT 9.9280 33.2235 9.9540 34.3170 ;
        RECT 9.8200 33.2235 9.8460 34.3170 ;
        RECT 9.7120 33.2235 9.7380 34.3170 ;
        RECT 9.6040 33.2235 9.6300 34.3170 ;
        RECT 9.4960 33.2235 9.5220 34.3170 ;
        RECT 9.3880 33.2235 9.4140 34.3170 ;
        RECT 9.2800 33.2235 9.3060 34.3170 ;
        RECT 9.1720 33.2235 9.1980 34.3170 ;
        RECT 9.0640 33.2235 9.0900 34.3170 ;
        RECT 8.9560 33.2235 8.9820 34.3170 ;
        RECT 8.8480 33.2235 8.8740 34.3170 ;
        RECT 8.7400 33.2235 8.7660 34.3170 ;
        RECT 8.6320 33.2235 8.6580 34.3170 ;
        RECT 8.5240 33.2235 8.5500 34.3170 ;
        RECT 8.4160 33.2235 8.4420 34.3170 ;
        RECT 8.3080 33.2235 8.3340 34.3170 ;
        RECT 8.2000 33.2235 8.2260 34.3170 ;
        RECT 8.0920 33.2235 8.1180 34.3170 ;
        RECT 7.9840 33.2235 8.0100 34.3170 ;
        RECT 7.8760 33.2235 7.9020 34.3170 ;
        RECT 7.7680 33.2235 7.7940 34.3170 ;
        RECT 7.6600 33.2235 7.6860 34.3170 ;
        RECT 7.5520 33.2235 7.5780 34.3170 ;
        RECT 7.4440 33.2235 7.4700 34.3170 ;
        RECT 7.3360 33.2235 7.3620 34.3170 ;
        RECT 7.2280 33.2235 7.2540 34.3170 ;
        RECT 7.1200 33.2235 7.1460 34.3170 ;
        RECT 7.0120 33.2235 7.0380 34.3170 ;
        RECT 6.9040 33.2235 6.9300 34.3170 ;
        RECT 6.7960 33.2235 6.8220 34.3170 ;
        RECT 6.6880 33.2235 6.7140 34.3170 ;
        RECT 6.5800 33.2235 6.6060 34.3170 ;
        RECT 6.4720 33.2235 6.4980 34.3170 ;
        RECT 6.3640 33.2235 6.3900 34.3170 ;
        RECT 6.2560 33.2235 6.2820 34.3170 ;
        RECT 6.1480 33.2235 6.1740 34.3170 ;
        RECT 6.0400 33.2235 6.0660 34.3170 ;
        RECT 5.9320 33.2235 5.9580 34.3170 ;
        RECT 5.8240 33.2235 5.8500 34.3170 ;
        RECT 5.7160 33.2235 5.7420 34.3170 ;
        RECT 5.6080 33.2235 5.6340 34.3170 ;
        RECT 5.5000 33.2235 5.5260 34.3170 ;
        RECT 5.3920 33.2235 5.4180 34.3170 ;
        RECT 5.2840 33.2235 5.3100 34.3170 ;
        RECT 5.1760 33.2235 5.2020 34.3170 ;
        RECT 5.0680 33.2235 5.0940 34.3170 ;
        RECT 4.9600 33.2235 4.9860 34.3170 ;
        RECT 4.8520 33.2235 4.8780 34.3170 ;
        RECT 4.7440 33.2235 4.7700 34.3170 ;
        RECT 4.6360 33.2235 4.6620 34.3170 ;
        RECT 4.5280 33.2235 4.5540 34.3170 ;
        RECT 4.4200 33.2235 4.4460 34.3170 ;
        RECT 4.3120 33.2235 4.3380 34.3170 ;
        RECT 4.2040 33.2235 4.2300 34.3170 ;
        RECT 4.0960 33.2235 4.1220 34.3170 ;
        RECT 3.9880 33.2235 4.0140 34.3170 ;
        RECT 3.8800 33.2235 3.9060 34.3170 ;
        RECT 3.7720 33.2235 3.7980 34.3170 ;
        RECT 3.6640 33.2235 3.6900 34.3170 ;
        RECT 3.5560 33.2235 3.5820 34.3170 ;
        RECT 3.4480 33.2235 3.4740 34.3170 ;
        RECT 3.3400 33.2235 3.3660 34.3170 ;
        RECT 3.2320 33.2235 3.2580 34.3170 ;
        RECT 3.1240 33.2235 3.1500 34.3170 ;
        RECT 3.0160 33.2235 3.0420 34.3170 ;
        RECT 2.9080 33.2235 2.9340 34.3170 ;
        RECT 2.8000 33.2235 2.8260 34.3170 ;
        RECT 2.6920 33.2235 2.7180 34.3170 ;
        RECT 2.5840 33.2235 2.6100 34.3170 ;
        RECT 2.4760 33.2235 2.5020 34.3170 ;
        RECT 2.3680 33.2235 2.3940 34.3170 ;
        RECT 2.2600 33.2235 2.2860 34.3170 ;
        RECT 2.1520 33.2235 2.1780 34.3170 ;
        RECT 2.0440 33.2235 2.0700 34.3170 ;
        RECT 1.9360 33.2235 1.9620 34.3170 ;
        RECT 1.8280 33.2235 1.8540 34.3170 ;
        RECT 1.7200 33.2235 1.7460 34.3170 ;
        RECT 1.6120 33.2235 1.6380 34.3170 ;
        RECT 1.5040 33.2235 1.5300 34.3170 ;
        RECT 1.3960 33.2235 1.4220 34.3170 ;
        RECT 1.2880 33.2235 1.3140 34.3170 ;
        RECT 1.1800 33.2235 1.2060 34.3170 ;
        RECT 1.0720 33.2235 1.0980 34.3170 ;
        RECT 0.9640 33.2235 0.9900 34.3170 ;
        RECT 0.8560 33.2235 0.8820 34.3170 ;
        RECT 0.7480 33.2235 0.7740 34.3170 ;
        RECT 0.6400 33.2235 0.6660 34.3170 ;
        RECT 0.5320 33.2235 0.5580 34.3170 ;
        RECT 0.4240 33.2235 0.4500 34.3170 ;
        RECT 0.3160 33.2235 0.3420 34.3170 ;
        RECT 0.2080 33.2235 0.2340 34.3170 ;
        RECT 0.0050 33.2235 0.0900 34.3170 ;
        RECT 15.5530 34.3035 15.6810 35.3970 ;
        RECT 15.5390 34.9690 15.6810 35.2915 ;
        RECT 15.3190 34.6960 15.4530 35.3970 ;
        RECT 15.2960 35.0310 15.4530 35.2890 ;
        RECT 15.3190 34.3035 15.4170 35.3970 ;
        RECT 15.3190 34.4245 15.4310 34.6640 ;
        RECT 15.3190 34.3035 15.4530 34.3925 ;
        RECT 15.0940 34.7540 15.2280 35.3970 ;
        RECT 15.0940 34.3035 15.1920 35.3970 ;
        RECT 14.6770 34.3035 14.7600 35.3970 ;
        RECT 14.6770 34.3920 14.7740 35.3275 ;
        RECT 30.2680 34.3035 30.3530 35.3970 ;
        RECT 30.1240 34.3035 30.1500 35.3970 ;
        RECT 30.0160 34.3035 30.0420 35.3970 ;
        RECT 29.9080 34.3035 29.9340 35.3970 ;
        RECT 29.8000 34.3035 29.8260 35.3970 ;
        RECT 29.6920 34.3035 29.7180 35.3970 ;
        RECT 29.5840 34.3035 29.6100 35.3970 ;
        RECT 29.4760 34.3035 29.5020 35.3970 ;
        RECT 29.3680 34.3035 29.3940 35.3970 ;
        RECT 29.2600 34.3035 29.2860 35.3970 ;
        RECT 29.1520 34.3035 29.1780 35.3970 ;
        RECT 29.0440 34.3035 29.0700 35.3970 ;
        RECT 28.9360 34.3035 28.9620 35.3970 ;
        RECT 28.8280 34.3035 28.8540 35.3970 ;
        RECT 28.7200 34.3035 28.7460 35.3970 ;
        RECT 28.6120 34.3035 28.6380 35.3970 ;
        RECT 28.5040 34.3035 28.5300 35.3970 ;
        RECT 28.3960 34.3035 28.4220 35.3970 ;
        RECT 28.2880 34.3035 28.3140 35.3970 ;
        RECT 28.1800 34.3035 28.2060 35.3970 ;
        RECT 28.0720 34.3035 28.0980 35.3970 ;
        RECT 27.9640 34.3035 27.9900 35.3970 ;
        RECT 27.8560 34.3035 27.8820 35.3970 ;
        RECT 27.7480 34.3035 27.7740 35.3970 ;
        RECT 27.6400 34.3035 27.6660 35.3970 ;
        RECT 27.5320 34.3035 27.5580 35.3970 ;
        RECT 27.4240 34.3035 27.4500 35.3970 ;
        RECT 27.3160 34.3035 27.3420 35.3970 ;
        RECT 27.2080 34.3035 27.2340 35.3970 ;
        RECT 27.1000 34.3035 27.1260 35.3970 ;
        RECT 26.9920 34.3035 27.0180 35.3970 ;
        RECT 26.8840 34.3035 26.9100 35.3970 ;
        RECT 26.7760 34.3035 26.8020 35.3970 ;
        RECT 26.6680 34.3035 26.6940 35.3970 ;
        RECT 26.5600 34.3035 26.5860 35.3970 ;
        RECT 26.4520 34.3035 26.4780 35.3970 ;
        RECT 26.3440 34.3035 26.3700 35.3970 ;
        RECT 26.2360 34.3035 26.2620 35.3970 ;
        RECT 26.1280 34.3035 26.1540 35.3970 ;
        RECT 26.0200 34.3035 26.0460 35.3970 ;
        RECT 25.9120 34.3035 25.9380 35.3970 ;
        RECT 25.8040 34.3035 25.8300 35.3970 ;
        RECT 25.6960 34.3035 25.7220 35.3970 ;
        RECT 25.5880 34.3035 25.6140 35.3970 ;
        RECT 25.4800 34.3035 25.5060 35.3970 ;
        RECT 25.3720 34.3035 25.3980 35.3970 ;
        RECT 25.2640 34.3035 25.2900 35.3970 ;
        RECT 25.1560 34.3035 25.1820 35.3970 ;
        RECT 25.0480 34.3035 25.0740 35.3970 ;
        RECT 24.9400 34.3035 24.9660 35.3970 ;
        RECT 24.8320 34.3035 24.8580 35.3970 ;
        RECT 24.7240 34.3035 24.7500 35.3970 ;
        RECT 24.6160 34.3035 24.6420 35.3970 ;
        RECT 24.5080 34.3035 24.5340 35.3970 ;
        RECT 24.4000 34.3035 24.4260 35.3970 ;
        RECT 24.2920 34.3035 24.3180 35.3970 ;
        RECT 24.1840 34.3035 24.2100 35.3970 ;
        RECT 24.0760 34.3035 24.1020 35.3970 ;
        RECT 23.9680 34.3035 23.9940 35.3970 ;
        RECT 23.8600 34.3035 23.8860 35.3970 ;
        RECT 23.7520 34.3035 23.7780 35.3970 ;
        RECT 23.6440 34.3035 23.6700 35.3970 ;
        RECT 23.5360 34.3035 23.5620 35.3970 ;
        RECT 23.4280 34.3035 23.4540 35.3970 ;
        RECT 23.3200 34.3035 23.3460 35.3970 ;
        RECT 23.2120 34.3035 23.2380 35.3970 ;
        RECT 23.1040 34.3035 23.1300 35.3970 ;
        RECT 22.9960 34.3035 23.0220 35.3970 ;
        RECT 22.8880 34.3035 22.9140 35.3970 ;
        RECT 22.7800 34.3035 22.8060 35.3970 ;
        RECT 22.6720 34.3035 22.6980 35.3970 ;
        RECT 22.5640 34.3035 22.5900 35.3970 ;
        RECT 22.4560 34.3035 22.4820 35.3970 ;
        RECT 22.3480 34.3035 22.3740 35.3970 ;
        RECT 22.2400 34.3035 22.2660 35.3970 ;
        RECT 22.1320 34.3035 22.1580 35.3970 ;
        RECT 22.0240 34.3035 22.0500 35.3970 ;
        RECT 21.9160 34.3035 21.9420 35.3970 ;
        RECT 21.8080 34.3035 21.8340 35.3970 ;
        RECT 21.7000 34.3035 21.7260 35.3970 ;
        RECT 21.5920 34.3035 21.6180 35.3970 ;
        RECT 21.4840 34.3035 21.5100 35.3970 ;
        RECT 21.3760 34.3035 21.4020 35.3970 ;
        RECT 21.2680 34.3035 21.2940 35.3970 ;
        RECT 21.1600 34.3035 21.1860 35.3970 ;
        RECT 21.0520 34.3035 21.0780 35.3970 ;
        RECT 20.9440 34.3035 20.9700 35.3970 ;
        RECT 20.8360 34.3035 20.8620 35.3970 ;
        RECT 20.7280 34.3035 20.7540 35.3970 ;
        RECT 20.6200 34.3035 20.6460 35.3970 ;
        RECT 20.5120 34.3035 20.5380 35.3970 ;
        RECT 20.4040 34.3035 20.4300 35.3970 ;
        RECT 20.2960 34.3035 20.3220 35.3970 ;
        RECT 20.1880 34.3035 20.2140 35.3970 ;
        RECT 20.0800 34.3035 20.1060 35.3970 ;
        RECT 19.9720 34.3035 19.9980 35.3970 ;
        RECT 19.8640 34.3035 19.8900 35.3970 ;
        RECT 19.7560 34.3035 19.7820 35.3970 ;
        RECT 19.6480 34.3035 19.6740 35.3970 ;
        RECT 19.5400 34.3035 19.5660 35.3970 ;
        RECT 19.4320 34.3035 19.4580 35.3970 ;
        RECT 19.3240 34.3035 19.3500 35.3970 ;
        RECT 19.2160 34.3035 19.2420 35.3970 ;
        RECT 19.1080 34.3035 19.1340 35.3970 ;
        RECT 19.0000 34.3035 19.0260 35.3970 ;
        RECT 18.8920 34.3035 18.9180 35.3970 ;
        RECT 18.7840 34.3035 18.8100 35.3970 ;
        RECT 18.6760 34.3035 18.7020 35.3970 ;
        RECT 18.5680 34.3035 18.5940 35.3970 ;
        RECT 18.4600 34.3035 18.4860 35.3970 ;
        RECT 18.3520 34.3035 18.3780 35.3970 ;
        RECT 18.2440 34.3035 18.2700 35.3970 ;
        RECT 18.1360 34.3035 18.1620 35.3970 ;
        RECT 18.0280 34.3035 18.0540 35.3970 ;
        RECT 17.9200 34.3035 17.9460 35.3970 ;
        RECT 17.8120 34.3035 17.8380 35.3970 ;
        RECT 17.7040 34.3035 17.7300 35.3970 ;
        RECT 17.5960 34.3035 17.6220 35.3970 ;
        RECT 17.4880 34.3035 17.5140 35.3970 ;
        RECT 17.3800 34.3035 17.4060 35.3970 ;
        RECT 17.2720 34.3035 17.2980 35.3970 ;
        RECT 17.1640 34.3035 17.1900 35.3970 ;
        RECT 17.0560 34.3035 17.0820 35.3970 ;
        RECT 16.9480 34.3035 16.9740 35.3970 ;
        RECT 16.8400 34.3035 16.8660 35.3970 ;
        RECT 16.7320 34.3035 16.7580 35.3970 ;
        RECT 16.6240 34.3035 16.6500 35.3970 ;
        RECT 16.5160 34.3035 16.5420 35.3970 ;
        RECT 16.4080 34.3035 16.4340 35.3970 ;
        RECT 16.3000 34.3035 16.3260 35.3970 ;
        RECT 16.0870 34.3035 16.1640 35.3970 ;
        RECT 14.1940 34.3035 14.2710 35.3970 ;
        RECT 14.0320 34.3035 14.0580 35.3970 ;
        RECT 13.9240 34.3035 13.9500 35.3970 ;
        RECT 13.8160 34.3035 13.8420 35.3970 ;
        RECT 13.7080 34.3035 13.7340 35.3970 ;
        RECT 13.6000 34.3035 13.6260 35.3970 ;
        RECT 13.4920 34.3035 13.5180 35.3970 ;
        RECT 13.3840 34.3035 13.4100 35.3970 ;
        RECT 13.2760 34.3035 13.3020 35.3970 ;
        RECT 13.1680 34.3035 13.1940 35.3970 ;
        RECT 13.0600 34.3035 13.0860 35.3970 ;
        RECT 12.9520 34.3035 12.9780 35.3970 ;
        RECT 12.8440 34.3035 12.8700 35.3970 ;
        RECT 12.7360 34.3035 12.7620 35.3970 ;
        RECT 12.6280 34.3035 12.6540 35.3970 ;
        RECT 12.5200 34.3035 12.5460 35.3970 ;
        RECT 12.4120 34.3035 12.4380 35.3970 ;
        RECT 12.3040 34.3035 12.3300 35.3970 ;
        RECT 12.1960 34.3035 12.2220 35.3970 ;
        RECT 12.0880 34.3035 12.1140 35.3970 ;
        RECT 11.9800 34.3035 12.0060 35.3970 ;
        RECT 11.8720 34.3035 11.8980 35.3970 ;
        RECT 11.7640 34.3035 11.7900 35.3970 ;
        RECT 11.6560 34.3035 11.6820 35.3970 ;
        RECT 11.5480 34.3035 11.5740 35.3970 ;
        RECT 11.4400 34.3035 11.4660 35.3970 ;
        RECT 11.3320 34.3035 11.3580 35.3970 ;
        RECT 11.2240 34.3035 11.2500 35.3970 ;
        RECT 11.1160 34.3035 11.1420 35.3970 ;
        RECT 11.0080 34.3035 11.0340 35.3970 ;
        RECT 10.9000 34.3035 10.9260 35.3970 ;
        RECT 10.7920 34.3035 10.8180 35.3970 ;
        RECT 10.6840 34.3035 10.7100 35.3970 ;
        RECT 10.5760 34.3035 10.6020 35.3970 ;
        RECT 10.4680 34.3035 10.4940 35.3970 ;
        RECT 10.3600 34.3035 10.3860 35.3970 ;
        RECT 10.2520 34.3035 10.2780 35.3970 ;
        RECT 10.1440 34.3035 10.1700 35.3970 ;
        RECT 10.0360 34.3035 10.0620 35.3970 ;
        RECT 9.9280 34.3035 9.9540 35.3970 ;
        RECT 9.8200 34.3035 9.8460 35.3970 ;
        RECT 9.7120 34.3035 9.7380 35.3970 ;
        RECT 9.6040 34.3035 9.6300 35.3970 ;
        RECT 9.4960 34.3035 9.5220 35.3970 ;
        RECT 9.3880 34.3035 9.4140 35.3970 ;
        RECT 9.2800 34.3035 9.3060 35.3970 ;
        RECT 9.1720 34.3035 9.1980 35.3970 ;
        RECT 9.0640 34.3035 9.0900 35.3970 ;
        RECT 8.9560 34.3035 8.9820 35.3970 ;
        RECT 8.8480 34.3035 8.8740 35.3970 ;
        RECT 8.7400 34.3035 8.7660 35.3970 ;
        RECT 8.6320 34.3035 8.6580 35.3970 ;
        RECT 8.5240 34.3035 8.5500 35.3970 ;
        RECT 8.4160 34.3035 8.4420 35.3970 ;
        RECT 8.3080 34.3035 8.3340 35.3970 ;
        RECT 8.2000 34.3035 8.2260 35.3970 ;
        RECT 8.0920 34.3035 8.1180 35.3970 ;
        RECT 7.9840 34.3035 8.0100 35.3970 ;
        RECT 7.8760 34.3035 7.9020 35.3970 ;
        RECT 7.7680 34.3035 7.7940 35.3970 ;
        RECT 7.6600 34.3035 7.6860 35.3970 ;
        RECT 7.5520 34.3035 7.5780 35.3970 ;
        RECT 7.4440 34.3035 7.4700 35.3970 ;
        RECT 7.3360 34.3035 7.3620 35.3970 ;
        RECT 7.2280 34.3035 7.2540 35.3970 ;
        RECT 7.1200 34.3035 7.1460 35.3970 ;
        RECT 7.0120 34.3035 7.0380 35.3970 ;
        RECT 6.9040 34.3035 6.9300 35.3970 ;
        RECT 6.7960 34.3035 6.8220 35.3970 ;
        RECT 6.6880 34.3035 6.7140 35.3970 ;
        RECT 6.5800 34.3035 6.6060 35.3970 ;
        RECT 6.4720 34.3035 6.4980 35.3970 ;
        RECT 6.3640 34.3035 6.3900 35.3970 ;
        RECT 6.2560 34.3035 6.2820 35.3970 ;
        RECT 6.1480 34.3035 6.1740 35.3970 ;
        RECT 6.0400 34.3035 6.0660 35.3970 ;
        RECT 5.9320 34.3035 5.9580 35.3970 ;
        RECT 5.8240 34.3035 5.8500 35.3970 ;
        RECT 5.7160 34.3035 5.7420 35.3970 ;
        RECT 5.6080 34.3035 5.6340 35.3970 ;
        RECT 5.5000 34.3035 5.5260 35.3970 ;
        RECT 5.3920 34.3035 5.4180 35.3970 ;
        RECT 5.2840 34.3035 5.3100 35.3970 ;
        RECT 5.1760 34.3035 5.2020 35.3970 ;
        RECT 5.0680 34.3035 5.0940 35.3970 ;
        RECT 4.9600 34.3035 4.9860 35.3970 ;
        RECT 4.8520 34.3035 4.8780 35.3970 ;
        RECT 4.7440 34.3035 4.7700 35.3970 ;
        RECT 4.6360 34.3035 4.6620 35.3970 ;
        RECT 4.5280 34.3035 4.5540 35.3970 ;
        RECT 4.4200 34.3035 4.4460 35.3970 ;
        RECT 4.3120 34.3035 4.3380 35.3970 ;
        RECT 4.2040 34.3035 4.2300 35.3970 ;
        RECT 4.0960 34.3035 4.1220 35.3970 ;
        RECT 3.9880 34.3035 4.0140 35.3970 ;
        RECT 3.8800 34.3035 3.9060 35.3970 ;
        RECT 3.7720 34.3035 3.7980 35.3970 ;
        RECT 3.6640 34.3035 3.6900 35.3970 ;
        RECT 3.5560 34.3035 3.5820 35.3970 ;
        RECT 3.4480 34.3035 3.4740 35.3970 ;
        RECT 3.3400 34.3035 3.3660 35.3970 ;
        RECT 3.2320 34.3035 3.2580 35.3970 ;
        RECT 3.1240 34.3035 3.1500 35.3970 ;
        RECT 3.0160 34.3035 3.0420 35.3970 ;
        RECT 2.9080 34.3035 2.9340 35.3970 ;
        RECT 2.8000 34.3035 2.8260 35.3970 ;
        RECT 2.6920 34.3035 2.7180 35.3970 ;
        RECT 2.5840 34.3035 2.6100 35.3970 ;
        RECT 2.4760 34.3035 2.5020 35.3970 ;
        RECT 2.3680 34.3035 2.3940 35.3970 ;
        RECT 2.2600 34.3035 2.2860 35.3970 ;
        RECT 2.1520 34.3035 2.1780 35.3970 ;
        RECT 2.0440 34.3035 2.0700 35.3970 ;
        RECT 1.9360 34.3035 1.9620 35.3970 ;
        RECT 1.8280 34.3035 1.8540 35.3970 ;
        RECT 1.7200 34.3035 1.7460 35.3970 ;
        RECT 1.6120 34.3035 1.6380 35.3970 ;
        RECT 1.5040 34.3035 1.5300 35.3970 ;
        RECT 1.3960 34.3035 1.4220 35.3970 ;
        RECT 1.2880 34.3035 1.3140 35.3970 ;
        RECT 1.1800 34.3035 1.2060 35.3970 ;
        RECT 1.0720 34.3035 1.0980 35.3970 ;
        RECT 0.9640 34.3035 0.9900 35.3970 ;
        RECT 0.8560 34.3035 0.8820 35.3970 ;
        RECT 0.7480 34.3035 0.7740 35.3970 ;
        RECT 0.6400 34.3035 0.6660 35.3970 ;
        RECT 0.5320 34.3035 0.5580 35.3970 ;
        RECT 0.4240 34.3035 0.4500 35.3970 ;
        RECT 0.3160 34.3035 0.3420 35.3970 ;
        RECT 0.2080 34.3035 0.2340 35.3970 ;
        RECT 0.0050 34.3035 0.0900 35.3970 ;
        RECT 15.5530 35.3835 15.6810 36.4770 ;
        RECT 15.5390 36.0490 15.6810 36.3715 ;
        RECT 15.3190 35.7760 15.4530 36.4770 ;
        RECT 15.2960 36.1110 15.4530 36.3690 ;
        RECT 15.3190 35.3835 15.4170 36.4770 ;
        RECT 15.3190 35.5045 15.4310 35.7440 ;
        RECT 15.3190 35.3835 15.4530 35.4725 ;
        RECT 15.0940 35.8340 15.2280 36.4770 ;
        RECT 15.0940 35.3835 15.1920 36.4770 ;
        RECT 14.6770 35.3835 14.7600 36.4770 ;
        RECT 14.6770 35.4720 14.7740 36.4075 ;
        RECT 30.2680 35.3835 30.3530 36.4770 ;
        RECT 30.1240 35.3835 30.1500 36.4770 ;
        RECT 30.0160 35.3835 30.0420 36.4770 ;
        RECT 29.9080 35.3835 29.9340 36.4770 ;
        RECT 29.8000 35.3835 29.8260 36.4770 ;
        RECT 29.6920 35.3835 29.7180 36.4770 ;
        RECT 29.5840 35.3835 29.6100 36.4770 ;
        RECT 29.4760 35.3835 29.5020 36.4770 ;
        RECT 29.3680 35.3835 29.3940 36.4770 ;
        RECT 29.2600 35.3835 29.2860 36.4770 ;
        RECT 29.1520 35.3835 29.1780 36.4770 ;
        RECT 29.0440 35.3835 29.0700 36.4770 ;
        RECT 28.9360 35.3835 28.9620 36.4770 ;
        RECT 28.8280 35.3835 28.8540 36.4770 ;
        RECT 28.7200 35.3835 28.7460 36.4770 ;
        RECT 28.6120 35.3835 28.6380 36.4770 ;
        RECT 28.5040 35.3835 28.5300 36.4770 ;
        RECT 28.3960 35.3835 28.4220 36.4770 ;
        RECT 28.2880 35.3835 28.3140 36.4770 ;
        RECT 28.1800 35.3835 28.2060 36.4770 ;
        RECT 28.0720 35.3835 28.0980 36.4770 ;
        RECT 27.9640 35.3835 27.9900 36.4770 ;
        RECT 27.8560 35.3835 27.8820 36.4770 ;
        RECT 27.7480 35.3835 27.7740 36.4770 ;
        RECT 27.6400 35.3835 27.6660 36.4770 ;
        RECT 27.5320 35.3835 27.5580 36.4770 ;
        RECT 27.4240 35.3835 27.4500 36.4770 ;
        RECT 27.3160 35.3835 27.3420 36.4770 ;
        RECT 27.2080 35.3835 27.2340 36.4770 ;
        RECT 27.1000 35.3835 27.1260 36.4770 ;
        RECT 26.9920 35.3835 27.0180 36.4770 ;
        RECT 26.8840 35.3835 26.9100 36.4770 ;
        RECT 26.7760 35.3835 26.8020 36.4770 ;
        RECT 26.6680 35.3835 26.6940 36.4770 ;
        RECT 26.5600 35.3835 26.5860 36.4770 ;
        RECT 26.4520 35.3835 26.4780 36.4770 ;
        RECT 26.3440 35.3835 26.3700 36.4770 ;
        RECT 26.2360 35.3835 26.2620 36.4770 ;
        RECT 26.1280 35.3835 26.1540 36.4770 ;
        RECT 26.0200 35.3835 26.0460 36.4770 ;
        RECT 25.9120 35.3835 25.9380 36.4770 ;
        RECT 25.8040 35.3835 25.8300 36.4770 ;
        RECT 25.6960 35.3835 25.7220 36.4770 ;
        RECT 25.5880 35.3835 25.6140 36.4770 ;
        RECT 25.4800 35.3835 25.5060 36.4770 ;
        RECT 25.3720 35.3835 25.3980 36.4770 ;
        RECT 25.2640 35.3835 25.2900 36.4770 ;
        RECT 25.1560 35.3835 25.1820 36.4770 ;
        RECT 25.0480 35.3835 25.0740 36.4770 ;
        RECT 24.9400 35.3835 24.9660 36.4770 ;
        RECT 24.8320 35.3835 24.8580 36.4770 ;
        RECT 24.7240 35.3835 24.7500 36.4770 ;
        RECT 24.6160 35.3835 24.6420 36.4770 ;
        RECT 24.5080 35.3835 24.5340 36.4770 ;
        RECT 24.4000 35.3835 24.4260 36.4770 ;
        RECT 24.2920 35.3835 24.3180 36.4770 ;
        RECT 24.1840 35.3835 24.2100 36.4770 ;
        RECT 24.0760 35.3835 24.1020 36.4770 ;
        RECT 23.9680 35.3835 23.9940 36.4770 ;
        RECT 23.8600 35.3835 23.8860 36.4770 ;
        RECT 23.7520 35.3835 23.7780 36.4770 ;
        RECT 23.6440 35.3835 23.6700 36.4770 ;
        RECT 23.5360 35.3835 23.5620 36.4770 ;
        RECT 23.4280 35.3835 23.4540 36.4770 ;
        RECT 23.3200 35.3835 23.3460 36.4770 ;
        RECT 23.2120 35.3835 23.2380 36.4770 ;
        RECT 23.1040 35.3835 23.1300 36.4770 ;
        RECT 22.9960 35.3835 23.0220 36.4770 ;
        RECT 22.8880 35.3835 22.9140 36.4770 ;
        RECT 22.7800 35.3835 22.8060 36.4770 ;
        RECT 22.6720 35.3835 22.6980 36.4770 ;
        RECT 22.5640 35.3835 22.5900 36.4770 ;
        RECT 22.4560 35.3835 22.4820 36.4770 ;
        RECT 22.3480 35.3835 22.3740 36.4770 ;
        RECT 22.2400 35.3835 22.2660 36.4770 ;
        RECT 22.1320 35.3835 22.1580 36.4770 ;
        RECT 22.0240 35.3835 22.0500 36.4770 ;
        RECT 21.9160 35.3835 21.9420 36.4770 ;
        RECT 21.8080 35.3835 21.8340 36.4770 ;
        RECT 21.7000 35.3835 21.7260 36.4770 ;
        RECT 21.5920 35.3835 21.6180 36.4770 ;
        RECT 21.4840 35.3835 21.5100 36.4770 ;
        RECT 21.3760 35.3835 21.4020 36.4770 ;
        RECT 21.2680 35.3835 21.2940 36.4770 ;
        RECT 21.1600 35.3835 21.1860 36.4770 ;
        RECT 21.0520 35.3835 21.0780 36.4770 ;
        RECT 20.9440 35.3835 20.9700 36.4770 ;
        RECT 20.8360 35.3835 20.8620 36.4770 ;
        RECT 20.7280 35.3835 20.7540 36.4770 ;
        RECT 20.6200 35.3835 20.6460 36.4770 ;
        RECT 20.5120 35.3835 20.5380 36.4770 ;
        RECT 20.4040 35.3835 20.4300 36.4770 ;
        RECT 20.2960 35.3835 20.3220 36.4770 ;
        RECT 20.1880 35.3835 20.2140 36.4770 ;
        RECT 20.0800 35.3835 20.1060 36.4770 ;
        RECT 19.9720 35.3835 19.9980 36.4770 ;
        RECT 19.8640 35.3835 19.8900 36.4770 ;
        RECT 19.7560 35.3835 19.7820 36.4770 ;
        RECT 19.6480 35.3835 19.6740 36.4770 ;
        RECT 19.5400 35.3835 19.5660 36.4770 ;
        RECT 19.4320 35.3835 19.4580 36.4770 ;
        RECT 19.3240 35.3835 19.3500 36.4770 ;
        RECT 19.2160 35.3835 19.2420 36.4770 ;
        RECT 19.1080 35.3835 19.1340 36.4770 ;
        RECT 19.0000 35.3835 19.0260 36.4770 ;
        RECT 18.8920 35.3835 18.9180 36.4770 ;
        RECT 18.7840 35.3835 18.8100 36.4770 ;
        RECT 18.6760 35.3835 18.7020 36.4770 ;
        RECT 18.5680 35.3835 18.5940 36.4770 ;
        RECT 18.4600 35.3835 18.4860 36.4770 ;
        RECT 18.3520 35.3835 18.3780 36.4770 ;
        RECT 18.2440 35.3835 18.2700 36.4770 ;
        RECT 18.1360 35.3835 18.1620 36.4770 ;
        RECT 18.0280 35.3835 18.0540 36.4770 ;
        RECT 17.9200 35.3835 17.9460 36.4770 ;
        RECT 17.8120 35.3835 17.8380 36.4770 ;
        RECT 17.7040 35.3835 17.7300 36.4770 ;
        RECT 17.5960 35.3835 17.6220 36.4770 ;
        RECT 17.4880 35.3835 17.5140 36.4770 ;
        RECT 17.3800 35.3835 17.4060 36.4770 ;
        RECT 17.2720 35.3835 17.2980 36.4770 ;
        RECT 17.1640 35.3835 17.1900 36.4770 ;
        RECT 17.0560 35.3835 17.0820 36.4770 ;
        RECT 16.9480 35.3835 16.9740 36.4770 ;
        RECT 16.8400 35.3835 16.8660 36.4770 ;
        RECT 16.7320 35.3835 16.7580 36.4770 ;
        RECT 16.6240 35.3835 16.6500 36.4770 ;
        RECT 16.5160 35.3835 16.5420 36.4770 ;
        RECT 16.4080 35.3835 16.4340 36.4770 ;
        RECT 16.3000 35.3835 16.3260 36.4770 ;
        RECT 16.0870 35.3835 16.1640 36.4770 ;
        RECT 14.1940 35.3835 14.2710 36.4770 ;
        RECT 14.0320 35.3835 14.0580 36.4770 ;
        RECT 13.9240 35.3835 13.9500 36.4770 ;
        RECT 13.8160 35.3835 13.8420 36.4770 ;
        RECT 13.7080 35.3835 13.7340 36.4770 ;
        RECT 13.6000 35.3835 13.6260 36.4770 ;
        RECT 13.4920 35.3835 13.5180 36.4770 ;
        RECT 13.3840 35.3835 13.4100 36.4770 ;
        RECT 13.2760 35.3835 13.3020 36.4770 ;
        RECT 13.1680 35.3835 13.1940 36.4770 ;
        RECT 13.0600 35.3835 13.0860 36.4770 ;
        RECT 12.9520 35.3835 12.9780 36.4770 ;
        RECT 12.8440 35.3835 12.8700 36.4770 ;
        RECT 12.7360 35.3835 12.7620 36.4770 ;
        RECT 12.6280 35.3835 12.6540 36.4770 ;
        RECT 12.5200 35.3835 12.5460 36.4770 ;
        RECT 12.4120 35.3835 12.4380 36.4770 ;
        RECT 12.3040 35.3835 12.3300 36.4770 ;
        RECT 12.1960 35.3835 12.2220 36.4770 ;
        RECT 12.0880 35.3835 12.1140 36.4770 ;
        RECT 11.9800 35.3835 12.0060 36.4770 ;
        RECT 11.8720 35.3835 11.8980 36.4770 ;
        RECT 11.7640 35.3835 11.7900 36.4770 ;
        RECT 11.6560 35.3835 11.6820 36.4770 ;
        RECT 11.5480 35.3835 11.5740 36.4770 ;
        RECT 11.4400 35.3835 11.4660 36.4770 ;
        RECT 11.3320 35.3835 11.3580 36.4770 ;
        RECT 11.2240 35.3835 11.2500 36.4770 ;
        RECT 11.1160 35.3835 11.1420 36.4770 ;
        RECT 11.0080 35.3835 11.0340 36.4770 ;
        RECT 10.9000 35.3835 10.9260 36.4770 ;
        RECT 10.7920 35.3835 10.8180 36.4770 ;
        RECT 10.6840 35.3835 10.7100 36.4770 ;
        RECT 10.5760 35.3835 10.6020 36.4770 ;
        RECT 10.4680 35.3835 10.4940 36.4770 ;
        RECT 10.3600 35.3835 10.3860 36.4770 ;
        RECT 10.2520 35.3835 10.2780 36.4770 ;
        RECT 10.1440 35.3835 10.1700 36.4770 ;
        RECT 10.0360 35.3835 10.0620 36.4770 ;
        RECT 9.9280 35.3835 9.9540 36.4770 ;
        RECT 9.8200 35.3835 9.8460 36.4770 ;
        RECT 9.7120 35.3835 9.7380 36.4770 ;
        RECT 9.6040 35.3835 9.6300 36.4770 ;
        RECT 9.4960 35.3835 9.5220 36.4770 ;
        RECT 9.3880 35.3835 9.4140 36.4770 ;
        RECT 9.2800 35.3835 9.3060 36.4770 ;
        RECT 9.1720 35.3835 9.1980 36.4770 ;
        RECT 9.0640 35.3835 9.0900 36.4770 ;
        RECT 8.9560 35.3835 8.9820 36.4770 ;
        RECT 8.8480 35.3835 8.8740 36.4770 ;
        RECT 8.7400 35.3835 8.7660 36.4770 ;
        RECT 8.6320 35.3835 8.6580 36.4770 ;
        RECT 8.5240 35.3835 8.5500 36.4770 ;
        RECT 8.4160 35.3835 8.4420 36.4770 ;
        RECT 8.3080 35.3835 8.3340 36.4770 ;
        RECT 8.2000 35.3835 8.2260 36.4770 ;
        RECT 8.0920 35.3835 8.1180 36.4770 ;
        RECT 7.9840 35.3835 8.0100 36.4770 ;
        RECT 7.8760 35.3835 7.9020 36.4770 ;
        RECT 7.7680 35.3835 7.7940 36.4770 ;
        RECT 7.6600 35.3835 7.6860 36.4770 ;
        RECT 7.5520 35.3835 7.5780 36.4770 ;
        RECT 7.4440 35.3835 7.4700 36.4770 ;
        RECT 7.3360 35.3835 7.3620 36.4770 ;
        RECT 7.2280 35.3835 7.2540 36.4770 ;
        RECT 7.1200 35.3835 7.1460 36.4770 ;
        RECT 7.0120 35.3835 7.0380 36.4770 ;
        RECT 6.9040 35.3835 6.9300 36.4770 ;
        RECT 6.7960 35.3835 6.8220 36.4770 ;
        RECT 6.6880 35.3835 6.7140 36.4770 ;
        RECT 6.5800 35.3835 6.6060 36.4770 ;
        RECT 6.4720 35.3835 6.4980 36.4770 ;
        RECT 6.3640 35.3835 6.3900 36.4770 ;
        RECT 6.2560 35.3835 6.2820 36.4770 ;
        RECT 6.1480 35.3835 6.1740 36.4770 ;
        RECT 6.0400 35.3835 6.0660 36.4770 ;
        RECT 5.9320 35.3835 5.9580 36.4770 ;
        RECT 5.8240 35.3835 5.8500 36.4770 ;
        RECT 5.7160 35.3835 5.7420 36.4770 ;
        RECT 5.6080 35.3835 5.6340 36.4770 ;
        RECT 5.5000 35.3835 5.5260 36.4770 ;
        RECT 5.3920 35.3835 5.4180 36.4770 ;
        RECT 5.2840 35.3835 5.3100 36.4770 ;
        RECT 5.1760 35.3835 5.2020 36.4770 ;
        RECT 5.0680 35.3835 5.0940 36.4770 ;
        RECT 4.9600 35.3835 4.9860 36.4770 ;
        RECT 4.8520 35.3835 4.8780 36.4770 ;
        RECT 4.7440 35.3835 4.7700 36.4770 ;
        RECT 4.6360 35.3835 4.6620 36.4770 ;
        RECT 4.5280 35.3835 4.5540 36.4770 ;
        RECT 4.4200 35.3835 4.4460 36.4770 ;
        RECT 4.3120 35.3835 4.3380 36.4770 ;
        RECT 4.2040 35.3835 4.2300 36.4770 ;
        RECT 4.0960 35.3835 4.1220 36.4770 ;
        RECT 3.9880 35.3835 4.0140 36.4770 ;
        RECT 3.8800 35.3835 3.9060 36.4770 ;
        RECT 3.7720 35.3835 3.7980 36.4770 ;
        RECT 3.6640 35.3835 3.6900 36.4770 ;
        RECT 3.5560 35.3835 3.5820 36.4770 ;
        RECT 3.4480 35.3835 3.4740 36.4770 ;
        RECT 3.3400 35.3835 3.3660 36.4770 ;
        RECT 3.2320 35.3835 3.2580 36.4770 ;
        RECT 3.1240 35.3835 3.1500 36.4770 ;
        RECT 3.0160 35.3835 3.0420 36.4770 ;
        RECT 2.9080 35.3835 2.9340 36.4770 ;
        RECT 2.8000 35.3835 2.8260 36.4770 ;
        RECT 2.6920 35.3835 2.7180 36.4770 ;
        RECT 2.5840 35.3835 2.6100 36.4770 ;
        RECT 2.4760 35.3835 2.5020 36.4770 ;
        RECT 2.3680 35.3835 2.3940 36.4770 ;
        RECT 2.2600 35.3835 2.2860 36.4770 ;
        RECT 2.1520 35.3835 2.1780 36.4770 ;
        RECT 2.0440 35.3835 2.0700 36.4770 ;
        RECT 1.9360 35.3835 1.9620 36.4770 ;
        RECT 1.8280 35.3835 1.8540 36.4770 ;
        RECT 1.7200 35.3835 1.7460 36.4770 ;
        RECT 1.6120 35.3835 1.6380 36.4770 ;
        RECT 1.5040 35.3835 1.5300 36.4770 ;
        RECT 1.3960 35.3835 1.4220 36.4770 ;
        RECT 1.2880 35.3835 1.3140 36.4770 ;
        RECT 1.1800 35.3835 1.2060 36.4770 ;
        RECT 1.0720 35.3835 1.0980 36.4770 ;
        RECT 0.9640 35.3835 0.9900 36.4770 ;
        RECT 0.8560 35.3835 0.8820 36.4770 ;
        RECT 0.7480 35.3835 0.7740 36.4770 ;
        RECT 0.6400 35.3835 0.6660 36.4770 ;
        RECT 0.5320 35.3835 0.5580 36.4770 ;
        RECT 0.4240 35.3835 0.4500 36.4770 ;
        RECT 0.3160 35.3835 0.3420 36.4770 ;
        RECT 0.2080 35.3835 0.2340 36.4770 ;
        RECT 0.0050 35.3835 0.0900 36.4770 ;
        RECT 15.5530 36.4635 15.6810 37.5570 ;
        RECT 15.5390 37.1290 15.6810 37.4515 ;
        RECT 15.3190 36.8560 15.4530 37.5570 ;
        RECT 15.2960 37.1910 15.4530 37.4490 ;
        RECT 15.3190 36.4635 15.4170 37.5570 ;
        RECT 15.3190 36.5845 15.4310 36.8240 ;
        RECT 15.3190 36.4635 15.4530 36.5525 ;
        RECT 15.0940 36.9140 15.2280 37.5570 ;
        RECT 15.0940 36.4635 15.1920 37.5570 ;
        RECT 14.6770 36.4635 14.7600 37.5570 ;
        RECT 14.6770 36.5520 14.7740 37.4875 ;
        RECT 30.2680 36.4635 30.3530 37.5570 ;
        RECT 30.1240 36.4635 30.1500 37.5570 ;
        RECT 30.0160 36.4635 30.0420 37.5570 ;
        RECT 29.9080 36.4635 29.9340 37.5570 ;
        RECT 29.8000 36.4635 29.8260 37.5570 ;
        RECT 29.6920 36.4635 29.7180 37.5570 ;
        RECT 29.5840 36.4635 29.6100 37.5570 ;
        RECT 29.4760 36.4635 29.5020 37.5570 ;
        RECT 29.3680 36.4635 29.3940 37.5570 ;
        RECT 29.2600 36.4635 29.2860 37.5570 ;
        RECT 29.1520 36.4635 29.1780 37.5570 ;
        RECT 29.0440 36.4635 29.0700 37.5570 ;
        RECT 28.9360 36.4635 28.9620 37.5570 ;
        RECT 28.8280 36.4635 28.8540 37.5570 ;
        RECT 28.7200 36.4635 28.7460 37.5570 ;
        RECT 28.6120 36.4635 28.6380 37.5570 ;
        RECT 28.5040 36.4635 28.5300 37.5570 ;
        RECT 28.3960 36.4635 28.4220 37.5570 ;
        RECT 28.2880 36.4635 28.3140 37.5570 ;
        RECT 28.1800 36.4635 28.2060 37.5570 ;
        RECT 28.0720 36.4635 28.0980 37.5570 ;
        RECT 27.9640 36.4635 27.9900 37.5570 ;
        RECT 27.8560 36.4635 27.8820 37.5570 ;
        RECT 27.7480 36.4635 27.7740 37.5570 ;
        RECT 27.6400 36.4635 27.6660 37.5570 ;
        RECT 27.5320 36.4635 27.5580 37.5570 ;
        RECT 27.4240 36.4635 27.4500 37.5570 ;
        RECT 27.3160 36.4635 27.3420 37.5570 ;
        RECT 27.2080 36.4635 27.2340 37.5570 ;
        RECT 27.1000 36.4635 27.1260 37.5570 ;
        RECT 26.9920 36.4635 27.0180 37.5570 ;
        RECT 26.8840 36.4635 26.9100 37.5570 ;
        RECT 26.7760 36.4635 26.8020 37.5570 ;
        RECT 26.6680 36.4635 26.6940 37.5570 ;
        RECT 26.5600 36.4635 26.5860 37.5570 ;
        RECT 26.4520 36.4635 26.4780 37.5570 ;
        RECT 26.3440 36.4635 26.3700 37.5570 ;
        RECT 26.2360 36.4635 26.2620 37.5570 ;
        RECT 26.1280 36.4635 26.1540 37.5570 ;
        RECT 26.0200 36.4635 26.0460 37.5570 ;
        RECT 25.9120 36.4635 25.9380 37.5570 ;
        RECT 25.8040 36.4635 25.8300 37.5570 ;
        RECT 25.6960 36.4635 25.7220 37.5570 ;
        RECT 25.5880 36.4635 25.6140 37.5570 ;
        RECT 25.4800 36.4635 25.5060 37.5570 ;
        RECT 25.3720 36.4635 25.3980 37.5570 ;
        RECT 25.2640 36.4635 25.2900 37.5570 ;
        RECT 25.1560 36.4635 25.1820 37.5570 ;
        RECT 25.0480 36.4635 25.0740 37.5570 ;
        RECT 24.9400 36.4635 24.9660 37.5570 ;
        RECT 24.8320 36.4635 24.8580 37.5570 ;
        RECT 24.7240 36.4635 24.7500 37.5570 ;
        RECT 24.6160 36.4635 24.6420 37.5570 ;
        RECT 24.5080 36.4635 24.5340 37.5570 ;
        RECT 24.4000 36.4635 24.4260 37.5570 ;
        RECT 24.2920 36.4635 24.3180 37.5570 ;
        RECT 24.1840 36.4635 24.2100 37.5570 ;
        RECT 24.0760 36.4635 24.1020 37.5570 ;
        RECT 23.9680 36.4635 23.9940 37.5570 ;
        RECT 23.8600 36.4635 23.8860 37.5570 ;
        RECT 23.7520 36.4635 23.7780 37.5570 ;
        RECT 23.6440 36.4635 23.6700 37.5570 ;
        RECT 23.5360 36.4635 23.5620 37.5570 ;
        RECT 23.4280 36.4635 23.4540 37.5570 ;
        RECT 23.3200 36.4635 23.3460 37.5570 ;
        RECT 23.2120 36.4635 23.2380 37.5570 ;
        RECT 23.1040 36.4635 23.1300 37.5570 ;
        RECT 22.9960 36.4635 23.0220 37.5570 ;
        RECT 22.8880 36.4635 22.9140 37.5570 ;
        RECT 22.7800 36.4635 22.8060 37.5570 ;
        RECT 22.6720 36.4635 22.6980 37.5570 ;
        RECT 22.5640 36.4635 22.5900 37.5570 ;
        RECT 22.4560 36.4635 22.4820 37.5570 ;
        RECT 22.3480 36.4635 22.3740 37.5570 ;
        RECT 22.2400 36.4635 22.2660 37.5570 ;
        RECT 22.1320 36.4635 22.1580 37.5570 ;
        RECT 22.0240 36.4635 22.0500 37.5570 ;
        RECT 21.9160 36.4635 21.9420 37.5570 ;
        RECT 21.8080 36.4635 21.8340 37.5570 ;
        RECT 21.7000 36.4635 21.7260 37.5570 ;
        RECT 21.5920 36.4635 21.6180 37.5570 ;
        RECT 21.4840 36.4635 21.5100 37.5570 ;
        RECT 21.3760 36.4635 21.4020 37.5570 ;
        RECT 21.2680 36.4635 21.2940 37.5570 ;
        RECT 21.1600 36.4635 21.1860 37.5570 ;
        RECT 21.0520 36.4635 21.0780 37.5570 ;
        RECT 20.9440 36.4635 20.9700 37.5570 ;
        RECT 20.8360 36.4635 20.8620 37.5570 ;
        RECT 20.7280 36.4635 20.7540 37.5570 ;
        RECT 20.6200 36.4635 20.6460 37.5570 ;
        RECT 20.5120 36.4635 20.5380 37.5570 ;
        RECT 20.4040 36.4635 20.4300 37.5570 ;
        RECT 20.2960 36.4635 20.3220 37.5570 ;
        RECT 20.1880 36.4635 20.2140 37.5570 ;
        RECT 20.0800 36.4635 20.1060 37.5570 ;
        RECT 19.9720 36.4635 19.9980 37.5570 ;
        RECT 19.8640 36.4635 19.8900 37.5570 ;
        RECT 19.7560 36.4635 19.7820 37.5570 ;
        RECT 19.6480 36.4635 19.6740 37.5570 ;
        RECT 19.5400 36.4635 19.5660 37.5570 ;
        RECT 19.4320 36.4635 19.4580 37.5570 ;
        RECT 19.3240 36.4635 19.3500 37.5570 ;
        RECT 19.2160 36.4635 19.2420 37.5570 ;
        RECT 19.1080 36.4635 19.1340 37.5570 ;
        RECT 19.0000 36.4635 19.0260 37.5570 ;
        RECT 18.8920 36.4635 18.9180 37.5570 ;
        RECT 18.7840 36.4635 18.8100 37.5570 ;
        RECT 18.6760 36.4635 18.7020 37.5570 ;
        RECT 18.5680 36.4635 18.5940 37.5570 ;
        RECT 18.4600 36.4635 18.4860 37.5570 ;
        RECT 18.3520 36.4635 18.3780 37.5570 ;
        RECT 18.2440 36.4635 18.2700 37.5570 ;
        RECT 18.1360 36.4635 18.1620 37.5570 ;
        RECT 18.0280 36.4635 18.0540 37.5570 ;
        RECT 17.9200 36.4635 17.9460 37.5570 ;
        RECT 17.8120 36.4635 17.8380 37.5570 ;
        RECT 17.7040 36.4635 17.7300 37.5570 ;
        RECT 17.5960 36.4635 17.6220 37.5570 ;
        RECT 17.4880 36.4635 17.5140 37.5570 ;
        RECT 17.3800 36.4635 17.4060 37.5570 ;
        RECT 17.2720 36.4635 17.2980 37.5570 ;
        RECT 17.1640 36.4635 17.1900 37.5570 ;
        RECT 17.0560 36.4635 17.0820 37.5570 ;
        RECT 16.9480 36.4635 16.9740 37.5570 ;
        RECT 16.8400 36.4635 16.8660 37.5570 ;
        RECT 16.7320 36.4635 16.7580 37.5570 ;
        RECT 16.6240 36.4635 16.6500 37.5570 ;
        RECT 16.5160 36.4635 16.5420 37.5570 ;
        RECT 16.4080 36.4635 16.4340 37.5570 ;
        RECT 16.3000 36.4635 16.3260 37.5570 ;
        RECT 16.0870 36.4635 16.1640 37.5570 ;
        RECT 14.1940 36.4635 14.2710 37.5570 ;
        RECT 14.0320 36.4635 14.0580 37.5570 ;
        RECT 13.9240 36.4635 13.9500 37.5570 ;
        RECT 13.8160 36.4635 13.8420 37.5570 ;
        RECT 13.7080 36.4635 13.7340 37.5570 ;
        RECT 13.6000 36.4635 13.6260 37.5570 ;
        RECT 13.4920 36.4635 13.5180 37.5570 ;
        RECT 13.3840 36.4635 13.4100 37.5570 ;
        RECT 13.2760 36.4635 13.3020 37.5570 ;
        RECT 13.1680 36.4635 13.1940 37.5570 ;
        RECT 13.0600 36.4635 13.0860 37.5570 ;
        RECT 12.9520 36.4635 12.9780 37.5570 ;
        RECT 12.8440 36.4635 12.8700 37.5570 ;
        RECT 12.7360 36.4635 12.7620 37.5570 ;
        RECT 12.6280 36.4635 12.6540 37.5570 ;
        RECT 12.5200 36.4635 12.5460 37.5570 ;
        RECT 12.4120 36.4635 12.4380 37.5570 ;
        RECT 12.3040 36.4635 12.3300 37.5570 ;
        RECT 12.1960 36.4635 12.2220 37.5570 ;
        RECT 12.0880 36.4635 12.1140 37.5570 ;
        RECT 11.9800 36.4635 12.0060 37.5570 ;
        RECT 11.8720 36.4635 11.8980 37.5570 ;
        RECT 11.7640 36.4635 11.7900 37.5570 ;
        RECT 11.6560 36.4635 11.6820 37.5570 ;
        RECT 11.5480 36.4635 11.5740 37.5570 ;
        RECT 11.4400 36.4635 11.4660 37.5570 ;
        RECT 11.3320 36.4635 11.3580 37.5570 ;
        RECT 11.2240 36.4635 11.2500 37.5570 ;
        RECT 11.1160 36.4635 11.1420 37.5570 ;
        RECT 11.0080 36.4635 11.0340 37.5570 ;
        RECT 10.9000 36.4635 10.9260 37.5570 ;
        RECT 10.7920 36.4635 10.8180 37.5570 ;
        RECT 10.6840 36.4635 10.7100 37.5570 ;
        RECT 10.5760 36.4635 10.6020 37.5570 ;
        RECT 10.4680 36.4635 10.4940 37.5570 ;
        RECT 10.3600 36.4635 10.3860 37.5570 ;
        RECT 10.2520 36.4635 10.2780 37.5570 ;
        RECT 10.1440 36.4635 10.1700 37.5570 ;
        RECT 10.0360 36.4635 10.0620 37.5570 ;
        RECT 9.9280 36.4635 9.9540 37.5570 ;
        RECT 9.8200 36.4635 9.8460 37.5570 ;
        RECT 9.7120 36.4635 9.7380 37.5570 ;
        RECT 9.6040 36.4635 9.6300 37.5570 ;
        RECT 9.4960 36.4635 9.5220 37.5570 ;
        RECT 9.3880 36.4635 9.4140 37.5570 ;
        RECT 9.2800 36.4635 9.3060 37.5570 ;
        RECT 9.1720 36.4635 9.1980 37.5570 ;
        RECT 9.0640 36.4635 9.0900 37.5570 ;
        RECT 8.9560 36.4635 8.9820 37.5570 ;
        RECT 8.8480 36.4635 8.8740 37.5570 ;
        RECT 8.7400 36.4635 8.7660 37.5570 ;
        RECT 8.6320 36.4635 8.6580 37.5570 ;
        RECT 8.5240 36.4635 8.5500 37.5570 ;
        RECT 8.4160 36.4635 8.4420 37.5570 ;
        RECT 8.3080 36.4635 8.3340 37.5570 ;
        RECT 8.2000 36.4635 8.2260 37.5570 ;
        RECT 8.0920 36.4635 8.1180 37.5570 ;
        RECT 7.9840 36.4635 8.0100 37.5570 ;
        RECT 7.8760 36.4635 7.9020 37.5570 ;
        RECT 7.7680 36.4635 7.7940 37.5570 ;
        RECT 7.6600 36.4635 7.6860 37.5570 ;
        RECT 7.5520 36.4635 7.5780 37.5570 ;
        RECT 7.4440 36.4635 7.4700 37.5570 ;
        RECT 7.3360 36.4635 7.3620 37.5570 ;
        RECT 7.2280 36.4635 7.2540 37.5570 ;
        RECT 7.1200 36.4635 7.1460 37.5570 ;
        RECT 7.0120 36.4635 7.0380 37.5570 ;
        RECT 6.9040 36.4635 6.9300 37.5570 ;
        RECT 6.7960 36.4635 6.8220 37.5570 ;
        RECT 6.6880 36.4635 6.7140 37.5570 ;
        RECT 6.5800 36.4635 6.6060 37.5570 ;
        RECT 6.4720 36.4635 6.4980 37.5570 ;
        RECT 6.3640 36.4635 6.3900 37.5570 ;
        RECT 6.2560 36.4635 6.2820 37.5570 ;
        RECT 6.1480 36.4635 6.1740 37.5570 ;
        RECT 6.0400 36.4635 6.0660 37.5570 ;
        RECT 5.9320 36.4635 5.9580 37.5570 ;
        RECT 5.8240 36.4635 5.8500 37.5570 ;
        RECT 5.7160 36.4635 5.7420 37.5570 ;
        RECT 5.6080 36.4635 5.6340 37.5570 ;
        RECT 5.5000 36.4635 5.5260 37.5570 ;
        RECT 5.3920 36.4635 5.4180 37.5570 ;
        RECT 5.2840 36.4635 5.3100 37.5570 ;
        RECT 5.1760 36.4635 5.2020 37.5570 ;
        RECT 5.0680 36.4635 5.0940 37.5570 ;
        RECT 4.9600 36.4635 4.9860 37.5570 ;
        RECT 4.8520 36.4635 4.8780 37.5570 ;
        RECT 4.7440 36.4635 4.7700 37.5570 ;
        RECT 4.6360 36.4635 4.6620 37.5570 ;
        RECT 4.5280 36.4635 4.5540 37.5570 ;
        RECT 4.4200 36.4635 4.4460 37.5570 ;
        RECT 4.3120 36.4635 4.3380 37.5570 ;
        RECT 4.2040 36.4635 4.2300 37.5570 ;
        RECT 4.0960 36.4635 4.1220 37.5570 ;
        RECT 3.9880 36.4635 4.0140 37.5570 ;
        RECT 3.8800 36.4635 3.9060 37.5570 ;
        RECT 3.7720 36.4635 3.7980 37.5570 ;
        RECT 3.6640 36.4635 3.6900 37.5570 ;
        RECT 3.5560 36.4635 3.5820 37.5570 ;
        RECT 3.4480 36.4635 3.4740 37.5570 ;
        RECT 3.3400 36.4635 3.3660 37.5570 ;
        RECT 3.2320 36.4635 3.2580 37.5570 ;
        RECT 3.1240 36.4635 3.1500 37.5570 ;
        RECT 3.0160 36.4635 3.0420 37.5570 ;
        RECT 2.9080 36.4635 2.9340 37.5570 ;
        RECT 2.8000 36.4635 2.8260 37.5570 ;
        RECT 2.6920 36.4635 2.7180 37.5570 ;
        RECT 2.5840 36.4635 2.6100 37.5570 ;
        RECT 2.4760 36.4635 2.5020 37.5570 ;
        RECT 2.3680 36.4635 2.3940 37.5570 ;
        RECT 2.2600 36.4635 2.2860 37.5570 ;
        RECT 2.1520 36.4635 2.1780 37.5570 ;
        RECT 2.0440 36.4635 2.0700 37.5570 ;
        RECT 1.9360 36.4635 1.9620 37.5570 ;
        RECT 1.8280 36.4635 1.8540 37.5570 ;
        RECT 1.7200 36.4635 1.7460 37.5570 ;
        RECT 1.6120 36.4635 1.6380 37.5570 ;
        RECT 1.5040 36.4635 1.5300 37.5570 ;
        RECT 1.3960 36.4635 1.4220 37.5570 ;
        RECT 1.2880 36.4635 1.3140 37.5570 ;
        RECT 1.1800 36.4635 1.2060 37.5570 ;
        RECT 1.0720 36.4635 1.0980 37.5570 ;
        RECT 0.9640 36.4635 0.9900 37.5570 ;
        RECT 0.8560 36.4635 0.8820 37.5570 ;
        RECT 0.7480 36.4635 0.7740 37.5570 ;
        RECT 0.6400 36.4635 0.6660 37.5570 ;
        RECT 0.5320 36.4635 0.5580 37.5570 ;
        RECT 0.4240 36.4635 0.4500 37.5570 ;
        RECT 0.3160 36.4635 0.3420 37.5570 ;
        RECT 0.2080 36.4635 0.2340 37.5570 ;
        RECT 0.0050 36.4635 0.0900 37.5570 ;
        RECT 15.5530 37.5435 15.6810 38.6370 ;
        RECT 15.5390 38.2090 15.6810 38.5315 ;
        RECT 15.3190 37.9360 15.4530 38.6370 ;
        RECT 15.2960 38.2710 15.4530 38.5290 ;
        RECT 15.3190 37.5435 15.4170 38.6370 ;
        RECT 15.3190 37.6645 15.4310 37.9040 ;
        RECT 15.3190 37.5435 15.4530 37.6325 ;
        RECT 15.0940 37.9940 15.2280 38.6370 ;
        RECT 15.0940 37.5435 15.1920 38.6370 ;
        RECT 14.6770 37.5435 14.7600 38.6370 ;
        RECT 14.6770 37.6320 14.7740 38.5675 ;
        RECT 30.2680 37.5435 30.3530 38.6370 ;
        RECT 30.1240 37.5435 30.1500 38.6370 ;
        RECT 30.0160 37.5435 30.0420 38.6370 ;
        RECT 29.9080 37.5435 29.9340 38.6370 ;
        RECT 29.8000 37.5435 29.8260 38.6370 ;
        RECT 29.6920 37.5435 29.7180 38.6370 ;
        RECT 29.5840 37.5435 29.6100 38.6370 ;
        RECT 29.4760 37.5435 29.5020 38.6370 ;
        RECT 29.3680 37.5435 29.3940 38.6370 ;
        RECT 29.2600 37.5435 29.2860 38.6370 ;
        RECT 29.1520 37.5435 29.1780 38.6370 ;
        RECT 29.0440 37.5435 29.0700 38.6370 ;
        RECT 28.9360 37.5435 28.9620 38.6370 ;
        RECT 28.8280 37.5435 28.8540 38.6370 ;
        RECT 28.7200 37.5435 28.7460 38.6370 ;
        RECT 28.6120 37.5435 28.6380 38.6370 ;
        RECT 28.5040 37.5435 28.5300 38.6370 ;
        RECT 28.3960 37.5435 28.4220 38.6370 ;
        RECT 28.2880 37.5435 28.3140 38.6370 ;
        RECT 28.1800 37.5435 28.2060 38.6370 ;
        RECT 28.0720 37.5435 28.0980 38.6370 ;
        RECT 27.9640 37.5435 27.9900 38.6370 ;
        RECT 27.8560 37.5435 27.8820 38.6370 ;
        RECT 27.7480 37.5435 27.7740 38.6370 ;
        RECT 27.6400 37.5435 27.6660 38.6370 ;
        RECT 27.5320 37.5435 27.5580 38.6370 ;
        RECT 27.4240 37.5435 27.4500 38.6370 ;
        RECT 27.3160 37.5435 27.3420 38.6370 ;
        RECT 27.2080 37.5435 27.2340 38.6370 ;
        RECT 27.1000 37.5435 27.1260 38.6370 ;
        RECT 26.9920 37.5435 27.0180 38.6370 ;
        RECT 26.8840 37.5435 26.9100 38.6370 ;
        RECT 26.7760 37.5435 26.8020 38.6370 ;
        RECT 26.6680 37.5435 26.6940 38.6370 ;
        RECT 26.5600 37.5435 26.5860 38.6370 ;
        RECT 26.4520 37.5435 26.4780 38.6370 ;
        RECT 26.3440 37.5435 26.3700 38.6370 ;
        RECT 26.2360 37.5435 26.2620 38.6370 ;
        RECT 26.1280 37.5435 26.1540 38.6370 ;
        RECT 26.0200 37.5435 26.0460 38.6370 ;
        RECT 25.9120 37.5435 25.9380 38.6370 ;
        RECT 25.8040 37.5435 25.8300 38.6370 ;
        RECT 25.6960 37.5435 25.7220 38.6370 ;
        RECT 25.5880 37.5435 25.6140 38.6370 ;
        RECT 25.4800 37.5435 25.5060 38.6370 ;
        RECT 25.3720 37.5435 25.3980 38.6370 ;
        RECT 25.2640 37.5435 25.2900 38.6370 ;
        RECT 25.1560 37.5435 25.1820 38.6370 ;
        RECT 25.0480 37.5435 25.0740 38.6370 ;
        RECT 24.9400 37.5435 24.9660 38.6370 ;
        RECT 24.8320 37.5435 24.8580 38.6370 ;
        RECT 24.7240 37.5435 24.7500 38.6370 ;
        RECT 24.6160 37.5435 24.6420 38.6370 ;
        RECT 24.5080 37.5435 24.5340 38.6370 ;
        RECT 24.4000 37.5435 24.4260 38.6370 ;
        RECT 24.2920 37.5435 24.3180 38.6370 ;
        RECT 24.1840 37.5435 24.2100 38.6370 ;
        RECT 24.0760 37.5435 24.1020 38.6370 ;
        RECT 23.9680 37.5435 23.9940 38.6370 ;
        RECT 23.8600 37.5435 23.8860 38.6370 ;
        RECT 23.7520 37.5435 23.7780 38.6370 ;
        RECT 23.6440 37.5435 23.6700 38.6370 ;
        RECT 23.5360 37.5435 23.5620 38.6370 ;
        RECT 23.4280 37.5435 23.4540 38.6370 ;
        RECT 23.3200 37.5435 23.3460 38.6370 ;
        RECT 23.2120 37.5435 23.2380 38.6370 ;
        RECT 23.1040 37.5435 23.1300 38.6370 ;
        RECT 22.9960 37.5435 23.0220 38.6370 ;
        RECT 22.8880 37.5435 22.9140 38.6370 ;
        RECT 22.7800 37.5435 22.8060 38.6370 ;
        RECT 22.6720 37.5435 22.6980 38.6370 ;
        RECT 22.5640 37.5435 22.5900 38.6370 ;
        RECT 22.4560 37.5435 22.4820 38.6370 ;
        RECT 22.3480 37.5435 22.3740 38.6370 ;
        RECT 22.2400 37.5435 22.2660 38.6370 ;
        RECT 22.1320 37.5435 22.1580 38.6370 ;
        RECT 22.0240 37.5435 22.0500 38.6370 ;
        RECT 21.9160 37.5435 21.9420 38.6370 ;
        RECT 21.8080 37.5435 21.8340 38.6370 ;
        RECT 21.7000 37.5435 21.7260 38.6370 ;
        RECT 21.5920 37.5435 21.6180 38.6370 ;
        RECT 21.4840 37.5435 21.5100 38.6370 ;
        RECT 21.3760 37.5435 21.4020 38.6370 ;
        RECT 21.2680 37.5435 21.2940 38.6370 ;
        RECT 21.1600 37.5435 21.1860 38.6370 ;
        RECT 21.0520 37.5435 21.0780 38.6370 ;
        RECT 20.9440 37.5435 20.9700 38.6370 ;
        RECT 20.8360 37.5435 20.8620 38.6370 ;
        RECT 20.7280 37.5435 20.7540 38.6370 ;
        RECT 20.6200 37.5435 20.6460 38.6370 ;
        RECT 20.5120 37.5435 20.5380 38.6370 ;
        RECT 20.4040 37.5435 20.4300 38.6370 ;
        RECT 20.2960 37.5435 20.3220 38.6370 ;
        RECT 20.1880 37.5435 20.2140 38.6370 ;
        RECT 20.0800 37.5435 20.1060 38.6370 ;
        RECT 19.9720 37.5435 19.9980 38.6370 ;
        RECT 19.8640 37.5435 19.8900 38.6370 ;
        RECT 19.7560 37.5435 19.7820 38.6370 ;
        RECT 19.6480 37.5435 19.6740 38.6370 ;
        RECT 19.5400 37.5435 19.5660 38.6370 ;
        RECT 19.4320 37.5435 19.4580 38.6370 ;
        RECT 19.3240 37.5435 19.3500 38.6370 ;
        RECT 19.2160 37.5435 19.2420 38.6370 ;
        RECT 19.1080 37.5435 19.1340 38.6370 ;
        RECT 19.0000 37.5435 19.0260 38.6370 ;
        RECT 18.8920 37.5435 18.9180 38.6370 ;
        RECT 18.7840 37.5435 18.8100 38.6370 ;
        RECT 18.6760 37.5435 18.7020 38.6370 ;
        RECT 18.5680 37.5435 18.5940 38.6370 ;
        RECT 18.4600 37.5435 18.4860 38.6370 ;
        RECT 18.3520 37.5435 18.3780 38.6370 ;
        RECT 18.2440 37.5435 18.2700 38.6370 ;
        RECT 18.1360 37.5435 18.1620 38.6370 ;
        RECT 18.0280 37.5435 18.0540 38.6370 ;
        RECT 17.9200 37.5435 17.9460 38.6370 ;
        RECT 17.8120 37.5435 17.8380 38.6370 ;
        RECT 17.7040 37.5435 17.7300 38.6370 ;
        RECT 17.5960 37.5435 17.6220 38.6370 ;
        RECT 17.4880 37.5435 17.5140 38.6370 ;
        RECT 17.3800 37.5435 17.4060 38.6370 ;
        RECT 17.2720 37.5435 17.2980 38.6370 ;
        RECT 17.1640 37.5435 17.1900 38.6370 ;
        RECT 17.0560 37.5435 17.0820 38.6370 ;
        RECT 16.9480 37.5435 16.9740 38.6370 ;
        RECT 16.8400 37.5435 16.8660 38.6370 ;
        RECT 16.7320 37.5435 16.7580 38.6370 ;
        RECT 16.6240 37.5435 16.6500 38.6370 ;
        RECT 16.5160 37.5435 16.5420 38.6370 ;
        RECT 16.4080 37.5435 16.4340 38.6370 ;
        RECT 16.3000 37.5435 16.3260 38.6370 ;
        RECT 16.0870 37.5435 16.1640 38.6370 ;
        RECT 14.1940 37.5435 14.2710 38.6370 ;
        RECT 14.0320 37.5435 14.0580 38.6370 ;
        RECT 13.9240 37.5435 13.9500 38.6370 ;
        RECT 13.8160 37.5435 13.8420 38.6370 ;
        RECT 13.7080 37.5435 13.7340 38.6370 ;
        RECT 13.6000 37.5435 13.6260 38.6370 ;
        RECT 13.4920 37.5435 13.5180 38.6370 ;
        RECT 13.3840 37.5435 13.4100 38.6370 ;
        RECT 13.2760 37.5435 13.3020 38.6370 ;
        RECT 13.1680 37.5435 13.1940 38.6370 ;
        RECT 13.0600 37.5435 13.0860 38.6370 ;
        RECT 12.9520 37.5435 12.9780 38.6370 ;
        RECT 12.8440 37.5435 12.8700 38.6370 ;
        RECT 12.7360 37.5435 12.7620 38.6370 ;
        RECT 12.6280 37.5435 12.6540 38.6370 ;
        RECT 12.5200 37.5435 12.5460 38.6370 ;
        RECT 12.4120 37.5435 12.4380 38.6370 ;
        RECT 12.3040 37.5435 12.3300 38.6370 ;
        RECT 12.1960 37.5435 12.2220 38.6370 ;
        RECT 12.0880 37.5435 12.1140 38.6370 ;
        RECT 11.9800 37.5435 12.0060 38.6370 ;
        RECT 11.8720 37.5435 11.8980 38.6370 ;
        RECT 11.7640 37.5435 11.7900 38.6370 ;
        RECT 11.6560 37.5435 11.6820 38.6370 ;
        RECT 11.5480 37.5435 11.5740 38.6370 ;
        RECT 11.4400 37.5435 11.4660 38.6370 ;
        RECT 11.3320 37.5435 11.3580 38.6370 ;
        RECT 11.2240 37.5435 11.2500 38.6370 ;
        RECT 11.1160 37.5435 11.1420 38.6370 ;
        RECT 11.0080 37.5435 11.0340 38.6370 ;
        RECT 10.9000 37.5435 10.9260 38.6370 ;
        RECT 10.7920 37.5435 10.8180 38.6370 ;
        RECT 10.6840 37.5435 10.7100 38.6370 ;
        RECT 10.5760 37.5435 10.6020 38.6370 ;
        RECT 10.4680 37.5435 10.4940 38.6370 ;
        RECT 10.3600 37.5435 10.3860 38.6370 ;
        RECT 10.2520 37.5435 10.2780 38.6370 ;
        RECT 10.1440 37.5435 10.1700 38.6370 ;
        RECT 10.0360 37.5435 10.0620 38.6370 ;
        RECT 9.9280 37.5435 9.9540 38.6370 ;
        RECT 9.8200 37.5435 9.8460 38.6370 ;
        RECT 9.7120 37.5435 9.7380 38.6370 ;
        RECT 9.6040 37.5435 9.6300 38.6370 ;
        RECT 9.4960 37.5435 9.5220 38.6370 ;
        RECT 9.3880 37.5435 9.4140 38.6370 ;
        RECT 9.2800 37.5435 9.3060 38.6370 ;
        RECT 9.1720 37.5435 9.1980 38.6370 ;
        RECT 9.0640 37.5435 9.0900 38.6370 ;
        RECT 8.9560 37.5435 8.9820 38.6370 ;
        RECT 8.8480 37.5435 8.8740 38.6370 ;
        RECT 8.7400 37.5435 8.7660 38.6370 ;
        RECT 8.6320 37.5435 8.6580 38.6370 ;
        RECT 8.5240 37.5435 8.5500 38.6370 ;
        RECT 8.4160 37.5435 8.4420 38.6370 ;
        RECT 8.3080 37.5435 8.3340 38.6370 ;
        RECT 8.2000 37.5435 8.2260 38.6370 ;
        RECT 8.0920 37.5435 8.1180 38.6370 ;
        RECT 7.9840 37.5435 8.0100 38.6370 ;
        RECT 7.8760 37.5435 7.9020 38.6370 ;
        RECT 7.7680 37.5435 7.7940 38.6370 ;
        RECT 7.6600 37.5435 7.6860 38.6370 ;
        RECT 7.5520 37.5435 7.5780 38.6370 ;
        RECT 7.4440 37.5435 7.4700 38.6370 ;
        RECT 7.3360 37.5435 7.3620 38.6370 ;
        RECT 7.2280 37.5435 7.2540 38.6370 ;
        RECT 7.1200 37.5435 7.1460 38.6370 ;
        RECT 7.0120 37.5435 7.0380 38.6370 ;
        RECT 6.9040 37.5435 6.9300 38.6370 ;
        RECT 6.7960 37.5435 6.8220 38.6370 ;
        RECT 6.6880 37.5435 6.7140 38.6370 ;
        RECT 6.5800 37.5435 6.6060 38.6370 ;
        RECT 6.4720 37.5435 6.4980 38.6370 ;
        RECT 6.3640 37.5435 6.3900 38.6370 ;
        RECT 6.2560 37.5435 6.2820 38.6370 ;
        RECT 6.1480 37.5435 6.1740 38.6370 ;
        RECT 6.0400 37.5435 6.0660 38.6370 ;
        RECT 5.9320 37.5435 5.9580 38.6370 ;
        RECT 5.8240 37.5435 5.8500 38.6370 ;
        RECT 5.7160 37.5435 5.7420 38.6370 ;
        RECT 5.6080 37.5435 5.6340 38.6370 ;
        RECT 5.5000 37.5435 5.5260 38.6370 ;
        RECT 5.3920 37.5435 5.4180 38.6370 ;
        RECT 5.2840 37.5435 5.3100 38.6370 ;
        RECT 5.1760 37.5435 5.2020 38.6370 ;
        RECT 5.0680 37.5435 5.0940 38.6370 ;
        RECT 4.9600 37.5435 4.9860 38.6370 ;
        RECT 4.8520 37.5435 4.8780 38.6370 ;
        RECT 4.7440 37.5435 4.7700 38.6370 ;
        RECT 4.6360 37.5435 4.6620 38.6370 ;
        RECT 4.5280 37.5435 4.5540 38.6370 ;
        RECT 4.4200 37.5435 4.4460 38.6370 ;
        RECT 4.3120 37.5435 4.3380 38.6370 ;
        RECT 4.2040 37.5435 4.2300 38.6370 ;
        RECT 4.0960 37.5435 4.1220 38.6370 ;
        RECT 3.9880 37.5435 4.0140 38.6370 ;
        RECT 3.8800 37.5435 3.9060 38.6370 ;
        RECT 3.7720 37.5435 3.7980 38.6370 ;
        RECT 3.6640 37.5435 3.6900 38.6370 ;
        RECT 3.5560 37.5435 3.5820 38.6370 ;
        RECT 3.4480 37.5435 3.4740 38.6370 ;
        RECT 3.3400 37.5435 3.3660 38.6370 ;
        RECT 3.2320 37.5435 3.2580 38.6370 ;
        RECT 3.1240 37.5435 3.1500 38.6370 ;
        RECT 3.0160 37.5435 3.0420 38.6370 ;
        RECT 2.9080 37.5435 2.9340 38.6370 ;
        RECT 2.8000 37.5435 2.8260 38.6370 ;
        RECT 2.6920 37.5435 2.7180 38.6370 ;
        RECT 2.5840 37.5435 2.6100 38.6370 ;
        RECT 2.4760 37.5435 2.5020 38.6370 ;
        RECT 2.3680 37.5435 2.3940 38.6370 ;
        RECT 2.2600 37.5435 2.2860 38.6370 ;
        RECT 2.1520 37.5435 2.1780 38.6370 ;
        RECT 2.0440 37.5435 2.0700 38.6370 ;
        RECT 1.9360 37.5435 1.9620 38.6370 ;
        RECT 1.8280 37.5435 1.8540 38.6370 ;
        RECT 1.7200 37.5435 1.7460 38.6370 ;
        RECT 1.6120 37.5435 1.6380 38.6370 ;
        RECT 1.5040 37.5435 1.5300 38.6370 ;
        RECT 1.3960 37.5435 1.4220 38.6370 ;
        RECT 1.2880 37.5435 1.3140 38.6370 ;
        RECT 1.1800 37.5435 1.2060 38.6370 ;
        RECT 1.0720 37.5435 1.0980 38.6370 ;
        RECT 0.9640 37.5435 0.9900 38.6370 ;
        RECT 0.8560 37.5435 0.8820 38.6370 ;
        RECT 0.7480 37.5435 0.7740 38.6370 ;
        RECT 0.6400 37.5435 0.6660 38.6370 ;
        RECT 0.5320 37.5435 0.5580 38.6370 ;
        RECT 0.4240 37.5435 0.4500 38.6370 ;
        RECT 0.3160 37.5435 0.3420 38.6370 ;
        RECT 0.2080 37.5435 0.2340 38.6370 ;
        RECT 0.0050 37.5435 0.0900 38.6370 ;
        RECT 15.5530 38.6235 15.6810 39.7170 ;
        RECT 15.5390 39.2890 15.6810 39.6115 ;
        RECT 15.3190 39.0160 15.4530 39.7170 ;
        RECT 15.2960 39.3510 15.4530 39.6090 ;
        RECT 15.3190 38.6235 15.4170 39.7170 ;
        RECT 15.3190 38.7445 15.4310 38.9840 ;
        RECT 15.3190 38.6235 15.4530 38.7125 ;
        RECT 15.0940 39.0740 15.2280 39.7170 ;
        RECT 15.0940 38.6235 15.1920 39.7170 ;
        RECT 14.6770 38.6235 14.7600 39.7170 ;
        RECT 14.6770 38.7120 14.7740 39.6475 ;
        RECT 30.2680 38.6235 30.3530 39.7170 ;
        RECT 30.1240 38.6235 30.1500 39.7170 ;
        RECT 30.0160 38.6235 30.0420 39.7170 ;
        RECT 29.9080 38.6235 29.9340 39.7170 ;
        RECT 29.8000 38.6235 29.8260 39.7170 ;
        RECT 29.6920 38.6235 29.7180 39.7170 ;
        RECT 29.5840 38.6235 29.6100 39.7170 ;
        RECT 29.4760 38.6235 29.5020 39.7170 ;
        RECT 29.3680 38.6235 29.3940 39.7170 ;
        RECT 29.2600 38.6235 29.2860 39.7170 ;
        RECT 29.1520 38.6235 29.1780 39.7170 ;
        RECT 29.0440 38.6235 29.0700 39.7170 ;
        RECT 28.9360 38.6235 28.9620 39.7170 ;
        RECT 28.8280 38.6235 28.8540 39.7170 ;
        RECT 28.7200 38.6235 28.7460 39.7170 ;
        RECT 28.6120 38.6235 28.6380 39.7170 ;
        RECT 28.5040 38.6235 28.5300 39.7170 ;
        RECT 28.3960 38.6235 28.4220 39.7170 ;
        RECT 28.2880 38.6235 28.3140 39.7170 ;
        RECT 28.1800 38.6235 28.2060 39.7170 ;
        RECT 28.0720 38.6235 28.0980 39.7170 ;
        RECT 27.9640 38.6235 27.9900 39.7170 ;
        RECT 27.8560 38.6235 27.8820 39.7170 ;
        RECT 27.7480 38.6235 27.7740 39.7170 ;
        RECT 27.6400 38.6235 27.6660 39.7170 ;
        RECT 27.5320 38.6235 27.5580 39.7170 ;
        RECT 27.4240 38.6235 27.4500 39.7170 ;
        RECT 27.3160 38.6235 27.3420 39.7170 ;
        RECT 27.2080 38.6235 27.2340 39.7170 ;
        RECT 27.1000 38.6235 27.1260 39.7170 ;
        RECT 26.9920 38.6235 27.0180 39.7170 ;
        RECT 26.8840 38.6235 26.9100 39.7170 ;
        RECT 26.7760 38.6235 26.8020 39.7170 ;
        RECT 26.6680 38.6235 26.6940 39.7170 ;
        RECT 26.5600 38.6235 26.5860 39.7170 ;
        RECT 26.4520 38.6235 26.4780 39.7170 ;
        RECT 26.3440 38.6235 26.3700 39.7170 ;
        RECT 26.2360 38.6235 26.2620 39.7170 ;
        RECT 26.1280 38.6235 26.1540 39.7170 ;
        RECT 26.0200 38.6235 26.0460 39.7170 ;
        RECT 25.9120 38.6235 25.9380 39.7170 ;
        RECT 25.8040 38.6235 25.8300 39.7170 ;
        RECT 25.6960 38.6235 25.7220 39.7170 ;
        RECT 25.5880 38.6235 25.6140 39.7170 ;
        RECT 25.4800 38.6235 25.5060 39.7170 ;
        RECT 25.3720 38.6235 25.3980 39.7170 ;
        RECT 25.2640 38.6235 25.2900 39.7170 ;
        RECT 25.1560 38.6235 25.1820 39.7170 ;
        RECT 25.0480 38.6235 25.0740 39.7170 ;
        RECT 24.9400 38.6235 24.9660 39.7170 ;
        RECT 24.8320 38.6235 24.8580 39.7170 ;
        RECT 24.7240 38.6235 24.7500 39.7170 ;
        RECT 24.6160 38.6235 24.6420 39.7170 ;
        RECT 24.5080 38.6235 24.5340 39.7170 ;
        RECT 24.4000 38.6235 24.4260 39.7170 ;
        RECT 24.2920 38.6235 24.3180 39.7170 ;
        RECT 24.1840 38.6235 24.2100 39.7170 ;
        RECT 24.0760 38.6235 24.1020 39.7170 ;
        RECT 23.9680 38.6235 23.9940 39.7170 ;
        RECT 23.8600 38.6235 23.8860 39.7170 ;
        RECT 23.7520 38.6235 23.7780 39.7170 ;
        RECT 23.6440 38.6235 23.6700 39.7170 ;
        RECT 23.5360 38.6235 23.5620 39.7170 ;
        RECT 23.4280 38.6235 23.4540 39.7170 ;
        RECT 23.3200 38.6235 23.3460 39.7170 ;
        RECT 23.2120 38.6235 23.2380 39.7170 ;
        RECT 23.1040 38.6235 23.1300 39.7170 ;
        RECT 22.9960 38.6235 23.0220 39.7170 ;
        RECT 22.8880 38.6235 22.9140 39.7170 ;
        RECT 22.7800 38.6235 22.8060 39.7170 ;
        RECT 22.6720 38.6235 22.6980 39.7170 ;
        RECT 22.5640 38.6235 22.5900 39.7170 ;
        RECT 22.4560 38.6235 22.4820 39.7170 ;
        RECT 22.3480 38.6235 22.3740 39.7170 ;
        RECT 22.2400 38.6235 22.2660 39.7170 ;
        RECT 22.1320 38.6235 22.1580 39.7170 ;
        RECT 22.0240 38.6235 22.0500 39.7170 ;
        RECT 21.9160 38.6235 21.9420 39.7170 ;
        RECT 21.8080 38.6235 21.8340 39.7170 ;
        RECT 21.7000 38.6235 21.7260 39.7170 ;
        RECT 21.5920 38.6235 21.6180 39.7170 ;
        RECT 21.4840 38.6235 21.5100 39.7170 ;
        RECT 21.3760 38.6235 21.4020 39.7170 ;
        RECT 21.2680 38.6235 21.2940 39.7170 ;
        RECT 21.1600 38.6235 21.1860 39.7170 ;
        RECT 21.0520 38.6235 21.0780 39.7170 ;
        RECT 20.9440 38.6235 20.9700 39.7170 ;
        RECT 20.8360 38.6235 20.8620 39.7170 ;
        RECT 20.7280 38.6235 20.7540 39.7170 ;
        RECT 20.6200 38.6235 20.6460 39.7170 ;
        RECT 20.5120 38.6235 20.5380 39.7170 ;
        RECT 20.4040 38.6235 20.4300 39.7170 ;
        RECT 20.2960 38.6235 20.3220 39.7170 ;
        RECT 20.1880 38.6235 20.2140 39.7170 ;
        RECT 20.0800 38.6235 20.1060 39.7170 ;
        RECT 19.9720 38.6235 19.9980 39.7170 ;
        RECT 19.8640 38.6235 19.8900 39.7170 ;
        RECT 19.7560 38.6235 19.7820 39.7170 ;
        RECT 19.6480 38.6235 19.6740 39.7170 ;
        RECT 19.5400 38.6235 19.5660 39.7170 ;
        RECT 19.4320 38.6235 19.4580 39.7170 ;
        RECT 19.3240 38.6235 19.3500 39.7170 ;
        RECT 19.2160 38.6235 19.2420 39.7170 ;
        RECT 19.1080 38.6235 19.1340 39.7170 ;
        RECT 19.0000 38.6235 19.0260 39.7170 ;
        RECT 18.8920 38.6235 18.9180 39.7170 ;
        RECT 18.7840 38.6235 18.8100 39.7170 ;
        RECT 18.6760 38.6235 18.7020 39.7170 ;
        RECT 18.5680 38.6235 18.5940 39.7170 ;
        RECT 18.4600 38.6235 18.4860 39.7170 ;
        RECT 18.3520 38.6235 18.3780 39.7170 ;
        RECT 18.2440 38.6235 18.2700 39.7170 ;
        RECT 18.1360 38.6235 18.1620 39.7170 ;
        RECT 18.0280 38.6235 18.0540 39.7170 ;
        RECT 17.9200 38.6235 17.9460 39.7170 ;
        RECT 17.8120 38.6235 17.8380 39.7170 ;
        RECT 17.7040 38.6235 17.7300 39.7170 ;
        RECT 17.5960 38.6235 17.6220 39.7170 ;
        RECT 17.4880 38.6235 17.5140 39.7170 ;
        RECT 17.3800 38.6235 17.4060 39.7170 ;
        RECT 17.2720 38.6235 17.2980 39.7170 ;
        RECT 17.1640 38.6235 17.1900 39.7170 ;
        RECT 17.0560 38.6235 17.0820 39.7170 ;
        RECT 16.9480 38.6235 16.9740 39.7170 ;
        RECT 16.8400 38.6235 16.8660 39.7170 ;
        RECT 16.7320 38.6235 16.7580 39.7170 ;
        RECT 16.6240 38.6235 16.6500 39.7170 ;
        RECT 16.5160 38.6235 16.5420 39.7170 ;
        RECT 16.4080 38.6235 16.4340 39.7170 ;
        RECT 16.3000 38.6235 16.3260 39.7170 ;
        RECT 16.0870 38.6235 16.1640 39.7170 ;
        RECT 14.1940 38.6235 14.2710 39.7170 ;
        RECT 14.0320 38.6235 14.0580 39.7170 ;
        RECT 13.9240 38.6235 13.9500 39.7170 ;
        RECT 13.8160 38.6235 13.8420 39.7170 ;
        RECT 13.7080 38.6235 13.7340 39.7170 ;
        RECT 13.6000 38.6235 13.6260 39.7170 ;
        RECT 13.4920 38.6235 13.5180 39.7170 ;
        RECT 13.3840 38.6235 13.4100 39.7170 ;
        RECT 13.2760 38.6235 13.3020 39.7170 ;
        RECT 13.1680 38.6235 13.1940 39.7170 ;
        RECT 13.0600 38.6235 13.0860 39.7170 ;
        RECT 12.9520 38.6235 12.9780 39.7170 ;
        RECT 12.8440 38.6235 12.8700 39.7170 ;
        RECT 12.7360 38.6235 12.7620 39.7170 ;
        RECT 12.6280 38.6235 12.6540 39.7170 ;
        RECT 12.5200 38.6235 12.5460 39.7170 ;
        RECT 12.4120 38.6235 12.4380 39.7170 ;
        RECT 12.3040 38.6235 12.3300 39.7170 ;
        RECT 12.1960 38.6235 12.2220 39.7170 ;
        RECT 12.0880 38.6235 12.1140 39.7170 ;
        RECT 11.9800 38.6235 12.0060 39.7170 ;
        RECT 11.8720 38.6235 11.8980 39.7170 ;
        RECT 11.7640 38.6235 11.7900 39.7170 ;
        RECT 11.6560 38.6235 11.6820 39.7170 ;
        RECT 11.5480 38.6235 11.5740 39.7170 ;
        RECT 11.4400 38.6235 11.4660 39.7170 ;
        RECT 11.3320 38.6235 11.3580 39.7170 ;
        RECT 11.2240 38.6235 11.2500 39.7170 ;
        RECT 11.1160 38.6235 11.1420 39.7170 ;
        RECT 11.0080 38.6235 11.0340 39.7170 ;
        RECT 10.9000 38.6235 10.9260 39.7170 ;
        RECT 10.7920 38.6235 10.8180 39.7170 ;
        RECT 10.6840 38.6235 10.7100 39.7170 ;
        RECT 10.5760 38.6235 10.6020 39.7170 ;
        RECT 10.4680 38.6235 10.4940 39.7170 ;
        RECT 10.3600 38.6235 10.3860 39.7170 ;
        RECT 10.2520 38.6235 10.2780 39.7170 ;
        RECT 10.1440 38.6235 10.1700 39.7170 ;
        RECT 10.0360 38.6235 10.0620 39.7170 ;
        RECT 9.9280 38.6235 9.9540 39.7170 ;
        RECT 9.8200 38.6235 9.8460 39.7170 ;
        RECT 9.7120 38.6235 9.7380 39.7170 ;
        RECT 9.6040 38.6235 9.6300 39.7170 ;
        RECT 9.4960 38.6235 9.5220 39.7170 ;
        RECT 9.3880 38.6235 9.4140 39.7170 ;
        RECT 9.2800 38.6235 9.3060 39.7170 ;
        RECT 9.1720 38.6235 9.1980 39.7170 ;
        RECT 9.0640 38.6235 9.0900 39.7170 ;
        RECT 8.9560 38.6235 8.9820 39.7170 ;
        RECT 8.8480 38.6235 8.8740 39.7170 ;
        RECT 8.7400 38.6235 8.7660 39.7170 ;
        RECT 8.6320 38.6235 8.6580 39.7170 ;
        RECT 8.5240 38.6235 8.5500 39.7170 ;
        RECT 8.4160 38.6235 8.4420 39.7170 ;
        RECT 8.3080 38.6235 8.3340 39.7170 ;
        RECT 8.2000 38.6235 8.2260 39.7170 ;
        RECT 8.0920 38.6235 8.1180 39.7170 ;
        RECT 7.9840 38.6235 8.0100 39.7170 ;
        RECT 7.8760 38.6235 7.9020 39.7170 ;
        RECT 7.7680 38.6235 7.7940 39.7170 ;
        RECT 7.6600 38.6235 7.6860 39.7170 ;
        RECT 7.5520 38.6235 7.5780 39.7170 ;
        RECT 7.4440 38.6235 7.4700 39.7170 ;
        RECT 7.3360 38.6235 7.3620 39.7170 ;
        RECT 7.2280 38.6235 7.2540 39.7170 ;
        RECT 7.1200 38.6235 7.1460 39.7170 ;
        RECT 7.0120 38.6235 7.0380 39.7170 ;
        RECT 6.9040 38.6235 6.9300 39.7170 ;
        RECT 6.7960 38.6235 6.8220 39.7170 ;
        RECT 6.6880 38.6235 6.7140 39.7170 ;
        RECT 6.5800 38.6235 6.6060 39.7170 ;
        RECT 6.4720 38.6235 6.4980 39.7170 ;
        RECT 6.3640 38.6235 6.3900 39.7170 ;
        RECT 6.2560 38.6235 6.2820 39.7170 ;
        RECT 6.1480 38.6235 6.1740 39.7170 ;
        RECT 6.0400 38.6235 6.0660 39.7170 ;
        RECT 5.9320 38.6235 5.9580 39.7170 ;
        RECT 5.8240 38.6235 5.8500 39.7170 ;
        RECT 5.7160 38.6235 5.7420 39.7170 ;
        RECT 5.6080 38.6235 5.6340 39.7170 ;
        RECT 5.5000 38.6235 5.5260 39.7170 ;
        RECT 5.3920 38.6235 5.4180 39.7170 ;
        RECT 5.2840 38.6235 5.3100 39.7170 ;
        RECT 5.1760 38.6235 5.2020 39.7170 ;
        RECT 5.0680 38.6235 5.0940 39.7170 ;
        RECT 4.9600 38.6235 4.9860 39.7170 ;
        RECT 4.8520 38.6235 4.8780 39.7170 ;
        RECT 4.7440 38.6235 4.7700 39.7170 ;
        RECT 4.6360 38.6235 4.6620 39.7170 ;
        RECT 4.5280 38.6235 4.5540 39.7170 ;
        RECT 4.4200 38.6235 4.4460 39.7170 ;
        RECT 4.3120 38.6235 4.3380 39.7170 ;
        RECT 4.2040 38.6235 4.2300 39.7170 ;
        RECT 4.0960 38.6235 4.1220 39.7170 ;
        RECT 3.9880 38.6235 4.0140 39.7170 ;
        RECT 3.8800 38.6235 3.9060 39.7170 ;
        RECT 3.7720 38.6235 3.7980 39.7170 ;
        RECT 3.6640 38.6235 3.6900 39.7170 ;
        RECT 3.5560 38.6235 3.5820 39.7170 ;
        RECT 3.4480 38.6235 3.4740 39.7170 ;
        RECT 3.3400 38.6235 3.3660 39.7170 ;
        RECT 3.2320 38.6235 3.2580 39.7170 ;
        RECT 3.1240 38.6235 3.1500 39.7170 ;
        RECT 3.0160 38.6235 3.0420 39.7170 ;
        RECT 2.9080 38.6235 2.9340 39.7170 ;
        RECT 2.8000 38.6235 2.8260 39.7170 ;
        RECT 2.6920 38.6235 2.7180 39.7170 ;
        RECT 2.5840 38.6235 2.6100 39.7170 ;
        RECT 2.4760 38.6235 2.5020 39.7170 ;
        RECT 2.3680 38.6235 2.3940 39.7170 ;
        RECT 2.2600 38.6235 2.2860 39.7170 ;
        RECT 2.1520 38.6235 2.1780 39.7170 ;
        RECT 2.0440 38.6235 2.0700 39.7170 ;
        RECT 1.9360 38.6235 1.9620 39.7170 ;
        RECT 1.8280 38.6235 1.8540 39.7170 ;
        RECT 1.7200 38.6235 1.7460 39.7170 ;
        RECT 1.6120 38.6235 1.6380 39.7170 ;
        RECT 1.5040 38.6235 1.5300 39.7170 ;
        RECT 1.3960 38.6235 1.4220 39.7170 ;
        RECT 1.2880 38.6235 1.3140 39.7170 ;
        RECT 1.1800 38.6235 1.2060 39.7170 ;
        RECT 1.0720 38.6235 1.0980 39.7170 ;
        RECT 0.9640 38.6235 0.9900 39.7170 ;
        RECT 0.8560 38.6235 0.8820 39.7170 ;
        RECT 0.7480 38.6235 0.7740 39.7170 ;
        RECT 0.6400 38.6235 0.6660 39.7170 ;
        RECT 0.5320 38.6235 0.5580 39.7170 ;
        RECT 0.4240 38.6235 0.4500 39.7170 ;
        RECT 0.3160 38.6235 0.3420 39.7170 ;
        RECT 0.2080 38.6235 0.2340 39.7170 ;
        RECT 0.0050 38.6235 0.0900 39.7170 ;
        RECT 15.5530 39.7035 15.6810 40.7970 ;
        RECT 15.5390 40.3690 15.6810 40.6915 ;
        RECT 15.3190 40.0960 15.4530 40.7970 ;
        RECT 15.2960 40.4310 15.4530 40.6890 ;
        RECT 15.3190 39.7035 15.4170 40.7970 ;
        RECT 15.3190 39.8245 15.4310 40.0640 ;
        RECT 15.3190 39.7035 15.4530 39.7925 ;
        RECT 15.0940 40.1540 15.2280 40.7970 ;
        RECT 15.0940 39.7035 15.1920 40.7970 ;
        RECT 14.6770 39.7035 14.7600 40.7970 ;
        RECT 14.6770 39.7920 14.7740 40.7275 ;
        RECT 30.2680 39.7035 30.3530 40.7970 ;
        RECT 30.1240 39.7035 30.1500 40.7970 ;
        RECT 30.0160 39.7035 30.0420 40.7970 ;
        RECT 29.9080 39.7035 29.9340 40.7970 ;
        RECT 29.8000 39.7035 29.8260 40.7970 ;
        RECT 29.6920 39.7035 29.7180 40.7970 ;
        RECT 29.5840 39.7035 29.6100 40.7970 ;
        RECT 29.4760 39.7035 29.5020 40.7970 ;
        RECT 29.3680 39.7035 29.3940 40.7970 ;
        RECT 29.2600 39.7035 29.2860 40.7970 ;
        RECT 29.1520 39.7035 29.1780 40.7970 ;
        RECT 29.0440 39.7035 29.0700 40.7970 ;
        RECT 28.9360 39.7035 28.9620 40.7970 ;
        RECT 28.8280 39.7035 28.8540 40.7970 ;
        RECT 28.7200 39.7035 28.7460 40.7970 ;
        RECT 28.6120 39.7035 28.6380 40.7970 ;
        RECT 28.5040 39.7035 28.5300 40.7970 ;
        RECT 28.3960 39.7035 28.4220 40.7970 ;
        RECT 28.2880 39.7035 28.3140 40.7970 ;
        RECT 28.1800 39.7035 28.2060 40.7970 ;
        RECT 28.0720 39.7035 28.0980 40.7970 ;
        RECT 27.9640 39.7035 27.9900 40.7970 ;
        RECT 27.8560 39.7035 27.8820 40.7970 ;
        RECT 27.7480 39.7035 27.7740 40.7970 ;
        RECT 27.6400 39.7035 27.6660 40.7970 ;
        RECT 27.5320 39.7035 27.5580 40.7970 ;
        RECT 27.4240 39.7035 27.4500 40.7970 ;
        RECT 27.3160 39.7035 27.3420 40.7970 ;
        RECT 27.2080 39.7035 27.2340 40.7970 ;
        RECT 27.1000 39.7035 27.1260 40.7970 ;
        RECT 26.9920 39.7035 27.0180 40.7970 ;
        RECT 26.8840 39.7035 26.9100 40.7970 ;
        RECT 26.7760 39.7035 26.8020 40.7970 ;
        RECT 26.6680 39.7035 26.6940 40.7970 ;
        RECT 26.5600 39.7035 26.5860 40.7970 ;
        RECT 26.4520 39.7035 26.4780 40.7970 ;
        RECT 26.3440 39.7035 26.3700 40.7970 ;
        RECT 26.2360 39.7035 26.2620 40.7970 ;
        RECT 26.1280 39.7035 26.1540 40.7970 ;
        RECT 26.0200 39.7035 26.0460 40.7970 ;
        RECT 25.9120 39.7035 25.9380 40.7970 ;
        RECT 25.8040 39.7035 25.8300 40.7970 ;
        RECT 25.6960 39.7035 25.7220 40.7970 ;
        RECT 25.5880 39.7035 25.6140 40.7970 ;
        RECT 25.4800 39.7035 25.5060 40.7970 ;
        RECT 25.3720 39.7035 25.3980 40.7970 ;
        RECT 25.2640 39.7035 25.2900 40.7970 ;
        RECT 25.1560 39.7035 25.1820 40.7970 ;
        RECT 25.0480 39.7035 25.0740 40.7970 ;
        RECT 24.9400 39.7035 24.9660 40.7970 ;
        RECT 24.8320 39.7035 24.8580 40.7970 ;
        RECT 24.7240 39.7035 24.7500 40.7970 ;
        RECT 24.6160 39.7035 24.6420 40.7970 ;
        RECT 24.5080 39.7035 24.5340 40.7970 ;
        RECT 24.4000 39.7035 24.4260 40.7970 ;
        RECT 24.2920 39.7035 24.3180 40.7970 ;
        RECT 24.1840 39.7035 24.2100 40.7970 ;
        RECT 24.0760 39.7035 24.1020 40.7970 ;
        RECT 23.9680 39.7035 23.9940 40.7970 ;
        RECT 23.8600 39.7035 23.8860 40.7970 ;
        RECT 23.7520 39.7035 23.7780 40.7970 ;
        RECT 23.6440 39.7035 23.6700 40.7970 ;
        RECT 23.5360 39.7035 23.5620 40.7970 ;
        RECT 23.4280 39.7035 23.4540 40.7970 ;
        RECT 23.3200 39.7035 23.3460 40.7970 ;
        RECT 23.2120 39.7035 23.2380 40.7970 ;
        RECT 23.1040 39.7035 23.1300 40.7970 ;
        RECT 22.9960 39.7035 23.0220 40.7970 ;
        RECT 22.8880 39.7035 22.9140 40.7970 ;
        RECT 22.7800 39.7035 22.8060 40.7970 ;
        RECT 22.6720 39.7035 22.6980 40.7970 ;
        RECT 22.5640 39.7035 22.5900 40.7970 ;
        RECT 22.4560 39.7035 22.4820 40.7970 ;
        RECT 22.3480 39.7035 22.3740 40.7970 ;
        RECT 22.2400 39.7035 22.2660 40.7970 ;
        RECT 22.1320 39.7035 22.1580 40.7970 ;
        RECT 22.0240 39.7035 22.0500 40.7970 ;
        RECT 21.9160 39.7035 21.9420 40.7970 ;
        RECT 21.8080 39.7035 21.8340 40.7970 ;
        RECT 21.7000 39.7035 21.7260 40.7970 ;
        RECT 21.5920 39.7035 21.6180 40.7970 ;
        RECT 21.4840 39.7035 21.5100 40.7970 ;
        RECT 21.3760 39.7035 21.4020 40.7970 ;
        RECT 21.2680 39.7035 21.2940 40.7970 ;
        RECT 21.1600 39.7035 21.1860 40.7970 ;
        RECT 21.0520 39.7035 21.0780 40.7970 ;
        RECT 20.9440 39.7035 20.9700 40.7970 ;
        RECT 20.8360 39.7035 20.8620 40.7970 ;
        RECT 20.7280 39.7035 20.7540 40.7970 ;
        RECT 20.6200 39.7035 20.6460 40.7970 ;
        RECT 20.5120 39.7035 20.5380 40.7970 ;
        RECT 20.4040 39.7035 20.4300 40.7970 ;
        RECT 20.2960 39.7035 20.3220 40.7970 ;
        RECT 20.1880 39.7035 20.2140 40.7970 ;
        RECT 20.0800 39.7035 20.1060 40.7970 ;
        RECT 19.9720 39.7035 19.9980 40.7970 ;
        RECT 19.8640 39.7035 19.8900 40.7970 ;
        RECT 19.7560 39.7035 19.7820 40.7970 ;
        RECT 19.6480 39.7035 19.6740 40.7970 ;
        RECT 19.5400 39.7035 19.5660 40.7970 ;
        RECT 19.4320 39.7035 19.4580 40.7970 ;
        RECT 19.3240 39.7035 19.3500 40.7970 ;
        RECT 19.2160 39.7035 19.2420 40.7970 ;
        RECT 19.1080 39.7035 19.1340 40.7970 ;
        RECT 19.0000 39.7035 19.0260 40.7970 ;
        RECT 18.8920 39.7035 18.9180 40.7970 ;
        RECT 18.7840 39.7035 18.8100 40.7970 ;
        RECT 18.6760 39.7035 18.7020 40.7970 ;
        RECT 18.5680 39.7035 18.5940 40.7970 ;
        RECT 18.4600 39.7035 18.4860 40.7970 ;
        RECT 18.3520 39.7035 18.3780 40.7970 ;
        RECT 18.2440 39.7035 18.2700 40.7970 ;
        RECT 18.1360 39.7035 18.1620 40.7970 ;
        RECT 18.0280 39.7035 18.0540 40.7970 ;
        RECT 17.9200 39.7035 17.9460 40.7970 ;
        RECT 17.8120 39.7035 17.8380 40.7970 ;
        RECT 17.7040 39.7035 17.7300 40.7970 ;
        RECT 17.5960 39.7035 17.6220 40.7970 ;
        RECT 17.4880 39.7035 17.5140 40.7970 ;
        RECT 17.3800 39.7035 17.4060 40.7970 ;
        RECT 17.2720 39.7035 17.2980 40.7970 ;
        RECT 17.1640 39.7035 17.1900 40.7970 ;
        RECT 17.0560 39.7035 17.0820 40.7970 ;
        RECT 16.9480 39.7035 16.9740 40.7970 ;
        RECT 16.8400 39.7035 16.8660 40.7970 ;
        RECT 16.7320 39.7035 16.7580 40.7970 ;
        RECT 16.6240 39.7035 16.6500 40.7970 ;
        RECT 16.5160 39.7035 16.5420 40.7970 ;
        RECT 16.4080 39.7035 16.4340 40.7970 ;
        RECT 16.3000 39.7035 16.3260 40.7970 ;
        RECT 16.0870 39.7035 16.1640 40.7970 ;
        RECT 14.1940 39.7035 14.2710 40.7970 ;
        RECT 14.0320 39.7035 14.0580 40.7970 ;
        RECT 13.9240 39.7035 13.9500 40.7970 ;
        RECT 13.8160 39.7035 13.8420 40.7970 ;
        RECT 13.7080 39.7035 13.7340 40.7970 ;
        RECT 13.6000 39.7035 13.6260 40.7970 ;
        RECT 13.4920 39.7035 13.5180 40.7970 ;
        RECT 13.3840 39.7035 13.4100 40.7970 ;
        RECT 13.2760 39.7035 13.3020 40.7970 ;
        RECT 13.1680 39.7035 13.1940 40.7970 ;
        RECT 13.0600 39.7035 13.0860 40.7970 ;
        RECT 12.9520 39.7035 12.9780 40.7970 ;
        RECT 12.8440 39.7035 12.8700 40.7970 ;
        RECT 12.7360 39.7035 12.7620 40.7970 ;
        RECT 12.6280 39.7035 12.6540 40.7970 ;
        RECT 12.5200 39.7035 12.5460 40.7970 ;
        RECT 12.4120 39.7035 12.4380 40.7970 ;
        RECT 12.3040 39.7035 12.3300 40.7970 ;
        RECT 12.1960 39.7035 12.2220 40.7970 ;
        RECT 12.0880 39.7035 12.1140 40.7970 ;
        RECT 11.9800 39.7035 12.0060 40.7970 ;
        RECT 11.8720 39.7035 11.8980 40.7970 ;
        RECT 11.7640 39.7035 11.7900 40.7970 ;
        RECT 11.6560 39.7035 11.6820 40.7970 ;
        RECT 11.5480 39.7035 11.5740 40.7970 ;
        RECT 11.4400 39.7035 11.4660 40.7970 ;
        RECT 11.3320 39.7035 11.3580 40.7970 ;
        RECT 11.2240 39.7035 11.2500 40.7970 ;
        RECT 11.1160 39.7035 11.1420 40.7970 ;
        RECT 11.0080 39.7035 11.0340 40.7970 ;
        RECT 10.9000 39.7035 10.9260 40.7970 ;
        RECT 10.7920 39.7035 10.8180 40.7970 ;
        RECT 10.6840 39.7035 10.7100 40.7970 ;
        RECT 10.5760 39.7035 10.6020 40.7970 ;
        RECT 10.4680 39.7035 10.4940 40.7970 ;
        RECT 10.3600 39.7035 10.3860 40.7970 ;
        RECT 10.2520 39.7035 10.2780 40.7970 ;
        RECT 10.1440 39.7035 10.1700 40.7970 ;
        RECT 10.0360 39.7035 10.0620 40.7970 ;
        RECT 9.9280 39.7035 9.9540 40.7970 ;
        RECT 9.8200 39.7035 9.8460 40.7970 ;
        RECT 9.7120 39.7035 9.7380 40.7970 ;
        RECT 9.6040 39.7035 9.6300 40.7970 ;
        RECT 9.4960 39.7035 9.5220 40.7970 ;
        RECT 9.3880 39.7035 9.4140 40.7970 ;
        RECT 9.2800 39.7035 9.3060 40.7970 ;
        RECT 9.1720 39.7035 9.1980 40.7970 ;
        RECT 9.0640 39.7035 9.0900 40.7970 ;
        RECT 8.9560 39.7035 8.9820 40.7970 ;
        RECT 8.8480 39.7035 8.8740 40.7970 ;
        RECT 8.7400 39.7035 8.7660 40.7970 ;
        RECT 8.6320 39.7035 8.6580 40.7970 ;
        RECT 8.5240 39.7035 8.5500 40.7970 ;
        RECT 8.4160 39.7035 8.4420 40.7970 ;
        RECT 8.3080 39.7035 8.3340 40.7970 ;
        RECT 8.2000 39.7035 8.2260 40.7970 ;
        RECT 8.0920 39.7035 8.1180 40.7970 ;
        RECT 7.9840 39.7035 8.0100 40.7970 ;
        RECT 7.8760 39.7035 7.9020 40.7970 ;
        RECT 7.7680 39.7035 7.7940 40.7970 ;
        RECT 7.6600 39.7035 7.6860 40.7970 ;
        RECT 7.5520 39.7035 7.5780 40.7970 ;
        RECT 7.4440 39.7035 7.4700 40.7970 ;
        RECT 7.3360 39.7035 7.3620 40.7970 ;
        RECT 7.2280 39.7035 7.2540 40.7970 ;
        RECT 7.1200 39.7035 7.1460 40.7970 ;
        RECT 7.0120 39.7035 7.0380 40.7970 ;
        RECT 6.9040 39.7035 6.9300 40.7970 ;
        RECT 6.7960 39.7035 6.8220 40.7970 ;
        RECT 6.6880 39.7035 6.7140 40.7970 ;
        RECT 6.5800 39.7035 6.6060 40.7970 ;
        RECT 6.4720 39.7035 6.4980 40.7970 ;
        RECT 6.3640 39.7035 6.3900 40.7970 ;
        RECT 6.2560 39.7035 6.2820 40.7970 ;
        RECT 6.1480 39.7035 6.1740 40.7970 ;
        RECT 6.0400 39.7035 6.0660 40.7970 ;
        RECT 5.9320 39.7035 5.9580 40.7970 ;
        RECT 5.8240 39.7035 5.8500 40.7970 ;
        RECT 5.7160 39.7035 5.7420 40.7970 ;
        RECT 5.6080 39.7035 5.6340 40.7970 ;
        RECT 5.5000 39.7035 5.5260 40.7970 ;
        RECT 5.3920 39.7035 5.4180 40.7970 ;
        RECT 5.2840 39.7035 5.3100 40.7970 ;
        RECT 5.1760 39.7035 5.2020 40.7970 ;
        RECT 5.0680 39.7035 5.0940 40.7970 ;
        RECT 4.9600 39.7035 4.9860 40.7970 ;
        RECT 4.8520 39.7035 4.8780 40.7970 ;
        RECT 4.7440 39.7035 4.7700 40.7970 ;
        RECT 4.6360 39.7035 4.6620 40.7970 ;
        RECT 4.5280 39.7035 4.5540 40.7970 ;
        RECT 4.4200 39.7035 4.4460 40.7970 ;
        RECT 4.3120 39.7035 4.3380 40.7970 ;
        RECT 4.2040 39.7035 4.2300 40.7970 ;
        RECT 4.0960 39.7035 4.1220 40.7970 ;
        RECT 3.9880 39.7035 4.0140 40.7970 ;
        RECT 3.8800 39.7035 3.9060 40.7970 ;
        RECT 3.7720 39.7035 3.7980 40.7970 ;
        RECT 3.6640 39.7035 3.6900 40.7970 ;
        RECT 3.5560 39.7035 3.5820 40.7970 ;
        RECT 3.4480 39.7035 3.4740 40.7970 ;
        RECT 3.3400 39.7035 3.3660 40.7970 ;
        RECT 3.2320 39.7035 3.2580 40.7970 ;
        RECT 3.1240 39.7035 3.1500 40.7970 ;
        RECT 3.0160 39.7035 3.0420 40.7970 ;
        RECT 2.9080 39.7035 2.9340 40.7970 ;
        RECT 2.8000 39.7035 2.8260 40.7970 ;
        RECT 2.6920 39.7035 2.7180 40.7970 ;
        RECT 2.5840 39.7035 2.6100 40.7970 ;
        RECT 2.4760 39.7035 2.5020 40.7970 ;
        RECT 2.3680 39.7035 2.3940 40.7970 ;
        RECT 2.2600 39.7035 2.2860 40.7970 ;
        RECT 2.1520 39.7035 2.1780 40.7970 ;
        RECT 2.0440 39.7035 2.0700 40.7970 ;
        RECT 1.9360 39.7035 1.9620 40.7970 ;
        RECT 1.8280 39.7035 1.8540 40.7970 ;
        RECT 1.7200 39.7035 1.7460 40.7970 ;
        RECT 1.6120 39.7035 1.6380 40.7970 ;
        RECT 1.5040 39.7035 1.5300 40.7970 ;
        RECT 1.3960 39.7035 1.4220 40.7970 ;
        RECT 1.2880 39.7035 1.3140 40.7970 ;
        RECT 1.1800 39.7035 1.2060 40.7970 ;
        RECT 1.0720 39.7035 1.0980 40.7970 ;
        RECT 0.9640 39.7035 0.9900 40.7970 ;
        RECT 0.8560 39.7035 0.8820 40.7970 ;
        RECT 0.7480 39.7035 0.7740 40.7970 ;
        RECT 0.6400 39.7035 0.6660 40.7970 ;
        RECT 0.5320 39.7035 0.5580 40.7970 ;
        RECT 0.4240 39.7035 0.4500 40.7970 ;
        RECT 0.3160 39.7035 0.3420 40.7970 ;
        RECT 0.2080 39.7035 0.2340 40.7970 ;
        RECT 0.0050 39.7035 0.0900 40.7970 ;
        RECT 15.5530 40.7835 15.6810 41.8770 ;
        RECT 15.5390 41.4490 15.6810 41.7715 ;
        RECT 15.3190 41.1760 15.4530 41.8770 ;
        RECT 15.2960 41.5110 15.4530 41.7690 ;
        RECT 15.3190 40.7835 15.4170 41.8770 ;
        RECT 15.3190 40.9045 15.4310 41.1440 ;
        RECT 15.3190 40.7835 15.4530 40.8725 ;
        RECT 15.0940 41.2340 15.2280 41.8770 ;
        RECT 15.0940 40.7835 15.1920 41.8770 ;
        RECT 14.6770 40.7835 14.7600 41.8770 ;
        RECT 14.6770 40.8720 14.7740 41.8075 ;
        RECT 30.2680 40.7835 30.3530 41.8770 ;
        RECT 30.1240 40.7835 30.1500 41.8770 ;
        RECT 30.0160 40.7835 30.0420 41.8770 ;
        RECT 29.9080 40.7835 29.9340 41.8770 ;
        RECT 29.8000 40.7835 29.8260 41.8770 ;
        RECT 29.6920 40.7835 29.7180 41.8770 ;
        RECT 29.5840 40.7835 29.6100 41.8770 ;
        RECT 29.4760 40.7835 29.5020 41.8770 ;
        RECT 29.3680 40.7835 29.3940 41.8770 ;
        RECT 29.2600 40.7835 29.2860 41.8770 ;
        RECT 29.1520 40.7835 29.1780 41.8770 ;
        RECT 29.0440 40.7835 29.0700 41.8770 ;
        RECT 28.9360 40.7835 28.9620 41.8770 ;
        RECT 28.8280 40.7835 28.8540 41.8770 ;
        RECT 28.7200 40.7835 28.7460 41.8770 ;
        RECT 28.6120 40.7835 28.6380 41.8770 ;
        RECT 28.5040 40.7835 28.5300 41.8770 ;
        RECT 28.3960 40.7835 28.4220 41.8770 ;
        RECT 28.2880 40.7835 28.3140 41.8770 ;
        RECT 28.1800 40.7835 28.2060 41.8770 ;
        RECT 28.0720 40.7835 28.0980 41.8770 ;
        RECT 27.9640 40.7835 27.9900 41.8770 ;
        RECT 27.8560 40.7835 27.8820 41.8770 ;
        RECT 27.7480 40.7835 27.7740 41.8770 ;
        RECT 27.6400 40.7835 27.6660 41.8770 ;
        RECT 27.5320 40.7835 27.5580 41.8770 ;
        RECT 27.4240 40.7835 27.4500 41.8770 ;
        RECT 27.3160 40.7835 27.3420 41.8770 ;
        RECT 27.2080 40.7835 27.2340 41.8770 ;
        RECT 27.1000 40.7835 27.1260 41.8770 ;
        RECT 26.9920 40.7835 27.0180 41.8770 ;
        RECT 26.8840 40.7835 26.9100 41.8770 ;
        RECT 26.7760 40.7835 26.8020 41.8770 ;
        RECT 26.6680 40.7835 26.6940 41.8770 ;
        RECT 26.5600 40.7835 26.5860 41.8770 ;
        RECT 26.4520 40.7835 26.4780 41.8770 ;
        RECT 26.3440 40.7835 26.3700 41.8770 ;
        RECT 26.2360 40.7835 26.2620 41.8770 ;
        RECT 26.1280 40.7835 26.1540 41.8770 ;
        RECT 26.0200 40.7835 26.0460 41.8770 ;
        RECT 25.9120 40.7835 25.9380 41.8770 ;
        RECT 25.8040 40.7835 25.8300 41.8770 ;
        RECT 25.6960 40.7835 25.7220 41.8770 ;
        RECT 25.5880 40.7835 25.6140 41.8770 ;
        RECT 25.4800 40.7835 25.5060 41.8770 ;
        RECT 25.3720 40.7835 25.3980 41.8770 ;
        RECT 25.2640 40.7835 25.2900 41.8770 ;
        RECT 25.1560 40.7835 25.1820 41.8770 ;
        RECT 25.0480 40.7835 25.0740 41.8770 ;
        RECT 24.9400 40.7835 24.9660 41.8770 ;
        RECT 24.8320 40.7835 24.8580 41.8770 ;
        RECT 24.7240 40.7835 24.7500 41.8770 ;
        RECT 24.6160 40.7835 24.6420 41.8770 ;
        RECT 24.5080 40.7835 24.5340 41.8770 ;
        RECT 24.4000 40.7835 24.4260 41.8770 ;
        RECT 24.2920 40.7835 24.3180 41.8770 ;
        RECT 24.1840 40.7835 24.2100 41.8770 ;
        RECT 24.0760 40.7835 24.1020 41.8770 ;
        RECT 23.9680 40.7835 23.9940 41.8770 ;
        RECT 23.8600 40.7835 23.8860 41.8770 ;
        RECT 23.7520 40.7835 23.7780 41.8770 ;
        RECT 23.6440 40.7835 23.6700 41.8770 ;
        RECT 23.5360 40.7835 23.5620 41.8770 ;
        RECT 23.4280 40.7835 23.4540 41.8770 ;
        RECT 23.3200 40.7835 23.3460 41.8770 ;
        RECT 23.2120 40.7835 23.2380 41.8770 ;
        RECT 23.1040 40.7835 23.1300 41.8770 ;
        RECT 22.9960 40.7835 23.0220 41.8770 ;
        RECT 22.8880 40.7835 22.9140 41.8770 ;
        RECT 22.7800 40.7835 22.8060 41.8770 ;
        RECT 22.6720 40.7835 22.6980 41.8770 ;
        RECT 22.5640 40.7835 22.5900 41.8770 ;
        RECT 22.4560 40.7835 22.4820 41.8770 ;
        RECT 22.3480 40.7835 22.3740 41.8770 ;
        RECT 22.2400 40.7835 22.2660 41.8770 ;
        RECT 22.1320 40.7835 22.1580 41.8770 ;
        RECT 22.0240 40.7835 22.0500 41.8770 ;
        RECT 21.9160 40.7835 21.9420 41.8770 ;
        RECT 21.8080 40.7835 21.8340 41.8770 ;
        RECT 21.7000 40.7835 21.7260 41.8770 ;
        RECT 21.5920 40.7835 21.6180 41.8770 ;
        RECT 21.4840 40.7835 21.5100 41.8770 ;
        RECT 21.3760 40.7835 21.4020 41.8770 ;
        RECT 21.2680 40.7835 21.2940 41.8770 ;
        RECT 21.1600 40.7835 21.1860 41.8770 ;
        RECT 21.0520 40.7835 21.0780 41.8770 ;
        RECT 20.9440 40.7835 20.9700 41.8770 ;
        RECT 20.8360 40.7835 20.8620 41.8770 ;
        RECT 20.7280 40.7835 20.7540 41.8770 ;
        RECT 20.6200 40.7835 20.6460 41.8770 ;
        RECT 20.5120 40.7835 20.5380 41.8770 ;
        RECT 20.4040 40.7835 20.4300 41.8770 ;
        RECT 20.2960 40.7835 20.3220 41.8770 ;
        RECT 20.1880 40.7835 20.2140 41.8770 ;
        RECT 20.0800 40.7835 20.1060 41.8770 ;
        RECT 19.9720 40.7835 19.9980 41.8770 ;
        RECT 19.8640 40.7835 19.8900 41.8770 ;
        RECT 19.7560 40.7835 19.7820 41.8770 ;
        RECT 19.6480 40.7835 19.6740 41.8770 ;
        RECT 19.5400 40.7835 19.5660 41.8770 ;
        RECT 19.4320 40.7835 19.4580 41.8770 ;
        RECT 19.3240 40.7835 19.3500 41.8770 ;
        RECT 19.2160 40.7835 19.2420 41.8770 ;
        RECT 19.1080 40.7835 19.1340 41.8770 ;
        RECT 19.0000 40.7835 19.0260 41.8770 ;
        RECT 18.8920 40.7835 18.9180 41.8770 ;
        RECT 18.7840 40.7835 18.8100 41.8770 ;
        RECT 18.6760 40.7835 18.7020 41.8770 ;
        RECT 18.5680 40.7835 18.5940 41.8770 ;
        RECT 18.4600 40.7835 18.4860 41.8770 ;
        RECT 18.3520 40.7835 18.3780 41.8770 ;
        RECT 18.2440 40.7835 18.2700 41.8770 ;
        RECT 18.1360 40.7835 18.1620 41.8770 ;
        RECT 18.0280 40.7835 18.0540 41.8770 ;
        RECT 17.9200 40.7835 17.9460 41.8770 ;
        RECT 17.8120 40.7835 17.8380 41.8770 ;
        RECT 17.7040 40.7835 17.7300 41.8770 ;
        RECT 17.5960 40.7835 17.6220 41.8770 ;
        RECT 17.4880 40.7835 17.5140 41.8770 ;
        RECT 17.3800 40.7835 17.4060 41.8770 ;
        RECT 17.2720 40.7835 17.2980 41.8770 ;
        RECT 17.1640 40.7835 17.1900 41.8770 ;
        RECT 17.0560 40.7835 17.0820 41.8770 ;
        RECT 16.9480 40.7835 16.9740 41.8770 ;
        RECT 16.8400 40.7835 16.8660 41.8770 ;
        RECT 16.7320 40.7835 16.7580 41.8770 ;
        RECT 16.6240 40.7835 16.6500 41.8770 ;
        RECT 16.5160 40.7835 16.5420 41.8770 ;
        RECT 16.4080 40.7835 16.4340 41.8770 ;
        RECT 16.3000 40.7835 16.3260 41.8770 ;
        RECT 16.0870 40.7835 16.1640 41.8770 ;
        RECT 14.1940 40.7835 14.2710 41.8770 ;
        RECT 14.0320 40.7835 14.0580 41.8770 ;
        RECT 13.9240 40.7835 13.9500 41.8770 ;
        RECT 13.8160 40.7835 13.8420 41.8770 ;
        RECT 13.7080 40.7835 13.7340 41.8770 ;
        RECT 13.6000 40.7835 13.6260 41.8770 ;
        RECT 13.4920 40.7835 13.5180 41.8770 ;
        RECT 13.3840 40.7835 13.4100 41.8770 ;
        RECT 13.2760 40.7835 13.3020 41.8770 ;
        RECT 13.1680 40.7835 13.1940 41.8770 ;
        RECT 13.0600 40.7835 13.0860 41.8770 ;
        RECT 12.9520 40.7835 12.9780 41.8770 ;
        RECT 12.8440 40.7835 12.8700 41.8770 ;
        RECT 12.7360 40.7835 12.7620 41.8770 ;
        RECT 12.6280 40.7835 12.6540 41.8770 ;
        RECT 12.5200 40.7835 12.5460 41.8770 ;
        RECT 12.4120 40.7835 12.4380 41.8770 ;
        RECT 12.3040 40.7835 12.3300 41.8770 ;
        RECT 12.1960 40.7835 12.2220 41.8770 ;
        RECT 12.0880 40.7835 12.1140 41.8770 ;
        RECT 11.9800 40.7835 12.0060 41.8770 ;
        RECT 11.8720 40.7835 11.8980 41.8770 ;
        RECT 11.7640 40.7835 11.7900 41.8770 ;
        RECT 11.6560 40.7835 11.6820 41.8770 ;
        RECT 11.5480 40.7835 11.5740 41.8770 ;
        RECT 11.4400 40.7835 11.4660 41.8770 ;
        RECT 11.3320 40.7835 11.3580 41.8770 ;
        RECT 11.2240 40.7835 11.2500 41.8770 ;
        RECT 11.1160 40.7835 11.1420 41.8770 ;
        RECT 11.0080 40.7835 11.0340 41.8770 ;
        RECT 10.9000 40.7835 10.9260 41.8770 ;
        RECT 10.7920 40.7835 10.8180 41.8770 ;
        RECT 10.6840 40.7835 10.7100 41.8770 ;
        RECT 10.5760 40.7835 10.6020 41.8770 ;
        RECT 10.4680 40.7835 10.4940 41.8770 ;
        RECT 10.3600 40.7835 10.3860 41.8770 ;
        RECT 10.2520 40.7835 10.2780 41.8770 ;
        RECT 10.1440 40.7835 10.1700 41.8770 ;
        RECT 10.0360 40.7835 10.0620 41.8770 ;
        RECT 9.9280 40.7835 9.9540 41.8770 ;
        RECT 9.8200 40.7835 9.8460 41.8770 ;
        RECT 9.7120 40.7835 9.7380 41.8770 ;
        RECT 9.6040 40.7835 9.6300 41.8770 ;
        RECT 9.4960 40.7835 9.5220 41.8770 ;
        RECT 9.3880 40.7835 9.4140 41.8770 ;
        RECT 9.2800 40.7835 9.3060 41.8770 ;
        RECT 9.1720 40.7835 9.1980 41.8770 ;
        RECT 9.0640 40.7835 9.0900 41.8770 ;
        RECT 8.9560 40.7835 8.9820 41.8770 ;
        RECT 8.8480 40.7835 8.8740 41.8770 ;
        RECT 8.7400 40.7835 8.7660 41.8770 ;
        RECT 8.6320 40.7835 8.6580 41.8770 ;
        RECT 8.5240 40.7835 8.5500 41.8770 ;
        RECT 8.4160 40.7835 8.4420 41.8770 ;
        RECT 8.3080 40.7835 8.3340 41.8770 ;
        RECT 8.2000 40.7835 8.2260 41.8770 ;
        RECT 8.0920 40.7835 8.1180 41.8770 ;
        RECT 7.9840 40.7835 8.0100 41.8770 ;
        RECT 7.8760 40.7835 7.9020 41.8770 ;
        RECT 7.7680 40.7835 7.7940 41.8770 ;
        RECT 7.6600 40.7835 7.6860 41.8770 ;
        RECT 7.5520 40.7835 7.5780 41.8770 ;
        RECT 7.4440 40.7835 7.4700 41.8770 ;
        RECT 7.3360 40.7835 7.3620 41.8770 ;
        RECT 7.2280 40.7835 7.2540 41.8770 ;
        RECT 7.1200 40.7835 7.1460 41.8770 ;
        RECT 7.0120 40.7835 7.0380 41.8770 ;
        RECT 6.9040 40.7835 6.9300 41.8770 ;
        RECT 6.7960 40.7835 6.8220 41.8770 ;
        RECT 6.6880 40.7835 6.7140 41.8770 ;
        RECT 6.5800 40.7835 6.6060 41.8770 ;
        RECT 6.4720 40.7835 6.4980 41.8770 ;
        RECT 6.3640 40.7835 6.3900 41.8770 ;
        RECT 6.2560 40.7835 6.2820 41.8770 ;
        RECT 6.1480 40.7835 6.1740 41.8770 ;
        RECT 6.0400 40.7835 6.0660 41.8770 ;
        RECT 5.9320 40.7835 5.9580 41.8770 ;
        RECT 5.8240 40.7835 5.8500 41.8770 ;
        RECT 5.7160 40.7835 5.7420 41.8770 ;
        RECT 5.6080 40.7835 5.6340 41.8770 ;
        RECT 5.5000 40.7835 5.5260 41.8770 ;
        RECT 5.3920 40.7835 5.4180 41.8770 ;
        RECT 5.2840 40.7835 5.3100 41.8770 ;
        RECT 5.1760 40.7835 5.2020 41.8770 ;
        RECT 5.0680 40.7835 5.0940 41.8770 ;
        RECT 4.9600 40.7835 4.9860 41.8770 ;
        RECT 4.8520 40.7835 4.8780 41.8770 ;
        RECT 4.7440 40.7835 4.7700 41.8770 ;
        RECT 4.6360 40.7835 4.6620 41.8770 ;
        RECT 4.5280 40.7835 4.5540 41.8770 ;
        RECT 4.4200 40.7835 4.4460 41.8770 ;
        RECT 4.3120 40.7835 4.3380 41.8770 ;
        RECT 4.2040 40.7835 4.2300 41.8770 ;
        RECT 4.0960 40.7835 4.1220 41.8770 ;
        RECT 3.9880 40.7835 4.0140 41.8770 ;
        RECT 3.8800 40.7835 3.9060 41.8770 ;
        RECT 3.7720 40.7835 3.7980 41.8770 ;
        RECT 3.6640 40.7835 3.6900 41.8770 ;
        RECT 3.5560 40.7835 3.5820 41.8770 ;
        RECT 3.4480 40.7835 3.4740 41.8770 ;
        RECT 3.3400 40.7835 3.3660 41.8770 ;
        RECT 3.2320 40.7835 3.2580 41.8770 ;
        RECT 3.1240 40.7835 3.1500 41.8770 ;
        RECT 3.0160 40.7835 3.0420 41.8770 ;
        RECT 2.9080 40.7835 2.9340 41.8770 ;
        RECT 2.8000 40.7835 2.8260 41.8770 ;
        RECT 2.6920 40.7835 2.7180 41.8770 ;
        RECT 2.5840 40.7835 2.6100 41.8770 ;
        RECT 2.4760 40.7835 2.5020 41.8770 ;
        RECT 2.3680 40.7835 2.3940 41.8770 ;
        RECT 2.2600 40.7835 2.2860 41.8770 ;
        RECT 2.1520 40.7835 2.1780 41.8770 ;
        RECT 2.0440 40.7835 2.0700 41.8770 ;
        RECT 1.9360 40.7835 1.9620 41.8770 ;
        RECT 1.8280 40.7835 1.8540 41.8770 ;
        RECT 1.7200 40.7835 1.7460 41.8770 ;
        RECT 1.6120 40.7835 1.6380 41.8770 ;
        RECT 1.5040 40.7835 1.5300 41.8770 ;
        RECT 1.3960 40.7835 1.4220 41.8770 ;
        RECT 1.2880 40.7835 1.3140 41.8770 ;
        RECT 1.1800 40.7835 1.2060 41.8770 ;
        RECT 1.0720 40.7835 1.0980 41.8770 ;
        RECT 0.9640 40.7835 0.9900 41.8770 ;
        RECT 0.8560 40.7835 0.8820 41.8770 ;
        RECT 0.7480 40.7835 0.7740 41.8770 ;
        RECT 0.6400 40.7835 0.6660 41.8770 ;
        RECT 0.5320 40.7835 0.5580 41.8770 ;
        RECT 0.4240 40.7835 0.4500 41.8770 ;
        RECT 0.3160 40.7835 0.3420 41.8770 ;
        RECT 0.2080 40.7835 0.2340 41.8770 ;
        RECT 0.0050 40.7835 0.0900 41.8770 ;
        RECT 15.5530 41.8635 15.6810 42.9570 ;
        RECT 15.5390 42.5290 15.6810 42.8515 ;
        RECT 15.3190 42.2560 15.4530 42.9570 ;
        RECT 15.2960 42.5910 15.4530 42.8490 ;
        RECT 15.3190 41.8635 15.4170 42.9570 ;
        RECT 15.3190 41.9845 15.4310 42.2240 ;
        RECT 15.3190 41.8635 15.4530 41.9525 ;
        RECT 15.0940 42.3140 15.2280 42.9570 ;
        RECT 15.0940 41.8635 15.1920 42.9570 ;
        RECT 14.6770 41.8635 14.7600 42.9570 ;
        RECT 14.6770 41.9520 14.7740 42.8875 ;
        RECT 30.2680 41.8635 30.3530 42.9570 ;
        RECT 30.1240 41.8635 30.1500 42.9570 ;
        RECT 30.0160 41.8635 30.0420 42.9570 ;
        RECT 29.9080 41.8635 29.9340 42.9570 ;
        RECT 29.8000 41.8635 29.8260 42.9570 ;
        RECT 29.6920 41.8635 29.7180 42.9570 ;
        RECT 29.5840 41.8635 29.6100 42.9570 ;
        RECT 29.4760 41.8635 29.5020 42.9570 ;
        RECT 29.3680 41.8635 29.3940 42.9570 ;
        RECT 29.2600 41.8635 29.2860 42.9570 ;
        RECT 29.1520 41.8635 29.1780 42.9570 ;
        RECT 29.0440 41.8635 29.0700 42.9570 ;
        RECT 28.9360 41.8635 28.9620 42.9570 ;
        RECT 28.8280 41.8635 28.8540 42.9570 ;
        RECT 28.7200 41.8635 28.7460 42.9570 ;
        RECT 28.6120 41.8635 28.6380 42.9570 ;
        RECT 28.5040 41.8635 28.5300 42.9570 ;
        RECT 28.3960 41.8635 28.4220 42.9570 ;
        RECT 28.2880 41.8635 28.3140 42.9570 ;
        RECT 28.1800 41.8635 28.2060 42.9570 ;
        RECT 28.0720 41.8635 28.0980 42.9570 ;
        RECT 27.9640 41.8635 27.9900 42.9570 ;
        RECT 27.8560 41.8635 27.8820 42.9570 ;
        RECT 27.7480 41.8635 27.7740 42.9570 ;
        RECT 27.6400 41.8635 27.6660 42.9570 ;
        RECT 27.5320 41.8635 27.5580 42.9570 ;
        RECT 27.4240 41.8635 27.4500 42.9570 ;
        RECT 27.3160 41.8635 27.3420 42.9570 ;
        RECT 27.2080 41.8635 27.2340 42.9570 ;
        RECT 27.1000 41.8635 27.1260 42.9570 ;
        RECT 26.9920 41.8635 27.0180 42.9570 ;
        RECT 26.8840 41.8635 26.9100 42.9570 ;
        RECT 26.7760 41.8635 26.8020 42.9570 ;
        RECT 26.6680 41.8635 26.6940 42.9570 ;
        RECT 26.5600 41.8635 26.5860 42.9570 ;
        RECT 26.4520 41.8635 26.4780 42.9570 ;
        RECT 26.3440 41.8635 26.3700 42.9570 ;
        RECT 26.2360 41.8635 26.2620 42.9570 ;
        RECT 26.1280 41.8635 26.1540 42.9570 ;
        RECT 26.0200 41.8635 26.0460 42.9570 ;
        RECT 25.9120 41.8635 25.9380 42.9570 ;
        RECT 25.8040 41.8635 25.8300 42.9570 ;
        RECT 25.6960 41.8635 25.7220 42.9570 ;
        RECT 25.5880 41.8635 25.6140 42.9570 ;
        RECT 25.4800 41.8635 25.5060 42.9570 ;
        RECT 25.3720 41.8635 25.3980 42.9570 ;
        RECT 25.2640 41.8635 25.2900 42.9570 ;
        RECT 25.1560 41.8635 25.1820 42.9570 ;
        RECT 25.0480 41.8635 25.0740 42.9570 ;
        RECT 24.9400 41.8635 24.9660 42.9570 ;
        RECT 24.8320 41.8635 24.8580 42.9570 ;
        RECT 24.7240 41.8635 24.7500 42.9570 ;
        RECT 24.6160 41.8635 24.6420 42.9570 ;
        RECT 24.5080 41.8635 24.5340 42.9570 ;
        RECT 24.4000 41.8635 24.4260 42.9570 ;
        RECT 24.2920 41.8635 24.3180 42.9570 ;
        RECT 24.1840 41.8635 24.2100 42.9570 ;
        RECT 24.0760 41.8635 24.1020 42.9570 ;
        RECT 23.9680 41.8635 23.9940 42.9570 ;
        RECT 23.8600 41.8635 23.8860 42.9570 ;
        RECT 23.7520 41.8635 23.7780 42.9570 ;
        RECT 23.6440 41.8635 23.6700 42.9570 ;
        RECT 23.5360 41.8635 23.5620 42.9570 ;
        RECT 23.4280 41.8635 23.4540 42.9570 ;
        RECT 23.3200 41.8635 23.3460 42.9570 ;
        RECT 23.2120 41.8635 23.2380 42.9570 ;
        RECT 23.1040 41.8635 23.1300 42.9570 ;
        RECT 22.9960 41.8635 23.0220 42.9570 ;
        RECT 22.8880 41.8635 22.9140 42.9570 ;
        RECT 22.7800 41.8635 22.8060 42.9570 ;
        RECT 22.6720 41.8635 22.6980 42.9570 ;
        RECT 22.5640 41.8635 22.5900 42.9570 ;
        RECT 22.4560 41.8635 22.4820 42.9570 ;
        RECT 22.3480 41.8635 22.3740 42.9570 ;
        RECT 22.2400 41.8635 22.2660 42.9570 ;
        RECT 22.1320 41.8635 22.1580 42.9570 ;
        RECT 22.0240 41.8635 22.0500 42.9570 ;
        RECT 21.9160 41.8635 21.9420 42.9570 ;
        RECT 21.8080 41.8635 21.8340 42.9570 ;
        RECT 21.7000 41.8635 21.7260 42.9570 ;
        RECT 21.5920 41.8635 21.6180 42.9570 ;
        RECT 21.4840 41.8635 21.5100 42.9570 ;
        RECT 21.3760 41.8635 21.4020 42.9570 ;
        RECT 21.2680 41.8635 21.2940 42.9570 ;
        RECT 21.1600 41.8635 21.1860 42.9570 ;
        RECT 21.0520 41.8635 21.0780 42.9570 ;
        RECT 20.9440 41.8635 20.9700 42.9570 ;
        RECT 20.8360 41.8635 20.8620 42.9570 ;
        RECT 20.7280 41.8635 20.7540 42.9570 ;
        RECT 20.6200 41.8635 20.6460 42.9570 ;
        RECT 20.5120 41.8635 20.5380 42.9570 ;
        RECT 20.4040 41.8635 20.4300 42.9570 ;
        RECT 20.2960 41.8635 20.3220 42.9570 ;
        RECT 20.1880 41.8635 20.2140 42.9570 ;
        RECT 20.0800 41.8635 20.1060 42.9570 ;
        RECT 19.9720 41.8635 19.9980 42.9570 ;
        RECT 19.8640 41.8635 19.8900 42.9570 ;
        RECT 19.7560 41.8635 19.7820 42.9570 ;
        RECT 19.6480 41.8635 19.6740 42.9570 ;
        RECT 19.5400 41.8635 19.5660 42.9570 ;
        RECT 19.4320 41.8635 19.4580 42.9570 ;
        RECT 19.3240 41.8635 19.3500 42.9570 ;
        RECT 19.2160 41.8635 19.2420 42.9570 ;
        RECT 19.1080 41.8635 19.1340 42.9570 ;
        RECT 19.0000 41.8635 19.0260 42.9570 ;
        RECT 18.8920 41.8635 18.9180 42.9570 ;
        RECT 18.7840 41.8635 18.8100 42.9570 ;
        RECT 18.6760 41.8635 18.7020 42.9570 ;
        RECT 18.5680 41.8635 18.5940 42.9570 ;
        RECT 18.4600 41.8635 18.4860 42.9570 ;
        RECT 18.3520 41.8635 18.3780 42.9570 ;
        RECT 18.2440 41.8635 18.2700 42.9570 ;
        RECT 18.1360 41.8635 18.1620 42.9570 ;
        RECT 18.0280 41.8635 18.0540 42.9570 ;
        RECT 17.9200 41.8635 17.9460 42.9570 ;
        RECT 17.8120 41.8635 17.8380 42.9570 ;
        RECT 17.7040 41.8635 17.7300 42.9570 ;
        RECT 17.5960 41.8635 17.6220 42.9570 ;
        RECT 17.4880 41.8635 17.5140 42.9570 ;
        RECT 17.3800 41.8635 17.4060 42.9570 ;
        RECT 17.2720 41.8635 17.2980 42.9570 ;
        RECT 17.1640 41.8635 17.1900 42.9570 ;
        RECT 17.0560 41.8635 17.0820 42.9570 ;
        RECT 16.9480 41.8635 16.9740 42.9570 ;
        RECT 16.8400 41.8635 16.8660 42.9570 ;
        RECT 16.7320 41.8635 16.7580 42.9570 ;
        RECT 16.6240 41.8635 16.6500 42.9570 ;
        RECT 16.5160 41.8635 16.5420 42.9570 ;
        RECT 16.4080 41.8635 16.4340 42.9570 ;
        RECT 16.3000 41.8635 16.3260 42.9570 ;
        RECT 16.0870 41.8635 16.1640 42.9570 ;
        RECT 14.1940 41.8635 14.2710 42.9570 ;
        RECT 14.0320 41.8635 14.0580 42.9570 ;
        RECT 13.9240 41.8635 13.9500 42.9570 ;
        RECT 13.8160 41.8635 13.8420 42.9570 ;
        RECT 13.7080 41.8635 13.7340 42.9570 ;
        RECT 13.6000 41.8635 13.6260 42.9570 ;
        RECT 13.4920 41.8635 13.5180 42.9570 ;
        RECT 13.3840 41.8635 13.4100 42.9570 ;
        RECT 13.2760 41.8635 13.3020 42.9570 ;
        RECT 13.1680 41.8635 13.1940 42.9570 ;
        RECT 13.0600 41.8635 13.0860 42.9570 ;
        RECT 12.9520 41.8635 12.9780 42.9570 ;
        RECT 12.8440 41.8635 12.8700 42.9570 ;
        RECT 12.7360 41.8635 12.7620 42.9570 ;
        RECT 12.6280 41.8635 12.6540 42.9570 ;
        RECT 12.5200 41.8635 12.5460 42.9570 ;
        RECT 12.4120 41.8635 12.4380 42.9570 ;
        RECT 12.3040 41.8635 12.3300 42.9570 ;
        RECT 12.1960 41.8635 12.2220 42.9570 ;
        RECT 12.0880 41.8635 12.1140 42.9570 ;
        RECT 11.9800 41.8635 12.0060 42.9570 ;
        RECT 11.8720 41.8635 11.8980 42.9570 ;
        RECT 11.7640 41.8635 11.7900 42.9570 ;
        RECT 11.6560 41.8635 11.6820 42.9570 ;
        RECT 11.5480 41.8635 11.5740 42.9570 ;
        RECT 11.4400 41.8635 11.4660 42.9570 ;
        RECT 11.3320 41.8635 11.3580 42.9570 ;
        RECT 11.2240 41.8635 11.2500 42.9570 ;
        RECT 11.1160 41.8635 11.1420 42.9570 ;
        RECT 11.0080 41.8635 11.0340 42.9570 ;
        RECT 10.9000 41.8635 10.9260 42.9570 ;
        RECT 10.7920 41.8635 10.8180 42.9570 ;
        RECT 10.6840 41.8635 10.7100 42.9570 ;
        RECT 10.5760 41.8635 10.6020 42.9570 ;
        RECT 10.4680 41.8635 10.4940 42.9570 ;
        RECT 10.3600 41.8635 10.3860 42.9570 ;
        RECT 10.2520 41.8635 10.2780 42.9570 ;
        RECT 10.1440 41.8635 10.1700 42.9570 ;
        RECT 10.0360 41.8635 10.0620 42.9570 ;
        RECT 9.9280 41.8635 9.9540 42.9570 ;
        RECT 9.8200 41.8635 9.8460 42.9570 ;
        RECT 9.7120 41.8635 9.7380 42.9570 ;
        RECT 9.6040 41.8635 9.6300 42.9570 ;
        RECT 9.4960 41.8635 9.5220 42.9570 ;
        RECT 9.3880 41.8635 9.4140 42.9570 ;
        RECT 9.2800 41.8635 9.3060 42.9570 ;
        RECT 9.1720 41.8635 9.1980 42.9570 ;
        RECT 9.0640 41.8635 9.0900 42.9570 ;
        RECT 8.9560 41.8635 8.9820 42.9570 ;
        RECT 8.8480 41.8635 8.8740 42.9570 ;
        RECT 8.7400 41.8635 8.7660 42.9570 ;
        RECT 8.6320 41.8635 8.6580 42.9570 ;
        RECT 8.5240 41.8635 8.5500 42.9570 ;
        RECT 8.4160 41.8635 8.4420 42.9570 ;
        RECT 8.3080 41.8635 8.3340 42.9570 ;
        RECT 8.2000 41.8635 8.2260 42.9570 ;
        RECT 8.0920 41.8635 8.1180 42.9570 ;
        RECT 7.9840 41.8635 8.0100 42.9570 ;
        RECT 7.8760 41.8635 7.9020 42.9570 ;
        RECT 7.7680 41.8635 7.7940 42.9570 ;
        RECT 7.6600 41.8635 7.6860 42.9570 ;
        RECT 7.5520 41.8635 7.5780 42.9570 ;
        RECT 7.4440 41.8635 7.4700 42.9570 ;
        RECT 7.3360 41.8635 7.3620 42.9570 ;
        RECT 7.2280 41.8635 7.2540 42.9570 ;
        RECT 7.1200 41.8635 7.1460 42.9570 ;
        RECT 7.0120 41.8635 7.0380 42.9570 ;
        RECT 6.9040 41.8635 6.9300 42.9570 ;
        RECT 6.7960 41.8635 6.8220 42.9570 ;
        RECT 6.6880 41.8635 6.7140 42.9570 ;
        RECT 6.5800 41.8635 6.6060 42.9570 ;
        RECT 6.4720 41.8635 6.4980 42.9570 ;
        RECT 6.3640 41.8635 6.3900 42.9570 ;
        RECT 6.2560 41.8635 6.2820 42.9570 ;
        RECT 6.1480 41.8635 6.1740 42.9570 ;
        RECT 6.0400 41.8635 6.0660 42.9570 ;
        RECT 5.9320 41.8635 5.9580 42.9570 ;
        RECT 5.8240 41.8635 5.8500 42.9570 ;
        RECT 5.7160 41.8635 5.7420 42.9570 ;
        RECT 5.6080 41.8635 5.6340 42.9570 ;
        RECT 5.5000 41.8635 5.5260 42.9570 ;
        RECT 5.3920 41.8635 5.4180 42.9570 ;
        RECT 5.2840 41.8635 5.3100 42.9570 ;
        RECT 5.1760 41.8635 5.2020 42.9570 ;
        RECT 5.0680 41.8635 5.0940 42.9570 ;
        RECT 4.9600 41.8635 4.9860 42.9570 ;
        RECT 4.8520 41.8635 4.8780 42.9570 ;
        RECT 4.7440 41.8635 4.7700 42.9570 ;
        RECT 4.6360 41.8635 4.6620 42.9570 ;
        RECT 4.5280 41.8635 4.5540 42.9570 ;
        RECT 4.4200 41.8635 4.4460 42.9570 ;
        RECT 4.3120 41.8635 4.3380 42.9570 ;
        RECT 4.2040 41.8635 4.2300 42.9570 ;
        RECT 4.0960 41.8635 4.1220 42.9570 ;
        RECT 3.9880 41.8635 4.0140 42.9570 ;
        RECT 3.8800 41.8635 3.9060 42.9570 ;
        RECT 3.7720 41.8635 3.7980 42.9570 ;
        RECT 3.6640 41.8635 3.6900 42.9570 ;
        RECT 3.5560 41.8635 3.5820 42.9570 ;
        RECT 3.4480 41.8635 3.4740 42.9570 ;
        RECT 3.3400 41.8635 3.3660 42.9570 ;
        RECT 3.2320 41.8635 3.2580 42.9570 ;
        RECT 3.1240 41.8635 3.1500 42.9570 ;
        RECT 3.0160 41.8635 3.0420 42.9570 ;
        RECT 2.9080 41.8635 2.9340 42.9570 ;
        RECT 2.8000 41.8635 2.8260 42.9570 ;
        RECT 2.6920 41.8635 2.7180 42.9570 ;
        RECT 2.5840 41.8635 2.6100 42.9570 ;
        RECT 2.4760 41.8635 2.5020 42.9570 ;
        RECT 2.3680 41.8635 2.3940 42.9570 ;
        RECT 2.2600 41.8635 2.2860 42.9570 ;
        RECT 2.1520 41.8635 2.1780 42.9570 ;
        RECT 2.0440 41.8635 2.0700 42.9570 ;
        RECT 1.9360 41.8635 1.9620 42.9570 ;
        RECT 1.8280 41.8635 1.8540 42.9570 ;
        RECT 1.7200 41.8635 1.7460 42.9570 ;
        RECT 1.6120 41.8635 1.6380 42.9570 ;
        RECT 1.5040 41.8635 1.5300 42.9570 ;
        RECT 1.3960 41.8635 1.4220 42.9570 ;
        RECT 1.2880 41.8635 1.3140 42.9570 ;
        RECT 1.1800 41.8635 1.2060 42.9570 ;
        RECT 1.0720 41.8635 1.0980 42.9570 ;
        RECT 0.9640 41.8635 0.9900 42.9570 ;
        RECT 0.8560 41.8635 0.8820 42.9570 ;
        RECT 0.7480 41.8635 0.7740 42.9570 ;
        RECT 0.6400 41.8635 0.6660 42.9570 ;
        RECT 0.5320 41.8635 0.5580 42.9570 ;
        RECT 0.4240 41.8635 0.4500 42.9570 ;
        RECT 0.3160 41.8635 0.3420 42.9570 ;
        RECT 0.2080 41.8635 0.2340 42.9570 ;
        RECT 0.0050 41.8635 0.0900 42.9570 ;
  LAYER V3 SPACING 0.018  ;
      RECT 0.0050 1.2200 30.3530 1.3500 ;
      RECT 30.2360 0.2565 30.3530 1.3500 ;
      RECT 16.2140 1.1240 30.2180 1.3500 ;
      RECT 14.8820 1.1240 16.1960 1.3500 ;
      RECT 14.1620 0.2565 14.7920 1.3500 ;
      RECT 0.1400 1.1240 14.1440 1.3500 ;
      RECT 0.0050 0.2565 0.1220 1.3500 ;
      RECT 30.2000 0.2565 30.3530 1.1720 ;
      RECT 16.2680 0.2565 30.1820 1.3500 ;
      RECT 15.5210 0.2565 16.2500 1.1720 ;
      RECT 15.2870 0.4520 15.4850 1.3500 ;
      RECT 14.1080 0.3560 15.2600 1.1720 ;
      RECT 0.1760 0.2565 14.0900 1.3500 ;
      RECT 0.0050 0.2565 0.1580 1.1720 ;
      RECT 15.4670 0.2565 30.3530 1.0760 ;
      RECT 0.0050 0.3560 15.4490 1.0760 ;
      RECT 15.2420 0.2565 30.3530 0.4280 ;
      RECT 0.0050 0.2565 15.2240 1.0760 ;
      RECT 0.0050 0.2565 30.3530 0.3320 ;
      RECT 0.0050 2.3000 30.3530 2.4300 ;
      RECT 30.2360 1.3365 30.3530 2.4300 ;
      RECT 16.2140 2.2040 30.2180 2.4300 ;
      RECT 14.8820 2.2040 16.1960 2.4300 ;
      RECT 14.1620 1.3365 14.7920 2.4300 ;
      RECT 0.1400 2.2040 14.1440 2.4300 ;
      RECT 0.0050 1.3365 0.1220 2.4300 ;
      RECT 30.2000 1.3365 30.3530 2.2520 ;
      RECT 16.2680 1.3365 30.1820 2.4300 ;
      RECT 15.5210 1.3365 16.2500 2.2520 ;
      RECT 15.2870 1.5320 15.4850 2.4300 ;
      RECT 14.1080 1.4360 15.2600 2.2520 ;
      RECT 0.1760 1.3365 14.0900 2.4300 ;
      RECT 0.0050 1.3365 0.1580 2.2520 ;
      RECT 15.4670 1.3365 30.3530 2.1560 ;
      RECT 0.0050 1.4360 15.4490 2.1560 ;
      RECT 15.2420 1.3365 30.3530 1.5080 ;
      RECT 0.0050 1.3365 15.2240 2.1560 ;
      RECT 0.0050 1.3365 30.3530 1.4120 ;
      RECT 0.0050 3.3800 30.3530 3.5100 ;
      RECT 30.2360 2.4165 30.3530 3.5100 ;
      RECT 16.2140 3.2840 30.2180 3.5100 ;
      RECT 14.8820 3.2840 16.1960 3.5100 ;
      RECT 14.1620 2.4165 14.7920 3.5100 ;
      RECT 0.1400 3.2840 14.1440 3.5100 ;
      RECT 0.0050 2.4165 0.1220 3.5100 ;
      RECT 30.2000 2.4165 30.3530 3.3320 ;
      RECT 16.2680 2.4165 30.1820 3.5100 ;
      RECT 15.5210 2.4165 16.2500 3.3320 ;
      RECT 15.2870 2.6120 15.4850 3.5100 ;
      RECT 14.1080 2.5160 15.2600 3.3320 ;
      RECT 0.1760 2.4165 14.0900 3.5100 ;
      RECT 0.0050 2.4165 0.1580 3.3320 ;
      RECT 15.4670 2.4165 30.3530 3.2360 ;
      RECT 0.0050 2.5160 15.4490 3.2360 ;
      RECT 15.2420 2.4165 30.3530 2.5880 ;
      RECT 0.0050 2.4165 15.2240 3.2360 ;
      RECT 0.0050 2.4165 30.3530 2.4920 ;
      RECT 0.0050 4.4600 30.3530 4.5900 ;
      RECT 30.2360 3.4965 30.3530 4.5900 ;
      RECT 16.2140 4.3640 30.2180 4.5900 ;
      RECT 14.8820 4.3640 16.1960 4.5900 ;
      RECT 14.1620 3.4965 14.7920 4.5900 ;
      RECT 0.1400 4.3640 14.1440 4.5900 ;
      RECT 0.0050 3.4965 0.1220 4.5900 ;
      RECT 30.2000 3.4965 30.3530 4.4120 ;
      RECT 16.2680 3.4965 30.1820 4.5900 ;
      RECT 15.5210 3.4965 16.2500 4.4120 ;
      RECT 15.2870 3.6920 15.4850 4.5900 ;
      RECT 14.1080 3.5960 15.2600 4.4120 ;
      RECT 0.1760 3.4965 14.0900 4.5900 ;
      RECT 0.0050 3.4965 0.1580 4.4120 ;
      RECT 15.4670 3.4965 30.3530 4.3160 ;
      RECT 0.0050 3.5960 15.4490 4.3160 ;
      RECT 15.2420 3.4965 30.3530 3.6680 ;
      RECT 0.0050 3.4965 15.2240 4.3160 ;
      RECT 0.0050 3.4965 30.3530 3.5720 ;
      RECT 0.0050 5.5400 30.3530 5.6700 ;
      RECT 30.2360 4.5765 30.3530 5.6700 ;
      RECT 16.2140 5.4440 30.2180 5.6700 ;
      RECT 14.8820 5.4440 16.1960 5.6700 ;
      RECT 14.1620 4.5765 14.7920 5.6700 ;
      RECT 0.1400 5.4440 14.1440 5.6700 ;
      RECT 0.0050 4.5765 0.1220 5.6700 ;
      RECT 30.2000 4.5765 30.3530 5.4920 ;
      RECT 16.2680 4.5765 30.1820 5.6700 ;
      RECT 15.5210 4.5765 16.2500 5.4920 ;
      RECT 15.2870 4.7720 15.4850 5.6700 ;
      RECT 14.1080 4.6760 15.2600 5.4920 ;
      RECT 0.1760 4.5765 14.0900 5.6700 ;
      RECT 0.0050 4.5765 0.1580 5.4920 ;
      RECT 15.4670 4.5765 30.3530 5.3960 ;
      RECT 0.0050 4.6760 15.4490 5.3960 ;
      RECT 15.2420 4.5765 30.3530 4.7480 ;
      RECT 0.0050 4.5765 15.2240 5.3960 ;
      RECT 0.0050 4.5765 30.3530 4.6520 ;
      RECT 0.0050 6.6200 30.3530 6.7500 ;
      RECT 30.2360 5.6565 30.3530 6.7500 ;
      RECT 16.2140 6.5240 30.2180 6.7500 ;
      RECT 14.8820 6.5240 16.1960 6.7500 ;
      RECT 14.1620 5.6565 14.7920 6.7500 ;
      RECT 0.1400 6.5240 14.1440 6.7500 ;
      RECT 0.0050 5.6565 0.1220 6.7500 ;
      RECT 30.2000 5.6565 30.3530 6.5720 ;
      RECT 16.2680 5.6565 30.1820 6.7500 ;
      RECT 15.5210 5.6565 16.2500 6.5720 ;
      RECT 15.2870 5.8520 15.4850 6.7500 ;
      RECT 14.1080 5.7560 15.2600 6.5720 ;
      RECT 0.1760 5.6565 14.0900 6.7500 ;
      RECT 0.0050 5.6565 0.1580 6.5720 ;
      RECT 15.4670 5.6565 30.3530 6.4760 ;
      RECT 0.0050 5.7560 15.4490 6.4760 ;
      RECT 15.2420 5.6565 30.3530 5.8280 ;
      RECT 0.0050 5.6565 15.2240 6.4760 ;
      RECT 0.0050 5.6565 30.3530 5.7320 ;
      RECT 0.0050 7.7000 30.3530 7.8300 ;
      RECT 30.2360 6.7365 30.3530 7.8300 ;
      RECT 16.2140 7.6040 30.2180 7.8300 ;
      RECT 14.8820 7.6040 16.1960 7.8300 ;
      RECT 14.1620 6.7365 14.7920 7.8300 ;
      RECT 0.1400 7.6040 14.1440 7.8300 ;
      RECT 0.0050 6.7365 0.1220 7.8300 ;
      RECT 30.2000 6.7365 30.3530 7.6520 ;
      RECT 16.2680 6.7365 30.1820 7.8300 ;
      RECT 15.5210 6.7365 16.2500 7.6520 ;
      RECT 15.2870 6.9320 15.4850 7.8300 ;
      RECT 14.1080 6.8360 15.2600 7.6520 ;
      RECT 0.1760 6.7365 14.0900 7.8300 ;
      RECT 0.0050 6.7365 0.1580 7.6520 ;
      RECT 15.4670 6.7365 30.3530 7.5560 ;
      RECT 0.0050 6.8360 15.4490 7.5560 ;
      RECT 15.2420 6.7365 30.3530 6.9080 ;
      RECT 0.0050 6.7365 15.2240 7.5560 ;
      RECT 0.0050 6.7365 30.3530 6.8120 ;
      RECT 0.0050 8.7800 30.3530 8.9100 ;
      RECT 30.2360 7.8165 30.3530 8.9100 ;
      RECT 16.2140 8.6840 30.2180 8.9100 ;
      RECT 14.8820 8.6840 16.1960 8.9100 ;
      RECT 14.1620 7.8165 14.7920 8.9100 ;
      RECT 0.1400 8.6840 14.1440 8.9100 ;
      RECT 0.0050 7.8165 0.1220 8.9100 ;
      RECT 30.2000 7.8165 30.3530 8.7320 ;
      RECT 16.2680 7.8165 30.1820 8.9100 ;
      RECT 15.5210 7.8165 16.2500 8.7320 ;
      RECT 15.2870 8.0120 15.4850 8.9100 ;
      RECT 14.1080 7.9160 15.2600 8.7320 ;
      RECT 0.1760 7.8165 14.0900 8.9100 ;
      RECT 0.0050 7.8165 0.1580 8.7320 ;
      RECT 15.4670 7.8165 30.3530 8.6360 ;
      RECT 0.0050 7.9160 15.4490 8.6360 ;
      RECT 15.2420 7.8165 30.3530 7.9880 ;
      RECT 0.0050 7.8165 15.2240 8.6360 ;
      RECT 0.0050 7.8165 30.3530 7.8920 ;
      RECT 0.0050 9.8600 30.3530 9.9900 ;
      RECT 30.2360 8.8965 30.3530 9.9900 ;
      RECT 16.2140 9.7640 30.2180 9.9900 ;
      RECT 14.8820 9.7640 16.1960 9.9900 ;
      RECT 14.1620 8.8965 14.7920 9.9900 ;
      RECT 0.1400 9.7640 14.1440 9.9900 ;
      RECT 0.0050 8.8965 0.1220 9.9900 ;
      RECT 30.2000 8.8965 30.3530 9.8120 ;
      RECT 16.2680 8.8965 30.1820 9.9900 ;
      RECT 15.5210 8.8965 16.2500 9.8120 ;
      RECT 15.2870 9.0920 15.4850 9.9900 ;
      RECT 14.1080 8.9960 15.2600 9.8120 ;
      RECT 0.1760 8.8965 14.0900 9.9900 ;
      RECT 0.0050 8.8965 0.1580 9.8120 ;
      RECT 15.4670 8.8965 30.3530 9.7160 ;
      RECT 0.0050 8.9960 15.4490 9.7160 ;
      RECT 15.2420 8.8965 30.3530 9.0680 ;
      RECT 0.0050 8.8965 15.2240 9.7160 ;
      RECT 0.0050 8.8965 30.3530 8.9720 ;
      RECT 0.0050 10.9400 30.3530 11.0700 ;
      RECT 30.2360 9.9765 30.3530 11.0700 ;
      RECT 16.2140 10.8440 30.2180 11.0700 ;
      RECT 14.8820 10.8440 16.1960 11.0700 ;
      RECT 14.1620 9.9765 14.7920 11.0700 ;
      RECT 0.1400 10.8440 14.1440 11.0700 ;
      RECT 0.0050 9.9765 0.1220 11.0700 ;
      RECT 30.2000 9.9765 30.3530 10.8920 ;
      RECT 16.2680 9.9765 30.1820 11.0700 ;
      RECT 15.5210 9.9765 16.2500 10.8920 ;
      RECT 15.2870 10.1720 15.4850 11.0700 ;
      RECT 14.1080 10.0760 15.2600 10.8920 ;
      RECT 0.1760 9.9765 14.0900 11.0700 ;
      RECT 0.0050 9.9765 0.1580 10.8920 ;
      RECT 15.4670 9.9765 30.3530 10.7960 ;
      RECT 0.0050 10.0760 15.4490 10.7960 ;
      RECT 15.2420 9.9765 30.3530 10.1480 ;
      RECT 0.0050 9.9765 15.2240 10.7960 ;
      RECT 0.0050 9.9765 30.3530 10.0520 ;
      RECT 0.0050 12.0200 30.3530 12.1500 ;
      RECT 30.2360 11.0565 30.3530 12.1500 ;
      RECT 16.2140 11.9240 30.2180 12.1500 ;
      RECT 14.8820 11.9240 16.1960 12.1500 ;
      RECT 14.1620 11.0565 14.7920 12.1500 ;
      RECT 0.1400 11.9240 14.1440 12.1500 ;
      RECT 0.0050 11.0565 0.1220 12.1500 ;
      RECT 30.2000 11.0565 30.3530 11.9720 ;
      RECT 16.2680 11.0565 30.1820 12.1500 ;
      RECT 15.5210 11.0565 16.2500 11.9720 ;
      RECT 15.2870 11.2520 15.4850 12.1500 ;
      RECT 14.1080 11.1560 15.2600 11.9720 ;
      RECT 0.1760 11.0565 14.0900 12.1500 ;
      RECT 0.0050 11.0565 0.1580 11.9720 ;
      RECT 15.4670 11.0565 30.3530 11.8760 ;
      RECT 0.0050 11.1560 15.4490 11.8760 ;
      RECT 15.2420 11.0565 30.3530 11.2280 ;
      RECT 0.0050 11.0565 15.2240 11.8760 ;
      RECT 0.0050 11.0565 30.3530 11.1320 ;
      RECT 0.0050 13.1000 30.3530 13.2300 ;
      RECT 30.2360 12.1365 30.3530 13.2300 ;
      RECT 16.2140 13.0040 30.2180 13.2300 ;
      RECT 14.8820 13.0040 16.1960 13.2300 ;
      RECT 14.1620 12.1365 14.7920 13.2300 ;
      RECT 0.1400 13.0040 14.1440 13.2300 ;
      RECT 0.0050 12.1365 0.1220 13.2300 ;
      RECT 30.2000 12.1365 30.3530 13.0520 ;
      RECT 16.2680 12.1365 30.1820 13.2300 ;
      RECT 15.5210 12.1365 16.2500 13.0520 ;
      RECT 15.2870 12.3320 15.4850 13.2300 ;
      RECT 14.1080 12.2360 15.2600 13.0520 ;
      RECT 0.1760 12.1365 14.0900 13.2300 ;
      RECT 0.0050 12.1365 0.1580 13.0520 ;
      RECT 15.4670 12.1365 30.3530 12.9560 ;
      RECT 0.0050 12.2360 15.4490 12.9560 ;
      RECT 15.2420 12.1365 30.3530 12.3080 ;
      RECT 0.0050 12.1365 15.2240 12.9560 ;
      RECT 0.0050 12.1365 30.3530 12.2120 ;
      RECT 0.0050 14.1800 30.3530 14.3100 ;
      RECT 30.2360 13.2165 30.3530 14.3100 ;
      RECT 16.2140 14.0840 30.2180 14.3100 ;
      RECT 14.8820 14.0840 16.1960 14.3100 ;
      RECT 14.1620 13.2165 14.7920 14.3100 ;
      RECT 0.1400 14.0840 14.1440 14.3100 ;
      RECT 0.0050 13.2165 0.1220 14.3100 ;
      RECT 30.2000 13.2165 30.3530 14.1320 ;
      RECT 16.2680 13.2165 30.1820 14.3100 ;
      RECT 15.5210 13.2165 16.2500 14.1320 ;
      RECT 15.2870 13.4120 15.4850 14.3100 ;
      RECT 14.1080 13.3160 15.2600 14.1320 ;
      RECT 0.1760 13.2165 14.0900 14.3100 ;
      RECT 0.0050 13.2165 0.1580 14.1320 ;
      RECT 15.4670 13.2165 30.3530 14.0360 ;
      RECT 0.0050 13.3160 15.4490 14.0360 ;
      RECT 15.2420 13.2165 30.3530 13.3880 ;
      RECT 0.0050 13.2165 15.2240 14.0360 ;
      RECT 0.0050 13.2165 30.3530 13.2920 ;
      RECT 0.0050 15.2600 30.3530 15.3900 ;
      RECT 30.2360 14.2965 30.3530 15.3900 ;
      RECT 16.2140 15.1640 30.2180 15.3900 ;
      RECT 14.8820 15.1640 16.1960 15.3900 ;
      RECT 14.1620 14.2965 14.7920 15.3900 ;
      RECT 0.1400 15.1640 14.1440 15.3900 ;
      RECT 0.0050 14.2965 0.1220 15.3900 ;
      RECT 30.2000 14.2965 30.3530 15.2120 ;
      RECT 16.2680 14.2965 30.1820 15.3900 ;
      RECT 15.5210 14.2965 16.2500 15.2120 ;
      RECT 15.2870 14.4920 15.4850 15.3900 ;
      RECT 14.1080 14.3960 15.2600 15.2120 ;
      RECT 0.1760 14.2965 14.0900 15.3900 ;
      RECT 0.0050 14.2965 0.1580 15.2120 ;
      RECT 15.4670 14.2965 30.3530 15.1160 ;
      RECT 0.0050 14.3960 15.4490 15.1160 ;
      RECT 15.2420 14.2965 30.3530 14.4680 ;
      RECT 0.0050 14.2965 15.2240 15.1160 ;
      RECT 0.0050 14.2965 30.3530 14.3720 ;
      RECT 0.0050 16.3400 30.3530 16.4700 ;
      RECT 30.2360 15.3765 30.3530 16.4700 ;
      RECT 16.2140 16.2440 30.2180 16.4700 ;
      RECT 14.8820 16.2440 16.1960 16.4700 ;
      RECT 14.1620 15.3765 14.7920 16.4700 ;
      RECT 0.1400 16.2440 14.1440 16.4700 ;
      RECT 0.0050 15.3765 0.1220 16.4700 ;
      RECT 30.2000 15.3765 30.3530 16.2920 ;
      RECT 16.2680 15.3765 30.1820 16.4700 ;
      RECT 15.5210 15.3765 16.2500 16.2920 ;
      RECT 15.2870 15.5720 15.4850 16.4700 ;
      RECT 14.1080 15.4760 15.2600 16.2920 ;
      RECT 0.1760 15.3765 14.0900 16.4700 ;
      RECT 0.0050 15.3765 0.1580 16.2920 ;
      RECT 15.4670 15.3765 30.3530 16.1960 ;
      RECT 0.0050 15.4760 15.4490 16.1960 ;
      RECT 15.2420 15.3765 30.3530 15.5480 ;
      RECT 0.0050 15.3765 15.2240 16.1960 ;
      RECT 0.0050 15.3765 30.3530 15.4520 ;
      RECT 0.0050 17.4200 30.3530 17.5500 ;
      RECT 30.2360 16.4565 30.3530 17.5500 ;
      RECT 16.2140 17.3240 30.2180 17.5500 ;
      RECT 14.8820 17.3240 16.1960 17.5500 ;
      RECT 14.1620 16.4565 14.7920 17.5500 ;
      RECT 0.1400 17.3240 14.1440 17.5500 ;
      RECT 0.0050 16.4565 0.1220 17.5500 ;
      RECT 30.2000 16.4565 30.3530 17.3720 ;
      RECT 16.2680 16.4565 30.1820 17.5500 ;
      RECT 15.5210 16.4565 16.2500 17.3720 ;
      RECT 15.2870 16.6520 15.4850 17.5500 ;
      RECT 14.1080 16.5560 15.2600 17.3720 ;
      RECT 0.1760 16.4565 14.0900 17.5500 ;
      RECT 0.0050 16.4565 0.1580 17.3720 ;
      RECT 15.4670 16.4565 30.3530 17.2760 ;
      RECT 0.0050 16.5560 15.4490 17.2760 ;
      RECT 15.2420 16.4565 30.3530 16.6280 ;
      RECT 0.0050 16.4565 15.2240 17.2760 ;
      RECT 0.0050 16.4565 30.3530 16.5320 ;
      RECT 0.0000 24.8935 30.3480 26.2270 ;
      RECT 17.7210 17.5735 30.3480 26.2270 ;
      RECT 15.5210 19.0375 30.3480 26.2270 ;
      RECT 16.4250 18.8455 30.3480 26.2270 ;
      RECT 15.4690 17.5735 15.5030 26.2270 ;
      RECT 15.4170 17.5735 15.4510 26.2270 ;
      RECT 15.3650 17.5735 15.3990 26.2270 ;
      RECT 15.3130 17.5735 15.3470 26.2270 ;
      RECT 0.0000 19.1335 15.2950 26.2270 ;
      RECT 0.0000 21.7255 30.3480 24.6775 ;
      RECT 14.1570 18.5575 15.8310 21.5095 ;
      RECT 0.0000 18.8455 14.1390 26.2270 ;
      RECT 0.0000 18.9415 16.4070 19.1095 ;
      RECT 16.2090 18.8455 30.3480 19.0135 ;
      RECT 0.0000 18.8455 16.1910 19.1095 ;
      RECT 17.5050 17.5735 17.7030 26.2270 ;
      RECT 13.7250 18.6535 17.4870 18.9175 ;
      RECT 12.8610 18.2695 13.7070 26.2270 ;
      RECT 0.0000 17.5735 12.8430 26.2270 ;
      RECT 17.2890 17.5735 30.3480 18.8215 ;
      RECT 17.0730 18.2695 30.3480 18.8215 ;
      RECT 15.8490 18.5575 17.0550 18.9175 ;
      RECT 0.0000 18.5575 15.8310 18.8215 ;
      RECT 16.8570 17.5735 17.2710 18.6295 ;
      RECT 16.2630 18.2695 30.3480 18.6295 ;
      RECT 15.5210 18.2695 16.2450 18.6295 ;
      RECT 14.1030 18.2695 15.2950 19.1095 ;
      RECT 0.0000 18.2695 14.0850 18.8215 ;
      RECT 15.5610 18.2215 16.8390 18.3415 ;
      RECT 14.3730 18.2215 15.5430 18.3415 ;
      RECT 13.5090 18.2215 14.3550 18.3415 ;
      RECT 13.0770 18.2215 13.4910 26.2270 ;
      RECT 0.0000 17.5735 13.0590 18.8215 ;
      RECT 16.6410 17.5735 30.3480 18.2455 ;
      RECT 15.1650 17.5735 16.6230 18.2455 ;
      RECT 14.1930 17.5735 15.1470 18.2455 ;
      RECT 13.2930 17.5735 14.1750 18.2455 ;
      RECT 0.0000 17.5735 13.2750 18.2455 ;
      RECT 0.0000 17.5735 30.3480 18.1975 ;
        RECT 0.0050 26.6270 30.3530 26.7570 ;
        RECT 30.2360 25.6635 30.3530 26.7570 ;
        RECT 16.2140 26.5310 30.2180 26.7570 ;
        RECT 14.8820 26.5310 16.1960 26.7570 ;
        RECT 14.1620 25.6635 14.7920 26.7570 ;
        RECT 0.1400 26.5310 14.1440 26.7570 ;
        RECT 0.0050 25.6635 0.1220 26.7570 ;
        RECT 30.2000 25.6635 30.3530 26.5790 ;
        RECT 16.2680 25.6635 30.1820 26.7570 ;
        RECT 15.5210 25.6635 16.2500 26.5790 ;
        RECT 15.2870 25.8590 15.4850 26.7570 ;
        RECT 14.1080 25.7630 15.2600 26.5790 ;
        RECT 0.1760 25.6635 14.0900 26.7570 ;
        RECT 0.0050 25.6635 0.1580 26.5790 ;
        RECT 15.4670 25.6635 30.3530 26.4830 ;
        RECT 0.0050 25.7630 15.4490 26.4830 ;
        RECT 15.2420 25.6635 30.3530 25.8350 ;
        RECT 0.0050 25.6635 15.2240 26.4830 ;
        RECT 0.0050 25.6635 30.3530 25.7390 ;
        RECT 0.0050 27.7070 30.3530 27.8370 ;
        RECT 30.2360 26.7435 30.3530 27.8370 ;
        RECT 16.2140 27.6110 30.2180 27.8370 ;
        RECT 14.8820 27.6110 16.1960 27.8370 ;
        RECT 14.1620 26.7435 14.7920 27.8370 ;
        RECT 0.1400 27.6110 14.1440 27.8370 ;
        RECT 0.0050 26.7435 0.1220 27.8370 ;
        RECT 30.2000 26.7435 30.3530 27.6590 ;
        RECT 16.2680 26.7435 30.1820 27.8370 ;
        RECT 15.5210 26.7435 16.2500 27.6590 ;
        RECT 15.2870 26.9390 15.4850 27.8370 ;
        RECT 14.1080 26.8430 15.2600 27.6590 ;
        RECT 0.1760 26.7435 14.0900 27.8370 ;
        RECT 0.0050 26.7435 0.1580 27.6590 ;
        RECT 15.4670 26.7435 30.3530 27.5630 ;
        RECT 0.0050 26.8430 15.4490 27.5630 ;
        RECT 15.2420 26.7435 30.3530 26.9150 ;
        RECT 0.0050 26.7435 15.2240 27.5630 ;
        RECT 0.0050 26.7435 30.3530 26.8190 ;
        RECT 0.0050 28.7870 30.3530 28.9170 ;
        RECT 30.2360 27.8235 30.3530 28.9170 ;
        RECT 16.2140 28.6910 30.2180 28.9170 ;
        RECT 14.8820 28.6910 16.1960 28.9170 ;
        RECT 14.1620 27.8235 14.7920 28.9170 ;
        RECT 0.1400 28.6910 14.1440 28.9170 ;
        RECT 0.0050 27.8235 0.1220 28.9170 ;
        RECT 30.2000 27.8235 30.3530 28.7390 ;
        RECT 16.2680 27.8235 30.1820 28.9170 ;
        RECT 15.5210 27.8235 16.2500 28.7390 ;
        RECT 15.2870 28.0190 15.4850 28.9170 ;
        RECT 14.1080 27.9230 15.2600 28.7390 ;
        RECT 0.1760 27.8235 14.0900 28.9170 ;
        RECT 0.0050 27.8235 0.1580 28.7390 ;
        RECT 15.4670 27.8235 30.3530 28.6430 ;
        RECT 0.0050 27.9230 15.4490 28.6430 ;
        RECT 15.2420 27.8235 30.3530 27.9950 ;
        RECT 0.0050 27.8235 15.2240 28.6430 ;
        RECT 0.0050 27.8235 30.3530 27.8990 ;
        RECT 0.0050 29.8670 30.3530 29.9970 ;
        RECT 30.2360 28.9035 30.3530 29.9970 ;
        RECT 16.2140 29.7710 30.2180 29.9970 ;
        RECT 14.8820 29.7710 16.1960 29.9970 ;
        RECT 14.1620 28.9035 14.7920 29.9970 ;
        RECT 0.1400 29.7710 14.1440 29.9970 ;
        RECT 0.0050 28.9035 0.1220 29.9970 ;
        RECT 30.2000 28.9035 30.3530 29.8190 ;
        RECT 16.2680 28.9035 30.1820 29.9970 ;
        RECT 15.5210 28.9035 16.2500 29.8190 ;
        RECT 15.2870 29.0990 15.4850 29.9970 ;
        RECT 14.1080 29.0030 15.2600 29.8190 ;
        RECT 0.1760 28.9035 14.0900 29.9970 ;
        RECT 0.0050 28.9035 0.1580 29.8190 ;
        RECT 15.4670 28.9035 30.3530 29.7230 ;
        RECT 0.0050 29.0030 15.4490 29.7230 ;
        RECT 15.2420 28.9035 30.3530 29.0750 ;
        RECT 0.0050 28.9035 15.2240 29.7230 ;
        RECT 0.0050 28.9035 30.3530 28.9790 ;
        RECT 0.0050 30.9470 30.3530 31.0770 ;
        RECT 30.2360 29.9835 30.3530 31.0770 ;
        RECT 16.2140 30.8510 30.2180 31.0770 ;
        RECT 14.8820 30.8510 16.1960 31.0770 ;
        RECT 14.1620 29.9835 14.7920 31.0770 ;
        RECT 0.1400 30.8510 14.1440 31.0770 ;
        RECT 0.0050 29.9835 0.1220 31.0770 ;
        RECT 30.2000 29.9835 30.3530 30.8990 ;
        RECT 16.2680 29.9835 30.1820 31.0770 ;
        RECT 15.5210 29.9835 16.2500 30.8990 ;
        RECT 15.2870 30.1790 15.4850 31.0770 ;
        RECT 14.1080 30.0830 15.2600 30.8990 ;
        RECT 0.1760 29.9835 14.0900 31.0770 ;
        RECT 0.0050 29.9835 0.1580 30.8990 ;
        RECT 15.4670 29.9835 30.3530 30.8030 ;
        RECT 0.0050 30.0830 15.4490 30.8030 ;
        RECT 15.2420 29.9835 30.3530 30.1550 ;
        RECT 0.0050 29.9835 15.2240 30.8030 ;
        RECT 0.0050 29.9835 30.3530 30.0590 ;
        RECT 0.0050 32.0270 30.3530 32.1570 ;
        RECT 30.2360 31.0635 30.3530 32.1570 ;
        RECT 16.2140 31.9310 30.2180 32.1570 ;
        RECT 14.8820 31.9310 16.1960 32.1570 ;
        RECT 14.1620 31.0635 14.7920 32.1570 ;
        RECT 0.1400 31.9310 14.1440 32.1570 ;
        RECT 0.0050 31.0635 0.1220 32.1570 ;
        RECT 30.2000 31.0635 30.3530 31.9790 ;
        RECT 16.2680 31.0635 30.1820 32.1570 ;
        RECT 15.5210 31.0635 16.2500 31.9790 ;
        RECT 15.2870 31.2590 15.4850 32.1570 ;
        RECT 14.1080 31.1630 15.2600 31.9790 ;
        RECT 0.1760 31.0635 14.0900 32.1570 ;
        RECT 0.0050 31.0635 0.1580 31.9790 ;
        RECT 15.4670 31.0635 30.3530 31.8830 ;
        RECT 0.0050 31.1630 15.4490 31.8830 ;
        RECT 15.2420 31.0635 30.3530 31.2350 ;
        RECT 0.0050 31.0635 15.2240 31.8830 ;
        RECT 0.0050 31.0635 30.3530 31.1390 ;
        RECT 0.0050 33.1070 30.3530 33.2370 ;
        RECT 30.2360 32.1435 30.3530 33.2370 ;
        RECT 16.2140 33.0110 30.2180 33.2370 ;
        RECT 14.8820 33.0110 16.1960 33.2370 ;
        RECT 14.1620 32.1435 14.7920 33.2370 ;
        RECT 0.1400 33.0110 14.1440 33.2370 ;
        RECT 0.0050 32.1435 0.1220 33.2370 ;
        RECT 30.2000 32.1435 30.3530 33.0590 ;
        RECT 16.2680 32.1435 30.1820 33.2370 ;
        RECT 15.5210 32.1435 16.2500 33.0590 ;
        RECT 15.2870 32.3390 15.4850 33.2370 ;
        RECT 14.1080 32.2430 15.2600 33.0590 ;
        RECT 0.1760 32.1435 14.0900 33.2370 ;
        RECT 0.0050 32.1435 0.1580 33.0590 ;
        RECT 15.4670 32.1435 30.3530 32.9630 ;
        RECT 0.0050 32.2430 15.4490 32.9630 ;
        RECT 15.2420 32.1435 30.3530 32.3150 ;
        RECT 0.0050 32.1435 15.2240 32.9630 ;
        RECT 0.0050 32.1435 30.3530 32.2190 ;
        RECT 0.0050 34.1870 30.3530 34.3170 ;
        RECT 30.2360 33.2235 30.3530 34.3170 ;
        RECT 16.2140 34.0910 30.2180 34.3170 ;
        RECT 14.8820 34.0910 16.1960 34.3170 ;
        RECT 14.1620 33.2235 14.7920 34.3170 ;
        RECT 0.1400 34.0910 14.1440 34.3170 ;
        RECT 0.0050 33.2235 0.1220 34.3170 ;
        RECT 30.2000 33.2235 30.3530 34.1390 ;
        RECT 16.2680 33.2235 30.1820 34.3170 ;
        RECT 15.5210 33.2235 16.2500 34.1390 ;
        RECT 15.2870 33.4190 15.4850 34.3170 ;
        RECT 14.1080 33.3230 15.2600 34.1390 ;
        RECT 0.1760 33.2235 14.0900 34.3170 ;
        RECT 0.0050 33.2235 0.1580 34.1390 ;
        RECT 15.4670 33.2235 30.3530 34.0430 ;
        RECT 0.0050 33.3230 15.4490 34.0430 ;
        RECT 15.2420 33.2235 30.3530 33.3950 ;
        RECT 0.0050 33.2235 15.2240 34.0430 ;
        RECT 0.0050 33.2235 30.3530 33.2990 ;
        RECT 0.0050 35.2670 30.3530 35.3970 ;
        RECT 30.2360 34.3035 30.3530 35.3970 ;
        RECT 16.2140 35.1710 30.2180 35.3970 ;
        RECT 14.8820 35.1710 16.1960 35.3970 ;
        RECT 14.1620 34.3035 14.7920 35.3970 ;
        RECT 0.1400 35.1710 14.1440 35.3970 ;
        RECT 0.0050 34.3035 0.1220 35.3970 ;
        RECT 30.2000 34.3035 30.3530 35.2190 ;
        RECT 16.2680 34.3035 30.1820 35.3970 ;
        RECT 15.5210 34.3035 16.2500 35.2190 ;
        RECT 15.2870 34.4990 15.4850 35.3970 ;
        RECT 14.1080 34.4030 15.2600 35.2190 ;
        RECT 0.1760 34.3035 14.0900 35.3970 ;
        RECT 0.0050 34.3035 0.1580 35.2190 ;
        RECT 15.4670 34.3035 30.3530 35.1230 ;
        RECT 0.0050 34.4030 15.4490 35.1230 ;
        RECT 15.2420 34.3035 30.3530 34.4750 ;
        RECT 0.0050 34.3035 15.2240 35.1230 ;
        RECT 0.0050 34.3035 30.3530 34.3790 ;
        RECT 0.0050 36.3470 30.3530 36.4770 ;
        RECT 30.2360 35.3835 30.3530 36.4770 ;
        RECT 16.2140 36.2510 30.2180 36.4770 ;
        RECT 14.8820 36.2510 16.1960 36.4770 ;
        RECT 14.1620 35.3835 14.7920 36.4770 ;
        RECT 0.1400 36.2510 14.1440 36.4770 ;
        RECT 0.0050 35.3835 0.1220 36.4770 ;
        RECT 30.2000 35.3835 30.3530 36.2990 ;
        RECT 16.2680 35.3835 30.1820 36.4770 ;
        RECT 15.5210 35.3835 16.2500 36.2990 ;
        RECT 15.2870 35.5790 15.4850 36.4770 ;
        RECT 14.1080 35.4830 15.2600 36.2990 ;
        RECT 0.1760 35.3835 14.0900 36.4770 ;
        RECT 0.0050 35.3835 0.1580 36.2990 ;
        RECT 15.4670 35.3835 30.3530 36.2030 ;
        RECT 0.0050 35.4830 15.4490 36.2030 ;
        RECT 15.2420 35.3835 30.3530 35.5550 ;
        RECT 0.0050 35.3835 15.2240 36.2030 ;
        RECT 0.0050 35.3835 30.3530 35.4590 ;
        RECT 0.0050 37.4270 30.3530 37.5570 ;
        RECT 30.2360 36.4635 30.3530 37.5570 ;
        RECT 16.2140 37.3310 30.2180 37.5570 ;
        RECT 14.8820 37.3310 16.1960 37.5570 ;
        RECT 14.1620 36.4635 14.7920 37.5570 ;
        RECT 0.1400 37.3310 14.1440 37.5570 ;
        RECT 0.0050 36.4635 0.1220 37.5570 ;
        RECT 30.2000 36.4635 30.3530 37.3790 ;
        RECT 16.2680 36.4635 30.1820 37.5570 ;
        RECT 15.5210 36.4635 16.2500 37.3790 ;
        RECT 15.2870 36.6590 15.4850 37.5570 ;
        RECT 14.1080 36.5630 15.2600 37.3790 ;
        RECT 0.1760 36.4635 14.0900 37.5570 ;
        RECT 0.0050 36.4635 0.1580 37.3790 ;
        RECT 15.4670 36.4635 30.3530 37.2830 ;
        RECT 0.0050 36.5630 15.4490 37.2830 ;
        RECT 15.2420 36.4635 30.3530 36.6350 ;
        RECT 0.0050 36.4635 15.2240 37.2830 ;
        RECT 0.0050 36.4635 30.3530 36.5390 ;
        RECT 0.0050 38.5070 30.3530 38.6370 ;
        RECT 30.2360 37.5435 30.3530 38.6370 ;
        RECT 16.2140 38.4110 30.2180 38.6370 ;
        RECT 14.8820 38.4110 16.1960 38.6370 ;
        RECT 14.1620 37.5435 14.7920 38.6370 ;
        RECT 0.1400 38.4110 14.1440 38.6370 ;
        RECT 0.0050 37.5435 0.1220 38.6370 ;
        RECT 30.2000 37.5435 30.3530 38.4590 ;
        RECT 16.2680 37.5435 30.1820 38.6370 ;
        RECT 15.5210 37.5435 16.2500 38.4590 ;
        RECT 15.2870 37.7390 15.4850 38.6370 ;
        RECT 14.1080 37.6430 15.2600 38.4590 ;
        RECT 0.1760 37.5435 14.0900 38.6370 ;
        RECT 0.0050 37.5435 0.1580 38.4590 ;
        RECT 15.4670 37.5435 30.3530 38.3630 ;
        RECT 0.0050 37.6430 15.4490 38.3630 ;
        RECT 15.2420 37.5435 30.3530 37.7150 ;
        RECT 0.0050 37.5435 15.2240 38.3630 ;
        RECT 0.0050 37.5435 30.3530 37.6190 ;
        RECT 0.0050 39.5870 30.3530 39.7170 ;
        RECT 30.2360 38.6235 30.3530 39.7170 ;
        RECT 16.2140 39.4910 30.2180 39.7170 ;
        RECT 14.8820 39.4910 16.1960 39.7170 ;
        RECT 14.1620 38.6235 14.7920 39.7170 ;
        RECT 0.1400 39.4910 14.1440 39.7170 ;
        RECT 0.0050 38.6235 0.1220 39.7170 ;
        RECT 30.2000 38.6235 30.3530 39.5390 ;
        RECT 16.2680 38.6235 30.1820 39.7170 ;
        RECT 15.5210 38.6235 16.2500 39.5390 ;
        RECT 15.2870 38.8190 15.4850 39.7170 ;
        RECT 14.1080 38.7230 15.2600 39.5390 ;
        RECT 0.1760 38.6235 14.0900 39.7170 ;
        RECT 0.0050 38.6235 0.1580 39.5390 ;
        RECT 15.4670 38.6235 30.3530 39.4430 ;
        RECT 0.0050 38.7230 15.4490 39.4430 ;
        RECT 15.2420 38.6235 30.3530 38.7950 ;
        RECT 0.0050 38.6235 15.2240 39.4430 ;
        RECT 0.0050 38.6235 30.3530 38.6990 ;
        RECT 0.0050 40.6670 30.3530 40.7970 ;
        RECT 30.2360 39.7035 30.3530 40.7970 ;
        RECT 16.2140 40.5710 30.2180 40.7970 ;
        RECT 14.8820 40.5710 16.1960 40.7970 ;
        RECT 14.1620 39.7035 14.7920 40.7970 ;
        RECT 0.1400 40.5710 14.1440 40.7970 ;
        RECT 0.0050 39.7035 0.1220 40.7970 ;
        RECT 30.2000 39.7035 30.3530 40.6190 ;
        RECT 16.2680 39.7035 30.1820 40.7970 ;
        RECT 15.5210 39.7035 16.2500 40.6190 ;
        RECT 15.2870 39.8990 15.4850 40.7970 ;
        RECT 14.1080 39.8030 15.2600 40.6190 ;
        RECT 0.1760 39.7035 14.0900 40.7970 ;
        RECT 0.0050 39.7035 0.1580 40.6190 ;
        RECT 15.4670 39.7035 30.3530 40.5230 ;
        RECT 0.0050 39.8030 15.4490 40.5230 ;
        RECT 15.2420 39.7035 30.3530 39.8750 ;
        RECT 0.0050 39.7035 15.2240 40.5230 ;
        RECT 0.0050 39.7035 30.3530 39.7790 ;
        RECT 0.0050 41.7470 30.3530 41.8770 ;
        RECT 30.2360 40.7835 30.3530 41.8770 ;
        RECT 16.2140 41.6510 30.2180 41.8770 ;
        RECT 14.8820 41.6510 16.1960 41.8770 ;
        RECT 14.1620 40.7835 14.7920 41.8770 ;
        RECT 0.1400 41.6510 14.1440 41.8770 ;
        RECT 0.0050 40.7835 0.1220 41.8770 ;
        RECT 30.2000 40.7835 30.3530 41.6990 ;
        RECT 16.2680 40.7835 30.1820 41.8770 ;
        RECT 15.5210 40.7835 16.2500 41.6990 ;
        RECT 15.2870 40.9790 15.4850 41.8770 ;
        RECT 14.1080 40.8830 15.2600 41.6990 ;
        RECT 0.1760 40.7835 14.0900 41.8770 ;
        RECT 0.0050 40.7835 0.1580 41.6990 ;
        RECT 15.4670 40.7835 30.3530 41.6030 ;
        RECT 0.0050 40.8830 15.4490 41.6030 ;
        RECT 15.2420 40.7835 30.3530 40.9550 ;
        RECT 0.0050 40.7835 15.2240 41.6030 ;
        RECT 0.0050 40.7835 30.3530 40.8590 ;
        RECT 0.0050 42.8270 30.3530 42.9570 ;
        RECT 30.2360 41.8635 30.3530 42.9570 ;
        RECT 16.2140 42.7310 30.2180 42.9570 ;
        RECT 14.8820 42.7310 16.1960 42.9570 ;
        RECT 14.1620 41.8635 14.7920 42.9570 ;
        RECT 0.1400 42.7310 14.1440 42.9570 ;
        RECT 0.0050 41.8635 0.1220 42.9570 ;
        RECT 30.2000 41.8635 30.3530 42.7790 ;
        RECT 16.2680 41.8635 30.1820 42.9570 ;
        RECT 15.5210 41.8635 16.2500 42.7790 ;
        RECT 15.2870 42.0590 15.4850 42.9570 ;
        RECT 14.1080 41.9630 15.2600 42.7790 ;
        RECT 0.1760 41.8635 14.0900 42.9570 ;
        RECT 0.0050 41.8635 0.1580 42.7790 ;
        RECT 15.4670 41.8635 30.3530 42.6830 ;
        RECT 0.0050 41.9630 15.4490 42.6830 ;
        RECT 15.2420 41.8635 30.3530 42.0350 ;
        RECT 0.0050 41.8635 15.2240 42.6830 ;
        RECT 0.0050 41.8635 30.3530 41.9390 ;
  LAYER M4  ;
      RECT 1.6000 19.2865 28.8355 19.3105 ;
      RECT 1.6000 19.5745 28.8355 19.5985 ;
      RECT 1.6000 19.9585 28.8355 19.9825 ;
      RECT 1.6000 20.0545 28.8355 20.0785 ;
      RECT 1.6000 20.3905 28.8355 20.4145 ;
      RECT 1.6000 20.7745 28.8355 20.7985 ;
      RECT 1.6000 20.8705 28.8355 20.8945 ;
      RECT 10.4760 17.9095 19.8720 18.1255 ;
      RECT 17.8670 18.2455 17.9510 18.2695 ;
      RECT 17.6785 18.6775 17.8085 18.7015 ;
      RECT 17.6870 19.6225 17.8040 19.6465 ;
      RECT 17.6865 19.3350 17.8035 19.3590 ;
      RECT 17.0375 18.6775 17.6085 18.7015 ;
      RECT 17.0975 19.4425 17.2055 19.4665 ;
      RECT 15.7750 19.8295 16.8680 19.8535 ;
      RECT 16.4630 19.3975 16.5470 19.4215 ;
      RECT 15.6790 20.5975 16.5470 20.6215 ;
      RECT 16.4630 20.6935 16.5470 20.7175 ;
      RECT 16.2850 18.9175 16.3690 18.9415 ;
      RECT 16.2470 20.2615 16.3310 20.2855 ;
      RECT 16.2470 20.9815 16.3310 21.0055 ;
      RECT 15.9780 17.6295 16.2410 17.6535 ;
      RECT 16.1090 21.4135 16.2210 21.4375 ;
      RECT 16.0690 18.8215 16.1530 18.8455 ;
      RECT 15.8550 17.5335 16.1180 17.5575 ;
      RECT 15.8550 26.1385 16.1180 26.1625 ;
      RECT 15.8710 20.3095 16.1150 20.3335 ;
      RECT 16.0310 20.4535 16.1150 20.4775 ;
      RECT 14.5750 20.6935 16.1150 20.7175 ;
      RECT 16.0310 20.9815 16.1150 21.0055 ;
      RECT 15.7970 26.0425 16.0600 26.0665 ;
      RECT 15.7960 17.4375 16.0590 17.4615 ;
      RECT 14.3100 21.0775 16.0380 21.2935 ;
      RECT 14.3100 24.2455 16.0380 24.4615 ;
      RECT 15.7580 17.3415 16.0210 17.3655 ;
      RECT 15.7580 25.8505 16.0210 25.8745 ;
      RECT 15.9230 21.4135 16.0070 21.4375 ;
      RECT 15.1510 21.7975 16.0070 21.8215 ;
      RECT 15.5350 24.0535 16.0070 24.0775 ;
      RECT 15.9230 24.1495 16.0070 24.1735 ;
      RECT 15.7100 17.2455 15.9730 17.2695 ;
      RECT 15.7100 25.7545 15.9730 25.7785 ;
      RECT 15.4870 23.1415 15.9320 23.1655 ;
      RECT 15.6660 17.1495 15.9290 17.1735 ;
      RECT 15.6660 26.0905 15.9290 26.1145 ;
      RECT 15.6170 17.4855 15.8800 17.5095 ;
      RECT 15.6170 25.9945 15.8800 26.0185 ;
      RECT 15.7480 20.4535 15.8690 20.4775 ;
      RECT 15.7270 22.5655 15.8600 22.5895 ;
      RECT 15.5700 17.3895 15.8330 17.4135 ;
      RECT 15.5700 25.8985 15.8330 25.9225 ;
      RECT 15.5350 17.1015 15.7980 17.1255 ;
      RECT 15.5350 25.8025 15.7980 25.8265 ;
      RECT 14.7190 24.1495 15.7880 24.1735 ;
      RECT 15.7040 25.3015 15.7880 25.3255 ;
      RECT 15.4790 16.9575 15.7420 16.9815 ;
      RECT 15.4790 25.7065 15.7420 25.7305 ;
      RECT 15.6310 21.4135 15.7160 21.4375 ;
      RECT 14.5270 21.9895 15.6440 22.0135 ;
      RECT 15.1720 19.8295 15.6290 19.8535 ;
      RECT 14.9990 17.6775 15.2660 17.7015 ;
      RECT 14.9990 25.5625 15.2660 25.5865 ;
      RECT 15.1360 21.3655 15.2450 21.3895 ;
      RECT 14.9760 17.5815 15.2180 17.6055 ;
      RECT 14.9760 26.1865 15.2180 26.2105 ;
      RECT 14.9200 17.1015 15.1620 17.1255 ;
      RECT 14.9490 26.2825 15.1620 26.3065 ;
      RECT 15.0650 20.9815 15.1490 21.0055 ;
      RECT 14.8660 17.1975 15.1140 17.2215 ;
      RECT 14.8660 26.1385 15.1140 26.1625 ;
      RECT 14.6320 23.5735 15.0530 23.5975 ;
      RECT 14.6000 17.5335 14.8670 17.5575 ;
      RECT 14.6000 26.2825 14.8670 26.3065 ;
      RECT 14.7400 22.1335 14.8610 22.1575 ;
      RECT 14.7320 25.3015 14.8160 25.3255 ;
      RECT 14.5660 17.4375 14.8130 17.4615 ;
      RECT 14.4990 25.8505 14.8130 25.8745 ;
      RECT 14.5400 17.3415 14.7700 17.3655 ;
      RECT 14.5280 26.1865 14.7700 26.2105 ;
      RECT 14.4870 17.2455 14.7170 17.2695 ;
      RECT 14.6330 23.7175 14.7170 23.7415 ;
      RECT 14.4370 25.7545 14.7170 25.7785 ;
      RECT 14.4420 17.1495 14.6720 17.1735 ;
      RECT 14.4420 26.0905 14.6720 26.1145 ;
      RECT 13.4800 20.9815 14.6690 21.0055 ;
      RECT 14.4040 17.3895 14.6340 17.4135 ;
      RECT 14.4040 25.9945 14.6340 26.0185 ;
      RECT 14.3860 17.2935 14.5790 17.3175 ;
      RECT 14.3860 25.8985 14.5790 25.9225 ;
      RECT 14.3370 17.1975 14.5300 17.2215 ;
      RECT 14.3370 25.8025 14.5300 25.8265 ;
      RECT 14.3410 21.8935 14.5250 21.9175 ;
      RECT 14.2850 17.1015 14.4780 17.1255 ;
      RECT 14.2850 25.7065 14.4780 25.7305 ;
      RECT 13.8010 19.2055 14.4770 19.2295 ;
      RECT 14.3410 21.9895 14.4250 22.0135 ;
      RECT 14.0720 17.6295 14.3350 17.6535 ;
      RECT 14.1950 19.8295 14.2790 19.8535 ;
      RECT 14.1260 21.4135 14.2380 21.4375 ;
      RECT 13.7630 19.3975 13.8470 19.4215 ;
  LAYER V4  ;
      RECT 17.9160 18.2455 17.9400 18.2695 ;
      RECT 17.9160 19.2865 17.9400 19.3105 ;
      RECT 17.7480 19.3350 17.7720 19.3590 ;
      RECT 17.7480 19.6225 17.7720 19.6465 ;
      RECT 17.7475 18.6775 17.7715 18.7015 ;
      RECT 17.1135 18.6775 17.1375 18.7015 ;
      RECT 17.1135 19.4425 17.1375 19.4665 ;
      RECT 16.5120 19.3975 16.5360 19.4215 ;
      RECT 16.5120 19.5745 16.5360 19.5985 ;
      RECT 16.5120 20.5975 16.5360 20.6215 ;
      RECT 16.5120 20.6935 16.5360 20.7175 ;
      RECT 16.2960 18.9175 16.3200 18.9415 ;
      RECT 16.2960 19.9585 16.3200 19.9825 ;
      RECT 16.2960 20.2615 16.3200 20.2855 ;
      RECT 16.2960 20.3905 16.3200 20.4145 ;
      RECT 16.2960 20.7745 16.3200 20.7985 ;
      RECT 16.2960 20.9815 16.3200 21.0055 ;
      RECT 16.1270 17.6295 16.1510 17.6535 ;
      RECT 16.1280 17.9095 16.1510 18.1255 ;
      RECT 16.1270 21.4135 16.1510 21.4375 ;
      RECT 16.0800 18.8215 16.1040 18.8455 ;
      RECT 16.0800 20.0545 16.1040 20.0785 ;
      RECT 16.0800 20.3095 16.1040 20.3335 ;
      RECT 16.0800 20.4535 16.1040 20.4775 ;
      RECT 16.0800 20.6935 16.1040 20.7175 ;
      RECT 16.0800 20.9815 16.1040 21.0055 ;
      RECT 15.9720 21.4135 15.9960 21.4375 ;
      RECT 15.9720 21.7975 15.9960 21.8215 ;
      RECT 15.9720 24.0535 15.9960 24.0775 ;
      RECT 15.9720 24.1495 15.9960 24.1735 ;
      RECT 15.8820 17.5335 15.9060 17.5575 ;
      RECT 15.8820 20.3095 15.9060 20.3335 ;
      RECT 15.8820 26.1385 15.9060 26.1625 ;
      RECT 15.8340 17.4375 15.8580 17.4615 ;
      RECT 15.8340 20.4535 15.8580 20.4775 ;
      RECT 15.8340 26.0425 15.8580 26.0665 ;
      RECT 15.7860 17.3415 15.8100 17.3655 ;
      RECT 15.7860 19.8295 15.8100 19.8535 ;
      RECT 15.7860 25.8505 15.8100 25.8745 ;
      RECT 15.7380 17.2455 15.7620 17.2695 ;
      RECT 15.7380 22.5655 15.7620 22.5895 ;
      RECT 15.7380 25.3015 15.7620 25.3255 ;
      RECT 15.7380 25.7545 15.7620 25.7785 ;
      RECT 15.6900 17.1495 15.7140 17.1735 ;
      RECT 15.6900 20.5975 15.7140 20.6215 ;
      RECT 15.6900 26.0905 15.7140 26.1145 ;
      RECT 15.6420 17.4855 15.6660 17.5095 ;
      RECT 15.6420 21.4135 15.6660 21.4375 ;
      RECT 15.6420 25.9945 15.6660 26.0185 ;
      RECT 15.5940 17.3895 15.6180 17.4135 ;
      RECT 15.5940 19.8295 15.6180 19.8535 ;
      RECT 15.5940 25.8985 15.6180 25.9225 ;
      RECT 15.5460 17.1015 15.5700 17.1255 ;
      RECT 15.5460 24.0535 15.5700 24.0775 ;
      RECT 15.5460 25.8025 15.5700 25.8265 ;
      RECT 15.4980 16.9575 15.5220 16.9815 ;
      RECT 15.4980 23.1415 15.5220 23.1655 ;
      RECT 15.4980 25.7065 15.5220 25.7305 ;
      RECT 15.2100 17.6775 15.2340 17.7015 ;
      RECT 15.2100 21.3655 15.2340 21.3895 ;
      RECT 15.2100 25.5625 15.2340 25.5865 ;
      RECT 15.1620 17.5815 15.1860 17.6055 ;
      RECT 15.1620 21.7975 15.1860 21.8215 ;
      RECT 15.1620 26.1865 15.1860 26.2105 ;
      RECT 15.1140 17.1015 15.1380 17.1255 ;
      RECT 15.1140 20.9815 15.1380 21.0055 ;
      RECT 15.1140 26.2825 15.1380 26.3065 ;
      RECT 15.0180 17.1975 15.0420 17.2215 ;
      RECT 15.0180 23.5735 15.0420 23.5975 ;
      RECT 15.0180 26.1385 15.0420 26.1625 ;
      RECT 14.8260 17.5335 14.8500 17.5575 ;
      RECT 14.8260 22.1335 14.8500 22.1575 ;
      RECT 14.8260 26.2825 14.8500 26.3065 ;
      RECT 14.7780 17.4375 14.8020 17.4615 ;
      RECT 14.7780 25.3015 14.8020 25.3255 ;
      RECT 14.7780 25.8505 14.8020 25.8745 ;
      RECT 14.7300 17.3415 14.7540 17.3655 ;
      RECT 14.7300 24.1495 14.7540 24.1735 ;
      RECT 14.7300 26.1865 14.7540 26.2105 ;
      RECT 14.6820 17.2455 14.7060 17.2695 ;
      RECT 14.6820 23.7175 14.7060 23.7415 ;
      RECT 14.6820 25.7545 14.7060 25.7785 ;
      RECT 14.6340 17.1495 14.6580 17.1735 ;
      RECT 14.6340 20.9815 14.6580 21.0055 ;
      RECT 14.6340 26.0905 14.6580 26.1145 ;
      RECT 14.5860 17.3895 14.6100 17.4135 ;
      RECT 14.5860 20.6935 14.6100 20.7175 ;
      RECT 14.5860 25.9945 14.6100 26.0185 ;
      RECT 14.5380 17.2935 14.5620 17.3175 ;
      RECT 14.5380 21.9895 14.5620 22.0135 ;
      RECT 14.5380 25.8985 14.5620 25.9225 ;
      RECT 14.4900 17.1975 14.5140 17.2215 ;
      RECT 14.4900 21.8935 14.5140 21.9175 ;
      RECT 14.4900 25.8025 14.5140 25.8265 ;
      RECT 14.4420 17.1015 14.4660 17.1255 ;
      RECT 14.4420 19.2055 14.4660 19.2295 ;
      RECT 14.4420 25.7065 14.4660 25.7305 ;
      RECT 14.3520 21.8935 14.3760 21.9175 ;
      RECT 14.3520 21.9895 14.3760 22.0135 ;
      RECT 14.2440 19.8295 14.2680 19.8535 ;
      RECT 14.2440 20.8705 14.2680 20.8945 ;
      RECT 14.1840 17.6295 14.2080 17.6535 ;
      RECT 14.1850 17.9095 14.2080 18.1255 ;
      RECT 14.1840 21.4135 14.2080 21.4375 ;
      RECT 13.8120 19.2055 13.8360 19.2295 ;
      RECT 13.8120 19.3975 13.8360 19.4215 ;
  LAYER M5  ;
      RECT 17.9160 18.2345 17.9400 19.3215 ;
      RECT 17.7475 18.6320 17.7715 19.6925 ;
      RECT 17.1135 18.6360 17.1375 19.5070 ;
      RECT 16.5120 19.3865 16.5360 19.6095 ;
      RECT 16.5120 20.5865 16.5360 20.7285 ;
      RECT 16.2960 18.9065 16.3200 19.9935 ;
      RECT 16.2960 20.2505 16.3200 20.4255 ;
      RECT 16.2960 20.7635 16.3200 21.0165 ;
      RECT 16.1270 17.6115 16.1510 21.4555 ;
      RECT 16.0800 18.8105 16.1040 20.0895 ;
      RECT 16.0800 20.2985 16.1040 20.4885 ;
      RECT 16.0800 20.6825 16.1040 21.0165 ;
      RECT 15.9720 21.4025 15.9960 21.8325 ;
      RECT 15.9720 24.0425 15.9960 24.1845 ;
      RECT 15.8820 16.8810 15.9060 26.3825 ;
      RECT 15.8340 16.8810 15.8580 26.3815 ;
      RECT 15.7860 16.8810 15.8100 26.3815 ;
      RECT 15.7380 16.8810 15.7620 26.3525 ;
      RECT 15.6900 16.8810 15.7140 26.3495 ;
      RECT 15.6420 16.8810 15.6660 26.3515 ;
      RECT 15.5940 16.8810 15.6180 26.3445 ;
      RECT 15.5460 16.8810 15.5700 26.3605 ;
      RECT 15.4980 16.8810 15.5220 26.3595 ;
      RECT 15.2100 17.0865 15.2340 26.4155 ;
      RECT 15.1620 17.0875 15.1860 26.4165 ;
      RECT 15.1140 17.0865 15.1380 26.4155 ;
      RECT 15.0180 17.1025 15.0420 26.4165 ;
      RECT 14.8260 17.1015 14.8500 26.3695 ;
      RECT 14.7780 17.1015 14.8020 26.3695 ;
      RECT 14.7300 17.1015 14.7540 26.3695 ;
      RECT 14.6820 17.1015 14.7060 26.3695 ;
      RECT 14.6340 17.1015 14.6580 26.3695 ;
      RECT 14.5860 17.0725 14.6100 26.3695 ;
      RECT 14.5380 17.0285 14.5620 26.0835 ;
      RECT 14.4900 16.9915 14.5140 26.0375 ;
      RECT 14.4420 16.9375 14.4660 25.9835 ;
      RECT 14.3520 21.8825 14.3760 22.0245 ;
      RECT 14.2440 19.8185 14.2680 20.9055 ;
      RECT 14.1840 17.6115 14.2080 21.4555 ;
      RECT 13.8120 19.1945 13.8360 19.4325 ;
  LAYER M2  ;
    RECT 0.108 0.036 30.2400 43.1640 ;
  LAYER M1  ;
    RECT 0.108 0.036 30.2400 43.1640 ;
  END
END srambank_256x4x32_6t122 
