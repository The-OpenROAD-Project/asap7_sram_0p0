VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_128x4x20_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_128x4x20_6t122 0 0 ;
  SIZE 16.0 BY 30.240000000000002 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.1720 16.4420 1.2200 ;
        RECT 0.0940 2.2520 16.4420 2.3000 ;
        RECT 0.0940 3.3320 16.4420 3.3800 ;
        RECT 0.0940 4.4120 16.4420 4.4600 ;
        RECT 0.0940 5.4920 16.4420 5.5400 ;
        RECT 0.0940 6.5720 16.4420 6.6200 ;
        RECT 0.0940 7.6520 16.4420 7.7000 ;
        RECT 0.0940 8.7320 16.4420 8.7800 ;
        RECT 0.0940 9.8120 16.4420 9.8600 ;
        RECT 0.0940 10.8920 16.4420 10.9400 ;
        RECT 3.5640 11.3730 12.9600 11.5890 ;
        RECT 9.1970 14.8770 9.3380 14.9010 ;
        RECT 9.0660 11.0930 9.3290 11.1170 ;
        RECT 7.3980 14.5410 9.1260 14.7570 ;
        RECT 7.3980 17.7090 9.1260 17.9250 ;
        RECT 0.0940 20.0990 16.4420 20.1470 ;
        RECT 0.0940 21.1790 16.4420 21.2270 ;
        RECT 0.0940 22.2590 16.4420 22.3070 ;
        RECT 0.0940 23.3390 16.4420 23.3870 ;
        RECT 0.0940 24.4190 16.4420 24.4670 ;
        RECT 0.0940 25.4990 16.4420 25.5470 ;
        RECT 0.0940 26.5790 16.4420 26.6270 ;
        RECT 0.0940 27.6590 16.4420 27.7070 ;
        RECT 0.0940 28.7390 16.4420 28.7870 ;
        RECT 0.0940 29.8190 16.4420 29.8670 ;
      LAYER M3  ;
        RECT 16.3940 0.2165 16.4120 1.3765 ;
        RECT 9.2840 0.2170 9.3020 1.3760 ;
        RECT 7.8800 0.2570 7.9700 1.3710 ;
        RECT 7.2320 0.2170 7.2500 1.3760 ;
        RECT 0.1220 0.2165 0.1400 1.3765 ;
        RECT 16.3940 1.2965 16.4120 2.4565 ;
        RECT 9.2840 1.2970 9.3020 2.4560 ;
        RECT 7.8800 1.3370 7.9700 2.4510 ;
        RECT 7.2320 1.2970 7.2500 2.4560 ;
        RECT 0.1220 1.2965 0.1400 2.4565 ;
        RECT 16.3940 2.3765 16.4120 3.5365 ;
        RECT 9.2840 2.3770 9.3020 3.5360 ;
        RECT 7.8800 2.4170 7.9700 3.5310 ;
        RECT 7.2320 2.3770 7.2500 3.5360 ;
        RECT 0.1220 2.3765 0.1400 3.5365 ;
        RECT 16.3940 3.4565 16.4120 4.6165 ;
        RECT 9.2840 3.4570 9.3020 4.6160 ;
        RECT 7.8800 3.4970 7.9700 4.6110 ;
        RECT 7.2320 3.4570 7.2500 4.6160 ;
        RECT 0.1220 3.4565 0.1400 4.6165 ;
        RECT 16.3940 4.5365 16.4120 5.6965 ;
        RECT 9.2840 4.5370 9.3020 5.6960 ;
        RECT 7.8800 4.5770 7.9700 5.6910 ;
        RECT 7.2320 4.5370 7.2500 5.6960 ;
        RECT 0.1220 4.5365 0.1400 5.6965 ;
        RECT 16.3940 5.6165 16.4120 6.7765 ;
        RECT 9.2840 5.6170 9.3020 6.7760 ;
        RECT 7.8800 5.6570 7.9700 6.7710 ;
        RECT 7.2320 5.6170 7.2500 6.7760 ;
        RECT 0.1220 5.6165 0.1400 6.7765 ;
        RECT 16.3940 6.6965 16.4120 7.8565 ;
        RECT 9.2840 6.6970 9.3020 7.8560 ;
        RECT 7.8800 6.7370 7.9700 7.8510 ;
        RECT 7.2320 6.6970 7.2500 7.8560 ;
        RECT 0.1220 6.6965 0.1400 7.8565 ;
        RECT 16.3940 7.7765 16.4120 8.9365 ;
        RECT 9.2840 7.7770 9.3020 8.9360 ;
        RECT 7.8800 7.8170 7.9700 8.9310 ;
        RECT 7.2320 7.7770 7.2500 8.9360 ;
        RECT 0.1220 7.7765 0.1400 8.9365 ;
        RECT 16.3940 8.8565 16.4120 10.0165 ;
        RECT 9.2840 8.8570 9.3020 10.0160 ;
        RECT 7.8800 8.8970 7.9700 10.0110 ;
        RECT 7.2320 8.8570 7.2500 10.0160 ;
        RECT 0.1220 8.8565 0.1400 10.0165 ;
        RECT 16.3940 9.9365 16.4120 11.0965 ;
        RECT 9.2840 9.9370 9.3020 11.0960 ;
        RECT 7.8800 9.9770 7.9700 11.0910 ;
        RECT 7.2320 9.9370 7.2500 11.0960 ;
        RECT 0.1220 9.9365 0.1400 11.0965 ;
        RECT 16.3890 11.0105 16.4070 19.2175 ;
        RECT 9.2970 14.8300 9.3150 19.1785 ;
        RECT 9.2790 11.0435 9.2970 11.1815 ;
        RECT 7.9110 11.3340 8.1450 18.9170 ;
        RECT 7.8750 18.8340 7.9650 19.2100 ;
        RECT 7.8750 11.0500 7.9650 11.4260 ;
        RECT 0.1170 11.0105 0.1350 19.2175 ;
        RECT 16.3940 19.1435 16.4120 20.3035 ;
        RECT 9.2840 19.1440 9.3020 20.3030 ;
        RECT 7.8800 19.1840 7.9700 20.2980 ;
        RECT 7.2320 19.1440 7.2500 20.3030 ;
        RECT 0.1220 19.1435 0.1400 20.3035 ;
        RECT 16.3940 20.2235 16.4120 21.3835 ;
        RECT 9.2840 20.2240 9.3020 21.3830 ;
        RECT 7.8800 20.2640 7.9700 21.3780 ;
        RECT 7.2320 20.2240 7.2500 21.3830 ;
        RECT 0.1220 20.2235 0.1400 21.3835 ;
        RECT 16.3940 21.3035 16.4120 22.4635 ;
        RECT 9.2840 21.3040 9.3020 22.4630 ;
        RECT 7.8800 21.3440 7.9700 22.4580 ;
        RECT 7.2320 21.3040 7.2500 22.4630 ;
        RECT 0.1220 21.3035 0.1400 22.4635 ;
        RECT 16.3940 22.3835 16.4120 23.5435 ;
        RECT 9.2840 22.3840 9.3020 23.5430 ;
        RECT 7.8800 22.4240 7.9700 23.5380 ;
        RECT 7.2320 22.3840 7.2500 23.5430 ;
        RECT 0.1220 22.3835 0.1400 23.5435 ;
        RECT 16.3940 23.4635 16.4120 24.6235 ;
        RECT 9.2840 23.4640 9.3020 24.6230 ;
        RECT 7.8800 23.5040 7.9700 24.6180 ;
        RECT 7.2320 23.4640 7.2500 24.6230 ;
        RECT 0.1220 23.4635 0.1400 24.6235 ;
        RECT 16.3940 24.5435 16.4120 25.7035 ;
        RECT 9.2840 24.5440 9.3020 25.7030 ;
        RECT 7.8800 24.5840 7.9700 25.6980 ;
        RECT 7.2320 24.5440 7.2500 25.7030 ;
        RECT 0.1220 24.5435 0.1400 25.7035 ;
        RECT 16.3940 25.6235 16.4120 26.7835 ;
        RECT 9.2840 25.6240 9.3020 26.7830 ;
        RECT 7.8800 25.6640 7.9700 26.7780 ;
        RECT 7.2320 25.6240 7.2500 26.7830 ;
        RECT 0.1220 25.6235 0.1400 26.7835 ;
        RECT 16.3940 26.7035 16.4120 27.8635 ;
        RECT 9.2840 26.7040 9.3020 27.8630 ;
        RECT 7.8800 26.7440 7.9700 27.8580 ;
        RECT 7.2320 26.7040 7.2500 27.8630 ;
        RECT 0.1220 26.7035 0.1400 27.8635 ;
        RECT 16.3940 27.7835 16.4120 28.9435 ;
        RECT 9.2840 27.7840 9.3020 28.9430 ;
        RECT 7.8800 27.8240 7.9700 28.9380 ;
        RECT 7.2320 27.7840 7.2500 28.9430 ;
        RECT 0.1220 27.7835 0.1400 28.9435 ;
        RECT 16.3940 28.8635 16.4120 30.0235 ;
        RECT 9.2840 28.8640 9.3020 30.0230 ;
        RECT 7.8800 28.9040 7.9700 30.0180 ;
        RECT 7.2320 28.8640 7.2500 30.0230 ;
        RECT 0.1220 28.8635 0.1400 30.0235 ;
      LAYER V3  ;
        RECT 0.1220 1.1720 0.1400 1.2200 ;
        RECT 7.2320 1.1720 7.2500 1.2200 ;
        RECT 7.8800 1.1720 7.9700 1.2200 ;
        RECT 9.2840 1.1720 9.3020 1.2200 ;
        RECT 16.3940 1.1720 16.4120 1.2200 ;
        RECT 0.1220 2.2520 0.1400 2.3000 ;
        RECT 7.2320 2.2520 7.2500 2.3000 ;
        RECT 7.8800 2.2520 7.9700 2.3000 ;
        RECT 9.2840 2.2520 9.3020 2.3000 ;
        RECT 16.3940 2.2520 16.4120 2.3000 ;
        RECT 0.1220 3.3320 0.1400 3.3800 ;
        RECT 7.2320 3.3320 7.2500 3.3800 ;
        RECT 7.8800 3.3320 7.9700 3.3800 ;
        RECT 9.2840 3.3320 9.3020 3.3800 ;
        RECT 16.3940 3.3320 16.4120 3.3800 ;
        RECT 0.1220 4.4120 0.1400 4.4600 ;
        RECT 7.2320 4.4120 7.2500 4.4600 ;
        RECT 7.8800 4.4120 7.9700 4.4600 ;
        RECT 9.2840 4.4120 9.3020 4.4600 ;
        RECT 16.3940 4.4120 16.4120 4.4600 ;
        RECT 0.1220 5.4920 0.1400 5.5400 ;
        RECT 7.2320 5.4920 7.2500 5.5400 ;
        RECT 7.8800 5.4920 7.9700 5.5400 ;
        RECT 9.2840 5.4920 9.3020 5.5400 ;
        RECT 16.3940 5.4920 16.4120 5.5400 ;
        RECT 0.1220 6.5720 0.1400 6.6200 ;
        RECT 7.2320 6.5720 7.2500 6.6200 ;
        RECT 7.8800 6.5720 7.9700 6.6200 ;
        RECT 9.2840 6.5720 9.3020 6.6200 ;
        RECT 16.3940 6.5720 16.4120 6.6200 ;
        RECT 0.1220 7.6520 0.1400 7.7000 ;
        RECT 7.2320 7.6520 7.2500 7.7000 ;
        RECT 7.8800 7.6520 7.9700 7.7000 ;
        RECT 9.2840 7.6520 9.3020 7.7000 ;
        RECT 16.3940 7.6520 16.4120 7.7000 ;
        RECT 0.1220 8.7320 0.1400 8.7800 ;
        RECT 7.2320 8.7320 7.2500 8.7800 ;
        RECT 7.8800 8.7320 7.9700 8.7800 ;
        RECT 9.2840 8.7320 9.3020 8.7800 ;
        RECT 16.3940 8.7320 16.4120 8.7800 ;
        RECT 0.1220 9.8120 0.1400 9.8600 ;
        RECT 7.2320 9.8120 7.2500 9.8600 ;
        RECT 7.8800 9.8120 7.9700 9.8600 ;
        RECT 9.2840 9.8120 9.3020 9.8600 ;
        RECT 16.3940 9.8120 16.4120 9.8600 ;
        RECT 0.1220 10.8920 0.1400 10.9400 ;
        RECT 7.2320 10.8920 7.2500 10.9400 ;
        RECT 7.8800 10.8920 7.9700 10.9400 ;
        RECT 9.2840 10.8920 9.3020 10.9400 ;
        RECT 16.3940 10.8920 16.4120 10.9400 ;
        RECT 7.9150 17.7090 7.9330 17.9250 ;
        RECT 7.9150 14.5410 7.9330 14.7570 ;
        RECT 7.9150 11.3730 7.9330 11.5890 ;
        RECT 7.9670 17.7090 7.9850 17.9250 ;
        RECT 7.9670 14.5410 7.9850 14.7570 ;
        RECT 7.9670 11.3730 7.9850 11.5890 ;
        RECT 8.0190 17.7090 8.0370 17.9250 ;
        RECT 8.0190 14.5410 8.0370 14.7570 ;
        RECT 8.0190 11.3730 8.0370 11.5890 ;
        RECT 8.0710 17.7090 8.0890 17.9250 ;
        RECT 8.0710 14.5410 8.0890 14.7570 ;
        RECT 8.0710 11.3730 8.0890 11.5890 ;
        RECT 8.1230 17.7090 8.1410 17.9250 ;
        RECT 8.1230 14.5410 8.1410 14.7570 ;
        RECT 8.1230 11.3730 8.1410 11.5890 ;
        RECT 9.2790 11.0930 9.2970 11.1170 ;
        RECT 9.2970 14.8770 9.3150 14.9010 ;
        RECT 0.1220 20.0990 0.1400 20.1470 ;
        RECT 7.2320 20.0990 7.2500 20.1470 ;
        RECT 7.8800 20.0990 7.9700 20.1470 ;
        RECT 9.2840 20.0990 9.3020 20.1470 ;
        RECT 16.3940 20.0990 16.4120 20.1470 ;
        RECT 0.1220 21.1790 0.1400 21.2270 ;
        RECT 7.2320 21.1790 7.2500 21.2270 ;
        RECT 7.8800 21.1790 7.9700 21.2270 ;
        RECT 9.2840 21.1790 9.3020 21.2270 ;
        RECT 16.3940 21.1790 16.4120 21.2270 ;
        RECT 0.1220 22.2590 0.1400 22.3070 ;
        RECT 7.2320 22.2590 7.2500 22.3070 ;
        RECT 7.8800 22.2590 7.9700 22.3070 ;
        RECT 9.2840 22.2590 9.3020 22.3070 ;
        RECT 16.3940 22.2590 16.4120 22.3070 ;
        RECT 0.1220 23.3390 0.1400 23.3870 ;
        RECT 7.2320 23.3390 7.2500 23.3870 ;
        RECT 7.8800 23.3390 7.9700 23.3870 ;
        RECT 9.2840 23.3390 9.3020 23.3870 ;
        RECT 16.3940 23.3390 16.4120 23.3870 ;
        RECT 0.1220 24.4190 0.1400 24.4670 ;
        RECT 7.2320 24.4190 7.2500 24.4670 ;
        RECT 7.8800 24.4190 7.9700 24.4670 ;
        RECT 9.2840 24.4190 9.3020 24.4670 ;
        RECT 16.3940 24.4190 16.4120 24.4670 ;
        RECT 0.1220 25.4990 0.1400 25.5470 ;
        RECT 7.2320 25.4990 7.2500 25.5470 ;
        RECT 7.8800 25.4990 7.9700 25.5470 ;
        RECT 9.2840 25.4990 9.3020 25.5470 ;
        RECT 16.3940 25.4990 16.4120 25.5470 ;
        RECT 0.1220 26.5790 0.1400 26.6270 ;
        RECT 7.2320 26.5790 7.2500 26.6270 ;
        RECT 7.8800 26.5790 7.9700 26.6270 ;
        RECT 9.2840 26.5790 9.3020 26.6270 ;
        RECT 16.3940 26.5790 16.4120 26.6270 ;
        RECT 0.1220 27.6590 0.1400 27.7070 ;
        RECT 7.2320 27.6590 7.2500 27.7070 ;
        RECT 7.8800 27.6590 7.9700 27.7070 ;
        RECT 9.2840 27.6590 9.3020 27.7070 ;
        RECT 16.3940 27.6590 16.4120 27.7070 ;
        RECT 0.1220 28.7390 0.1400 28.7870 ;
        RECT 7.2320 28.7390 7.2500 28.7870 ;
        RECT 7.8800 28.7390 7.9700 28.7870 ;
        RECT 9.2840 28.7390 9.3020 28.7870 ;
        RECT 16.3940 28.7390 16.4120 28.7870 ;
        RECT 0.1220 29.8190 0.1400 29.8670 ;
        RECT 7.2320 29.8190 7.2500 29.8670 ;
        RECT 7.8800 29.8190 7.9700 29.8670 ;
        RECT 9.2840 29.8190 9.3020 29.8670 ;
        RECT 16.3940 29.8190 16.4120 29.8670 ;
      LAYER M5  ;
        RECT 9.2160 11.0750 9.2400 14.9190 ;
      LAYER V4  ;
        RECT 9.2160 14.8770 9.2400 14.9010 ;
        RECT 9.2160 11.3730 9.2400 11.5890 ;
        RECT 9.2160 11.0930 9.2400 11.1170 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.0760 16.4370 1.1240 ;
        RECT 0.0940 2.1560 16.4370 2.2040 ;
        RECT 0.0940 3.2360 16.4370 3.2840 ;
        RECT 0.0940 4.3160 16.4370 4.3640 ;
        RECT 0.0940 5.3960 16.4370 5.4440 ;
        RECT 0.0940 6.4760 16.4370 6.5240 ;
        RECT 0.0940 7.5560 16.4370 7.6040 ;
        RECT 0.0940 8.6360 16.4370 8.6840 ;
        RECT 0.0940 9.7160 16.4370 9.7640 ;
        RECT 0.0940 10.7960 16.4370 10.8440 ;
        RECT 3.5640 11.8050 12.9600 12.0210 ;
        RECT 7.3980 14.9730 9.1260 15.1890 ;
        RECT 7.3980 18.1410 9.1260 18.3570 ;
        RECT 0.0940 20.0030 16.4370 20.0510 ;
        RECT 0.0940 21.0830 16.4370 21.1310 ;
        RECT 0.0940 22.1630 16.4370 22.2110 ;
        RECT 0.0940 23.2430 16.4370 23.2910 ;
        RECT 0.0940 24.3230 16.4370 24.3710 ;
        RECT 0.0940 25.4030 16.4370 25.4510 ;
        RECT 0.0940 26.4830 16.4370 26.5310 ;
        RECT 0.0940 27.5630 16.4370 27.6110 ;
        RECT 0.0940 28.6430 16.4370 28.6910 ;
        RECT 0.0940 29.7230 16.4370 29.7710 ;
      LAYER M3  ;
        RECT 16.3580 0.2165 16.3760 1.3765 ;
        RECT 9.3380 0.2165 9.3560 1.3765 ;
        RECT 8.5730 0.2530 8.6090 1.3670 ;
        RECT 8.4200 0.2530 8.4470 1.3670 ;
        RECT 7.1780 0.2165 7.1960 1.3765 ;
        RECT 0.1580 0.2165 0.1760 1.3765 ;
        RECT 16.3580 1.2965 16.3760 2.4565 ;
        RECT 9.3380 1.2965 9.3560 2.4565 ;
        RECT 8.5730 1.3330 8.6090 2.4470 ;
        RECT 8.4200 1.3330 8.4470 2.4470 ;
        RECT 7.1780 1.2965 7.1960 2.4565 ;
        RECT 0.1580 1.2965 0.1760 2.4565 ;
        RECT 16.3580 2.3765 16.3760 3.5365 ;
        RECT 9.3380 2.3765 9.3560 3.5365 ;
        RECT 8.5730 2.4130 8.6090 3.5270 ;
        RECT 8.4200 2.4130 8.4470 3.5270 ;
        RECT 7.1780 2.3765 7.1960 3.5365 ;
        RECT 0.1580 2.3765 0.1760 3.5365 ;
        RECT 16.3580 3.4565 16.3760 4.6165 ;
        RECT 9.3380 3.4565 9.3560 4.6165 ;
        RECT 8.5730 3.4930 8.6090 4.6070 ;
        RECT 8.4200 3.4930 8.4470 4.6070 ;
        RECT 7.1780 3.4565 7.1960 4.6165 ;
        RECT 0.1580 3.4565 0.1760 4.6165 ;
        RECT 16.3580 4.5365 16.3760 5.6965 ;
        RECT 9.3380 4.5365 9.3560 5.6965 ;
        RECT 8.5730 4.5730 8.6090 5.6870 ;
        RECT 8.4200 4.5730 8.4470 5.6870 ;
        RECT 7.1780 4.5365 7.1960 5.6965 ;
        RECT 0.1580 4.5365 0.1760 5.6965 ;
        RECT 16.3580 5.6165 16.3760 6.7765 ;
        RECT 9.3380 5.6165 9.3560 6.7765 ;
        RECT 8.5730 5.6530 8.6090 6.7670 ;
        RECT 8.4200 5.6530 8.4470 6.7670 ;
        RECT 7.1780 5.6165 7.1960 6.7765 ;
        RECT 0.1580 5.6165 0.1760 6.7765 ;
        RECT 16.3580 6.6965 16.3760 7.8565 ;
        RECT 9.3380 6.6965 9.3560 7.8565 ;
        RECT 8.5730 6.7330 8.6090 7.8470 ;
        RECT 8.4200 6.7330 8.4470 7.8470 ;
        RECT 7.1780 6.6965 7.1960 7.8565 ;
        RECT 0.1580 6.6965 0.1760 7.8565 ;
        RECT 16.3580 7.7765 16.3760 8.9365 ;
        RECT 9.3380 7.7765 9.3560 8.9365 ;
        RECT 8.5730 7.8130 8.6090 8.9270 ;
        RECT 8.4200 7.8130 8.4470 8.9270 ;
        RECT 7.1780 7.7765 7.1960 8.9365 ;
        RECT 0.1580 7.7765 0.1760 8.9365 ;
        RECT 16.3580 8.8565 16.3760 10.0165 ;
        RECT 9.3380 8.8565 9.3560 10.0165 ;
        RECT 8.5730 8.8930 8.6090 10.0070 ;
        RECT 8.4200 8.8930 8.4470 10.0070 ;
        RECT 7.1780 8.8565 7.1960 10.0165 ;
        RECT 0.1580 8.8565 0.1760 10.0165 ;
        RECT 16.3580 9.9365 16.3760 11.0965 ;
        RECT 9.3380 9.9365 9.3560 11.0965 ;
        RECT 8.5730 9.9730 8.6090 11.0870 ;
        RECT 8.4200 9.9730 8.4470 11.0870 ;
        RECT 7.1780 9.9365 7.1960 11.0965 ;
        RECT 0.1580 9.9365 0.1760 11.0965 ;
        RECT 16.3530 11.0105 16.3710 19.2175 ;
        RECT 9.3330 11.0105 9.3510 19.2175 ;
        RECT 8.3790 11.2340 8.6130 18.9170 ;
        RECT 8.5680 11.0545 8.6040 19.1740 ;
        RECT 8.4150 11.0540 8.4420 19.1740 ;
        RECT 7.1730 11.0105 7.1910 19.2175 ;
        RECT 0.1530 11.0105 0.1710 19.2175 ;
        RECT 16.3580 19.1435 16.3760 20.3035 ;
        RECT 9.3380 19.1435 9.3560 20.3035 ;
        RECT 8.5730 19.1800 8.6090 20.2940 ;
        RECT 8.4200 19.1800 8.4470 20.2940 ;
        RECT 7.1780 19.1435 7.1960 20.3035 ;
        RECT 0.1580 19.1435 0.1760 20.3035 ;
        RECT 16.3580 20.2235 16.3760 21.3835 ;
        RECT 9.3380 20.2235 9.3560 21.3835 ;
        RECT 8.5730 20.2600 8.6090 21.3740 ;
        RECT 8.4200 20.2600 8.4470 21.3740 ;
        RECT 7.1780 20.2235 7.1960 21.3835 ;
        RECT 0.1580 20.2235 0.1760 21.3835 ;
        RECT 16.3580 21.3035 16.3760 22.4635 ;
        RECT 9.3380 21.3035 9.3560 22.4635 ;
        RECT 8.5730 21.3400 8.6090 22.4540 ;
        RECT 8.4200 21.3400 8.4470 22.4540 ;
        RECT 7.1780 21.3035 7.1960 22.4635 ;
        RECT 0.1580 21.3035 0.1760 22.4635 ;
        RECT 16.3580 22.3835 16.3760 23.5435 ;
        RECT 9.3380 22.3835 9.3560 23.5435 ;
        RECT 8.5730 22.4200 8.6090 23.5340 ;
        RECT 8.4200 22.4200 8.4470 23.5340 ;
        RECT 7.1780 22.3835 7.1960 23.5435 ;
        RECT 0.1580 22.3835 0.1760 23.5435 ;
        RECT 16.3580 23.4635 16.3760 24.6235 ;
        RECT 9.3380 23.4635 9.3560 24.6235 ;
        RECT 8.5730 23.5000 8.6090 24.6140 ;
        RECT 8.4200 23.5000 8.4470 24.6140 ;
        RECT 7.1780 23.4635 7.1960 24.6235 ;
        RECT 0.1580 23.4635 0.1760 24.6235 ;
        RECT 16.3580 24.5435 16.3760 25.7035 ;
        RECT 9.3380 24.5435 9.3560 25.7035 ;
        RECT 8.5730 24.5800 8.6090 25.6940 ;
        RECT 8.4200 24.5800 8.4470 25.6940 ;
        RECT 7.1780 24.5435 7.1960 25.7035 ;
        RECT 0.1580 24.5435 0.1760 25.7035 ;
        RECT 16.3580 25.6235 16.3760 26.7835 ;
        RECT 9.3380 25.6235 9.3560 26.7835 ;
        RECT 8.5730 25.6600 8.6090 26.7740 ;
        RECT 8.4200 25.6600 8.4470 26.7740 ;
        RECT 7.1780 25.6235 7.1960 26.7835 ;
        RECT 0.1580 25.6235 0.1760 26.7835 ;
        RECT 16.3580 26.7035 16.3760 27.8635 ;
        RECT 9.3380 26.7035 9.3560 27.8635 ;
        RECT 8.5730 26.7400 8.6090 27.8540 ;
        RECT 8.4200 26.7400 8.4470 27.8540 ;
        RECT 7.1780 26.7035 7.1960 27.8635 ;
        RECT 0.1580 26.7035 0.1760 27.8635 ;
        RECT 16.3580 27.7835 16.3760 28.9435 ;
        RECT 9.3380 27.7835 9.3560 28.9435 ;
        RECT 8.5730 27.8200 8.6090 28.9340 ;
        RECT 8.4200 27.8200 8.4470 28.9340 ;
        RECT 7.1780 27.7835 7.1960 28.9435 ;
        RECT 0.1580 27.7835 0.1760 28.9435 ;
        RECT 16.3580 28.8635 16.3760 30.0235 ;
        RECT 9.3380 28.8635 9.3560 30.0235 ;
        RECT 8.5730 28.9000 8.6090 30.0140 ;
        RECT 8.4200 28.9000 8.4470 30.0140 ;
        RECT 7.1780 28.8635 7.1960 30.0235 ;
        RECT 0.1580 28.8635 0.1760 30.0235 ;
      LAYER V3  ;
        RECT 0.1580 1.0760 0.1760 1.1240 ;
        RECT 7.1780 1.0760 7.1960 1.1240 ;
        RECT 8.4200 1.0760 8.4470 1.1240 ;
        RECT 8.5730 1.0760 8.6090 1.1240 ;
        RECT 9.3380 1.0760 9.3560 1.1240 ;
        RECT 16.3580 1.0760 16.3760 1.1240 ;
        RECT 0.1580 2.1560 0.1760 2.2040 ;
        RECT 7.1780 2.1560 7.1960 2.2040 ;
        RECT 8.4200 2.1560 8.4470 2.2040 ;
        RECT 8.5730 2.1560 8.6090 2.2040 ;
        RECT 9.3380 2.1560 9.3560 2.2040 ;
        RECT 16.3580 2.1560 16.3760 2.2040 ;
        RECT 0.1580 3.2360 0.1760 3.2840 ;
        RECT 7.1780 3.2360 7.1960 3.2840 ;
        RECT 8.4200 3.2360 8.4470 3.2840 ;
        RECT 8.5730 3.2360 8.6090 3.2840 ;
        RECT 9.3380 3.2360 9.3560 3.2840 ;
        RECT 16.3580 3.2360 16.3760 3.2840 ;
        RECT 0.1580 4.3160 0.1760 4.3640 ;
        RECT 7.1780 4.3160 7.1960 4.3640 ;
        RECT 8.4200 4.3160 8.4470 4.3640 ;
        RECT 8.5730 4.3160 8.6090 4.3640 ;
        RECT 9.3380 4.3160 9.3560 4.3640 ;
        RECT 16.3580 4.3160 16.3760 4.3640 ;
        RECT 0.1580 5.3960 0.1760 5.4440 ;
        RECT 7.1780 5.3960 7.1960 5.4440 ;
        RECT 8.4200 5.3960 8.4470 5.4440 ;
        RECT 8.5730 5.3960 8.6090 5.4440 ;
        RECT 9.3380 5.3960 9.3560 5.4440 ;
        RECT 16.3580 5.3960 16.3760 5.4440 ;
        RECT 0.1580 6.4760 0.1760 6.5240 ;
        RECT 7.1780 6.4760 7.1960 6.5240 ;
        RECT 8.4200 6.4760 8.4470 6.5240 ;
        RECT 8.5730 6.4760 8.6090 6.5240 ;
        RECT 9.3380 6.4760 9.3560 6.5240 ;
        RECT 16.3580 6.4760 16.3760 6.5240 ;
        RECT 0.1580 7.5560 0.1760 7.6040 ;
        RECT 7.1780 7.5560 7.1960 7.6040 ;
        RECT 8.4200 7.5560 8.4470 7.6040 ;
        RECT 8.5730 7.5560 8.6090 7.6040 ;
        RECT 9.3380 7.5560 9.3560 7.6040 ;
        RECT 16.3580 7.5560 16.3760 7.6040 ;
        RECT 0.1580 8.6360 0.1760 8.6840 ;
        RECT 7.1780 8.6360 7.1960 8.6840 ;
        RECT 8.4200 8.6360 8.4470 8.6840 ;
        RECT 8.5730 8.6360 8.6090 8.6840 ;
        RECT 9.3380 8.6360 9.3560 8.6840 ;
        RECT 16.3580 8.6360 16.3760 8.6840 ;
        RECT 0.1580 9.7160 0.1760 9.7640 ;
        RECT 7.1780 9.7160 7.1960 9.7640 ;
        RECT 8.4200 9.7160 8.4470 9.7640 ;
        RECT 8.5730 9.7160 8.6090 9.7640 ;
        RECT 9.3380 9.7160 9.3560 9.7640 ;
        RECT 16.3580 9.7160 16.3760 9.7640 ;
        RECT 0.1580 10.7960 0.1760 10.8440 ;
        RECT 7.1780 10.7960 7.1960 10.8440 ;
        RECT 8.4200 10.7960 8.4470 10.8440 ;
        RECT 8.5730 10.7960 8.6090 10.8440 ;
        RECT 9.3380 10.7960 9.3560 10.8440 ;
        RECT 16.3580 10.7960 16.3760 10.8440 ;
        RECT 8.3830 18.1410 8.4010 18.3570 ;
        RECT 8.3830 14.9730 8.4010 15.1890 ;
        RECT 8.3830 11.8050 8.4010 12.0210 ;
        RECT 8.4350 18.1410 8.4530 18.3570 ;
        RECT 8.4350 14.9730 8.4530 15.1890 ;
        RECT 8.4350 11.8050 8.4530 12.0210 ;
        RECT 8.4870 18.1410 8.5050 18.3570 ;
        RECT 8.4870 14.9730 8.5050 15.1890 ;
        RECT 8.4870 11.8050 8.5050 12.0210 ;
        RECT 8.5390 18.1410 8.5570 18.3570 ;
        RECT 8.5390 14.9730 8.5570 15.1890 ;
        RECT 8.5390 11.8050 8.5570 12.0210 ;
        RECT 8.5910 18.1410 8.6090 18.3570 ;
        RECT 8.5910 14.9730 8.6090 15.1890 ;
        RECT 8.5910 11.8050 8.6090 12.0210 ;
        RECT 9.3330 11.8055 9.3510 12.0215 ;
        RECT 0.1580 20.0030 0.1760 20.0510 ;
        RECT 7.1780 20.0030 7.1960 20.0510 ;
        RECT 8.4200 20.0030 8.4470 20.0510 ;
        RECT 8.5730 20.0030 8.6090 20.0510 ;
        RECT 9.3380 20.0030 9.3560 20.0510 ;
        RECT 16.3580 20.0030 16.3760 20.0510 ;
        RECT 0.1580 21.0830 0.1760 21.1310 ;
        RECT 7.1780 21.0830 7.1960 21.1310 ;
        RECT 8.4200 21.0830 8.4470 21.1310 ;
        RECT 8.5730 21.0830 8.6090 21.1310 ;
        RECT 9.3380 21.0830 9.3560 21.1310 ;
        RECT 16.3580 21.0830 16.3760 21.1310 ;
        RECT 0.1580 22.1630 0.1760 22.2110 ;
        RECT 7.1780 22.1630 7.1960 22.2110 ;
        RECT 8.4200 22.1630 8.4470 22.2110 ;
        RECT 8.5730 22.1630 8.6090 22.2110 ;
        RECT 9.3380 22.1630 9.3560 22.2110 ;
        RECT 16.3580 22.1630 16.3760 22.2110 ;
        RECT 0.1580 23.2430 0.1760 23.2910 ;
        RECT 7.1780 23.2430 7.1960 23.2910 ;
        RECT 8.4200 23.2430 8.4470 23.2910 ;
        RECT 8.5730 23.2430 8.6090 23.2910 ;
        RECT 9.3380 23.2430 9.3560 23.2910 ;
        RECT 16.3580 23.2430 16.3760 23.2910 ;
        RECT 0.1580 24.3230 0.1760 24.3710 ;
        RECT 7.1780 24.3230 7.1960 24.3710 ;
        RECT 8.4200 24.3230 8.4470 24.3710 ;
        RECT 8.5730 24.3230 8.6090 24.3710 ;
        RECT 9.3380 24.3230 9.3560 24.3710 ;
        RECT 16.3580 24.3230 16.3760 24.3710 ;
        RECT 0.1580 25.4030 0.1760 25.4510 ;
        RECT 7.1780 25.4030 7.1960 25.4510 ;
        RECT 8.4200 25.4030 8.4470 25.4510 ;
        RECT 8.5730 25.4030 8.6090 25.4510 ;
        RECT 9.3380 25.4030 9.3560 25.4510 ;
        RECT 16.3580 25.4030 16.3760 25.4510 ;
        RECT 0.1580 26.4830 0.1760 26.5310 ;
        RECT 7.1780 26.4830 7.1960 26.5310 ;
        RECT 8.4200 26.4830 8.4470 26.5310 ;
        RECT 8.5730 26.4830 8.6090 26.5310 ;
        RECT 9.3380 26.4830 9.3560 26.5310 ;
        RECT 16.3580 26.4830 16.3760 26.5310 ;
        RECT 0.1580 27.5630 0.1760 27.6110 ;
        RECT 7.1780 27.5630 7.1960 27.6110 ;
        RECT 8.4200 27.5630 8.4470 27.6110 ;
        RECT 8.5730 27.5630 8.6090 27.6110 ;
        RECT 9.3380 27.5630 9.3560 27.6110 ;
        RECT 16.3580 27.5630 16.3760 27.6110 ;
        RECT 0.1580 28.6430 0.1760 28.6910 ;
        RECT 7.1780 28.6430 7.1960 28.6910 ;
        RECT 8.4200 28.6430 8.4470 28.6910 ;
        RECT 8.5730 28.6430 8.6090 28.6910 ;
        RECT 9.3380 28.6430 9.3560 28.6910 ;
        RECT 16.3580 28.6430 16.3760 28.6910 ;
        RECT 0.1580 29.7230 0.1760 29.7710 ;
        RECT 7.1780 29.7230 7.1960 29.7710 ;
        RECT 8.4200 29.7230 8.4470 29.7710 ;
        RECT 8.5730 29.7230 8.6090 29.7710 ;
        RECT 9.3380 29.7230 9.3560 29.7710 ;
        RECT 16.3580 29.7230 16.3760 29.7710 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.7910 12.2770 10.8090 12.3140 ;
      LAYER M4  ;
        RECT 10.7390 12.2850 10.8230 12.3090 ;
      LAYER M5  ;
        RECT 10.7880 11.3340 10.8120 14.5740 ;
      LAYER V3  ;
        RECT 10.7910 12.2850 10.8090 12.3090 ;
      LAYER V4  ;
        RECT 10.7880 12.2850 10.8120 12.3090 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.5750 12.2800 10.5930 12.3170 ;
      LAYER M4  ;
        RECT 10.5230 12.2850 10.6070 12.3090 ;
      LAYER M5  ;
        RECT 10.5720 11.3340 10.5960 14.5740 ;
      LAYER V3  ;
        RECT 10.5750 12.2850 10.5930 12.3090 ;
      LAYER V4  ;
        RECT 10.5720 12.2850 10.5960 12.3090 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.3590 11.7010 10.3770 11.7380 ;
      LAYER M4  ;
        RECT 10.3070 11.7090 10.3910 11.7330 ;
      LAYER M5  ;
        RECT 10.3560 11.3340 10.3800 14.5740 ;
      LAYER V3  ;
        RECT 10.3590 11.7090 10.3770 11.7330 ;
      LAYER V4  ;
        RECT 10.3560 11.7090 10.3800 11.7330 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.1430 11.9410 10.1610 12.1220 ;
      LAYER M4  ;
        RECT 10.0910 12.0930 10.1750 12.1170 ;
      LAYER M5  ;
        RECT 10.1400 11.3340 10.1640 14.5740 ;
      LAYER V3  ;
        RECT 10.1430 12.0930 10.1610 12.1170 ;
      LAYER V4  ;
        RECT 10.1400 12.0930 10.1640 12.1170 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.9270 11.7040 9.9450 11.7710 ;
      LAYER M4  ;
        RECT 9.8750 11.7090 9.9590 11.7330 ;
      LAYER M5  ;
        RECT 9.9240 11.3340 9.9480 14.5740 ;
      LAYER V3  ;
        RECT 9.9270 11.7090 9.9450 11.7330 ;
      LAYER V4  ;
        RECT 9.9240 11.7090 9.9480 11.7330 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.7110 11.4370 9.7290 11.6900 ;
      LAYER M4  ;
        RECT 9.6590 11.6610 9.7430 11.6850 ;
      LAYER M5  ;
        RECT 9.7080 11.3340 9.7320 14.5740 ;
      LAYER V3  ;
        RECT 9.7110 11.6610 9.7290 11.6850 ;
      LAYER V4  ;
        RECT 9.7080 11.6610 9.7320 11.6850 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.4950 12.4720 9.5130 12.5090 ;
      LAYER M4  ;
        RECT 9.4430 12.4770 9.5270 12.5010 ;
      LAYER M5  ;
        RECT 9.4920 11.3340 9.5160 14.5740 ;
      LAYER V3  ;
        RECT 9.4950 12.4770 9.5130 12.5010 ;
      LAYER V4  ;
        RECT 9.4920 12.4770 9.5160 12.5010 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.2790 12.3190 9.2970 12.4100 ;
      LAYER M4  ;
        RECT 9.2270 12.3810 9.3110 12.4050 ;
      LAYER M5  ;
        RECT 9.2760 11.3340 9.3000 14.5740 ;
      LAYER V3  ;
        RECT 9.2790 12.3810 9.2970 12.4050 ;
      LAYER V4  ;
        RECT 9.2760 12.3810 9.3000 12.4050 ;
    END
  END ADDRESS[7]
  PIN ADDRESS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.6310 11.7040 8.6490 11.7710 ;
      LAYER M4  ;
        RECT 8.3470 11.7090 8.6600 11.7330 ;
      LAYER M5  ;
        RECT 8.3580 11.3340 8.3820 14.5740 ;
      LAYER V3  ;
        RECT 8.6310 11.7090 8.6490 11.7330 ;
      LAYER V4  ;
        RECT 8.3580 11.7090 8.3820 11.7330 ;
    END
  END ADDRESS[8]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.2350 11.4370 8.2530 11.6900 ;
      LAYER M4  ;
        RECT 8.0230 11.6610 8.2640 11.6850 ;
      LAYER M5  ;
        RECT 8.0340 11.3340 8.0580 14.5740 ;
      LAYER V3  ;
        RECT 8.2350 11.6610 8.2530 11.6850 ;
      LAYER V4  ;
        RECT 8.0340 11.6610 8.0580 11.6850 ;
    END
  END banksel
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.4430 11.7040 7.4610 11.7710 ;
      LAYER M4  ;
        RECT 7.3910 11.7090 7.4750 11.7330 ;
      LAYER M5  ;
        RECT 7.4400 11.3340 7.4640 14.5740 ;
      LAYER V3  ;
        RECT 7.4430 11.7090 7.4610 11.7330 ;
      LAYER V4  ;
        RECT 7.4400 11.7090 7.4640 11.7330 ;
    END
  END write
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2270 12.5680 7.2450 12.6170 ;
      LAYER M4  ;
        RECT 7.1750 12.5730 7.2590 12.5970 ;
      LAYER M5  ;
        RECT 7.2240 11.3340 7.2480 14.5740 ;
      LAYER V3  ;
        RECT 7.2270 12.5730 7.2450 12.5970 ;
      LAYER V4  ;
        RECT 7.2240 12.5730 7.2480 12.5970 ;
    END
  END clk
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2630 11.4370 7.2810 11.6900 ;
      LAYER M4  ;
        RECT 6.9970 11.6610 7.2920 11.6850 ;
      LAYER M5  ;
        RECT 7.0080 11.3340 7.0320 14.5740 ;
      LAYER V3  ;
        RECT 7.2630 11.6610 7.2810 11.6850 ;
      LAYER V4  ;
        RECT 7.0080 11.6610 7.0320 11.6850 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.7950 12.2770 6.8130 12.3140 ;
      LAYER M4  ;
        RECT 6.7430 12.2850 6.8270 12.3090 ;
      LAYER M5  ;
        RECT 6.7920 11.3340 6.8160 14.5740 ;
      LAYER V3  ;
        RECT 6.7950 12.2850 6.8130 12.3090 ;
      LAYER V4  ;
        RECT 6.7920 12.2850 6.8160 12.3090 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.5790 11.7040 6.5970 11.9330 ;
      LAYER M4  ;
        RECT 6.5270 11.7090 6.6110 11.7330 ;
      LAYER M5  ;
        RECT 6.5760 11.3340 6.6000 14.5740 ;
      LAYER V3  ;
        RECT 6.5790 11.7090 6.5970 11.7330 ;
      LAYER V4  ;
        RECT 6.5760 11.7090 6.6000 11.7330 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.3630 11.4370 6.3810 11.6900 ;
      LAYER M4  ;
        RECT 6.3110 11.6610 6.3950 11.6850 ;
      LAYER M5  ;
        RECT 6.3600 11.3340 6.3840 14.5740 ;
      LAYER V3  ;
        RECT 6.3630 11.6610 6.3810 11.6850 ;
      LAYER V4  ;
        RECT 6.3600 11.6610 6.3840 11.6850 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.1470 11.7010 6.1650 11.7380 ;
      LAYER M4  ;
        RECT 6.0950 11.7090 6.1790 11.7330 ;
      LAYER M5  ;
        RECT 6.1440 11.3340 6.1680 14.5740 ;
      LAYER V3  ;
        RECT 6.1470 11.7090 6.1650 11.7330 ;
      LAYER V4  ;
        RECT 6.1440 11.7090 6.1680 11.7330 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 5.9310 12.2770 5.9490 12.3140 ;
      LAYER M4  ;
        RECT 5.8790 12.2850 5.9630 12.3090 ;
      LAYER M5  ;
        RECT 5.9280 11.3340 5.9520 14.5740 ;
      LAYER V3  ;
        RECT 5.9310 12.2850 5.9490 12.3090 ;
      LAYER V4  ;
        RECT 5.9280 12.2850 5.9520 12.3090 ;
    END
  END sdel[4]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.4280 8.5970 0.4520 ;
      LAYER M3  ;
        RECT 8.5370 0.3775 8.5550 0.6170 ;
      LAYER V3  ;
        RECT 8.5370 0.4280 8.5550 0.4520 ;
    END
  END dataout[0]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.3320 8.6650 0.3560 ;
      LAYER M3  ;
        RECT 8.3120 0.2700 8.3300 0.6750 ;
      LAYER V3  ;
        RECT 8.3120 0.3320 8.3300 0.3560 ;
    END
  END wd[0]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.5080 8.5970 1.5320 ;
      LAYER M3  ;
        RECT 8.5370 1.4575 8.5550 1.6970 ;
      LAYER V3  ;
        RECT 8.5370 1.5080 8.5550 1.5320 ;
    END
  END dataout[1]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.4120 8.6650 1.4360 ;
      LAYER M3  ;
        RECT 8.3120 1.3500 8.3300 1.7550 ;
      LAYER V3  ;
        RECT 8.3120 1.4120 8.3300 1.4360 ;
    END
  END wd[1]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.5880 8.5970 2.6120 ;
      LAYER M3  ;
        RECT 8.5370 2.5375 8.5550 2.7770 ;
      LAYER V3  ;
        RECT 8.5370 2.5880 8.5550 2.6120 ;
    END
  END dataout[2]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.4920 8.6650 2.5160 ;
      LAYER M3  ;
        RECT 8.3120 2.4300 8.3300 2.8350 ;
      LAYER V3  ;
        RECT 8.3120 2.4920 8.3300 2.5160 ;
    END
  END wd[2]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.6680 8.5970 3.6920 ;
      LAYER M3  ;
        RECT 8.5370 3.6175 8.5550 3.8570 ;
      LAYER V3  ;
        RECT 8.5370 3.6680 8.5550 3.6920 ;
    END
  END dataout[3]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.5720 8.6650 3.5960 ;
      LAYER M3  ;
        RECT 8.3120 3.5100 8.3300 3.9150 ;
      LAYER V3  ;
        RECT 8.3120 3.5720 8.3300 3.5960 ;
    END
  END wd[3]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.7480 8.5970 4.7720 ;
      LAYER M3  ;
        RECT 8.5370 4.6975 8.5550 4.9370 ;
      LAYER V3  ;
        RECT 8.5370 4.7480 8.5550 4.7720 ;
    END
  END dataout[4]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.6520 8.6650 4.6760 ;
      LAYER M3  ;
        RECT 8.3120 4.5900 8.3300 4.9950 ;
      LAYER V3  ;
        RECT 8.3120 4.6520 8.3300 4.6760 ;
    END
  END wd[4]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.8280 8.5970 5.8520 ;
      LAYER M3  ;
        RECT 8.5370 5.7775 8.5550 6.0170 ;
      LAYER V3  ;
        RECT 8.5370 5.8280 8.5550 5.8520 ;
    END
  END dataout[5]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.7320 8.6650 5.7560 ;
      LAYER M3  ;
        RECT 8.3120 5.6700 8.3300 6.0750 ;
      LAYER V3  ;
        RECT 8.3120 5.7320 8.3300 5.7560 ;
    END
  END wd[5]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.9080 8.5970 6.9320 ;
      LAYER M3  ;
        RECT 8.5370 6.8575 8.5550 7.0970 ;
      LAYER V3  ;
        RECT 8.5370 6.9080 8.5550 6.9320 ;
    END
  END dataout[6]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.8120 8.6650 6.8360 ;
      LAYER M3  ;
        RECT 8.3120 6.7500 8.3300 7.1550 ;
      LAYER V3  ;
        RECT 8.3120 6.8120 8.3300 6.8360 ;
    END
  END wd[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.9880 8.5970 8.0120 ;
      LAYER M3  ;
        RECT 8.5370 7.9375 8.5550 8.1770 ;
      LAYER V3  ;
        RECT 8.5370 7.9880 8.5550 8.0120 ;
    END
  END dataout[7]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.8920 8.6650 7.9160 ;
      LAYER M3  ;
        RECT 8.3120 7.8300 8.3300 8.2350 ;
      LAYER V3  ;
        RECT 8.3120 7.8920 8.3300 7.9160 ;
    END
  END wd[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 9.0680 8.5970 9.0920 ;
      LAYER M3  ;
        RECT 8.5370 9.0175 8.5550 9.2570 ;
      LAYER V3  ;
        RECT 8.5370 9.0680 8.5550 9.0920 ;
    END
  END dataout[8]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 8.9720 8.6650 8.9960 ;
      LAYER M3  ;
        RECT 8.3120 8.9100 8.3300 9.3150 ;
      LAYER V3  ;
        RECT 8.3120 8.9720 8.3300 8.9960 ;
    END
  END wd[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 10.1480 8.5970 10.1720 ;
      LAYER M3  ;
        RECT 8.5370 10.0975 8.5550 10.3370 ;
      LAYER V3  ;
        RECT 8.5370 10.1480 8.5550 10.1720 ;
    END
  END dataout[9]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 10.0520 8.6650 10.0760 ;
      LAYER M3  ;
        RECT 8.3120 9.9900 8.3300 10.3950 ;
      LAYER V3  ;
        RECT 8.3120 10.0520 8.3300 10.0760 ;
    END
  END wd[9]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.3550 8.5970 19.3790 ;
      LAYER M3  ;
        RECT 8.5370 19.3045 8.5550 19.5440 ;
      LAYER V3  ;
        RECT 8.5370 19.3550 8.5550 19.3790 ;
    END
  END dataout[10]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.2590 8.6650 19.2830 ;
      LAYER M3  ;
        RECT 8.3120 19.1970 8.3300 19.6020 ;
      LAYER V3  ;
        RECT 8.3120 19.2590 8.3300 19.2830 ;
    END
  END wd[10]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.4350 8.5970 20.4590 ;
      LAYER M3  ;
        RECT 8.5370 20.3845 8.5550 20.6240 ;
      LAYER V3  ;
        RECT 8.5370 20.4350 8.5550 20.4590 ;
    END
  END dataout[11]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.3390 8.6650 20.3630 ;
      LAYER M3  ;
        RECT 8.3120 20.2770 8.3300 20.6820 ;
      LAYER V3  ;
        RECT 8.3120 20.3390 8.3300 20.3630 ;
    END
  END wd[11]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 21.5150 8.5970 21.5390 ;
      LAYER M3  ;
        RECT 8.5370 21.4645 8.5550 21.7040 ;
      LAYER V3  ;
        RECT 8.5370 21.5150 8.5550 21.5390 ;
    END
  END dataout[12]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 21.4190 8.6650 21.4430 ;
      LAYER M3  ;
        RECT 8.3120 21.3570 8.3300 21.7620 ;
      LAYER V3  ;
        RECT 8.3120 21.4190 8.3300 21.4430 ;
    END
  END wd[12]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 22.5950 8.5970 22.6190 ;
      LAYER M3  ;
        RECT 8.5370 22.5445 8.5550 22.7840 ;
      LAYER V3  ;
        RECT 8.5370 22.5950 8.5550 22.6190 ;
    END
  END dataout[13]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 22.4990 8.6650 22.5230 ;
      LAYER M3  ;
        RECT 8.3120 22.4370 8.3300 22.8420 ;
      LAYER V3  ;
        RECT 8.3120 22.4990 8.3300 22.5230 ;
    END
  END wd[13]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.6750 8.5970 23.6990 ;
      LAYER M3  ;
        RECT 8.5370 23.6245 8.5550 23.8640 ;
      LAYER V3  ;
        RECT 8.5370 23.6750 8.5550 23.6990 ;
    END
  END dataout[14]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.5790 8.6650 23.6030 ;
      LAYER M3  ;
        RECT 8.3120 23.5170 8.3300 23.9220 ;
      LAYER V3  ;
        RECT 8.3120 23.5790 8.3300 23.6030 ;
    END
  END wd[14]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.7550 8.5970 24.7790 ;
      LAYER M3  ;
        RECT 8.5370 24.7045 8.5550 24.9440 ;
      LAYER V3  ;
        RECT 8.5370 24.7550 8.5550 24.7790 ;
    END
  END dataout[15]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.6590 8.6650 24.6830 ;
      LAYER M3  ;
        RECT 8.3120 24.5970 8.3300 25.0020 ;
      LAYER V3  ;
        RECT 8.3120 24.6590 8.3300 24.6830 ;
    END
  END wd[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.8350 8.5970 25.8590 ;
      LAYER M3  ;
        RECT 8.5370 25.7845 8.5550 26.0240 ;
      LAYER V3  ;
        RECT 8.5370 25.8350 8.5550 25.8590 ;
    END
  END dataout[16]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.7390 8.6650 25.7630 ;
      LAYER M3  ;
        RECT 8.3120 25.6770 8.3300 26.0820 ;
      LAYER V3  ;
        RECT 8.3120 25.7390 8.3300 25.7630 ;
    END
  END wd[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 26.9150 8.5970 26.9390 ;
      LAYER M3  ;
        RECT 8.5370 26.8645 8.5550 27.1040 ;
      LAYER V3  ;
        RECT 8.5370 26.9150 8.5550 26.9390 ;
    END
  END dataout[17]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 26.8190 8.6650 26.8430 ;
      LAYER M3  ;
        RECT 8.3120 26.7570 8.3300 27.1620 ;
      LAYER V3  ;
        RECT 8.3120 26.8190 8.3300 26.8430 ;
    END
  END wd[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 27.9950 8.5970 28.0190 ;
      LAYER M3  ;
        RECT 8.5370 27.9445 8.5550 28.1840 ;
      LAYER V3  ;
        RECT 8.5370 27.9950 8.5550 28.0190 ;
    END
  END dataout[18]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 27.8990 8.6650 27.9230 ;
      LAYER M3  ;
        RECT 8.3120 27.8370 8.3300 28.2420 ;
      LAYER V3  ;
        RECT 8.3120 27.8990 8.3300 27.9230 ;
    END
  END wd[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 29.0750 8.5970 29.0990 ;
      LAYER M3  ;
        RECT 8.5370 29.0245 8.5550 29.2640 ;
      LAYER V3  ;
        RECT 8.5370 29.0750 8.5550 29.0990 ;
    END
  END dataout[19]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 28.9790 8.6650 29.0030 ;
      LAYER M3  ;
        RECT 8.3120 28.9170 8.3300 29.3220 ;
      LAYER V3  ;
        RECT 8.3120 28.9790 8.3300 29.0030 ;
    END
  END wd[19]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0000 11.0370 16.5240 19.6905 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
        RECT 0.0050 27.8235 16.5290 28.9170 ;
        RECT 0.0050 28.9035 16.5290 29.9970 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0000 11.0370 16.5240 19.6905 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
        RECT 0.0050 27.8235 16.5290 28.9170 ;
        RECT 0.0050 28.9035 16.5290 29.9970 ;
  LAYER V1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0000 11.0370 16.5240 19.6905 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
        RECT 0.0050 27.8235 16.5290 28.9170 ;
        RECT 0.0050 28.9035 16.5290 29.9970 ;
  LAYER V2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0000 11.0370 16.5240 19.6905 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
        RECT 0.0050 27.8235 16.5290 28.9170 ;
        RECT 0.0050 28.9035 16.5290 29.9970 ;
  LAYER M3  ;
      RECT 8.6990 0.3450 8.7170 1.2805 ;
      RECT 8.6630 0.3450 8.6810 1.2805 ;
      RECT 8.6270 0.9220 8.6450 1.2445 ;
      RECT 8.5100 1.1190 8.5280 1.2285 ;
      RECT 8.5010 0.3775 8.5190 0.6170 ;
      RECT 8.4650 0.9585 8.4830 1.1120 ;
      RECT 8.3840 0.9840 8.4020 1.2420 ;
      RECT 7.8440 0.3450 7.8620 1.2805 ;
      RECT 7.8080 0.3450 7.8260 1.2805 ;
      RECT 7.7720 0.5260 7.7900 1.0940 ;
      RECT 8.6990 1.4250 8.7170 2.3605 ;
      RECT 8.6630 1.4250 8.6810 2.3605 ;
      RECT 8.6270 2.0020 8.6450 2.3245 ;
      RECT 8.5100 2.1990 8.5280 2.3085 ;
      RECT 8.5010 1.4575 8.5190 1.6970 ;
      RECT 8.4650 2.0385 8.4830 2.1920 ;
      RECT 8.3840 2.0640 8.4020 2.3220 ;
      RECT 7.8440 1.4250 7.8620 2.3605 ;
      RECT 7.8080 1.4250 7.8260 2.3605 ;
      RECT 7.7720 1.6060 7.7900 2.1740 ;
      RECT 8.6990 2.5050 8.7170 3.4405 ;
      RECT 8.6630 2.5050 8.6810 3.4405 ;
      RECT 8.6270 3.0820 8.6450 3.4045 ;
      RECT 8.5100 3.2790 8.5280 3.3885 ;
      RECT 8.5010 2.5375 8.5190 2.7770 ;
      RECT 8.4650 3.1185 8.4830 3.2720 ;
      RECT 8.3840 3.1440 8.4020 3.4020 ;
      RECT 7.8440 2.5050 7.8620 3.4405 ;
      RECT 7.8080 2.5050 7.8260 3.4405 ;
      RECT 7.7720 2.6860 7.7900 3.2540 ;
      RECT 8.6990 3.5850 8.7170 4.5205 ;
      RECT 8.6630 3.5850 8.6810 4.5205 ;
      RECT 8.6270 4.1620 8.6450 4.4845 ;
      RECT 8.5100 4.3590 8.5280 4.4685 ;
      RECT 8.5010 3.6175 8.5190 3.8570 ;
      RECT 8.4650 4.1985 8.4830 4.3520 ;
      RECT 8.3840 4.2240 8.4020 4.4820 ;
      RECT 7.8440 3.5850 7.8620 4.5205 ;
      RECT 7.8080 3.5850 7.8260 4.5205 ;
      RECT 7.7720 3.7660 7.7900 4.3340 ;
      RECT 8.6990 4.6650 8.7170 5.6005 ;
      RECT 8.6630 4.6650 8.6810 5.6005 ;
      RECT 8.6270 5.2420 8.6450 5.5645 ;
      RECT 8.5100 5.4390 8.5280 5.5485 ;
      RECT 8.5010 4.6975 8.5190 4.9370 ;
      RECT 8.4650 5.2785 8.4830 5.4320 ;
      RECT 8.3840 5.3040 8.4020 5.5620 ;
      RECT 7.8440 4.6650 7.8620 5.6005 ;
      RECT 7.8080 4.6650 7.8260 5.6005 ;
      RECT 7.7720 4.8460 7.7900 5.4140 ;
      RECT 8.6990 5.7450 8.7170 6.6805 ;
      RECT 8.6630 5.7450 8.6810 6.6805 ;
      RECT 8.6270 6.3220 8.6450 6.6445 ;
      RECT 8.5100 6.5190 8.5280 6.6285 ;
      RECT 8.5010 5.7775 8.5190 6.0170 ;
      RECT 8.4650 6.3585 8.4830 6.5120 ;
      RECT 8.3840 6.3840 8.4020 6.6420 ;
      RECT 7.8440 5.7450 7.8620 6.6805 ;
      RECT 7.8080 5.7450 7.8260 6.6805 ;
      RECT 7.7720 5.9260 7.7900 6.4940 ;
      RECT 8.6990 6.8250 8.7170 7.7605 ;
      RECT 8.6630 6.8250 8.6810 7.7605 ;
      RECT 8.6270 7.4020 8.6450 7.7245 ;
      RECT 8.5100 7.5990 8.5280 7.7085 ;
      RECT 8.5010 6.8575 8.5190 7.0970 ;
      RECT 8.4650 7.4385 8.4830 7.5920 ;
      RECT 8.3840 7.4640 8.4020 7.7220 ;
      RECT 7.8440 6.8250 7.8620 7.7605 ;
      RECT 7.8080 6.8250 7.8260 7.7605 ;
      RECT 7.7720 7.0060 7.7900 7.5740 ;
      RECT 8.6990 7.9050 8.7170 8.8405 ;
      RECT 8.6630 7.9050 8.6810 8.8405 ;
      RECT 8.6270 8.4820 8.6450 8.8045 ;
      RECT 8.5100 8.6790 8.5280 8.7885 ;
      RECT 8.5010 7.9375 8.5190 8.1770 ;
      RECT 8.4650 8.5185 8.4830 8.6720 ;
      RECT 8.3840 8.5440 8.4020 8.8020 ;
      RECT 7.8440 7.9050 7.8620 8.8405 ;
      RECT 7.8080 7.9050 7.8260 8.8405 ;
      RECT 7.7720 8.0860 7.7900 8.6540 ;
      RECT 8.6990 8.9850 8.7170 9.9205 ;
      RECT 8.6630 8.9850 8.6810 9.9205 ;
      RECT 8.6270 9.5620 8.6450 9.8845 ;
      RECT 8.5100 9.7590 8.5280 9.8685 ;
      RECT 8.5010 9.0175 8.5190 9.2570 ;
      RECT 8.4650 9.5985 8.4830 9.7520 ;
      RECT 8.3840 9.6240 8.4020 9.8820 ;
      RECT 7.8440 8.9850 7.8620 9.9205 ;
      RECT 7.8080 8.9850 7.8260 9.9205 ;
      RECT 7.7720 9.1660 7.7900 9.7340 ;
      RECT 8.6990 10.0650 8.7170 11.0005 ;
      RECT 8.6630 10.0650 8.6810 11.0005 ;
      RECT 8.6270 10.6420 8.6450 10.9645 ;
      RECT 8.5100 10.8390 8.5280 10.9485 ;
      RECT 8.5010 10.0975 8.5190 10.3370 ;
      RECT 8.4650 10.6785 8.4830 10.8320 ;
      RECT 8.3840 10.7040 8.4020 10.9620 ;
      RECT 7.8440 10.0650 7.8620 11.0005 ;
      RECT 7.8080 10.0650 7.8260 11.0005 ;
      RECT 7.7720 10.2460 7.7900 10.8140 ;
      RECT 16.3170 14.8300 16.3350 19.1840 ;
      RECT 16.2810 13.5150 16.2990 13.5840 ;
      RECT 16.2810 15.1350 16.2990 15.2180 ;
      RECT 16.2450 11.0105 16.2630 19.2175 ;
      RECT 16.2090 14.8625 16.2270 15.5525 ;
      RECT 16.2090 15.6035 16.2270 16.5900 ;
      RECT 16.2090 16.6300 16.2270 17.2470 ;
      RECT 16.1730 14.7990 16.1910 15.5038 ;
      RECT 16.1730 16.2570 16.1910 17.4270 ;
      RECT 16.1370 11.0105 16.1550 14.6070 ;
      RECT 16.0290 11.0105 16.0470 14.6070 ;
      RECT 15.9210 11.0105 15.9390 14.6070 ;
      RECT 15.8130 11.0105 15.8310 14.6070 ;
      RECT 15.7050 11.0105 15.7230 14.6070 ;
      RECT 15.5970 11.0105 15.6150 14.6070 ;
      RECT 15.4890 11.0105 15.5070 14.6070 ;
      RECT 15.3810 11.0105 15.3990 14.6070 ;
      RECT 15.2730 11.0105 15.2910 14.6070 ;
      RECT 15.1650 11.0105 15.1830 14.6070 ;
      RECT 15.0570 11.0105 15.0750 14.6070 ;
      RECT 14.9490 11.0105 14.9670 14.6070 ;
      RECT 14.8410 11.0105 14.8590 14.6070 ;
      RECT 14.7330 11.0105 14.7510 14.6070 ;
      RECT 14.6250 11.0105 14.6430 14.6070 ;
      RECT 14.5170 11.0105 14.5350 14.6070 ;
      RECT 14.4090 11.0105 14.4270 14.6070 ;
      RECT 14.3010 11.0105 14.3190 14.6070 ;
      RECT 14.1930 11.0105 14.2110 14.6070 ;
      RECT 14.0850 11.0105 14.1030 14.6070 ;
      RECT 13.9770 11.0105 13.9950 14.6070 ;
      RECT 13.8690 11.0105 13.8870 14.6070 ;
      RECT 13.7610 11.0105 13.7790 14.6070 ;
      RECT 13.6530 11.0105 13.6710 14.6070 ;
      RECT 13.5450 11.0105 13.5630 14.6070 ;
      RECT 13.4370 11.0105 13.4550 14.6070 ;
      RECT 13.3290 11.0105 13.3470 14.6070 ;
      RECT 13.2210 11.0105 13.2390 14.6070 ;
      RECT 13.1130 11.0105 13.1310 14.6070 ;
      RECT 13.0050 11.0105 13.0230 14.6070 ;
      RECT 12.8970 11.0105 12.9150 14.6070 ;
      RECT 12.7890 11.0105 12.8070 14.6070 ;
      RECT 12.6810 11.0105 12.6990 14.6070 ;
      RECT 12.5730 11.0105 12.5910 14.6070 ;
      RECT 12.4650 11.0105 12.4830 14.6070 ;
      RECT 12.3570 11.0105 12.3750 14.6070 ;
      RECT 12.2490 11.0105 12.2670 14.6070 ;
      RECT 12.1410 11.0105 12.1590 14.6070 ;
      RECT 12.0330 11.0105 12.0510 14.6070 ;
      RECT 11.9250 11.0105 11.9430 14.6070 ;
      RECT 11.8170 11.0105 11.8350 14.6070 ;
      RECT 11.7090 11.0105 11.7270 14.6070 ;
      RECT 11.6010 11.0105 11.6190 14.6070 ;
      RECT 11.4930 11.0105 11.5110 14.6070 ;
      RECT 11.3850 11.0105 11.4030 14.6070 ;
      RECT 11.2770 11.0105 11.2950 14.6070 ;
      RECT 11.1690 11.0105 11.1870 14.6070 ;
      RECT 11.0610 11.0105 11.0790 14.6070 ;
      RECT 10.9530 11.0105 10.9710 14.6070 ;
      RECT 10.8450 11.0105 10.8630 14.6070 ;
      RECT 10.7370 11.0105 10.7550 14.6070 ;
      RECT 10.6290 11.0105 10.6470 14.6070 ;
      RECT 10.5210 11.0105 10.5390 14.6070 ;
      RECT 10.4130 11.0105 10.4310 14.6070 ;
      RECT 10.3050 11.0105 10.3230 14.6070 ;
      RECT 10.1970 11.0105 10.2150 14.6070 ;
      RECT 10.0890 11.0105 10.1070 14.6070 ;
      RECT 9.9810 11.0105 9.9990 14.6070 ;
      RECT 9.8730 11.0105 9.8910 14.6070 ;
      RECT 9.7650 11.0105 9.7830 14.6070 ;
      RECT 9.6570 11.0105 9.6750 14.6070 ;
      RECT 9.5490 11.0105 9.5670 14.6070 ;
      RECT 9.5130 14.8655 9.5310 15.5075 ;
      RECT 9.5130 16.1850 9.5310 16.7170 ;
      RECT 9.4950 11.6710 9.5130 12.3470 ;
      RECT 9.4950 13.0930 9.5130 13.3910 ;
      RECT 9.4950 14.2090 9.5130 14.4710 ;
      RECT 9.4770 14.7800 9.4950 15.5525 ;
      RECT 9.4770 15.6037 9.4950 16.0950 ;
      RECT 9.4770 16.1400 9.4950 16.5110 ;
      RECT 9.4770 16.5870 9.4950 17.2470 ;
      RECT 9.4410 11.0105 9.4590 19.2175 ;
      RECT 9.4050 15.3230 9.4230 15.7875 ;
      RECT 9.3870 11.7790 9.4050 12.4100 ;
      RECT 9.3870 12.8230 9.4050 13.0130 ;
      RECT 9.3870 13.7050 9.4050 13.7540 ;
      RECT 9.3870 14.4370 9.4050 14.4740 ;
      RECT 9.3690 14.8300 9.3870 19.1795 ;
      RECT 9.2790 11.4010 9.2970 12.2030 ;
      RECT 9.2790 12.7510 9.2970 13.3190 ;
      RECT 9.2430 12.8230 9.2610 13.1930 ;
      RECT 9.2070 12.1750 9.2250 12.3110 ;
      RECT 9.2070 13.1650 9.2250 13.3910 ;
      RECT 9.2070 14.4070 9.2250 14.4710 ;
      RECT 9.1710 12.2770 9.1890 12.3140 ;
      RECT 9.1710 13.9030 9.1890 13.9460 ;
      RECT 9.1710 14.4370 9.1890 14.4740 ;
      RECT 9.1350 12.5890 9.1530 13.0850 ;
      RECT 9.1350 13.1290 9.1530 13.3190 ;
      RECT 9.1350 14.0890 9.1530 14.3990 ;
      RECT 9.0990 12.4810 9.1170 13.7280 ;
      RECT 9.0990 16.3690 9.1170 17.0990 ;
      RECT 9.0990 17.4490 9.1170 18.1790 ;
      RECT 8.7750 12.2110 8.7930 12.5090 ;
      RECT 8.7750 13.3990 8.7930 13.4630 ;
      RECT 8.7750 13.6690 8.7930 14.1290 ;
      RECT 8.7750 14.8690 8.7930 14.9060 ;
      RECT 8.7750 16.9090 8.7930 17.2070 ;
      RECT 8.7390 12.2830 8.7570 12.7880 ;
      RECT 8.7390 13.0570 8.7570 13.8590 ;
      RECT 8.7390 14.9020 8.7570 15.1730 ;
      RECT 8.7390 15.2530 8.7570 15.4790 ;
      RECT 8.7030 12.2110 8.7210 12.8870 ;
      RECT 8.7030 12.9850 8.7210 13.3190 ;
      RECT 8.7030 13.5250 8.7210 13.6610 ;
      RECT 8.7030 14.2090 8.7210 15.0110 ;
      RECT 8.7030 15.4450 8.7210 15.4820 ;
      RECT 8.7030 17.6110 8.7210 17.9450 ;
      RECT 8.6670 12.4450 8.6850 12.5810 ;
      RECT 8.6670 14.3350 8.6850 15.3170 ;
      RECT 8.6670 15.7570 8.6850 16.0550 ;
      RECT 8.6670 17.4490 8.6850 17.7110 ;
      RECT 8.6310 11.5090 8.6490 11.6630 ;
      RECT 8.6310 12.3190 8.6490 14.1050 ;
      RECT 8.6310 15.1450 8.6490 17.4770 ;
      RECT 8.6310 17.6830 8.6490 18.7910 ;
      RECT 8.3430 11.7790 8.3610 12.0410 ;
      RECT 8.3430 12.1750 8.3610 12.2390 ;
      RECT 8.3430 12.3190 8.3610 12.5450 ;
      RECT 8.3430 12.5890 8.3610 12.7790 ;
      RECT 8.3430 12.8590 8.3610 15.4790 ;
      RECT 8.3430 15.5230 8.3610 16.8290 ;
      RECT 8.3430 17.9170 8.3610 18.1790 ;
      RECT 8.3070 12.7780 8.3250 13.0490 ;
      RECT 8.3070 13.1290 8.3250 13.9670 ;
      RECT 8.3070 14.1370 8.3250 14.9750 ;
      RECT 8.3070 15.0190 8.3250 16.2890 ;
      RECT 8.3070 16.4950 8.3250 16.6670 ;
      RECT 8.3070 17.3770 8.3250 18.4490 ;
      RECT 8.2710 12.8590 8.2890 13.1300 ;
      RECT 8.2710 13.2850 8.2890 13.3220 ;
      RECT 8.2710 14.0650 8.2890 15.0470 ;
      RECT 8.2710 15.2890 8.2890 15.7490 ;
      RECT 8.2710 16.0990 8.2890 16.8380 ;
      RECT 8.2350 11.9770 8.2530 13.0490 ;
      RECT 8.2350 14.6410 8.2530 14.8580 ;
      RECT 8.2350 16.0270 8.2530 16.3250 ;
      RECT 8.1990 12.6250 8.2170 13.0850 ;
      RECT 8.1990 14.2090 8.2170 14.3990 ;
      RECT 8.1990 14.4400 8.2170 14.4770 ;
      RECT 8.1990 14.7130 8.2170 15.0470 ;
      RECT 8.1990 15.1810 8.2170 16.5230 ;
      RECT 8.1990 16.6300 8.2170 17.7470 ;
      RECT 8.1630 12.0490 8.1810 12.2390 ;
      RECT 8.1630 12.4450 8.1810 12.5810 ;
      RECT 8.1630 12.8590 8.1810 16.0190 ;
      RECT 8.1630 16.0990 8.1810 16.5590 ;
      RECT 8.1630 17.1790 8.1810 17.6390 ;
      RECT 8.1630 18.4930 8.1810 18.7190 ;
      RECT 8.1270 11.0370 8.1450 11.1910 ;
      RECT 8.1270 19.0320 8.1450 19.1980 ;
      RECT 8.0910 11.0370 8.1090 11.0870 ;
      RECT 8.0190 11.0370 8.0370 11.1085 ;
      RECT 8.0190 19.1015 8.0370 19.2175 ;
      RECT 7.8750 12.5530 7.8930 12.7430 ;
      RECT 7.8750 13.2910 7.8930 13.6610 ;
      RECT 7.8750 15.2530 7.8930 15.4790 ;
      RECT 7.8750 15.7930 7.8930 16.9370 ;
      RECT 7.8750 17.7190 7.8930 18.1790 ;
      RECT 7.8750 18.7570 7.8930 18.7940 ;
      RECT 7.8390 11.5090 7.8570 12.0050 ;
      RECT 7.8390 15.5890 7.8570 15.6260 ;
      RECT 7.8390 16.6660 7.8570 17.4770 ;
      RECT 7.8030 11.9770 7.8210 12.2390 ;
      RECT 7.8030 12.5170 7.8210 12.8510 ;
      RECT 7.8030 13.0570 7.8210 13.1570 ;
      RECT 7.8030 13.9390 7.8210 16.7030 ;
      RECT 7.8030 16.8370 7.8210 17.0630 ;
      RECT 7.7670 11.6350 7.7850 12.7790 ;
      RECT 7.7670 16.3690 7.7850 16.5590 ;
      RECT 7.7670 17.1730 7.7850 17.2100 ;
      RECT 7.7670 17.4490 7.7850 18.2510 ;
      RECT 7.7310 12.5890 7.7490 13.5890 ;
      RECT 7.7310 17.0290 7.7490 17.0660 ;
      RECT 7.3710 12.1750 7.3890 12.5810 ;
      RECT 7.2990 12.2110 7.3170 12.8150 ;
      RECT 7.2630 12.0490 7.2810 12.1130 ;
      RECT 7.2270 11.0900 7.2450 11.1410 ;
      RECT 7.2270 14.2090 7.2450 14.3990 ;
      RECT 7.2090 14.8300 7.2270 19.1785 ;
      RECT 7.1370 14.8300 7.1550 19.1795 ;
      RECT 7.1190 11.5090 7.1370 11.6990 ;
      RECT 7.1190 12.2830 7.1370 14.5430 ;
      RECT 7.1010 15.3230 7.1190 15.7875 ;
      RECT 7.0650 11.0105 7.0830 19.2175 ;
      RECT 7.0290 14.7800 7.0470 15.5525 ;
      RECT 7.0290 15.6037 7.0470 16.0950 ;
      RECT 7.0290 16.1400 7.0470 16.5110 ;
      RECT 7.0290 16.5870 7.0470 17.2470 ;
      RECT 7.0110 11.5090 7.0290 12.0050 ;
      RECT 7.0110 12.7870 7.0290 13.3550 ;
      RECT 7.0110 13.6690 7.0290 14.3990 ;
      RECT 6.9930 14.8655 7.0110 15.5075 ;
      RECT 6.9930 16.1850 7.0110 16.7170 ;
      RECT 6.9570 11.0105 6.9750 14.6070 ;
      RECT 6.8490 11.0105 6.8670 14.6070 ;
      RECT 6.7410 11.0105 6.7590 14.6070 ;
      RECT 6.6330 11.0105 6.6510 14.6070 ;
      RECT 6.5250 11.0105 6.5430 14.6070 ;
      RECT 6.4170 11.0105 6.4350 14.6070 ;
      RECT 6.3090 11.0105 6.3270 14.6070 ;
      RECT 6.2010 11.0105 6.2190 14.6070 ;
      RECT 6.0930 11.0105 6.1110 14.6070 ;
      RECT 5.9850 11.0105 6.0030 14.6070 ;
      RECT 5.8770 11.0105 5.8950 14.6070 ;
      RECT 5.7690 11.0105 5.7870 14.6070 ;
      RECT 5.6610 11.0105 5.6790 14.6070 ;
      RECT 5.5530 11.0105 5.5710 14.6070 ;
      RECT 5.4450 11.0105 5.4630 14.6070 ;
      RECT 5.3370 11.0105 5.3550 14.6070 ;
      RECT 5.2290 11.0105 5.2470 14.6070 ;
      RECT 5.1210 11.0105 5.1390 14.6070 ;
      RECT 5.0130 11.0105 5.0310 14.6070 ;
      RECT 4.9050 11.0105 4.9230 14.6070 ;
      RECT 4.7970 11.0105 4.8150 14.6070 ;
      RECT 4.6890 11.0105 4.7070 14.6070 ;
      RECT 4.5810 11.0105 4.5990 14.6070 ;
      RECT 4.4730 11.0105 4.4910 14.6070 ;
      RECT 4.3650 11.0105 4.3830 14.6070 ;
      RECT 4.2570 11.0105 4.2750 14.6070 ;
      RECT 4.1490 11.0105 4.1670 14.6070 ;
      RECT 4.0410 11.0105 4.0590 14.6070 ;
      RECT 3.9330 11.0105 3.9510 14.6070 ;
      RECT 3.8250 11.0105 3.8430 14.6070 ;
      RECT 3.7170 11.0105 3.7350 14.6070 ;
      RECT 3.6090 11.0105 3.6270 14.6070 ;
      RECT 3.5010 11.0105 3.5190 14.6070 ;
      RECT 3.3930 11.0105 3.4110 14.6070 ;
      RECT 3.2850 11.0105 3.3030 14.6070 ;
      RECT 3.1770 11.0105 3.1950 14.6070 ;
      RECT 3.0690 11.0105 3.0870 14.6070 ;
      RECT 2.9610 11.0105 2.9790 14.6070 ;
      RECT 2.8530 11.0105 2.8710 14.6070 ;
      RECT 2.7450 11.0105 2.7630 14.6070 ;
      RECT 2.6370 11.0105 2.6550 14.6070 ;
      RECT 2.5290 11.0105 2.5470 14.6070 ;
      RECT 2.4210 11.0105 2.4390 14.6070 ;
      RECT 2.3130 11.0105 2.3310 14.6070 ;
      RECT 2.2050 11.0105 2.2230 14.6070 ;
      RECT 2.0970 11.0105 2.1150 14.6070 ;
      RECT 1.9890 11.0105 2.0070 14.6070 ;
      RECT 1.8810 11.0105 1.8990 14.6070 ;
      RECT 1.7730 11.0105 1.7910 14.6070 ;
      RECT 1.6650 11.0105 1.6830 14.6070 ;
      RECT 1.5570 11.0105 1.5750 14.6070 ;
      RECT 1.4490 11.0105 1.4670 14.6070 ;
      RECT 1.3410 11.0105 1.3590 14.6070 ;
      RECT 1.2330 11.0105 1.2510 14.6070 ;
      RECT 1.1250 11.0105 1.1430 14.6070 ;
      RECT 1.0170 11.0105 1.0350 14.6070 ;
      RECT 0.9090 11.0105 0.9270 14.6070 ;
      RECT 0.8010 11.0105 0.8190 14.6070 ;
      RECT 0.6930 11.0105 0.7110 14.6070 ;
      RECT 0.5850 11.0105 0.6030 14.6070 ;
      RECT 0.4770 11.0105 0.4950 14.6070 ;
      RECT 0.3690 11.0105 0.3870 14.6070 ;
      RECT 0.3330 14.7990 0.3510 15.5038 ;
      RECT 0.3330 16.2570 0.3510 17.4270 ;
      RECT 0.2970 14.8625 0.3150 15.5525 ;
      RECT 0.2970 15.6035 0.3150 16.5900 ;
      RECT 0.2970 16.6300 0.3150 17.2470 ;
      RECT 0.2610 11.0105 0.2790 19.2175 ;
      RECT 0.2250 13.5150 0.2430 13.5840 ;
      RECT 0.2250 15.1350 0.2430 15.2180 ;
      RECT 0.1890 14.8300 0.2070 19.1840 ;
        RECT 8.6990 19.2720 8.7170 20.2075 ;
        RECT 8.6630 19.2720 8.6810 20.2075 ;
        RECT 8.6270 19.8490 8.6450 20.1715 ;
        RECT 8.5100 20.0460 8.5280 20.1555 ;
        RECT 8.5010 19.3045 8.5190 19.5440 ;
        RECT 8.4650 19.8855 8.4830 20.0390 ;
        RECT 8.3840 19.9110 8.4020 20.1690 ;
        RECT 7.8440 19.2720 7.8620 20.2075 ;
        RECT 7.8080 19.2720 7.8260 20.2075 ;
        RECT 7.7720 19.4530 7.7900 20.0210 ;
        RECT 8.6990 20.3520 8.7170 21.2875 ;
        RECT 8.6630 20.3520 8.6810 21.2875 ;
        RECT 8.6270 20.9290 8.6450 21.2515 ;
        RECT 8.5100 21.1260 8.5280 21.2355 ;
        RECT 8.5010 20.3845 8.5190 20.6240 ;
        RECT 8.4650 20.9655 8.4830 21.1190 ;
        RECT 8.3840 20.9910 8.4020 21.2490 ;
        RECT 7.8440 20.3520 7.8620 21.2875 ;
        RECT 7.8080 20.3520 7.8260 21.2875 ;
        RECT 7.7720 20.5330 7.7900 21.1010 ;
        RECT 8.6990 21.4320 8.7170 22.3675 ;
        RECT 8.6630 21.4320 8.6810 22.3675 ;
        RECT 8.6270 22.0090 8.6450 22.3315 ;
        RECT 8.5100 22.2060 8.5280 22.3155 ;
        RECT 8.5010 21.4645 8.5190 21.7040 ;
        RECT 8.4650 22.0455 8.4830 22.1990 ;
        RECT 8.3840 22.0710 8.4020 22.3290 ;
        RECT 7.8440 21.4320 7.8620 22.3675 ;
        RECT 7.8080 21.4320 7.8260 22.3675 ;
        RECT 7.7720 21.6130 7.7900 22.1810 ;
        RECT 8.6990 22.5120 8.7170 23.4475 ;
        RECT 8.6630 22.5120 8.6810 23.4475 ;
        RECT 8.6270 23.0890 8.6450 23.4115 ;
        RECT 8.5100 23.2860 8.5280 23.3955 ;
        RECT 8.5010 22.5445 8.5190 22.7840 ;
        RECT 8.4650 23.1255 8.4830 23.2790 ;
        RECT 8.3840 23.1510 8.4020 23.4090 ;
        RECT 7.8440 22.5120 7.8620 23.4475 ;
        RECT 7.8080 22.5120 7.8260 23.4475 ;
        RECT 7.7720 22.6930 7.7900 23.2610 ;
        RECT 8.6990 23.5920 8.7170 24.5275 ;
        RECT 8.6630 23.5920 8.6810 24.5275 ;
        RECT 8.6270 24.1690 8.6450 24.4915 ;
        RECT 8.5100 24.3660 8.5280 24.4755 ;
        RECT 8.5010 23.6245 8.5190 23.8640 ;
        RECT 8.4650 24.2055 8.4830 24.3590 ;
        RECT 8.3840 24.2310 8.4020 24.4890 ;
        RECT 7.8440 23.5920 7.8620 24.5275 ;
        RECT 7.8080 23.5920 7.8260 24.5275 ;
        RECT 7.7720 23.7730 7.7900 24.3410 ;
        RECT 8.6990 24.6720 8.7170 25.6075 ;
        RECT 8.6630 24.6720 8.6810 25.6075 ;
        RECT 8.6270 25.2490 8.6450 25.5715 ;
        RECT 8.5100 25.4460 8.5280 25.5555 ;
        RECT 8.5010 24.7045 8.5190 24.9440 ;
        RECT 8.4650 25.2855 8.4830 25.4390 ;
        RECT 8.3840 25.3110 8.4020 25.5690 ;
        RECT 7.8440 24.6720 7.8620 25.6075 ;
        RECT 7.8080 24.6720 7.8260 25.6075 ;
        RECT 7.7720 24.8530 7.7900 25.4210 ;
        RECT 8.6990 25.7520 8.7170 26.6875 ;
        RECT 8.6630 25.7520 8.6810 26.6875 ;
        RECT 8.6270 26.3290 8.6450 26.6515 ;
        RECT 8.5100 26.5260 8.5280 26.6355 ;
        RECT 8.5010 25.7845 8.5190 26.0240 ;
        RECT 8.4650 26.3655 8.4830 26.5190 ;
        RECT 8.3840 26.3910 8.4020 26.6490 ;
        RECT 7.8440 25.7520 7.8620 26.6875 ;
        RECT 7.8080 25.7520 7.8260 26.6875 ;
        RECT 7.7720 25.9330 7.7900 26.5010 ;
        RECT 8.6990 26.8320 8.7170 27.7675 ;
        RECT 8.6630 26.8320 8.6810 27.7675 ;
        RECT 8.6270 27.4090 8.6450 27.7315 ;
        RECT 8.5100 27.6060 8.5280 27.7155 ;
        RECT 8.5010 26.8645 8.5190 27.1040 ;
        RECT 8.4650 27.4455 8.4830 27.5990 ;
        RECT 8.3840 27.4710 8.4020 27.7290 ;
        RECT 7.8440 26.8320 7.8620 27.7675 ;
        RECT 7.8080 26.8320 7.8260 27.7675 ;
        RECT 7.7720 27.0130 7.7900 27.5810 ;
        RECT 8.6990 27.9120 8.7170 28.8475 ;
        RECT 8.6630 27.9120 8.6810 28.8475 ;
        RECT 8.6270 28.4890 8.6450 28.8115 ;
        RECT 8.5100 28.6860 8.5280 28.7955 ;
        RECT 8.5010 27.9445 8.5190 28.1840 ;
        RECT 8.4650 28.5255 8.4830 28.6790 ;
        RECT 8.3840 28.5510 8.4020 28.8090 ;
        RECT 7.8440 27.9120 7.8620 28.8475 ;
        RECT 7.8080 27.9120 7.8260 28.8475 ;
        RECT 7.7720 28.0930 7.7900 28.6610 ;
        RECT 8.6990 28.9920 8.7170 29.9275 ;
        RECT 8.6630 28.9920 8.6810 29.9275 ;
        RECT 8.6270 29.5690 8.6450 29.8915 ;
        RECT 8.5100 29.7660 8.5280 29.8755 ;
        RECT 8.5010 29.0245 8.5190 29.2640 ;
        RECT 8.4650 29.6055 8.4830 29.7590 ;
        RECT 8.3840 29.6310 8.4020 29.8890 ;
        RECT 7.8440 28.9920 7.8620 29.9275 ;
        RECT 7.8080 28.9920 7.8260 29.9275 ;
        RECT 7.7720 29.1730 7.7900 29.7410 ;
  LAYER M3 SPACING 0.018  ;
      RECT 8.6410 0.2565 8.7690 1.3500 ;
      RECT 8.6270 0.9220 8.7690 1.2445 ;
      RECT 8.4790 0.6490 8.5410 1.3500 ;
      RECT 8.4650 0.9585 8.5410 1.1120 ;
      RECT 8.4790 0.2565 8.5050 1.3500 ;
      RECT 8.4790 0.3775 8.5190 0.6170 ;
      RECT 8.4790 0.2565 8.5410 0.3455 ;
      RECT 8.1820 0.7070 8.3880 1.3500 ;
      RECT 8.3620 0.2565 8.3880 1.3500 ;
      RECT 8.1820 0.9840 8.4020 1.2420 ;
      RECT 8.1820 0.2565 8.2800 1.3500 ;
      RECT 7.7650 0.2565 7.8480 1.3500 ;
      RECT 7.7650 0.3450 7.8620 1.2805 ;
      RECT 16.4440 0.2565 16.5290 1.3500 ;
      RECT 16.3000 0.2565 16.3260 1.3500 ;
      RECT 16.1920 0.2565 16.2180 1.3500 ;
      RECT 16.0840 0.2565 16.1100 1.3500 ;
      RECT 15.9760 0.2565 16.0020 1.3500 ;
      RECT 15.8680 0.2565 15.8940 1.3500 ;
      RECT 15.7600 0.2565 15.7860 1.3500 ;
      RECT 15.6520 0.2565 15.6780 1.3500 ;
      RECT 15.5440 0.2565 15.5700 1.3500 ;
      RECT 15.4360 0.2565 15.4620 1.3500 ;
      RECT 15.3280 0.2565 15.3540 1.3500 ;
      RECT 15.2200 0.2565 15.2460 1.3500 ;
      RECT 15.1120 0.2565 15.1380 1.3500 ;
      RECT 15.0040 0.2565 15.0300 1.3500 ;
      RECT 14.8960 0.2565 14.9220 1.3500 ;
      RECT 14.7880 0.2565 14.8140 1.3500 ;
      RECT 14.6800 0.2565 14.7060 1.3500 ;
      RECT 14.5720 0.2565 14.5980 1.3500 ;
      RECT 14.4640 0.2565 14.4900 1.3500 ;
      RECT 14.3560 0.2565 14.3820 1.3500 ;
      RECT 14.2480 0.2565 14.2740 1.3500 ;
      RECT 14.1400 0.2565 14.1660 1.3500 ;
      RECT 14.0320 0.2565 14.0580 1.3500 ;
      RECT 13.9240 0.2565 13.9500 1.3500 ;
      RECT 13.8160 0.2565 13.8420 1.3500 ;
      RECT 13.7080 0.2565 13.7340 1.3500 ;
      RECT 13.6000 0.2565 13.6260 1.3500 ;
      RECT 13.4920 0.2565 13.5180 1.3500 ;
      RECT 13.3840 0.2565 13.4100 1.3500 ;
      RECT 13.2760 0.2565 13.3020 1.3500 ;
      RECT 13.1680 0.2565 13.1940 1.3500 ;
      RECT 13.0600 0.2565 13.0860 1.3500 ;
      RECT 12.9520 0.2565 12.9780 1.3500 ;
      RECT 12.8440 0.2565 12.8700 1.3500 ;
      RECT 12.7360 0.2565 12.7620 1.3500 ;
      RECT 12.6280 0.2565 12.6540 1.3500 ;
      RECT 12.5200 0.2565 12.5460 1.3500 ;
      RECT 12.4120 0.2565 12.4380 1.3500 ;
      RECT 12.3040 0.2565 12.3300 1.3500 ;
      RECT 12.1960 0.2565 12.2220 1.3500 ;
      RECT 12.0880 0.2565 12.1140 1.3500 ;
      RECT 11.9800 0.2565 12.0060 1.3500 ;
      RECT 11.8720 0.2565 11.8980 1.3500 ;
      RECT 11.7640 0.2565 11.7900 1.3500 ;
      RECT 11.6560 0.2565 11.6820 1.3500 ;
      RECT 11.5480 0.2565 11.5740 1.3500 ;
      RECT 11.4400 0.2565 11.4660 1.3500 ;
      RECT 11.3320 0.2565 11.3580 1.3500 ;
      RECT 11.2240 0.2565 11.2500 1.3500 ;
      RECT 11.1160 0.2565 11.1420 1.3500 ;
      RECT 11.0080 0.2565 11.0340 1.3500 ;
      RECT 10.9000 0.2565 10.9260 1.3500 ;
      RECT 10.7920 0.2565 10.8180 1.3500 ;
      RECT 10.6840 0.2565 10.7100 1.3500 ;
      RECT 10.5760 0.2565 10.6020 1.3500 ;
      RECT 10.4680 0.2565 10.4940 1.3500 ;
      RECT 10.3600 0.2565 10.3860 1.3500 ;
      RECT 10.2520 0.2565 10.2780 1.3500 ;
      RECT 10.1440 0.2565 10.1700 1.3500 ;
      RECT 10.0360 0.2565 10.0620 1.3500 ;
      RECT 9.9280 0.2565 9.9540 1.3500 ;
      RECT 9.8200 0.2565 9.8460 1.3500 ;
      RECT 9.7120 0.2565 9.7380 1.3500 ;
      RECT 9.6040 0.2565 9.6300 1.3500 ;
      RECT 9.4960 0.2565 9.5220 1.3500 ;
      RECT 9.3880 0.2565 9.4140 1.3500 ;
      RECT 9.1750 0.2565 9.2520 1.3500 ;
      RECT 7.2820 0.2565 7.3590 1.3500 ;
      RECT 7.1200 0.2565 7.1460 1.3500 ;
      RECT 7.0120 0.2565 7.0380 1.3500 ;
      RECT 6.9040 0.2565 6.9300 1.3500 ;
      RECT 6.7960 0.2565 6.8220 1.3500 ;
      RECT 6.6880 0.2565 6.7140 1.3500 ;
      RECT 6.5800 0.2565 6.6060 1.3500 ;
      RECT 6.4720 0.2565 6.4980 1.3500 ;
      RECT 6.3640 0.2565 6.3900 1.3500 ;
      RECT 6.2560 0.2565 6.2820 1.3500 ;
      RECT 6.1480 0.2565 6.1740 1.3500 ;
      RECT 6.0400 0.2565 6.0660 1.3500 ;
      RECT 5.9320 0.2565 5.9580 1.3500 ;
      RECT 5.8240 0.2565 5.8500 1.3500 ;
      RECT 5.7160 0.2565 5.7420 1.3500 ;
      RECT 5.6080 0.2565 5.6340 1.3500 ;
      RECT 5.5000 0.2565 5.5260 1.3500 ;
      RECT 5.3920 0.2565 5.4180 1.3500 ;
      RECT 5.2840 0.2565 5.3100 1.3500 ;
      RECT 5.1760 0.2565 5.2020 1.3500 ;
      RECT 5.0680 0.2565 5.0940 1.3500 ;
      RECT 4.9600 0.2565 4.9860 1.3500 ;
      RECT 4.8520 0.2565 4.8780 1.3500 ;
      RECT 4.7440 0.2565 4.7700 1.3500 ;
      RECT 4.6360 0.2565 4.6620 1.3500 ;
      RECT 4.5280 0.2565 4.5540 1.3500 ;
      RECT 4.4200 0.2565 4.4460 1.3500 ;
      RECT 4.3120 0.2565 4.3380 1.3500 ;
      RECT 4.2040 0.2565 4.2300 1.3500 ;
      RECT 4.0960 0.2565 4.1220 1.3500 ;
      RECT 3.9880 0.2565 4.0140 1.3500 ;
      RECT 3.8800 0.2565 3.9060 1.3500 ;
      RECT 3.7720 0.2565 3.7980 1.3500 ;
      RECT 3.6640 0.2565 3.6900 1.3500 ;
      RECT 3.5560 0.2565 3.5820 1.3500 ;
      RECT 3.4480 0.2565 3.4740 1.3500 ;
      RECT 3.3400 0.2565 3.3660 1.3500 ;
      RECT 3.2320 0.2565 3.2580 1.3500 ;
      RECT 3.1240 0.2565 3.1500 1.3500 ;
      RECT 3.0160 0.2565 3.0420 1.3500 ;
      RECT 2.9080 0.2565 2.9340 1.3500 ;
      RECT 2.8000 0.2565 2.8260 1.3500 ;
      RECT 2.6920 0.2565 2.7180 1.3500 ;
      RECT 2.5840 0.2565 2.6100 1.3500 ;
      RECT 2.4760 0.2565 2.5020 1.3500 ;
      RECT 2.3680 0.2565 2.3940 1.3500 ;
      RECT 2.2600 0.2565 2.2860 1.3500 ;
      RECT 2.1520 0.2565 2.1780 1.3500 ;
      RECT 2.0440 0.2565 2.0700 1.3500 ;
      RECT 1.9360 0.2565 1.9620 1.3500 ;
      RECT 1.8280 0.2565 1.8540 1.3500 ;
      RECT 1.7200 0.2565 1.7460 1.3500 ;
      RECT 1.6120 0.2565 1.6380 1.3500 ;
      RECT 1.5040 0.2565 1.5300 1.3500 ;
      RECT 1.3960 0.2565 1.4220 1.3500 ;
      RECT 1.2880 0.2565 1.3140 1.3500 ;
      RECT 1.1800 0.2565 1.2060 1.3500 ;
      RECT 1.0720 0.2565 1.0980 1.3500 ;
      RECT 0.9640 0.2565 0.9900 1.3500 ;
      RECT 0.8560 0.2565 0.8820 1.3500 ;
      RECT 0.7480 0.2565 0.7740 1.3500 ;
      RECT 0.6400 0.2565 0.6660 1.3500 ;
      RECT 0.5320 0.2565 0.5580 1.3500 ;
      RECT 0.4240 0.2565 0.4500 1.3500 ;
      RECT 0.3160 0.2565 0.3420 1.3500 ;
      RECT 0.2080 0.2565 0.2340 1.3500 ;
      RECT 0.0050 0.2565 0.0900 1.3500 ;
      RECT 8.6410 1.3365 8.7690 2.4300 ;
      RECT 8.6270 2.0020 8.7690 2.3245 ;
      RECT 8.4790 1.7290 8.5410 2.4300 ;
      RECT 8.4650 2.0385 8.5410 2.1920 ;
      RECT 8.4790 1.3365 8.5050 2.4300 ;
      RECT 8.4790 1.4575 8.5190 1.6970 ;
      RECT 8.4790 1.3365 8.5410 1.4255 ;
      RECT 8.1820 1.7870 8.3880 2.4300 ;
      RECT 8.3620 1.3365 8.3880 2.4300 ;
      RECT 8.1820 2.0640 8.4020 2.3220 ;
      RECT 8.1820 1.3365 8.2800 2.4300 ;
      RECT 7.7650 1.3365 7.8480 2.4300 ;
      RECT 7.7650 1.4250 7.8620 2.3605 ;
      RECT 16.4440 1.3365 16.5290 2.4300 ;
      RECT 16.3000 1.3365 16.3260 2.4300 ;
      RECT 16.1920 1.3365 16.2180 2.4300 ;
      RECT 16.0840 1.3365 16.1100 2.4300 ;
      RECT 15.9760 1.3365 16.0020 2.4300 ;
      RECT 15.8680 1.3365 15.8940 2.4300 ;
      RECT 15.7600 1.3365 15.7860 2.4300 ;
      RECT 15.6520 1.3365 15.6780 2.4300 ;
      RECT 15.5440 1.3365 15.5700 2.4300 ;
      RECT 15.4360 1.3365 15.4620 2.4300 ;
      RECT 15.3280 1.3365 15.3540 2.4300 ;
      RECT 15.2200 1.3365 15.2460 2.4300 ;
      RECT 15.1120 1.3365 15.1380 2.4300 ;
      RECT 15.0040 1.3365 15.0300 2.4300 ;
      RECT 14.8960 1.3365 14.9220 2.4300 ;
      RECT 14.7880 1.3365 14.8140 2.4300 ;
      RECT 14.6800 1.3365 14.7060 2.4300 ;
      RECT 14.5720 1.3365 14.5980 2.4300 ;
      RECT 14.4640 1.3365 14.4900 2.4300 ;
      RECT 14.3560 1.3365 14.3820 2.4300 ;
      RECT 14.2480 1.3365 14.2740 2.4300 ;
      RECT 14.1400 1.3365 14.1660 2.4300 ;
      RECT 14.0320 1.3365 14.0580 2.4300 ;
      RECT 13.9240 1.3365 13.9500 2.4300 ;
      RECT 13.8160 1.3365 13.8420 2.4300 ;
      RECT 13.7080 1.3365 13.7340 2.4300 ;
      RECT 13.6000 1.3365 13.6260 2.4300 ;
      RECT 13.4920 1.3365 13.5180 2.4300 ;
      RECT 13.3840 1.3365 13.4100 2.4300 ;
      RECT 13.2760 1.3365 13.3020 2.4300 ;
      RECT 13.1680 1.3365 13.1940 2.4300 ;
      RECT 13.0600 1.3365 13.0860 2.4300 ;
      RECT 12.9520 1.3365 12.9780 2.4300 ;
      RECT 12.8440 1.3365 12.8700 2.4300 ;
      RECT 12.7360 1.3365 12.7620 2.4300 ;
      RECT 12.6280 1.3365 12.6540 2.4300 ;
      RECT 12.5200 1.3365 12.5460 2.4300 ;
      RECT 12.4120 1.3365 12.4380 2.4300 ;
      RECT 12.3040 1.3365 12.3300 2.4300 ;
      RECT 12.1960 1.3365 12.2220 2.4300 ;
      RECT 12.0880 1.3365 12.1140 2.4300 ;
      RECT 11.9800 1.3365 12.0060 2.4300 ;
      RECT 11.8720 1.3365 11.8980 2.4300 ;
      RECT 11.7640 1.3365 11.7900 2.4300 ;
      RECT 11.6560 1.3365 11.6820 2.4300 ;
      RECT 11.5480 1.3365 11.5740 2.4300 ;
      RECT 11.4400 1.3365 11.4660 2.4300 ;
      RECT 11.3320 1.3365 11.3580 2.4300 ;
      RECT 11.2240 1.3365 11.2500 2.4300 ;
      RECT 11.1160 1.3365 11.1420 2.4300 ;
      RECT 11.0080 1.3365 11.0340 2.4300 ;
      RECT 10.9000 1.3365 10.9260 2.4300 ;
      RECT 10.7920 1.3365 10.8180 2.4300 ;
      RECT 10.6840 1.3365 10.7100 2.4300 ;
      RECT 10.5760 1.3365 10.6020 2.4300 ;
      RECT 10.4680 1.3365 10.4940 2.4300 ;
      RECT 10.3600 1.3365 10.3860 2.4300 ;
      RECT 10.2520 1.3365 10.2780 2.4300 ;
      RECT 10.1440 1.3365 10.1700 2.4300 ;
      RECT 10.0360 1.3365 10.0620 2.4300 ;
      RECT 9.9280 1.3365 9.9540 2.4300 ;
      RECT 9.8200 1.3365 9.8460 2.4300 ;
      RECT 9.7120 1.3365 9.7380 2.4300 ;
      RECT 9.6040 1.3365 9.6300 2.4300 ;
      RECT 9.4960 1.3365 9.5220 2.4300 ;
      RECT 9.3880 1.3365 9.4140 2.4300 ;
      RECT 9.1750 1.3365 9.2520 2.4300 ;
      RECT 7.2820 1.3365 7.3590 2.4300 ;
      RECT 7.1200 1.3365 7.1460 2.4300 ;
      RECT 7.0120 1.3365 7.0380 2.4300 ;
      RECT 6.9040 1.3365 6.9300 2.4300 ;
      RECT 6.7960 1.3365 6.8220 2.4300 ;
      RECT 6.6880 1.3365 6.7140 2.4300 ;
      RECT 6.5800 1.3365 6.6060 2.4300 ;
      RECT 6.4720 1.3365 6.4980 2.4300 ;
      RECT 6.3640 1.3365 6.3900 2.4300 ;
      RECT 6.2560 1.3365 6.2820 2.4300 ;
      RECT 6.1480 1.3365 6.1740 2.4300 ;
      RECT 6.0400 1.3365 6.0660 2.4300 ;
      RECT 5.9320 1.3365 5.9580 2.4300 ;
      RECT 5.8240 1.3365 5.8500 2.4300 ;
      RECT 5.7160 1.3365 5.7420 2.4300 ;
      RECT 5.6080 1.3365 5.6340 2.4300 ;
      RECT 5.5000 1.3365 5.5260 2.4300 ;
      RECT 5.3920 1.3365 5.4180 2.4300 ;
      RECT 5.2840 1.3365 5.3100 2.4300 ;
      RECT 5.1760 1.3365 5.2020 2.4300 ;
      RECT 5.0680 1.3365 5.0940 2.4300 ;
      RECT 4.9600 1.3365 4.9860 2.4300 ;
      RECT 4.8520 1.3365 4.8780 2.4300 ;
      RECT 4.7440 1.3365 4.7700 2.4300 ;
      RECT 4.6360 1.3365 4.6620 2.4300 ;
      RECT 4.5280 1.3365 4.5540 2.4300 ;
      RECT 4.4200 1.3365 4.4460 2.4300 ;
      RECT 4.3120 1.3365 4.3380 2.4300 ;
      RECT 4.2040 1.3365 4.2300 2.4300 ;
      RECT 4.0960 1.3365 4.1220 2.4300 ;
      RECT 3.9880 1.3365 4.0140 2.4300 ;
      RECT 3.8800 1.3365 3.9060 2.4300 ;
      RECT 3.7720 1.3365 3.7980 2.4300 ;
      RECT 3.6640 1.3365 3.6900 2.4300 ;
      RECT 3.5560 1.3365 3.5820 2.4300 ;
      RECT 3.4480 1.3365 3.4740 2.4300 ;
      RECT 3.3400 1.3365 3.3660 2.4300 ;
      RECT 3.2320 1.3365 3.2580 2.4300 ;
      RECT 3.1240 1.3365 3.1500 2.4300 ;
      RECT 3.0160 1.3365 3.0420 2.4300 ;
      RECT 2.9080 1.3365 2.9340 2.4300 ;
      RECT 2.8000 1.3365 2.8260 2.4300 ;
      RECT 2.6920 1.3365 2.7180 2.4300 ;
      RECT 2.5840 1.3365 2.6100 2.4300 ;
      RECT 2.4760 1.3365 2.5020 2.4300 ;
      RECT 2.3680 1.3365 2.3940 2.4300 ;
      RECT 2.2600 1.3365 2.2860 2.4300 ;
      RECT 2.1520 1.3365 2.1780 2.4300 ;
      RECT 2.0440 1.3365 2.0700 2.4300 ;
      RECT 1.9360 1.3365 1.9620 2.4300 ;
      RECT 1.8280 1.3365 1.8540 2.4300 ;
      RECT 1.7200 1.3365 1.7460 2.4300 ;
      RECT 1.6120 1.3365 1.6380 2.4300 ;
      RECT 1.5040 1.3365 1.5300 2.4300 ;
      RECT 1.3960 1.3365 1.4220 2.4300 ;
      RECT 1.2880 1.3365 1.3140 2.4300 ;
      RECT 1.1800 1.3365 1.2060 2.4300 ;
      RECT 1.0720 1.3365 1.0980 2.4300 ;
      RECT 0.9640 1.3365 0.9900 2.4300 ;
      RECT 0.8560 1.3365 0.8820 2.4300 ;
      RECT 0.7480 1.3365 0.7740 2.4300 ;
      RECT 0.6400 1.3365 0.6660 2.4300 ;
      RECT 0.5320 1.3365 0.5580 2.4300 ;
      RECT 0.4240 1.3365 0.4500 2.4300 ;
      RECT 0.3160 1.3365 0.3420 2.4300 ;
      RECT 0.2080 1.3365 0.2340 2.4300 ;
      RECT 0.0050 1.3365 0.0900 2.4300 ;
      RECT 8.6410 2.4165 8.7690 3.5100 ;
      RECT 8.6270 3.0820 8.7690 3.4045 ;
      RECT 8.4790 2.8090 8.5410 3.5100 ;
      RECT 8.4650 3.1185 8.5410 3.2720 ;
      RECT 8.4790 2.4165 8.5050 3.5100 ;
      RECT 8.4790 2.5375 8.5190 2.7770 ;
      RECT 8.4790 2.4165 8.5410 2.5055 ;
      RECT 8.1820 2.8670 8.3880 3.5100 ;
      RECT 8.3620 2.4165 8.3880 3.5100 ;
      RECT 8.1820 3.1440 8.4020 3.4020 ;
      RECT 8.1820 2.4165 8.2800 3.5100 ;
      RECT 7.7650 2.4165 7.8480 3.5100 ;
      RECT 7.7650 2.5050 7.8620 3.4405 ;
      RECT 16.4440 2.4165 16.5290 3.5100 ;
      RECT 16.3000 2.4165 16.3260 3.5100 ;
      RECT 16.1920 2.4165 16.2180 3.5100 ;
      RECT 16.0840 2.4165 16.1100 3.5100 ;
      RECT 15.9760 2.4165 16.0020 3.5100 ;
      RECT 15.8680 2.4165 15.8940 3.5100 ;
      RECT 15.7600 2.4165 15.7860 3.5100 ;
      RECT 15.6520 2.4165 15.6780 3.5100 ;
      RECT 15.5440 2.4165 15.5700 3.5100 ;
      RECT 15.4360 2.4165 15.4620 3.5100 ;
      RECT 15.3280 2.4165 15.3540 3.5100 ;
      RECT 15.2200 2.4165 15.2460 3.5100 ;
      RECT 15.1120 2.4165 15.1380 3.5100 ;
      RECT 15.0040 2.4165 15.0300 3.5100 ;
      RECT 14.8960 2.4165 14.9220 3.5100 ;
      RECT 14.7880 2.4165 14.8140 3.5100 ;
      RECT 14.6800 2.4165 14.7060 3.5100 ;
      RECT 14.5720 2.4165 14.5980 3.5100 ;
      RECT 14.4640 2.4165 14.4900 3.5100 ;
      RECT 14.3560 2.4165 14.3820 3.5100 ;
      RECT 14.2480 2.4165 14.2740 3.5100 ;
      RECT 14.1400 2.4165 14.1660 3.5100 ;
      RECT 14.0320 2.4165 14.0580 3.5100 ;
      RECT 13.9240 2.4165 13.9500 3.5100 ;
      RECT 13.8160 2.4165 13.8420 3.5100 ;
      RECT 13.7080 2.4165 13.7340 3.5100 ;
      RECT 13.6000 2.4165 13.6260 3.5100 ;
      RECT 13.4920 2.4165 13.5180 3.5100 ;
      RECT 13.3840 2.4165 13.4100 3.5100 ;
      RECT 13.2760 2.4165 13.3020 3.5100 ;
      RECT 13.1680 2.4165 13.1940 3.5100 ;
      RECT 13.0600 2.4165 13.0860 3.5100 ;
      RECT 12.9520 2.4165 12.9780 3.5100 ;
      RECT 12.8440 2.4165 12.8700 3.5100 ;
      RECT 12.7360 2.4165 12.7620 3.5100 ;
      RECT 12.6280 2.4165 12.6540 3.5100 ;
      RECT 12.5200 2.4165 12.5460 3.5100 ;
      RECT 12.4120 2.4165 12.4380 3.5100 ;
      RECT 12.3040 2.4165 12.3300 3.5100 ;
      RECT 12.1960 2.4165 12.2220 3.5100 ;
      RECT 12.0880 2.4165 12.1140 3.5100 ;
      RECT 11.9800 2.4165 12.0060 3.5100 ;
      RECT 11.8720 2.4165 11.8980 3.5100 ;
      RECT 11.7640 2.4165 11.7900 3.5100 ;
      RECT 11.6560 2.4165 11.6820 3.5100 ;
      RECT 11.5480 2.4165 11.5740 3.5100 ;
      RECT 11.4400 2.4165 11.4660 3.5100 ;
      RECT 11.3320 2.4165 11.3580 3.5100 ;
      RECT 11.2240 2.4165 11.2500 3.5100 ;
      RECT 11.1160 2.4165 11.1420 3.5100 ;
      RECT 11.0080 2.4165 11.0340 3.5100 ;
      RECT 10.9000 2.4165 10.9260 3.5100 ;
      RECT 10.7920 2.4165 10.8180 3.5100 ;
      RECT 10.6840 2.4165 10.7100 3.5100 ;
      RECT 10.5760 2.4165 10.6020 3.5100 ;
      RECT 10.4680 2.4165 10.4940 3.5100 ;
      RECT 10.3600 2.4165 10.3860 3.5100 ;
      RECT 10.2520 2.4165 10.2780 3.5100 ;
      RECT 10.1440 2.4165 10.1700 3.5100 ;
      RECT 10.0360 2.4165 10.0620 3.5100 ;
      RECT 9.9280 2.4165 9.9540 3.5100 ;
      RECT 9.8200 2.4165 9.8460 3.5100 ;
      RECT 9.7120 2.4165 9.7380 3.5100 ;
      RECT 9.6040 2.4165 9.6300 3.5100 ;
      RECT 9.4960 2.4165 9.5220 3.5100 ;
      RECT 9.3880 2.4165 9.4140 3.5100 ;
      RECT 9.1750 2.4165 9.2520 3.5100 ;
      RECT 7.2820 2.4165 7.3590 3.5100 ;
      RECT 7.1200 2.4165 7.1460 3.5100 ;
      RECT 7.0120 2.4165 7.0380 3.5100 ;
      RECT 6.9040 2.4165 6.9300 3.5100 ;
      RECT 6.7960 2.4165 6.8220 3.5100 ;
      RECT 6.6880 2.4165 6.7140 3.5100 ;
      RECT 6.5800 2.4165 6.6060 3.5100 ;
      RECT 6.4720 2.4165 6.4980 3.5100 ;
      RECT 6.3640 2.4165 6.3900 3.5100 ;
      RECT 6.2560 2.4165 6.2820 3.5100 ;
      RECT 6.1480 2.4165 6.1740 3.5100 ;
      RECT 6.0400 2.4165 6.0660 3.5100 ;
      RECT 5.9320 2.4165 5.9580 3.5100 ;
      RECT 5.8240 2.4165 5.8500 3.5100 ;
      RECT 5.7160 2.4165 5.7420 3.5100 ;
      RECT 5.6080 2.4165 5.6340 3.5100 ;
      RECT 5.5000 2.4165 5.5260 3.5100 ;
      RECT 5.3920 2.4165 5.4180 3.5100 ;
      RECT 5.2840 2.4165 5.3100 3.5100 ;
      RECT 5.1760 2.4165 5.2020 3.5100 ;
      RECT 5.0680 2.4165 5.0940 3.5100 ;
      RECT 4.9600 2.4165 4.9860 3.5100 ;
      RECT 4.8520 2.4165 4.8780 3.5100 ;
      RECT 4.7440 2.4165 4.7700 3.5100 ;
      RECT 4.6360 2.4165 4.6620 3.5100 ;
      RECT 4.5280 2.4165 4.5540 3.5100 ;
      RECT 4.4200 2.4165 4.4460 3.5100 ;
      RECT 4.3120 2.4165 4.3380 3.5100 ;
      RECT 4.2040 2.4165 4.2300 3.5100 ;
      RECT 4.0960 2.4165 4.1220 3.5100 ;
      RECT 3.9880 2.4165 4.0140 3.5100 ;
      RECT 3.8800 2.4165 3.9060 3.5100 ;
      RECT 3.7720 2.4165 3.7980 3.5100 ;
      RECT 3.6640 2.4165 3.6900 3.5100 ;
      RECT 3.5560 2.4165 3.5820 3.5100 ;
      RECT 3.4480 2.4165 3.4740 3.5100 ;
      RECT 3.3400 2.4165 3.3660 3.5100 ;
      RECT 3.2320 2.4165 3.2580 3.5100 ;
      RECT 3.1240 2.4165 3.1500 3.5100 ;
      RECT 3.0160 2.4165 3.0420 3.5100 ;
      RECT 2.9080 2.4165 2.9340 3.5100 ;
      RECT 2.8000 2.4165 2.8260 3.5100 ;
      RECT 2.6920 2.4165 2.7180 3.5100 ;
      RECT 2.5840 2.4165 2.6100 3.5100 ;
      RECT 2.4760 2.4165 2.5020 3.5100 ;
      RECT 2.3680 2.4165 2.3940 3.5100 ;
      RECT 2.2600 2.4165 2.2860 3.5100 ;
      RECT 2.1520 2.4165 2.1780 3.5100 ;
      RECT 2.0440 2.4165 2.0700 3.5100 ;
      RECT 1.9360 2.4165 1.9620 3.5100 ;
      RECT 1.8280 2.4165 1.8540 3.5100 ;
      RECT 1.7200 2.4165 1.7460 3.5100 ;
      RECT 1.6120 2.4165 1.6380 3.5100 ;
      RECT 1.5040 2.4165 1.5300 3.5100 ;
      RECT 1.3960 2.4165 1.4220 3.5100 ;
      RECT 1.2880 2.4165 1.3140 3.5100 ;
      RECT 1.1800 2.4165 1.2060 3.5100 ;
      RECT 1.0720 2.4165 1.0980 3.5100 ;
      RECT 0.9640 2.4165 0.9900 3.5100 ;
      RECT 0.8560 2.4165 0.8820 3.5100 ;
      RECT 0.7480 2.4165 0.7740 3.5100 ;
      RECT 0.6400 2.4165 0.6660 3.5100 ;
      RECT 0.5320 2.4165 0.5580 3.5100 ;
      RECT 0.4240 2.4165 0.4500 3.5100 ;
      RECT 0.3160 2.4165 0.3420 3.5100 ;
      RECT 0.2080 2.4165 0.2340 3.5100 ;
      RECT 0.0050 2.4165 0.0900 3.5100 ;
      RECT 8.6410 3.4965 8.7690 4.5900 ;
      RECT 8.6270 4.1620 8.7690 4.4845 ;
      RECT 8.4790 3.8890 8.5410 4.5900 ;
      RECT 8.4650 4.1985 8.5410 4.3520 ;
      RECT 8.4790 3.4965 8.5050 4.5900 ;
      RECT 8.4790 3.6175 8.5190 3.8570 ;
      RECT 8.4790 3.4965 8.5410 3.5855 ;
      RECT 8.1820 3.9470 8.3880 4.5900 ;
      RECT 8.3620 3.4965 8.3880 4.5900 ;
      RECT 8.1820 4.2240 8.4020 4.4820 ;
      RECT 8.1820 3.4965 8.2800 4.5900 ;
      RECT 7.7650 3.4965 7.8480 4.5900 ;
      RECT 7.7650 3.5850 7.8620 4.5205 ;
      RECT 16.4440 3.4965 16.5290 4.5900 ;
      RECT 16.3000 3.4965 16.3260 4.5900 ;
      RECT 16.1920 3.4965 16.2180 4.5900 ;
      RECT 16.0840 3.4965 16.1100 4.5900 ;
      RECT 15.9760 3.4965 16.0020 4.5900 ;
      RECT 15.8680 3.4965 15.8940 4.5900 ;
      RECT 15.7600 3.4965 15.7860 4.5900 ;
      RECT 15.6520 3.4965 15.6780 4.5900 ;
      RECT 15.5440 3.4965 15.5700 4.5900 ;
      RECT 15.4360 3.4965 15.4620 4.5900 ;
      RECT 15.3280 3.4965 15.3540 4.5900 ;
      RECT 15.2200 3.4965 15.2460 4.5900 ;
      RECT 15.1120 3.4965 15.1380 4.5900 ;
      RECT 15.0040 3.4965 15.0300 4.5900 ;
      RECT 14.8960 3.4965 14.9220 4.5900 ;
      RECT 14.7880 3.4965 14.8140 4.5900 ;
      RECT 14.6800 3.4965 14.7060 4.5900 ;
      RECT 14.5720 3.4965 14.5980 4.5900 ;
      RECT 14.4640 3.4965 14.4900 4.5900 ;
      RECT 14.3560 3.4965 14.3820 4.5900 ;
      RECT 14.2480 3.4965 14.2740 4.5900 ;
      RECT 14.1400 3.4965 14.1660 4.5900 ;
      RECT 14.0320 3.4965 14.0580 4.5900 ;
      RECT 13.9240 3.4965 13.9500 4.5900 ;
      RECT 13.8160 3.4965 13.8420 4.5900 ;
      RECT 13.7080 3.4965 13.7340 4.5900 ;
      RECT 13.6000 3.4965 13.6260 4.5900 ;
      RECT 13.4920 3.4965 13.5180 4.5900 ;
      RECT 13.3840 3.4965 13.4100 4.5900 ;
      RECT 13.2760 3.4965 13.3020 4.5900 ;
      RECT 13.1680 3.4965 13.1940 4.5900 ;
      RECT 13.0600 3.4965 13.0860 4.5900 ;
      RECT 12.9520 3.4965 12.9780 4.5900 ;
      RECT 12.8440 3.4965 12.8700 4.5900 ;
      RECT 12.7360 3.4965 12.7620 4.5900 ;
      RECT 12.6280 3.4965 12.6540 4.5900 ;
      RECT 12.5200 3.4965 12.5460 4.5900 ;
      RECT 12.4120 3.4965 12.4380 4.5900 ;
      RECT 12.3040 3.4965 12.3300 4.5900 ;
      RECT 12.1960 3.4965 12.2220 4.5900 ;
      RECT 12.0880 3.4965 12.1140 4.5900 ;
      RECT 11.9800 3.4965 12.0060 4.5900 ;
      RECT 11.8720 3.4965 11.8980 4.5900 ;
      RECT 11.7640 3.4965 11.7900 4.5900 ;
      RECT 11.6560 3.4965 11.6820 4.5900 ;
      RECT 11.5480 3.4965 11.5740 4.5900 ;
      RECT 11.4400 3.4965 11.4660 4.5900 ;
      RECT 11.3320 3.4965 11.3580 4.5900 ;
      RECT 11.2240 3.4965 11.2500 4.5900 ;
      RECT 11.1160 3.4965 11.1420 4.5900 ;
      RECT 11.0080 3.4965 11.0340 4.5900 ;
      RECT 10.9000 3.4965 10.9260 4.5900 ;
      RECT 10.7920 3.4965 10.8180 4.5900 ;
      RECT 10.6840 3.4965 10.7100 4.5900 ;
      RECT 10.5760 3.4965 10.6020 4.5900 ;
      RECT 10.4680 3.4965 10.4940 4.5900 ;
      RECT 10.3600 3.4965 10.3860 4.5900 ;
      RECT 10.2520 3.4965 10.2780 4.5900 ;
      RECT 10.1440 3.4965 10.1700 4.5900 ;
      RECT 10.0360 3.4965 10.0620 4.5900 ;
      RECT 9.9280 3.4965 9.9540 4.5900 ;
      RECT 9.8200 3.4965 9.8460 4.5900 ;
      RECT 9.7120 3.4965 9.7380 4.5900 ;
      RECT 9.6040 3.4965 9.6300 4.5900 ;
      RECT 9.4960 3.4965 9.5220 4.5900 ;
      RECT 9.3880 3.4965 9.4140 4.5900 ;
      RECT 9.1750 3.4965 9.2520 4.5900 ;
      RECT 7.2820 3.4965 7.3590 4.5900 ;
      RECT 7.1200 3.4965 7.1460 4.5900 ;
      RECT 7.0120 3.4965 7.0380 4.5900 ;
      RECT 6.9040 3.4965 6.9300 4.5900 ;
      RECT 6.7960 3.4965 6.8220 4.5900 ;
      RECT 6.6880 3.4965 6.7140 4.5900 ;
      RECT 6.5800 3.4965 6.6060 4.5900 ;
      RECT 6.4720 3.4965 6.4980 4.5900 ;
      RECT 6.3640 3.4965 6.3900 4.5900 ;
      RECT 6.2560 3.4965 6.2820 4.5900 ;
      RECT 6.1480 3.4965 6.1740 4.5900 ;
      RECT 6.0400 3.4965 6.0660 4.5900 ;
      RECT 5.9320 3.4965 5.9580 4.5900 ;
      RECT 5.8240 3.4965 5.8500 4.5900 ;
      RECT 5.7160 3.4965 5.7420 4.5900 ;
      RECT 5.6080 3.4965 5.6340 4.5900 ;
      RECT 5.5000 3.4965 5.5260 4.5900 ;
      RECT 5.3920 3.4965 5.4180 4.5900 ;
      RECT 5.2840 3.4965 5.3100 4.5900 ;
      RECT 5.1760 3.4965 5.2020 4.5900 ;
      RECT 5.0680 3.4965 5.0940 4.5900 ;
      RECT 4.9600 3.4965 4.9860 4.5900 ;
      RECT 4.8520 3.4965 4.8780 4.5900 ;
      RECT 4.7440 3.4965 4.7700 4.5900 ;
      RECT 4.6360 3.4965 4.6620 4.5900 ;
      RECT 4.5280 3.4965 4.5540 4.5900 ;
      RECT 4.4200 3.4965 4.4460 4.5900 ;
      RECT 4.3120 3.4965 4.3380 4.5900 ;
      RECT 4.2040 3.4965 4.2300 4.5900 ;
      RECT 4.0960 3.4965 4.1220 4.5900 ;
      RECT 3.9880 3.4965 4.0140 4.5900 ;
      RECT 3.8800 3.4965 3.9060 4.5900 ;
      RECT 3.7720 3.4965 3.7980 4.5900 ;
      RECT 3.6640 3.4965 3.6900 4.5900 ;
      RECT 3.5560 3.4965 3.5820 4.5900 ;
      RECT 3.4480 3.4965 3.4740 4.5900 ;
      RECT 3.3400 3.4965 3.3660 4.5900 ;
      RECT 3.2320 3.4965 3.2580 4.5900 ;
      RECT 3.1240 3.4965 3.1500 4.5900 ;
      RECT 3.0160 3.4965 3.0420 4.5900 ;
      RECT 2.9080 3.4965 2.9340 4.5900 ;
      RECT 2.8000 3.4965 2.8260 4.5900 ;
      RECT 2.6920 3.4965 2.7180 4.5900 ;
      RECT 2.5840 3.4965 2.6100 4.5900 ;
      RECT 2.4760 3.4965 2.5020 4.5900 ;
      RECT 2.3680 3.4965 2.3940 4.5900 ;
      RECT 2.2600 3.4965 2.2860 4.5900 ;
      RECT 2.1520 3.4965 2.1780 4.5900 ;
      RECT 2.0440 3.4965 2.0700 4.5900 ;
      RECT 1.9360 3.4965 1.9620 4.5900 ;
      RECT 1.8280 3.4965 1.8540 4.5900 ;
      RECT 1.7200 3.4965 1.7460 4.5900 ;
      RECT 1.6120 3.4965 1.6380 4.5900 ;
      RECT 1.5040 3.4965 1.5300 4.5900 ;
      RECT 1.3960 3.4965 1.4220 4.5900 ;
      RECT 1.2880 3.4965 1.3140 4.5900 ;
      RECT 1.1800 3.4965 1.2060 4.5900 ;
      RECT 1.0720 3.4965 1.0980 4.5900 ;
      RECT 0.9640 3.4965 0.9900 4.5900 ;
      RECT 0.8560 3.4965 0.8820 4.5900 ;
      RECT 0.7480 3.4965 0.7740 4.5900 ;
      RECT 0.6400 3.4965 0.6660 4.5900 ;
      RECT 0.5320 3.4965 0.5580 4.5900 ;
      RECT 0.4240 3.4965 0.4500 4.5900 ;
      RECT 0.3160 3.4965 0.3420 4.5900 ;
      RECT 0.2080 3.4965 0.2340 4.5900 ;
      RECT 0.0050 3.4965 0.0900 4.5900 ;
      RECT 8.6410 4.5765 8.7690 5.6700 ;
      RECT 8.6270 5.2420 8.7690 5.5645 ;
      RECT 8.4790 4.9690 8.5410 5.6700 ;
      RECT 8.4650 5.2785 8.5410 5.4320 ;
      RECT 8.4790 4.5765 8.5050 5.6700 ;
      RECT 8.4790 4.6975 8.5190 4.9370 ;
      RECT 8.4790 4.5765 8.5410 4.6655 ;
      RECT 8.1820 5.0270 8.3880 5.6700 ;
      RECT 8.3620 4.5765 8.3880 5.6700 ;
      RECT 8.1820 5.3040 8.4020 5.5620 ;
      RECT 8.1820 4.5765 8.2800 5.6700 ;
      RECT 7.7650 4.5765 7.8480 5.6700 ;
      RECT 7.7650 4.6650 7.8620 5.6005 ;
      RECT 16.4440 4.5765 16.5290 5.6700 ;
      RECT 16.3000 4.5765 16.3260 5.6700 ;
      RECT 16.1920 4.5765 16.2180 5.6700 ;
      RECT 16.0840 4.5765 16.1100 5.6700 ;
      RECT 15.9760 4.5765 16.0020 5.6700 ;
      RECT 15.8680 4.5765 15.8940 5.6700 ;
      RECT 15.7600 4.5765 15.7860 5.6700 ;
      RECT 15.6520 4.5765 15.6780 5.6700 ;
      RECT 15.5440 4.5765 15.5700 5.6700 ;
      RECT 15.4360 4.5765 15.4620 5.6700 ;
      RECT 15.3280 4.5765 15.3540 5.6700 ;
      RECT 15.2200 4.5765 15.2460 5.6700 ;
      RECT 15.1120 4.5765 15.1380 5.6700 ;
      RECT 15.0040 4.5765 15.0300 5.6700 ;
      RECT 14.8960 4.5765 14.9220 5.6700 ;
      RECT 14.7880 4.5765 14.8140 5.6700 ;
      RECT 14.6800 4.5765 14.7060 5.6700 ;
      RECT 14.5720 4.5765 14.5980 5.6700 ;
      RECT 14.4640 4.5765 14.4900 5.6700 ;
      RECT 14.3560 4.5765 14.3820 5.6700 ;
      RECT 14.2480 4.5765 14.2740 5.6700 ;
      RECT 14.1400 4.5765 14.1660 5.6700 ;
      RECT 14.0320 4.5765 14.0580 5.6700 ;
      RECT 13.9240 4.5765 13.9500 5.6700 ;
      RECT 13.8160 4.5765 13.8420 5.6700 ;
      RECT 13.7080 4.5765 13.7340 5.6700 ;
      RECT 13.6000 4.5765 13.6260 5.6700 ;
      RECT 13.4920 4.5765 13.5180 5.6700 ;
      RECT 13.3840 4.5765 13.4100 5.6700 ;
      RECT 13.2760 4.5765 13.3020 5.6700 ;
      RECT 13.1680 4.5765 13.1940 5.6700 ;
      RECT 13.0600 4.5765 13.0860 5.6700 ;
      RECT 12.9520 4.5765 12.9780 5.6700 ;
      RECT 12.8440 4.5765 12.8700 5.6700 ;
      RECT 12.7360 4.5765 12.7620 5.6700 ;
      RECT 12.6280 4.5765 12.6540 5.6700 ;
      RECT 12.5200 4.5765 12.5460 5.6700 ;
      RECT 12.4120 4.5765 12.4380 5.6700 ;
      RECT 12.3040 4.5765 12.3300 5.6700 ;
      RECT 12.1960 4.5765 12.2220 5.6700 ;
      RECT 12.0880 4.5765 12.1140 5.6700 ;
      RECT 11.9800 4.5765 12.0060 5.6700 ;
      RECT 11.8720 4.5765 11.8980 5.6700 ;
      RECT 11.7640 4.5765 11.7900 5.6700 ;
      RECT 11.6560 4.5765 11.6820 5.6700 ;
      RECT 11.5480 4.5765 11.5740 5.6700 ;
      RECT 11.4400 4.5765 11.4660 5.6700 ;
      RECT 11.3320 4.5765 11.3580 5.6700 ;
      RECT 11.2240 4.5765 11.2500 5.6700 ;
      RECT 11.1160 4.5765 11.1420 5.6700 ;
      RECT 11.0080 4.5765 11.0340 5.6700 ;
      RECT 10.9000 4.5765 10.9260 5.6700 ;
      RECT 10.7920 4.5765 10.8180 5.6700 ;
      RECT 10.6840 4.5765 10.7100 5.6700 ;
      RECT 10.5760 4.5765 10.6020 5.6700 ;
      RECT 10.4680 4.5765 10.4940 5.6700 ;
      RECT 10.3600 4.5765 10.3860 5.6700 ;
      RECT 10.2520 4.5765 10.2780 5.6700 ;
      RECT 10.1440 4.5765 10.1700 5.6700 ;
      RECT 10.0360 4.5765 10.0620 5.6700 ;
      RECT 9.9280 4.5765 9.9540 5.6700 ;
      RECT 9.8200 4.5765 9.8460 5.6700 ;
      RECT 9.7120 4.5765 9.7380 5.6700 ;
      RECT 9.6040 4.5765 9.6300 5.6700 ;
      RECT 9.4960 4.5765 9.5220 5.6700 ;
      RECT 9.3880 4.5765 9.4140 5.6700 ;
      RECT 9.1750 4.5765 9.2520 5.6700 ;
      RECT 7.2820 4.5765 7.3590 5.6700 ;
      RECT 7.1200 4.5765 7.1460 5.6700 ;
      RECT 7.0120 4.5765 7.0380 5.6700 ;
      RECT 6.9040 4.5765 6.9300 5.6700 ;
      RECT 6.7960 4.5765 6.8220 5.6700 ;
      RECT 6.6880 4.5765 6.7140 5.6700 ;
      RECT 6.5800 4.5765 6.6060 5.6700 ;
      RECT 6.4720 4.5765 6.4980 5.6700 ;
      RECT 6.3640 4.5765 6.3900 5.6700 ;
      RECT 6.2560 4.5765 6.2820 5.6700 ;
      RECT 6.1480 4.5765 6.1740 5.6700 ;
      RECT 6.0400 4.5765 6.0660 5.6700 ;
      RECT 5.9320 4.5765 5.9580 5.6700 ;
      RECT 5.8240 4.5765 5.8500 5.6700 ;
      RECT 5.7160 4.5765 5.7420 5.6700 ;
      RECT 5.6080 4.5765 5.6340 5.6700 ;
      RECT 5.5000 4.5765 5.5260 5.6700 ;
      RECT 5.3920 4.5765 5.4180 5.6700 ;
      RECT 5.2840 4.5765 5.3100 5.6700 ;
      RECT 5.1760 4.5765 5.2020 5.6700 ;
      RECT 5.0680 4.5765 5.0940 5.6700 ;
      RECT 4.9600 4.5765 4.9860 5.6700 ;
      RECT 4.8520 4.5765 4.8780 5.6700 ;
      RECT 4.7440 4.5765 4.7700 5.6700 ;
      RECT 4.6360 4.5765 4.6620 5.6700 ;
      RECT 4.5280 4.5765 4.5540 5.6700 ;
      RECT 4.4200 4.5765 4.4460 5.6700 ;
      RECT 4.3120 4.5765 4.3380 5.6700 ;
      RECT 4.2040 4.5765 4.2300 5.6700 ;
      RECT 4.0960 4.5765 4.1220 5.6700 ;
      RECT 3.9880 4.5765 4.0140 5.6700 ;
      RECT 3.8800 4.5765 3.9060 5.6700 ;
      RECT 3.7720 4.5765 3.7980 5.6700 ;
      RECT 3.6640 4.5765 3.6900 5.6700 ;
      RECT 3.5560 4.5765 3.5820 5.6700 ;
      RECT 3.4480 4.5765 3.4740 5.6700 ;
      RECT 3.3400 4.5765 3.3660 5.6700 ;
      RECT 3.2320 4.5765 3.2580 5.6700 ;
      RECT 3.1240 4.5765 3.1500 5.6700 ;
      RECT 3.0160 4.5765 3.0420 5.6700 ;
      RECT 2.9080 4.5765 2.9340 5.6700 ;
      RECT 2.8000 4.5765 2.8260 5.6700 ;
      RECT 2.6920 4.5765 2.7180 5.6700 ;
      RECT 2.5840 4.5765 2.6100 5.6700 ;
      RECT 2.4760 4.5765 2.5020 5.6700 ;
      RECT 2.3680 4.5765 2.3940 5.6700 ;
      RECT 2.2600 4.5765 2.2860 5.6700 ;
      RECT 2.1520 4.5765 2.1780 5.6700 ;
      RECT 2.0440 4.5765 2.0700 5.6700 ;
      RECT 1.9360 4.5765 1.9620 5.6700 ;
      RECT 1.8280 4.5765 1.8540 5.6700 ;
      RECT 1.7200 4.5765 1.7460 5.6700 ;
      RECT 1.6120 4.5765 1.6380 5.6700 ;
      RECT 1.5040 4.5765 1.5300 5.6700 ;
      RECT 1.3960 4.5765 1.4220 5.6700 ;
      RECT 1.2880 4.5765 1.3140 5.6700 ;
      RECT 1.1800 4.5765 1.2060 5.6700 ;
      RECT 1.0720 4.5765 1.0980 5.6700 ;
      RECT 0.9640 4.5765 0.9900 5.6700 ;
      RECT 0.8560 4.5765 0.8820 5.6700 ;
      RECT 0.7480 4.5765 0.7740 5.6700 ;
      RECT 0.6400 4.5765 0.6660 5.6700 ;
      RECT 0.5320 4.5765 0.5580 5.6700 ;
      RECT 0.4240 4.5765 0.4500 5.6700 ;
      RECT 0.3160 4.5765 0.3420 5.6700 ;
      RECT 0.2080 4.5765 0.2340 5.6700 ;
      RECT 0.0050 4.5765 0.0900 5.6700 ;
      RECT 8.6410 5.6565 8.7690 6.7500 ;
      RECT 8.6270 6.3220 8.7690 6.6445 ;
      RECT 8.4790 6.0490 8.5410 6.7500 ;
      RECT 8.4650 6.3585 8.5410 6.5120 ;
      RECT 8.4790 5.6565 8.5050 6.7500 ;
      RECT 8.4790 5.7775 8.5190 6.0170 ;
      RECT 8.4790 5.6565 8.5410 5.7455 ;
      RECT 8.1820 6.1070 8.3880 6.7500 ;
      RECT 8.3620 5.6565 8.3880 6.7500 ;
      RECT 8.1820 6.3840 8.4020 6.6420 ;
      RECT 8.1820 5.6565 8.2800 6.7500 ;
      RECT 7.7650 5.6565 7.8480 6.7500 ;
      RECT 7.7650 5.7450 7.8620 6.6805 ;
      RECT 16.4440 5.6565 16.5290 6.7500 ;
      RECT 16.3000 5.6565 16.3260 6.7500 ;
      RECT 16.1920 5.6565 16.2180 6.7500 ;
      RECT 16.0840 5.6565 16.1100 6.7500 ;
      RECT 15.9760 5.6565 16.0020 6.7500 ;
      RECT 15.8680 5.6565 15.8940 6.7500 ;
      RECT 15.7600 5.6565 15.7860 6.7500 ;
      RECT 15.6520 5.6565 15.6780 6.7500 ;
      RECT 15.5440 5.6565 15.5700 6.7500 ;
      RECT 15.4360 5.6565 15.4620 6.7500 ;
      RECT 15.3280 5.6565 15.3540 6.7500 ;
      RECT 15.2200 5.6565 15.2460 6.7500 ;
      RECT 15.1120 5.6565 15.1380 6.7500 ;
      RECT 15.0040 5.6565 15.0300 6.7500 ;
      RECT 14.8960 5.6565 14.9220 6.7500 ;
      RECT 14.7880 5.6565 14.8140 6.7500 ;
      RECT 14.6800 5.6565 14.7060 6.7500 ;
      RECT 14.5720 5.6565 14.5980 6.7500 ;
      RECT 14.4640 5.6565 14.4900 6.7500 ;
      RECT 14.3560 5.6565 14.3820 6.7500 ;
      RECT 14.2480 5.6565 14.2740 6.7500 ;
      RECT 14.1400 5.6565 14.1660 6.7500 ;
      RECT 14.0320 5.6565 14.0580 6.7500 ;
      RECT 13.9240 5.6565 13.9500 6.7500 ;
      RECT 13.8160 5.6565 13.8420 6.7500 ;
      RECT 13.7080 5.6565 13.7340 6.7500 ;
      RECT 13.6000 5.6565 13.6260 6.7500 ;
      RECT 13.4920 5.6565 13.5180 6.7500 ;
      RECT 13.3840 5.6565 13.4100 6.7500 ;
      RECT 13.2760 5.6565 13.3020 6.7500 ;
      RECT 13.1680 5.6565 13.1940 6.7500 ;
      RECT 13.0600 5.6565 13.0860 6.7500 ;
      RECT 12.9520 5.6565 12.9780 6.7500 ;
      RECT 12.8440 5.6565 12.8700 6.7500 ;
      RECT 12.7360 5.6565 12.7620 6.7500 ;
      RECT 12.6280 5.6565 12.6540 6.7500 ;
      RECT 12.5200 5.6565 12.5460 6.7500 ;
      RECT 12.4120 5.6565 12.4380 6.7500 ;
      RECT 12.3040 5.6565 12.3300 6.7500 ;
      RECT 12.1960 5.6565 12.2220 6.7500 ;
      RECT 12.0880 5.6565 12.1140 6.7500 ;
      RECT 11.9800 5.6565 12.0060 6.7500 ;
      RECT 11.8720 5.6565 11.8980 6.7500 ;
      RECT 11.7640 5.6565 11.7900 6.7500 ;
      RECT 11.6560 5.6565 11.6820 6.7500 ;
      RECT 11.5480 5.6565 11.5740 6.7500 ;
      RECT 11.4400 5.6565 11.4660 6.7500 ;
      RECT 11.3320 5.6565 11.3580 6.7500 ;
      RECT 11.2240 5.6565 11.2500 6.7500 ;
      RECT 11.1160 5.6565 11.1420 6.7500 ;
      RECT 11.0080 5.6565 11.0340 6.7500 ;
      RECT 10.9000 5.6565 10.9260 6.7500 ;
      RECT 10.7920 5.6565 10.8180 6.7500 ;
      RECT 10.6840 5.6565 10.7100 6.7500 ;
      RECT 10.5760 5.6565 10.6020 6.7500 ;
      RECT 10.4680 5.6565 10.4940 6.7500 ;
      RECT 10.3600 5.6565 10.3860 6.7500 ;
      RECT 10.2520 5.6565 10.2780 6.7500 ;
      RECT 10.1440 5.6565 10.1700 6.7500 ;
      RECT 10.0360 5.6565 10.0620 6.7500 ;
      RECT 9.9280 5.6565 9.9540 6.7500 ;
      RECT 9.8200 5.6565 9.8460 6.7500 ;
      RECT 9.7120 5.6565 9.7380 6.7500 ;
      RECT 9.6040 5.6565 9.6300 6.7500 ;
      RECT 9.4960 5.6565 9.5220 6.7500 ;
      RECT 9.3880 5.6565 9.4140 6.7500 ;
      RECT 9.1750 5.6565 9.2520 6.7500 ;
      RECT 7.2820 5.6565 7.3590 6.7500 ;
      RECT 7.1200 5.6565 7.1460 6.7500 ;
      RECT 7.0120 5.6565 7.0380 6.7500 ;
      RECT 6.9040 5.6565 6.9300 6.7500 ;
      RECT 6.7960 5.6565 6.8220 6.7500 ;
      RECT 6.6880 5.6565 6.7140 6.7500 ;
      RECT 6.5800 5.6565 6.6060 6.7500 ;
      RECT 6.4720 5.6565 6.4980 6.7500 ;
      RECT 6.3640 5.6565 6.3900 6.7500 ;
      RECT 6.2560 5.6565 6.2820 6.7500 ;
      RECT 6.1480 5.6565 6.1740 6.7500 ;
      RECT 6.0400 5.6565 6.0660 6.7500 ;
      RECT 5.9320 5.6565 5.9580 6.7500 ;
      RECT 5.8240 5.6565 5.8500 6.7500 ;
      RECT 5.7160 5.6565 5.7420 6.7500 ;
      RECT 5.6080 5.6565 5.6340 6.7500 ;
      RECT 5.5000 5.6565 5.5260 6.7500 ;
      RECT 5.3920 5.6565 5.4180 6.7500 ;
      RECT 5.2840 5.6565 5.3100 6.7500 ;
      RECT 5.1760 5.6565 5.2020 6.7500 ;
      RECT 5.0680 5.6565 5.0940 6.7500 ;
      RECT 4.9600 5.6565 4.9860 6.7500 ;
      RECT 4.8520 5.6565 4.8780 6.7500 ;
      RECT 4.7440 5.6565 4.7700 6.7500 ;
      RECT 4.6360 5.6565 4.6620 6.7500 ;
      RECT 4.5280 5.6565 4.5540 6.7500 ;
      RECT 4.4200 5.6565 4.4460 6.7500 ;
      RECT 4.3120 5.6565 4.3380 6.7500 ;
      RECT 4.2040 5.6565 4.2300 6.7500 ;
      RECT 4.0960 5.6565 4.1220 6.7500 ;
      RECT 3.9880 5.6565 4.0140 6.7500 ;
      RECT 3.8800 5.6565 3.9060 6.7500 ;
      RECT 3.7720 5.6565 3.7980 6.7500 ;
      RECT 3.6640 5.6565 3.6900 6.7500 ;
      RECT 3.5560 5.6565 3.5820 6.7500 ;
      RECT 3.4480 5.6565 3.4740 6.7500 ;
      RECT 3.3400 5.6565 3.3660 6.7500 ;
      RECT 3.2320 5.6565 3.2580 6.7500 ;
      RECT 3.1240 5.6565 3.1500 6.7500 ;
      RECT 3.0160 5.6565 3.0420 6.7500 ;
      RECT 2.9080 5.6565 2.9340 6.7500 ;
      RECT 2.8000 5.6565 2.8260 6.7500 ;
      RECT 2.6920 5.6565 2.7180 6.7500 ;
      RECT 2.5840 5.6565 2.6100 6.7500 ;
      RECT 2.4760 5.6565 2.5020 6.7500 ;
      RECT 2.3680 5.6565 2.3940 6.7500 ;
      RECT 2.2600 5.6565 2.2860 6.7500 ;
      RECT 2.1520 5.6565 2.1780 6.7500 ;
      RECT 2.0440 5.6565 2.0700 6.7500 ;
      RECT 1.9360 5.6565 1.9620 6.7500 ;
      RECT 1.8280 5.6565 1.8540 6.7500 ;
      RECT 1.7200 5.6565 1.7460 6.7500 ;
      RECT 1.6120 5.6565 1.6380 6.7500 ;
      RECT 1.5040 5.6565 1.5300 6.7500 ;
      RECT 1.3960 5.6565 1.4220 6.7500 ;
      RECT 1.2880 5.6565 1.3140 6.7500 ;
      RECT 1.1800 5.6565 1.2060 6.7500 ;
      RECT 1.0720 5.6565 1.0980 6.7500 ;
      RECT 0.9640 5.6565 0.9900 6.7500 ;
      RECT 0.8560 5.6565 0.8820 6.7500 ;
      RECT 0.7480 5.6565 0.7740 6.7500 ;
      RECT 0.6400 5.6565 0.6660 6.7500 ;
      RECT 0.5320 5.6565 0.5580 6.7500 ;
      RECT 0.4240 5.6565 0.4500 6.7500 ;
      RECT 0.3160 5.6565 0.3420 6.7500 ;
      RECT 0.2080 5.6565 0.2340 6.7500 ;
      RECT 0.0050 5.6565 0.0900 6.7500 ;
      RECT 8.6410 6.7365 8.7690 7.8300 ;
      RECT 8.6270 7.4020 8.7690 7.7245 ;
      RECT 8.4790 7.1290 8.5410 7.8300 ;
      RECT 8.4650 7.4385 8.5410 7.5920 ;
      RECT 8.4790 6.7365 8.5050 7.8300 ;
      RECT 8.4790 6.8575 8.5190 7.0970 ;
      RECT 8.4790 6.7365 8.5410 6.8255 ;
      RECT 8.1820 7.1870 8.3880 7.8300 ;
      RECT 8.3620 6.7365 8.3880 7.8300 ;
      RECT 8.1820 7.4640 8.4020 7.7220 ;
      RECT 8.1820 6.7365 8.2800 7.8300 ;
      RECT 7.7650 6.7365 7.8480 7.8300 ;
      RECT 7.7650 6.8250 7.8620 7.7605 ;
      RECT 16.4440 6.7365 16.5290 7.8300 ;
      RECT 16.3000 6.7365 16.3260 7.8300 ;
      RECT 16.1920 6.7365 16.2180 7.8300 ;
      RECT 16.0840 6.7365 16.1100 7.8300 ;
      RECT 15.9760 6.7365 16.0020 7.8300 ;
      RECT 15.8680 6.7365 15.8940 7.8300 ;
      RECT 15.7600 6.7365 15.7860 7.8300 ;
      RECT 15.6520 6.7365 15.6780 7.8300 ;
      RECT 15.5440 6.7365 15.5700 7.8300 ;
      RECT 15.4360 6.7365 15.4620 7.8300 ;
      RECT 15.3280 6.7365 15.3540 7.8300 ;
      RECT 15.2200 6.7365 15.2460 7.8300 ;
      RECT 15.1120 6.7365 15.1380 7.8300 ;
      RECT 15.0040 6.7365 15.0300 7.8300 ;
      RECT 14.8960 6.7365 14.9220 7.8300 ;
      RECT 14.7880 6.7365 14.8140 7.8300 ;
      RECT 14.6800 6.7365 14.7060 7.8300 ;
      RECT 14.5720 6.7365 14.5980 7.8300 ;
      RECT 14.4640 6.7365 14.4900 7.8300 ;
      RECT 14.3560 6.7365 14.3820 7.8300 ;
      RECT 14.2480 6.7365 14.2740 7.8300 ;
      RECT 14.1400 6.7365 14.1660 7.8300 ;
      RECT 14.0320 6.7365 14.0580 7.8300 ;
      RECT 13.9240 6.7365 13.9500 7.8300 ;
      RECT 13.8160 6.7365 13.8420 7.8300 ;
      RECT 13.7080 6.7365 13.7340 7.8300 ;
      RECT 13.6000 6.7365 13.6260 7.8300 ;
      RECT 13.4920 6.7365 13.5180 7.8300 ;
      RECT 13.3840 6.7365 13.4100 7.8300 ;
      RECT 13.2760 6.7365 13.3020 7.8300 ;
      RECT 13.1680 6.7365 13.1940 7.8300 ;
      RECT 13.0600 6.7365 13.0860 7.8300 ;
      RECT 12.9520 6.7365 12.9780 7.8300 ;
      RECT 12.8440 6.7365 12.8700 7.8300 ;
      RECT 12.7360 6.7365 12.7620 7.8300 ;
      RECT 12.6280 6.7365 12.6540 7.8300 ;
      RECT 12.5200 6.7365 12.5460 7.8300 ;
      RECT 12.4120 6.7365 12.4380 7.8300 ;
      RECT 12.3040 6.7365 12.3300 7.8300 ;
      RECT 12.1960 6.7365 12.2220 7.8300 ;
      RECT 12.0880 6.7365 12.1140 7.8300 ;
      RECT 11.9800 6.7365 12.0060 7.8300 ;
      RECT 11.8720 6.7365 11.8980 7.8300 ;
      RECT 11.7640 6.7365 11.7900 7.8300 ;
      RECT 11.6560 6.7365 11.6820 7.8300 ;
      RECT 11.5480 6.7365 11.5740 7.8300 ;
      RECT 11.4400 6.7365 11.4660 7.8300 ;
      RECT 11.3320 6.7365 11.3580 7.8300 ;
      RECT 11.2240 6.7365 11.2500 7.8300 ;
      RECT 11.1160 6.7365 11.1420 7.8300 ;
      RECT 11.0080 6.7365 11.0340 7.8300 ;
      RECT 10.9000 6.7365 10.9260 7.8300 ;
      RECT 10.7920 6.7365 10.8180 7.8300 ;
      RECT 10.6840 6.7365 10.7100 7.8300 ;
      RECT 10.5760 6.7365 10.6020 7.8300 ;
      RECT 10.4680 6.7365 10.4940 7.8300 ;
      RECT 10.3600 6.7365 10.3860 7.8300 ;
      RECT 10.2520 6.7365 10.2780 7.8300 ;
      RECT 10.1440 6.7365 10.1700 7.8300 ;
      RECT 10.0360 6.7365 10.0620 7.8300 ;
      RECT 9.9280 6.7365 9.9540 7.8300 ;
      RECT 9.8200 6.7365 9.8460 7.8300 ;
      RECT 9.7120 6.7365 9.7380 7.8300 ;
      RECT 9.6040 6.7365 9.6300 7.8300 ;
      RECT 9.4960 6.7365 9.5220 7.8300 ;
      RECT 9.3880 6.7365 9.4140 7.8300 ;
      RECT 9.1750 6.7365 9.2520 7.8300 ;
      RECT 7.2820 6.7365 7.3590 7.8300 ;
      RECT 7.1200 6.7365 7.1460 7.8300 ;
      RECT 7.0120 6.7365 7.0380 7.8300 ;
      RECT 6.9040 6.7365 6.9300 7.8300 ;
      RECT 6.7960 6.7365 6.8220 7.8300 ;
      RECT 6.6880 6.7365 6.7140 7.8300 ;
      RECT 6.5800 6.7365 6.6060 7.8300 ;
      RECT 6.4720 6.7365 6.4980 7.8300 ;
      RECT 6.3640 6.7365 6.3900 7.8300 ;
      RECT 6.2560 6.7365 6.2820 7.8300 ;
      RECT 6.1480 6.7365 6.1740 7.8300 ;
      RECT 6.0400 6.7365 6.0660 7.8300 ;
      RECT 5.9320 6.7365 5.9580 7.8300 ;
      RECT 5.8240 6.7365 5.8500 7.8300 ;
      RECT 5.7160 6.7365 5.7420 7.8300 ;
      RECT 5.6080 6.7365 5.6340 7.8300 ;
      RECT 5.5000 6.7365 5.5260 7.8300 ;
      RECT 5.3920 6.7365 5.4180 7.8300 ;
      RECT 5.2840 6.7365 5.3100 7.8300 ;
      RECT 5.1760 6.7365 5.2020 7.8300 ;
      RECT 5.0680 6.7365 5.0940 7.8300 ;
      RECT 4.9600 6.7365 4.9860 7.8300 ;
      RECT 4.8520 6.7365 4.8780 7.8300 ;
      RECT 4.7440 6.7365 4.7700 7.8300 ;
      RECT 4.6360 6.7365 4.6620 7.8300 ;
      RECT 4.5280 6.7365 4.5540 7.8300 ;
      RECT 4.4200 6.7365 4.4460 7.8300 ;
      RECT 4.3120 6.7365 4.3380 7.8300 ;
      RECT 4.2040 6.7365 4.2300 7.8300 ;
      RECT 4.0960 6.7365 4.1220 7.8300 ;
      RECT 3.9880 6.7365 4.0140 7.8300 ;
      RECT 3.8800 6.7365 3.9060 7.8300 ;
      RECT 3.7720 6.7365 3.7980 7.8300 ;
      RECT 3.6640 6.7365 3.6900 7.8300 ;
      RECT 3.5560 6.7365 3.5820 7.8300 ;
      RECT 3.4480 6.7365 3.4740 7.8300 ;
      RECT 3.3400 6.7365 3.3660 7.8300 ;
      RECT 3.2320 6.7365 3.2580 7.8300 ;
      RECT 3.1240 6.7365 3.1500 7.8300 ;
      RECT 3.0160 6.7365 3.0420 7.8300 ;
      RECT 2.9080 6.7365 2.9340 7.8300 ;
      RECT 2.8000 6.7365 2.8260 7.8300 ;
      RECT 2.6920 6.7365 2.7180 7.8300 ;
      RECT 2.5840 6.7365 2.6100 7.8300 ;
      RECT 2.4760 6.7365 2.5020 7.8300 ;
      RECT 2.3680 6.7365 2.3940 7.8300 ;
      RECT 2.2600 6.7365 2.2860 7.8300 ;
      RECT 2.1520 6.7365 2.1780 7.8300 ;
      RECT 2.0440 6.7365 2.0700 7.8300 ;
      RECT 1.9360 6.7365 1.9620 7.8300 ;
      RECT 1.8280 6.7365 1.8540 7.8300 ;
      RECT 1.7200 6.7365 1.7460 7.8300 ;
      RECT 1.6120 6.7365 1.6380 7.8300 ;
      RECT 1.5040 6.7365 1.5300 7.8300 ;
      RECT 1.3960 6.7365 1.4220 7.8300 ;
      RECT 1.2880 6.7365 1.3140 7.8300 ;
      RECT 1.1800 6.7365 1.2060 7.8300 ;
      RECT 1.0720 6.7365 1.0980 7.8300 ;
      RECT 0.9640 6.7365 0.9900 7.8300 ;
      RECT 0.8560 6.7365 0.8820 7.8300 ;
      RECT 0.7480 6.7365 0.7740 7.8300 ;
      RECT 0.6400 6.7365 0.6660 7.8300 ;
      RECT 0.5320 6.7365 0.5580 7.8300 ;
      RECT 0.4240 6.7365 0.4500 7.8300 ;
      RECT 0.3160 6.7365 0.3420 7.8300 ;
      RECT 0.2080 6.7365 0.2340 7.8300 ;
      RECT 0.0050 6.7365 0.0900 7.8300 ;
      RECT 8.6410 7.8165 8.7690 8.9100 ;
      RECT 8.6270 8.4820 8.7690 8.8045 ;
      RECT 8.4790 8.2090 8.5410 8.9100 ;
      RECT 8.4650 8.5185 8.5410 8.6720 ;
      RECT 8.4790 7.8165 8.5050 8.9100 ;
      RECT 8.4790 7.9375 8.5190 8.1770 ;
      RECT 8.4790 7.8165 8.5410 7.9055 ;
      RECT 8.1820 8.2670 8.3880 8.9100 ;
      RECT 8.3620 7.8165 8.3880 8.9100 ;
      RECT 8.1820 8.5440 8.4020 8.8020 ;
      RECT 8.1820 7.8165 8.2800 8.9100 ;
      RECT 7.7650 7.8165 7.8480 8.9100 ;
      RECT 7.7650 7.9050 7.8620 8.8405 ;
      RECT 16.4440 7.8165 16.5290 8.9100 ;
      RECT 16.3000 7.8165 16.3260 8.9100 ;
      RECT 16.1920 7.8165 16.2180 8.9100 ;
      RECT 16.0840 7.8165 16.1100 8.9100 ;
      RECT 15.9760 7.8165 16.0020 8.9100 ;
      RECT 15.8680 7.8165 15.8940 8.9100 ;
      RECT 15.7600 7.8165 15.7860 8.9100 ;
      RECT 15.6520 7.8165 15.6780 8.9100 ;
      RECT 15.5440 7.8165 15.5700 8.9100 ;
      RECT 15.4360 7.8165 15.4620 8.9100 ;
      RECT 15.3280 7.8165 15.3540 8.9100 ;
      RECT 15.2200 7.8165 15.2460 8.9100 ;
      RECT 15.1120 7.8165 15.1380 8.9100 ;
      RECT 15.0040 7.8165 15.0300 8.9100 ;
      RECT 14.8960 7.8165 14.9220 8.9100 ;
      RECT 14.7880 7.8165 14.8140 8.9100 ;
      RECT 14.6800 7.8165 14.7060 8.9100 ;
      RECT 14.5720 7.8165 14.5980 8.9100 ;
      RECT 14.4640 7.8165 14.4900 8.9100 ;
      RECT 14.3560 7.8165 14.3820 8.9100 ;
      RECT 14.2480 7.8165 14.2740 8.9100 ;
      RECT 14.1400 7.8165 14.1660 8.9100 ;
      RECT 14.0320 7.8165 14.0580 8.9100 ;
      RECT 13.9240 7.8165 13.9500 8.9100 ;
      RECT 13.8160 7.8165 13.8420 8.9100 ;
      RECT 13.7080 7.8165 13.7340 8.9100 ;
      RECT 13.6000 7.8165 13.6260 8.9100 ;
      RECT 13.4920 7.8165 13.5180 8.9100 ;
      RECT 13.3840 7.8165 13.4100 8.9100 ;
      RECT 13.2760 7.8165 13.3020 8.9100 ;
      RECT 13.1680 7.8165 13.1940 8.9100 ;
      RECT 13.0600 7.8165 13.0860 8.9100 ;
      RECT 12.9520 7.8165 12.9780 8.9100 ;
      RECT 12.8440 7.8165 12.8700 8.9100 ;
      RECT 12.7360 7.8165 12.7620 8.9100 ;
      RECT 12.6280 7.8165 12.6540 8.9100 ;
      RECT 12.5200 7.8165 12.5460 8.9100 ;
      RECT 12.4120 7.8165 12.4380 8.9100 ;
      RECT 12.3040 7.8165 12.3300 8.9100 ;
      RECT 12.1960 7.8165 12.2220 8.9100 ;
      RECT 12.0880 7.8165 12.1140 8.9100 ;
      RECT 11.9800 7.8165 12.0060 8.9100 ;
      RECT 11.8720 7.8165 11.8980 8.9100 ;
      RECT 11.7640 7.8165 11.7900 8.9100 ;
      RECT 11.6560 7.8165 11.6820 8.9100 ;
      RECT 11.5480 7.8165 11.5740 8.9100 ;
      RECT 11.4400 7.8165 11.4660 8.9100 ;
      RECT 11.3320 7.8165 11.3580 8.9100 ;
      RECT 11.2240 7.8165 11.2500 8.9100 ;
      RECT 11.1160 7.8165 11.1420 8.9100 ;
      RECT 11.0080 7.8165 11.0340 8.9100 ;
      RECT 10.9000 7.8165 10.9260 8.9100 ;
      RECT 10.7920 7.8165 10.8180 8.9100 ;
      RECT 10.6840 7.8165 10.7100 8.9100 ;
      RECT 10.5760 7.8165 10.6020 8.9100 ;
      RECT 10.4680 7.8165 10.4940 8.9100 ;
      RECT 10.3600 7.8165 10.3860 8.9100 ;
      RECT 10.2520 7.8165 10.2780 8.9100 ;
      RECT 10.1440 7.8165 10.1700 8.9100 ;
      RECT 10.0360 7.8165 10.0620 8.9100 ;
      RECT 9.9280 7.8165 9.9540 8.9100 ;
      RECT 9.8200 7.8165 9.8460 8.9100 ;
      RECT 9.7120 7.8165 9.7380 8.9100 ;
      RECT 9.6040 7.8165 9.6300 8.9100 ;
      RECT 9.4960 7.8165 9.5220 8.9100 ;
      RECT 9.3880 7.8165 9.4140 8.9100 ;
      RECT 9.1750 7.8165 9.2520 8.9100 ;
      RECT 7.2820 7.8165 7.3590 8.9100 ;
      RECT 7.1200 7.8165 7.1460 8.9100 ;
      RECT 7.0120 7.8165 7.0380 8.9100 ;
      RECT 6.9040 7.8165 6.9300 8.9100 ;
      RECT 6.7960 7.8165 6.8220 8.9100 ;
      RECT 6.6880 7.8165 6.7140 8.9100 ;
      RECT 6.5800 7.8165 6.6060 8.9100 ;
      RECT 6.4720 7.8165 6.4980 8.9100 ;
      RECT 6.3640 7.8165 6.3900 8.9100 ;
      RECT 6.2560 7.8165 6.2820 8.9100 ;
      RECT 6.1480 7.8165 6.1740 8.9100 ;
      RECT 6.0400 7.8165 6.0660 8.9100 ;
      RECT 5.9320 7.8165 5.9580 8.9100 ;
      RECT 5.8240 7.8165 5.8500 8.9100 ;
      RECT 5.7160 7.8165 5.7420 8.9100 ;
      RECT 5.6080 7.8165 5.6340 8.9100 ;
      RECT 5.5000 7.8165 5.5260 8.9100 ;
      RECT 5.3920 7.8165 5.4180 8.9100 ;
      RECT 5.2840 7.8165 5.3100 8.9100 ;
      RECT 5.1760 7.8165 5.2020 8.9100 ;
      RECT 5.0680 7.8165 5.0940 8.9100 ;
      RECT 4.9600 7.8165 4.9860 8.9100 ;
      RECT 4.8520 7.8165 4.8780 8.9100 ;
      RECT 4.7440 7.8165 4.7700 8.9100 ;
      RECT 4.6360 7.8165 4.6620 8.9100 ;
      RECT 4.5280 7.8165 4.5540 8.9100 ;
      RECT 4.4200 7.8165 4.4460 8.9100 ;
      RECT 4.3120 7.8165 4.3380 8.9100 ;
      RECT 4.2040 7.8165 4.2300 8.9100 ;
      RECT 4.0960 7.8165 4.1220 8.9100 ;
      RECT 3.9880 7.8165 4.0140 8.9100 ;
      RECT 3.8800 7.8165 3.9060 8.9100 ;
      RECT 3.7720 7.8165 3.7980 8.9100 ;
      RECT 3.6640 7.8165 3.6900 8.9100 ;
      RECT 3.5560 7.8165 3.5820 8.9100 ;
      RECT 3.4480 7.8165 3.4740 8.9100 ;
      RECT 3.3400 7.8165 3.3660 8.9100 ;
      RECT 3.2320 7.8165 3.2580 8.9100 ;
      RECT 3.1240 7.8165 3.1500 8.9100 ;
      RECT 3.0160 7.8165 3.0420 8.9100 ;
      RECT 2.9080 7.8165 2.9340 8.9100 ;
      RECT 2.8000 7.8165 2.8260 8.9100 ;
      RECT 2.6920 7.8165 2.7180 8.9100 ;
      RECT 2.5840 7.8165 2.6100 8.9100 ;
      RECT 2.4760 7.8165 2.5020 8.9100 ;
      RECT 2.3680 7.8165 2.3940 8.9100 ;
      RECT 2.2600 7.8165 2.2860 8.9100 ;
      RECT 2.1520 7.8165 2.1780 8.9100 ;
      RECT 2.0440 7.8165 2.0700 8.9100 ;
      RECT 1.9360 7.8165 1.9620 8.9100 ;
      RECT 1.8280 7.8165 1.8540 8.9100 ;
      RECT 1.7200 7.8165 1.7460 8.9100 ;
      RECT 1.6120 7.8165 1.6380 8.9100 ;
      RECT 1.5040 7.8165 1.5300 8.9100 ;
      RECT 1.3960 7.8165 1.4220 8.9100 ;
      RECT 1.2880 7.8165 1.3140 8.9100 ;
      RECT 1.1800 7.8165 1.2060 8.9100 ;
      RECT 1.0720 7.8165 1.0980 8.9100 ;
      RECT 0.9640 7.8165 0.9900 8.9100 ;
      RECT 0.8560 7.8165 0.8820 8.9100 ;
      RECT 0.7480 7.8165 0.7740 8.9100 ;
      RECT 0.6400 7.8165 0.6660 8.9100 ;
      RECT 0.5320 7.8165 0.5580 8.9100 ;
      RECT 0.4240 7.8165 0.4500 8.9100 ;
      RECT 0.3160 7.8165 0.3420 8.9100 ;
      RECT 0.2080 7.8165 0.2340 8.9100 ;
      RECT 0.0050 7.8165 0.0900 8.9100 ;
      RECT 8.6410 8.8965 8.7690 9.9900 ;
      RECT 8.6270 9.5620 8.7690 9.8845 ;
      RECT 8.4790 9.2890 8.5410 9.9900 ;
      RECT 8.4650 9.5985 8.5410 9.7520 ;
      RECT 8.4790 8.8965 8.5050 9.9900 ;
      RECT 8.4790 9.0175 8.5190 9.2570 ;
      RECT 8.4790 8.8965 8.5410 8.9855 ;
      RECT 8.1820 9.3470 8.3880 9.9900 ;
      RECT 8.3620 8.8965 8.3880 9.9900 ;
      RECT 8.1820 9.6240 8.4020 9.8820 ;
      RECT 8.1820 8.8965 8.2800 9.9900 ;
      RECT 7.7650 8.8965 7.8480 9.9900 ;
      RECT 7.7650 8.9850 7.8620 9.9205 ;
      RECT 16.4440 8.8965 16.5290 9.9900 ;
      RECT 16.3000 8.8965 16.3260 9.9900 ;
      RECT 16.1920 8.8965 16.2180 9.9900 ;
      RECT 16.0840 8.8965 16.1100 9.9900 ;
      RECT 15.9760 8.8965 16.0020 9.9900 ;
      RECT 15.8680 8.8965 15.8940 9.9900 ;
      RECT 15.7600 8.8965 15.7860 9.9900 ;
      RECT 15.6520 8.8965 15.6780 9.9900 ;
      RECT 15.5440 8.8965 15.5700 9.9900 ;
      RECT 15.4360 8.8965 15.4620 9.9900 ;
      RECT 15.3280 8.8965 15.3540 9.9900 ;
      RECT 15.2200 8.8965 15.2460 9.9900 ;
      RECT 15.1120 8.8965 15.1380 9.9900 ;
      RECT 15.0040 8.8965 15.0300 9.9900 ;
      RECT 14.8960 8.8965 14.9220 9.9900 ;
      RECT 14.7880 8.8965 14.8140 9.9900 ;
      RECT 14.6800 8.8965 14.7060 9.9900 ;
      RECT 14.5720 8.8965 14.5980 9.9900 ;
      RECT 14.4640 8.8965 14.4900 9.9900 ;
      RECT 14.3560 8.8965 14.3820 9.9900 ;
      RECT 14.2480 8.8965 14.2740 9.9900 ;
      RECT 14.1400 8.8965 14.1660 9.9900 ;
      RECT 14.0320 8.8965 14.0580 9.9900 ;
      RECT 13.9240 8.8965 13.9500 9.9900 ;
      RECT 13.8160 8.8965 13.8420 9.9900 ;
      RECT 13.7080 8.8965 13.7340 9.9900 ;
      RECT 13.6000 8.8965 13.6260 9.9900 ;
      RECT 13.4920 8.8965 13.5180 9.9900 ;
      RECT 13.3840 8.8965 13.4100 9.9900 ;
      RECT 13.2760 8.8965 13.3020 9.9900 ;
      RECT 13.1680 8.8965 13.1940 9.9900 ;
      RECT 13.0600 8.8965 13.0860 9.9900 ;
      RECT 12.9520 8.8965 12.9780 9.9900 ;
      RECT 12.8440 8.8965 12.8700 9.9900 ;
      RECT 12.7360 8.8965 12.7620 9.9900 ;
      RECT 12.6280 8.8965 12.6540 9.9900 ;
      RECT 12.5200 8.8965 12.5460 9.9900 ;
      RECT 12.4120 8.8965 12.4380 9.9900 ;
      RECT 12.3040 8.8965 12.3300 9.9900 ;
      RECT 12.1960 8.8965 12.2220 9.9900 ;
      RECT 12.0880 8.8965 12.1140 9.9900 ;
      RECT 11.9800 8.8965 12.0060 9.9900 ;
      RECT 11.8720 8.8965 11.8980 9.9900 ;
      RECT 11.7640 8.8965 11.7900 9.9900 ;
      RECT 11.6560 8.8965 11.6820 9.9900 ;
      RECT 11.5480 8.8965 11.5740 9.9900 ;
      RECT 11.4400 8.8965 11.4660 9.9900 ;
      RECT 11.3320 8.8965 11.3580 9.9900 ;
      RECT 11.2240 8.8965 11.2500 9.9900 ;
      RECT 11.1160 8.8965 11.1420 9.9900 ;
      RECT 11.0080 8.8965 11.0340 9.9900 ;
      RECT 10.9000 8.8965 10.9260 9.9900 ;
      RECT 10.7920 8.8965 10.8180 9.9900 ;
      RECT 10.6840 8.8965 10.7100 9.9900 ;
      RECT 10.5760 8.8965 10.6020 9.9900 ;
      RECT 10.4680 8.8965 10.4940 9.9900 ;
      RECT 10.3600 8.8965 10.3860 9.9900 ;
      RECT 10.2520 8.8965 10.2780 9.9900 ;
      RECT 10.1440 8.8965 10.1700 9.9900 ;
      RECT 10.0360 8.8965 10.0620 9.9900 ;
      RECT 9.9280 8.8965 9.9540 9.9900 ;
      RECT 9.8200 8.8965 9.8460 9.9900 ;
      RECT 9.7120 8.8965 9.7380 9.9900 ;
      RECT 9.6040 8.8965 9.6300 9.9900 ;
      RECT 9.4960 8.8965 9.5220 9.9900 ;
      RECT 9.3880 8.8965 9.4140 9.9900 ;
      RECT 9.1750 8.8965 9.2520 9.9900 ;
      RECT 7.2820 8.8965 7.3590 9.9900 ;
      RECT 7.1200 8.8965 7.1460 9.9900 ;
      RECT 7.0120 8.8965 7.0380 9.9900 ;
      RECT 6.9040 8.8965 6.9300 9.9900 ;
      RECT 6.7960 8.8965 6.8220 9.9900 ;
      RECT 6.6880 8.8965 6.7140 9.9900 ;
      RECT 6.5800 8.8965 6.6060 9.9900 ;
      RECT 6.4720 8.8965 6.4980 9.9900 ;
      RECT 6.3640 8.8965 6.3900 9.9900 ;
      RECT 6.2560 8.8965 6.2820 9.9900 ;
      RECT 6.1480 8.8965 6.1740 9.9900 ;
      RECT 6.0400 8.8965 6.0660 9.9900 ;
      RECT 5.9320 8.8965 5.9580 9.9900 ;
      RECT 5.8240 8.8965 5.8500 9.9900 ;
      RECT 5.7160 8.8965 5.7420 9.9900 ;
      RECT 5.6080 8.8965 5.6340 9.9900 ;
      RECT 5.5000 8.8965 5.5260 9.9900 ;
      RECT 5.3920 8.8965 5.4180 9.9900 ;
      RECT 5.2840 8.8965 5.3100 9.9900 ;
      RECT 5.1760 8.8965 5.2020 9.9900 ;
      RECT 5.0680 8.8965 5.0940 9.9900 ;
      RECT 4.9600 8.8965 4.9860 9.9900 ;
      RECT 4.8520 8.8965 4.8780 9.9900 ;
      RECT 4.7440 8.8965 4.7700 9.9900 ;
      RECT 4.6360 8.8965 4.6620 9.9900 ;
      RECT 4.5280 8.8965 4.5540 9.9900 ;
      RECT 4.4200 8.8965 4.4460 9.9900 ;
      RECT 4.3120 8.8965 4.3380 9.9900 ;
      RECT 4.2040 8.8965 4.2300 9.9900 ;
      RECT 4.0960 8.8965 4.1220 9.9900 ;
      RECT 3.9880 8.8965 4.0140 9.9900 ;
      RECT 3.8800 8.8965 3.9060 9.9900 ;
      RECT 3.7720 8.8965 3.7980 9.9900 ;
      RECT 3.6640 8.8965 3.6900 9.9900 ;
      RECT 3.5560 8.8965 3.5820 9.9900 ;
      RECT 3.4480 8.8965 3.4740 9.9900 ;
      RECT 3.3400 8.8965 3.3660 9.9900 ;
      RECT 3.2320 8.8965 3.2580 9.9900 ;
      RECT 3.1240 8.8965 3.1500 9.9900 ;
      RECT 3.0160 8.8965 3.0420 9.9900 ;
      RECT 2.9080 8.8965 2.9340 9.9900 ;
      RECT 2.8000 8.8965 2.8260 9.9900 ;
      RECT 2.6920 8.8965 2.7180 9.9900 ;
      RECT 2.5840 8.8965 2.6100 9.9900 ;
      RECT 2.4760 8.8965 2.5020 9.9900 ;
      RECT 2.3680 8.8965 2.3940 9.9900 ;
      RECT 2.2600 8.8965 2.2860 9.9900 ;
      RECT 2.1520 8.8965 2.1780 9.9900 ;
      RECT 2.0440 8.8965 2.0700 9.9900 ;
      RECT 1.9360 8.8965 1.9620 9.9900 ;
      RECT 1.8280 8.8965 1.8540 9.9900 ;
      RECT 1.7200 8.8965 1.7460 9.9900 ;
      RECT 1.6120 8.8965 1.6380 9.9900 ;
      RECT 1.5040 8.8965 1.5300 9.9900 ;
      RECT 1.3960 8.8965 1.4220 9.9900 ;
      RECT 1.2880 8.8965 1.3140 9.9900 ;
      RECT 1.1800 8.8965 1.2060 9.9900 ;
      RECT 1.0720 8.8965 1.0980 9.9900 ;
      RECT 0.9640 8.8965 0.9900 9.9900 ;
      RECT 0.8560 8.8965 0.8820 9.9900 ;
      RECT 0.7480 8.8965 0.7740 9.9900 ;
      RECT 0.6400 8.8965 0.6660 9.9900 ;
      RECT 0.5320 8.8965 0.5580 9.9900 ;
      RECT 0.4240 8.8965 0.4500 9.9900 ;
      RECT 0.3160 8.8965 0.3420 9.9900 ;
      RECT 0.2080 8.8965 0.2340 9.9900 ;
      RECT 0.0050 8.8965 0.0900 9.9900 ;
      RECT 8.6410 9.9765 8.7690 11.0700 ;
      RECT 8.6270 10.6420 8.7690 10.9645 ;
      RECT 8.4790 10.3690 8.5410 11.0700 ;
      RECT 8.4650 10.6785 8.5410 10.8320 ;
      RECT 8.4790 9.9765 8.5050 11.0700 ;
      RECT 8.4790 10.0975 8.5190 10.3370 ;
      RECT 8.4790 9.9765 8.5410 10.0655 ;
      RECT 8.1820 10.4270 8.3880 11.0700 ;
      RECT 8.3620 9.9765 8.3880 11.0700 ;
      RECT 8.1820 10.7040 8.4020 10.9620 ;
      RECT 8.1820 9.9765 8.2800 11.0700 ;
      RECT 7.7650 9.9765 7.8480 11.0700 ;
      RECT 7.7650 10.0650 7.8620 11.0005 ;
      RECT 16.4440 9.9765 16.5290 11.0700 ;
      RECT 16.3000 9.9765 16.3260 11.0700 ;
      RECT 16.1920 9.9765 16.2180 11.0700 ;
      RECT 16.0840 9.9765 16.1100 11.0700 ;
      RECT 15.9760 9.9765 16.0020 11.0700 ;
      RECT 15.8680 9.9765 15.8940 11.0700 ;
      RECT 15.7600 9.9765 15.7860 11.0700 ;
      RECT 15.6520 9.9765 15.6780 11.0700 ;
      RECT 15.5440 9.9765 15.5700 11.0700 ;
      RECT 15.4360 9.9765 15.4620 11.0700 ;
      RECT 15.3280 9.9765 15.3540 11.0700 ;
      RECT 15.2200 9.9765 15.2460 11.0700 ;
      RECT 15.1120 9.9765 15.1380 11.0700 ;
      RECT 15.0040 9.9765 15.0300 11.0700 ;
      RECT 14.8960 9.9765 14.9220 11.0700 ;
      RECT 14.7880 9.9765 14.8140 11.0700 ;
      RECT 14.6800 9.9765 14.7060 11.0700 ;
      RECT 14.5720 9.9765 14.5980 11.0700 ;
      RECT 14.4640 9.9765 14.4900 11.0700 ;
      RECT 14.3560 9.9765 14.3820 11.0700 ;
      RECT 14.2480 9.9765 14.2740 11.0700 ;
      RECT 14.1400 9.9765 14.1660 11.0700 ;
      RECT 14.0320 9.9765 14.0580 11.0700 ;
      RECT 13.9240 9.9765 13.9500 11.0700 ;
      RECT 13.8160 9.9765 13.8420 11.0700 ;
      RECT 13.7080 9.9765 13.7340 11.0700 ;
      RECT 13.6000 9.9765 13.6260 11.0700 ;
      RECT 13.4920 9.9765 13.5180 11.0700 ;
      RECT 13.3840 9.9765 13.4100 11.0700 ;
      RECT 13.2760 9.9765 13.3020 11.0700 ;
      RECT 13.1680 9.9765 13.1940 11.0700 ;
      RECT 13.0600 9.9765 13.0860 11.0700 ;
      RECT 12.9520 9.9765 12.9780 11.0700 ;
      RECT 12.8440 9.9765 12.8700 11.0700 ;
      RECT 12.7360 9.9765 12.7620 11.0700 ;
      RECT 12.6280 9.9765 12.6540 11.0700 ;
      RECT 12.5200 9.9765 12.5460 11.0700 ;
      RECT 12.4120 9.9765 12.4380 11.0700 ;
      RECT 12.3040 9.9765 12.3300 11.0700 ;
      RECT 12.1960 9.9765 12.2220 11.0700 ;
      RECT 12.0880 9.9765 12.1140 11.0700 ;
      RECT 11.9800 9.9765 12.0060 11.0700 ;
      RECT 11.8720 9.9765 11.8980 11.0700 ;
      RECT 11.7640 9.9765 11.7900 11.0700 ;
      RECT 11.6560 9.9765 11.6820 11.0700 ;
      RECT 11.5480 9.9765 11.5740 11.0700 ;
      RECT 11.4400 9.9765 11.4660 11.0700 ;
      RECT 11.3320 9.9765 11.3580 11.0700 ;
      RECT 11.2240 9.9765 11.2500 11.0700 ;
      RECT 11.1160 9.9765 11.1420 11.0700 ;
      RECT 11.0080 9.9765 11.0340 11.0700 ;
      RECT 10.9000 9.9765 10.9260 11.0700 ;
      RECT 10.7920 9.9765 10.8180 11.0700 ;
      RECT 10.6840 9.9765 10.7100 11.0700 ;
      RECT 10.5760 9.9765 10.6020 11.0700 ;
      RECT 10.4680 9.9765 10.4940 11.0700 ;
      RECT 10.3600 9.9765 10.3860 11.0700 ;
      RECT 10.2520 9.9765 10.2780 11.0700 ;
      RECT 10.1440 9.9765 10.1700 11.0700 ;
      RECT 10.0360 9.9765 10.0620 11.0700 ;
      RECT 9.9280 9.9765 9.9540 11.0700 ;
      RECT 9.8200 9.9765 9.8460 11.0700 ;
      RECT 9.7120 9.9765 9.7380 11.0700 ;
      RECT 9.6040 9.9765 9.6300 11.0700 ;
      RECT 9.4960 9.9765 9.5220 11.0700 ;
      RECT 9.3880 9.9765 9.4140 11.0700 ;
      RECT 9.1750 9.9765 9.2520 11.0700 ;
      RECT 7.2820 9.9765 7.3590 11.0700 ;
      RECT 7.1200 9.9765 7.1460 11.0700 ;
      RECT 7.0120 9.9765 7.0380 11.0700 ;
      RECT 6.9040 9.9765 6.9300 11.0700 ;
      RECT 6.7960 9.9765 6.8220 11.0700 ;
      RECT 6.6880 9.9765 6.7140 11.0700 ;
      RECT 6.5800 9.9765 6.6060 11.0700 ;
      RECT 6.4720 9.9765 6.4980 11.0700 ;
      RECT 6.3640 9.9765 6.3900 11.0700 ;
      RECT 6.2560 9.9765 6.2820 11.0700 ;
      RECT 6.1480 9.9765 6.1740 11.0700 ;
      RECT 6.0400 9.9765 6.0660 11.0700 ;
      RECT 5.9320 9.9765 5.9580 11.0700 ;
      RECT 5.8240 9.9765 5.8500 11.0700 ;
      RECT 5.7160 9.9765 5.7420 11.0700 ;
      RECT 5.6080 9.9765 5.6340 11.0700 ;
      RECT 5.5000 9.9765 5.5260 11.0700 ;
      RECT 5.3920 9.9765 5.4180 11.0700 ;
      RECT 5.2840 9.9765 5.3100 11.0700 ;
      RECT 5.1760 9.9765 5.2020 11.0700 ;
      RECT 5.0680 9.9765 5.0940 11.0700 ;
      RECT 4.9600 9.9765 4.9860 11.0700 ;
      RECT 4.8520 9.9765 4.8780 11.0700 ;
      RECT 4.7440 9.9765 4.7700 11.0700 ;
      RECT 4.6360 9.9765 4.6620 11.0700 ;
      RECT 4.5280 9.9765 4.5540 11.0700 ;
      RECT 4.4200 9.9765 4.4460 11.0700 ;
      RECT 4.3120 9.9765 4.3380 11.0700 ;
      RECT 4.2040 9.9765 4.2300 11.0700 ;
      RECT 4.0960 9.9765 4.1220 11.0700 ;
      RECT 3.9880 9.9765 4.0140 11.0700 ;
      RECT 3.8800 9.9765 3.9060 11.0700 ;
      RECT 3.7720 9.9765 3.7980 11.0700 ;
      RECT 3.6640 9.9765 3.6900 11.0700 ;
      RECT 3.5560 9.9765 3.5820 11.0700 ;
      RECT 3.4480 9.9765 3.4740 11.0700 ;
      RECT 3.3400 9.9765 3.3660 11.0700 ;
      RECT 3.2320 9.9765 3.2580 11.0700 ;
      RECT 3.1240 9.9765 3.1500 11.0700 ;
      RECT 3.0160 9.9765 3.0420 11.0700 ;
      RECT 2.9080 9.9765 2.9340 11.0700 ;
      RECT 2.8000 9.9765 2.8260 11.0700 ;
      RECT 2.6920 9.9765 2.7180 11.0700 ;
      RECT 2.5840 9.9765 2.6100 11.0700 ;
      RECT 2.4760 9.9765 2.5020 11.0700 ;
      RECT 2.3680 9.9765 2.3940 11.0700 ;
      RECT 2.2600 9.9765 2.2860 11.0700 ;
      RECT 2.1520 9.9765 2.1780 11.0700 ;
      RECT 2.0440 9.9765 2.0700 11.0700 ;
      RECT 1.9360 9.9765 1.9620 11.0700 ;
      RECT 1.8280 9.9765 1.8540 11.0700 ;
      RECT 1.7200 9.9765 1.7460 11.0700 ;
      RECT 1.6120 9.9765 1.6380 11.0700 ;
      RECT 1.5040 9.9765 1.5300 11.0700 ;
      RECT 1.3960 9.9765 1.4220 11.0700 ;
      RECT 1.2880 9.9765 1.3140 11.0700 ;
      RECT 1.1800 9.9765 1.2060 11.0700 ;
      RECT 1.0720 9.9765 1.0980 11.0700 ;
      RECT 0.9640 9.9765 0.9900 11.0700 ;
      RECT 0.8560 9.9765 0.8820 11.0700 ;
      RECT 0.7480 9.9765 0.7740 11.0700 ;
      RECT 0.6400 9.9765 0.6660 11.0700 ;
      RECT 0.5320 9.9765 0.5580 11.0700 ;
      RECT 0.4240 9.9765 0.4500 11.0700 ;
      RECT 0.3160 9.9765 0.3420 11.0700 ;
      RECT 0.2080 9.9765 0.2340 11.0700 ;
      RECT 0.0050 9.9765 0.0900 11.0700 ;
      RECT 0.0000 19.2495 16.5240 19.6905 ;
      RECT 16.4390 11.0370 16.5240 19.6905 ;
      RECT 9.3830 12.5410 16.3210 19.6905 ;
      RECT 10.8410 11.0370 16.3210 19.6905 ;
      RECT 7.2230 19.2420 9.3010 19.6905 ;
      RECT 7.9970 19.2105 9.3010 19.6905 ;
      RECT 0.2030 12.3460 7.1410 19.6905 ;
      RECT 6.8450 11.0370 7.1410 19.6905 ;
      RECT 0.0000 11.0370 0.0850 19.6905 ;
      RECT 7.2230 12.6490 7.8430 19.6905 ;
      RECT 7.9970 19.2060 9.2650 19.6905 ;
      RECT 8.6450 12.4420 9.2650 19.6905 ;
      RECT 8.6360 18.9490 9.2650 19.6905 ;
      RECT 8.4740 18.9490 8.5360 19.6905 ;
      RECT 7.9970 18.9490 8.3830 19.6905 ;
      RECT 9.3830 14.8300 16.3350 19.1840 ;
      RECT 0.1890 14.8300 7.1410 19.1840 ;
      RECT 9.3690 14.8300 16.3350 19.1795 ;
      RECT 0.1890 14.8300 7.1550 19.1795 ;
      RECT 7.2090 14.8300 7.8430 19.1785 ;
      RECT 8.1770 11.7220 8.3470 19.6905 ;
      RECT 8.2850 11.0370 8.3470 19.6905 ;
      RECT 7.4930 11.4580 7.8790 18.8020 ;
      RECT 7.2090 18.7570 7.8930 18.7940 ;
      RECT 8.6310 17.6830 9.2650 18.7910 ;
      RECT 8.1630 18.4930 8.3470 18.7190 ;
      RECT 8.1770 17.9170 8.3610 18.1790 ;
      RECT 7.2090 17.7190 7.8930 18.1790 ;
      RECT 8.1630 17.1790 8.3470 17.6390 ;
      RECT 8.6310 15.1450 9.2650 17.4770 ;
      RECT 7.2090 15.7930 7.8930 16.9370 ;
      RECT 8.1770 15.5230 8.3610 16.8290 ;
      RECT 8.1630 16.0990 8.3610 16.5590 ;
      RECT 8.1630 12.8590 8.3470 16.0190 ;
      RECT 8.1630 12.8590 8.3610 15.4790 ;
      RECT 7.2090 15.2530 7.8930 15.4790 ;
      RECT 8.6450 12.4420 9.3010 14.7980 ;
      RECT 8.6310 12.3190 9.2470 14.1050 ;
      RECT 7.2230 13.2910 7.8930 13.6610 ;
      RECT 8.1770 12.5890 8.3610 12.7790 ;
      RECT 7.2770 12.5530 7.8930 12.7430 ;
      RECT 8.1630 12.4450 8.3470 12.5810 ;
      RECT 7.2770 11.8030 7.8790 18.8020 ;
      RECT 8.1770 12.3190 8.3610 12.5450 ;
      RECT 9.5450 12.3490 16.3210 19.6905 ;
      RECT 10.6250 12.3460 16.3210 19.6905 ;
      RECT 9.3830 11.0370 9.4630 19.6905 ;
      RECT 7.2230 11.7220 7.4110 12.5360 ;
      RECT 9.3830 11.0370 9.6790 12.4400 ;
      RECT 9.3830 12.1540 10.5430 12.4400 ;
      RECT 10.6250 11.0370 10.7590 19.6905 ;
      RECT 5.9810 11.9650 6.7630 19.6905 ;
      RECT 0.2030 11.0370 5.8990 19.6905 ;
      RECT 8.6450 11.8030 9.2470 19.6905 ;
      RECT 8.6810 11.2135 9.3010 12.2870 ;
      RECT 9.3830 12.1540 10.7590 12.2480 ;
      RECT 10.4090 11.0370 16.3210 12.2450 ;
      RECT 6.6290 11.0370 7.1410 12.2450 ;
      RECT 8.1630 12.1750 8.3610 12.2390 ;
      RECT 8.1630 12.0490 8.3470 12.2390 ;
      RECT 10.1930 11.7700 16.3210 12.2450 ;
      RECT 9.3830 11.8030 10.1110 12.4400 ;
      RECT 8.1770 11.7790 8.3610 12.0410 ;
      RECT 0.2030 11.7700 6.5470 12.2450 ;
      RECT 6.4130 11.0370 6.5470 19.6905 ;
      RECT 9.9770 11.0370 10.3270 11.9090 ;
      RECT 9.3830 11.7220 9.8950 12.4400 ;
      RECT 9.7610 11.0370 9.8950 19.6905 ;
      RECT 6.1970 11.7220 6.5470 19.6905 ;
      RECT 0.2030 11.0370 6.1150 12.2450 ;
      RECT 8.1770 11.0370 8.2030 19.6905 ;
      RECT 7.3130 11.0370 7.4110 19.6905 ;
      RECT 6.1970 11.0370 6.3310 19.6905 ;
      RECT 9.7610 11.0370 10.3270 11.6720 ;
      RECT 8.6450 11.0370 9.2470 11.6720 ;
      RECT 7.3130 11.0370 7.8430 11.6720 ;
      RECT 6.4130 11.0370 7.1410 11.6720 ;
      RECT 9.7610 11.0370 16.3210 11.6690 ;
      RECT 0.2030 11.0370 6.3310 11.6690 ;
      RECT 8.6310 11.5090 9.3010 11.6630 ;
      RECT 9.3830 11.0370 16.3210 11.4050 ;
      RECT 8.1770 11.0370 8.3470 11.4050 ;
      RECT 7.2230 11.0370 7.8430 11.4050 ;
      RECT 0.2030 11.0370 7.1410 11.4050 ;
      RECT 7.9970 11.0370 8.3470 11.3020 ;
      RECT 8.6360 11.0370 9.2470 11.2020 ;
      RECT 7.9970 11.0370 8.3830 11.2020 ;
      RECT 9.7650 11.0105 9.7830 19.6905 ;
      RECT 9.6570 11.0105 9.6750 19.6905 ;
      RECT 6.8490 11.0230 6.8670 19.6905 ;
      RECT 6.7410 11.0230 6.7590 19.6905 ;
      RECT 6.6330 11.0230 6.6510 19.6905 ;
      RECT 6.5250 11.0230 6.5430 19.6905 ;
      RECT 6.4170 11.0105 6.4350 19.6905 ;
      RECT 6.3090 11.0105 6.3270 19.6905 ;
      RECT 6.2010 11.0230 6.2190 19.6905 ;
      RECT 6.0930 11.0230 6.1110 19.6905 ;
      RECT 5.9850 11.0230 6.0030 19.6905 ;
      RECT 5.8770 11.0230 5.8950 19.6905 ;
      RECT 8.4740 11.0370 8.5360 11.2020 ;
        RECT 8.6410 19.1835 8.7690 20.2770 ;
        RECT 8.6270 19.8490 8.7690 20.1715 ;
        RECT 8.4790 19.5760 8.5410 20.2770 ;
        RECT 8.4650 19.8855 8.5410 20.0390 ;
        RECT 8.4790 19.1835 8.5050 20.2770 ;
        RECT 8.4790 19.3045 8.5190 19.5440 ;
        RECT 8.4790 19.1835 8.5410 19.2725 ;
        RECT 8.1820 19.6340 8.3880 20.2770 ;
        RECT 8.3620 19.1835 8.3880 20.2770 ;
        RECT 8.1820 19.9110 8.4020 20.1690 ;
        RECT 8.1820 19.1835 8.2800 20.2770 ;
        RECT 7.7650 19.1835 7.8480 20.2770 ;
        RECT 7.7650 19.2720 7.8620 20.2075 ;
        RECT 16.4440 19.1835 16.5290 20.2770 ;
        RECT 16.3000 19.1835 16.3260 20.2770 ;
        RECT 16.1920 19.1835 16.2180 20.2770 ;
        RECT 16.0840 19.1835 16.1100 20.2770 ;
        RECT 15.9760 19.1835 16.0020 20.2770 ;
        RECT 15.8680 19.1835 15.8940 20.2770 ;
        RECT 15.7600 19.1835 15.7860 20.2770 ;
        RECT 15.6520 19.1835 15.6780 20.2770 ;
        RECT 15.5440 19.1835 15.5700 20.2770 ;
        RECT 15.4360 19.1835 15.4620 20.2770 ;
        RECT 15.3280 19.1835 15.3540 20.2770 ;
        RECT 15.2200 19.1835 15.2460 20.2770 ;
        RECT 15.1120 19.1835 15.1380 20.2770 ;
        RECT 15.0040 19.1835 15.0300 20.2770 ;
        RECT 14.8960 19.1835 14.9220 20.2770 ;
        RECT 14.7880 19.1835 14.8140 20.2770 ;
        RECT 14.6800 19.1835 14.7060 20.2770 ;
        RECT 14.5720 19.1835 14.5980 20.2770 ;
        RECT 14.4640 19.1835 14.4900 20.2770 ;
        RECT 14.3560 19.1835 14.3820 20.2770 ;
        RECT 14.2480 19.1835 14.2740 20.2770 ;
        RECT 14.1400 19.1835 14.1660 20.2770 ;
        RECT 14.0320 19.1835 14.0580 20.2770 ;
        RECT 13.9240 19.1835 13.9500 20.2770 ;
        RECT 13.8160 19.1835 13.8420 20.2770 ;
        RECT 13.7080 19.1835 13.7340 20.2770 ;
        RECT 13.6000 19.1835 13.6260 20.2770 ;
        RECT 13.4920 19.1835 13.5180 20.2770 ;
        RECT 13.3840 19.1835 13.4100 20.2770 ;
        RECT 13.2760 19.1835 13.3020 20.2770 ;
        RECT 13.1680 19.1835 13.1940 20.2770 ;
        RECT 13.0600 19.1835 13.0860 20.2770 ;
        RECT 12.9520 19.1835 12.9780 20.2770 ;
        RECT 12.8440 19.1835 12.8700 20.2770 ;
        RECT 12.7360 19.1835 12.7620 20.2770 ;
        RECT 12.6280 19.1835 12.6540 20.2770 ;
        RECT 12.5200 19.1835 12.5460 20.2770 ;
        RECT 12.4120 19.1835 12.4380 20.2770 ;
        RECT 12.3040 19.1835 12.3300 20.2770 ;
        RECT 12.1960 19.1835 12.2220 20.2770 ;
        RECT 12.0880 19.1835 12.1140 20.2770 ;
        RECT 11.9800 19.1835 12.0060 20.2770 ;
        RECT 11.8720 19.1835 11.8980 20.2770 ;
        RECT 11.7640 19.1835 11.7900 20.2770 ;
        RECT 11.6560 19.1835 11.6820 20.2770 ;
        RECT 11.5480 19.1835 11.5740 20.2770 ;
        RECT 11.4400 19.1835 11.4660 20.2770 ;
        RECT 11.3320 19.1835 11.3580 20.2770 ;
        RECT 11.2240 19.1835 11.2500 20.2770 ;
        RECT 11.1160 19.1835 11.1420 20.2770 ;
        RECT 11.0080 19.1835 11.0340 20.2770 ;
        RECT 10.9000 19.1835 10.9260 20.2770 ;
        RECT 10.7920 19.1835 10.8180 20.2770 ;
        RECT 10.6840 19.1835 10.7100 20.2770 ;
        RECT 10.5760 19.1835 10.6020 20.2770 ;
        RECT 10.4680 19.1835 10.4940 20.2770 ;
        RECT 10.3600 19.1835 10.3860 20.2770 ;
        RECT 10.2520 19.1835 10.2780 20.2770 ;
        RECT 10.1440 19.1835 10.1700 20.2770 ;
        RECT 10.0360 19.1835 10.0620 20.2770 ;
        RECT 9.9280 19.1835 9.9540 20.2770 ;
        RECT 9.8200 19.1835 9.8460 20.2770 ;
        RECT 9.7120 19.1835 9.7380 20.2770 ;
        RECT 9.6040 19.1835 9.6300 20.2770 ;
        RECT 9.4960 19.1835 9.5220 20.2770 ;
        RECT 9.3880 19.1835 9.4140 20.2770 ;
        RECT 9.1750 19.1835 9.2520 20.2770 ;
        RECT 7.2820 19.1835 7.3590 20.2770 ;
        RECT 7.1200 19.1835 7.1460 20.2770 ;
        RECT 7.0120 19.1835 7.0380 20.2770 ;
        RECT 6.9040 19.1835 6.9300 20.2770 ;
        RECT 6.7960 19.1835 6.8220 20.2770 ;
        RECT 6.6880 19.1835 6.7140 20.2770 ;
        RECT 6.5800 19.1835 6.6060 20.2770 ;
        RECT 6.4720 19.1835 6.4980 20.2770 ;
        RECT 6.3640 19.1835 6.3900 20.2770 ;
        RECT 6.2560 19.1835 6.2820 20.2770 ;
        RECT 6.1480 19.1835 6.1740 20.2770 ;
        RECT 6.0400 19.1835 6.0660 20.2770 ;
        RECT 5.9320 19.1835 5.9580 20.2770 ;
        RECT 5.8240 19.1835 5.8500 20.2770 ;
        RECT 5.7160 19.1835 5.7420 20.2770 ;
        RECT 5.6080 19.1835 5.6340 20.2770 ;
        RECT 5.5000 19.1835 5.5260 20.2770 ;
        RECT 5.3920 19.1835 5.4180 20.2770 ;
        RECT 5.2840 19.1835 5.3100 20.2770 ;
        RECT 5.1760 19.1835 5.2020 20.2770 ;
        RECT 5.0680 19.1835 5.0940 20.2770 ;
        RECT 4.9600 19.1835 4.9860 20.2770 ;
        RECT 4.8520 19.1835 4.8780 20.2770 ;
        RECT 4.7440 19.1835 4.7700 20.2770 ;
        RECT 4.6360 19.1835 4.6620 20.2770 ;
        RECT 4.5280 19.1835 4.5540 20.2770 ;
        RECT 4.4200 19.1835 4.4460 20.2770 ;
        RECT 4.3120 19.1835 4.3380 20.2770 ;
        RECT 4.2040 19.1835 4.2300 20.2770 ;
        RECT 4.0960 19.1835 4.1220 20.2770 ;
        RECT 3.9880 19.1835 4.0140 20.2770 ;
        RECT 3.8800 19.1835 3.9060 20.2770 ;
        RECT 3.7720 19.1835 3.7980 20.2770 ;
        RECT 3.6640 19.1835 3.6900 20.2770 ;
        RECT 3.5560 19.1835 3.5820 20.2770 ;
        RECT 3.4480 19.1835 3.4740 20.2770 ;
        RECT 3.3400 19.1835 3.3660 20.2770 ;
        RECT 3.2320 19.1835 3.2580 20.2770 ;
        RECT 3.1240 19.1835 3.1500 20.2770 ;
        RECT 3.0160 19.1835 3.0420 20.2770 ;
        RECT 2.9080 19.1835 2.9340 20.2770 ;
        RECT 2.8000 19.1835 2.8260 20.2770 ;
        RECT 2.6920 19.1835 2.7180 20.2770 ;
        RECT 2.5840 19.1835 2.6100 20.2770 ;
        RECT 2.4760 19.1835 2.5020 20.2770 ;
        RECT 2.3680 19.1835 2.3940 20.2770 ;
        RECT 2.2600 19.1835 2.2860 20.2770 ;
        RECT 2.1520 19.1835 2.1780 20.2770 ;
        RECT 2.0440 19.1835 2.0700 20.2770 ;
        RECT 1.9360 19.1835 1.9620 20.2770 ;
        RECT 1.8280 19.1835 1.8540 20.2770 ;
        RECT 1.7200 19.1835 1.7460 20.2770 ;
        RECT 1.6120 19.1835 1.6380 20.2770 ;
        RECT 1.5040 19.1835 1.5300 20.2770 ;
        RECT 1.3960 19.1835 1.4220 20.2770 ;
        RECT 1.2880 19.1835 1.3140 20.2770 ;
        RECT 1.1800 19.1835 1.2060 20.2770 ;
        RECT 1.0720 19.1835 1.0980 20.2770 ;
        RECT 0.9640 19.1835 0.9900 20.2770 ;
        RECT 0.8560 19.1835 0.8820 20.2770 ;
        RECT 0.7480 19.1835 0.7740 20.2770 ;
        RECT 0.6400 19.1835 0.6660 20.2770 ;
        RECT 0.5320 19.1835 0.5580 20.2770 ;
        RECT 0.4240 19.1835 0.4500 20.2770 ;
        RECT 0.3160 19.1835 0.3420 20.2770 ;
        RECT 0.2080 19.1835 0.2340 20.2770 ;
        RECT 0.0050 19.1835 0.0900 20.2770 ;
        RECT 8.6410 20.2635 8.7690 21.3570 ;
        RECT 8.6270 20.9290 8.7690 21.2515 ;
        RECT 8.4790 20.6560 8.5410 21.3570 ;
        RECT 8.4650 20.9655 8.5410 21.1190 ;
        RECT 8.4790 20.2635 8.5050 21.3570 ;
        RECT 8.4790 20.3845 8.5190 20.6240 ;
        RECT 8.4790 20.2635 8.5410 20.3525 ;
        RECT 8.1820 20.7140 8.3880 21.3570 ;
        RECT 8.3620 20.2635 8.3880 21.3570 ;
        RECT 8.1820 20.9910 8.4020 21.2490 ;
        RECT 8.1820 20.2635 8.2800 21.3570 ;
        RECT 7.7650 20.2635 7.8480 21.3570 ;
        RECT 7.7650 20.3520 7.8620 21.2875 ;
        RECT 16.4440 20.2635 16.5290 21.3570 ;
        RECT 16.3000 20.2635 16.3260 21.3570 ;
        RECT 16.1920 20.2635 16.2180 21.3570 ;
        RECT 16.0840 20.2635 16.1100 21.3570 ;
        RECT 15.9760 20.2635 16.0020 21.3570 ;
        RECT 15.8680 20.2635 15.8940 21.3570 ;
        RECT 15.7600 20.2635 15.7860 21.3570 ;
        RECT 15.6520 20.2635 15.6780 21.3570 ;
        RECT 15.5440 20.2635 15.5700 21.3570 ;
        RECT 15.4360 20.2635 15.4620 21.3570 ;
        RECT 15.3280 20.2635 15.3540 21.3570 ;
        RECT 15.2200 20.2635 15.2460 21.3570 ;
        RECT 15.1120 20.2635 15.1380 21.3570 ;
        RECT 15.0040 20.2635 15.0300 21.3570 ;
        RECT 14.8960 20.2635 14.9220 21.3570 ;
        RECT 14.7880 20.2635 14.8140 21.3570 ;
        RECT 14.6800 20.2635 14.7060 21.3570 ;
        RECT 14.5720 20.2635 14.5980 21.3570 ;
        RECT 14.4640 20.2635 14.4900 21.3570 ;
        RECT 14.3560 20.2635 14.3820 21.3570 ;
        RECT 14.2480 20.2635 14.2740 21.3570 ;
        RECT 14.1400 20.2635 14.1660 21.3570 ;
        RECT 14.0320 20.2635 14.0580 21.3570 ;
        RECT 13.9240 20.2635 13.9500 21.3570 ;
        RECT 13.8160 20.2635 13.8420 21.3570 ;
        RECT 13.7080 20.2635 13.7340 21.3570 ;
        RECT 13.6000 20.2635 13.6260 21.3570 ;
        RECT 13.4920 20.2635 13.5180 21.3570 ;
        RECT 13.3840 20.2635 13.4100 21.3570 ;
        RECT 13.2760 20.2635 13.3020 21.3570 ;
        RECT 13.1680 20.2635 13.1940 21.3570 ;
        RECT 13.0600 20.2635 13.0860 21.3570 ;
        RECT 12.9520 20.2635 12.9780 21.3570 ;
        RECT 12.8440 20.2635 12.8700 21.3570 ;
        RECT 12.7360 20.2635 12.7620 21.3570 ;
        RECT 12.6280 20.2635 12.6540 21.3570 ;
        RECT 12.5200 20.2635 12.5460 21.3570 ;
        RECT 12.4120 20.2635 12.4380 21.3570 ;
        RECT 12.3040 20.2635 12.3300 21.3570 ;
        RECT 12.1960 20.2635 12.2220 21.3570 ;
        RECT 12.0880 20.2635 12.1140 21.3570 ;
        RECT 11.9800 20.2635 12.0060 21.3570 ;
        RECT 11.8720 20.2635 11.8980 21.3570 ;
        RECT 11.7640 20.2635 11.7900 21.3570 ;
        RECT 11.6560 20.2635 11.6820 21.3570 ;
        RECT 11.5480 20.2635 11.5740 21.3570 ;
        RECT 11.4400 20.2635 11.4660 21.3570 ;
        RECT 11.3320 20.2635 11.3580 21.3570 ;
        RECT 11.2240 20.2635 11.2500 21.3570 ;
        RECT 11.1160 20.2635 11.1420 21.3570 ;
        RECT 11.0080 20.2635 11.0340 21.3570 ;
        RECT 10.9000 20.2635 10.9260 21.3570 ;
        RECT 10.7920 20.2635 10.8180 21.3570 ;
        RECT 10.6840 20.2635 10.7100 21.3570 ;
        RECT 10.5760 20.2635 10.6020 21.3570 ;
        RECT 10.4680 20.2635 10.4940 21.3570 ;
        RECT 10.3600 20.2635 10.3860 21.3570 ;
        RECT 10.2520 20.2635 10.2780 21.3570 ;
        RECT 10.1440 20.2635 10.1700 21.3570 ;
        RECT 10.0360 20.2635 10.0620 21.3570 ;
        RECT 9.9280 20.2635 9.9540 21.3570 ;
        RECT 9.8200 20.2635 9.8460 21.3570 ;
        RECT 9.7120 20.2635 9.7380 21.3570 ;
        RECT 9.6040 20.2635 9.6300 21.3570 ;
        RECT 9.4960 20.2635 9.5220 21.3570 ;
        RECT 9.3880 20.2635 9.4140 21.3570 ;
        RECT 9.1750 20.2635 9.2520 21.3570 ;
        RECT 7.2820 20.2635 7.3590 21.3570 ;
        RECT 7.1200 20.2635 7.1460 21.3570 ;
        RECT 7.0120 20.2635 7.0380 21.3570 ;
        RECT 6.9040 20.2635 6.9300 21.3570 ;
        RECT 6.7960 20.2635 6.8220 21.3570 ;
        RECT 6.6880 20.2635 6.7140 21.3570 ;
        RECT 6.5800 20.2635 6.6060 21.3570 ;
        RECT 6.4720 20.2635 6.4980 21.3570 ;
        RECT 6.3640 20.2635 6.3900 21.3570 ;
        RECT 6.2560 20.2635 6.2820 21.3570 ;
        RECT 6.1480 20.2635 6.1740 21.3570 ;
        RECT 6.0400 20.2635 6.0660 21.3570 ;
        RECT 5.9320 20.2635 5.9580 21.3570 ;
        RECT 5.8240 20.2635 5.8500 21.3570 ;
        RECT 5.7160 20.2635 5.7420 21.3570 ;
        RECT 5.6080 20.2635 5.6340 21.3570 ;
        RECT 5.5000 20.2635 5.5260 21.3570 ;
        RECT 5.3920 20.2635 5.4180 21.3570 ;
        RECT 5.2840 20.2635 5.3100 21.3570 ;
        RECT 5.1760 20.2635 5.2020 21.3570 ;
        RECT 5.0680 20.2635 5.0940 21.3570 ;
        RECT 4.9600 20.2635 4.9860 21.3570 ;
        RECT 4.8520 20.2635 4.8780 21.3570 ;
        RECT 4.7440 20.2635 4.7700 21.3570 ;
        RECT 4.6360 20.2635 4.6620 21.3570 ;
        RECT 4.5280 20.2635 4.5540 21.3570 ;
        RECT 4.4200 20.2635 4.4460 21.3570 ;
        RECT 4.3120 20.2635 4.3380 21.3570 ;
        RECT 4.2040 20.2635 4.2300 21.3570 ;
        RECT 4.0960 20.2635 4.1220 21.3570 ;
        RECT 3.9880 20.2635 4.0140 21.3570 ;
        RECT 3.8800 20.2635 3.9060 21.3570 ;
        RECT 3.7720 20.2635 3.7980 21.3570 ;
        RECT 3.6640 20.2635 3.6900 21.3570 ;
        RECT 3.5560 20.2635 3.5820 21.3570 ;
        RECT 3.4480 20.2635 3.4740 21.3570 ;
        RECT 3.3400 20.2635 3.3660 21.3570 ;
        RECT 3.2320 20.2635 3.2580 21.3570 ;
        RECT 3.1240 20.2635 3.1500 21.3570 ;
        RECT 3.0160 20.2635 3.0420 21.3570 ;
        RECT 2.9080 20.2635 2.9340 21.3570 ;
        RECT 2.8000 20.2635 2.8260 21.3570 ;
        RECT 2.6920 20.2635 2.7180 21.3570 ;
        RECT 2.5840 20.2635 2.6100 21.3570 ;
        RECT 2.4760 20.2635 2.5020 21.3570 ;
        RECT 2.3680 20.2635 2.3940 21.3570 ;
        RECT 2.2600 20.2635 2.2860 21.3570 ;
        RECT 2.1520 20.2635 2.1780 21.3570 ;
        RECT 2.0440 20.2635 2.0700 21.3570 ;
        RECT 1.9360 20.2635 1.9620 21.3570 ;
        RECT 1.8280 20.2635 1.8540 21.3570 ;
        RECT 1.7200 20.2635 1.7460 21.3570 ;
        RECT 1.6120 20.2635 1.6380 21.3570 ;
        RECT 1.5040 20.2635 1.5300 21.3570 ;
        RECT 1.3960 20.2635 1.4220 21.3570 ;
        RECT 1.2880 20.2635 1.3140 21.3570 ;
        RECT 1.1800 20.2635 1.2060 21.3570 ;
        RECT 1.0720 20.2635 1.0980 21.3570 ;
        RECT 0.9640 20.2635 0.9900 21.3570 ;
        RECT 0.8560 20.2635 0.8820 21.3570 ;
        RECT 0.7480 20.2635 0.7740 21.3570 ;
        RECT 0.6400 20.2635 0.6660 21.3570 ;
        RECT 0.5320 20.2635 0.5580 21.3570 ;
        RECT 0.4240 20.2635 0.4500 21.3570 ;
        RECT 0.3160 20.2635 0.3420 21.3570 ;
        RECT 0.2080 20.2635 0.2340 21.3570 ;
        RECT 0.0050 20.2635 0.0900 21.3570 ;
        RECT 8.6410 21.3435 8.7690 22.4370 ;
        RECT 8.6270 22.0090 8.7690 22.3315 ;
        RECT 8.4790 21.7360 8.5410 22.4370 ;
        RECT 8.4650 22.0455 8.5410 22.1990 ;
        RECT 8.4790 21.3435 8.5050 22.4370 ;
        RECT 8.4790 21.4645 8.5190 21.7040 ;
        RECT 8.4790 21.3435 8.5410 21.4325 ;
        RECT 8.1820 21.7940 8.3880 22.4370 ;
        RECT 8.3620 21.3435 8.3880 22.4370 ;
        RECT 8.1820 22.0710 8.4020 22.3290 ;
        RECT 8.1820 21.3435 8.2800 22.4370 ;
        RECT 7.7650 21.3435 7.8480 22.4370 ;
        RECT 7.7650 21.4320 7.8620 22.3675 ;
        RECT 16.4440 21.3435 16.5290 22.4370 ;
        RECT 16.3000 21.3435 16.3260 22.4370 ;
        RECT 16.1920 21.3435 16.2180 22.4370 ;
        RECT 16.0840 21.3435 16.1100 22.4370 ;
        RECT 15.9760 21.3435 16.0020 22.4370 ;
        RECT 15.8680 21.3435 15.8940 22.4370 ;
        RECT 15.7600 21.3435 15.7860 22.4370 ;
        RECT 15.6520 21.3435 15.6780 22.4370 ;
        RECT 15.5440 21.3435 15.5700 22.4370 ;
        RECT 15.4360 21.3435 15.4620 22.4370 ;
        RECT 15.3280 21.3435 15.3540 22.4370 ;
        RECT 15.2200 21.3435 15.2460 22.4370 ;
        RECT 15.1120 21.3435 15.1380 22.4370 ;
        RECT 15.0040 21.3435 15.0300 22.4370 ;
        RECT 14.8960 21.3435 14.9220 22.4370 ;
        RECT 14.7880 21.3435 14.8140 22.4370 ;
        RECT 14.6800 21.3435 14.7060 22.4370 ;
        RECT 14.5720 21.3435 14.5980 22.4370 ;
        RECT 14.4640 21.3435 14.4900 22.4370 ;
        RECT 14.3560 21.3435 14.3820 22.4370 ;
        RECT 14.2480 21.3435 14.2740 22.4370 ;
        RECT 14.1400 21.3435 14.1660 22.4370 ;
        RECT 14.0320 21.3435 14.0580 22.4370 ;
        RECT 13.9240 21.3435 13.9500 22.4370 ;
        RECT 13.8160 21.3435 13.8420 22.4370 ;
        RECT 13.7080 21.3435 13.7340 22.4370 ;
        RECT 13.6000 21.3435 13.6260 22.4370 ;
        RECT 13.4920 21.3435 13.5180 22.4370 ;
        RECT 13.3840 21.3435 13.4100 22.4370 ;
        RECT 13.2760 21.3435 13.3020 22.4370 ;
        RECT 13.1680 21.3435 13.1940 22.4370 ;
        RECT 13.0600 21.3435 13.0860 22.4370 ;
        RECT 12.9520 21.3435 12.9780 22.4370 ;
        RECT 12.8440 21.3435 12.8700 22.4370 ;
        RECT 12.7360 21.3435 12.7620 22.4370 ;
        RECT 12.6280 21.3435 12.6540 22.4370 ;
        RECT 12.5200 21.3435 12.5460 22.4370 ;
        RECT 12.4120 21.3435 12.4380 22.4370 ;
        RECT 12.3040 21.3435 12.3300 22.4370 ;
        RECT 12.1960 21.3435 12.2220 22.4370 ;
        RECT 12.0880 21.3435 12.1140 22.4370 ;
        RECT 11.9800 21.3435 12.0060 22.4370 ;
        RECT 11.8720 21.3435 11.8980 22.4370 ;
        RECT 11.7640 21.3435 11.7900 22.4370 ;
        RECT 11.6560 21.3435 11.6820 22.4370 ;
        RECT 11.5480 21.3435 11.5740 22.4370 ;
        RECT 11.4400 21.3435 11.4660 22.4370 ;
        RECT 11.3320 21.3435 11.3580 22.4370 ;
        RECT 11.2240 21.3435 11.2500 22.4370 ;
        RECT 11.1160 21.3435 11.1420 22.4370 ;
        RECT 11.0080 21.3435 11.0340 22.4370 ;
        RECT 10.9000 21.3435 10.9260 22.4370 ;
        RECT 10.7920 21.3435 10.8180 22.4370 ;
        RECT 10.6840 21.3435 10.7100 22.4370 ;
        RECT 10.5760 21.3435 10.6020 22.4370 ;
        RECT 10.4680 21.3435 10.4940 22.4370 ;
        RECT 10.3600 21.3435 10.3860 22.4370 ;
        RECT 10.2520 21.3435 10.2780 22.4370 ;
        RECT 10.1440 21.3435 10.1700 22.4370 ;
        RECT 10.0360 21.3435 10.0620 22.4370 ;
        RECT 9.9280 21.3435 9.9540 22.4370 ;
        RECT 9.8200 21.3435 9.8460 22.4370 ;
        RECT 9.7120 21.3435 9.7380 22.4370 ;
        RECT 9.6040 21.3435 9.6300 22.4370 ;
        RECT 9.4960 21.3435 9.5220 22.4370 ;
        RECT 9.3880 21.3435 9.4140 22.4370 ;
        RECT 9.1750 21.3435 9.2520 22.4370 ;
        RECT 7.2820 21.3435 7.3590 22.4370 ;
        RECT 7.1200 21.3435 7.1460 22.4370 ;
        RECT 7.0120 21.3435 7.0380 22.4370 ;
        RECT 6.9040 21.3435 6.9300 22.4370 ;
        RECT 6.7960 21.3435 6.8220 22.4370 ;
        RECT 6.6880 21.3435 6.7140 22.4370 ;
        RECT 6.5800 21.3435 6.6060 22.4370 ;
        RECT 6.4720 21.3435 6.4980 22.4370 ;
        RECT 6.3640 21.3435 6.3900 22.4370 ;
        RECT 6.2560 21.3435 6.2820 22.4370 ;
        RECT 6.1480 21.3435 6.1740 22.4370 ;
        RECT 6.0400 21.3435 6.0660 22.4370 ;
        RECT 5.9320 21.3435 5.9580 22.4370 ;
        RECT 5.8240 21.3435 5.8500 22.4370 ;
        RECT 5.7160 21.3435 5.7420 22.4370 ;
        RECT 5.6080 21.3435 5.6340 22.4370 ;
        RECT 5.5000 21.3435 5.5260 22.4370 ;
        RECT 5.3920 21.3435 5.4180 22.4370 ;
        RECT 5.2840 21.3435 5.3100 22.4370 ;
        RECT 5.1760 21.3435 5.2020 22.4370 ;
        RECT 5.0680 21.3435 5.0940 22.4370 ;
        RECT 4.9600 21.3435 4.9860 22.4370 ;
        RECT 4.8520 21.3435 4.8780 22.4370 ;
        RECT 4.7440 21.3435 4.7700 22.4370 ;
        RECT 4.6360 21.3435 4.6620 22.4370 ;
        RECT 4.5280 21.3435 4.5540 22.4370 ;
        RECT 4.4200 21.3435 4.4460 22.4370 ;
        RECT 4.3120 21.3435 4.3380 22.4370 ;
        RECT 4.2040 21.3435 4.2300 22.4370 ;
        RECT 4.0960 21.3435 4.1220 22.4370 ;
        RECT 3.9880 21.3435 4.0140 22.4370 ;
        RECT 3.8800 21.3435 3.9060 22.4370 ;
        RECT 3.7720 21.3435 3.7980 22.4370 ;
        RECT 3.6640 21.3435 3.6900 22.4370 ;
        RECT 3.5560 21.3435 3.5820 22.4370 ;
        RECT 3.4480 21.3435 3.4740 22.4370 ;
        RECT 3.3400 21.3435 3.3660 22.4370 ;
        RECT 3.2320 21.3435 3.2580 22.4370 ;
        RECT 3.1240 21.3435 3.1500 22.4370 ;
        RECT 3.0160 21.3435 3.0420 22.4370 ;
        RECT 2.9080 21.3435 2.9340 22.4370 ;
        RECT 2.8000 21.3435 2.8260 22.4370 ;
        RECT 2.6920 21.3435 2.7180 22.4370 ;
        RECT 2.5840 21.3435 2.6100 22.4370 ;
        RECT 2.4760 21.3435 2.5020 22.4370 ;
        RECT 2.3680 21.3435 2.3940 22.4370 ;
        RECT 2.2600 21.3435 2.2860 22.4370 ;
        RECT 2.1520 21.3435 2.1780 22.4370 ;
        RECT 2.0440 21.3435 2.0700 22.4370 ;
        RECT 1.9360 21.3435 1.9620 22.4370 ;
        RECT 1.8280 21.3435 1.8540 22.4370 ;
        RECT 1.7200 21.3435 1.7460 22.4370 ;
        RECT 1.6120 21.3435 1.6380 22.4370 ;
        RECT 1.5040 21.3435 1.5300 22.4370 ;
        RECT 1.3960 21.3435 1.4220 22.4370 ;
        RECT 1.2880 21.3435 1.3140 22.4370 ;
        RECT 1.1800 21.3435 1.2060 22.4370 ;
        RECT 1.0720 21.3435 1.0980 22.4370 ;
        RECT 0.9640 21.3435 0.9900 22.4370 ;
        RECT 0.8560 21.3435 0.8820 22.4370 ;
        RECT 0.7480 21.3435 0.7740 22.4370 ;
        RECT 0.6400 21.3435 0.6660 22.4370 ;
        RECT 0.5320 21.3435 0.5580 22.4370 ;
        RECT 0.4240 21.3435 0.4500 22.4370 ;
        RECT 0.3160 21.3435 0.3420 22.4370 ;
        RECT 0.2080 21.3435 0.2340 22.4370 ;
        RECT 0.0050 21.3435 0.0900 22.4370 ;
        RECT 8.6410 22.4235 8.7690 23.5170 ;
        RECT 8.6270 23.0890 8.7690 23.4115 ;
        RECT 8.4790 22.8160 8.5410 23.5170 ;
        RECT 8.4650 23.1255 8.5410 23.2790 ;
        RECT 8.4790 22.4235 8.5050 23.5170 ;
        RECT 8.4790 22.5445 8.5190 22.7840 ;
        RECT 8.4790 22.4235 8.5410 22.5125 ;
        RECT 8.1820 22.8740 8.3880 23.5170 ;
        RECT 8.3620 22.4235 8.3880 23.5170 ;
        RECT 8.1820 23.1510 8.4020 23.4090 ;
        RECT 8.1820 22.4235 8.2800 23.5170 ;
        RECT 7.7650 22.4235 7.8480 23.5170 ;
        RECT 7.7650 22.5120 7.8620 23.4475 ;
        RECT 16.4440 22.4235 16.5290 23.5170 ;
        RECT 16.3000 22.4235 16.3260 23.5170 ;
        RECT 16.1920 22.4235 16.2180 23.5170 ;
        RECT 16.0840 22.4235 16.1100 23.5170 ;
        RECT 15.9760 22.4235 16.0020 23.5170 ;
        RECT 15.8680 22.4235 15.8940 23.5170 ;
        RECT 15.7600 22.4235 15.7860 23.5170 ;
        RECT 15.6520 22.4235 15.6780 23.5170 ;
        RECT 15.5440 22.4235 15.5700 23.5170 ;
        RECT 15.4360 22.4235 15.4620 23.5170 ;
        RECT 15.3280 22.4235 15.3540 23.5170 ;
        RECT 15.2200 22.4235 15.2460 23.5170 ;
        RECT 15.1120 22.4235 15.1380 23.5170 ;
        RECT 15.0040 22.4235 15.0300 23.5170 ;
        RECT 14.8960 22.4235 14.9220 23.5170 ;
        RECT 14.7880 22.4235 14.8140 23.5170 ;
        RECT 14.6800 22.4235 14.7060 23.5170 ;
        RECT 14.5720 22.4235 14.5980 23.5170 ;
        RECT 14.4640 22.4235 14.4900 23.5170 ;
        RECT 14.3560 22.4235 14.3820 23.5170 ;
        RECT 14.2480 22.4235 14.2740 23.5170 ;
        RECT 14.1400 22.4235 14.1660 23.5170 ;
        RECT 14.0320 22.4235 14.0580 23.5170 ;
        RECT 13.9240 22.4235 13.9500 23.5170 ;
        RECT 13.8160 22.4235 13.8420 23.5170 ;
        RECT 13.7080 22.4235 13.7340 23.5170 ;
        RECT 13.6000 22.4235 13.6260 23.5170 ;
        RECT 13.4920 22.4235 13.5180 23.5170 ;
        RECT 13.3840 22.4235 13.4100 23.5170 ;
        RECT 13.2760 22.4235 13.3020 23.5170 ;
        RECT 13.1680 22.4235 13.1940 23.5170 ;
        RECT 13.0600 22.4235 13.0860 23.5170 ;
        RECT 12.9520 22.4235 12.9780 23.5170 ;
        RECT 12.8440 22.4235 12.8700 23.5170 ;
        RECT 12.7360 22.4235 12.7620 23.5170 ;
        RECT 12.6280 22.4235 12.6540 23.5170 ;
        RECT 12.5200 22.4235 12.5460 23.5170 ;
        RECT 12.4120 22.4235 12.4380 23.5170 ;
        RECT 12.3040 22.4235 12.3300 23.5170 ;
        RECT 12.1960 22.4235 12.2220 23.5170 ;
        RECT 12.0880 22.4235 12.1140 23.5170 ;
        RECT 11.9800 22.4235 12.0060 23.5170 ;
        RECT 11.8720 22.4235 11.8980 23.5170 ;
        RECT 11.7640 22.4235 11.7900 23.5170 ;
        RECT 11.6560 22.4235 11.6820 23.5170 ;
        RECT 11.5480 22.4235 11.5740 23.5170 ;
        RECT 11.4400 22.4235 11.4660 23.5170 ;
        RECT 11.3320 22.4235 11.3580 23.5170 ;
        RECT 11.2240 22.4235 11.2500 23.5170 ;
        RECT 11.1160 22.4235 11.1420 23.5170 ;
        RECT 11.0080 22.4235 11.0340 23.5170 ;
        RECT 10.9000 22.4235 10.9260 23.5170 ;
        RECT 10.7920 22.4235 10.8180 23.5170 ;
        RECT 10.6840 22.4235 10.7100 23.5170 ;
        RECT 10.5760 22.4235 10.6020 23.5170 ;
        RECT 10.4680 22.4235 10.4940 23.5170 ;
        RECT 10.3600 22.4235 10.3860 23.5170 ;
        RECT 10.2520 22.4235 10.2780 23.5170 ;
        RECT 10.1440 22.4235 10.1700 23.5170 ;
        RECT 10.0360 22.4235 10.0620 23.5170 ;
        RECT 9.9280 22.4235 9.9540 23.5170 ;
        RECT 9.8200 22.4235 9.8460 23.5170 ;
        RECT 9.7120 22.4235 9.7380 23.5170 ;
        RECT 9.6040 22.4235 9.6300 23.5170 ;
        RECT 9.4960 22.4235 9.5220 23.5170 ;
        RECT 9.3880 22.4235 9.4140 23.5170 ;
        RECT 9.1750 22.4235 9.2520 23.5170 ;
        RECT 7.2820 22.4235 7.3590 23.5170 ;
        RECT 7.1200 22.4235 7.1460 23.5170 ;
        RECT 7.0120 22.4235 7.0380 23.5170 ;
        RECT 6.9040 22.4235 6.9300 23.5170 ;
        RECT 6.7960 22.4235 6.8220 23.5170 ;
        RECT 6.6880 22.4235 6.7140 23.5170 ;
        RECT 6.5800 22.4235 6.6060 23.5170 ;
        RECT 6.4720 22.4235 6.4980 23.5170 ;
        RECT 6.3640 22.4235 6.3900 23.5170 ;
        RECT 6.2560 22.4235 6.2820 23.5170 ;
        RECT 6.1480 22.4235 6.1740 23.5170 ;
        RECT 6.0400 22.4235 6.0660 23.5170 ;
        RECT 5.9320 22.4235 5.9580 23.5170 ;
        RECT 5.8240 22.4235 5.8500 23.5170 ;
        RECT 5.7160 22.4235 5.7420 23.5170 ;
        RECT 5.6080 22.4235 5.6340 23.5170 ;
        RECT 5.5000 22.4235 5.5260 23.5170 ;
        RECT 5.3920 22.4235 5.4180 23.5170 ;
        RECT 5.2840 22.4235 5.3100 23.5170 ;
        RECT 5.1760 22.4235 5.2020 23.5170 ;
        RECT 5.0680 22.4235 5.0940 23.5170 ;
        RECT 4.9600 22.4235 4.9860 23.5170 ;
        RECT 4.8520 22.4235 4.8780 23.5170 ;
        RECT 4.7440 22.4235 4.7700 23.5170 ;
        RECT 4.6360 22.4235 4.6620 23.5170 ;
        RECT 4.5280 22.4235 4.5540 23.5170 ;
        RECT 4.4200 22.4235 4.4460 23.5170 ;
        RECT 4.3120 22.4235 4.3380 23.5170 ;
        RECT 4.2040 22.4235 4.2300 23.5170 ;
        RECT 4.0960 22.4235 4.1220 23.5170 ;
        RECT 3.9880 22.4235 4.0140 23.5170 ;
        RECT 3.8800 22.4235 3.9060 23.5170 ;
        RECT 3.7720 22.4235 3.7980 23.5170 ;
        RECT 3.6640 22.4235 3.6900 23.5170 ;
        RECT 3.5560 22.4235 3.5820 23.5170 ;
        RECT 3.4480 22.4235 3.4740 23.5170 ;
        RECT 3.3400 22.4235 3.3660 23.5170 ;
        RECT 3.2320 22.4235 3.2580 23.5170 ;
        RECT 3.1240 22.4235 3.1500 23.5170 ;
        RECT 3.0160 22.4235 3.0420 23.5170 ;
        RECT 2.9080 22.4235 2.9340 23.5170 ;
        RECT 2.8000 22.4235 2.8260 23.5170 ;
        RECT 2.6920 22.4235 2.7180 23.5170 ;
        RECT 2.5840 22.4235 2.6100 23.5170 ;
        RECT 2.4760 22.4235 2.5020 23.5170 ;
        RECT 2.3680 22.4235 2.3940 23.5170 ;
        RECT 2.2600 22.4235 2.2860 23.5170 ;
        RECT 2.1520 22.4235 2.1780 23.5170 ;
        RECT 2.0440 22.4235 2.0700 23.5170 ;
        RECT 1.9360 22.4235 1.9620 23.5170 ;
        RECT 1.8280 22.4235 1.8540 23.5170 ;
        RECT 1.7200 22.4235 1.7460 23.5170 ;
        RECT 1.6120 22.4235 1.6380 23.5170 ;
        RECT 1.5040 22.4235 1.5300 23.5170 ;
        RECT 1.3960 22.4235 1.4220 23.5170 ;
        RECT 1.2880 22.4235 1.3140 23.5170 ;
        RECT 1.1800 22.4235 1.2060 23.5170 ;
        RECT 1.0720 22.4235 1.0980 23.5170 ;
        RECT 0.9640 22.4235 0.9900 23.5170 ;
        RECT 0.8560 22.4235 0.8820 23.5170 ;
        RECT 0.7480 22.4235 0.7740 23.5170 ;
        RECT 0.6400 22.4235 0.6660 23.5170 ;
        RECT 0.5320 22.4235 0.5580 23.5170 ;
        RECT 0.4240 22.4235 0.4500 23.5170 ;
        RECT 0.3160 22.4235 0.3420 23.5170 ;
        RECT 0.2080 22.4235 0.2340 23.5170 ;
        RECT 0.0050 22.4235 0.0900 23.5170 ;
        RECT 8.6410 23.5035 8.7690 24.5970 ;
        RECT 8.6270 24.1690 8.7690 24.4915 ;
        RECT 8.4790 23.8960 8.5410 24.5970 ;
        RECT 8.4650 24.2055 8.5410 24.3590 ;
        RECT 8.4790 23.5035 8.5050 24.5970 ;
        RECT 8.4790 23.6245 8.5190 23.8640 ;
        RECT 8.4790 23.5035 8.5410 23.5925 ;
        RECT 8.1820 23.9540 8.3880 24.5970 ;
        RECT 8.3620 23.5035 8.3880 24.5970 ;
        RECT 8.1820 24.2310 8.4020 24.4890 ;
        RECT 8.1820 23.5035 8.2800 24.5970 ;
        RECT 7.7650 23.5035 7.8480 24.5970 ;
        RECT 7.7650 23.5920 7.8620 24.5275 ;
        RECT 16.4440 23.5035 16.5290 24.5970 ;
        RECT 16.3000 23.5035 16.3260 24.5970 ;
        RECT 16.1920 23.5035 16.2180 24.5970 ;
        RECT 16.0840 23.5035 16.1100 24.5970 ;
        RECT 15.9760 23.5035 16.0020 24.5970 ;
        RECT 15.8680 23.5035 15.8940 24.5970 ;
        RECT 15.7600 23.5035 15.7860 24.5970 ;
        RECT 15.6520 23.5035 15.6780 24.5970 ;
        RECT 15.5440 23.5035 15.5700 24.5970 ;
        RECT 15.4360 23.5035 15.4620 24.5970 ;
        RECT 15.3280 23.5035 15.3540 24.5970 ;
        RECT 15.2200 23.5035 15.2460 24.5970 ;
        RECT 15.1120 23.5035 15.1380 24.5970 ;
        RECT 15.0040 23.5035 15.0300 24.5970 ;
        RECT 14.8960 23.5035 14.9220 24.5970 ;
        RECT 14.7880 23.5035 14.8140 24.5970 ;
        RECT 14.6800 23.5035 14.7060 24.5970 ;
        RECT 14.5720 23.5035 14.5980 24.5970 ;
        RECT 14.4640 23.5035 14.4900 24.5970 ;
        RECT 14.3560 23.5035 14.3820 24.5970 ;
        RECT 14.2480 23.5035 14.2740 24.5970 ;
        RECT 14.1400 23.5035 14.1660 24.5970 ;
        RECT 14.0320 23.5035 14.0580 24.5970 ;
        RECT 13.9240 23.5035 13.9500 24.5970 ;
        RECT 13.8160 23.5035 13.8420 24.5970 ;
        RECT 13.7080 23.5035 13.7340 24.5970 ;
        RECT 13.6000 23.5035 13.6260 24.5970 ;
        RECT 13.4920 23.5035 13.5180 24.5970 ;
        RECT 13.3840 23.5035 13.4100 24.5970 ;
        RECT 13.2760 23.5035 13.3020 24.5970 ;
        RECT 13.1680 23.5035 13.1940 24.5970 ;
        RECT 13.0600 23.5035 13.0860 24.5970 ;
        RECT 12.9520 23.5035 12.9780 24.5970 ;
        RECT 12.8440 23.5035 12.8700 24.5970 ;
        RECT 12.7360 23.5035 12.7620 24.5970 ;
        RECT 12.6280 23.5035 12.6540 24.5970 ;
        RECT 12.5200 23.5035 12.5460 24.5970 ;
        RECT 12.4120 23.5035 12.4380 24.5970 ;
        RECT 12.3040 23.5035 12.3300 24.5970 ;
        RECT 12.1960 23.5035 12.2220 24.5970 ;
        RECT 12.0880 23.5035 12.1140 24.5970 ;
        RECT 11.9800 23.5035 12.0060 24.5970 ;
        RECT 11.8720 23.5035 11.8980 24.5970 ;
        RECT 11.7640 23.5035 11.7900 24.5970 ;
        RECT 11.6560 23.5035 11.6820 24.5970 ;
        RECT 11.5480 23.5035 11.5740 24.5970 ;
        RECT 11.4400 23.5035 11.4660 24.5970 ;
        RECT 11.3320 23.5035 11.3580 24.5970 ;
        RECT 11.2240 23.5035 11.2500 24.5970 ;
        RECT 11.1160 23.5035 11.1420 24.5970 ;
        RECT 11.0080 23.5035 11.0340 24.5970 ;
        RECT 10.9000 23.5035 10.9260 24.5970 ;
        RECT 10.7920 23.5035 10.8180 24.5970 ;
        RECT 10.6840 23.5035 10.7100 24.5970 ;
        RECT 10.5760 23.5035 10.6020 24.5970 ;
        RECT 10.4680 23.5035 10.4940 24.5970 ;
        RECT 10.3600 23.5035 10.3860 24.5970 ;
        RECT 10.2520 23.5035 10.2780 24.5970 ;
        RECT 10.1440 23.5035 10.1700 24.5970 ;
        RECT 10.0360 23.5035 10.0620 24.5970 ;
        RECT 9.9280 23.5035 9.9540 24.5970 ;
        RECT 9.8200 23.5035 9.8460 24.5970 ;
        RECT 9.7120 23.5035 9.7380 24.5970 ;
        RECT 9.6040 23.5035 9.6300 24.5970 ;
        RECT 9.4960 23.5035 9.5220 24.5970 ;
        RECT 9.3880 23.5035 9.4140 24.5970 ;
        RECT 9.1750 23.5035 9.2520 24.5970 ;
        RECT 7.2820 23.5035 7.3590 24.5970 ;
        RECT 7.1200 23.5035 7.1460 24.5970 ;
        RECT 7.0120 23.5035 7.0380 24.5970 ;
        RECT 6.9040 23.5035 6.9300 24.5970 ;
        RECT 6.7960 23.5035 6.8220 24.5970 ;
        RECT 6.6880 23.5035 6.7140 24.5970 ;
        RECT 6.5800 23.5035 6.6060 24.5970 ;
        RECT 6.4720 23.5035 6.4980 24.5970 ;
        RECT 6.3640 23.5035 6.3900 24.5970 ;
        RECT 6.2560 23.5035 6.2820 24.5970 ;
        RECT 6.1480 23.5035 6.1740 24.5970 ;
        RECT 6.0400 23.5035 6.0660 24.5970 ;
        RECT 5.9320 23.5035 5.9580 24.5970 ;
        RECT 5.8240 23.5035 5.8500 24.5970 ;
        RECT 5.7160 23.5035 5.7420 24.5970 ;
        RECT 5.6080 23.5035 5.6340 24.5970 ;
        RECT 5.5000 23.5035 5.5260 24.5970 ;
        RECT 5.3920 23.5035 5.4180 24.5970 ;
        RECT 5.2840 23.5035 5.3100 24.5970 ;
        RECT 5.1760 23.5035 5.2020 24.5970 ;
        RECT 5.0680 23.5035 5.0940 24.5970 ;
        RECT 4.9600 23.5035 4.9860 24.5970 ;
        RECT 4.8520 23.5035 4.8780 24.5970 ;
        RECT 4.7440 23.5035 4.7700 24.5970 ;
        RECT 4.6360 23.5035 4.6620 24.5970 ;
        RECT 4.5280 23.5035 4.5540 24.5970 ;
        RECT 4.4200 23.5035 4.4460 24.5970 ;
        RECT 4.3120 23.5035 4.3380 24.5970 ;
        RECT 4.2040 23.5035 4.2300 24.5970 ;
        RECT 4.0960 23.5035 4.1220 24.5970 ;
        RECT 3.9880 23.5035 4.0140 24.5970 ;
        RECT 3.8800 23.5035 3.9060 24.5970 ;
        RECT 3.7720 23.5035 3.7980 24.5970 ;
        RECT 3.6640 23.5035 3.6900 24.5970 ;
        RECT 3.5560 23.5035 3.5820 24.5970 ;
        RECT 3.4480 23.5035 3.4740 24.5970 ;
        RECT 3.3400 23.5035 3.3660 24.5970 ;
        RECT 3.2320 23.5035 3.2580 24.5970 ;
        RECT 3.1240 23.5035 3.1500 24.5970 ;
        RECT 3.0160 23.5035 3.0420 24.5970 ;
        RECT 2.9080 23.5035 2.9340 24.5970 ;
        RECT 2.8000 23.5035 2.8260 24.5970 ;
        RECT 2.6920 23.5035 2.7180 24.5970 ;
        RECT 2.5840 23.5035 2.6100 24.5970 ;
        RECT 2.4760 23.5035 2.5020 24.5970 ;
        RECT 2.3680 23.5035 2.3940 24.5970 ;
        RECT 2.2600 23.5035 2.2860 24.5970 ;
        RECT 2.1520 23.5035 2.1780 24.5970 ;
        RECT 2.0440 23.5035 2.0700 24.5970 ;
        RECT 1.9360 23.5035 1.9620 24.5970 ;
        RECT 1.8280 23.5035 1.8540 24.5970 ;
        RECT 1.7200 23.5035 1.7460 24.5970 ;
        RECT 1.6120 23.5035 1.6380 24.5970 ;
        RECT 1.5040 23.5035 1.5300 24.5970 ;
        RECT 1.3960 23.5035 1.4220 24.5970 ;
        RECT 1.2880 23.5035 1.3140 24.5970 ;
        RECT 1.1800 23.5035 1.2060 24.5970 ;
        RECT 1.0720 23.5035 1.0980 24.5970 ;
        RECT 0.9640 23.5035 0.9900 24.5970 ;
        RECT 0.8560 23.5035 0.8820 24.5970 ;
        RECT 0.7480 23.5035 0.7740 24.5970 ;
        RECT 0.6400 23.5035 0.6660 24.5970 ;
        RECT 0.5320 23.5035 0.5580 24.5970 ;
        RECT 0.4240 23.5035 0.4500 24.5970 ;
        RECT 0.3160 23.5035 0.3420 24.5970 ;
        RECT 0.2080 23.5035 0.2340 24.5970 ;
        RECT 0.0050 23.5035 0.0900 24.5970 ;
        RECT 8.6410 24.5835 8.7690 25.6770 ;
        RECT 8.6270 25.2490 8.7690 25.5715 ;
        RECT 8.4790 24.9760 8.5410 25.6770 ;
        RECT 8.4650 25.2855 8.5410 25.4390 ;
        RECT 8.4790 24.5835 8.5050 25.6770 ;
        RECT 8.4790 24.7045 8.5190 24.9440 ;
        RECT 8.4790 24.5835 8.5410 24.6725 ;
        RECT 8.1820 25.0340 8.3880 25.6770 ;
        RECT 8.3620 24.5835 8.3880 25.6770 ;
        RECT 8.1820 25.3110 8.4020 25.5690 ;
        RECT 8.1820 24.5835 8.2800 25.6770 ;
        RECT 7.7650 24.5835 7.8480 25.6770 ;
        RECT 7.7650 24.6720 7.8620 25.6075 ;
        RECT 16.4440 24.5835 16.5290 25.6770 ;
        RECT 16.3000 24.5835 16.3260 25.6770 ;
        RECT 16.1920 24.5835 16.2180 25.6770 ;
        RECT 16.0840 24.5835 16.1100 25.6770 ;
        RECT 15.9760 24.5835 16.0020 25.6770 ;
        RECT 15.8680 24.5835 15.8940 25.6770 ;
        RECT 15.7600 24.5835 15.7860 25.6770 ;
        RECT 15.6520 24.5835 15.6780 25.6770 ;
        RECT 15.5440 24.5835 15.5700 25.6770 ;
        RECT 15.4360 24.5835 15.4620 25.6770 ;
        RECT 15.3280 24.5835 15.3540 25.6770 ;
        RECT 15.2200 24.5835 15.2460 25.6770 ;
        RECT 15.1120 24.5835 15.1380 25.6770 ;
        RECT 15.0040 24.5835 15.0300 25.6770 ;
        RECT 14.8960 24.5835 14.9220 25.6770 ;
        RECT 14.7880 24.5835 14.8140 25.6770 ;
        RECT 14.6800 24.5835 14.7060 25.6770 ;
        RECT 14.5720 24.5835 14.5980 25.6770 ;
        RECT 14.4640 24.5835 14.4900 25.6770 ;
        RECT 14.3560 24.5835 14.3820 25.6770 ;
        RECT 14.2480 24.5835 14.2740 25.6770 ;
        RECT 14.1400 24.5835 14.1660 25.6770 ;
        RECT 14.0320 24.5835 14.0580 25.6770 ;
        RECT 13.9240 24.5835 13.9500 25.6770 ;
        RECT 13.8160 24.5835 13.8420 25.6770 ;
        RECT 13.7080 24.5835 13.7340 25.6770 ;
        RECT 13.6000 24.5835 13.6260 25.6770 ;
        RECT 13.4920 24.5835 13.5180 25.6770 ;
        RECT 13.3840 24.5835 13.4100 25.6770 ;
        RECT 13.2760 24.5835 13.3020 25.6770 ;
        RECT 13.1680 24.5835 13.1940 25.6770 ;
        RECT 13.0600 24.5835 13.0860 25.6770 ;
        RECT 12.9520 24.5835 12.9780 25.6770 ;
        RECT 12.8440 24.5835 12.8700 25.6770 ;
        RECT 12.7360 24.5835 12.7620 25.6770 ;
        RECT 12.6280 24.5835 12.6540 25.6770 ;
        RECT 12.5200 24.5835 12.5460 25.6770 ;
        RECT 12.4120 24.5835 12.4380 25.6770 ;
        RECT 12.3040 24.5835 12.3300 25.6770 ;
        RECT 12.1960 24.5835 12.2220 25.6770 ;
        RECT 12.0880 24.5835 12.1140 25.6770 ;
        RECT 11.9800 24.5835 12.0060 25.6770 ;
        RECT 11.8720 24.5835 11.8980 25.6770 ;
        RECT 11.7640 24.5835 11.7900 25.6770 ;
        RECT 11.6560 24.5835 11.6820 25.6770 ;
        RECT 11.5480 24.5835 11.5740 25.6770 ;
        RECT 11.4400 24.5835 11.4660 25.6770 ;
        RECT 11.3320 24.5835 11.3580 25.6770 ;
        RECT 11.2240 24.5835 11.2500 25.6770 ;
        RECT 11.1160 24.5835 11.1420 25.6770 ;
        RECT 11.0080 24.5835 11.0340 25.6770 ;
        RECT 10.9000 24.5835 10.9260 25.6770 ;
        RECT 10.7920 24.5835 10.8180 25.6770 ;
        RECT 10.6840 24.5835 10.7100 25.6770 ;
        RECT 10.5760 24.5835 10.6020 25.6770 ;
        RECT 10.4680 24.5835 10.4940 25.6770 ;
        RECT 10.3600 24.5835 10.3860 25.6770 ;
        RECT 10.2520 24.5835 10.2780 25.6770 ;
        RECT 10.1440 24.5835 10.1700 25.6770 ;
        RECT 10.0360 24.5835 10.0620 25.6770 ;
        RECT 9.9280 24.5835 9.9540 25.6770 ;
        RECT 9.8200 24.5835 9.8460 25.6770 ;
        RECT 9.7120 24.5835 9.7380 25.6770 ;
        RECT 9.6040 24.5835 9.6300 25.6770 ;
        RECT 9.4960 24.5835 9.5220 25.6770 ;
        RECT 9.3880 24.5835 9.4140 25.6770 ;
        RECT 9.1750 24.5835 9.2520 25.6770 ;
        RECT 7.2820 24.5835 7.3590 25.6770 ;
        RECT 7.1200 24.5835 7.1460 25.6770 ;
        RECT 7.0120 24.5835 7.0380 25.6770 ;
        RECT 6.9040 24.5835 6.9300 25.6770 ;
        RECT 6.7960 24.5835 6.8220 25.6770 ;
        RECT 6.6880 24.5835 6.7140 25.6770 ;
        RECT 6.5800 24.5835 6.6060 25.6770 ;
        RECT 6.4720 24.5835 6.4980 25.6770 ;
        RECT 6.3640 24.5835 6.3900 25.6770 ;
        RECT 6.2560 24.5835 6.2820 25.6770 ;
        RECT 6.1480 24.5835 6.1740 25.6770 ;
        RECT 6.0400 24.5835 6.0660 25.6770 ;
        RECT 5.9320 24.5835 5.9580 25.6770 ;
        RECT 5.8240 24.5835 5.8500 25.6770 ;
        RECT 5.7160 24.5835 5.7420 25.6770 ;
        RECT 5.6080 24.5835 5.6340 25.6770 ;
        RECT 5.5000 24.5835 5.5260 25.6770 ;
        RECT 5.3920 24.5835 5.4180 25.6770 ;
        RECT 5.2840 24.5835 5.3100 25.6770 ;
        RECT 5.1760 24.5835 5.2020 25.6770 ;
        RECT 5.0680 24.5835 5.0940 25.6770 ;
        RECT 4.9600 24.5835 4.9860 25.6770 ;
        RECT 4.8520 24.5835 4.8780 25.6770 ;
        RECT 4.7440 24.5835 4.7700 25.6770 ;
        RECT 4.6360 24.5835 4.6620 25.6770 ;
        RECT 4.5280 24.5835 4.5540 25.6770 ;
        RECT 4.4200 24.5835 4.4460 25.6770 ;
        RECT 4.3120 24.5835 4.3380 25.6770 ;
        RECT 4.2040 24.5835 4.2300 25.6770 ;
        RECT 4.0960 24.5835 4.1220 25.6770 ;
        RECT 3.9880 24.5835 4.0140 25.6770 ;
        RECT 3.8800 24.5835 3.9060 25.6770 ;
        RECT 3.7720 24.5835 3.7980 25.6770 ;
        RECT 3.6640 24.5835 3.6900 25.6770 ;
        RECT 3.5560 24.5835 3.5820 25.6770 ;
        RECT 3.4480 24.5835 3.4740 25.6770 ;
        RECT 3.3400 24.5835 3.3660 25.6770 ;
        RECT 3.2320 24.5835 3.2580 25.6770 ;
        RECT 3.1240 24.5835 3.1500 25.6770 ;
        RECT 3.0160 24.5835 3.0420 25.6770 ;
        RECT 2.9080 24.5835 2.9340 25.6770 ;
        RECT 2.8000 24.5835 2.8260 25.6770 ;
        RECT 2.6920 24.5835 2.7180 25.6770 ;
        RECT 2.5840 24.5835 2.6100 25.6770 ;
        RECT 2.4760 24.5835 2.5020 25.6770 ;
        RECT 2.3680 24.5835 2.3940 25.6770 ;
        RECT 2.2600 24.5835 2.2860 25.6770 ;
        RECT 2.1520 24.5835 2.1780 25.6770 ;
        RECT 2.0440 24.5835 2.0700 25.6770 ;
        RECT 1.9360 24.5835 1.9620 25.6770 ;
        RECT 1.8280 24.5835 1.8540 25.6770 ;
        RECT 1.7200 24.5835 1.7460 25.6770 ;
        RECT 1.6120 24.5835 1.6380 25.6770 ;
        RECT 1.5040 24.5835 1.5300 25.6770 ;
        RECT 1.3960 24.5835 1.4220 25.6770 ;
        RECT 1.2880 24.5835 1.3140 25.6770 ;
        RECT 1.1800 24.5835 1.2060 25.6770 ;
        RECT 1.0720 24.5835 1.0980 25.6770 ;
        RECT 0.9640 24.5835 0.9900 25.6770 ;
        RECT 0.8560 24.5835 0.8820 25.6770 ;
        RECT 0.7480 24.5835 0.7740 25.6770 ;
        RECT 0.6400 24.5835 0.6660 25.6770 ;
        RECT 0.5320 24.5835 0.5580 25.6770 ;
        RECT 0.4240 24.5835 0.4500 25.6770 ;
        RECT 0.3160 24.5835 0.3420 25.6770 ;
        RECT 0.2080 24.5835 0.2340 25.6770 ;
        RECT 0.0050 24.5835 0.0900 25.6770 ;
        RECT 8.6410 25.6635 8.7690 26.7570 ;
        RECT 8.6270 26.3290 8.7690 26.6515 ;
        RECT 8.4790 26.0560 8.5410 26.7570 ;
        RECT 8.4650 26.3655 8.5410 26.5190 ;
        RECT 8.4790 25.6635 8.5050 26.7570 ;
        RECT 8.4790 25.7845 8.5190 26.0240 ;
        RECT 8.4790 25.6635 8.5410 25.7525 ;
        RECT 8.1820 26.1140 8.3880 26.7570 ;
        RECT 8.3620 25.6635 8.3880 26.7570 ;
        RECT 8.1820 26.3910 8.4020 26.6490 ;
        RECT 8.1820 25.6635 8.2800 26.7570 ;
        RECT 7.7650 25.6635 7.8480 26.7570 ;
        RECT 7.7650 25.7520 7.8620 26.6875 ;
        RECT 16.4440 25.6635 16.5290 26.7570 ;
        RECT 16.3000 25.6635 16.3260 26.7570 ;
        RECT 16.1920 25.6635 16.2180 26.7570 ;
        RECT 16.0840 25.6635 16.1100 26.7570 ;
        RECT 15.9760 25.6635 16.0020 26.7570 ;
        RECT 15.8680 25.6635 15.8940 26.7570 ;
        RECT 15.7600 25.6635 15.7860 26.7570 ;
        RECT 15.6520 25.6635 15.6780 26.7570 ;
        RECT 15.5440 25.6635 15.5700 26.7570 ;
        RECT 15.4360 25.6635 15.4620 26.7570 ;
        RECT 15.3280 25.6635 15.3540 26.7570 ;
        RECT 15.2200 25.6635 15.2460 26.7570 ;
        RECT 15.1120 25.6635 15.1380 26.7570 ;
        RECT 15.0040 25.6635 15.0300 26.7570 ;
        RECT 14.8960 25.6635 14.9220 26.7570 ;
        RECT 14.7880 25.6635 14.8140 26.7570 ;
        RECT 14.6800 25.6635 14.7060 26.7570 ;
        RECT 14.5720 25.6635 14.5980 26.7570 ;
        RECT 14.4640 25.6635 14.4900 26.7570 ;
        RECT 14.3560 25.6635 14.3820 26.7570 ;
        RECT 14.2480 25.6635 14.2740 26.7570 ;
        RECT 14.1400 25.6635 14.1660 26.7570 ;
        RECT 14.0320 25.6635 14.0580 26.7570 ;
        RECT 13.9240 25.6635 13.9500 26.7570 ;
        RECT 13.8160 25.6635 13.8420 26.7570 ;
        RECT 13.7080 25.6635 13.7340 26.7570 ;
        RECT 13.6000 25.6635 13.6260 26.7570 ;
        RECT 13.4920 25.6635 13.5180 26.7570 ;
        RECT 13.3840 25.6635 13.4100 26.7570 ;
        RECT 13.2760 25.6635 13.3020 26.7570 ;
        RECT 13.1680 25.6635 13.1940 26.7570 ;
        RECT 13.0600 25.6635 13.0860 26.7570 ;
        RECT 12.9520 25.6635 12.9780 26.7570 ;
        RECT 12.8440 25.6635 12.8700 26.7570 ;
        RECT 12.7360 25.6635 12.7620 26.7570 ;
        RECT 12.6280 25.6635 12.6540 26.7570 ;
        RECT 12.5200 25.6635 12.5460 26.7570 ;
        RECT 12.4120 25.6635 12.4380 26.7570 ;
        RECT 12.3040 25.6635 12.3300 26.7570 ;
        RECT 12.1960 25.6635 12.2220 26.7570 ;
        RECT 12.0880 25.6635 12.1140 26.7570 ;
        RECT 11.9800 25.6635 12.0060 26.7570 ;
        RECT 11.8720 25.6635 11.8980 26.7570 ;
        RECT 11.7640 25.6635 11.7900 26.7570 ;
        RECT 11.6560 25.6635 11.6820 26.7570 ;
        RECT 11.5480 25.6635 11.5740 26.7570 ;
        RECT 11.4400 25.6635 11.4660 26.7570 ;
        RECT 11.3320 25.6635 11.3580 26.7570 ;
        RECT 11.2240 25.6635 11.2500 26.7570 ;
        RECT 11.1160 25.6635 11.1420 26.7570 ;
        RECT 11.0080 25.6635 11.0340 26.7570 ;
        RECT 10.9000 25.6635 10.9260 26.7570 ;
        RECT 10.7920 25.6635 10.8180 26.7570 ;
        RECT 10.6840 25.6635 10.7100 26.7570 ;
        RECT 10.5760 25.6635 10.6020 26.7570 ;
        RECT 10.4680 25.6635 10.4940 26.7570 ;
        RECT 10.3600 25.6635 10.3860 26.7570 ;
        RECT 10.2520 25.6635 10.2780 26.7570 ;
        RECT 10.1440 25.6635 10.1700 26.7570 ;
        RECT 10.0360 25.6635 10.0620 26.7570 ;
        RECT 9.9280 25.6635 9.9540 26.7570 ;
        RECT 9.8200 25.6635 9.8460 26.7570 ;
        RECT 9.7120 25.6635 9.7380 26.7570 ;
        RECT 9.6040 25.6635 9.6300 26.7570 ;
        RECT 9.4960 25.6635 9.5220 26.7570 ;
        RECT 9.3880 25.6635 9.4140 26.7570 ;
        RECT 9.1750 25.6635 9.2520 26.7570 ;
        RECT 7.2820 25.6635 7.3590 26.7570 ;
        RECT 7.1200 25.6635 7.1460 26.7570 ;
        RECT 7.0120 25.6635 7.0380 26.7570 ;
        RECT 6.9040 25.6635 6.9300 26.7570 ;
        RECT 6.7960 25.6635 6.8220 26.7570 ;
        RECT 6.6880 25.6635 6.7140 26.7570 ;
        RECT 6.5800 25.6635 6.6060 26.7570 ;
        RECT 6.4720 25.6635 6.4980 26.7570 ;
        RECT 6.3640 25.6635 6.3900 26.7570 ;
        RECT 6.2560 25.6635 6.2820 26.7570 ;
        RECT 6.1480 25.6635 6.1740 26.7570 ;
        RECT 6.0400 25.6635 6.0660 26.7570 ;
        RECT 5.9320 25.6635 5.9580 26.7570 ;
        RECT 5.8240 25.6635 5.8500 26.7570 ;
        RECT 5.7160 25.6635 5.7420 26.7570 ;
        RECT 5.6080 25.6635 5.6340 26.7570 ;
        RECT 5.5000 25.6635 5.5260 26.7570 ;
        RECT 5.3920 25.6635 5.4180 26.7570 ;
        RECT 5.2840 25.6635 5.3100 26.7570 ;
        RECT 5.1760 25.6635 5.2020 26.7570 ;
        RECT 5.0680 25.6635 5.0940 26.7570 ;
        RECT 4.9600 25.6635 4.9860 26.7570 ;
        RECT 4.8520 25.6635 4.8780 26.7570 ;
        RECT 4.7440 25.6635 4.7700 26.7570 ;
        RECT 4.6360 25.6635 4.6620 26.7570 ;
        RECT 4.5280 25.6635 4.5540 26.7570 ;
        RECT 4.4200 25.6635 4.4460 26.7570 ;
        RECT 4.3120 25.6635 4.3380 26.7570 ;
        RECT 4.2040 25.6635 4.2300 26.7570 ;
        RECT 4.0960 25.6635 4.1220 26.7570 ;
        RECT 3.9880 25.6635 4.0140 26.7570 ;
        RECT 3.8800 25.6635 3.9060 26.7570 ;
        RECT 3.7720 25.6635 3.7980 26.7570 ;
        RECT 3.6640 25.6635 3.6900 26.7570 ;
        RECT 3.5560 25.6635 3.5820 26.7570 ;
        RECT 3.4480 25.6635 3.4740 26.7570 ;
        RECT 3.3400 25.6635 3.3660 26.7570 ;
        RECT 3.2320 25.6635 3.2580 26.7570 ;
        RECT 3.1240 25.6635 3.1500 26.7570 ;
        RECT 3.0160 25.6635 3.0420 26.7570 ;
        RECT 2.9080 25.6635 2.9340 26.7570 ;
        RECT 2.8000 25.6635 2.8260 26.7570 ;
        RECT 2.6920 25.6635 2.7180 26.7570 ;
        RECT 2.5840 25.6635 2.6100 26.7570 ;
        RECT 2.4760 25.6635 2.5020 26.7570 ;
        RECT 2.3680 25.6635 2.3940 26.7570 ;
        RECT 2.2600 25.6635 2.2860 26.7570 ;
        RECT 2.1520 25.6635 2.1780 26.7570 ;
        RECT 2.0440 25.6635 2.0700 26.7570 ;
        RECT 1.9360 25.6635 1.9620 26.7570 ;
        RECT 1.8280 25.6635 1.8540 26.7570 ;
        RECT 1.7200 25.6635 1.7460 26.7570 ;
        RECT 1.6120 25.6635 1.6380 26.7570 ;
        RECT 1.5040 25.6635 1.5300 26.7570 ;
        RECT 1.3960 25.6635 1.4220 26.7570 ;
        RECT 1.2880 25.6635 1.3140 26.7570 ;
        RECT 1.1800 25.6635 1.2060 26.7570 ;
        RECT 1.0720 25.6635 1.0980 26.7570 ;
        RECT 0.9640 25.6635 0.9900 26.7570 ;
        RECT 0.8560 25.6635 0.8820 26.7570 ;
        RECT 0.7480 25.6635 0.7740 26.7570 ;
        RECT 0.6400 25.6635 0.6660 26.7570 ;
        RECT 0.5320 25.6635 0.5580 26.7570 ;
        RECT 0.4240 25.6635 0.4500 26.7570 ;
        RECT 0.3160 25.6635 0.3420 26.7570 ;
        RECT 0.2080 25.6635 0.2340 26.7570 ;
        RECT 0.0050 25.6635 0.0900 26.7570 ;
        RECT 8.6410 26.7435 8.7690 27.8370 ;
        RECT 8.6270 27.4090 8.7690 27.7315 ;
        RECT 8.4790 27.1360 8.5410 27.8370 ;
        RECT 8.4650 27.4455 8.5410 27.5990 ;
        RECT 8.4790 26.7435 8.5050 27.8370 ;
        RECT 8.4790 26.8645 8.5190 27.1040 ;
        RECT 8.4790 26.7435 8.5410 26.8325 ;
        RECT 8.1820 27.1940 8.3880 27.8370 ;
        RECT 8.3620 26.7435 8.3880 27.8370 ;
        RECT 8.1820 27.4710 8.4020 27.7290 ;
        RECT 8.1820 26.7435 8.2800 27.8370 ;
        RECT 7.7650 26.7435 7.8480 27.8370 ;
        RECT 7.7650 26.8320 7.8620 27.7675 ;
        RECT 16.4440 26.7435 16.5290 27.8370 ;
        RECT 16.3000 26.7435 16.3260 27.8370 ;
        RECT 16.1920 26.7435 16.2180 27.8370 ;
        RECT 16.0840 26.7435 16.1100 27.8370 ;
        RECT 15.9760 26.7435 16.0020 27.8370 ;
        RECT 15.8680 26.7435 15.8940 27.8370 ;
        RECT 15.7600 26.7435 15.7860 27.8370 ;
        RECT 15.6520 26.7435 15.6780 27.8370 ;
        RECT 15.5440 26.7435 15.5700 27.8370 ;
        RECT 15.4360 26.7435 15.4620 27.8370 ;
        RECT 15.3280 26.7435 15.3540 27.8370 ;
        RECT 15.2200 26.7435 15.2460 27.8370 ;
        RECT 15.1120 26.7435 15.1380 27.8370 ;
        RECT 15.0040 26.7435 15.0300 27.8370 ;
        RECT 14.8960 26.7435 14.9220 27.8370 ;
        RECT 14.7880 26.7435 14.8140 27.8370 ;
        RECT 14.6800 26.7435 14.7060 27.8370 ;
        RECT 14.5720 26.7435 14.5980 27.8370 ;
        RECT 14.4640 26.7435 14.4900 27.8370 ;
        RECT 14.3560 26.7435 14.3820 27.8370 ;
        RECT 14.2480 26.7435 14.2740 27.8370 ;
        RECT 14.1400 26.7435 14.1660 27.8370 ;
        RECT 14.0320 26.7435 14.0580 27.8370 ;
        RECT 13.9240 26.7435 13.9500 27.8370 ;
        RECT 13.8160 26.7435 13.8420 27.8370 ;
        RECT 13.7080 26.7435 13.7340 27.8370 ;
        RECT 13.6000 26.7435 13.6260 27.8370 ;
        RECT 13.4920 26.7435 13.5180 27.8370 ;
        RECT 13.3840 26.7435 13.4100 27.8370 ;
        RECT 13.2760 26.7435 13.3020 27.8370 ;
        RECT 13.1680 26.7435 13.1940 27.8370 ;
        RECT 13.0600 26.7435 13.0860 27.8370 ;
        RECT 12.9520 26.7435 12.9780 27.8370 ;
        RECT 12.8440 26.7435 12.8700 27.8370 ;
        RECT 12.7360 26.7435 12.7620 27.8370 ;
        RECT 12.6280 26.7435 12.6540 27.8370 ;
        RECT 12.5200 26.7435 12.5460 27.8370 ;
        RECT 12.4120 26.7435 12.4380 27.8370 ;
        RECT 12.3040 26.7435 12.3300 27.8370 ;
        RECT 12.1960 26.7435 12.2220 27.8370 ;
        RECT 12.0880 26.7435 12.1140 27.8370 ;
        RECT 11.9800 26.7435 12.0060 27.8370 ;
        RECT 11.8720 26.7435 11.8980 27.8370 ;
        RECT 11.7640 26.7435 11.7900 27.8370 ;
        RECT 11.6560 26.7435 11.6820 27.8370 ;
        RECT 11.5480 26.7435 11.5740 27.8370 ;
        RECT 11.4400 26.7435 11.4660 27.8370 ;
        RECT 11.3320 26.7435 11.3580 27.8370 ;
        RECT 11.2240 26.7435 11.2500 27.8370 ;
        RECT 11.1160 26.7435 11.1420 27.8370 ;
        RECT 11.0080 26.7435 11.0340 27.8370 ;
        RECT 10.9000 26.7435 10.9260 27.8370 ;
        RECT 10.7920 26.7435 10.8180 27.8370 ;
        RECT 10.6840 26.7435 10.7100 27.8370 ;
        RECT 10.5760 26.7435 10.6020 27.8370 ;
        RECT 10.4680 26.7435 10.4940 27.8370 ;
        RECT 10.3600 26.7435 10.3860 27.8370 ;
        RECT 10.2520 26.7435 10.2780 27.8370 ;
        RECT 10.1440 26.7435 10.1700 27.8370 ;
        RECT 10.0360 26.7435 10.0620 27.8370 ;
        RECT 9.9280 26.7435 9.9540 27.8370 ;
        RECT 9.8200 26.7435 9.8460 27.8370 ;
        RECT 9.7120 26.7435 9.7380 27.8370 ;
        RECT 9.6040 26.7435 9.6300 27.8370 ;
        RECT 9.4960 26.7435 9.5220 27.8370 ;
        RECT 9.3880 26.7435 9.4140 27.8370 ;
        RECT 9.1750 26.7435 9.2520 27.8370 ;
        RECT 7.2820 26.7435 7.3590 27.8370 ;
        RECT 7.1200 26.7435 7.1460 27.8370 ;
        RECT 7.0120 26.7435 7.0380 27.8370 ;
        RECT 6.9040 26.7435 6.9300 27.8370 ;
        RECT 6.7960 26.7435 6.8220 27.8370 ;
        RECT 6.6880 26.7435 6.7140 27.8370 ;
        RECT 6.5800 26.7435 6.6060 27.8370 ;
        RECT 6.4720 26.7435 6.4980 27.8370 ;
        RECT 6.3640 26.7435 6.3900 27.8370 ;
        RECT 6.2560 26.7435 6.2820 27.8370 ;
        RECT 6.1480 26.7435 6.1740 27.8370 ;
        RECT 6.0400 26.7435 6.0660 27.8370 ;
        RECT 5.9320 26.7435 5.9580 27.8370 ;
        RECT 5.8240 26.7435 5.8500 27.8370 ;
        RECT 5.7160 26.7435 5.7420 27.8370 ;
        RECT 5.6080 26.7435 5.6340 27.8370 ;
        RECT 5.5000 26.7435 5.5260 27.8370 ;
        RECT 5.3920 26.7435 5.4180 27.8370 ;
        RECT 5.2840 26.7435 5.3100 27.8370 ;
        RECT 5.1760 26.7435 5.2020 27.8370 ;
        RECT 5.0680 26.7435 5.0940 27.8370 ;
        RECT 4.9600 26.7435 4.9860 27.8370 ;
        RECT 4.8520 26.7435 4.8780 27.8370 ;
        RECT 4.7440 26.7435 4.7700 27.8370 ;
        RECT 4.6360 26.7435 4.6620 27.8370 ;
        RECT 4.5280 26.7435 4.5540 27.8370 ;
        RECT 4.4200 26.7435 4.4460 27.8370 ;
        RECT 4.3120 26.7435 4.3380 27.8370 ;
        RECT 4.2040 26.7435 4.2300 27.8370 ;
        RECT 4.0960 26.7435 4.1220 27.8370 ;
        RECT 3.9880 26.7435 4.0140 27.8370 ;
        RECT 3.8800 26.7435 3.9060 27.8370 ;
        RECT 3.7720 26.7435 3.7980 27.8370 ;
        RECT 3.6640 26.7435 3.6900 27.8370 ;
        RECT 3.5560 26.7435 3.5820 27.8370 ;
        RECT 3.4480 26.7435 3.4740 27.8370 ;
        RECT 3.3400 26.7435 3.3660 27.8370 ;
        RECT 3.2320 26.7435 3.2580 27.8370 ;
        RECT 3.1240 26.7435 3.1500 27.8370 ;
        RECT 3.0160 26.7435 3.0420 27.8370 ;
        RECT 2.9080 26.7435 2.9340 27.8370 ;
        RECT 2.8000 26.7435 2.8260 27.8370 ;
        RECT 2.6920 26.7435 2.7180 27.8370 ;
        RECT 2.5840 26.7435 2.6100 27.8370 ;
        RECT 2.4760 26.7435 2.5020 27.8370 ;
        RECT 2.3680 26.7435 2.3940 27.8370 ;
        RECT 2.2600 26.7435 2.2860 27.8370 ;
        RECT 2.1520 26.7435 2.1780 27.8370 ;
        RECT 2.0440 26.7435 2.0700 27.8370 ;
        RECT 1.9360 26.7435 1.9620 27.8370 ;
        RECT 1.8280 26.7435 1.8540 27.8370 ;
        RECT 1.7200 26.7435 1.7460 27.8370 ;
        RECT 1.6120 26.7435 1.6380 27.8370 ;
        RECT 1.5040 26.7435 1.5300 27.8370 ;
        RECT 1.3960 26.7435 1.4220 27.8370 ;
        RECT 1.2880 26.7435 1.3140 27.8370 ;
        RECT 1.1800 26.7435 1.2060 27.8370 ;
        RECT 1.0720 26.7435 1.0980 27.8370 ;
        RECT 0.9640 26.7435 0.9900 27.8370 ;
        RECT 0.8560 26.7435 0.8820 27.8370 ;
        RECT 0.7480 26.7435 0.7740 27.8370 ;
        RECT 0.6400 26.7435 0.6660 27.8370 ;
        RECT 0.5320 26.7435 0.5580 27.8370 ;
        RECT 0.4240 26.7435 0.4500 27.8370 ;
        RECT 0.3160 26.7435 0.3420 27.8370 ;
        RECT 0.2080 26.7435 0.2340 27.8370 ;
        RECT 0.0050 26.7435 0.0900 27.8370 ;
        RECT 8.6410 27.8235 8.7690 28.9170 ;
        RECT 8.6270 28.4890 8.7690 28.8115 ;
        RECT 8.4790 28.2160 8.5410 28.9170 ;
        RECT 8.4650 28.5255 8.5410 28.6790 ;
        RECT 8.4790 27.8235 8.5050 28.9170 ;
        RECT 8.4790 27.9445 8.5190 28.1840 ;
        RECT 8.4790 27.8235 8.5410 27.9125 ;
        RECT 8.1820 28.2740 8.3880 28.9170 ;
        RECT 8.3620 27.8235 8.3880 28.9170 ;
        RECT 8.1820 28.5510 8.4020 28.8090 ;
        RECT 8.1820 27.8235 8.2800 28.9170 ;
        RECT 7.7650 27.8235 7.8480 28.9170 ;
        RECT 7.7650 27.9120 7.8620 28.8475 ;
        RECT 16.4440 27.8235 16.5290 28.9170 ;
        RECT 16.3000 27.8235 16.3260 28.9170 ;
        RECT 16.1920 27.8235 16.2180 28.9170 ;
        RECT 16.0840 27.8235 16.1100 28.9170 ;
        RECT 15.9760 27.8235 16.0020 28.9170 ;
        RECT 15.8680 27.8235 15.8940 28.9170 ;
        RECT 15.7600 27.8235 15.7860 28.9170 ;
        RECT 15.6520 27.8235 15.6780 28.9170 ;
        RECT 15.5440 27.8235 15.5700 28.9170 ;
        RECT 15.4360 27.8235 15.4620 28.9170 ;
        RECT 15.3280 27.8235 15.3540 28.9170 ;
        RECT 15.2200 27.8235 15.2460 28.9170 ;
        RECT 15.1120 27.8235 15.1380 28.9170 ;
        RECT 15.0040 27.8235 15.0300 28.9170 ;
        RECT 14.8960 27.8235 14.9220 28.9170 ;
        RECT 14.7880 27.8235 14.8140 28.9170 ;
        RECT 14.6800 27.8235 14.7060 28.9170 ;
        RECT 14.5720 27.8235 14.5980 28.9170 ;
        RECT 14.4640 27.8235 14.4900 28.9170 ;
        RECT 14.3560 27.8235 14.3820 28.9170 ;
        RECT 14.2480 27.8235 14.2740 28.9170 ;
        RECT 14.1400 27.8235 14.1660 28.9170 ;
        RECT 14.0320 27.8235 14.0580 28.9170 ;
        RECT 13.9240 27.8235 13.9500 28.9170 ;
        RECT 13.8160 27.8235 13.8420 28.9170 ;
        RECT 13.7080 27.8235 13.7340 28.9170 ;
        RECT 13.6000 27.8235 13.6260 28.9170 ;
        RECT 13.4920 27.8235 13.5180 28.9170 ;
        RECT 13.3840 27.8235 13.4100 28.9170 ;
        RECT 13.2760 27.8235 13.3020 28.9170 ;
        RECT 13.1680 27.8235 13.1940 28.9170 ;
        RECT 13.0600 27.8235 13.0860 28.9170 ;
        RECT 12.9520 27.8235 12.9780 28.9170 ;
        RECT 12.8440 27.8235 12.8700 28.9170 ;
        RECT 12.7360 27.8235 12.7620 28.9170 ;
        RECT 12.6280 27.8235 12.6540 28.9170 ;
        RECT 12.5200 27.8235 12.5460 28.9170 ;
        RECT 12.4120 27.8235 12.4380 28.9170 ;
        RECT 12.3040 27.8235 12.3300 28.9170 ;
        RECT 12.1960 27.8235 12.2220 28.9170 ;
        RECT 12.0880 27.8235 12.1140 28.9170 ;
        RECT 11.9800 27.8235 12.0060 28.9170 ;
        RECT 11.8720 27.8235 11.8980 28.9170 ;
        RECT 11.7640 27.8235 11.7900 28.9170 ;
        RECT 11.6560 27.8235 11.6820 28.9170 ;
        RECT 11.5480 27.8235 11.5740 28.9170 ;
        RECT 11.4400 27.8235 11.4660 28.9170 ;
        RECT 11.3320 27.8235 11.3580 28.9170 ;
        RECT 11.2240 27.8235 11.2500 28.9170 ;
        RECT 11.1160 27.8235 11.1420 28.9170 ;
        RECT 11.0080 27.8235 11.0340 28.9170 ;
        RECT 10.9000 27.8235 10.9260 28.9170 ;
        RECT 10.7920 27.8235 10.8180 28.9170 ;
        RECT 10.6840 27.8235 10.7100 28.9170 ;
        RECT 10.5760 27.8235 10.6020 28.9170 ;
        RECT 10.4680 27.8235 10.4940 28.9170 ;
        RECT 10.3600 27.8235 10.3860 28.9170 ;
        RECT 10.2520 27.8235 10.2780 28.9170 ;
        RECT 10.1440 27.8235 10.1700 28.9170 ;
        RECT 10.0360 27.8235 10.0620 28.9170 ;
        RECT 9.9280 27.8235 9.9540 28.9170 ;
        RECT 9.8200 27.8235 9.8460 28.9170 ;
        RECT 9.7120 27.8235 9.7380 28.9170 ;
        RECT 9.6040 27.8235 9.6300 28.9170 ;
        RECT 9.4960 27.8235 9.5220 28.9170 ;
        RECT 9.3880 27.8235 9.4140 28.9170 ;
        RECT 9.1750 27.8235 9.2520 28.9170 ;
        RECT 7.2820 27.8235 7.3590 28.9170 ;
        RECT 7.1200 27.8235 7.1460 28.9170 ;
        RECT 7.0120 27.8235 7.0380 28.9170 ;
        RECT 6.9040 27.8235 6.9300 28.9170 ;
        RECT 6.7960 27.8235 6.8220 28.9170 ;
        RECT 6.6880 27.8235 6.7140 28.9170 ;
        RECT 6.5800 27.8235 6.6060 28.9170 ;
        RECT 6.4720 27.8235 6.4980 28.9170 ;
        RECT 6.3640 27.8235 6.3900 28.9170 ;
        RECT 6.2560 27.8235 6.2820 28.9170 ;
        RECT 6.1480 27.8235 6.1740 28.9170 ;
        RECT 6.0400 27.8235 6.0660 28.9170 ;
        RECT 5.9320 27.8235 5.9580 28.9170 ;
        RECT 5.8240 27.8235 5.8500 28.9170 ;
        RECT 5.7160 27.8235 5.7420 28.9170 ;
        RECT 5.6080 27.8235 5.6340 28.9170 ;
        RECT 5.5000 27.8235 5.5260 28.9170 ;
        RECT 5.3920 27.8235 5.4180 28.9170 ;
        RECT 5.2840 27.8235 5.3100 28.9170 ;
        RECT 5.1760 27.8235 5.2020 28.9170 ;
        RECT 5.0680 27.8235 5.0940 28.9170 ;
        RECT 4.9600 27.8235 4.9860 28.9170 ;
        RECT 4.8520 27.8235 4.8780 28.9170 ;
        RECT 4.7440 27.8235 4.7700 28.9170 ;
        RECT 4.6360 27.8235 4.6620 28.9170 ;
        RECT 4.5280 27.8235 4.5540 28.9170 ;
        RECT 4.4200 27.8235 4.4460 28.9170 ;
        RECT 4.3120 27.8235 4.3380 28.9170 ;
        RECT 4.2040 27.8235 4.2300 28.9170 ;
        RECT 4.0960 27.8235 4.1220 28.9170 ;
        RECT 3.9880 27.8235 4.0140 28.9170 ;
        RECT 3.8800 27.8235 3.9060 28.9170 ;
        RECT 3.7720 27.8235 3.7980 28.9170 ;
        RECT 3.6640 27.8235 3.6900 28.9170 ;
        RECT 3.5560 27.8235 3.5820 28.9170 ;
        RECT 3.4480 27.8235 3.4740 28.9170 ;
        RECT 3.3400 27.8235 3.3660 28.9170 ;
        RECT 3.2320 27.8235 3.2580 28.9170 ;
        RECT 3.1240 27.8235 3.1500 28.9170 ;
        RECT 3.0160 27.8235 3.0420 28.9170 ;
        RECT 2.9080 27.8235 2.9340 28.9170 ;
        RECT 2.8000 27.8235 2.8260 28.9170 ;
        RECT 2.6920 27.8235 2.7180 28.9170 ;
        RECT 2.5840 27.8235 2.6100 28.9170 ;
        RECT 2.4760 27.8235 2.5020 28.9170 ;
        RECT 2.3680 27.8235 2.3940 28.9170 ;
        RECT 2.2600 27.8235 2.2860 28.9170 ;
        RECT 2.1520 27.8235 2.1780 28.9170 ;
        RECT 2.0440 27.8235 2.0700 28.9170 ;
        RECT 1.9360 27.8235 1.9620 28.9170 ;
        RECT 1.8280 27.8235 1.8540 28.9170 ;
        RECT 1.7200 27.8235 1.7460 28.9170 ;
        RECT 1.6120 27.8235 1.6380 28.9170 ;
        RECT 1.5040 27.8235 1.5300 28.9170 ;
        RECT 1.3960 27.8235 1.4220 28.9170 ;
        RECT 1.2880 27.8235 1.3140 28.9170 ;
        RECT 1.1800 27.8235 1.2060 28.9170 ;
        RECT 1.0720 27.8235 1.0980 28.9170 ;
        RECT 0.9640 27.8235 0.9900 28.9170 ;
        RECT 0.8560 27.8235 0.8820 28.9170 ;
        RECT 0.7480 27.8235 0.7740 28.9170 ;
        RECT 0.6400 27.8235 0.6660 28.9170 ;
        RECT 0.5320 27.8235 0.5580 28.9170 ;
        RECT 0.4240 27.8235 0.4500 28.9170 ;
        RECT 0.3160 27.8235 0.3420 28.9170 ;
        RECT 0.2080 27.8235 0.2340 28.9170 ;
        RECT 0.0050 27.8235 0.0900 28.9170 ;
        RECT 8.6410 28.9035 8.7690 29.9970 ;
        RECT 8.6270 29.5690 8.7690 29.8915 ;
        RECT 8.4790 29.2960 8.5410 29.9970 ;
        RECT 8.4650 29.6055 8.5410 29.7590 ;
        RECT 8.4790 28.9035 8.5050 29.9970 ;
        RECT 8.4790 29.0245 8.5190 29.2640 ;
        RECT 8.4790 28.9035 8.5410 28.9925 ;
        RECT 8.1820 29.3540 8.3880 29.9970 ;
        RECT 8.3620 28.9035 8.3880 29.9970 ;
        RECT 8.1820 29.6310 8.4020 29.8890 ;
        RECT 8.1820 28.9035 8.2800 29.9970 ;
        RECT 7.7650 28.9035 7.8480 29.9970 ;
        RECT 7.7650 28.9920 7.8620 29.9275 ;
        RECT 16.4440 28.9035 16.5290 29.9970 ;
        RECT 16.3000 28.9035 16.3260 29.9970 ;
        RECT 16.1920 28.9035 16.2180 29.9970 ;
        RECT 16.0840 28.9035 16.1100 29.9970 ;
        RECT 15.9760 28.9035 16.0020 29.9970 ;
        RECT 15.8680 28.9035 15.8940 29.9970 ;
        RECT 15.7600 28.9035 15.7860 29.9970 ;
        RECT 15.6520 28.9035 15.6780 29.9970 ;
        RECT 15.5440 28.9035 15.5700 29.9970 ;
        RECT 15.4360 28.9035 15.4620 29.9970 ;
        RECT 15.3280 28.9035 15.3540 29.9970 ;
        RECT 15.2200 28.9035 15.2460 29.9970 ;
        RECT 15.1120 28.9035 15.1380 29.9970 ;
        RECT 15.0040 28.9035 15.0300 29.9970 ;
        RECT 14.8960 28.9035 14.9220 29.9970 ;
        RECT 14.7880 28.9035 14.8140 29.9970 ;
        RECT 14.6800 28.9035 14.7060 29.9970 ;
        RECT 14.5720 28.9035 14.5980 29.9970 ;
        RECT 14.4640 28.9035 14.4900 29.9970 ;
        RECT 14.3560 28.9035 14.3820 29.9970 ;
        RECT 14.2480 28.9035 14.2740 29.9970 ;
        RECT 14.1400 28.9035 14.1660 29.9970 ;
        RECT 14.0320 28.9035 14.0580 29.9970 ;
        RECT 13.9240 28.9035 13.9500 29.9970 ;
        RECT 13.8160 28.9035 13.8420 29.9970 ;
        RECT 13.7080 28.9035 13.7340 29.9970 ;
        RECT 13.6000 28.9035 13.6260 29.9970 ;
        RECT 13.4920 28.9035 13.5180 29.9970 ;
        RECT 13.3840 28.9035 13.4100 29.9970 ;
        RECT 13.2760 28.9035 13.3020 29.9970 ;
        RECT 13.1680 28.9035 13.1940 29.9970 ;
        RECT 13.0600 28.9035 13.0860 29.9970 ;
        RECT 12.9520 28.9035 12.9780 29.9970 ;
        RECT 12.8440 28.9035 12.8700 29.9970 ;
        RECT 12.7360 28.9035 12.7620 29.9970 ;
        RECT 12.6280 28.9035 12.6540 29.9970 ;
        RECT 12.5200 28.9035 12.5460 29.9970 ;
        RECT 12.4120 28.9035 12.4380 29.9970 ;
        RECT 12.3040 28.9035 12.3300 29.9970 ;
        RECT 12.1960 28.9035 12.2220 29.9970 ;
        RECT 12.0880 28.9035 12.1140 29.9970 ;
        RECT 11.9800 28.9035 12.0060 29.9970 ;
        RECT 11.8720 28.9035 11.8980 29.9970 ;
        RECT 11.7640 28.9035 11.7900 29.9970 ;
        RECT 11.6560 28.9035 11.6820 29.9970 ;
        RECT 11.5480 28.9035 11.5740 29.9970 ;
        RECT 11.4400 28.9035 11.4660 29.9970 ;
        RECT 11.3320 28.9035 11.3580 29.9970 ;
        RECT 11.2240 28.9035 11.2500 29.9970 ;
        RECT 11.1160 28.9035 11.1420 29.9970 ;
        RECT 11.0080 28.9035 11.0340 29.9970 ;
        RECT 10.9000 28.9035 10.9260 29.9970 ;
        RECT 10.7920 28.9035 10.8180 29.9970 ;
        RECT 10.6840 28.9035 10.7100 29.9970 ;
        RECT 10.5760 28.9035 10.6020 29.9970 ;
        RECT 10.4680 28.9035 10.4940 29.9970 ;
        RECT 10.3600 28.9035 10.3860 29.9970 ;
        RECT 10.2520 28.9035 10.2780 29.9970 ;
        RECT 10.1440 28.9035 10.1700 29.9970 ;
        RECT 10.0360 28.9035 10.0620 29.9970 ;
        RECT 9.9280 28.9035 9.9540 29.9970 ;
        RECT 9.8200 28.9035 9.8460 29.9970 ;
        RECT 9.7120 28.9035 9.7380 29.9970 ;
        RECT 9.6040 28.9035 9.6300 29.9970 ;
        RECT 9.4960 28.9035 9.5220 29.9970 ;
        RECT 9.3880 28.9035 9.4140 29.9970 ;
        RECT 9.1750 28.9035 9.2520 29.9970 ;
        RECT 7.2820 28.9035 7.3590 29.9970 ;
        RECT 7.1200 28.9035 7.1460 29.9970 ;
        RECT 7.0120 28.9035 7.0380 29.9970 ;
        RECT 6.9040 28.9035 6.9300 29.9970 ;
        RECT 6.7960 28.9035 6.8220 29.9970 ;
        RECT 6.6880 28.9035 6.7140 29.9970 ;
        RECT 6.5800 28.9035 6.6060 29.9970 ;
        RECT 6.4720 28.9035 6.4980 29.9970 ;
        RECT 6.3640 28.9035 6.3900 29.9970 ;
        RECT 6.2560 28.9035 6.2820 29.9970 ;
        RECT 6.1480 28.9035 6.1740 29.9970 ;
        RECT 6.0400 28.9035 6.0660 29.9970 ;
        RECT 5.9320 28.9035 5.9580 29.9970 ;
        RECT 5.8240 28.9035 5.8500 29.9970 ;
        RECT 5.7160 28.9035 5.7420 29.9970 ;
        RECT 5.6080 28.9035 5.6340 29.9970 ;
        RECT 5.5000 28.9035 5.5260 29.9970 ;
        RECT 5.3920 28.9035 5.4180 29.9970 ;
        RECT 5.2840 28.9035 5.3100 29.9970 ;
        RECT 5.1760 28.9035 5.2020 29.9970 ;
        RECT 5.0680 28.9035 5.0940 29.9970 ;
        RECT 4.9600 28.9035 4.9860 29.9970 ;
        RECT 4.8520 28.9035 4.8780 29.9970 ;
        RECT 4.7440 28.9035 4.7700 29.9970 ;
        RECT 4.6360 28.9035 4.6620 29.9970 ;
        RECT 4.5280 28.9035 4.5540 29.9970 ;
        RECT 4.4200 28.9035 4.4460 29.9970 ;
        RECT 4.3120 28.9035 4.3380 29.9970 ;
        RECT 4.2040 28.9035 4.2300 29.9970 ;
        RECT 4.0960 28.9035 4.1220 29.9970 ;
        RECT 3.9880 28.9035 4.0140 29.9970 ;
        RECT 3.8800 28.9035 3.9060 29.9970 ;
        RECT 3.7720 28.9035 3.7980 29.9970 ;
        RECT 3.6640 28.9035 3.6900 29.9970 ;
        RECT 3.5560 28.9035 3.5820 29.9970 ;
        RECT 3.4480 28.9035 3.4740 29.9970 ;
        RECT 3.3400 28.9035 3.3660 29.9970 ;
        RECT 3.2320 28.9035 3.2580 29.9970 ;
        RECT 3.1240 28.9035 3.1500 29.9970 ;
        RECT 3.0160 28.9035 3.0420 29.9970 ;
        RECT 2.9080 28.9035 2.9340 29.9970 ;
        RECT 2.8000 28.9035 2.8260 29.9970 ;
        RECT 2.6920 28.9035 2.7180 29.9970 ;
        RECT 2.5840 28.9035 2.6100 29.9970 ;
        RECT 2.4760 28.9035 2.5020 29.9970 ;
        RECT 2.3680 28.9035 2.3940 29.9970 ;
        RECT 2.2600 28.9035 2.2860 29.9970 ;
        RECT 2.1520 28.9035 2.1780 29.9970 ;
        RECT 2.0440 28.9035 2.0700 29.9970 ;
        RECT 1.9360 28.9035 1.9620 29.9970 ;
        RECT 1.8280 28.9035 1.8540 29.9970 ;
        RECT 1.7200 28.9035 1.7460 29.9970 ;
        RECT 1.6120 28.9035 1.6380 29.9970 ;
        RECT 1.5040 28.9035 1.5300 29.9970 ;
        RECT 1.3960 28.9035 1.4220 29.9970 ;
        RECT 1.2880 28.9035 1.3140 29.9970 ;
        RECT 1.1800 28.9035 1.2060 29.9970 ;
        RECT 1.0720 28.9035 1.0980 29.9970 ;
        RECT 0.9640 28.9035 0.9900 29.9970 ;
        RECT 0.8560 28.9035 0.8820 29.9970 ;
        RECT 0.7480 28.9035 0.7740 29.9970 ;
        RECT 0.6400 28.9035 0.6660 29.9970 ;
        RECT 0.5320 28.9035 0.5580 29.9970 ;
        RECT 0.4240 28.9035 0.4500 29.9970 ;
        RECT 0.3160 28.9035 0.3420 29.9970 ;
        RECT 0.2080 28.9035 0.2340 29.9970 ;
        RECT 0.0050 28.9035 0.0900 29.9970 ;
  LAYER V3 SPACING 0.018  ;
      RECT 0.0050 1.2200 16.5290 1.3500 ;
      RECT 16.4120 0.2565 16.5290 1.3500 ;
      RECT 9.3020 1.1240 16.3940 1.3500 ;
      RECT 7.9700 1.1240 9.2840 1.3500 ;
      RECT 7.2500 0.2565 7.8800 1.3500 ;
      RECT 0.1400 1.1240 7.2320 1.3500 ;
      RECT 0.0050 0.2565 0.1220 1.3500 ;
      RECT 16.3760 0.2565 16.5290 1.1720 ;
      RECT 9.3560 0.2565 16.3580 1.3500 ;
      RECT 8.6090 0.2565 9.3380 1.1720 ;
      RECT 8.4470 0.4520 8.5730 1.3500 ;
      RECT 7.1960 0.3560 8.4200 1.1720 ;
      RECT 0.1760 0.2565 7.1780 1.3500 ;
      RECT 0.0050 0.2565 0.1580 1.1720 ;
      RECT 8.5550 0.2565 16.5290 1.0760 ;
      RECT 0.0050 0.3560 8.5370 1.0760 ;
      RECT 8.3300 0.2565 16.5290 0.4280 ;
      RECT 0.0050 0.2565 8.3120 1.0760 ;
      RECT 0.0050 0.2565 16.5290 0.3320 ;
      RECT 0.0050 2.3000 16.5290 2.4300 ;
      RECT 16.4120 1.3365 16.5290 2.4300 ;
      RECT 9.3020 2.2040 16.3940 2.4300 ;
      RECT 7.9700 2.2040 9.2840 2.4300 ;
      RECT 7.2500 1.3365 7.8800 2.4300 ;
      RECT 0.1400 2.2040 7.2320 2.4300 ;
      RECT 0.0050 1.3365 0.1220 2.4300 ;
      RECT 16.3760 1.3365 16.5290 2.2520 ;
      RECT 9.3560 1.3365 16.3580 2.4300 ;
      RECT 8.6090 1.3365 9.3380 2.2520 ;
      RECT 8.4470 1.5320 8.5730 2.4300 ;
      RECT 7.1960 1.4360 8.4200 2.2520 ;
      RECT 0.1760 1.3365 7.1780 2.4300 ;
      RECT 0.0050 1.3365 0.1580 2.2520 ;
      RECT 8.5550 1.3365 16.5290 2.1560 ;
      RECT 0.0050 1.4360 8.5370 2.1560 ;
      RECT 8.3300 1.3365 16.5290 1.5080 ;
      RECT 0.0050 1.3365 8.3120 2.1560 ;
      RECT 0.0050 1.3365 16.5290 1.4120 ;
      RECT 0.0050 3.3800 16.5290 3.5100 ;
      RECT 16.4120 2.4165 16.5290 3.5100 ;
      RECT 9.3020 3.2840 16.3940 3.5100 ;
      RECT 7.9700 3.2840 9.2840 3.5100 ;
      RECT 7.2500 2.4165 7.8800 3.5100 ;
      RECT 0.1400 3.2840 7.2320 3.5100 ;
      RECT 0.0050 2.4165 0.1220 3.5100 ;
      RECT 16.3760 2.4165 16.5290 3.3320 ;
      RECT 9.3560 2.4165 16.3580 3.5100 ;
      RECT 8.6090 2.4165 9.3380 3.3320 ;
      RECT 8.4470 2.6120 8.5730 3.5100 ;
      RECT 7.1960 2.5160 8.4200 3.3320 ;
      RECT 0.1760 2.4165 7.1780 3.5100 ;
      RECT 0.0050 2.4165 0.1580 3.3320 ;
      RECT 8.5550 2.4165 16.5290 3.2360 ;
      RECT 0.0050 2.5160 8.5370 3.2360 ;
      RECT 8.3300 2.4165 16.5290 2.5880 ;
      RECT 0.0050 2.4165 8.3120 3.2360 ;
      RECT 0.0050 2.4165 16.5290 2.4920 ;
      RECT 0.0050 4.4600 16.5290 4.5900 ;
      RECT 16.4120 3.4965 16.5290 4.5900 ;
      RECT 9.3020 4.3640 16.3940 4.5900 ;
      RECT 7.9700 4.3640 9.2840 4.5900 ;
      RECT 7.2500 3.4965 7.8800 4.5900 ;
      RECT 0.1400 4.3640 7.2320 4.5900 ;
      RECT 0.0050 3.4965 0.1220 4.5900 ;
      RECT 16.3760 3.4965 16.5290 4.4120 ;
      RECT 9.3560 3.4965 16.3580 4.5900 ;
      RECT 8.6090 3.4965 9.3380 4.4120 ;
      RECT 8.4470 3.6920 8.5730 4.5900 ;
      RECT 7.1960 3.5960 8.4200 4.4120 ;
      RECT 0.1760 3.4965 7.1780 4.5900 ;
      RECT 0.0050 3.4965 0.1580 4.4120 ;
      RECT 8.5550 3.4965 16.5290 4.3160 ;
      RECT 0.0050 3.5960 8.5370 4.3160 ;
      RECT 8.3300 3.4965 16.5290 3.6680 ;
      RECT 0.0050 3.4965 8.3120 4.3160 ;
      RECT 0.0050 3.4965 16.5290 3.5720 ;
      RECT 0.0050 5.5400 16.5290 5.6700 ;
      RECT 16.4120 4.5765 16.5290 5.6700 ;
      RECT 9.3020 5.4440 16.3940 5.6700 ;
      RECT 7.9700 5.4440 9.2840 5.6700 ;
      RECT 7.2500 4.5765 7.8800 5.6700 ;
      RECT 0.1400 5.4440 7.2320 5.6700 ;
      RECT 0.0050 4.5765 0.1220 5.6700 ;
      RECT 16.3760 4.5765 16.5290 5.4920 ;
      RECT 9.3560 4.5765 16.3580 5.6700 ;
      RECT 8.6090 4.5765 9.3380 5.4920 ;
      RECT 8.4470 4.7720 8.5730 5.6700 ;
      RECT 7.1960 4.6760 8.4200 5.4920 ;
      RECT 0.1760 4.5765 7.1780 5.6700 ;
      RECT 0.0050 4.5765 0.1580 5.4920 ;
      RECT 8.5550 4.5765 16.5290 5.3960 ;
      RECT 0.0050 4.6760 8.5370 5.3960 ;
      RECT 8.3300 4.5765 16.5290 4.7480 ;
      RECT 0.0050 4.5765 8.3120 5.3960 ;
      RECT 0.0050 4.5765 16.5290 4.6520 ;
      RECT 0.0050 6.6200 16.5290 6.7500 ;
      RECT 16.4120 5.6565 16.5290 6.7500 ;
      RECT 9.3020 6.5240 16.3940 6.7500 ;
      RECT 7.9700 6.5240 9.2840 6.7500 ;
      RECT 7.2500 5.6565 7.8800 6.7500 ;
      RECT 0.1400 6.5240 7.2320 6.7500 ;
      RECT 0.0050 5.6565 0.1220 6.7500 ;
      RECT 16.3760 5.6565 16.5290 6.5720 ;
      RECT 9.3560 5.6565 16.3580 6.7500 ;
      RECT 8.6090 5.6565 9.3380 6.5720 ;
      RECT 8.4470 5.8520 8.5730 6.7500 ;
      RECT 7.1960 5.7560 8.4200 6.5720 ;
      RECT 0.1760 5.6565 7.1780 6.7500 ;
      RECT 0.0050 5.6565 0.1580 6.5720 ;
      RECT 8.5550 5.6565 16.5290 6.4760 ;
      RECT 0.0050 5.7560 8.5370 6.4760 ;
      RECT 8.3300 5.6565 16.5290 5.8280 ;
      RECT 0.0050 5.6565 8.3120 6.4760 ;
      RECT 0.0050 5.6565 16.5290 5.7320 ;
      RECT 0.0050 7.7000 16.5290 7.8300 ;
      RECT 16.4120 6.7365 16.5290 7.8300 ;
      RECT 9.3020 7.6040 16.3940 7.8300 ;
      RECT 7.9700 7.6040 9.2840 7.8300 ;
      RECT 7.2500 6.7365 7.8800 7.8300 ;
      RECT 0.1400 7.6040 7.2320 7.8300 ;
      RECT 0.0050 6.7365 0.1220 7.8300 ;
      RECT 16.3760 6.7365 16.5290 7.6520 ;
      RECT 9.3560 6.7365 16.3580 7.8300 ;
      RECT 8.6090 6.7365 9.3380 7.6520 ;
      RECT 8.4470 6.9320 8.5730 7.8300 ;
      RECT 7.1960 6.8360 8.4200 7.6520 ;
      RECT 0.1760 6.7365 7.1780 7.8300 ;
      RECT 0.0050 6.7365 0.1580 7.6520 ;
      RECT 8.5550 6.7365 16.5290 7.5560 ;
      RECT 0.0050 6.8360 8.5370 7.5560 ;
      RECT 8.3300 6.7365 16.5290 6.9080 ;
      RECT 0.0050 6.7365 8.3120 7.5560 ;
      RECT 0.0050 6.7365 16.5290 6.8120 ;
      RECT 0.0050 8.7800 16.5290 8.9100 ;
      RECT 16.4120 7.8165 16.5290 8.9100 ;
      RECT 9.3020 8.6840 16.3940 8.9100 ;
      RECT 7.9700 8.6840 9.2840 8.9100 ;
      RECT 7.2500 7.8165 7.8800 8.9100 ;
      RECT 0.1400 8.6840 7.2320 8.9100 ;
      RECT 0.0050 7.8165 0.1220 8.9100 ;
      RECT 16.3760 7.8165 16.5290 8.7320 ;
      RECT 9.3560 7.8165 16.3580 8.9100 ;
      RECT 8.6090 7.8165 9.3380 8.7320 ;
      RECT 8.4470 8.0120 8.5730 8.9100 ;
      RECT 7.1960 7.9160 8.4200 8.7320 ;
      RECT 0.1760 7.8165 7.1780 8.9100 ;
      RECT 0.0050 7.8165 0.1580 8.7320 ;
      RECT 8.5550 7.8165 16.5290 8.6360 ;
      RECT 0.0050 7.9160 8.5370 8.6360 ;
      RECT 8.3300 7.8165 16.5290 7.9880 ;
      RECT 0.0050 7.8165 8.3120 8.6360 ;
      RECT 0.0050 7.8165 16.5290 7.8920 ;
      RECT 0.0050 9.8600 16.5290 9.9900 ;
      RECT 16.4120 8.8965 16.5290 9.9900 ;
      RECT 9.3020 9.7640 16.3940 9.9900 ;
      RECT 7.9700 9.7640 9.2840 9.9900 ;
      RECT 7.2500 8.8965 7.8800 9.9900 ;
      RECT 0.1400 9.7640 7.2320 9.9900 ;
      RECT 0.0050 8.8965 0.1220 9.9900 ;
      RECT 16.3760 8.8965 16.5290 9.8120 ;
      RECT 9.3560 8.8965 16.3580 9.9900 ;
      RECT 8.6090 8.8965 9.3380 9.8120 ;
      RECT 8.4470 9.0920 8.5730 9.9900 ;
      RECT 7.1960 8.9960 8.4200 9.8120 ;
      RECT 0.1760 8.8965 7.1780 9.9900 ;
      RECT 0.0050 8.8965 0.1580 9.8120 ;
      RECT 8.5550 8.8965 16.5290 9.7160 ;
      RECT 0.0050 8.9960 8.5370 9.7160 ;
      RECT 8.3300 8.8965 16.5290 9.0680 ;
      RECT 0.0050 8.8965 8.3120 9.7160 ;
      RECT 0.0050 8.8965 16.5290 8.9720 ;
      RECT 0.0050 10.9400 16.5290 11.0700 ;
      RECT 16.4120 9.9765 16.5290 11.0700 ;
      RECT 9.3020 10.8440 16.3940 11.0700 ;
      RECT 7.9700 10.8440 9.2840 11.0700 ;
      RECT 7.2500 9.9765 7.8800 11.0700 ;
      RECT 0.1400 10.8440 7.2320 11.0700 ;
      RECT 0.0050 9.9765 0.1220 11.0700 ;
      RECT 16.3760 9.9765 16.5290 10.8920 ;
      RECT 9.3560 9.9765 16.3580 11.0700 ;
      RECT 8.6090 9.9765 9.3380 10.8920 ;
      RECT 8.4470 10.1720 8.5730 11.0700 ;
      RECT 7.1960 10.0760 8.4200 10.8920 ;
      RECT 0.1760 9.9765 7.1780 11.0700 ;
      RECT 0.0050 9.9765 0.1580 10.8920 ;
      RECT 8.5550 9.9765 16.5290 10.7960 ;
      RECT 0.0050 10.0760 8.5370 10.7960 ;
      RECT 8.3300 9.9765 16.5290 10.1480 ;
      RECT 0.0050 9.9765 8.3120 10.7960 ;
      RECT 0.0050 9.9765 16.5290 10.0520 ;
      RECT 0.0000 18.3570 16.5240 19.6905 ;
      RECT 10.8090 11.0370 16.5240 19.6905 ;
      RECT 8.6090 14.9010 16.5240 19.6905 ;
      RECT 9.5130 12.3090 16.5240 19.6905 ;
      RECT 8.5570 11.0370 8.5910 19.6905 ;
      RECT 8.5050 11.0370 8.5390 19.6905 ;
      RECT 8.4530 11.0370 8.4870 19.6905 ;
      RECT 8.4010 11.0370 8.4350 19.6905 ;
      RECT 0.0000 17.9250 8.3830 19.6905 ;
      RECT 8.1410 15.1890 16.5240 18.1410 ;
      RECT 8.0890 11.0370 8.1230 19.6905 ;
      RECT 8.0370 11.0370 8.0710 19.6905 ;
      RECT 7.9850 11.0370 8.0190 19.6905 ;
      RECT 7.9330 11.0370 7.9670 19.6905 ;
      RECT 0.0000 12.5970 7.9150 19.6905 ;
      RECT 0.0000 14.7570 8.3830 17.7090 ;
      RECT 8.1410 12.0210 9.2790 14.9730 ;
      RECT 9.3150 12.5010 16.5240 19.6905 ;
      RECT 0.0000 14.7570 9.2970 14.9730 ;
      RECT 8.1410 12.5010 16.5240 14.8770 ;
      RECT 7.4610 11.5890 8.2350 14.5410 ;
      RECT 7.2450 11.7330 7.9150 19.6905 ;
      RECT 0.0000 12.3090 7.2270 19.6905 ;
      RECT 6.8130 11.0370 7.2630 12.5730 ;
      RECT 0.0000 12.4050 9.4950 12.5730 ;
      RECT 9.2970 12.3090 16.5240 12.4770 ;
      RECT 10.5930 11.0370 10.7910 19.6905 ;
      RECT 6.8130 12.1170 10.5750 12.3810 ;
      RECT 5.9490 11.7330 6.7950 19.6905 ;
      RECT 0.0000 11.0370 5.9310 19.6905 ;
      RECT 10.3770 11.0370 16.5240 12.2850 ;
      RECT 10.1610 11.7330 16.5240 12.2850 ;
      RECT 0.0000 12.0215 10.1430 12.2850 ;
      RECT 9.9450 11.0370 10.3590 12.0930 ;
      RECT 9.3510 11.7330 16.5240 12.0930 ;
      RECT 8.6090 11.7330 9.3330 12.3810 ;
      RECT 8.1410 11.6850 8.3830 19.6905 ;
      RECT 8.2530 11.0370 8.6310 11.8050 ;
      RECT 8.6490 11.6850 9.9270 11.8055 ;
      RECT 6.5970 11.6850 7.4430 12.2850 ;
      RECT 6.1650 11.6850 6.5790 19.6905 ;
      RECT 0.0000 11.0370 6.1470 12.2850 ;
      RECT 9.7290 11.0370 16.5240 11.7090 ;
      RECT 8.2530 11.1170 9.7110 11.7090 ;
      RECT 7.2810 11.5890 8.2350 11.7090 ;
      RECT 6.3810 11.0370 7.2630 11.7090 ;
      RECT 0.0000 11.0370 6.3630 11.7090 ;
      RECT 9.2970 11.0370 16.5240 11.6610 ;
      RECT 8.1410 11.1170 16.5240 11.6610 ;
      RECT 0.0000 11.0370 7.9150 11.6610 ;
      RECT 0.0000 11.0370 9.2790 11.3730 ;
      RECT 0.0000 11.0370 16.5240 11.0930 ;
        RECT 0.0050 20.1470 16.5290 20.2770 ;
        RECT 16.4120 19.1835 16.5290 20.2770 ;
        RECT 9.3020 20.0510 16.3940 20.2770 ;
        RECT 7.9700 20.0510 9.2840 20.2770 ;
        RECT 7.2500 19.1835 7.8800 20.2770 ;
        RECT 0.1400 20.0510 7.2320 20.2770 ;
        RECT 0.0050 19.1835 0.1220 20.2770 ;
        RECT 16.3760 19.1835 16.5290 20.0990 ;
        RECT 9.3560 19.1835 16.3580 20.2770 ;
        RECT 8.6090 19.1835 9.3380 20.0990 ;
        RECT 8.4470 19.3790 8.5730 20.2770 ;
        RECT 7.1960 19.2830 8.4200 20.0990 ;
        RECT 0.1760 19.1835 7.1780 20.2770 ;
        RECT 0.0050 19.1835 0.1580 20.0990 ;
        RECT 8.5550 19.1835 16.5290 20.0030 ;
        RECT 0.0050 19.2830 8.5370 20.0030 ;
        RECT 8.3300 19.1835 16.5290 19.3550 ;
        RECT 0.0050 19.1835 8.3120 20.0030 ;
        RECT 0.0050 19.1835 16.5290 19.2590 ;
        RECT 0.0050 21.2270 16.5290 21.3570 ;
        RECT 16.4120 20.2635 16.5290 21.3570 ;
        RECT 9.3020 21.1310 16.3940 21.3570 ;
        RECT 7.9700 21.1310 9.2840 21.3570 ;
        RECT 7.2500 20.2635 7.8800 21.3570 ;
        RECT 0.1400 21.1310 7.2320 21.3570 ;
        RECT 0.0050 20.2635 0.1220 21.3570 ;
        RECT 16.3760 20.2635 16.5290 21.1790 ;
        RECT 9.3560 20.2635 16.3580 21.3570 ;
        RECT 8.6090 20.2635 9.3380 21.1790 ;
        RECT 8.4470 20.4590 8.5730 21.3570 ;
        RECT 7.1960 20.3630 8.4200 21.1790 ;
        RECT 0.1760 20.2635 7.1780 21.3570 ;
        RECT 0.0050 20.2635 0.1580 21.1790 ;
        RECT 8.5550 20.2635 16.5290 21.0830 ;
        RECT 0.0050 20.3630 8.5370 21.0830 ;
        RECT 8.3300 20.2635 16.5290 20.4350 ;
        RECT 0.0050 20.2635 8.3120 21.0830 ;
        RECT 0.0050 20.2635 16.5290 20.3390 ;
        RECT 0.0050 22.3070 16.5290 22.4370 ;
        RECT 16.4120 21.3435 16.5290 22.4370 ;
        RECT 9.3020 22.2110 16.3940 22.4370 ;
        RECT 7.9700 22.2110 9.2840 22.4370 ;
        RECT 7.2500 21.3435 7.8800 22.4370 ;
        RECT 0.1400 22.2110 7.2320 22.4370 ;
        RECT 0.0050 21.3435 0.1220 22.4370 ;
        RECT 16.3760 21.3435 16.5290 22.2590 ;
        RECT 9.3560 21.3435 16.3580 22.4370 ;
        RECT 8.6090 21.3435 9.3380 22.2590 ;
        RECT 8.4470 21.5390 8.5730 22.4370 ;
        RECT 7.1960 21.4430 8.4200 22.2590 ;
        RECT 0.1760 21.3435 7.1780 22.4370 ;
        RECT 0.0050 21.3435 0.1580 22.2590 ;
        RECT 8.5550 21.3435 16.5290 22.1630 ;
        RECT 0.0050 21.4430 8.5370 22.1630 ;
        RECT 8.3300 21.3435 16.5290 21.5150 ;
        RECT 0.0050 21.3435 8.3120 22.1630 ;
        RECT 0.0050 21.3435 16.5290 21.4190 ;
        RECT 0.0050 23.3870 16.5290 23.5170 ;
        RECT 16.4120 22.4235 16.5290 23.5170 ;
        RECT 9.3020 23.2910 16.3940 23.5170 ;
        RECT 7.9700 23.2910 9.2840 23.5170 ;
        RECT 7.2500 22.4235 7.8800 23.5170 ;
        RECT 0.1400 23.2910 7.2320 23.5170 ;
        RECT 0.0050 22.4235 0.1220 23.5170 ;
        RECT 16.3760 22.4235 16.5290 23.3390 ;
        RECT 9.3560 22.4235 16.3580 23.5170 ;
        RECT 8.6090 22.4235 9.3380 23.3390 ;
        RECT 8.4470 22.6190 8.5730 23.5170 ;
        RECT 7.1960 22.5230 8.4200 23.3390 ;
        RECT 0.1760 22.4235 7.1780 23.5170 ;
        RECT 0.0050 22.4235 0.1580 23.3390 ;
        RECT 8.5550 22.4235 16.5290 23.2430 ;
        RECT 0.0050 22.5230 8.5370 23.2430 ;
        RECT 8.3300 22.4235 16.5290 22.5950 ;
        RECT 0.0050 22.4235 8.3120 23.2430 ;
        RECT 0.0050 22.4235 16.5290 22.4990 ;
        RECT 0.0050 24.4670 16.5290 24.5970 ;
        RECT 16.4120 23.5035 16.5290 24.5970 ;
        RECT 9.3020 24.3710 16.3940 24.5970 ;
        RECT 7.9700 24.3710 9.2840 24.5970 ;
        RECT 7.2500 23.5035 7.8800 24.5970 ;
        RECT 0.1400 24.3710 7.2320 24.5970 ;
        RECT 0.0050 23.5035 0.1220 24.5970 ;
        RECT 16.3760 23.5035 16.5290 24.4190 ;
        RECT 9.3560 23.5035 16.3580 24.5970 ;
        RECT 8.6090 23.5035 9.3380 24.4190 ;
        RECT 8.4470 23.6990 8.5730 24.5970 ;
        RECT 7.1960 23.6030 8.4200 24.4190 ;
        RECT 0.1760 23.5035 7.1780 24.5970 ;
        RECT 0.0050 23.5035 0.1580 24.4190 ;
        RECT 8.5550 23.5035 16.5290 24.3230 ;
        RECT 0.0050 23.6030 8.5370 24.3230 ;
        RECT 8.3300 23.5035 16.5290 23.6750 ;
        RECT 0.0050 23.5035 8.3120 24.3230 ;
        RECT 0.0050 23.5035 16.5290 23.5790 ;
        RECT 0.0050 25.5470 16.5290 25.6770 ;
        RECT 16.4120 24.5835 16.5290 25.6770 ;
        RECT 9.3020 25.4510 16.3940 25.6770 ;
        RECT 7.9700 25.4510 9.2840 25.6770 ;
        RECT 7.2500 24.5835 7.8800 25.6770 ;
        RECT 0.1400 25.4510 7.2320 25.6770 ;
        RECT 0.0050 24.5835 0.1220 25.6770 ;
        RECT 16.3760 24.5835 16.5290 25.4990 ;
        RECT 9.3560 24.5835 16.3580 25.6770 ;
        RECT 8.6090 24.5835 9.3380 25.4990 ;
        RECT 8.4470 24.7790 8.5730 25.6770 ;
        RECT 7.1960 24.6830 8.4200 25.4990 ;
        RECT 0.1760 24.5835 7.1780 25.6770 ;
        RECT 0.0050 24.5835 0.1580 25.4990 ;
        RECT 8.5550 24.5835 16.5290 25.4030 ;
        RECT 0.0050 24.6830 8.5370 25.4030 ;
        RECT 8.3300 24.5835 16.5290 24.7550 ;
        RECT 0.0050 24.5835 8.3120 25.4030 ;
        RECT 0.0050 24.5835 16.5290 24.6590 ;
        RECT 0.0050 26.6270 16.5290 26.7570 ;
        RECT 16.4120 25.6635 16.5290 26.7570 ;
        RECT 9.3020 26.5310 16.3940 26.7570 ;
        RECT 7.9700 26.5310 9.2840 26.7570 ;
        RECT 7.2500 25.6635 7.8800 26.7570 ;
        RECT 0.1400 26.5310 7.2320 26.7570 ;
        RECT 0.0050 25.6635 0.1220 26.7570 ;
        RECT 16.3760 25.6635 16.5290 26.5790 ;
        RECT 9.3560 25.6635 16.3580 26.7570 ;
        RECT 8.6090 25.6635 9.3380 26.5790 ;
        RECT 8.4470 25.8590 8.5730 26.7570 ;
        RECT 7.1960 25.7630 8.4200 26.5790 ;
        RECT 0.1760 25.6635 7.1780 26.7570 ;
        RECT 0.0050 25.6635 0.1580 26.5790 ;
        RECT 8.5550 25.6635 16.5290 26.4830 ;
        RECT 0.0050 25.7630 8.5370 26.4830 ;
        RECT 8.3300 25.6635 16.5290 25.8350 ;
        RECT 0.0050 25.6635 8.3120 26.4830 ;
        RECT 0.0050 25.6635 16.5290 25.7390 ;
        RECT 0.0050 27.7070 16.5290 27.8370 ;
        RECT 16.4120 26.7435 16.5290 27.8370 ;
        RECT 9.3020 27.6110 16.3940 27.8370 ;
        RECT 7.9700 27.6110 9.2840 27.8370 ;
        RECT 7.2500 26.7435 7.8800 27.8370 ;
        RECT 0.1400 27.6110 7.2320 27.8370 ;
        RECT 0.0050 26.7435 0.1220 27.8370 ;
        RECT 16.3760 26.7435 16.5290 27.6590 ;
        RECT 9.3560 26.7435 16.3580 27.8370 ;
        RECT 8.6090 26.7435 9.3380 27.6590 ;
        RECT 8.4470 26.9390 8.5730 27.8370 ;
        RECT 7.1960 26.8430 8.4200 27.6590 ;
        RECT 0.1760 26.7435 7.1780 27.8370 ;
        RECT 0.0050 26.7435 0.1580 27.6590 ;
        RECT 8.5550 26.7435 16.5290 27.5630 ;
        RECT 0.0050 26.8430 8.5370 27.5630 ;
        RECT 8.3300 26.7435 16.5290 26.9150 ;
        RECT 0.0050 26.7435 8.3120 27.5630 ;
        RECT 0.0050 26.7435 16.5290 26.8190 ;
        RECT 0.0050 28.7870 16.5290 28.9170 ;
        RECT 16.4120 27.8235 16.5290 28.9170 ;
        RECT 9.3020 28.6910 16.3940 28.9170 ;
        RECT 7.9700 28.6910 9.2840 28.9170 ;
        RECT 7.2500 27.8235 7.8800 28.9170 ;
        RECT 0.1400 28.6910 7.2320 28.9170 ;
        RECT 0.0050 27.8235 0.1220 28.9170 ;
        RECT 16.3760 27.8235 16.5290 28.7390 ;
        RECT 9.3560 27.8235 16.3580 28.9170 ;
        RECT 8.6090 27.8235 9.3380 28.7390 ;
        RECT 8.4470 28.0190 8.5730 28.9170 ;
        RECT 7.1960 27.9230 8.4200 28.7390 ;
        RECT 0.1760 27.8235 7.1780 28.9170 ;
        RECT 0.0050 27.8235 0.1580 28.7390 ;
        RECT 8.5550 27.8235 16.5290 28.6430 ;
        RECT 0.0050 27.9230 8.5370 28.6430 ;
        RECT 8.3300 27.8235 16.5290 27.9950 ;
        RECT 0.0050 27.8235 8.3120 28.6430 ;
        RECT 0.0050 27.8235 16.5290 27.8990 ;
        RECT 0.0050 29.8670 16.5290 29.9970 ;
        RECT 16.4120 28.9035 16.5290 29.9970 ;
        RECT 9.3020 29.7710 16.3940 29.9970 ;
        RECT 7.9700 29.7710 9.2840 29.9970 ;
        RECT 7.2500 28.9035 7.8800 29.9970 ;
        RECT 0.1400 29.7710 7.2320 29.9970 ;
        RECT 0.0050 28.9035 0.1220 29.9970 ;
        RECT 16.3760 28.9035 16.5290 29.8190 ;
        RECT 9.3560 28.9035 16.3580 29.9970 ;
        RECT 8.6090 28.9035 9.3380 29.8190 ;
        RECT 8.4470 29.0990 8.5730 29.9970 ;
        RECT 7.1960 29.0030 8.4200 29.8190 ;
        RECT 0.1760 28.9035 7.1780 29.9970 ;
        RECT 0.0050 28.9035 0.1580 29.8190 ;
        RECT 8.5550 28.9035 16.5290 29.7230 ;
        RECT 0.0050 29.0030 8.5370 29.7230 ;
        RECT 8.3300 28.9035 16.5290 29.0750 ;
        RECT 0.0050 28.9035 8.3120 29.7230 ;
        RECT 0.0050 28.9035 16.5290 28.9790 ;
  LAYER M4  ;
      RECT 1.5690 12.7500 15.0095 12.7740 ;
      RECT 1.5690 13.0380 15.0095 13.0620 ;
      RECT 1.5690 13.4220 15.0095 13.4460 ;
      RECT 1.5690 13.5180 15.0095 13.5420 ;
      RECT 1.5690 13.8540 15.0095 13.8780 ;
      RECT 1.5690 14.2380 15.0095 14.2620 ;
      RECT 10.9550 11.7090 11.0390 11.7330 ;
      RECT 10.7670 12.1410 10.8970 12.1650 ;
      RECT 10.7750 12.7985 10.8920 12.8225 ;
      RECT 10.7750 13.0860 10.8920 13.1100 ;
      RECT 10.1360 12.1410 10.7070 12.1650 ;
      RECT 10.1960 12.9180 10.3040 12.9420 ;
      RECT 8.8630 13.2930 9.9560 13.3170 ;
      RECT 9.5510 12.8610 9.6350 12.8850 ;
      RECT 8.7670 14.0610 9.6350 14.0850 ;
      RECT 9.5510 14.1570 9.6350 14.1810 ;
      RECT 9.3730 12.3810 9.4570 12.4050 ;
      RECT 9.3350 13.7250 9.4190 13.7490 ;
      RECT 9.3350 14.4450 9.4190 14.4690 ;
      RECT 9.1570 12.2850 9.2410 12.3090 ;
      RECT 8.9430 10.9970 9.2060 11.0210 ;
      RECT 8.9430 19.6210 9.2060 19.6450 ;
      RECT 8.9590 13.7730 9.2030 13.7970 ;
      RECT 9.1190 13.9170 9.2030 13.9410 ;
      RECT 7.6630 14.1570 9.2030 14.1810 ;
      RECT 9.1190 14.4450 9.2030 14.4690 ;
      RECT 8.8850 19.5250 9.1480 19.5490 ;
      RECT 8.8840 10.9010 9.1470 10.9250 ;
      RECT 8.8460 10.8050 9.1090 10.8290 ;
      RECT 8.8460 19.3330 9.1090 19.3570 ;
      RECT 9.0110 14.8770 9.0950 14.9010 ;
      RECT 8.2390 15.2610 9.0950 15.2850 ;
      RECT 8.6230 17.5170 9.0950 17.5410 ;
      RECT 9.0110 17.6130 9.0950 17.6370 ;
      RECT 8.7980 10.7090 9.0610 10.7330 ;
      RECT 8.7980 19.2370 9.0610 19.2610 ;
      RECT 8.5750 16.6050 9.0200 16.6290 ;
      RECT 8.7540 10.6130 9.0170 10.6370 ;
      RECT 8.7540 19.5730 9.0170 19.5970 ;
      RECT 8.7050 10.9490 8.9680 10.9730 ;
      RECT 8.7050 19.4770 8.9680 19.5010 ;
      RECT 8.8360 13.9170 8.9570 13.9410 ;
      RECT 8.8150 16.0290 8.9480 16.0530 ;
      RECT 8.6580 10.8530 8.9210 10.8770 ;
      RECT 8.6580 19.3810 8.9210 19.4050 ;
      RECT 8.6230 10.5650 8.8860 10.5890 ;
      RECT 8.6230 19.2850 8.8860 19.3090 ;
      RECT 7.8070 17.6130 8.8760 17.6370 ;
      RECT 8.7920 18.7650 8.8760 18.7890 ;
      RECT 8.5670 10.4210 8.8300 10.4450 ;
      RECT 8.5670 19.1890 8.8300 19.2130 ;
      RECT 8.7190 14.8770 8.8040 14.9010 ;
      RECT 7.6150 15.4530 8.7320 15.4770 ;
      RECT 8.2600 13.2930 8.7170 13.3170 ;
      RECT 8.0870 11.1410 8.3540 11.1650 ;
      RECT 8.0870 19.0450 8.3540 19.0690 ;
      RECT 8.2240 14.8290 8.3330 14.8530 ;
      RECT 8.0640 11.0450 8.3060 11.0690 ;
      RECT 8.0640 19.6690 8.3060 19.6930 ;
      RECT 8.0080 10.5650 8.2500 10.5890 ;
      RECT 8.0370 19.7650 8.2500 19.7890 ;
      RECT 8.1530 14.4450 8.2370 14.4690 ;
      RECT 7.9540 10.6610 8.2020 10.6850 ;
      RECT 7.9540 19.6210 8.2020 19.6450 ;
      RECT 7.7200 17.0370 8.1410 17.0610 ;
      RECT 7.6880 10.9970 7.9550 11.0210 ;
      RECT 7.6880 19.7650 7.9550 19.7890 ;
      RECT 7.8280 15.5970 7.9490 15.6210 ;
      RECT 7.8200 18.7650 7.9040 18.7890 ;
      RECT 7.6540 10.9010 7.9010 10.9250 ;
      RECT 7.5870 19.3330 7.9010 19.3570 ;
      RECT 7.6280 10.8050 7.8580 10.8290 ;
      RECT 7.6160 19.6690 7.8580 19.6930 ;
      RECT 7.5750 10.7090 7.8050 10.7330 ;
      RECT 7.7210 17.1810 7.8050 17.2050 ;
      RECT 7.5250 19.2370 7.8050 19.2610 ;
      RECT 7.5300 10.6130 7.7600 10.6370 ;
      RECT 7.5300 19.5730 7.7600 19.5970 ;
      RECT 6.5680 14.4450 7.7570 14.4690 ;
      RECT 7.4920 10.8530 7.7220 10.8770 ;
      RECT 7.4920 19.4770 7.7220 19.5010 ;
      RECT 7.4740 10.7570 7.6670 10.7810 ;
      RECT 7.4740 19.3810 7.6670 19.4050 ;
      RECT 7.4250 10.6610 7.6180 10.6850 ;
      RECT 7.4250 19.2850 7.6180 19.3090 ;
      RECT 7.4290 15.3570 7.6130 15.3810 ;
      RECT 7.3730 10.5650 7.5660 10.5890 ;
      RECT 7.3730 19.1890 7.5660 19.2130 ;
      RECT 6.8890 12.6690 7.5650 12.6930 ;
      RECT 7.4290 15.4530 7.5130 15.4770 ;
      RECT 7.1600 11.0930 7.4230 11.1170 ;
      RECT 7.1925 14.8770 7.3260 14.9010 ;
      RECT 6.8510 12.8610 6.9350 12.8850 ;
  LAYER V4  ;
      RECT 11.0040 11.7090 11.0280 11.7330 ;
      RECT 11.0040 12.7500 11.0280 12.7740 ;
      RECT 10.8360 12.1410 10.8600 12.1650 ;
      RECT 10.8360 12.7985 10.8600 12.8225 ;
      RECT 10.8360 13.0860 10.8600 13.1100 ;
      RECT 10.2120 12.1410 10.2360 12.1650 ;
      RECT 10.2120 12.9180 10.2360 12.9420 ;
      RECT 9.6000 12.8610 9.6240 12.8850 ;
      RECT 9.6000 13.0380 9.6240 13.0620 ;
      RECT 9.6000 14.0610 9.6240 14.0850 ;
      RECT 9.6000 14.1570 9.6240 14.1810 ;
      RECT 9.3840 12.3810 9.4080 12.4050 ;
      RECT 9.3840 13.4220 9.4080 13.4460 ;
      RECT 9.3840 13.7250 9.4080 13.7490 ;
      RECT 9.3840 13.8540 9.4080 13.8780 ;
      RECT 9.3840 14.2380 9.4080 14.2620 ;
      RECT 9.3840 14.4450 9.4080 14.4690 ;
      RECT 9.1680 12.2850 9.1920 12.3090 ;
      RECT 9.1680 13.5180 9.1920 13.5420 ;
      RECT 9.1680 13.7730 9.1920 13.7970 ;
      RECT 9.1680 13.9170 9.1920 13.9410 ;
      RECT 9.1680 14.1570 9.1920 14.1810 ;
      RECT 9.1680 14.4450 9.1920 14.4690 ;
      RECT 9.0600 14.8770 9.0840 14.9010 ;
      RECT 9.0600 15.2610 9.0840 15.2850 ;
      RECT 9.0600 17.5170 9.0840 17.5410 ;
      RECT 9.0600 17.6130 9.0840 17.6370 ;
      RECT 8.9700 10.9970 8.9940 11.0210 ;
      RECT 8.9700 13.7730 8.9940 13.7970 ;
      RECT 8.9700 19.6210 8.9940 19.6450 ;
      RECT 8.9220 10.9010 8.9460 10.9250 ;
      RECT 8.9220 13.9170 8.9460 13.9410 ;
      RECT 8.9220 19.5250 8.9460 19.5490 ;
      RECT 8.8740 10.8050 8.8980 10.8290 ;
      RECT 8.8740 13.2930 8.8980 13.3170 ;
      RECT 8.8740 19.3330 8.8980 19.3570 ;
      RECT 8.8260 10.7090 8.8500 10.7330 ;
      RECT 8.8260 16.0290 8.8500 16.0530 ;
      RECT 8.8260 18.7650 8.8500 18.7890 ;
      RECT 8.8260 19.2370 8.8500 19.2610 ;
      RECT 8.7780 10.6130 8.8020 10.6370 ;
      RECT 8.7780 14.0610 8.8020 14.0850 ;
      RECT 8.7780 19.5730 8.8020 19.5970 ;
      RECT 8.7300 10.9490 8.7540 10.9730 ;
      RECT 8.7300 14.8770 8.7540 14.9010 ;
      RECT 8.7300 19.4770 8.7540 19.5010 ;
      RECT 8.6820 10.8530 8.7060 10.8770 ;
      RECT 8.6820 13.2930 8.7060 13.3170 ;
      RECT 8.6820 19.3810 8.7060 19.4050 ;
      RECT 8.6340 10.5650 8.6580 10.5890 ;
      RECT 8.6340 17.5170 8.6580 17.5410 ;
      RECT 8.6340 19.2850 8.6580 19.3090 ;
      RECT 8.5860 10.4210 8.6100 10.4450 ;
      RECT 8.5860 16.6050 8.6100 16.6290 ;
      RECT 8.5860 19.1890 8.6100 19.2130 ;
      RECT 8.2980 11.1410 8.3220 11.1650 ;
      RECT 8.2980 14.8290 8.3220 14.8530 ;
      RECT 8.2980 19.0450 8.3220 19.0690 ;
      RECT 8.2500 11.0450 8.2740 11.0690 ;
      RECT 8.2500 15.2610 8.2740 15.2850 ;
      RECT 8.2500 19.6690 8.2740 19.6930 ;
      RECT 8.2020 10.5650 8.2260 10.5890 ;
      RECT 8.2020 14.4450 8.2260 14.4690 ;
      RECT 8.2020 19.7650 8.2260 19.7890 ;
      RECT 8.1060 10.6610 8.1300 10.6850 ;
      RECT 8.1060 17.0370 8.1300 17.0610 ;
      RECT 8.1060 19.6210 8.1300 19.6450 ;
      RECT 7.9140 10.9970 7.9380 11.0210 ;
      RECT 7.9140 15.5970 7.9380 15.6210 ;
      RECT 7.9140 19.7650 7.9380 19.7890 ;
      RECT 7.8660 10.9010 7.8900 10.9250 ;
      RECT 7.8660 18.7650 7.8900 18.7890 ;
      RECT 7.8660 19.3330 7.8900 19.3570 ;
      RECT 7.8180 10.8050 7.8420 10.8290 ;
      RECT 7.8180 17.6130 7.8420 17.6370 ;
      RECT 7.8180 19.6690 7.8420 19.6930 ;
      RECT 7.7700 10.7090 7.7940 10.7330 ;
      RECT 7.7700 17.1810 7.7940 17.2050 ;
      RECT 7.7700 19.2370 7.7940 19.2610 ;
      RECT 7.7220 10.6130 7.7460 10.6370 ;
      RECT 7.7220 14.4450 7.7460 14.4690 ;
      RECT 7.7220 19.5730 7.7460 19.5970 ;
      RECT 7.6740 10.8530 7.6980 10.8770 ;
      RECT 7.6740 14.1570 7.6980 14.1810 ;
      RECT 7.6740 19.4770 7.6980 19.5010 ;
      RECT 7.6260 10.7570 7.6500 10.7810 ;
      RECT 7.6260 15.4530 7.6500 15.4770 ;
      RECT 7.6260 19.3810 7.6500 19.4050 ;
      RECT 7.5780 10.6610 7.6020 10.6850 ;
      RECT 7.5780 15.3570 7.6020 15.3810 ;
      RECT 7.5780 19.2850 7.6020 19.3090 ;
      RECT 7.5300 10.5650 7.5540 10.5890 ;
      RECT 7.5300 12.6690 7.5540 12.6930 ;
      RECT 7.5300 19.1890 7.5540 19.2130 ;
      RECT 7.4400 15.3570 7.4640 15.3810 ;
      RECT 7.4400 15.4530 7.4640 15.4770 ;
      RECT 7.2720 11.0930 7.2960 11.1170 ;
      RECT 7.2720 14.8770 7.2960 14.9010 ;
      RECT 6.9000 12.6690 6.9240 12.6930 ;
      RECT 6.9000 12.8610 6.9240 12.8850 ;
  LAYER M5  ;
      RECT 11.0040 11.6980 11.0280 12.7850 ;
      RECT 10.8360 12.1130 10.8600 13.1735 ;
      RECT 10.2120 12.1215 10.2360 12.9540 ;
      RECT 9.6000 12.8500 9.6240 13.0730 ;
      RECT 9.6000 14.0500 9.6240 14.1920 ;
      RECT 9.3840 12.3700 9.4080 13.4570 ;
      RECT 9.3840 13.7140 9.4080 13.8890 ;
      RECT 9.3840 14.2270 9.4080 14.4800 ;
      RECT 9.1680 12.2740 9.1920 13.5530 ;
      RECT 9.1680 13.7620 9.1920 13.9520 ;
      RECT 9.1680 14.1460 9.1920 14.4800 ;
      RECT 9.0600 14.8660 9.0840 15.2960 ;
      RECT 9.0600 17.5060 9.0840 17.6480 ;
      RECT 8.9700 11.3340 8.9940 18.9170 ;
      RECT 8.9220 11.3340 8.9460 18.9170 ;
      RECT 8.8740 11.3340 8.8980 18.9170 ;
      RECT 8.8260 11.3340 8.8500 18.9170 ;
      RECT 8.7780 11.3340 8.8020 18.9170 ;
      RECT 8.7300 11.3340 8.7540 18.9170 ;
      RECT 8.6820 11.3340 8.7060 18.9170 ;
      RECT 8.6340 11.3340 8.6580 18.9170 ;
      RECT 8.5860 11.3340 8.6100 18.9170 ;
      RECT 8.2980 11.3340 8.3220 18.9170 ;
      RECT 8.2500 11.3340 8.2740 18.9170 ;
      RECT 8.2020 11.3340 8.2260 18.9170 ;
      RECT 8.1060 11.3340 8.1300 18.9170 ;
      RECT 7.9140 11.3340 7.9380 18.9170 ;
      RECT 7.8660 11.3340 7.8900 18.9170 ;
      RECT 7.8180 11.3340 7.8420 18.9170 ;
      RECT 7.7700 11.3340 7.7940 18.9170 ;
      RECT 7.7220 11.3340 7.7460 18.9170 ;
      RECT 7.6740 11.3340 7.6980 18.9170 ;
      RECT 7.6260 10.4920 7.6500 19.5470 ;
      RECT 7.5780 10.4550 7.6020 19.5010 ;
      RECT 7.5300 10.4010 7.5540 19.4470 ;
      RECT 7.4400 15.3460 7.4640 15.4880 ;
      RECT 7.2720 11.0750 7.2960 14.9190 ;
      RECT 6.9000 12.6580 6.9240 12.8960 ;
  LAYER M2  ;
    RECT 0.108 0.036 15.8920 30.2040 ;
  LAYER M1  ;
    RECT 0.108 0.036 15.8920 30.2040 ;
  END
END srambank_128x4x20_6t122 
