VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_128x4x74_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_128x4x74_6t122 0 0 ; 
  SIZE 64 BY 354.24 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.688 65.768 4.88 ; 
        RECT 0.376 9.008 65.768 9.2 ; 
        RECT 0.376 13.328 65.768 13.52 ; 
        RECT 0.376 17.648 65.768 17.84 ; 
        RECT 0.376 21.968 65.768 22.16 ; 
        RECT 0.376 26.288 65.768 26.48 ; 
        RECT 0.376 30.608 65.768 30.8 ; 
        RECT 0.376 34.928 65.768 35.12 ; 
        RECT 0.376 39.248 65.768 39.44 ; 
        RECT 0.376 43.568 65.768 43.76 ; 
        RECT 0.376 47.888 65.768 48.08 ; 
        RECT 0.376 52.208 65.768 52.4 ; 
        RECT 0.376 56.528 65.768 56.72 ; 
        RECT 0.376 60.848 65.768 61.04 ; 
        RECT 0.376 65.168 65.768 65.36 ; 
        RECT 0.376 69.488 65.768 69.68 ; 
        RECT 0.376 73.808 65.768 74 ; 
        RECT 0.376 78.128 65.768 78.32 ; 
        RECT 0.376 82.448 65.768 82.64 ; 
        RECT 0.376 86.768 65.768 86.96 ; 
        RECT 0.376 91.088 65.768 91.28 ; 
        RECT 0.376 95.408 65.768 95.6 ; 
        RECT 0.376 99.728 65.768 99.92 ; 
        RECT 0.376 104.048 65.768 104.24 ; 
        RECT 0.376 108.368 65.768 108.56 ; 
        RECT 0.376 112.688 65.768 112.88 ; 
        RECT 0.376 117.008 65.768 117.2 ; 
        RECT 0.376 121.328 65.768 121.52 ; 
        RECT 0.376 125.648 65.768 125.84 ; 
        RECT 0.376 129.968 65.768 130.16 ; 
        RECT 0.376 134.288 65.768 134.48 ; 
        RECT 0.376 138.608 65.768 138.8 ; 
        RECT 0.376 142.928 65.768 143.12 ; 
        RECT 0.376 147.248 65.768 147.44 ; 
        RECT 0.376 151.568 65.768 151.76 ; 
        RECT 0.376 155.888 65.768 156.08 ; 
        RECT 0.376 160.208 65.768 160.4 ; 
        RECT 14.256 162.132 51.84 162.996 ; 
        RECT 36.788 176.148 37.352 176.244 ; 
        RECT 36.264 161.012 37.316 161.108 ; 
        RECT 29.592 174.804 36.504 175.668 ; 
        RECT 29.592 187.476 36.504 188.34 ; 
        RECT 0.376 197.036 65.768 197.228 ; 
        RECT 0.376 201.356 65.768 201.548 ; 
        RECT 0.376 205.676 65.768 205.868 ; 
        RECT 0.376 209.996 65.768 210.188 ; 
        RECT 0.376 214.316 65.768 214.508 ; 
        RECT 0.376 218.636 65.768 218.828 ; 
        RECT 0.376 222.956 65.768 223.148 ; 
        RECT 0.376 227.276 65.768 227.468 ; 
        RECT 0.376 231.596 65.768 231.788 ; 
        RECT 0.376 235.916 65.768 236.108 ; 
        RECT 0.376 240.236 65.768 240.428 ; 
        RECT 0.376 244.556 65.768 244.748 ; 
        RECT 0.376 248.876 65.768 249.068 ; 
        RECT 0.376 253.196 65.768 253.388 ; 
        RECT 0.376 257.516 65.768 257.708 ; 
        RECT 0.376 261.836 65.768 262.028 ; 
        RECT 0.376 266.156 65.768 266.348 ; 
        RECT 0.376 270.476 65.768 270.668 ; 
        RECT 0.376 274.796 65.768 274.988 ; 
        RECT 0.376 279.116 65.768 279.308 ; 
        RECT 0.376 283.436 65.768 283.628 ; 
        RECT 0.376 287.756 65.768 287.948 ; 
        RECT 0.376 292.076 65.768 292.268 ; 
        RECT 0.376 296.396 65.768 296.588 ; 
        RECT 0.376 300.716 65.768 300.908 ; 
        RECT 0.376 305.036 65.768 305.228 ; 
        RECT 0.376 309.356 65.768 309.548 ; 
        RECT 0.376 313.676 65.768 313.868 ; 
        RECT 0.376 317.996 65.768 318.188 ; 
        RECT 0.376 322.316 65.768 322.508 ; 
        RECT 0.376 326.636 65.768 326.828 ; 
        RECT 0.376 330.956 65.768 331.148 ; 
        RECT 0.376 335.276 65.768 335.468 ; 
        RECT 0.376 339.596 65.768 339.788 ; 
        RECT 0.376 343.916 65.768 344.108 ; 
        RECT 0.376 348.236 65.768 348.428 ; 
        RECT 0.376 352.556 65.768 352.748 ; 
      LAYER M3 ; 
        RECT 65.576 0.866 65.648 5.506 ; 
        RECT 37.136 0.868 37.208 5.504 ; 
        RECT 31.52 1.028 31.88 5.484 ; 
        RECT 28.928 0.868 29 5.504 ; 
        RECT 0.488 0.866 0.56 5.506 ; 
        RECT 65.576 5.186 65.648 9.826 ; 
        RECT 37.136 5.188 37.208 9.824 ; 
        RECT 31.52 5.348 31.88 9.804 ; 
        RECT 28.928 5.188 29 9.824 ; 
        RECT 0.488 5.186 0.56 9.826 ; 
        RECT 65.576 9.506 65.648 14.146 ; 
        RECT 37.136 9.508 37.208 14.144 ; 
        RECT 31.52 9.668 31.88 14.124 ; 
        RECT 28.928 9.508 29 14.144 ; 
        RECT 0.488 9.506 0.56 14.146 ; 
        RECT 65.576 13.826 65.648 18.466 ; 
        RECT 37.136 13.828 37.208 18.464 ; 
        RECT 31.52 13.988 31.88 18.444 ; 
        RECT 28.928 13.828 29 18.464 ; 
        RECT 0.488 13.826 0.56 18.466 ; 
        RECT 65.576 18.146 65.648 22.786 ; 
        RECT 37.136 18.148 37.208 22.784 ; 
        RECT 31.52 18.308 31.88 22.764 ; 
        RECT 28.928 18.148 29 22.784 ; 
        RECT 0.488 18.146 0.56 22.786 ; 
        RECT 65.576 22.466 65.648 27.106 ; 
        RECT 37.136 22.468 37.208 27.104 ; 
        RECT 31.52 22.628 31.88 27.084 ; 
        RECT 28.928 22.468 29 27.104 ; 
        RECT 0.488 22.466 0.56 27.106 ; 
        RECT 65.576 26.786 65.648 31.426 ; 
        RECT 37.136 26.788 37.208 31.424 ; 
        RECT 31.52 26.948 31.88 31.404 ; 
        RECT 28.928 26.788 29 31.424 ; 
        RECT 0.488 26.786 0.56 31.426 ; 
        RECT 65.576 31.106 65.648 35.746 ; 
        RECT 37.136 31.108 37.208 35.744 ; 
        RECT 31.52 31.268 31.88 35.724 ; 
        RECT 28.928 31.108 29 35.744 ; 
        RECT 0.488 31.106 0.56 35.746 ; 
        RECT 65.576 35.426 65.648 40.066 ; 
        RECT 37.136 35.428 37.208 40.064 ; 
        RECT 31.52 35.588 31.88 40.044 ; 
        RECT 28.928 35.428 29 40.064 ; 
        RECT 0.488 35.426 0.56 40.066 ; 
        RECT 65.576 39.746 65.648 44.386 ; 
        RECT 37.136 39.748 37.208 44.384 ; 
        RECT 31.52 39.908 31.88 44.364 ; 
        RECT 28.928 39.748 29 44.384 ; 
        RECT 0.488 39.746 0.56 44.386 ; 
        RECT 65.576 44.066 65.648 48.706 ; 
        RECT 37.136 44.068 37.208 48.704 ; 
        RECT 31.52 44.228 31.88 48.684 ; 
        RECT 28.928 44.068 29 48.704 ; 
        RECT 0.488 44.066 0.56 48.706 ; 
        RECT 65.576 48.386 65.648 53.026 ; 
        RECT 37.136 48.388 37.208 53.024 ; 
        RECT 31.52 48.548 31.88 53.004 ; 
        RECT 28.928 48.388 29 53.024 ; 
        RECT 0.488 48.386 0.56 53.026 ; 
        RECT 65.576 52.706 65.648 57.346 ; 
        RECT 37.136 52.708 37.208 57.344 ; 
        RECT 31.52 52.868 31.88 57.324 ; 
        RECT 28.928 52.708 29 57.344 ; 
        RECT 0.488 52.706 0.56 57.346 ; 
        RECT 65.576 57.026 65.648 61.666 ; 
        RECT 37.136 57.028 37.208 61.664 ; 
        RECT 31.52 57.188 31.88 61.644 ; 
        RECT 28.928 57.028 29 61.664 ; 
        RECT 0.488 57.026 0.56 61.666 ; 
        RECT 65.576 61.346 65.648 65.986 ; 
        RECT 37.136 61.348 37.208 65.984 ; 
        RECT 31.52 61.508 31.88 65.964 ; 
        RECT 28.928 61.348 29 65.984 ; 
        RECT 0.488 61.346 0.56 65.986 ; 
        RECT 65.576 65.666 65.648 70.306 ; 
        RECT 37.136 65.668 37.208 70.304 ; 
        RECT 31.52 65.828 31.88 70.284 ; 
        RECT 28.928 65.668 29 70.304 ; 
        RECT 0.488 65.666 0.56 70.306 ; 
        RECT 65.576 69.986 65.648 74.626 ; 
        RECT 37.136 69.988 37.208 74.624 ; 
        RECT 31.52 70.148 31.88 74.604 ; 
        RECT 28.928 69.988 29 74.624 ; 
        RECT 0.488 69.986 0.56 74.626 ; 
        RECT 65.576 74.306 65.648 78.946 ; 
        RECT 37.136 74.308 37.208 78.944 ; 
        RECT 31.52 74.468 31.88 78.924 ; 
        RECT 28.928 74.308 29 78.944 ; 
        RECT 0.488 74.306 0.56 78.946 ; 
        RECT 65.576 78.626 65.648 83.266 ; 
        RECT 37.136 78.628 37.208 83.264 ; 
        RECT 31.52 78.788 31.88 83.244 ; 
        RECT 28.928 78.628 29 83.264 ; 
        RECT 0.488 78.626 0.56 83.266 ; 
        RECT 65.576 82.946 65.648 87.586 ; 
        RECT 37.136 82.948 37.208 87.584 ; 
        RECT 31.52 83.108 31.88 87.564 ; 
        RECT 28.928 82.948 29 87.584 ; 
        RECT 0.488 82.946 0.56 87.586 ; 
        RECT 65.576 87.266 65.648 91.906 ; 
        RECT 37.136 87.268 37.208 91.904 ; 
        RECT 31.52 87.428 31.88 91.884 ; 
        RECT 28.928 87.268 29 91.904 ; 
        RECT 0.488 87.266 0.56 91.906 ; 
        RECT 65.576 91.586 65.648 96.226 ; 
        RECT 37.136 91.588 37.208 96.224 ; 
        RECT 31.52 91.748 31.88 96.204 ; 
        RECT 28.928 91.588 29 96.224 ; 
        RECT 0.488 91.586 0.56 96.226 ; 
        RECT 65.576 95.906 65.648 100.546 ; 
        RECT 37.136 95.908 37.208 100.544 ; 
        RECT 31.52 96.068 31.88 100.524 ; 
        RECT 28.928 95.908 29 100.544 ; 
        RECT 0.488 95.906 0.56 100.546 ; 
        RECT 65.576 100.226 65.648 104.866 ; 
        RECT 37.136 100.228 37.208 104.864 ; 
        RECT 31.52 100.388 31.88 104.844 ; 
        RECT 28.928 100.228 29 104.864 ; 
        RECT 0.488 100.226 0.56 104.866 ; 
        RECT 65.576 104.546 65.648 109.186 ; 
        RECT 37.136 104.548 37.208 109.184 ; 
        RECT 31.52 104.708 31.88 109.164 ; 
        RECT 28.928 104.548 29 109.184 ; 
        RECT 0.488 104.546 0.56 109.186 ; 
        RECT 65.576 108.866 65.648 113.506 ; 
        RECT 37.136 108.868 37.208 113.504 ; 
        RECT 31.52 109.028 31.88 113.484 ; 
        RECT 28.928 108.868 29 113.504 ; 
        RECT 0.488 108.866 0.56 113.506 ; 
        RECT 65.576 113.186 65.648 117.826 ; 
        RECT 37.136 113.188 37.208 117.824 ; 
        RECT 31.52 113.348 31.88 117.804 ; 
        RECT 28.928 113.188 29 117.824 ; 
        RECT 0.488 113.186 0.56 117.826 ; 
        RECT 65.576 117.506 65.648 122.146 ; 
        RECT 37.136 117.508 37.208 122.144 ; 
        RECT 31.52 117.668 31.88 122.124 ; 
        RECT 28.928 117.508 29 122.144 ; 
        RECT 0.488 117.506 0.56 122.146 ; 
        RECT 65.576 121.826 65.648 126.466 ; 
        RECT 37.136 121.828 37.208 126.464 ; 
        RECT 31.52 121.988 31.88 126.444 ; 
        RECT 28.928 121.828 29 126.464 ; 
        RECT 0.488 121.826 0.56 126.466 ; 
        RECT 65.576 126.146 65.648 130.786 ; 
        RECT 37.136 126.148 37.208 130.784 ; 
        RECT 31.52 126.308 31.88 130.764 ; 
        RECT 28.928 126.148 29 130.784 ; 
        RECT 0.488 126.146 0.56 130.786 ; 
        RECT 65.576 130.466 65.648 135.106 ; 
        RECT 37.136 130.468 37.208 135.104 ; 
        RECT 31.52 130.628 31.88 135.084 ; 
        RECT 28.928 130.468 29 135.104 ; 
        RECT 0.488 130.466 0.56 135.106 ; 
        RECT 65.576 134.786 65.648 139.426 ; 
        RECT 37.136 134.788 37.208 139.424 ; 
        RECT 31.52 134.948 31.88 139.404 ; 
        RECT 28.928 134.788 29 139.424 ; 
        RECT 0.488 134.786 0.56 139.426 ; 
        RECT 65.576 139.106 65.648 143.746 ; 
        RECT 37.136 139.108 37.208 143.744 ; 
        RECT 31.52 139.268 31.88 143.724 ; 
        RECT 28.928 139.108 29 143.744 ; 
        RECT 0.488 139.106 0.56 143.746 ; 
        RECT 65.576 143.426 65.648 148.066 ; 
        RECT 37.136 143.428 37.208 148.064 ; 
        RECT 31.52 143.588 31.88 148.044 ; 
        RECT 28.928 143.428 29 148.064 ; 
        RECT 0.488 143.426 0.56 148.066 ; 
        RECT 65.576 147.746 65.648 152.386 ; 
        RECT 37.136 147.748 37.208 152.384 ; 
        RECT 31.52 147.908 31.88 152.364 ; 
        RECT 28.928 147.748 29 152.384 ; 
        RECT 0.488 147.746 0.56 152.386 ; 
        RECT 65.576 152.066 65.648 156.706 ; 
        RECT 37.136 152.068 37.208 156.704 ; 
        RECT 31.52 152.228 31.88 156.684 ; 
        RECT 28.928 152.068 29 156.704 ; 
        RECT 0.488 152.066 0.56 156.706 ; 
        RECT 65.576 156.386 65.648 161.026 ; 
        RECT 37.136 156.388 37.208 161.024 ; 
        RECT 31.52 156.548 31.88 161.004 ; 
        RECT 28.928 156.388 29 161.024 ; 
        RECT 0.488 156.386 0.56 161.026 ; 
        RECT 65.556 160.682 65.628 193.51 ; 
        RECT 37.188 175.96 37.26 193.354 ; 
        RECT 37.116 160.814 37.188 161.366 ; 
        RECT 31.644 161.976 32.58 192.308 ; 
        RECT 31.5 191.976 31.86 193.48 ; 
        RECT 31.5 160.84 31.86 162.344 ; 
        RECT 0.468 160.682 0.54 193.51 ; 
        RECT 65.576 193.214 65.648 197.854 ; 
        RECT 37.136 193.216 37.208 197.852 ; 
        RECT 31.52 193.376 31.88 197.832 ; 
        RECT 28.928 193.216 29 197.852 ; 
        RECT 0.488 193.214 0.56 197.854 ; 
        RECT 65.576 197.534 65.648 202.174 ; 
        RECT 37.136 197.536 37.208 202.172 ; 
        RECT 31.52 197.696 31.88 202.152 ; 
        RECT 28.928 197.536 29 202.172 ; 
        RECT 0.488 197.534 0.56 202.174 ; 
        RECT 65.576 201.854 65.648 206.494 ; 
        RECT 37.136 201.856 37.208 206.492 ; 
        RECT 31.52 202.016 31.88 206.472 ; 
        RECT 28.928 201.856 29 206.492 ; 
        RECT 0.488 201.854 0.56 206.494 ; 
        RECT 65.576 206.174 65.648 210.814 ; 
        RECT 37.136 206.176 37.208 210.812 ; 
        RECT 31.52 206.336 31.88 210.792 ; 
        RECT 28.928 206.176 29 210.812 ; 
        RECT 0.488 206.174 0.56 210.814 ; 
        RECT 65.576 210.494 65.648 215.134 ; 
        RECT 37.136 210.496 37.208 215.132 ; 
        RECT 31.52 210.656 31.88 215.112 ; 
        RECT 28.928 210.496 29 215.132 ; 
        RECT 0.488 210.494 0.56 215.134 ; 
        RECT 65.576 214.814 65.648 219.454 ; 
        RECT 37.136 214.816 37.208 219.452 ; 
        RECT 31.52 214.976 31.88 219.432 ; 
        RECT 28.928 214.816 29 219.452 ; 
        RECT 0.488 214.814 0.56 219.454 ; 
        RECT 65.576 219.134 65.648 223.774 ; 
        RECT 37.136 219.136 37.208 223.772 ; 
        RECT 31.52 219.296 31.88 223.752 ; 
        RECT 28.928 219.136 29 223.772 ; 
        RECT 0.488 219.134 0.56 223.774 ; 
        RECT 65.576 223.454 65.648 228.094 ; 
        RECT 37.136 223.456 37.208 228.092 ; 
        RECT 31.52 223.616 31.88 228.072 ; 
        RECT 28.928 223.456 29 228.092 ; 
        RECT 0.488 223.454 0.56 228.094 ; 
        RECT 65.576 227.774 65.648 232.414 ; 
        RECT 37.136 227.776 37.208 232.412 ; 
        RECT 31.52 227.936 31.88 232.392 ; 
        RECT 28.928 227.776 29 232.412 ; 
        RECT 0.488 227.774 0.56 232.414 ; 
        RECT 65.576 232.094 65.648 236.734 ; 
        RECT 37.136 232.096 37.208 236.732 ; 
        RECT 31.52 232.256 31.88 236.712 ; 
        RECT 28.928 232.096 29 236.732 ; 
        RECT 0.488 232.094 0.56 236.734 ; 
        RECT 65.576 236.414 65.648 241.054 ; 
        RECT 37.136 236.416 37.208 241.052 ; 
        RECT 31.52 236.576 31.88 241.032 ; 
        RECT 28.928 236.416 29 241.052 ; 
        RECT 0.488 236.414 0.56 241.054 ; 
        RECT 65.576 240.734 65.648 245.374 ; 
        RECT 37.136 240.736 37.208 245.372 ; 
        RECT 31.52 240.896 31.88 245.352 ; 
        RECT 28.928 240.736 29 245.372 ; 
        RECT 0.488 240.734 0.56 245.374 ; 
        RECT 65.576 245.054 65.648 249.694 ; 
        RECT 37.136 245.056 37.208 249.692 ; 
        RECT 31.52 245.216 31.88 249.672 ; 
        RECT 28.928 245.056 29 249.692 ; 
        RECT 0.488 245.054 0.56 249.694 ; 
        RECT 65.576 249.374 65.648 254.014 ; 
        RECT 37.136 249.376 37.208 254.012 ; 
        RECT 31.52 249.536 31.88 253.992 ; 
        RECT 28.928 249.376 29 254.012 ; 
        RECT 0.488 249.374 0.56 254.014 ; 
        RECT 65.576 253.694 65.648 258.334 ; 
        RECT 37.136 253.696 37.208 258.332 ; 
        RECT 31.52 253.856 31.88 258.312 ; 
        RECT 28.928 253.696 29 258.332 ; 
        RECT 0.488 253.694 0.56 258.334 ; 
        RECT 65.576 258.014 65.648 262.654 ; 
        RECT 37.136 258.016 37.208 262.652 ; 
        RECT 31.52 258.176 31.88 262.632 ; 
        RECT 28.928 258.016 29 262.652 ; 
        RECT 0.488 258.014 0.56 262.654 ; 
        RECT 65.576 262.334 65.648 266.974 ; 
        RECT 37.136 262.336 37.208 266.972 ; 
        RECT 31.52 262.496 31.88 266.952 ; 
        RECT 28.928 262.336 29 266.972 ; 
        RECT 0.488 262.334 0.56 266.974 ; 
        RECT 65.576 266.654 65.648 271.294 ; 
        RECT 37.136 266.656 37.208 271.292 ; 
        RECT 31.52 266.816 31.88 271.272 ; 
        RECT 28.928 266.656 29 271.292 ; 
        RECT 0.488 266.654 0.56 271.294 ; 
        RECT 65.576 270.974 65.648 275.614 ; 
        RECT 37.136 270.976 37.208 275.612 ; 
        RECT 31.52 271.136 31.88 275.592 ; 
        RECT 28.928 270.976 29 275.612 ; 
        RECT 0.488 270.974 0.56 275.614 ; 
        RECT 65.576 275.294 65.648 279.934 ; 
        RECT 37.136 275.296 37.208 279.932 ; 
        RECT 31.52 275.456 31.88 279.912 ; 
        RECT 28.928 275.296 29 279.932 ; 
        RECT 0.488 275.294 0.56 279.934 ; 
        RECT 65.576 279.614 65.648 284.254 ; 
        RECT 37.136 279.616 37.208 284.252 ; 
        RECT 31.52 279.776 31.88 284.232 ; 
        RECT 28.928 279.616 29 284.252 ; 
        RECT 0.488 279.614 0.56 284.254 ; 
        RECT 65.576 283.934 65.648 288.574 ; 
        RECT 37.136 283.936 37.208 288.572 ; 
        RECT 31.52 284.096 31.88 288.552 ; 
        RECT 28.928 283.936 29 288.572 ; 
        RECT 0.488 283.934 0.56 288.574 ; 
        RECT 65.576 288.254 65.648 292.894 ; 
        RECT 37.136 288.256 37.208 292.892 ; 
        RECT 31.52 288.416 31.88 292.872 ; 
        RECT 28.928 288.256 29 292.892 ; 
        RECT 0.488 288.254 0.56 292.894 ; 
        RECT 65.576 292.574 65.648 297.214 ; 
        RECT 37.136 292.576 37.208 297.212 ; 
        RECT 31.52 292.736 31.88 297.192 ; 
        RECT 28.928 292.576 29 297.212 ; 
        RECT 0.488 292.574 0.56 297.214 ; 
        RECT 65.576 296.894 65.648 301.534 ; 
        RECT 37.136 296.896 37.208 301.532 ; 
        RECT 31.52 297.056 31.88 301.512 ; 
        RECT 28.928 296.896 29 301.532 ; 
        RECT 0.488 296.894 0.56 301.534 ; 
        RECT 65.576 301.214 65.648 305.854 ; 
        RECT 37.136 301.216 37.208 305.852 ; 
        RECT 31.52 301.376 31.88 305.832 ; 
        RECT 28.928 301.216 29 305.852 ; 
        RECT 0.488 301.214 0.56 305.854 ; 
        RECT 65.576 305.534 65.648 310.174 ; 
        RECT 37.136 305.536 37.208 310.172 ; 
        RECT 31.52 305.696 31.88 310.152 ; 
        RECT 28.928 305.536 29 310.172 ; 
        RECT 0.488 305.534 0.56 310.174 ; 
        RECT 65.576 309.854 65.648 314.494 ; 
        RECT 37.136 309.856 37.208 314.492 ; 
        RECT 31.52 310.016 31.88 314.472 ; 
        RECT 28.928 309.856 29 314.492 ; 
        RECT 0.488 309.854 0.56 314.494 ; 
        RECT 65.576 314.174 65.648 318.814 ; 
        RECT 37.136 314.176 37.208 318.812 ; 
        RECT 31.52 314.336 31.88 318.792 ; 
        RECT 28.928 314.176 29 318.812 ; 
        RECT 0.488 314.174 0.56 318.814 ; 
        RECT 65.576 318.494 65.648 323.134 ; 
        RECT 37.136 318.496 37.208 323.132 ; 
        RECT 31.52 318.656 31.88 323.112 ; 
        RECT 28.928 318.496 29 323.132 ; 
        RECT 0.488 318.494 0.56 323.134 ; 
        RECT 65.576 322.814 65.648 327.454 ; 
        RECT 37.136 322.816 37.208 327.452 ; 
        RECT 31.52 322.976 31.88 327.432 ; 
        RECT 28.928 322.816 29 327.452 ; 
        RECT 0.488 322.814 0.56 327.454 ; 
        RECT 65.576 327.134 65.648 331.774 ; 
        RECT 37.136 327.136 37.208 331.772 ; 
        RECT 31.52 327.296 31.88 331.752 ; 
        RECT 28.928 327.136 29 331.772 ; 
        RECT 0.488 327.134 0.56 331.774 ; 
        RECT 65.576 331.454 65.648 336.094 ; 
        RECT 37.136 331.456 37.208 336.092 ; 
        RECT 31.52 331.616 31.88 336.072 ; 
        RECT 28.928 331.456 29 336.092 ; 
        RECT 0.488 331.454 0.56 336.094 ; 
        RECT 65.576 335.774 65.648 340.414 ; 
        RECT 37.136 335.776 37.208 340.412 ; 
        RECT 31.52 335.936 31.88 340.392 ; 
        RECT 28.928 335.776 29 340.412 ; 
        RECT 0.488 335.774 0.56 340.414 ; 
        RECT 65.576 340.094 65.648 344.734 ; 
        RECT 37.136 340.096 37.208 344.732 ; 
        RECT 31.52 340.256 31.88 344.712 ; 
        RECT 28.928 340.096 29 344.732 ; 
        RECT 0.488 340.094 0.56 344.734 ; 
        RECT 65.576 344.414 65.648 349.054 ; 
        RECT 37.136 344.416 37.208 349.052 ; 
        RECT 31.52 344.576 31.88 349.032 ; 
        RECT 28.928 344.416 29 349.052 ; 
        RECT 0.488 344.414 0.56 349.054 ; 
        RECT 65.576 348.734 65.648 353.374 ; 
        RECT 37.136 348.736 37.208 353.372 ; 
        RECT 31.52 348.896 31.88 353.352 ; 
        RECT 28.928 348.736 29 353.372 ; 
        RECT 0.488 348.734 0.56 353.374 ; 
      LAYER V3 ; 
        RECT 0.488 4.688 0.56 4.88 ; 
        RECT 28.928 4.688 29 4.88 ; 
        RECT 31.52 4.688 31.88 4.88 ; 
        RECT 37.136 4.688 37.208 4.88 ; 
        RECT 65.576 4.688 65.648 4.88 ; 
        RECT 0.488 9.008 0.56 9.2 ; 
        RECT 28.928 9.008 29 9.2 ; 
        RECT 31.52 9.008 31.88 9.2 ; 
        RECT 37.136 9.008 37.208 9.2 ; 
        RECT 65.576 9.008 65.648 9.2 ; 
        RECT 0.488 13.328 0.56 13.52 ; 
        RECT 28.928 13.328 29 13.52 ; 
        RECT 31.52 13.328 31.88 13.52 ; 
        RECT 37.136 13.328 37.208 13.52 ; 
        RECT 65.576 13.328 65.648 13.52 ; 
        RECT 0.488 17.648 0.56 17.84 ; 
        RECT 28.928 17.648 29 17.84 ; 
        RECT 31.52 17.648 31.88 17.84 ; 
        RECT 37.136 17.648 37.208 17.84 ; 
        RECT 65.576 17.648 65.648 17.84 ; 
        RECT 0.488 21.968 0.56 22.16 ; 
        RECT 28.928 21.968 29 22.16 ; 
        RECT 31.52 21.968 31.88 22.16 ; 
        RECT 37.136 21.968 37.208 22.16 ; 
        RECT 65.576 21.968 65.648 22.16 ; 
        RECT 0.488 26.288 0.56 26.48 ; 
        RECT 28.928 26.288 29 26.48 ; 
        RECT 31.52 26.288 31.88 26.48 ; 
        RECT 37.136 26.288 37.208 26.48 ; 
        RECT 65.576 26.288 65.648 26.48 ; 
        RECT 0.488 30.608 0.56 30.8 ; 
        RECT 28.928 30.608 29 30.8 ; 
        RECT 31.52 30.608 31.88 30.8 ; 
        RECT 37.136 30.608 37.208 30.8 ; 
        RECT 65.576 30.608 65.648 30.8 ; 
        RECT 0.488 34.928 0.56 35.12 ; 
        RECT 28.928 34.928 29 35.12 ; 
        RECT 31.52 34.928 31.88 35.12 ; 
        RECT 37.136 34.928 37.208 35.12 ; 
        RECT 65.576 34.928 65.648 35.12 ; 
        RECT 0.488 39.248 0.56 39.44 ; 
        RECT 28.928 39.248 29 39.44 ; 
        RECT 31.52 39.248 31.88 39.44 ; 
        RECT 37.136 39.248 37.208 39.44 ; 
        RECT 65.576 39.248 65.648 39.44 ; 
        RECT 0.488 43.568 0.56 43.76 ; 
        RECT 28.928 43.568 29 43.76 ; 
        RECT 31.52 43.568 31.88 43.76 ; 
        RECT 37.136 43.568 37.208 43.76 ; 
        RECT 65.576 43.568 65.648 43.76 ; 
        RECT 0.488 47.888 0.56 48.08 ; 
        RECT 28.928 47.888 29 48.08 ; 
        RECT 31.52 47.888 31.88 48.08 ; 
        RECT 37.136 47.888 37.208 48.08 ; 
        RECT 65.576 47.888 65.648 48.08 ; 
        RECT 0.488 52.208 0.56 52.4 ; 
        RECT 28.928 52.208 29 52.4 ; 
        RECT 31.52 52.208 31.88 52.4 ; 
        RECT 37.136 52.208 37.208 52.4 ; 
        RECT 65.576 52.208 65.648 52.4 ; 
        RECT 0.488 56.528 0.56 56.72 ; 
        RECT 28.928 56.528 29 56.72 ; 
        RECT 31.52 56.528 31.88 56.72 ; 
        RECT 37.136 56.528 37.208 56.72 ; 
        RECT 65.576 56.528 65.648 56.72 ; 
        RECT 0.488 60.848 0.56 61.04 ; 
        RECT 28.928 60.848 29 61.04 ; 
        RECT 31.52 60.848 31.88 61.04 ; 
        RECT 37.136 60.848 37.208 61.04 ; 
        RECT 65.576 60.848 65.648 61.04 ; 
        RECT 0.488 65.168 0.56 65.36 ; 
        RECT 28.928 65.168 29 65.36 ; 
        RECT 31.52 65.168 31.88 65.36 ; 
        RECT 37.136 65.168 37.208 65.36 ; 
        RECT 65.576 65.168 65.648 65.36 ; 
        RECT 0.488 69.488 0.56 69.68 ; 
        RECT 28.928 69.488 29 69.68 ; 
        RECT 31.52 69.488 31.88 69.68 ; 
        RECT 37.136 69.488 37.208 69.68 ; 
        RECT 65.576 69.488 65.648 69.68 ; 
        RECT 0.488 73.808 0.56 74 ; 
        RECT 28.928 73.808 29 74 ; 
        RECT 31.52 73.808 31.88 74 ; 
        RECT 37.136 73.808 37.208 74 ; 
        RECT 65.576 73.808 65.648 74 ; 
        RECT 0.488 78.128 0.56 78.32 ; 
        RECT 28.928 78.128 29 78.32 ; 
        RECT 31.52 78.128 31.88 78.32 ; 
        RECT 37.136 78.128 37.208 78.32 ; 
        RECT 65.576 78.128 65.648 78.32 ; 
        RECT 0.488 82.448 0.56 82.64 ; 
        RECT 28.928 82.448 29 82.64 ; 
        RECT 31.52 82.448 31.88 82.64 ; 
        RECT 37.136 82.448 37.208 82.64 ; 
        RECT 65.576 82.448 65.648 82.64 ; 
        RECT 0.488 86.768 0.56 86.96 ; 
        RECT 28.928 86.768 29 86.96 ; 
        RECT 31.52 86.768 31.88 86.96 ; 
        RECT 37.136 86.768 37.208 86.96 ; 
        RECT 65.576 86.768 65.648 86.96 ; 
        RECT 0.488 91.088 0.56 91.28 ; 
        RECT 28.928 91.088 29 91.28 ; 
        RECT 31.52 91.088 31.88 91.28 ; 
        RECT 37.136 91.088 37.208 91.28 ; 
        RECT 65.576 91.088 65.648 91.28 ; 
        RECT 0.488 95.408 0.56 95.6 ; 
        RECT 28.928 95.408 29 95.6 ; 
        RECT 31.52 95.408 31.88 95.6 ; 
        RECT 37.136 95.408 37.208 95.6 ; 
        RECT 65.576 95.408 65.648 95.6 ; 
        RECT 0.488 99.728 0.56 99.92 ; 
        RECT 28.928 99.728 29 99.92 ; 
        RECT 31.52 99.728 31.88 99.92 ; 
        RECT 37.136 99.728 37.208 99.92 ; 
        RECT 65.576 99.728 65.648 99.92 ; 
        RECT 0.488 104.048 0.56 104.24 ; 
        RECT 28.928 104.048 29 104.24 ; 
        RECT 31.52 104.048 31.88 104.24 ; 
        RECT 37.136 104.048 37.208 104.24 ; 
        RECT 65.576 104.048 65.648 104.24 ; 
        RECT 0.488 108.368 0.56 108.56 ; 
        RECT 28.928 108.368 29 108.56 ; 
        RECT 31.52 108.368 31.88 108.56 ; 
        RECT 37.136 108.368 37.208 108.56 ; 
        RECT 65.576 108.368 65.648 108.56 ; 
        RECT 0.488 112.688 0.56 112.88 ; 
        RECT 28.928 112.688 29 112.88 ; 
        RECT 31.52 112.688 31.88 112.88 ; 
        RECT 37.136 112.688 37.208 112.88 ; 
        RECT 65.576 112.688 65.648 112.88 ; 
        RECT 0.488 117.008 0.56 117.2 ; 
        RECT 28.928 117.008 29 117.2 ; 
        RECT 31.52 117.008 31.88 117.2 ; 
        RECT 37.136 117.008 37.208 117.2 ; 
        RECT 65.576 117.008 65.648 117.2 ; 
        RECT 0.488 121.328 0.56 121.52 ; 
        RECT 28.928 121.328 29 121.52 ; 
        RECT 31.52 121.328 31.88 121.52 ; 
        RECT 37.136 121.328 37.208 121.52 ; 
        RECT 65.576 121.328 65.648 121.52 ; 
        RECT 0.488 125.648 0.56 125.84 ; 
        RECT 28.928 125.648 29 125.84 ; 
        RECT 31.52 125.648 31.88 125.84 ; 
        RECT 37.136 125.648 37.208 125.84 ; 
        RECT 65.576 125.648 65.648 125.84 ; 
        RECT 0.488 129.968 0.56 130.16 ; 
        RECT 28.928 129.968 29 130.16 ; 
        RECT 31.52 129.968 31.88 130.16 ; 
        RECT 37.136 129.968 37.208 130.16 ; 
        RECT 65.576 129.968 65.648 130.16 ; 
        RECT 0.488 134.288 0.56 134.48 ; 
        RECT 28.928 134.288 29 134.48 ; 
        RECT 31.52 134.288 31.88 134.48 ; 
        RECT 37.136 134.288 37.208 134.48 ; 
        RECT 65.576 134.288 65.648 134.48 ; 
        RECT 0.488 138.608 0.56 138.8 ; 
        RECT 28.928 138.608 29 138.8 ; 
        RECT 31.52 138.608 31.88 138.8 ; 
        RECT 37.136 138.608 37.208 138.8 ; 
        RECT 65.576 138.608 65.648 138.8 ; 
        RECT 0.488 142.928 0.56 143.12 ; 
        RECT 28.928 142.928 29 143.12 ; 
        RECT 31.52 142.928 31.88 143.12 ; 
        RECT 37.136 142.928 37.208 143.12 ; 
        RECT 65.576 142.928 65.648 143.12 ; 
        RECT 0.488 147.248 0.56 147.44 ; 
        RECT 28.928 147.248 29 147.44 ; 
        RECT 31.52 147.248 31.88 147.44 ; 
        RECT 37.136 147.248 37.208 147.44 ; 
        RECT 65.576 147.248 65.648 147.44 ; 
        RECT 0.488 151.568 0.56 151.76 ; 
        RECT 28.928 151.568 29 151.76 ; 
        RECT 31.52 151.568 31.88 151.76 ; 
        RECT 37.136 151.568 37.208 151.76 ; 
        RECT 65.576 151.568 65.648 151.76 ; 
        RECT 0.488 155.888 0.56 156.08 ; 
        RECT 28.928 155.888 29 156.08 ; 
        RECT 31.52 155.888 31.88 156.08 ; 
        RECT 37.136 155.888 37.208 156.08 ; 
        RECT 65.576 155.888 65.648 156.08 ; 
        RECT 0.488 160.208 0.56 160.4 ; 
        RECT 28.928 160.208 29 160.4 ; 
        RECT 31.52 160.208 31.88 160.4 ; 
        RECT 37.136 160.208 37.208 160.4 ; 
        RECT 65.576 160.208 65.648 160.4 ; 
        RECT 31.66 187.476 31.732 188.34 ; 
        RECT 31.66 174.804 31.732 175.668 ; 
        RECT 31.66 162.132 31.732 162.996 ; 
        RECT 31.868 187.476 31.94 188.34 ; 
        RECT 31.868 174.804 31.94 175.668 ; 
        RECT 31.868 162.132 31.94 162.996 ; 
        RECT 32.076 187.476 32.148 188.34 ; 
        RECT 32.076 174.804 32.148 175.668 ; 
        RECT 32.076 162.132 32.148 162.996 ; 
        RECT 32.284 187.476 32.356 188.34 ; 
        RECT 32.284 174.804 32.356 175.668 ; 
        RECT 32.284 162.132 32.356 162.996 ; 
        RECT 32.492 187.476 32.564 188.34 ; 
        RECT 32.492 174.804 32.564 175.668 ; 
        RECT 32.492 162.132 32.564 162.996 ; 
        RECT 37.116 161.012 37.188 161.108 ; 
        RECT 37.188 176.148 37.26 176.244 ; 
        RECT 0.488 197.036 0.56 197.228 ; 
        RECT 28.928 197.036 29 197.228 ; 
        RECT 31.52 197.036 31.88 197.228 ; 
        RECT 37.136 197.036 37.208 197.228 ; 
        RECT 65.576 197.036 65.648 197.228 ; 
        RECT 0.488 201.356 0.56 201.548 ; 
        RECT 28.928 201.356 29 201.548 ; 
        RECT 31.52 201.356 31.88 201.548 ; 
        RECT 37.136 201.356 37.208 201.548 ; 
        RECT 65.576 201.356 65.648 201.548 ; 
        RECT 0.488 205.676 0.56 205.868 ; 
        RECT 28.928 205.676 29 205.868 ; 
        RECT 31.52 205.676 31.88 205.868 ; 
        RECT 37.136 205.676 37.208 205.868 ; 
        RECT 65.576 205.676 65.648 205.868 ; 
        RECT 0.488 209.996 0.56 210.188 ; 
        RECT 28.928 209.996 29 210.188 ; 
        RECT 31.52 209.996 31.88 210.188 ; 
        RECT 37.136 209.996 37.208 210.188 ; 
        RECT 65.576 209.996 65.648 210.188 ; 
        RECT 0.488 214.316 0.56 214.508 ; 
        RECT 28.928 214.316 29 214.508 ; 
        RECT 31.52 214.316 31.88 214.508 ; 
        RECT 37.136 214.316 37.208 214.508 ; 
        RECT 65.576 214.316 65.648 214.508 ; 
        RECT 0.488 218.636 0.56 218.828 ; 
        RECT 28.928 218.636 29 218.828 ; 
        RECT 31.52 218.636 31.88 218.828 ; 
        RECT 37.136 218.636 37.208 218.828 ; 
        RECT 65.576 218.636 65.648 218.828 ; 
        RECT 0.488 222.956 0.56 223.148 ; 
        RECT 28.928 222.956 29 223.148 ; 
        RECT 31.52 222.956 31.88 223.148 ; 
        RECT 37.136 222.956 37.208 223.148 ; 
        RECT 65.576 222.956 65.648 223.148 ; 
        RECT 0.488 227.276 0.56 227.468 ; 
        RECT 28.928 227.276 29 227.468 ; 
        RECT 31.52 227.276 31.88 227.468 ; 
        RECT 37.136 227.276 37.208 227.468 ; 
        RECT 65.576 227.276 65.648 227.468 ; 
        RECT 0.488 231.596 0.56 231.788 ; 
        RECT 28.928 231.596 29 231.788 ; 
        RECT 31.52 231.596 31.88 231.788 ; 
        RECT 37.136 231.596 37.208 231.788 ; 
        RECT 65.576 231.596 65.648 231.788 ; 
        RECT 0.488 235.916 0.56 236.108 ; 
        RECT 28.928 235.916 29 236.108 ; 
        RECT 31.52 235.916 31.88 236.108 ; 
        RECT 37.136 235.916 37.208 236.108 ; 
        RECT 65.576 235.916 65.648 236.108 ; 
        RECT 0.488 240.236 0.56 240.428 ; 
        RECT 28.928 240.236 29 240.428 ; 
        RECT 31.52 240.236 31.88 240.428 ; 
        RECT 37.136 240.236 37.208 240.428 ; 
        RECT 65.576 240.236 65.648 240.428 ; 
        RECT 0.488 244.556 0.56 244.748 ; 
        RECT 28.928 244.556 29 244.748 ; 
        RECT 31.52 244.556 31.88 244.748 ; 
        RECT 37.136 244.556 37.208 244.748 ; 
        RECT 65.576 244.556 65.648 244.748 ; 
        RECT 0.488 248.876 0.56 249.068 ; 
        RECT 28.928 248.876 29 249.068 ; 
        RECT 31.52 248.876 31.88 249.068 ; 
        RECT 37.136 248.876 37.208 249.068 ; 
        RECT 65.576 248.876 65.648 249.068 ; 
        RECT 0.488 253.196 0.56 253.388 ; 
        RECT 28.928 253.196 29 253.388 ; 
        RECT 31.52 253.196 31.88 253.388 ; 
        RECT 37.136 253.196 37.208 253.388 ; 
        RECT 65.576 253.196 65.648 253.388 ; 
        RECT 0.488 257.516 0.56 257.708 ; 
        RECT 28.928 257.516 29 257.708 ; 
        RECT 31.52 257.516 31.88 257.708 ; 
        RECT 37.136 257.516 37.208 257.708 ; 
        RECT 65.576 257.516 65.648 257.708 ; 
        RECT 0.488 261.836 0.56 262.028 ; 
        RECT 28.928 261.836 29 262.028 ; 
        RECT 31.52 261.836 31.88 262.028 ; 
        RECT 37.136 261.836 37.208 262.028 ; 
        RECT 65.576 261.836 65.648 262.028 ; 
        RECT 0.488 266.156 0.56 266.348 ; 
        RECT 28.928 266.156 29 266.348 ; 
        RECT 31.52 266.156 31.88 266.348 ; 
        RECT 37.136 266.156 37.208 266.348 ; 
        RECT 65.576 266.156 65.648 266.348 ; 
        RECT 0.488 270.476 0.56 270.668 ; 
        RECT 28.928 270.476 29 270.668 ; 
        RECT 31.52 270.476 31.88 270.668 ; 
        RECT 37.136 270.476 37.208 270.668 ; 
        RECT 65.576 270.476 65.648 270.668 ; 
        RECT 0.488 274.796 0.56 274.988 ; 
        RECT 28.928 274.796 29 274.988 ; 
        RECT 31.52 274.796 31.88 274.988 ; 
        RECT 37.136 274.796 37.208 274.988 ; 
        RECT 65.576 274.796 65.648 274.988 ; 
        RECT 0.488 279.116 0.56 279.308 ; 
        RECT 28.928 279.116 29 279.308 ; 
        RECT 31.52 279.116 31.88 279.308 ; 
        RECT 37.136 279.116 37.208 279.308 ; 
        RECT 65.576 279.116 65.648 279.308 ; 
        RECT 0.488 283.436 0.56 283.628 ; 
        RECT 28.928 283.436 29 283.628 ; 
        RECT 31.52 283.436 31.88 283.628 ; 
        RECT 37.136 283.436 37.208 283.628 ; 
        RECT 65.576 283.436 65.648 283.628 ; 
        RECT 0.488 287.756 0.56 287.948 ; 
        RECT 28.928 287.756 29 287.948 ; 
        RECT 31.52 287.756 31.88 287.948 ; 
        RECT 37.136 287.756 37.208 287.948 ; 
        RECT 65.576 287.756 65.648 287.948 ; 
        RECT 0.488 292.076 0.56 292.268 ; 
        RECT 28.928 292.076 29 292.268 ; 
        RECT 31.52 292.076 31.88 292.268 ; 
        RECT 37.136 292.076 37.208 292.268 ; 
        RECT 65.576 292.076 65.648 292.268 ; 
        RECT 0.488 296.396 0.56 296.588 ; 
        RECT 28.928 296.396 29 296.588 ; 
        RECT 31.52 296.396 31.88 296.588 ; 
        RECT 37.136 296.396 37.208 296.588 ; 
        RECT 65.576 296.396 65.648 296.588 ; 
        RECT 0.488 300.716 0.56 300.908 ; 
        RECT 28.928 300.716 29 300.908 ; 
        RECT 31.52 300.716 31.88 300.908 ; 
        RECT 37.136 300.716 37.208 300.908 ; 
        RECT 65.576 300.716 65.648 300.908 ; 
        RECT 0.488 305.036 0.56 305.228 ; 
        RECT 28.928 305.036 29 305.228 ; 
        RECT 31.52 305.036 31.88 305.228 ; 
        RECT 37.136 305.036 37.208 305.228 ; 
        RECT 65.576 305.036 65.648 305.228 ; 
        RECT 0.488 309.356 0.56 309.548 ; 
        RECT 28.928 309.356 29 309.548 ; 
        RECT 31.52 309.356 31.88 309.548 ; 
        RECT 37.136 309.356 37.208 309.548 ; 
        RECT 65.576 309.356 65.648 309.548 ; 
        RECT 0.488 313.676 0.56 313.868 ; 
        RECT 28.928 313.676 29 313.868 ; 
        RECT 31.52 313.676 31.88 313.868 ; 
        RECT 37.136 313.676 37.208 313.868 ; 
        RECT 65.576 313.676 65.648 313.868 ; 
        RECT 0.488 317.996 0.56 318.188 ; 
        RECT 28.928 317.996 29 318.188 ; 
        RECT 31.52 317.996 31.88 318.188 ; 
        RECT 37.136 317.996 37.208 318.188 ; 
        RECT 65.576 317.996 65.648 318.188 ; 
        RECT 0.488 322.316 0.56 322.508 ; 
        RECT 28.928 322.316 29 322.508 ; 
        RECT 31.52 322.316 31.88 322.508 ; 
        RECT 37.136 322.316 37.208 322.508 ; 
        RECT 65.576 322.316 65.648 322.508 ; 
        RECT 0.488 326.636 0.56 326.828 ; 
        RECT 28.928 326.636 29 326.828 ; 
        RECT 31.52 326.636 31.88 326.828 ; 
        RECT 37.136 326.636 37.208 326.828 ; 
        RECT 65.576 326.636 65.648 326.828 ; 
        RECT 0.488 330.956 0.56 331.148 ; 
        RECT 28.928 330.956 29 331.148 ; 
        RECT 31.52 330.956 31.88 331.148 ; 
        RECT 37.136 330.956 37.208 331.148 ; 
        RECT 65.576 330.956 65.648 331.148 ; 
        RECT 0.488 335.276 0.56 335.468 ; 
        RECT 28.928 335.276 29 335.468 ; 
        RECT 31.52 335.276 31.88 335.468 ; 
        RECT 37.136 335.276 37.208 335.468 ; 
        RECT 65.576 335.276 65.648 335.468 ; 
        RECT 0.488 339.596 0.56 339.788 ; 
        RECT 28.928 339.596 29 339.788 ; 
        RECT 31.52 339.596 31.88 339.788 ; 
        RECT 37.136 339.596 37.208 339.788 ; 
        RECT 65.576 339.596 65.648 339.788 ; 
        RECT 0.488 343.916 0.56 344.108 ; 
        RECT 28.928 343.916 29 344.108 ; 
        RECT 31.52 343.916 31.88 344.108 ; 
        RECT 37.136 343.916 37.208 344.108 ; 
        RECT 65.576 343.916 65.648 344.108 ; 
        RECT 0.488 348.236 0.56 348.428 ; 
        RECT 28.928 348.236 29 348.428 ; 
        RECT 31.52 348.236 31.88 348.428 ; 
        RECT 37.136 348.236 37.208 348.428 ; 
        RECT 65.576 348.236 65.648 348.428 ; 
        RECT 0.488 352.556 0.56 352.748 ; 
        RECT 28.928 352.556 29 352.748 ; 
        RECT 31.52 352.556 31.88 352.748 ; 
        RECT 37.136 352.556 37.208 352.748 ; 
        RECT 65.576 352.556 65.648 352.748 ; 
      LAYER M5 ; 
        RECT 36.864 160.94 36.96 176.316 ; 
      LAYER V4 ; 
        RECT 36.864 176.148 36.96 176.244 ; 
        RECT 36.864 162.132 36.96 162.996 ; 
        RECT 36.864 161.012 36.96 161.108 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.304 65.748 4.496 ; 
        RECT 0.376 8.624 65.748 8.816 ; 
        RECT 0.376 12.944 65.748 13.136 ; 
        RECT 0.376 17.264 65.748 17.456 ; 
        RECT 0.376 21.584 65.748 21.776 ; 
        RECT 0.376 25.904 65.748 26.096 ; 
        RECT 0.376 30.224 65.748 30.416 ; 
        RECT 0.376 34.544 65.748 34.736 ; 
        RECT 0.376 38.864 65.748 39.056 ; 
        RECT 0.376 43.184 65.748 43.376 ; 
        RECT 0.376 47.504 65.748 47.696 ; 
        RECT 0.376 51.824 65.748 52.016 ; 
        RECT 0.376 56.144 65.748 56.336 ; 
        RECT 0.376 60.464 65.748 60.656 ; 
        RECT 0.376 64.784 65.748 64.976 ; 
        RECT 0.376 69.104 65.748 69.296 ; 
        RECT 0.376 73.424 65.748 73.616 ; 
        RECT 0.376 77.744 65.748 77.936 ; 
        RECT 0.376 82.064 65.748 82.256 ; 
        RECT 0.376 86.384 65.748 86.576 ; 
        RECT 0.376 90.704 65.748 90.896 ; 
        RECT 0.376 95.024 65.748 95.216 ; 
        RECT 0.376 99.344 65.748 99.536 ; 
        RECT 0.376 103.664 65.748 103.856 ; 
        RECT 0.376 107.984 65.748 108.176 ; 
        RECT 0.376 112.304 65.748 112.496 ; 
        RECT 0.376 116.624 65.748 116.816 ; 
        RECT 0.376 120.944 65.748 121.136 ; 
        RECT 0.376 125.264 65.748 125.456 ; 
        RECT 0.376 129.584 65.748 129.776 ; 
        RECT 0.376 133.904 65.748 134.096 ; 
        RECT 0.376 138.224 65.748 138.416 ; 
        RECT 0.376 142.544 65.748 142.736 ; 
        RECT 0.376 146.864 65.748 147.056 ; 
        RECT 0.376 151.184 65.748 151.376 ; 
        RECT 0.376 155.504 65.748 155.696 ; 
        RECT 0.376 159.824 65.748 160.016 ; 
        RECT 14.256 163.86 51.84 164.724 ; 
        RECT 29.592 176.532 36.504 177.396 ; 
        RECT 29.592 189.204 36.504 190.068 ; 
        RECT 0.376 196.652 65.748 196.844 ; 
        RECT 0.376 200.972 65.748 201.164 ; 
        RECT 0.376 205.292 65.748 205.484 ; 
        RECT 0.376 209.612 65.748 209.804 ; 
        RECT 0.376 213.932 65.748 214.124 ; 
        RECT 0.376 218.252 65.748 218.444 ; 
        RECT 0.376 222.572 65.748 222.764 ; 
        RECT 0.376 226.892 65.748 227.084 ; 
        RECT 0.376 231.212 65.748 231.404 ; 
        RECT 0.376 235.532 65.748 235.724 ; 
        RECT 0.376 239.852 65.748 240.044 ; 
        RECT 0.376 244.172 65.748 244.364 ; 
        RECT 0.376 248.492 65.748 248.684 ; 
        RECT 0.376 252.812 65.748 253.004 ; 
        RECT 0.376 257.132 65.748 257.324 ; 
        RECT 0.376 261.452 65.748 261.644 ; 
        RECT 0.376 265.772 65.748 265.964 ; 
        RECT 0.376 270.092 65.748 270.284 ; 
        RECT 0.376 274.412 65.748 274.604 ; 
        RECT 0.376 278.732 65.748 278.924 ; 
        RECT 0.376 283.052 65.748 283.244 ; 
        RECT 0.376 287.372 65.748 287.564 ; 
        RECT 0.376 291.692 65.748 291.884 ; 
        RECT 0.376 296.012 65.748 296.204 ; 
        RECT 0.376 300.332 65.748 300.524 ; 
        RECT 0.376 304.652 65.748 304.844 ; 
        RECT 0.376 308.972 65.748 309.164 ; 
        RECT 0.376 313.292 65.748 313.484 ; 
        RECT 0.376 317.612 65.748 317.804 ; 
        RECT 0.376 321.932 65.748 322.124 ; 
        RECT 0.376 326.252 65.748 326.444 ; 
        RECT 0.376 330.572 65.748 330.764 ; 
        RECT 0.376 334.892 65.748 335.084 ; 
        RECT 0.376 339.212 65.748 339.404 ; 
        RECT 0.376 343.532 65.748 343.724 ; 
        RECT 0.376 347.852 65.748 348.044 ; 
        RECT 0.376 352.172 65.748 352.364 ; 
      LAYER M3 ; 
        RECT 65.432 0.866 65.504 5.506 ; 
        RECT 37.352 0.866 37.424 5.506 ; 
        RECT 34.292 1.012 34.436 5.468 ; 
        RECT 33.68 1.012 33.788 5.468 ; 
        RECT 28.712 0.866 28.784 5.506 ; 
        RECT 0.632 0.866 0.704 5.506 ; 
        RECT 65.432 5.186 65.504 9.826 ; 
        RECT 37.352 5.186 37.424 9.826 ; 
        RECT 34.292 5.332 34.436 9.788 ; 
        RECT 33.68 5.332 33.788 9.788 ; 
        RECT 28.712 5.186 28.784 9.826 ; 
        RECT 0.632 5.186 0.704 9.826 ; 
        RECT 65.432 9.506 65.504 14.146 ; 
        RECT 37.352 9.506 37.424 14.146 ; 
        RECT 34.292 9.652 34.436 14.108 ; 
        RECT 33.68 9.652 33.788 14.108 ; 
        RECT 28.712 9.506 28.784 14.146 ; 
        RECT 0.632 9.506 0.704 14.146 ; 
        RECT 65.432 13.826 65.504 18.466 ; 
        RECT 37.352 13.826 37.424 18.466 ; 
        RECT 34.292 13.972 34.436 18.428 ; 
        RECT 33.68 13.972 33.788 18.428 ; 
        RECT 28.712 13.826 28.784 18.466 ; 
        RECT 0.632 13.826 0.704 18.466 ; 
        RECT 65.432 18.146 65.504 22.786 ; 
        RECT 37.352 18.146 37.424 22.786 ; 
        RECT 34.292 18.292 34.436 22.748 ; 
        RECT 33.68 18.292 33.788 22.748 ; 
        RECT 28.712 18.146 28.784 22.786 ; 
        RECT 0.632 18.146 0.704 22.786 ; 
        RECT 65.432 22.466 65.504 27.106 ; 
        RECT 37.352 22.466 37.424 27.106 ; 
        RECT 34.292 22.612 34.436 27.068 ; 
        RECT 33.68 22.612 33.788 27.068 ; 
        RECT 28.712 22.466 28.784 27.106 ; 
        RECT 0.632 22.466 0.704 27.106 ; 
        RECT 65.432 26.786 65.504 31.426 ; 
        RECT 37.352 26.786 37.424 31.426 ; 
        RECT 34.292 26.932 34.436 31.388 ; 
        RECT 33.68 26.932 33.788 31.388 ; 
        RECT 28.712 26.786 28.784 31.426 ; 
        RECT 0.632 26.786 0.704 31.426 ; 
        RECT 65.432 31.106 65.504 35.746 ; 
        RECT 37.352 31.106 37.424 35.746 ; 
        RECT 34.292 31.252 34.436 35.708 ; 
        RECT 33.68 31.252 33.788 35.708 ; 
        RECT 28.712 31.106 28.784 35.746 ; 
        RECT 0.632 31.106 0.704 35.746 ; 
        RECT 65.432 35.426 65.504 40.066 ; 
        RECT 37.352 35.426 37.424 40.066 ; 
        RECT 34.292 35.572 34.436 40.028 ; 
        RECT 33.68 35.572 33.788 40.028 ; 
        RECT 28.712 35.426 28.784 40.066 ; 
        RECT 0.632 35.426 0.704 40.066 ; 
        RECT 65.432 39.746 65.504 44.386 ; 
        RECT 37.352 39.746 37.424 44.386 ; 
        RECT 34.292 39.892 34.436 44.348 ; 
        RECT 33.68 39.892 33.788 44.348 ; 
        RECT 28.712 39.746 28.784 44.386 ; 
        RECT 0.632 39.746 0.704 44.386 ; 
        RECT 65.432 44.066 65.504 48.706 ; 
        RECT 37.352 44.066 37.424 48.706 ; 
        RECT 34.292 44.212 34.436 48.668 ; 
        RECT 33.68 44.212 33.788 48.668 ; 
        RECT 28.712 44.066 28.784 48.706 ; 
        RECT 0.632 44.066 0.704 48.706 ; 
        RECT 65.432 48.386 65.504 53.026 ; 
        RECT 37.352 48.386 37.424 53.026 ; 
        RECT 34.292 48.532 34.436 52.988 ; 
        RECT 33.68 48.532 33.788 52.988 ; 
        RECT 28.712 48.386 28.784 53.026 ; 
        RECT 0.632 48.386 0.704 53.026 ; 
        RECT 65.432 52.706 65.504 57.346 ; 
        RECT 37.352 52.706 37.424 57.346 ; 
        RECT 34.292 52.852 34.436 57.308 ; 
        RECT 33.68 52.852 33.788 57.308 ; 
        RECT 28.712 52.706 28.784 57.346 ; 
        RECT 0.632 52.706 0.704 57.346 ; 
        RECT 65.432 57.026 65.504 61.666 ; 
        RECT 37.352 57.026 37.424 61.666 ; 
        RECT 34.292 57.172 34.436 61.628 ; 
        RECT 33.68 57.172 33.788 61.628 ; 
        RECT 28.712 57.026 28.784 61.666 ; 
        RECT 0.632 57.026 0.704 61.666 ; 
        RECT 65.432 61.346 65.504 65.986 ; 
        RECT 37.352 61.346 37.424 65.986 ; 
        RECT 34.292 61.492 34.436 65.948 ; 
        RECT 33.68 61.492 33.788 65.948 ; 
        RECT 28.712 61.346 28.784 65.986 ; 
        RECT 0.632 61.346 0.704 65.986 ; 
        RECT 65.432 65.666 65.504 70.306 ; 
        RECT 37.352 65.666 37.424 70.306 ; 
        RECT 34.292 65.812 34.436 70.268 ; 
        RECT 33.68 65.812 33.788 70.268 ; 
        RECT 28.712 65.666 28.784 70.306 ; 
        RECT 0.632 65.666 0.704 70.306 ; 
        RECT 65.432 69.986 65.504 74.626 ; 
        RECT 37.352 69.986 37.424 74.626 ; 
        RECT 34.292 70.132 34.436 74.588 ; 
        RECT 33.68 70.132 33.788 74.588 ; 
        RECT 28.712 69.986 28.784 74.626 ; 
        RECT 0.632 69.986 0.704 74.626 ; 
        RECT 65.432 74.306 65.504 78.946 ; 
        RECT 37.352 74.306 37.424 78.946 ; 
        RECT 34.292 74.452 34.436 78.908 ; 
        RECT 33.68 74.452 33.788 78.908 ; 
        RECT 28.712 74.306 28.784 78.946 ; 
        RECT 0.632 74.306 0.704 78.946 ; 
        RECT 65.432 78.626 65.504 83.266 ; 
        RECT 37.352 78.626 37.424 83.266 ; 
        RECT 34.292 78.772 34.436 83.228 ; 
        RECT 33.68 78.772 33.788 83.228 ; 
        RECT 28.712 78.626 28.784 83.266 ; 
        RECT 0.632 78.626 0.704 83.266 ; 
        RECT 65.432 82.946 65.504 87.586 ; 
        RECT 37.352 82.946 37.424 87.586 ; 
        RECT 34.292 83.092 34.436 87.548 ; 
        RECT 33.68 83.092 33.788 87.548 ; 
        RECT 28.712 82.946 28.784 87.586 ; 
        RECT 0.632 82.946 0.704 87.586 ; 
        RECT 65.432 87.266 65.504 91.906 ; 
        RECT 37.352 87.266 37.424 91.906 ; 
        RECT 34.292 87.412 34.436 91.868 ; 
        RECT 33.68 87.412 33.788 91.868 ; 
        RECT 28.712 87.266 28.784 91.906 ; 
        RECT 0.632 87.266 0.704 91.906 ; 
        RECT 65.432 91.586 65.504 96.226 ; 
        RECT 37.352 91.586 37.424 96.226 ; 
        RECT 34.292 91.732 34.436 96.188 ; 
        RECT 33.68 91.732 33.788 96.188 ; 
        RECT 28.712 91.586 28.784 96.226 ; 
        RECT 0.632 91.586 0.704 96.226 ; 
        RECT 65.432 95.906 65.504 100.546 ; 
        RECT 37.352 95.906 37.424 100.546 ; 
        RECT 34.292 96.052 34.436 100.508 ; 
        RECT 33.68 96.052 33.788 100.508 ; 
        RECT 28.712 95.906 28.784 100.546 ; 
        RECT 0.632 95.906 0.704 100.546 ; 
        RECT 65.432 100.226 65.504 104.866 ; 
        RECT 37.352 100.226 37.424 104.866 ; 
        RECT 34.292 100.372 34.436 104.828 ; 
        RECT 33.68 100.372 33.788 104.828 ; 
        RECT 28.712 100.226 28.784 104.866 ; 
        RECT 0.632 100.226 0.704 104.866 ; 
        RECT 65.432 104.546 65.504 109.186 ; 
        RECT 37.352 104.546 37.424 109.186 ; 
        RECT 34.292 104.692 34.436 109.148 ; 
        RECT 33.68 104.692 33.788 109.148 ; 
        RECT 28.712 104.546 28.784 109.186 ; 
        RECT 0.632 104.546 0.704 109.186 ; 
        RECT 65.432 108.866 65.504 113.506 ; 
        RECT 37.352 108.866 37.424 113.506 ; 
        RECT 34.292 109.012 34.436 113.468 ; 
        RECT 33.68 109.012 33.788 113.468 ; 
        RECT 28.712 108.866 28.784 113.506 ; 
        RECT 0.632 108.866 0.704 113.506 ; 
        RECT 65.432 113.186 65.504 117.826 ; 
        RECT 37.352 113.186 37.424 117.826 ; 
        RECT 34.292 113.332 34.436 117.788 ; 
        RECT 33.68 113.332 33.788 117.788 ; 
        RECT 28.712 113.186 28.784 117.826 ; 
        RECT 0.632 113.186 0.704 117.826 ; 
        RECT 65.432 117.506 65.504 122.146 ; 
        RECT 37.352 117.506 37.424 122.146 ; 
        RECT 34.292 117.652 34.436 122.108 ; 
        RECT 33.68 117.652 33.788 122.108 ; 
        RECT 28.712 117.506 28.784 122.146 ; 
        RECT 0.632 117.506 0.704 122.146 ; 
        RECT 65.432 121.826 65.504 126.466 ; 
        RECT 37.352 121.826 37.424 126.466 ; 
        RECT 34.292 121.972 34.436 126.428 ; 
        RECT 33.68 121.972 33.788 126.428 ; 
        RECT 28.712 121.826 28.784 126.466 ; 
        RECT 0.632 121.826 0.704 126.466 ; 
        RECT 65.432 126.146 65.504 130.786 ; 
        RECT 37.352 126.146 37.424 130.786 ; 
        RECT 34.292 126.292 34.436 130.748 ; 
        RECT 33.68 126.292 33.788 130.748 ; 
        RECT 28.712 126.146 28.784 130.786 ; 
        RECT 0.632 126.146 0.704 130.786 ; 
        RECT 65.432 130.466 65.504 135.106 ; 
        RECT 37.352 130.466 37.424 135.106 ; 
        RECT 34.292 130.612 34.436 135.068 ; 
        RECT 33.68 130.612 33.788 135.068 ; 
        RECT 28.712 130.466 28.784 135.106 ; 
        RECT 0.632 130.466 0.704 135.106 ; 
        RECT 65.432 134.786 65.504 139.426 ; 
        RECT 37.352 134.786 37.424 139.426 ; 
        RECT 34.292 134.932 34.436 139.388 ; 
        RECT 33.68 134.932 33.788 139.388 ; 
        RECT 28.712 134.786 28.784 139.426 ; 
        RECT 0.632 134.786 0.704 139.426 ; 
        RECT 65.432 139.106 65.504 143.746 ; 
        RECT 37.352 139.106 37.424 143.746 ; 
        RECT 34.292 139.252 34.436 143.708 ; 
        RECT 33.68 139.252 33.788 143.708 ; 
        RECT 28.712 139.106 28.784 143.746 ; 
        RECT 0.632 139.106 0.704 143.746 ; 
        RECT 65.432 143.426 65.504 148.066 ; 
        RECT 37.352 143.426 37.424 148.066 ; 
        RECT 34.292 143.572 34.436 148.028 ; 
        RECT 33.68 143.572 33.788 148.028 ; 
        RECT 28.712 143.426 28.784 148.066 ; 
        RECT 0.632 143.426 0.704 148.066 ; 
        RECT 65.432 147.746 65.504 152.386 ; 
        RECT 37.352 147.746 37.424 152.386 ; 
        RECT 34.292 147.892 34.436 152.348 ; 
        RECT 33.68 147.892 33.788 152.348 ; 
        RECT 28.712 147.746 28.784 152.386 ; 
        RECT 0.632 147.746 0.704 152.386 ; 
        RECT 65.432 152.066 65.504 156.706 ; 
        RECT 37.352 152.066 37.424 156.706 ; 
        RECT 34.292 152.212 34.436 156.668 ; 
        RECT 33.68 152.212 33.788 156.668 ; 
        RECT 28.712 152.066 28.784 156.706 ; 
        RECT 0.632 152.066 0.704 156.706 ; 
        RECT 65.432 156.386 65.504 161.026 ; 
        RECT 37.352 156.386 37.424 161.026 ; 
        RECT 34.292 156.532 34.436 160.988 ; 
        RECT 33.68 156.532 33.788 160.988 ; 
        RECT 28.712 156.386 28.784 161.026 ; 
        RECT 0.632 156.386 0.704 161.026 ; 
        RECT 65.412 160.682 65.484 193.51 ; 
        RECT 37.332 160.682 37.404 193.51 ; 
        RECT 33.516 161.576 34.452 192.308 ; 
        RECT 34.272 160.858 34.416 193.336 ; 
        RECT 33.66 160.856 33.768 193.336 ; 
        RECT 28.692 160.682 28.764 193.51 ; 
        RECT 0.612 160.682 0.684 193.51 ; 
        RECT 65.432 193.214 65.504 197.854 ; 
        RECT 37.352 193.214 37.424 197.854 ; 
        RECT 34.292 193.36 34.436 197.816 ; 
        RECT 33.68 193.36 33.788 197.816 ; 
        RECT 28.712 193.214 28.784 197.854 ; 
        RECT 0.632 193.214 0.704 197.854 ; 
        RECT 65.432 197.534 65.504 202.174 ; 
        RECT 37.352 197.534 37.424 202.174 ; 
        RECT 34.292 197.68 34.436 202.136 ; 
        RECT 33.68 197.68 33.788 202.136 ; 
        RECT 28.712 197.534 28.784 202.174 ; 
        RECT 0.632 197.534 0.704 202.174 ; 
        RECT 65.432 201.854 65.504 206.494 ; 
        RECT 37.352 201.854 37.424 206.494 ; 
        RECT 34.292 202 34.436 206.456 ; 
        RECT 33.68 202 33.788 206.456 ; 
        RECT 28.712 201.854 28.784 206.494 ; 
        RECT 0.632 201.854 0.704 206.494 ; 
        RECT 65.432 206.174 65.504 210.814 ; 
        RECT 37.352 206.174 37.424 210.814 ; 
        RECT 34.292 206.32 34.436 210.776 ; 
        RECT 33.68 206.32 33.788 210.776 ; 
        RECT 28.712 206.174 28.784 210.814 ; 
        RECT 0.632 206.174 0.704 210.814 ; 
        RECT 65.432 210.494 65.504 215.134 ; 
        RECT 37.352 210.494 37.424 215.134 ; 
        RECT 34.292 210.64 34.436 215.096 ; 
        RECT 33.68 210.64 33.788 215.096 ; 
        RECT 28.712 210.494 28.784 215.134 ; 
        RECT 0.632 210.494 0.704 215.134 ; 
        RECT 65.432 214.814 65.504 219.454 ; 
        RECT 37.352 214.814 37.424 219.454 ; 
        RECT 34.292 214.96 34.436 219.416 ; 
        RECT 33.68 214.96 33.788 219.416 ; 
        RECT 28.712 214.814 28.784 219.454 ; 
        RECT 0.632 214.814 0.704 219.454 ; 
        RECT 65.432 219.134 65.504 223.774 ; 
        RECT 37.352 219.134 37.424 223.774 ; 
        RECT 34.292 219.28 34.436 223.736 ; 
        RECT 33.68 219.28 33.788 223.736 ; 
        RECT 28.712 219.134 28.784 223.774 ; 
        RECT 0.632 219.134 0.704 223.774 ; 
        RECT 65.432 223.454 65.504 228.094 ; 
        RECT 37.352 223.454 37.424 228.094 ; 
        RECT 34.292 223.6 34.436 228.056 ; 
        RECT 33.68 223.6 33.788 228.056 ; 
        RECT 28.712 223.454 28.784 228.094 ; 
        RECT 0.632 223.454 0.704 228.094 ; 
        RECT 65.432 227.774 65.504 232.414 ; 
        RECT 37.352 227.774 37.424 232.414 ; 
        RECT 34.292 227.92 34.436 232.376 ; 
        RECT 33.68 227.92 33.788 232.376 ; 
        RECT 28.712 227.774 28.784 232.414 ; 
        RECT 0.632 227.774 0.704 232.414 ; 
        RECT 65.432 232.094 65.504 236.734 ; 
        RECT 37.352 232.094 37.424 236.734 ; 
        RECT 34.292 232.24 34.436 236.696 ; 
        RECT 33.68 232.24 33.788 236.696 ; 
        RECT 28.712 232.094 28.784 236.734 ; 
        RECT 0.632 232.094 0.704 236.734 ; 
        RECT 65.432 236.414 65.504 241.054 ; 
        RECT 37.352 236.414 37.424 241.054 ; 
        RECT 34.292 236.56 34.436 241.016 ; 
        RECT 33.68 236.56 33.788 241.016 ; 
        RECT 28.712 236.414 28.784 241.054 ; 
        RECT 0.632 236.414 0.704 241.054 ; 
        RECT 65.432 240.734 65.504 245.374 ; 
        RECT 37.352 240.734 37.424 245.374 ; 
        RECT 34.292 240.88 34.436 245.336 ; 
        RECT 33.68 240.88 33.788 245.336 ; 
        RECT 28.712 240.734 28.784 245.374 ; 
        RECT 0.632 240.734 0.704 245.374 ; 
        RECT 65.432 245.054 65.504 249.694 ; 
        RECT 37.352 245.054 37.424 249.694 ; 
        RECT 34.292 245.2 34.436 249.656 ; 
        RECT 33.68 245.2 33.788 249.656 ; 
        RECT 28.712 245.054 28.784 249.694 ; 
        RECT 0.632 245.054 0.704 249.694 ; 
        RECT 65.432 249.374 65.504 254.014 ; 
        RECT 37.352 249.374 37.424 254.014 ; 
        RECT 34.292 249.52 34.436 253.976 ; 
        RECT 33.68 249.52 33.788 253.976 ; 
        RECT 28.712 249.374 28.784 254.014 ; 
        RECT 0.632 249.374 0.704 254.014 ; 
        RECT 65.432 253.694 65.504 258.334 ; 
        RECT 37.352 253.694 37.424 258.334 ; 
        RECT 34.292 253.84 34.436 258.296 ; 
        RECT 33.68 253.84 33.788 258.296 ; 
        RECT 28.712 253.694 28.784 258.334 ; 
        RECT 0.632 253.694 0.704 258.334 ; 
        RECT 65.432 258.014 65.504 262.654 ; 
        RECT 37.352 258.014 37.424 262.654 ; 
        RECT 34.292 258.16 34.436 262.616 ; 
        RECT 33.68 258.16 33.788 262.616 ; 
        RECT 28.712 258.014 28.784 262.654 ; 
        RECT 0.632 258.014 0.704 262.654 ; 
        RECT 65.432 262.334 65.504 266.974 ; 
        RECT 37.352 262.334 37.424 266.974 ; 
        RECT 34.292 262.48 34.436 266.936 ; 
        RECT 33.68 262.48 33.788 266.936 ; 
        RECT 28.712 262.334 28.784 266.974 ; 
        RECT 0.632 262.334 0.704 266.974 ; 
        RECT 65.432 266.654 65.504 271.294 ; 
        RECT 37.352 266.654 37.424 271.294 ; 
        RECT 34.292 266.8 34.436 271.256 ; 
        RECT 33.68 266.8 33.788 271.256 ; 
        RECT 28.712 266.654 28.784 271.294 ; 
        RECT 0.632 266.654 0.704 271.294 ; 
        RECT 65.432 270.974 65.504 275.614 ; 
        RECT 37.352 270.974 37.424 275.614 ; 
        RECT 34.292 271.12 34.436 275.576 ; 
        RECT 33.68 271.12 33.788 275.576 ; 
        RECT 28.712 270.974 28.784 275.614 ; 
        RECT 0.632 270.974 0.704 275.614 ; 
        RECT 65.432 275.294 65.504 279.934 ; 
        RECT 37.352 275.294 37.424 279.934 ; 
        RECT 34.292 275.44 34.436 279.896 ; 
        RECT 33.68 275.44 33.788 279.896 ; 
        RECT 28.712 275.294 28.784 279.934 ; 
        RECT 0.632 275.294 0.704 279.934 ; 
        RECT 65.432 279.614 65.504 284.254 ; 
        RECT 37.352 279.614 37.424 284.254 ; 
        RECT 34.292 279.76 34.436 284.216 ; 
        RECT 33.68 279.76 33.788 284.216 ; 
        RECT 28.712 279.614 28.784 284.254 ; 
        RECT 0.632 279.614 0.704 284.254 ; 
        RECT 65.432 283.934 65.504 288.574 ; 
        RECT 37.352 283.934 37.424 288.574 ; 
        RECT 34.292 284.08 34.436 288.536 ; 
        RECT 33.68 284.08 33.788 288.536 ; 
        RECT 28.712 283.934 28.784 288.574 ; 
        RECT 0.632 283.934 0.704 288.574 ; 
        RECT 65.432 288.254 65.504 292.894 ; 
        RECT 37.352 288.254 37.424 292.894 ; 
        RECT 34.292 288.4 34.436 292.856 ; 
        RECT 33.68 288.4 33.788 292.856 ; 
        RECT 28.712 288.254 28.784 292.894 ; 
        RECT 0.632 288.254 0.704 292.894 ; 
        RECT 65.432 292.574 65.504 297.214 ; 
        RECT 37.352 292.574 37.424 297.214 ; 
        RECT 34.292 292.72 34.436 297.176 ; 
        RECT 33.68 292.72 33.788 297.176 ; 
        RECT 28.712 292.574 28.784 297.214 ; 
        RECT 0.632 292.574 0.704 297.214 ; 
        RECT 65.432 296.894 65.504 301.534 ; 
        RECT 37.352 296.894 37.424 301.534 ; 
        RECT 34.292 297.04 34.436 301.496 ; 
        RECT 33.68 297.04 33.788 301.496 ; 
        RECT 28.712 296.894 28.784 301.534 ; 
        RECT 0.632 296.894 0.704 301.534 ; 
        RECT 65.432 301.214 65.504 305.854 ; 
        RECT 37.352 301.214 37.424 305.854 ; 
        RECT 34.292 301.36 34.436 305.816 ; 
        RECT 33.68 301.36 33.788 305.816 ; 
        RECT 28.712 301.214 28.784 305.854 ; 
        RECT 0.632 301.214 0.704 305.854 ; 
        RECT 65.432 305.534 65.504 310.174 ; 
        RECT 37.352 305.534 37.424 310.174 ; 
        RECT 34.292 305.68 34.436 310.136 ; 
        RECT 33.68 305.68 33.788 310.136 ; 
        RECT 28.712 305.534 28.784 310.174 ; 
        RECT 0.632 305.534 0.704 310.174 ; 
        RECT 65.432 309.854 65.504 314.494 ; 
        RECT 37.352 309.854 37.424 314.494 ; 
        RECT 34.292 310 34.436 314.456 ; 
        RECT 33.68 310 33.788 314.456 ; 
        RECT 28.712 309.854 28.784 314.494 ; 
        RECT 0.632 309.854 0.704 314.494 ; 
        RECT 65.432 314.174 65.504 318.814 ; 
        RECT 37.352 314.174 37.424 318.814 ; 
        RECT 34.292 314.32 34.436 318.776 ; 
        RECT 33.68 314.32 33.788 318.776 ; 
        RECT 28.712 314.174 28.784 318.814 ; 
        RECT 0.632 314.174 0.704 318.814 ; 
        RECT 65.432 318.494 65.504 323.134 ; 
        RECT 37.352 318.494 37.424 323.134 ; 
        RECT 34.292 318.64 34.436 323.096 ; 
        RECT 33.68 318.64 33.788 323.096 ; 
        RECT 28.712 318.494 28.784 323.134 ; 
        RECT 0.632 318.494 0.704 323.134 ; 
        RECT 65.432 322.814 65.504 327.454 ; 
        RECT 37.352 322.814 37.424 327.454 ; 
        RECT 34.292 322.96 34.436 327.416 ; 
        RECT 33.68 322.96 33.788 327.416 ; 
        RECT 28.712 322.814 28.784 327.454 ; 
        RECT 0.632 322.814 0.704 327.454 ; 
        RECT 65.432 327.134 65.504 331.774 ; 
        RECT 37.352 327.134 37.424 331.774 ; 
        RECT 34.292 327.28 34.436 331.736 ; 
        RECT 33.68 327.28 33.788 331.736 ; 
        RECT 28.712 327.134 28.784 331.774 ; 
        RECT 0.632 327.134 0.704 331.774 ; 
        RECT 65.432 331.454 65.504 336.094 ; 
        RECT 37.352 331.454 37.424 336.094 ; 
        RECT 34.292 331.6 34.436 336.056 ; 
        RECT 33.68 331.6 33.788 336.056 ; 
        RECT 28.712 331.454 28.784 336.094 ; 
        RECT 0.632 331.454 0.704 336.094 ; 
        RECT 65.432 335.774 65.504 340.414 ; 
        RECT 37.352 335.774 37.424 340.414 ; 
        RECT 34.292 335.92 34.436 340.376 ; 
        RECT 33.68 335.92 33.788 340.376 ; 
        RECT 28.712 335.774 28.784 340.414 ; 
        RECT 0.632 335.774 0.704 340.414 ; 
        RECT 65.432 340.094 65.504 344.734 ; 
        RECT 37.352 340.094 37.424 344.734 ; 
        RECT 34.292 340.24 34.436 344.696 ; 
        RECT 33.68 340.24 33.788 344.696 ; 
        RECT 28.712 340.094 28.784 344.734 ; 
        RECT 0.632 340.094 0.704 344.734 ; 
        RECT 65.432 344.414 65.504 349.054 ; 
        RECT 37.352 344.414 37.424 349.054 ; 
        RECT 34.292 344.56 34.436 349.016 ; 
        RECT 33.68 344.56 33.788 349.016 ; 
        RECT 28.712 344.414 28.784 349.054 ; 
        RECT 0.632 344.414 0.704 349.054 ; 
        RECT 65.432 348.734 65.504 353.374 ; 
        RECT 37.352 348.734 37.424 353.374 ; 
        RECT 34.292 348.88 34.436 353.336 ; 
        RECT 33.68 348.88 33.788 353.336 ; 
        RECT 28.712 348.734 28.784 353.374 ; 
        RECT 0.632 348.734 0.704 353.374 ; 
      LAYER V3 ; 
        RECT 0.632 4.304 0.704 4.496 ; 
        RECT 28.712 4.304 28.784 4.496 ; 
        RECT 33.68 4.304 33.788 4.496 ; 
        RECT 34.292 4.304 34.436 4.496 ; 
        RECT 37.352 4.304 37.424 4.496 ; 
        RECT 65.432 4.304 65.504 4.496 ; 
        RECT 0.632 8.624 0.704 8.816 ; 
        RECT 28.712 8.624 28.784 8.816 ; 
        RECT 33.68 8.624 33.788 8.816 ; 
        RECT 34.292 8.624 34.436 8.816 ; 
        RECT 37.352 8.624 37.424 8.816 ; 
        RECT 65.432 8.624 65.504 8.816 ; 
        RECT 0.632 12.944 0.704 13.136 ; 
        RECT 28.712 12.944 28.784 13.136 ; 
        RECT 33.68 12.944 33.788 13.136 ; 
        RECT 34.292 12.944 34.436 13.136 ; 
        RECT 37.352 12.944 37.424 13.136 ; 
        RECT 65.432 12.944 65.504 13.136 ; 
        RECT 0.632 17.264 0.704 17.456 ; 
        RECT 28.712 17.264 28.784 17.456 ; 
        RECT 33.68 17.264 33.788 17.456 ; 
        RECT 34.292 17.264 34.436 17.456 ; 
        RECT 37.352 17.264 37.424 17.456 ; 
        RECT 65.432 17.264 65.504 17.456 ; 
        RECT 0.632 21.584 0.704 21.776 ; 
        RECT 28.712 21.584 28.784 21.776 ; 
        RECT 33.68 21.584 33.788 21.776 ; 
        RECT 34.292 21.584 34.436 21.776 ; 
        RECT 37.352 21.584 37.424 21.776 ; 
        RECT 65.432 21.584 65.504 21.776 ; 
        RECT 0.632 25.904 0.704 26.096 ; 
        RECT 28.712 25.904 28.784 26.096 ; 
        RECT 33.68 25.904 33.788 26.096 ; 
        RECT 34.292 25.904 34.436 26.096 ; 
        RECT 37.352 25.904 37.424 26.096 ; 
        RECT 65.432 25.904 65.504 26.096 ; 
        RECT 0.632 30.224 0.704 30.416 ; 
        RECT 28.712 30.224 28.784 30.416 ; 
        RECT 33.68 30.224 33.788 30.416 ; 
        RECT 34.292 30.224 34.436 30.416 ; 
        RECT 37.352 30.224 37.424 30.416 ; 
        RECT 65.432 30.224 65.504 30.416 ; 
        RECT 0.632 34.544 0.704 34.736 ; 
        RECT 28.712 34.544 28.784 34.736 ; 
        RECT 33.68 34.544 33.788 34.736 ; 
        RECT 34.292 34.544 34.436 34.736 ; 
        RECT 37.352 34.544 37.424 34.736 ; 
        RECT 65.432 34.544 65.504 34.736 ; 
        RECT 0.632 38.864 0.704 39.056 ; 
        RECT 28.712 38.864 28.784 39.056 ; 
        RECT 33.68 38.864 33.788 39.056 ; 
        RECT 34.292 38.864 34.436 39.056 ; 
        RECT 37.352 38.864 37.424 39.056 ; 
        RECT 65.432 38.864 65.504 39.056 ; 
        RECT 0.632 43.184 0.704 43.376 ; 
        RECT 28.712 43.184 28.784 43.376 ; 
        RECT 33.68 43.184 33.788 43.376 ; 
        RECT 34.292 43.184 34.436 43.376 ; 
        RECT 37.352 43.184 37.424 43.376 ; 
        RECT 65.432 43.184 65.504 43.376 ; 
        RECT 0.632 47.504 0.704 47.696 ; 
        RECT 28.712 47.504 28.784 47.696 ; 
        RECT 33.68 47.504 33.788 47.696 ; 
        RECT 34.292 47.504 34.436 47.696 ; 
        RECT 37.352 47.504 37.424 47.696 ; 
        RECT 65.432 47.504 65.504 47.696 ; 
        RECT 0.632 51.824 0.704 52.016 ; 
        RECT 28.712 51.824 28.784 52.016 ; 
        RECT 33.68 51.824 33.788 52.016 ; 
        RECT 34.292 51.824 34.436 52.016 ; 
        RECT 37.352 51.824 37.424 52.016 ; 
        RECT 65.432 51.824 65.504 52.016 ; 
        RECT 0.632 56.144 0.704 56.336 ; 
        RECT 28.712 56.144 28.784 56.336 ; 
        RECT 33.68 56.144 33.788 56.336 ; 
        RECT 34.292 56.144 34.436 56.336 ; 
        RECT 37.352 56.144 37.424 56.336 ; 
        RECT 65.432 56.144 65.504 56.336 ; 
        RECT 0.632 60.464 0.704 60.656 ; 
        RECT 28.712 60.464 28.784 60.656 ; 
        RECT 33.68 60.464 33.788 60.656 ; 
        RECT 34.292 60.464 34.436 60.656 ; 
        RECT 37.352 60.464 37.424 60.656 ; 
        RECT 65.432 60.464 65.504 60.656 ; 
        RECT 0.632 64.784 0.704 64.976 ; 
        RECT 28.712 64.784 28.784 64.976 ; 
        RECT 33.68 64.784 33.788 64.976 ; 
        RECT 34.292 64.784 34.436 64.976 ; 
        RECT 37.352 64.784 37.424 64.976 ; 
        RECT 65.432 64.784 65.504 64.976 ; 
        RECT 0.632 69.104 0.704 69.296 ; 
        RECT 28.712 69.104 28.784 69.296 ; 
        RECT 33.68 69.104 33.788 69.296 ; 
        RECT 34.292 69.104 34.436 69.296 ; 
        RECT 37.352 69.104 37.424 69.296 ; 
        RECT 65.432 69.104 65.504 69.296 ; 
        RECT 0.632 73.424 0.704 73.616 ; 
        RECT 28.712 73.424 28.784 73.616 ; 
        RECT 33.68 73.424 33.788 73.616 ; 
        RECT 34.292 73.424 34.436 73.616 ; 
        RECT 37.352 73.424 37.424 73.616 ; 
        RECT 65.432 73.424 65.504 73.616 ; 
        RECT 0.632 77.744 0.704 77.936 ; 
        RECT 28.712 77.744 28.784 77.936 ; 
        RECT 33.68 77.744 33.788 77.936 ; 
        RECT 34.292 77.744 34.436 77.936 ; 
        RECT 37.352 77.744 37.424 77.936 ; 
        RECT 65.432 77.744 65.504 77.936 ; 
        RECT 0.632 82.064 0.704 82.256 ; 
        RECT 28.712 82.064 28.784 82.256 ; 
        RECT 33.68 82.064 33.788 82.256 ; 
        RECT 34.292 82.064 34.436 82.256 ; 
        RECT 37.352 82.064 37.424 82.256 ; 
        RECT 65.432 82.064 65.504 82.256 ; 
        RECT 0.632 86.384 0.704 86.576 ; 
        RECT 28.712 86.384 28.784 86.576 ; 
        RECT 33.68 86.384 33.788 86.576 ; 
        RECT 34.292 86.384 34.436 86.576 ; 
        RECT 37.352 86.384 37.424 86.576 ; 
        RECT 65.432 86.384 65.504 86.576 ; 
        RECT 0.632 90.704 0.704 90.896 ; 
        RECT 28.712 90.704 28.784 90.896 ; 
        RECT 33.68 90.704 33.788 90.896 ; 
        RECT 34.292 90.704 34.436 90.896 ; 
        RECT 37.352 90.704 37.424 90.896 ; 
        RECT 65.432 90.704 65.504 90.896 ; 
        RECT 0.632 95.024 0.704 95.216 ; 
        RECT 28.712 95.024 28.784 95.216 ; 
        RECT 33.68 95.024 33.788 95.216 ; 
        RECT 34.292 95.024 34.436 95.216 ; 
        RECT 37.352 95.024 37.424 95.216 ; 
        RECT 65.432 95.024 65.504 95.216 ; 
        RECT 0.632 99.344 0.704 99.536 ; 
        RECT 28.712 99.344 28.784 99.536 ; 
        RECT 33.68 99.344 33.788 99.536 ; 
        RECT 34.292 99.344 34.436 99.536 ; 
        RECT 37.352 99.344 37.424 99.536 ; 
        RECT 65.432 99.344 65.504 99.536 ; 
        RECT 0.632 103.664 0.704 103.856 ; 
        RECT 28.712 103.664 28.784 103.856 ; 
        RECT 33.68 103.664 33.788 103.856 ; 
        RECT 34.292 103.664 34.436 103.856 ; 
        RECT 37.352 103.664 37.424 103.856 ; 
        RECT 65.432 103.664 65.504 103.856 ; 
        RECT 0.632 107.984 0.704 108.176 ; 
        RECT 28.712 107.984 28.784 108.176 ; 
        RECT 33.68 107.984 33.788 108.176 ; 
        RECT 34.292 107.984 34.436 108.176 ; 
        RECT 37.352 107.984 37.424 108.176 ; 
        RECT 65.432 107.984 65.504 108.176 ; 
        RECT 0.632 112.304 0.704 112.496 ; 
        RECT 28.712 112.304 28.784 112.496 ; 
        RECT 33.68 112.304 33.788 112.496 ; 
        RECT 34.292 112.304 34.436 112.496 ; 
        RECT 37.352 112.304 37.424 112.496 ; 
        RECT 65.432 112.304 65.504 112.496 ; 
        RECT 0.632 116.624 0.704 116.816 ; 
        RECT 28.712 116.624 28.784 116.816 ; 
        RECT 33.68 116.624 33.788 116.816 ; 
        RECT 34.292 116.624 34.436 116.816 ; 
        RECT 37.352 116.624 37.424 116.816 ; 
        RECT 65.432 116.624 65.504 116.816 ; 
        RECT 0.632 120.944 0.704 121.136 ; 
        RECT 28.712 120.944 28.784 121.136 ; 
        RECT 33.68 120.944 33.788 121.136 ; 
        RECT 34.292 120.944 34.436 121.136 ; 
        RECT 37.352 120.944 37.424 121.136 ; 
        RECT 65.432 120.944 65.504 121.136 ; 
        RECT 0.632 125.264 0.704 125.456 ; 
        RECT 28.712 125.264 28.784 125.456 ; 
        RECT 33.68 125.264 33.788 125.456 ; 
        RECT 34.292 125.264 34.436 125.456 ; 
        RECT 37.352 125.264 37.424 125.456 ; 
        RECT 65.432 125.264 65.504 125.456 ; 
        RECT 0.632 129.584 0.704 129.776 ; 
        RECT 28.712 129.584 28.784 129.776 ; 
        RECT 33.68 129.584 33.788 129.776 ; 
        RECT 34.292 129.584 34.436 129.776 ; 
        RECT 37.352 129.584 37.424 129.776 ; 
        RECT 65.432 129.584 65.504 129.776 ; 
        RECT 0.632 133.904 0.704 134.096 ; 
        RECT 28.712 133.904 28.784 134.096 ; 
        RECT 33.68 133.904 33.788 134.096 ; 
        RECT 34.292 133.904 34.436 134.096 ; 
        RECT 37.352 133.904 37.424 134.096 ; 
        RECT 65.432 133.904 65.504 134.096 ; 
        RECT 0.632 138.224 0.704 138.416 ; 
        RECT 28.712 138.224 28.784 138.416 ; 
        RECT 33.68 138.224 33.788 138.416 ; 
        RECT 34.292 138.224 34.436 138.416 ; 
        RECT 37.352 138.224 37.424 138.416 ; 
        RECT 65.432 138.224 65.504 138.416 ; 
        RECT 0.632 142.544 0.704 142.736 ; 
        RECT 28.712 142.544 28.784 142.736 ; 
        RECT 33.68 142.544 33.788 142.736 ; 
        RECT 34.292 142.544 34.436 142.736 ; 
        RECT 37.352 142.544 37.424 142.736 ; 
        RECT 65.432 142.544 65.504 142.736 ; 
        RECT 0.632 146.864 0.704 147.056 ; 
        RECT 28.712 146.864 28.784 147.056 ; 
        RECT 33.68 146.864 33.788 147.056 ; 
        RECT 34.292 146.864 34.436 147.056 ; 
        RECT 37.352 146.864 37.424 147.056 ; 
        RECT 65.432 146.864 65.504 147.056 ; 
        RECT 0.632 151.184 0.704 151.376 ; 
        RECT 28.712 151.184 28.784 151.376 ; 
        RECT 33.68 151.184 33.788 151.376 ; 
        RECT 34.292 151.184 34.436 151.376 ; 
        RECT 37.352 151.184 37.424 151.376 ; 
        RECT 65.432 151.184 65.504 151.376 ; 
        RECT 0.632 155.504 0.704 155.696 ; 
        RECT 28.712 155.504 28.784 155.696 ; 
        RECT 33.68 155.504 33.788 155.696 ; 
        RECT 34.292 155.504 34.436 155.696 ; 
        RECT 37.352 155.504 37.424 155.696 ; 
        RECT 65.432 155.504 65.504 155.696 ; 
        RECT 0.632 159.824 0.704 160.016 ; 
        RECT 28.712 159.824 28.784 160.016 ; 
        RECT 33.68 159.824 33.788 160.016 ; 
        RECT 34.292 159.824 34.436 160.016 ; 
        RECT 37.352 159.824 37.424 160.016 ; 
        RECT 65.432 159.824 65.504 160.016 ; 
        RECT 33.532 189.204 33.604 190.068 ; 
        RECT 33.532 176.532 33.604 177.396 ; 
        RECT 33.532 163.86 33.604 164.724 ; 
        RECT 33.74 189.204 33.812 190.068 ; 
        RECT 33.74 176.532 33.812 177.396 ; 
        RECT 33.74 163.86 33.812 164.724 ; 
        RECT 33.948 189.204 34.02 190.068 ; 
        RECT 33.948 176.532 34.02 177.396 ; 
        RECT 33.948 163.86 34.02 164.724 ; 
        RECT 34.156 189.204 34.228 190.068 ; 
        RECT 34.156 176.532 34.228 177.396 ; 
        RECT 34.156 163.86 34.228 164.724 ; 
        RECT 34.364 189.204 34.436 190.068 ; 
        RECT 34.364 176.532 34.436 177.396 ; 
        RECT 34.364 163.86 34.436 164.724 ; 
        RECT 37.332 163.862 37.404 164.726 ; 
        RECT 0.632 196.652 0.704 196.844 ; 
        RECT 28.712 196.652 28.784 196.844 ; 
        RECT 33.68 196.652 33.788 196.844 ; 
        RECT 34.292 196.652 34.436 196.844 ; 
        RECT 37.352 196.652 37.424 196.844 ; 
        RECT 65.432 196.652 65.504 196.844 ; 
        RECT 0.632 200.972 0.704 201.164 ; 
        RECT 28.712 200.972 28.784 201.164 ; 
        RECT 33.68 200.972 33.788 201.164 ; 
        RECT 34.292 200.972 34.436 201.164 ; 
        RECT 37.352 200.972 37.424 201.164 ; 
        RECT 65.432 200.972 65.504 201.164 ; 
        RECT 0.632 205.292 0.704 205.484 ; 
        RECT 28.712 205.292 28.784 205.484 ; 
        RECT 33.68 205.292 33.788 205.484 ; 
        RECT 34.292 205.292 34.436 205.484 ; 
        RECT 37.352 205.292 37.424 205.484 ; 
        RECT 65.432 205.292 65.504 205.484 ; 
        RECT 0.632 209.612 0.704 209.804 ; 
        RECT 28.712 209.612 28.784 209.804 ; 
        RECT 33.68 209.612 33.788 209.804 ; 
        RECT 34.292 209.612 34.436 209.804 ; 
        RECT 37.352 209.612 37.424 209.804 ; 
        RECT 65.432 209.612 65.504 209.804 ; 
        RECT 0.632 213.932 0.704 214.124 ; 
        RECT 28.712 213.932 28.784 214.124 ; 
        RECT 33.68 213.932 33.788 214.124 ; 
        RECT 34.292 213.932 34.436 214.124 ; 
        RECT 37.352 213.932 37.424 214.124 ; 
        RECT 65.432 213.932 65.504 214.124 ; 
        RECT 0.632 218.252 0.704 218.444 ; 
        RECT 28.712 218.252 28.784 218.444 ; 
        RECT 33.68 218.252 33.788 218.444 ; 
        RECT 34.292 218.252 34.436 218.444 ; 
        RECT 37.352 218.252 37.424 218.444 ; 
        RECT 65.432 218.252 65.504 218.444 ; 
        RECT 0.632 222.572 0.704 222.764 ; 
        RECT 28.712 222.572 28.784 222.764 ; 
        RECT 33.68 222.572 33.788 222.764 ; 
        RECT 34.292 222.572 34.436 222.764 ; 
        RECT 37.352 222.572 37.424 222.764 ; 
        RECT 65.432 222.572 65.504 222.764 ; 
        RECT 0.632 226.892 0.704 227.084 ; 
        RECT 28.712 226.892 28.784 227.084 ; 
        RECT 33.68 226.892 33.788 227.084 ; 
        RECT 34.292 226.892 34.436 227.084 ; 
        RECT 37.352 226.892 37.424 227.084 ; 
        RECT 65.432 226.892 65.504 227.084 ; 
        RECT 0.632 231.212 0.704 231.404 ; 
        RECT 28.712 231.212 28.784 231.404 ; 
        RECT 33.68 231.212 33.788 231.404 ; 
        RECT 34.292 231.212 34.436 231.404 ; 
        RECT 37.352 231.212 37.424 231.404 ; 
        RECT 65.432 231.212 65.504 231.404 ; 
        RECT 0.632 235.532 0.704 235.724 ; 
        RECT 28.712 235.532 28.784 235.724 ; 
        RECT 33.68 235.532 33.788 235.724 ; 
        RECT 34.292 235.532 34.436 235.724 ; 
        RECT 37.352 235.532 37.424 235.724 ; 
        RECT 65.432 235.532 65.504 235.724 ; 
        RECT 0.632 239.852 0.704 240.044 ; 
        RECT 28.712 239.852 28.784 240.044 ; 
        RECT 33.68 239.852 33.788 240.044 ; 
        RECT 34.292 239.852 34.436 240.044 ; 
        RECT 37.352 239.852 37.424 240.044 ; 
        RECT 65.432 239.852 65.504 240.044 ; 
        RECT 0.632 244.172 0.704 244.364 ; 
        RECT 28.712 244.172 28.784 244.364 ; 
        RECT 33.68 244.172 33.788 244.364 ; 
        RECT 34.292 244.172 34.436 244.364 ; 
        RECT 37.352 244.172 37.424 244.364 ; 
        RECT 65.432 244.172 65.504 244.364 ; 
        RECT 0.632 248.492 0.704 248.684 ; 
        RECT 28.712 248.492 28.784 248.684 ; 
        RECT 33.68 248.492 33.788 248.684 ; 
        RECT 34.292 248.492 34.436 248.684 ; 
        RECT 37.352 248.492 37.424 248.684 ; 
        RECT 65.432 248.492 65.504 248.684 ; 
        RECT 0.632 252.812 0.704 253.004 ; 
        RECT 28.712 252.812 28.784 253.004 ; 
        RECT 33.68 252.812 33.788 253.004 ; 
        RECT 34.292 252.812 34.436 253.004 ; 
        RECT 37.352 252.812 37.424 253.004 ; 
        RECT 65.432 252.812 65.504 253.004 ; 
        RECT 0.632 257.132 0.704 257.324 ; 
        RECT 28.712 257.132 28.784 257.324 ; 
        RECT 33.68 257.132 33.788 257.324 ; 
        RECT 34.292 257.132 34.436 257.324 ; 
        RECT 37.352 257.132 37.424 257.324 ; 
        RECT 65.432 257.132 65.504 257.324 ; 
        RECT 0.632 261.452 0.704 261.644 ; 
        RECT 28.712 261.452 28.784 261.644 ; 
        RECT 33.68 261.452 33.788 261.644 ; 
        RECT 34.292 261.452 34.436 261.644 ; 
        RECT 37.352 261.452 37.424 261.644 ; 
        RECT 65.432 261.452 65.504 261.644 ; 
        RECT 0.632 265.772 0.704 265.964 ; 
        RECT 28.712 265.772 28.784 265.964 ; 
        RECT 33.68 265.772 33.788 265.964 ; 
        RECT 34.292 265.772 34.436 265.964 ; 
        RECT 37.352 265.772 37.424 265.964 ; 
        RECT 65.432 265.772 65.504 265.964 ; 
        RECT 0.632 270.092 0.704 270.284 ; 
        RECT 28.712 270.092 28.784 270.284 ; 
        RECT 33.68 270.092 33.788 270.284 ; 
        RECT 34.292 270.092 34.436 270.284 ; 
        RECT 37.352 270.092 37.424 270.284 ; 
        RECT 65.432 270.092 65.504 270.284 ; 
        RECT 0.632 274.412 0.704 274.604 ; 
        RECT 28.712 274.412 28.784 274.604 ; 
        RECT 33.68 274.412 33.788 274.604 ; 
        RECT 34.292 274.412 34.436 274.604 ; 
        RECT 37.352 274.412 37.424 274.604 ; 
        RECT 65.432 274.412 65.504 274.604 ; 
        RECT 0.632 278.732 0.704 278.924 ; 
        RECT 28.712 278.732 28.784 278.924 ; 
        RECT 33.68 278.732 33.788 278.924 ; 
        RECT 34.292 278.732 34.436 278.924 ; 
        RECT 37.352 278.732 37.424 278.924 ; 
        RECT 65.432 278.732 65.504 278.924 ; 
        RECT 0.632 283.052 0.704 283.244 ; 
        RECT 28.712 283.052 28.784 283.244 ; 
        RECT 33.68 283.052 33.788 283.244 ; 
        RECT 34.292 283.052 34.436 283.244 ; 
        RECT 37.352 283.052 37.424 283.244 ; 
        RECT 65.432 283.052 65.504 283.244 ; 
        RECT 0.632 287.372 0.704 287.564 ; 
        RECT 28.712 287.372 28.784 287.564 ; 
        RECT 33.68 287.372 33.788 287.564 ; 
        RECT 34.292 287.372 34.436 287.564 ; 
        RECT 37.352 287.372 37.424 287.564 ; 
        RECT 65.432 287.372 65.504 287.564 ; 
        RECT 0.632 291.692 0.704 291.884 ; 
        RECT 28.712 291.692 28.784 291.884 ; 
        RECT 33.68 291.692 33.788 291.884 ; 
        RECT 34.292 291.692 34.436 291.884 ; 
        RECT 37.352 291.692 37.424 291.884 ; 
        RECT 65.432 291.692 65.504 291.884 ; 
        RECT 0.632 296.012 0.704 296.204 ; 
        RECT 28.712 296.012 28.784 296.204 ; 
        RECT 33.68 296.012 33.788 296.204 ; 
        RECT 34.292 296.012 34.436 296.204 ; 
        RECT 37.352 296.012 37.424 296.204 ; 
        RECT 65.432 296.012 65.504 296.204 ; 
        RECT 0.632 300.332 0.704 300.524 ; 
        RECT 28.712 300.332 28.784 300.524 ; 
        RECT 33.68 300.332 33.788 300.524 ; 
        RECT 34.292 300.332 34.436 300.524 ; 
        RECT 37.352 300.332 37.424 300.524 ; 
        RECT 65.432 300.332 65.504 300.524 ; 
        RECT 0.632 304.652 0.704 304.844 ; 
        RECT 28.712 304.652 28.784 304.844 ; 
        RECT 33.68 304.652 33.788 304.844 ; 
        RECT 34.292 304.652 34.436 304.844 ; 
        RECT 37.352 304.652 37.424 304.844 ; 
        RECT 65.432 304.652 65.504 304.844 ; 
        RECT 0.632 308.972 0.704 309.164 ; 
        RECT 28.712 308.972 28.784 309.164 ; 
        RECT 33.68 308.972 33.788 309.164 ; 
        RECT 34.292 308.972 34.436 309.164 ; 
        RECT 37.352 308.972 37.424 309.164 ; 
        RECT 65.432 308.972 65.504 309.164 ; 
        RECT 0.632 313.292 0.704 313.484 ; 
        RECT 28.712 313.292 28.784 313.484 ; 
        RECT 33.68 313.292 33.788 313.484 ; 
        RECT 34.292 313.292 34.436 313.484 ; 
        RECT 37.352 313.292 37.424 313.484 ; 
        RECT 65.432 313.292 65.504 313.484 ; 
        RECT 0.632 317.612 0.704 317.804 ; 
        RECT 28.712 317.612 28.784 317.804 ; 
        RECT 33.68 317.612 33.788 317.804 ; 
        RECT 34.292 317.612 34.436 317.804 ; 
        RECT 37.352 317.612 37.424 317.804 ; 
        RECT 65.432 317.612 65.504 317.804 ; 
        RECT 0.632 321.932 0.704 322.124 ; 
        RECT 28.712 321.932 28.784 322.124 ; 
        RECT 33.68 321.932 33.788 322.124 ; 
        RECT 34.292 321.932 34.436 322.124 ; 
        RECT 37.352 321.932 37.424 322.124 ; 
        RECT 65.432 321.932 65.504 322.124 ; 
        RECT 0.632 326.252 0.704 326.444 ; 
        RECT 28.712 326.252 28.784 326.444 ; 
        RECT 33.68 326.252 33.788 326.444 ; 
        RECT 34.292 326.252 34.436 326.444 ; 
        RECT 37.352 326.252 37.424 326.444 ; 
        RECT 65.432 326.252 65.504 326.444 ; 
        RECT 0.632 330.572 0.704 330.764 ; 
        RECT 28.712 330.572 28.784 330.764 ; 
        RECT 33.68 330.572 33.788 330.764 ; 
        RECT 34.292 330.572 34.436 330.764 ; 
        RECT 37.352 330.572 37.424 330.764 ; 
        RECT 65.432 330.572 65.504 330.764 ; 
        RECT 0.632 334.892 0.704 335.084 ; 
        RECT 28.712 334.892 28.784 335.084 ; 
        RECT 33.68 334.892 33.788 335.084 ; 
        RECT 34.292 334.892 34.436 335.084 ; 
        RECT 37.352 334.892 37.424 335.084 ; 
        RECT 65.432 334.892 65.504 335.084 ; 
        RECT 0.632 339.212 0.704 339.404 ; 
        RECT 28.712 339.212 28.784 339.404 ; 
        RECT 33.68 339.212 33.788 339.404 ; 
        RECT 34.292 339.212 34.436 339.404 ; 
        RECT 37.352 339.212 37.424 339.404 ; 
        RECT 65.432 339.212 65.504 339.404 ; 
        RECT 0.632 343.532 0.704 343.724 ; 
        RECT 28.712 343.532 28.784 343.724 ; 
        RECT 33.68 343.532 33.788 343.724 ; 
        RECT 34.292 343.532 34.436 343.724 ; 
        RECT 37.352 343.532 37.424 343.724 ; 
        RECT 65.432 343.532 65.504 343.724 ; 
        RECT 0.632 347.852 0.704 348.044 ; 
        RECT 28.712 347.852 28.784 348.044 ; 
        RECT 33.68 347.852 33.788 348.044 ; 
        RECT 34.292 347.852 34.436 348.044 ; 
        RECT 37.352 347.852 37.424 348.044 ; 
        RECT 65.432 347.852 65.504 348.044 ; 
        RECT 0.632 352.172 0.704 352.364 ; 
        RECT 28.712 352.172 28.784 352.364 ; 
        RECT 33.68 352.172 33.788 352.364 ; 
        RECT 34.292 352.172 34.436 352.364 ; 
        RECT 37.352 352.172 37.424 352.364 ; 
        RECT 65.432 352.172 65.504 352.364 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 43.164 165.748 43.236 165.896 ; 
      LAYER M4 ; 
        RECT 42.956 165.78 43.292 165.876 ; 
      LAYER M5 ; 
        RECT 43.152 161.976 43.248 174.936 ; 
      LAYER V3 ; 
        RECT 43.164 165.78 43.236 165.876 ; 
      LAYER V4 ; 
        RECT 43.152 165.78 43.248 165.876 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 42.3 165.76 42.372 165.908 ; 
      LAYER M4 ; 
        RECT 42.092 165.78 42.428 165.876 ; 
      LAYER M5 ; 
        RECT 42.288 161.976 42.384 174.936 ; 
      LAYER V3 ; 
        RECT 42.3 165.78 42.372 165.876 ; 
      LAYER V4 ; 
        RECT 42.288 165.78 42.384 165.876 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 41.436 163.444 41.508 163.592 ; 
      LAYER M4 ; 
        RECT 41.228 163.476 41.564 163.572 ; 
      LAYER M5 ; 
        RECT 41.424 161.976 41.52 174.936 ; 
      LAYER V3 ; 
        RECT 41.436 163.476 41.508 163.572 ; 
      LAYER V4 ; 
        RECT 41.424 163.476 41.52 163.572 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 40.572 164.404 40.644 165.128 ; 
      LAYER M4 ; 
        RECT 40.364 165.012 40.7 165.108 ; 
      LAYER M5 ; 
        RECT 40.56 161.976 40.656 174.936 ; 
      LAYER V3 ; 
        RECT 40.572 165.012 40.644 165.108 ; 
      LAYER V4 ; 
        RECT 40.56 165.012 40.656 165.108 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 39.708 163.456 39.78 163.724 ; 
      LAYER M4 ; 
        RECT 39.5 163.476 39.836 163.572 ; 
      LAYER M5 ; 
        RECT 39.696 161.976 39.792 174.936 ; 
      LAYER V3 ; 
        RECT 39.708 163.476 39.78 163.572 ; 
      LAYER V4 ; 
        RECT 39.696 163.476 39.792 163.572 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 38.844 162.388 38.916 163.4 ; 
      LAYER M4 ; 
        RECT 38.636 163.284 38.972 163.38 ; 
      LAYER M5 ; 
        RECT 38.832 161.976 38.928 174.936 ; 
      LAYER V3 ; 
        RECT 38.844 163.284 38.916 163.38 ; 
      LAYER V4 ; 
        RECT 38.832 163.284 38.928 163.38 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.98 166.528 38.052 166.676 ; 
      LAYER M4 ; 
        RECT 37.772 166.548 38.108 166.644 ; 
      LAYER M5 ; 
        RECT 37.968 161.976 38.064 174.936 ; 
      LAYER V3 ; 
        RECT 37.98 166.548 38.052 166.644 ; 
      LAYER V4 ; 
        RECT 37.968 166.548 38.064 166.644 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.116 165.916 37.188 166.28 ; 
      LAYER M4 ; 
        RECT 36.908 166.164 37.244 166.26 ; 
      LAYER M5 ; 
        RECT 37.104 161.976 37.2 174.936 ; 
      LAYER V3 ; 
        RECT 37.116 166.164 37.188 166.26 ; 
      LAYER V4 ; 
        RECT 37.104 166.164 37.2 166.26 ; 
    END 
  END ADDRESS[7] 
  PIN ADDRESS[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 34.524 163.456 34.596 163.724 ; 
      LAYER M4 ; 
        RECT 33.388 163.476 34.64 163.572 ; 
      LAYER M5 ; 
        RECT 33.432 161.976 33.528 174.936 ; 
      LAYER V3 ; 
        RECT 34.524 163.476 34.596 163.572 ; 
      LAYER V4 ; 
        RECT 33.432 163.476 33.528 163.572 ; 
    END 
  END ADDRESS[8] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 32.94 162.388 33.012 163.4 ; 
      LAYER M4 ; 
        RECT 32.092 163.284 33.056 163.38 ; 
      LAYER M5 ; 
        RECT 32.136 161.976 32.232 174.936 ; 
      LAYER V3 ; 
        RECT 32.94 163.284 33.012 163.38 ; 
      LAYER V4 ; 
        RECT 32.136 163.284 32.232 163.38 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.772 163.456 29.844 163.724 ; 
      LAYER M4 ; 
        RECT 29.564 163.476 29.9 163.572 ; 
      LAYER M5 ; 
        RECT 29.76 161.976 29.856 174.936 ; 
      LAYER V3 ; 
        RECT 29.772 163.476 29.844 163.572 ; 
      LAYER V4 ; 
        RECT 29.76 163.476 29.856 163.572 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.908 166.912 28.98 167.108 ; 
      LAYER M4 ; 
        RECT 28.7 166.932 29.036 167.028 ; 
      LAYER M5 ; 
        RECT 28.896 161.976 28.992 174.936 ; 
      LAYER V3 ; 
        RECT 28.908 166.932 28.98 167.028 ; 
      LAYER V4 ; 
        RECT 28.896 166.932 28.992 167.028 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.052 162.388 29.124 163.4 ; 
      LAYER M4 ; 
        RECT 27.988 163.284 29.168 163.38 ; 
      LAYER M5 ; 
        RECT 28.032 161.976 28.128 174.936 ; 
      LAYER V3 ; 
        RECT 29.052 163.284 29.124 163.38 ; 
      LAYER V4 ; 
        RECT 28.032 163.284 28.128 163.38 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.18 165.748 27.252 165.896 ; 
      LAYER M4 ; 
        RECT 26.972 165.78 27.308 165.876 ; 
      LAYER M5 ; 
        RECT 27.168 161.976 27.264 174.936 ; 
      LAYER V3 ; 
        RECT 27.18 165.78 27.252 165.876 ; 
      LAYER V4 ; 
        RECT 27.168 165.78 27.264 165.876 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.316 163.456 26.388 164.372 ; 
      LAYER M4 ; 
        RECT 26.108 163.476 26.444 163.572 ; 
      LAYER M5 ; 
        RECT 26.304 161.976 26.4 174.936 ; 
      LAYER V3 ; 
        RECT 26.316 163.476 26.388 163.572 ; 
      LAYER V4 ; 
        RECT 26.304 163.476 26.4 163.572 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.452 162.388 25.524 163.4 ; 
      LAYER M4 ; 
        RECT 25.244 163.284 25.58 163.38 ; 
      LAYER M5 ; 
        RECT 25.44 161.976 25.536 174.936 ; 
      LAYER V3 ; 
        RECT 25.452 163.284 25.524 163.38 ; 
      LAYER V4 ; 
        RECT 25.44 163.284 25.536 163.38 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.588 163.444 24.66 163.592 ; 
      LAYER M4 ; 
        RECT 24.38 163.476 24.716 163.572 ; 
      LAYER M5 ; 
        RECT 24.576 161.976 24.672 174.936 ; 
      LAYER V3 ; 
        RECT 24.588 163.476 24.66 163.572 ; 
      LAYER V4 ; 
        RECT 24.576 163.476 24.672 163.572 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 23.724 165.748 23.796 165.896 ; 
      LAYER M4 ; 
        RECT 23.516 165.78 23.852 165.876 ; 
      LAYER M5 ; 
        RECT 23.712 161.976 23.808 174.936 ; 
      LAYER V3 ; 
        RECT 23.724 165.78 23.796 165.876 ; 
      LAYER V4 ; 
        RECT 23.712 165.78 23.808 165.876 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.712 34.388 1.808 ; 
      LAYER M3 ; 
        RECT 34.148 1.51 34.22 2.468 ; 
      LAYER V3 ; 
        RECT 34.148 1.712 34.22 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.328 34.66 1.424 ; 
      LAYER M3 ; 
        RECT 33.248 1.08 33.32 2.7 ; 
      LAYER V3 ; 
        RECT 33.248 1.328 33.32 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 6.032 34.388 6.128 ; 
      LAYER M3 ; 
        RECT 34.148 5.83 34.22 6.788 ; 
      LAYER V3 ; 
        RECT 34.148 6.032 34.22 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 5.648 34.66 5.744 ; 
      LAYER M3 ; 
        RECT 33.248 5.4 33.32 7.02 ; 
      LAYER V3 ; 
        RECT 33.248 5.648 33.32 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 10.352 34.388 10.448 ; 
      LAYER M3 ; 
        RECT 34.148 10.15 34.22 11.108 ; 
      LAYER V3 ; 
        RECT 34.148 10.352 34.22 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 9.968 34.66 10.064 ; 
      LAYER M3 ; 
        RECT 33.248 9.72 33.32 11.34 ; 
      LAYER V3 ; 
        RECT 33.248 9.968 33.32 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.672 34.388 14.768 ; 
      LAYER M3 ; 
        RECT 34.148 14.47 34.22 15.428 ; 
      LAYER V3 ; 
        RECT 34.148 14.672 34.22 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.288 34.66 14.384 ; 
      LAYER M3 ; 
        RECT 33.248 14.04 33.32 15.66 ; 
      LAYER V3 ; 
        RECT 33.248 14.288 33.32 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.992 34.388 19.088 ; 
      LAYER M3 ; 
        RECT 34.148 18.79 34.22 19.748 ; 
      LAYER V3 ; 
        RECT 34.148 18.992 34.22 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.608 34.66 18.704 ; 
      LAYER M3 ; 
        RECT 33.248 18.36 33.32 19.98 ; 
      LAYER V3 ; 
        RECT 33.248 18.608 33.32 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 23.312 34.388 23.408 ; 
      LAYER M3 ; 
        RECT 34.148 23.11 34.22 24.068 ; 
      LAYER V3 ; 
        RECT 34.148 23.312 34.22 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 22.928 34.66 23.024 ; 
      LAYER M3 ; 
        RECT 33.248 22.68 33.32 24.3 ; 
      LAYER V3 ; 
        RECT 33.248 22.928 33.32 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.632 34.388 27.728 ; 
      LAYER M3 ; 
        RECT 34.148 27.43 34.22 28.388 ; 
      LAYER V3 ; 
        RECT 34.148 27.632 34.22 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.248 34.66 27.344 ; 
      LAYER M3 ; 
        RECT 33.248 27 33.32 28.62 ; 
      LAYER V3 ; 
        RECT 33.248 27.248 33.32 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.952 34.388 32.048 ; 
      LAYER M3 ; 
        RECT 34.148 31.75 34.22 32.708 ; 
      LAYER V3 ; 
        RECT 34.148 31.952 34.22 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.568 34.66 31.664 ; 
      LAYER M3 ; 
        RECT 33.248 31.32 33.32 32.94 ; 
      LAYER V3 ; 
        RECT 33.248 31.568 33.32 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 36.272 34.388 36.368 ; 
      LAYER M3 ; 
        RECT 34.148 36.07 34.22 37.028 ; 
      LAYER V3 ; 
        RECT 34.148 36.272 34.22 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 35.888 34.66 35.984 ; 
      LAYER M3 ; 
        RECT 33.248 35.64 33.32 37.26 ; 
      LAYER V3 ; 
        RECT 33.248 35.888 33.32 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.592 34.388 40.688 ; 
      LAYER M3 ; 
        RECT 34.148 40.39 34.22 41.348 ; 
      LAYER V3 ; 
        RECT 34.148 40.592 34.22 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.208 34.66 40.304 ; 
      LAYER M3 ; 
        RECT 33.248 39.96 33.32 41.58 ; 
      LAYER V3 ; 
        RECT 33.248 40.208 33.32 40.304 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 44.912 34.388 45.008 ; 
      LAYER M3 ; 
        RECT 34.148 44.71 34.22 45.668 ; 
      LAYER V3 ; 
        RECT 34.148 44.912 34.22 45.008 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 44.528 34.66 44.624 ; 
      LAYER M3 ; 
        RECT 33.248 44.28 33.32 45.9 ; 
      LAYER V3 ; 
        RECT 33.248 44.528 33.32 44.624 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 49.232 34.388 49.328 ; 
      LAYER M3 ; 
        RECT 34.148 49.03 34.22 49.988 ; 
      LAYER V3 ; 
        RECT 34.148 49.232 34.22 49.328 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 48.848 34.66 48.944 ; 
      LAYER M3 ; 
        RECT 33.248 48.6 33.32 50.22 ; 
      LAYER V3 ; 
        RECT 33.248 48.848 33.32 48.944 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 53.552 34.388 53.648 ; 
      LAYER M3 ; 
        RECT 34.148 53.35 34.22 54.308 ; 
      LAYER V3 ; 
        RECT 34.148 53.552 34.22 53.648 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 53.168 34.66 53.264 ; 
      LAYER M3 ; 
        RECT 33.248 52.92 33.32 54.54 ; 
      LAYER V3 ; 
        RECT 33.248 53.168 33.32 53.264 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 57.872 34.388 57.968 ; 
      LAYER M3 ; 
        RECT 34.148 57.67 34.22 58.628 ; 
      LAYER V3 ; 
        RECT 34.148 57.872 34.22 57.968 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 57.488 34.66 57.584 ; 
      LAYER M3 ; 
        RECT 33.248 57.24 33.32 58.86 ; 
      LAYER V3 ; 
        RECT 33.248 57.488 33.32 57.584 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 62.192 34.388 62.288 ; 
      LAYER M3 ; 
        RECT 34.148 61.99 34.22 62.948 ; 
      LAYER V3 ; 
        RECT 34.148 62.192 34.22 62.288 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 61.808 34.66 61.904 ; 
      LAYER M3 ; 
        RECT 33.248 61.56 33.32 63.18 ; 
      LAYER V3 ; 
        RECT 33.248 61.808 33.32 61.904 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 66.512 34.388 66.608 ; 
      LAYER M3 ; 
        RECT 34.148 66.31 34.22 67.268 ; 
      LAYER V3 ; 
        RECT 34.148 66.512 34.22 66.608 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 66.128 34.66 66.224 ; 
      LAYER M3 ; 
        RECT 33.248 65.88 33.32 67.5 ; 
      LAYER V3 ; 
        RECT 33.248 66.128 33.32 66.224 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 70.832 34.388 70.928 ; 
      LAYER M3 ; 
        RECT 34.148 70.63 34.22 71.588 ; 
      LAYER V3 ; 
        RECT 34.148 70.832 34.22 70.928 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 70.448 34.66 70.544 ; 
      LAYER M3 ; 
        RECT 33.248 70.2 33.32 71.82 ; 
      LAYER V3 ; 
        RECT 33.248 70.448 33.32 70.544 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 75.152 34.388 75.248 ; 
      LAYER M3 ; 
        RECT 34.148 74.95 34.22 75.908 ; 
      LAYER V3 ; 
        RECT 34.148 75.152 34.22 75.248 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 74.768 34.66 74.864 ; 
      LAYER M3 ; 
        RECT 33.248 74.52 33.32 76.14 ; 
      LAYER V3 ; 
        RECT 33.248 74.768 33.32 74.864 ; 
    END 
  END wd[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 79.472 34.388 79.568 ; 
      LAYER M3 ; 
        RECT 34.148 79.27 34.22 80.228 ; 
      LAYER V3 ; 
        RECT 34.148 79.472 34.22 79.568 ; 
    END 
  END dataout[18] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 79.088 34.66 79.184 ; 
      LAYER M3 ; 
        RECT 33.248 78.84 33.32 80.46 ; 
      LAYER V3 ; 
        RECT 33.248 79.088 33.32 79.184 ; 
    END 
  END wd[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 83.792 34.388 83.888 ; 
      LAYER M3 ; 
        RECT 34.148 83.59 34.22 84.548 ; 
      LAYER V3 ; 
        RECT 34.148 83.792 34.22 83.888 ; 
    END 
  END dataout[19] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 83.408 34.66 83.504 ; 
      LAYER M3 ; 
        RECT 33.248 83.16 33.32 84.78 ; 
      LAYER V3 ; 
        RECT 33.248 83.408 33.32 83.504 ; 
    END 
  END wd[19] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 88.112 34.388 88.208 ; 
      LAYER M3 ; 
        RECT 34.148 87.91 34.22 88.868 ; 
      LAYER V3 ; 
        RECT 34.148 88.112 34.22 88.208 ; 
    END 
  END dataout[20] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 87.728 34.66 87.824 ; 
      LAYER M3 ; 
        RECT 33.248 87.48 33.32 89.1 ; 
      LAYER V3 ; 
        RECT 33.248 87.728 33.32 87.824 ; 
    END 
  END wd[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 92.432 34.388 92.528 ; 
      LAYER M3 ; 
        RECT 34.148 92.23 34.22 93.188 ; 
      LAYER V3 ; 
        RECT 34.148 92.432 34.22 92.528 ; 
    END 
  END dataout[21] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 92.048 34.66 92.144 ; 
      LAYER M3 ; 
        RECT 33.248 91.8 33.32 93.42 ; 
      LAYER V3 ; 
        RECT 33.248 92.048 33.32 92.144 ; 
    END 
  END wd[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 96.752 34.388 96.848 ; 
      LAYER M3 ; 
        RECT 34.148 96.55 34.22 97.508 ; 
      LAYER V3 ; 
        RECT 34.148 96.752 34.22 96.848 ; 
    END 
  END dataout[22] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 96.368 34.66 96.464 ; 
      LAYER M3 ; 
        RECT 33.248 96.12 33.32 97.74 ; 
      LAYER V3 ; 
        RECT 33.248 96.368 33.32 96.464 ; 
    END 
  END wd[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 101.072 34.388 101.168 ; 
      LAYER M3 ; 
        RECT 34.148 100.87 34.22 101.828 ; 
      LAYER V3 ; 
        RECT 34.148 101.072 34.22 101.168 ; 
    END 
  END dataout[23] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 100.688 34.66 100.784 ; 
      LAYER M3 ; 
        RECT 33.248 100.44 33.32 102.06 ; 
      LAYER V3 ; 
        RECT 33.248 100.688 33.32 100.784 ; 
    END 
  END wd[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 105.392 34.388 105.488 ; 
      LAYER M3 ; 
        RECT 34.148 105.19 34.22 106.148 ; 
      LAYER V3 ; 
        RECT 34.148 105.392 34.22 105.488 ; 
    END 
  END dataout[24] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 105.008 34.66 105.104 ; 
      LAYER M3 ; 
        RECT 33.248 104.76 33.32 106.38 ; 
      LAYER V3 ; 
        RECT 33.248 105.008 33.32 105.104 ; 
    END 
  END wd[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 109.712 34.388 109.808 ; 
      LAYER M3 ; 
        RECT 34.148 109.51 34.22 110.468 ; 
      LAYER V3 ; 
        RECT 34.148 109.712 34.22 109.808 ; 
    END 
  END dataout[25] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 109.328 34.66 109.424 ; 
      LAYER M3 ; 
        RECT 33.248 109.08 33.32 110.7 ; 
      LAYER V3 ; 
        RECT 33.248 109.328 33.32 109.424 ; 
    END 
  END wd[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 114.032 34.388 114.128 ; 
      LAYER M3 ; 
        RECT 34.148 113.83 34.22 114.788 ; 
      LAYER V3 ; 
        RECT 34.148 114.032 34.22 114.128 ; 
    END 
  END dataout[26] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 113.648 34.66 113.744 ; 
      LAYER M3 ; 
        RECT 33.248 113.4 33.32 115.02 ; 
      LAYER V3 ; 
        RECT 33.248 113.648 33.32 113.744 ; 
    END 
  END wd[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 118.352 34.388 118.448 ; 
      LAYER M3 ; 
        RECT 34.148 118.15 34.22 119.108 ; 
      LAYER V3 ; 
        RECT 34.148 118.352 34.22 118.448 ; 
    END 
  END dataout[27] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 117.968 34.66 118.064 ; 
      LAYER M3 ; 
        RECT 33.248 117.72 33.32 119.34 ; 
      LAYER V3 ; 
        RECT 33.248 117.968 33.32 118.064 ; 
    END 
  END wd[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 122.672 34.388 122.768 ; 
      LAYER M3 ; 
        RECT 34.148 122.47 34.22 123.428 ; 
      LAYER V3 ; 
        RECT 34.148 122.672 34.22 122.768 ; 
    END 
  END dataout[28] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 122.288 34.66 122.384 ; 
      LAYER M3 ; 
        RECT 33.248 122.04 33.32 123.66 ; 
      LAYER V3 ; 
        RECT 33.248 122.288 33.32 122.384 ; 
    END 
  END wd[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 126.992 34.388 127.088 ; 
      LAYER M3 ; 
        RECT 34.148 126.79 34.22 127.748 ; 
      LAYER V3 ; 
        RECT 34.148 126.992 34.22 127.088 ; 
    END 
  END dataout[29] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 126.608 34.66 126.704 ; 
      LAYER M3 ; 
        RECT 33.248 126.36 33.32 127.98 ; 
      LAYER V3 ; 
        RECT 33.248 126.608 33.32 126.704 ; 
    END 
  END wd[29] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 131.312 34.388 131.408 ; 
      LAYER M3 ; 
        RECT 34.148 131.11 34.22 132.068 ; 
      LAYER V3 ; 
        RECT 34.148 131.312 34.22 131.408 ; 
    END 
  END dataout[30] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 130.928 34.66 131.024 ; 
      LAYER M3 ; 
        RECT 33.248 130.68 33.32 132.3 ; 
      LAYER V3 ; 
        RECT 33.248 130.928 33.32 131.024 ; 
    END 
  END wd[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 135.632 34.388 135.728 ; 
      LAYER M3 ; 
        RECT 34.148 135.43 34.22 136.388 ; 
      LAYER V3 ; 
        RECT 34.148 135.632 34.22 135.728 ; 
    END 
  END dataout[31] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 135.248 34.66 135.344 ; 
      LAYER M3 ; 
        RECT 33.248 135 33.32 136.62 ; 
      LAYER V3 ; 
        RECT 33.248 135.248 33.32 135.344 ; 
    END 
  END wd[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 139.952 34.388 140.048 ; 
      LAYER M3 ; 
        RECT 34.148 139.75 34.22 140.708 ; 
      LAYER V3 ; 
        RECT 34.148 139.952 34.22 140.048 ; 
    END 
  END dataout[32] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 139.568 34.66 139.664 ; 
      LAYER M3 ; 
        RECT 33.248 139.32 33.32 140.94 ; 
      LAYER V3 ; 
        RECT 33.248 139.568 33.32 139.664 ; 
    END 
  END wd[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 144.272 34.388 144.368 ; 
      LAYER M3 ; 
        RECT 34.148 144.07 34.22 145.028 ; 
      LAYER V3 ; 
        RECT 34.148 144.272 34.22 144.368 ; 
    END 
  END dataout[33] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 143.888 34.66 143.984 ; 
      LAYER M3 ; 
        RECT 33.248 143.64 33.32 145.26 ; 
      LAYER V3 ; 
        RECT 33.248 143.888 33.32 143.984 ; 
    END 
  END wd[33] 
  PIN dataout[34] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 148.592 34.388 148.688 ; 
      LAYER M3 ; 
        RECT 34.148 148.39 34.22 149.348 ; 
      LAYER V3 ; 
        RECT 34.148 148.592 34.22 148.688 ; 
    END 
  END dataout[34] 
  PIN wd[34] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 148.208 34.66 148.304 ; 
      LAYER M3 ; 
        RECT 33.248 147.96 33.32 149.58 ; 
      LAYER V3 ; 
        RECT 33.248 148.208 33.32 148.304 ; 
    END 
  END wd[34] 
  PIN dataout[35] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 152.912 34.388 153.008 ; 
      LAYER M3 ; 
        RECT 34.148 152.71 34.22 153.668 ; 
      LAYER V3 ; 
        RECT 34.148 152.912 34.22 153.008 ; 
    END 
  END dataout[35] 
  PIN wd[35] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 152.528 34.66 152.624 ; 
      LAYER M3 ; 
        RECT 33.248 152.28 33.32 153.9 ; 
      LAYER V3 ; 
        RECT 33.248 152.528 33.32 152.624 ; 
    END 
  END wd[35] 
  PIN dataout[36] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 157.232 34.388 157.328 ; 
      LAYER M3 ; 
        RECT 34.148 157.03 34.22 157.988 ; 
      LAYER V3 ; 
        RECT 34.148 157.232 34.22 157.328 ; 
    END 
  END dataout[36] 
  PIN wd[36] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 156.848 34.66 156.944 ; 
      LAYER M3 ; 
        RECT 33.248 156.6 33.32 158.22 ; 
      LAYER V3 ; 
        RECT 33.248 156.848 33.32 156.944 ; 
    END 
  END wd[36] 
  PIN dataout[37] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 194.06 34.388 194.156 ; 
      LAYER M3 ; 
        RECT 34.148 193.858 34.22 194.816 ; 
      LAYER V3 ; 
        RECT 34.148 194.06 34.22 194.156 ; 
    END 
  END dataout[37] 
  PIN wd[37] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 193.676 34.66 193.772 ; 
      LAYER M3 ; 
        RECT 33.248 193.428 33.32 195.048 ; 
      LAYER V3 ; 
        RECT 33.248 193.676 33.32 193.772 ; 
    END 
  END wd[37] 
  PIN dataout[38] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 198.38 34.388 198.476 ; 
      LAYER M3 ; 
        RECT 34.148 198.178 34.22 199.136 ; 
      LAYER V3 ; 
        RECT 34.148 198.38 34.22 198.476 ; 
    END 
  END dataout[38] 
  PIN wd[38] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 197.996 34.66 198.092 ; 
      LAYER M3 ; 
        RECT 33.248 197.748 33.32 199.368 ; 
      LAYER V3 ; 
        RECT 33.248 197.996 33.32 198.092 ; 
    END 
  END wd[38] 
  PIN dataout[39] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 202.7 34.388 202.796 ; 
      LAYER M3 ; 
        RECT 34.148 202.498 34.22 203.456 ; 
      LAYER V3 ; 
        RECT 34.148 202.7 34.22 202.796 ; 
    END 
  END dataout[39] 
  PIN wd[39] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 202.316 34.66 202.412 ; 
      LAYER M3 ; 
        RECT 33.248 202.068 33.32 203.688 ; 
      LAYER V3 ; 
        RECT 33.248 202.316 33.32 202.412 ; 
    END 
  END wd[39] 
  PIN dataout[40] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 207.02 34.388 207.116 ; 
      LAYER M3 ; 
        RECT 34.148 206.818 34.22 207.776 ; 
      LAYER V3 ; 
        RECT 34.148 207.02 34.22 207.116 ; 
    END 
  END dataout[40] 
  PIN wd[40] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 206.636 34.66 206.732 ; 
      LAYER M3 ; 
        RECT 33.248 206.388 33.32 208.008 ; 
      LAYER V3 ; 
        RECT 33.248 206.636 33.32 206.732 ; 
    END 
  END wd[40] 
  PIN dataout[41] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 211.34 34.388 211.436 ; 
      LAYER M3 ; 
        RECT 34.148 211.138 34.22 212.096 ; 
      LAYER V3 ; 
        RECT 34.148 211.34 34.22 211.436 ; 
    END 
  END dataout[41] 
  PIN wd[41] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 210.956 34.66 211.052 ; 
      LAYER M3 ; 
        RECT 33.248 210.708 33.32 212.328 ; 
      LAYER V3 ; 
        RECT 33.248 210.956 33.32 211.052 ; 
    END 
  END wd[41] 
  PIN dataout[42] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 215.66 34.388 215.756 ; 
      LAYER M3 ; 
        RECT 34.148 215.458 34.22 216.416 ; 
      LAYER V3 ; 
        RECT 34.148 215.66 34.22 215.756 ; 
    END 
  END dataout[42] 
  PIN wd[42] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 215.276 34.66 215.372 ; 
      LAYER M3 ; 
        RECT 33.248 215.028 33.32 216.648 ; 
      LAYER V3 ; 
        RECT 33.248 215.276 33.32 215.372 ; 
    END 
  END wd[42] 
  PIN dataout[43] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 219.98 34.388 220.076 ; 
      LAYER M3 ; 
        RECT 34.148 219.778 34.22 220.736 ; 
      LAYER V3 ; 
        RECT 34.148 219.98 34.22 220.076 ; 
    END 
  END dataout[43] 
  PIN wd[43] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 219.596 34.66 219.692 ; 
      LAYER M3 ; 
        RECT 33.248 219.348 33.32 220.968 ; 
      LAYER V3 ; 
        RECT 33.248 219.596 33.32 219.692 ; 
    END 
  END wd[43] 
  PIN dataout[44] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 224.3 34.388 224.396 ; 
      LAYER M3 ; 
        RECT 34.148 224.098 34.22 225.056 ; 
      LAYER V3 ; 
        RECT 34.148 224.3 34.22 224.396 ; 
    END 
  END dataout[44] 
  PIN wd[44] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 223.916 34.66 224.012 ; 
      LAYER M3 ; 
        RECT 33.248 223.668 33.32 225.288 ; 
      LAYER V3 ; 
        RECT 33.248 223.916 33.32 224.012 ; 
    END 
  END wd[44] 
  PIN dataout[45] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 228.62 34.388 228.716 ; 
      LAYER M3 ; 
        RECT 34.148 228.418 34.22 229.376 ; 
      LAYER V3 ; 
        RECT 34.148 228.62 34.22 228.716 ; 
    END 
  END dataout[45] 
  PIN wd[45] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 228.236 34.66 228.332 ; 
      LAYER M3 ; 
        RECT 33.248 227.988 33.32 229.608 ; 
      LAYER V3 ; 
        RECT 33.248 228.236 33.32 228.332 ; 
    END 
  END wd[45] 
  PIN dataout[46] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 232.94 34.388 233.036 ; 
      LAYER M3 ; 
        RECT 34.148 232.738 34.22 233.696 ; 
      LAYER V3 ; 
        RECT 34.148 232.94 34.22 233.036 ; 
    END 
  END dataout[46] 
  PIN wd[46] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 232.556 34.66 232.652 ; 
      LAYER M3 ; 
        RECT 33.248 232.308 33.32 233.928 ; 
      LAYER V3 ; 
        RECT 33.248 232.556 33.32 232.652 ; 
    END 
  END wd[46] 
  PIN dataout[47] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 237.26 34.388 237.356 ; 
      LAYER M3 ; 
        RECT 34.148 237.058 34.22 238.016 ; 
      LAYER V3 ; 
        RECT 34.148 237.26 34.22 237.356 ; 
    END 
  END dataout[47] 
  PIN wd[47] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 236.876 34.66 236.972 ; 
      LAYER M3 ; 
        RECT 33.248 236.628 33.32 238.248 ; 
      LAYER V3 ; 
        RECT 33.248 236.876 33.32 236.972 ; 
    END 
  END wd[47] 
  PIN dataout[48] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 241.58 34.388 241.676 ; 
      LAYER M3 ; 
        RECT 34.148 241.378 34.22 242.336 ; 
      LAYER V3 ; 
        RECT 34.148 241.58 34.22 241.676 ; 
    END 
  END dataout[48] 
  PIN wd[48] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 241.196 34.66 241.292 ; 
      LAYER M3 ; 
        RECT 33.248 240.948 33.32 242.568 ; 
      LAYER V3 ; 
        RECT 33.248 241.196 33.32 241.292 ; 
    END 
  END wd[48] 
  PIN dataout[49] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 245.9 34.388 245.996 ; 
      LAYER M3 ; 
        RECT 34.148 245.698 34.22 246.656 ; 
      LAYER V3 ; 
        RECT 34.148 245.9 34.22 245.996 ; 
    END 
  END dataout[49] 
  PIN wd[49] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 245.516 34.66 245.612 ; 
      LAYER M3 ; 
        RECT 33.248 245.268 33.32 246.888 ; 
      LAYER V3 ; 
        RECT 33.248 245.516 33.32 245.612 ; 
    END 
  END wd[49] 
  PIN dataout[50] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 250.22 34.388 250.316 ; 
      LAYER M3 ; 
        RECT 34.148 250.018 34.22 250.976 ; 
      LAYER V3 ; 
        RECT 34.148 250.22 34.22 250.316 ; 
    END 
  END dataout[50] 
  PIN wd[50] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 249.836 34.66 249.932 ; 
      LAYER M3 ; 
        RECT 33.248 249.588 33.32 251.208 ; 
      LAYER V3 ; 
        RECT 33.248 249.836 33.32 249.932 ; 
    END 
  END wd[50] 
  PIN dataout[51] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 254.54 34.388 254.636 ; 
      LAYER M3 ; 
        RECT 34.148 254.338 34.22 255.296 ; 
      LAYER V3 ; 
        RECT 34.148 254.54 34.22 254.636 ; 
    END 
  END dataout[51] 
  PIN wd[51] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 254.156 34.66 254.252 ; 
      LAYER M3 ; 
        RECT 33.248 253.908 33.32 255.528 ; 
      LAYER V3 ; 
        RECT 33.248 254.156 33.32 254.252 ; 
    END 
  END wd[51] 
  PIN dataout[52] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 258.86 34.388 258.956 ; 
      LAYER M3 ; 
        RECT 34.148 258.658 34.22 259.616 ; 
      LAYER V3 ; 
        RECT 34.148 258.86 34.22 258.956 ; 
    END 
  END dataout[52] 
  PIN wd[52] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 258.476 34.66 258.572 ; 
      LAYER M3 ; 
        RECT 33.248 258.228 33.32 259.848 ; 
      LAYER V3 ; 
        RECT 33.248 258.476 33.32 258.572 ; 
    END 
  END wd[52] 
  PIN dataout[53] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 263.18 34.388 263.276 ; 
      LAYER M3 ; 
        RECT 34.148 262.978 34.22 263.936 ; 
      LAYER V3 ; 
        RECT 34.148 263.18 34.22 263.276 ; 
    END 
  END dataout[53] 
  PIN wd[53] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 262.796 34.66 262.892 ; 
      LAYER M3 ; 
        RECT 33.248 262.548 33.32 264.168 ; 
      LAYER V3 ; 
        RECT 33.248 262.796 33.32 262.892 ; 
    END 
  END wd[53] 
  PIN dataout[54] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 267.5 34.388 267.596 ; 
      LAYER M3 ; 
        RECT 34.148 267.298 34.22 268.256 ; 
      LAYER V3 ; 
        RECT 34.148 267.5 34.22 267.596 ; 
    END 
  END dataout[54] 
  PIN wd[54] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 267.116 34.66 267.212 ; 
      LAYER M3 ; 
        RECT 33.248 266.868 33.32 268.488 ; 
      LAYER V3 ; 
        RECT 33.248 267.116 33.32 267.212 ; 
    END 
  END wd[54] 
  PIN dataout[55] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 271.82 34.388 271.916 ; 
      LAYER M3 ; 
        RECT 34.148 271.618 34.22 272.576 ; 
      LAYER V3 ; 
        RECT 34.148 271.82 34.22 271.916 ; 
    END 
  END dataout[55] 
  PIN wd[55] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 271.436 34.66 271.532 ; 
      LAYER M3 ; 
        RECT 33.248 271.188 33.32 272.808 ; 
      LAYER V3 ; 
        RECT 33.248 271.436 33.32 271.532 ; 
    END 
  END wd[55] 
  PIN dataout[56] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 276.14 34.388 276.236 ; 
      LAYER M3 ; 
        RECT 34.148 275.938 34.22 276.896 ; 
      LAYER V3 ; 
        RECT 34.148 276.14 34.22 276.236 ; 
    END 
  END dataout[56] 
  PIN wd[56] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 275.756 34.66 275.852 ; 
      LAYER M3 ; 
        RECT 33.248 275.508 33.32 277.128 ; 
      LAYER V3 ; 
        RECT 33.248 275.756 33.32 275.852 ; 
    END 
  END wd[56] 
  PIN dataout[57] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 280.46 34.388 280.556 ; 
      LAYER M3 ; 
        RECT 34.148 280.258 34.22 281.216 ; 
      LAYER V3 ; 
        RECT 34.148 280.46 34.22 280.556 ; 
    END 
  END dataout[57] 
  PIN wd[57] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 280.076 34.66 280.172 ; 
      LAYER M3 ; 
        RECT 33.248 279.828 33.32 281.448 ; 
      LAYER V3 ; 
        RECT 33.248 280.076 33.32 280.172 ; 
    END 
  END wd[57] 
  PIN dataout[58] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 284.78 34.388 284.876 ; 
      LAYER M3 ; 
        RECT 34.148 284.578 34.22 285.536 ; 
      LAYER V3 ; 
        RECT 34.148 284.78 34.22 284.876 ; 
    END 
  END dataout[58] 
  PIN wd[58] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 284.396 34.66 284.492 ; 
      LAYER M3 ; 
        RECT 33.248 284.148 33.32 285.768 ; 
      LAYER V3 ; 
        RECT 33.248 284.396 33.32 284.492 ; 
    END 
  END wd[58] 
  PIN dataout[59] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 289.1 34.388 289.196 ; 
      LAYER M3 ; 
        RECT 34.148 288.898 34.22 289.856 ; 
      LAYER V3 ; 
        RECT 34.148 289.1 34.22 289.196 ; 
    END 
  END dataout[59] 
  PIN wd[59] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 288.716 34.66 288.812 ; 
      LAYER M3 ; 
        RECT 33.248 288.468 33.32 290.088 ; 
      LAYER V3 ; 
        RECT 33.248 288.716 33.32 288.812 ; 
    END 
  END wd[59] 
  PIN dataout[60] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 293.42 34.388 293.516 ; 
      LAYER M3 ; 
        RECT 34.148 293.218 34.22 294.176 ; 
      LAYER V3 ; 
        RECT 34.148 293.42 34.22 293.516 ; 
    END 
  END dataout[60] 
  PIN wd[60] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 293.036 34.66 293.132 ; 
      LAYER M3 ; 
        RECT 33.248 292.788 33.32 294.408 ; 
      LAYER V3 ; 
        RECT 33.248 293.036 33.32 293.132 ; 
    END 
  END wd[60] 
  PIN dataout[61] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 297.74 34.388 297.836 ; 
      LAYER M3 ; 
        RECT 34.148 297.538 34.22 298.496 ; 
      LAYER V3 ; 
        RECT 34.148 297.74 34.22 297.836 ; 
    END 
  END dataout[61] 
  PIN wd[61] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 297.356 34.66 297.452 ; 
      LAYER M3 ; 
        RECT 33.248 297.108 33.32 298.728 ; 
      LAYER V3 ; 
        RECT 33.248 297.356 33.32 297.452 ; 
    END 
  END wd[61] 
  PIN dataout[62] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 302.06 34.388 302.156 ; 
      LAYER M3 ; 
        RECT 34.148 301.858 34.22 302.816 ; 
      LAYER V3 ; 
        RECT 34.148 302.06 34.22 302.156 ; 
    END 
  END dataout[62] 
  PIN wd[62] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 301.676 34.66 301.772 ; 
      LAYER M3 ; 
        RECT 33.248 301.428 33.32 303.048 ; 
      LAYER V3 ; 
        RECT 33.248 301.676 33.32 301.772 ; 
    END 
  END wd[62] 
  PIN dataout[63] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 306.38 34.388 306.476 ; 
      LAYER M3 ; 
        RECT 34.148 306.178 34.22 307.136 ; 
      LAYER V3 ; 
        RECT 34.148 306.38 34.22 306.476 ; 
    END 
  END dataout[63] 
  PIN wd[63] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 305.996 34.66 306.092 ; 
      LAYER M3 ; 
        RECT 33.248 305.748 33.32 307.368 ; 
      LAYER V3 ; 
        RECT 33.248 305.996 33.32 306.092 ; 
    END 
  END wd[63] 
  PIN dataout[64] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 310.7 34.388 310.796 ; 
      LAYER M3 ; 
        RECT 34.148 310.498 34.22 311.456 ; 
      LAYER V3 ; 
        RECT 34.148 310.7 34.22 310.796 ; 
    END 
  END dataout[64] 
  PIN wd[64] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 310.316 34.66 310.412 ; 
      LAYER M3 ; 
        RECT 33.248 310.068 33.32 311.688 ; 
      LAYER V3 ; 
        RECT 33.248 310.316 33.32 310.412 ; 
    END 
  END wd[64] 
  PIN dataout[65] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 315.02 34.388 315.116 ; 
      LAYER M3 ; 
        RECT 34.148 314.818 34.22 315.776 ; 
      LAYER V3 ; 
        RECT 34.148 315.02 34.22 315.116 ; 
    END 
  END dataout[65] 
  PIN wd[65] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 314.636 34.66 314.732 ; 
      LAYER M3 ; 
        RECT 33.248 314.388 33.32 316.008 ; 
      LAYER V3 ; 
        RECT 33.248 314.636 33.32 314.732 ; 
    END 
  END wd[65] 
  PIN dataout[66] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 319.34 34.388 319.436 ; 
      LAYER M3 ; 
        RECT 34.148 319.138 34.22 320.096 ; 
      LAYER V3 ; 
        RECT 34.148 319.34 34.22 319.436 ; 
    END 
  END dataout[66] 
  PIN wd[66] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 318.956 34.66 319.052 ; 
      LAYER M3 ; 
        RECT 33.248 318.708 33.32 320.328 ; 
      LAYER V3 ; 
        RECT 33.248 318.956 33.32 319.052 ; 
    END 
  END wd[66] 
  PIN dataout[67] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 323.66 34.388 323.756 ; 
      LAYER M3 ; 
        RECT 34.148 323.458 34.22 324.416 ; 
      LAYER V3 ; 
        RECT 34.148 323.66 34.22 323.756 ; 
    END 
  END dataout[67] 
  PIN wd[67] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 323.276 34.66 323.372 ; 
      LAYER M3 ; 
        RECT 33.248 323.028 33.32 324.648 ; 
      LAYER V3 ; 
        RECT 33.248 323.276 33.32 323.372 ; 
    END 
  END wd[67] 
  PIN dataout[68] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 327.98 34.388 328.076 ; 
      LAYER M3 ; 
        RECT 34.148 327.778 34.22 328.736 ; 
      LAYER V3 ; 
        RECT 34.148 327.98 34.22 328.076 ; 
    END 
  END dataout[68] 
  PIN wd[68] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 327.596 34.66 327.692 ; 
      LAYER M3 ; 
        RECT 33.248 327.348 33.32 328.968 ; 
      LAYER V3 ; 
        RECT 33.248 327.596 33.32 327.692 ; 
    END 
  END wd[68] 
  PIN dataout[69] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 332.3 34.388 332.396 ; 
      LAYER M3 ; 
        RECT 34.148 332.098 34.22 333.056 ; 
      LAYER V3 ; 
        RECT 34.148 332.3 34.22 332.396 ; 
    END 
  END dataout[69] 
  PIN wd[69] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 331.916 34.66 332.012 ; 
      LAYER M3 ; 
        RECT 33.248 331.668 33.32 333.288 ; 
      LAYER V3 ; 
        RECT 33.248 331.916 33.32 332.012 ; 
    END 
  END wd[69] 
  PIN dataout[70] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 336.62 34.388 336.716 ; 
      LAYER M3 ; 
        RECT 34.148 336.418 34.22 337.376 ; 
      LAYER V3 ; 
        RECT 34.148 336.62 34.22 336.716 ; 
    END 
  END dataout[70] 
  PIN wd[70] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 336.236 34.66 336.332 ; 
      LAYER M3 ; 
        RECT 33.248 335.988 33.32 337.608 ; 
      LAYER V3 ; 
        RECT 33.248 336.236 33.32 336.332 ; 
    END 
  END wd[70] 
  PIN dataout[71] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 340.94 34.388 341.036 ; 
      LAYER M3 ; 
        RECT 34.148 340.738 34.22 341.696 ; 
      LAYER V3 ; 
        RECT 34.148 340.94 34.22 341.036 ; 
    END 
  END dataout[71] 
  PIN wd[71] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 340.556 34.66 340.652 ; 
      LAYER M3 ; 
        RECT 33.248 340.308 33.32 341.928 ; 
      LAYER V3 ; 
        RECT 33.248 340.556 33.32 340.652 ; 
    END 
  END wd[71] 
  PIN dataout[72] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 345.26 34.388 345.356 ; 
      LAYER M3 ; 
        RECT 34.148 345.058 34.22 346.016 ; 
      LAYER V3 ; 
        RECT 34.148 345.26 34.22 345.356 ; 
    END 
  END dataout[72] 
  PIN wd[72] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 344.876 34.66 344.972 ; 
      LAYER M3 ; 
        RECT 33.248 344.628 33.32 346.248 ; 
      LAYER V3 ; 
        RECT 33.248 344.876 33.32 344.972 ; 
    END 
  END wd[72] 
  PIN dataout[73] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 349.58 34.388 349.676 ; 
      LAYER M3 ; 
        RECT 34.148 349.378 34.22 350.336 ; 
      LAYER V3 ; 
        RECT 34.148 349.58 34.22 349.676 ; 
    END 
  END dataout[73] 
  PIN wd[73] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 349.196 34.66 349.292 ; 
      LAYER M3 ; 
        RECT 33.248 348.948 33.32 350.568 ; 
      LAYER V3 ; 
        RECT 33.248 349.196 33.32 349.292 ; 
    END 
  END wd[73] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0.02 104.706 66.116 109.08 ; 
      RECT 0.02 109.026 66.116 113.4 ; 
      RECT 0.02 113.346 66.116 117.72 ; 
      RECT 0.02 117.666 66.116 122.04 ; 
      RECT 0.02 121.986 66.116 126.36 ; 
      RECT 0.02 126.306 66.116 130.68 ; 
      RECT 0.02 130.626 66.116 135 ; 
      RECT 0.02 134.946 66.116 139.32 ; 
      RECT 0.02 139.266 66.116 143.64 ; 
      RECT 0.02 143.586 66.116 147.96 ; 
      RECT 0.02 147.906 66.116 152.28 ; 
      RECT 0.02 152.226 66.116 156.6 ; 
      RECT 0.02 156.546 66.116 160.92 ; 
      RECT 0 160.788 66.096 195.402 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
        RECT 0.02 240.894 66.116 245.268 ; 
        RECT 0.02 245.214 66.116 249.588 ; 
        RECT 0.02 249.534 66.116 253.908 ; 
        RECT 0.02 253.854 66.116 258.228 ; 
        RECT 0.02 258.174 66.116 262.548 ; 
        RECT 0.02 262.494 66.116 266.868 ; 
        RECT 0.02 266.814 66.116 271.188 ; 
        RECT 0.02 271.134 66.116 275.508 ; 
        RECT 0.02 275.454 66.116 279.828 ; 
        RECT 0.02 279.774 66.116 284.148 ; 
        RECT 0.02 284.094 66.116 288.468 ; 
        RECT 0.02 288.414 66.116 292.788 ; 
        RECT 0.02 292.734 66.116 297.108 ; 
        RECT 0.02 297.054 66.116 301.428 ; 
        RECT 0.02 301.374 66.116 305.748 ; 
        RECT 0.02 305.694 66.116 310.068 ; 
        RECT 0.02 310.014 66.116 314.388 ; 
        RECT 0.02 314.334 66.116 318.708 ; 
        RECT 0.02 318.654 66.116 323.028 ; 
        RECT 0.02 322.974 66.116 327.348 ; 
        RECT 0.02 327.294 66.116 331.668 ; 
        RECT 0.02 331.614 66.116 335.988 ; 
        RECT 0.02 335.934 66.116 340.308 ; 
        RECT 0.02 340.254 66.116 344.628 ; 
        RECT 0.02 344.574 66.116 348.948 ; 
        RECT 0.02 348.894 66.116 353.268 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0.02 104.706 66.116 109.08 ; 
      RECT 0.02 109.026 66.116 113.4 ; 
      RECT 0.02 113.346 66.116 117.72 ; 
      RECT 0.02 117.666 66.116 122.04 ; 
      RECT 0.02 121.986 66.116 126.36 ; 
      RECT 0.02 126.306 66.116 130.68 ; 
      RECT 0.02 130.626 66.116 135 ; 
      RECT 0.02 134.946 66.116 139.32 ; 
      RECT 0.02 139.266 66.116 143.64 ; 
      RECT 0.02 143.586 66.116 147.96 ; 
      RECT 0.02 147.906 66.116 152.28 ; 
      RECT 0.02 152.226 66.116 156.6 ; 
      RECT 0.02 156.546 66.116 160.92 ; 
      RECT 0 160.788 66.096 195.402 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
        RECT 0.02 240.894 66.116 245.268 ; 
        RECT 0.02 245.214 66.116 249.588 ; 
        RECT 0.02 249.534 66.116 253.908 ; 
        RECT 0.02 253.854 66.116 258.228 ; 
        RECT 0.02 258.174 66.116 262.548 ; 
        RECT 0.02 262.494 66.116 266.868 ; 
        RECT 0.02 266.814 66.116 271.188 ; 
        RECT 0.02 271.134 66.116 275.508 ; 
        RECT 0.02 275.454 66.116 279.828 ; 
        RECT 0.02 279.774 66.116 284.148 ; 
        RECT 0.02 284.094 66.116 288.468 ; 
        RECT 0.02 288.414 66.116 292.788 ; 
        RECT 0.02 292.734 66.116 297.108 ; 
        RECT 0.02 297.054 66.116 301.428 ; 
        RECT 0.02 301.374 66.116 305.748 ; 
        RECT 0.02 305.694 66.116 310.068 ; 
        RECT 0.02 310.014 66.116 314.388 ; 
        RECT 0.02 314.334 66.116 318.708 ; 
        RECT 0.02 318.654 66.116 323.028 ; 
        RECT 0.02 322.974 66.116 327.348 ; 
        RECT 0.02 327.294 66.116 331.668 ; 
        RECT 0.02 331.614 66.116 335.988 ; 
        RECT 0.02 335.934 66.116 340.308 ; 
        RECT 0.02 340.254 66.116 344.628 ; 
        RECT 0.02 344.574 66.116 348.948 ; 
        RECT 0.02 348.894 66.116 353.268 ; 
  LAYER V1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0.02 104.706 66.116 109.08 ; 
      RECT 0.02 109.026 66.116 113.4 ; 
      RECT 0.02 113.346 66.116 117.72 ; 
      RECT 0.02 117.666 66.116 122.04 ; 
      RECT 0.02 121.986 66.116 126.36 ; 
      RECT 0.02 126.306 66.116 130.68 ; 
      RECT 0.02 130.626 66.116 135 ; 
      RECT 0.02 134.946 66.116 139.32 ; 
      RECT 0.02 139.266 66.116 143.64 ; 
      RECT 0.02 143.586 66.116 147.96 ; 
      RECT 0.02 147.906 66.116 152.28 ; 
      RECT 0.02 152.226 66.116 156.6 ; 
      RECT 0.02 156.546 66.116 160.92 ; 
      RECT 0 160.788 66.096 195.402 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
        RECT 0.02 240.894 66.116 245.268 ; 
        RECT 0.02 245.214 66.116 249.588 ; 
        RECT 0.02 249.534 66.116 253.908 ; 
        RECT 0.02 253.854 66.116 258.228 ; 
        RECT 0.02 258.174 66.116 262.548 ; 
        RECT 0.02 262.494 66.116 266.868 ; 
        RECT 0.02 266.814 66.116 271.188 ; 
        RECT 0.02 271.134 66.116 275.508 ; 
        RECT 0.02 275.454 66.116 279.828 ; 
        RECT 0.02 279.774 66.116 284.148 ; 
        RECT 0.02 284.094 66.116 288.468 ; 
        RECT 0.02 288.414 66.116 292.788 ; 
        RECT 0.02 292.734 66.116 297.108 ; 
        RECT 0.02 297.054 66.116 301.428 ; 
        RECT 0.02 301.374 66.116 305.748 ; 
        RECT 0.02 305.694 66.116 310.068 ; 
        RECT 0.02 310.014 66.116 314.388 ; 
        RECT 0.02 314.334 66.116 318.708 ; 
        RECT 0.02 318.654 66.116 323.028 ; 
        RECT 0.02 322.974 66.116 327.348 ; 
        RECT 0.02 327.294 66.116 331.668 ; 
        RECT 0.02 331.614 66.116 335.988 ; 
        RECT 0.02 335.934 66.116 340.308 ; 
        RECT 0.02 340.254 66.116 344.628 ; 
        RECT 0.02 344.574 66.116 348.948 ; 
        RECT 0.02 348.894 66.116 353.268 ; 
  LAYER V2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0.02 104.706 66.116 109.08 ; 
      RECT 0.02 109.026 66.116 113.4 ; 
      RECT 0.02 113.346 66.116 117.72 ; 
      RECT 0.02 117.666 66.116 122.04 ; 
      RECT 0.02 121.986 66.116 126.36 ; 
      RECT 0.02 126.306 66.116 130.68 ; 
      RECT 0.02 130.626 66.116 135 ; 
      RECT 0.02 134.946 66.116 139.32 ; 
      RECT 0.02 139.266 66.116 143.64 ; 
      RECT 0.02 143.586 66.116 147.96 ; 
      RECT 0.02 147.906 66.116 152.28 ; 
      RECT 0.02 152.226 66.116 156.6 ; 
      RECT 0.02 156.546 66.116 160.92 ; 
      RECT 0 160.788 66.096 195.402 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
        RECT 0.02 240.894 66.116 245.268 ; 
        RECT 0.02 245.214 66.116 249.588 ; 
        RECT 0.02 249.534 66.116 253.908 ; 
        RECT 0.02 253.854 66.116 258.228 ; 
        RECT 0.02 258.174 66.116 262.548 ; 
        RECT 0.02 262.494 66.116 266.868 ; 
        RECT 0.02 266.814 66.116 271.188 ; 
        RECT 0.02 271.134 66.116 275.508 ; 
        RECT 0.02 275.454 66.116 279.828 ; 
        RECT 0.02 279.774 66.116 284.148 ; 
        RECT 0.02 284.094 66.116 288.468 ; 
        RECT 0.02 288.414 66.116 292.788 ; 
        RECT 0.02 292.734 66.116 297.108 ; 
        RECT 0.02 297.054 66.116 301.428 ; 
        RECT 0.02 301.374 66.116 305.748 ; 
        RECT 0.02 305.694 66.116 310.068 ; 
        RECT 0.02 310.014 66.116 314.388 ; 
        RECT 0.02 314.334 66.116 318.708 ; 
        RECT 0.02 318.654 66.116 323.028 ; 
        RECT 0.02 322.974 66.116 327.348 ; 
        RECT 0.02 327.294 66.116 331.668 ; 
        RECT 0.02 331.614 66.116 335.988 ; 
        RECT 0.02 335.934 66.116 340.308 ; 
        RECT 0.02 340.254 66.116 344.628 ; 
        RECT 0.02 344.574 66.116 348.948 ; 
        RECT 0.02 348.894 66.116 353.268 ; 
  LAYER M3 ; 
      RECT 34.796 1.38 34.868 5.122 ; 
      RECT 34.652 1.38 34.724 5.122 ; 
      RECT 34.508 3.688 34.58 4.978 ; 
      RECT 34.04 4.476 34.112 4.914 ; 
      RECT 34.004 1.51 34.076 2.468 ; 
      RECT 33.86 3.834 33.932 4.448 ; 
      RECT 33.536 3.936 33.608 4.968 ; 
      RECT 31.376 1.38 31.448 5.122 ; 
      RECT 31.232 1.38 31.304 5.122 ; 
      RECT 31.088 2.104 31.16 4.376 ; 
      RECT 34.796 5.7 34.868 9.442 ; 
      RECT 34.652 5.7 34.724 9.442 ; 
      RECT 34.508 8.008 34.58 9.298 ; 
      RECT 34.04 8.796 34.112 9.234 ; 
      RECT 34.004 5.83 34.076 6.788 ; 
      RECT 33.86 8.154 33.932 8.768 ; 
      RECT 33.536 8.256 33.608 9.288 ; 
      RECT 31.376 5.7 31.448 9.442 ; 
      RECT 31.232 5.7 31.304 9.442 ; 
      RECT 31.088 6.424 31.16 8.696 ; 
      RECT 34.796 10.02 34.868 13.762 ; 
      RECT 34.652 10.02 34.724 13.762 ; 
      RECT 34.508 12.328 34.58 13.618 ; 
      RECT 34.04 13.116 34.112 13.554 ; 
      RECT 34.004 10.15 34.076 11.108 ; 
      RECT 33.86 12.474 33.932 13.088 ; 
      RECT 33.536 12.576 33.608 13.608 ; 
      RECT 31.376 10.02 31.448 13.762 ; 
      RECT 31.232 10.02 31.304 13.762 ; 
      RECT 31.088 10.744 31.16 13.016 ; 
      RECT 34.796 14.34 34.868 18.082 ; 
      RECT 34.652 14.34 34.724 18.082 ; 
      RECT 34.508 16.648 34.58 17.938 ; 
      RECT 34.04 17.436 34.112 17.874 ; 
      RECT 34.004 14.47 34.076 15.428 ; 
      RECT 33.86 16.794 33.932 17.408 ; 
      RECT 33.536 16.896 33.608 17.928 ; 
      RECT 31.376 14.34 31.448 18.082 ; 
      RECT 31.232 14.34 31.304 18.082 ; 
      RECT 31.088 15.064 31.16 17.336 ; 
      RECT 34.796 18.66 34.868 22.402 ; 
      RECT 34.652 18.66 34.724 22.402 ; 
      RECT 34.508 20.968 34.58 22.258 ; 
      RECT 34.04 21.756 34.112 22.194 ; 
      RECT 34.004 18.79 34.076 19.748 ; 
      RECT 33.86 21.114 33.932 21.728 ; 
      RECT 33.536 21.216 33.608 22.248 ; 
      RECT 31.376 18.66 31.448 22.402 ; 
      RECT 31.232 18.66 31.304 22.402 ; 
      RECT 31.088 19.384 31.16 21.656 ; 
      RECT 34.796 22.98 34.868 26.722 ; 
      RECT 34.652 22.98 34.724 26.722 ; 
      RECT 34.508 25.288 34.58 26.578 ; 
      RECT 34.04 26.076 34.112 26.514 ; 
      RECT 34.004 23.11 34.076 24.068 ; 
      RECT 33.86 25.434 33.932 26.048 ; 
      RECT 33.536 25.536 33.608 26.568 ; 
      RECT 31.376 22.98 31.448 26.722 ; 
      RECT 31.232 22.98 31.304 26.722 ; 
      RECT 31.088 23.704 31.16 25.976 ; 
      RECT 34.796 27.3 34.868 31.042 ; 
      RECT 34.652 27.3 34.724 31.042 ; 
      RECT 34.508 29.608 34.58 30.898 ; 
      RECT 34.04 30.396 34.112 30.834 ; 
      RECT 34.004 27.43 34.076 28.388 ; 
      RECT 33.86 29.754 33.932 30.368 ; 
      RECT 33.536 29.856 33.608 30.888 ; 
      RECT 31.376 27.3 31.448 31.042 ; 
      RECT 31.232 27.3 31.304 31.042 ; 
      RECT 31.088 28.024 31.16 30.296 ; 
      RECT 34.796 31.62 34.868 35.362 ; 
      RECT 34.652 31.62 34.724 35.362 ; 
      RECT 34.508 33.928 34.58 35.218 ; 
      RECT 34.04 34.716 34.112 35.154 ; 
      RECT 34.004 31.75 34.076 32.708 ; 
      RECT 33.86 34.074 33.932 34.688 ; 
      RECT 33.536 34.176 33.608 35.208 ; 
      RECT 31.376 31.62 31.448 35.362 ; 
      RECT 31.232 31.62 31.304 35.362 ; 
      RECT 31.088 32.344 31.16 34.616 ; 
      RECT 34.796 35.94 34.868 39.682 ; 
      RECT 34.652 35.94 34.724 39.682 ; 
      RECT 34.508 38.248 34.58 39.538 ; 
      RECT 34.04 39.036 34.112 39.474 ; 
      RECT 34.004 36.07 34.076 37.028 ; 
      RECT 33.86 38.394 33.932 39.008 ; 
      RECT 33.536 38.496 33.608 39.528 ; 
      RECT 31.376 35.94 31.448 39.682 ; 
      RECT 31.232 35.94 31.304 39.682 ; 
      RECT 31.088 36.664 31.16 38.936 ; 
      RECT 34.796 40.26 34.868 44.002 ; 
      RECT 34.652 40.26 34.724 44.002 ; 
      RECT 34.508 42.568 34.58 43.858 ; 
      RECT 34.04 43.356 34.112 43.794 ; 
      RECT 34.004 40.39 34.076 41.348 ; 
      RECT 33.86 42.714 33.932 43.328 ; 
      RECT 33.536 42.816 33.608 43.848 ; 
      RECT 31.376 40.26 31.448 44.002 ; 
      RECT 31.232 40.26 31.304 44.002 ; 
      RECT 31.088 40.984 31.16 43.256 ; 
      RECT 34.796 44.58 34.868 48.322 ; 
      RECT 34.652 44.58 34.724 48.322 ; 
      RECT 34.508 46.888 34.58 48.178 ; 
      RECT 34.04 47.676 34.112 48.114 ; 
      RECT 34.004 44.71 34.076 45.668 ; 
      RECT 33.86 47.034 33.932 47.648 ; 
      RECT 33.536 47.136 33.608 48.168 ; 
      RECT 31.376 44.58 31.448 48.322 ; 
      RECT 31.232 44.58 31.304 48.322 ; 
      RECT 31.088 45.304 31.16 47.576 ; 
      RECT 34.796 48.9 34.868 52.642 ; 
      RECT 34.652 48.9 34.724 52.642 ; 
      RECT 34.508 51.208 34.58 52.498 ; 
      RECT 34.04 51.996 34.112 52.434 ; 
      RECT 34.004 49.03 34.076 49.988 ; 
      RECT 33.86 51.354 33.932 51.968 ; 
      RECT 33.536 51.456 33.608 52.488 ; 
      RECT 31.376 48.9 31.448 52.642 ; 
      RECT 31.232 48.9 31.304 52.642 ; 
      RECT 31.088 49.624 31.16 51.896 ; 
      RECT 34.796 53.22 34.868 56.962 ; 
      RECT 34.652 53.22 34.724 56.962 ; 
      RECT 34.508 55.528 34.58 56.818 ; 
      RECT 34.04 56.316 34.112 56.754 ; 
      RECT 34.004 53.35 34.076 54.308 ; 
      RECT 33.86 55.674 33.932 56.288 ; 
      RECT 33.536 55.776 33.608 56.808 ; 
      RECT 31.376 53.22 31.448 56.962 ; 
      RECT 31.232 53.22 31.304 56.962 ; 
      RECT 31.088 53.944 31.16 56.216 ; 
      RECT 34.796 57.54 34.868 61.282 ; 
      RECT 34.652 57.54 34.724 61.282 ; 
      RECT 34.508 59.848 34.58 61.138 ; 
      RECT 34.04 60.636 34.112 61.074 ; 
      RECT 34.004 57.67 34.076 58.628 ; 
      RECT 33.86 59.994 33.932 60.608 ; 
      RECT 33.536 60.096 33.608 61.128 ; 
      RECT 31.376 57.54 31.448 61.282 ; 
      RECT 31.232 57.54 31.304 61.282 ; 
      RECT 31.088 58.264 31.16 60.536 ; 
      RECT 34.796 61.86 34.868 65.602 ; 
      RECT 34.652 61.86 34.724 65.602 ; 
      RECT 34.508 64.168 34.58 65.458 ; 
      RECT 34.04 64.956 34.112 65.394 ; 
      RECT 34.004 61.99 34.076 62.948 ; 
      RECT 33.86 64.314 33.932 64.928 ; 
      RECT 33.536 64.416 33.608 65.448 ; 
      RECT 31.376 61.86 31.448 65.602 ; 
      RECT 31.232 61.86 31.304 65.602 ; 
      RECT 31.088 62.584 31.16 64.856 ; 
      RECT 34.796 66.18 34.868 69.922 ; 
      RECT 34.652 66.18 34.724 69.922 ; 
      RECT 34.508 68.488 34.58 69.778 ; 
      RECT 34.04 69.276 34.112 69.714 ; 
      RECT 34.004 66.31 34.076 67.268 ; 
      RECT 33.86 68.634 33.932 69.248 ; 
      RECT 33.536 68.736 33.608 69.768 ; 
      RECT 31.376 66.18 31.448 69.922 ; 
      RECT 31.232 66.18 31.304 69.922 ; 
      RECT 31.088 66.904 31.16 69.176 ; 
      RECT 34.796 70.5 34.868 74.242 ; 
      RECT 34.652 70.5 34.724 74.242 ; 
      RECT 34.508 72.808 34.58 74.098 ; 
      RECT 34.04 73.596 34.112 74.034 ; 
      RECT 34.004 70.63 34.076 71.588 ; 
      RECT 33.86 72.954 33.932 73.568 ; 
      RECT 33.536 73.056 33.608 74.088 ; 
      RECT 31.376 70.5 31.448 74.242 ; 
      RECT 31.232 70.5 31.304 74.242 ; 
      RECT 31.088 71.224 31.16 73.496 ; 
      RECT 34.796 74.82 34.868 78.562 ; 
      RECT 34.652 74.82 34.724 78.562 ; 
      RECT 34.508 77.128 34.58 78.418 ; 
      RECT 34.04 77.916 34.112 78.354 ; 
      RECT 34.004 74.95 34.076 75.908 ; 
      RECT 33.86 77.274 33.932 77.888 ; 
      RECT 33.536 77.376 33.608 78.408 ; 
      RECT 31.376 74.82 31.448 78.562 ; 
      RECT 31.232 74.82 31.304 78.562 ; 
      RECT 31.088 75.544 31.16 77.816 ; 
      RECT 34.796 79.14 34.868 82.882 ; 
      RECT 34.652 79.14 34.724 82.882 ; 
      RECT 34.508 81.448 34.58 82.738 ; 
      RECT 34.04 82.236 34.112 82.674 ; 
      RECT 34.004 79.27 34.076 80.228 ; 
      RECT 33.86 81.594 33.932 82.208 ; 
      RECT 33.536 81.696 33.608 82.728 ; 
      RECT 31.376 79.14 31.448 82.882 ; 
      RECT 31.232 79.14 31.304 82.882 ; 
      RECT 31.088 79.864 31.16 82.136 ; 
      RECT 34.796 83.46 34.868 87.202 ; 
      RECT 34.652 83.46 34.724 87.202 ; 
      RECT 34.508 85.768 34.58 87.058 ; 
      RECT 34.04 86.556 34.112 86.994 ; 
      RECT 34.004 83.59 34.076 84.548 ; 
      RECT 33.86 85.914 33.932 86.528 ; 
      RECT 33.536 86.016 33.608 87.048 ; 
      RECT 31.376 83.46 31.448 87.202 ; 
      RECT 31.232 83.46 31.304 87.202 ; 
      RECT 31.088 84.184 31.16 86.456 ; 
      RECT 34.796 87.78 34.868 91.522 ; 
      RECT 34.652 87.78 34.724 91.522 ; 
      RECT 34.508 90.088 34.58 91.378 ; 
      RECT 34.04 90.876 34.112 91.314 ; 
      RECT 34.004 87.91 34.076 88.868 ; 
      RECT 33.86 90.234 33.932 90.848 ; 
      RECT 33.536 90.336 33.608 91.368 ; 
      RECT 31.376 87.78 31.448 91.522 ; 
      RECT 31.232 87.78 31.304 91.522 ; 
      RECT 31.088 88.504 31.16 90.776 ; 
      RECT 34.796 92.1 34.868 95.842 ; 
      RECT 34.652 92.1 34.724 95.842 ; 
      RECT 34.508 94.408 34.58 95.698 ; 
      RECT 34.04 95.196 34.112 95.634 ; 
      RECT 34.004 92.23 34.076 93.188 ; 
      RECT 33.86 94.554 33.932 95.168 ; 
      RECT 33.536 94.656 33.608 95.688 ; 
      RECT 31.376 92.1 31.448 95.842 ; 
      RECT 31.232 92.1 31.304 95.842 ; 
      RECT 31.088 92.824 31.16 95.096 ; 
      RECT 34.796 96.42 34.868 100.162 ; 
      RECT 34.652 96.42 34.724 100.162 ; 
      RECT 34.508 98.728 34.58 100.018 ; 
      RECT 34.04 99.516 34.112 99.954 ; 
      RECT 34.004 96.55 34.076 97.508 ; 
      RECT 33.86 98.874 33.932 99.488 ; 
      RECT 33.536 98.976 33.608 100.008 ; 
      RECT 31.376 96.42 31.448 100.162 ; 
      RECT 31.232 96.42 31.304 100.162 ; 
      RECT 31.088 97.144 31.16 99.416 ; 
      RECT 34.796 100.74 34.868 104.482 ; 
      RECT 34.652 100.74 34.724 104.482 ; 
      RECT 34.508 103.048 34.58 104.338 ; 
      RECT 34.04 103.836 34.112 104.274 ; 
      RECT 34.004 100.87 34.076 101.828 ; 
      RECT 33.86 103.194 33.932 103.808 ; 
      RECT 33.536 103.296 33.608 104.328 ; 
      RECT 31.376 100.74 31.448 104.482 ; 
      RECT 31.232 100.74 31.304 104.482 ; 
      RECT 31.088 101.464 31.16 103.736 ; 
      RECT 34.796 105.06 34.868 108.802 ; 
      RECT 34.652 105.06 34.724 108.802 ; 
      RECT 34.508 107.368 34.58 108.658 ; 
      RECT 34.04 108.156 34.112 108.594 ; 
      RECT 34.004 105.19 34.076 106.148 ; 
      RECT 33.86 107.514 33.932 108.128 ; 
      RECT 33.536 107.616 33.608 108.648 ; 
      RECT 31.376 105.06 31.448 108.802 ; 
      RECT 31.232 105.06 31.304 108.802 ; 
      RECT 31.088 105.784 31.16 108.056 ; 
      RECT 34.796 109.38 34.868 113.122 ; 
      RECT 34.652 109.38 34.724 113.122 ; 
      RECT 34.508 111.688 34.58 112.978 ; 
      RECT 34.04 112.476 34.112 112.914 ; 
      RECT 34.004 109.51 34.076 110.468 ; 
      RECT 33.86 111.834 33.932 112.448 ; 
      RECT 33.536 111.936 33.608 112.968 ; 
      RECT 31.376 109.38 31.448 113.122 ; 
      RECT 31.232 109.38 31.304 113.122 ; 
      RECT 31.088 110.104 31.16 112.376 ; 
      RECT 34.796 113.7 34.868 117.442 ; 
      RECT 34.652 113.7 34.724 117.442 ; 
      RECT 34.508 116.008 34.58 117.298 ; 
      RECT 34.04 116.796 34.112 117.234 ; 
      RECT 34.004 113.83 34.076 114.788 ; 
      RECT 33.86 116.154 33.932 116.768 ; 
      RECT 33.536 116.256 33.608 117.288 ; 
      RECT 31.376 113.7 31.448 117.442 ; 
      RECT 31.232 113.7 31.304 117.442 ; 
      RECT 31.088 114.424 31.16 116.696 ; 
      RECT 34.796 118.02 34.868 121.762 ; 
      RECT 34.652 118.02 34.724 121.762 ; 
      RECT 34.508 120.328 34.58 121.618 ; 
      RECT 34.04 121.116 34.112 121.554 ; 
      RECT 34.004 118.15 34.076 119.108 ; 
      RECT 33.86 120.474 33.932 121.088 ; 
      RECT 33.536 120.576 33.608 121.608 ; 
      RECT 31.376 118.02 31.448 121.762 ; 
      RECT 31.232 118.02 31.304 121.762 ; 
      RECT 31.088 118.744 31.16 121.016 ; 
      RECT 34.796 122.34 34.868 126.082 ; 
      RECT 34.652 122.34 34.724 126.082 ; 
      RECT 34.508 124.648 34.58 125.938 ; 
      RECT 34.04 125.436 34.112 125.874 ; 
      RECT 34.004 122.47 34.076 123.428 ; 
      RECT 33.86 124.794 33.932 125.408 ; 
      RECT 33.536 124.896 33.608 125.928 ; 
      RECT 31.376 122.34 31.448 126.082 ; 
      RECT 31.232 122.34 31.304 126.082 ; 
      RECT 31.088 123.064 31.16 125.336 ; 
      RECT 34.796 126.66 34.868 130.402 ; 
      RECT 34.652 126.66 34.724 130.402 ; 
      RECT 34.508 128.968 34.58 130.258 ; 
      RECT 34.04 129.756 34.112 130.194 ; 
      RECT 34.004 126.79 34.076 127.748 ; 
      RECT 33.86 129.114 33.932 129.728 ; 
      RECT 33.536 129.216 33.608 130.248 ; 
      RECT 31.376 126.66 31.448 130.402 ; 
      RECT 31.232 126.66 31.304 130.402 ; 
      RECT 31.088 127.384 31.16 129.656 ; 
      RECT 34.796 130.98 34.868 134.722 ; 
      RECT 34.652 130.98 34.724 134.722 ; 
      RECT 34.508 133.288 34.58 134.578 ; 
      RECT 34.04 134.076 34.112 134.514 ; 
      RECT 34.004 131.11 34.076 132.068 ; 
      RECT 33.86 133.434 33.932 134.048 ; 
      RECT 33.536 133.536 33.608 134.568 ; 
      RECT 31.376 130.98 31.448 134.722 ; 
      RECT 31.232 130.98 31.304 134.722 ; 
      RECT 31.088 131.704 31.16 133.976 ; 
      RECT 34.796 135.3 34.868 139.042 ; 
      RECT 34.652 135.3 34.724 139.042 ; 
      RECT 34.508 137.608 34.58 138.898 ; 
      RECT 34.04 138.396 34.112 138.834 ; 
      RECT 34.004 135.43 34.076 136.388 ; 
      RECT 33.86 137.754 33.932 138.368 ; 
      RECT 33.536 137.856 33.608 138.888 ; 
      RECT 31.376 135.3 31.448 139.042 ; 
      RECT 31.232 135.3 31.304 139.042 ; 
      RECT 31.088 136.024 31.16 138.296 ; 
      RECT 34.796 139.62 34.868 143.362 ; 
      RECT 34.652 139.62 34.724 143.362 ; 
      RECT 34.508 141.928 34.58 143.218 ; 
      RECT 34.04 142.716 34.112 143.154 ; 
      RECT 34.004 139.75 34.076 140.708 ; 
      RECT 33.86 142.074 33.932 142.688 ; 
      RECT 33.536 142.176 33.608 143.208 ; 
      RECT 31.376 139.62 31.448 143.362 ; 
      RECT 31.232 139.62 31.304 143.362 ; 
      RECT 31.088 140.344 31.16 142.616 ; 
      RECT 34.796 143.94 34.868 147.682 ; 
      RECT 34.652 143.94 34.724 147.682 ; 
      RECT 34.508 146.248 34.58 147.538 ; 
      RECT 34.04 147.036 34.112 147.474 ; 
      RECT 34.004 144.07 34.076 145.028 ; 
      RECT 33.86 146.394 33.932 147.008 ; 
      RECT 33.536 146.496 33.608 147.528 ; 
      RECT 31.376 143.94 31.448 147.682 ; 
      RECT 31.232 143.94 31.304 147.682 ; 
      RECT 31.088 144.664 31.16 146.936 ; 
      RECT 34.796 148.26 34.868 152.002 ; 
      RECT 34.652 148.26 34.724 152.002 ; 
      RECT 34.508 150.568 34.58 151.858 ; 
      RECT 34.04 151.356 34.112 151.794 ; 
      RECT 34.004 148.39 34.076 149.348 ; 
      RECT 33.86 150.714 33.932 151.328 ; 
      RECT 33.536 150.816 33.608 151.848 ; 
      RECT 31.376 148.26 31.448 152.002 ; 
      RECT 31.232 148.26 31.304 152.002 ; 
      RECT 31.088 148.984 31.16 151.256 ; 
      RECT 34.796 152.58 34.868 156.322 ; 
      RECT 34.652 152.58 34.724 156.322 ; 
      RECT 34.508 154.888 34.58 156.178 ; 
      RECT 34.04 155.676 34.112 156.114 ; 
      RECT 34.004 152.71 34.076 153.668 ; 
      RECT 33.86 155.034 33.932 155.648 ; 
      RECT 33.536 155.136 33.608 156.168 ; 
      RECT 31.376 152.58 31.448 156.322 ; 
      RECT 31.232 152.58 31.304 156.322 ; 
      RECT 31.088 153.304 31.16 155.576 ; 
      RECT 34.796 156.9 34.868 160.642 ; 
      RECT 34.652 156.9 34.724 160.642 ; 
      RECT 34.508 159.208 34.58 160.498 ; 
      RECT 34.04 159.996 34.112 160.434 ; 
      RECT 34.004 157.03 34.076 157.988 ; 
      RECT 33.86 159.354 33.932 159.968 ; 
      RECT 33.536 159.456 33.608 160.488 ; 
      RECT 31.376 156.9 31.448 160.642 ; 
      RECT 31.232 156.9 31.304 160.642 ; 
      RECT 31.088 157.624 31.16 159.896 ; 
      RECT 65.268 175.96 65.34 193.376 ; 
      RECT 65.124 170.7 65.196 170.976 ; 
      RECT 65.124 177.18 65.196 177.512 ; 
      RECT 64.98 160.682 65.052 193.51 ; 
      RECT 64.836 176.09 64.908 178.85 ; 
      RECT 64.836 179.054 64.908 183 ; 
      RECT 64.836 183.16 64.908 185.628 ; 
      RECT 64.692 175.836 64.764 178.6548 ; 
      RECT 64.692 181.668 64.764 186.348 ; 
      RECT 64.548 160.682 64.62 175.068 ; 
      RECT 64.116 160.682 64.188 175.068 ; 
      RECT 63.684 160.682 63.756 175.068 ; 
      RECT 63.252 160.682 63.324 175.068 ; 
      RECT 62.82 160.682 62.892 175.068 ; 
      RECT 62.388 160.682 62.46 175.068 ; 
      RECT 61.956 160.682 62.028 175.068 ; 
      RECT 61.524 160.682 61.596 175.068 ; 
      RECT 61.092 160.682 61.164 175.068 ; 
      RECT 60.66 160.682 60.732 175.068 ; 
      RECT 60.228 160.682 60.3 175.068 ; 
      RECT 59.796 160.682 59.868 175.068 ; 
      RECT 59.364 160.682 59.436 175.068 ; 
      RECT 58.932 160.682 59.004 175.068 ; 
      RECT 58.5 160.682 58.572 175.068 ; 
      RECT 58.068 160.682 58.14 175.068 ; 
      RECT 57.636 160.682 57.708 175.068 ; 
      RECT 57.204 160.682 57.276 175.068 ; 
      RECT 56.772 160.682 56.844 175.068 ; 
      RECT 56.34 160.682 56.412 175.068 ; 
      RECT 55.908 160.682 55.98 175.068 ; 
      RECT 55.476 160.682 55.548 175.068 ; 
      RECT 55.044 160.682 55.116 175.068 ; 
      RECT 54.612 160.682 54.684 175.068 ; 
      RECT 54.18 160.682 54.252 175.068 ; 
      RECT 53.748 160.682 53.82 175.068 ; 
      RECT 53.316 160.682 53.388 175.068 ; 
      RECT 52.884 160.682 52.956 175.068 ; 
      RECT 52.452 160.682 52.524 175.068 ; 
      RECT 52.02 160.682 52.092 175.068 ; 
      RECT 51.588 160.682 51.66 175.068 ; 
      RECT 51.156 160.682 51.228 175.068 ; 
      RECT 50.724 160.682 50.796 175.068 ; 
      RECT 50.292 160.682 50.364 175.068 ; 
      RECT 49.86 160.682 49.932 175.068 ; 
      RECT 49.428 160.682 49.5 175.068 ; 
      RECT 48.996 160.682 49.068 175.068 ; 
      RECT 48.564 160.682 48.636 175.068 ; 
      RECT 48.132 160.682 48.204 175.068 ; 
      RECT 47.7 160.682 47.772 175.068 ; 
      RECT 47.268 160.682 47.34 175.068 ; 
      RECT 46.836 160.682 46.908 175.068 ; 
      RECT 46.404 160.682 46.476 175.068 ; 
      RECT 45.972 160.682 46.044 175.068 ; 
      RECT 45.54 160.682 45.612 175.068 ; 
      RECT 45.108 160.682 45.18 175.068 ; 
      RECT 44.676 160.682 44.748 175.068 ; 
      RECT 44.244 160.682 44.316 175.068 ; 
      RECT 43.812 160.682 43.884 175.068 ; 
      RECT 43.38 160.682 43.452 175.068 ; 
      RECT 42.948 160.682 43.02 175.068 ; 
      RECT 42.516 160.682 42.588 175.068 ; 
      RECT 42.084 160.682 42.156 175.068 ; 
      RECT 41.652 160.682 41.724 175.068 ; 
      RECT 41.22 160.682 41.292 175.068 ; 
      RECT 40.788 160.682 40.86 175.068 ; 
      RECT 40.356 160.682 40.428 175.068 ; 
      RECT 39.924 160.682 39.996 175.068 ; 
      RECT 39.492 160.682 39.564 175.068 ; 
      RECT 39.06 160.682 39.132 175.068 ; 
      RECT 38.628 160.682 38.7 175.068 ; 
      RECT 38.196 160.682 38.268 175.068 ; 
      RECT 38.052 176.102 38.124 178.67 ; 
      RECT 38.052 181.38 38.124 183.508 ; 
      RECT 37.98 163.324 38.052 166.028 ; 
      RECT 37.98 169.012 38.052 170.204 ; 
      RECT 37.98 173.476 38.052 174.524 ; 
      RECT 37.908 175.76 37.98 178.85 ; 
      RECT 37.908 179.0548 37.98 181.02 ; 
      RECT 37.908 181.2 37.98 182.684 ; 
      RECT 37.908 182.988 37.98 185.628 ; 
      RECT 37.764 160.682 37.836 193.51 ; 
      RECT 37.62 177.932 37.692 179.79 ; 
      RECT 37.548 163.756 37.62 166.28 ; 
      RECT 37.548 167.932 37.62 168.692 ; 
      RECT 37.548 171.46 37.62 171.656 ; 
      RECT 37.548 174.388 37.62 174.536 ; 
      RECT 37.476 175.96 37.548 193.358 ; 
      RECT 37.116 162.244 37.188 165.452 ; 
      RECT 37.116 167.644 37.188 169.916 ; 
      RECT 36.972 167.932 37.044 169.412 ; 
      RECT 36.828 165.34 36.9 165.884 ; 
      RECT 36.828 169.3 36.9 170.204 ; 
      RECT 36.828 174.268 36.9 174.524 ; 
      RECT 36.684 165.748 36.756 165.896 ; 
      RECT 36.684 172.252 36.756 172.424 ; 
      RECT 36.684 174.388 36.756 174.536 ; 
      RECT 36.54 166.996 36.612 168.98 ; 
      RECT 36.54 169.156 36.612 169.916 ; 
      RECT 36.54 172.996 36.612 174.236 ; 
      RECT 36.396 166.564 36.468 171.552 ; 
      RECT 36.396 182.116 36.468 185.036 ; 
      RECT 36.396 186.436 36.468 189.356 ; 
      RECT 35.1 165.484 35.172 166.676 ; 
      RECT 35.1 170.236 35.172 170.492 ; 
      RECT 35.1 171.316 35.172 173.156 ; 
      RECT 35.1 176.116 35.172 176.264 ; 
      RECT 35.1 184.276 35.172 185.468 ; 
      RECT 34.956 165.772 35.028 167.792 ; 
      RECT 34.956 168.868 35.028 172.076 ; 
      RECT 34.956 176.248 35.028 177.332 ; 
      RECT 34.956 177.652 35.028 178.556 ; 
      RECT 34.812 165.484 34.884 168.188 ; 
      RECT 34.812 168.58 34.884 169.916 ; 
      RECT 34.812 170.74 34.884 171.284 ; 
      RECT 34.812 173.476 34.884 176.684 ; 
      RECT 34.812 178.42 34.884 178.568 ; 
      RECT 34.812 187.084 34.884 188.42 ; 
      RECT 34.668 166.42 34.74 166.964 ; 
      RECT 34.668 173.98 34.74 177.908 ; 
      RECT 34.668 179.668 34.74 180.86 ; 
      RECT 34.668 186.436 34.74 187.484 ; 
      RECT 34.524 162.676 34.596 163.292 ; 
      RECT 34.524 165.916 34.596 173.06 ; 
      RECT 34.524 177.22 34.596 186.548 ; 
      RECT 34.524 187.372 34.596 191.804 ; 
      RECT 33.372 163.756 33.444 164.804 ; 
      RECT 33.372 165.34 33.444 165.596 ; 
      RECT 33.372 165.916 33.444 166.82 ; 
      RECT 33.372 166.996 33.444 167.756 ; 
      RECT 33.372 168.076 33.444 178.556 ; 
      RECT 33.372 178.732 33.444 183.956 ; 
      RECT 33.372 188.308 33.444 189.356 ; 
      RECT 33.228 167.752 33.3 168.836 ; 
      RECT 33.228 169.156 33.3 172.508 ; 
      RECT 33.228 173.188 33.3 176.54 ; 
      RECT 33.228 176.716 33.3 181.796 ; 
      RECT 33.228 182.62 33.3 183.308 ; 
      RECT 33.228 186.148 33.3 190.436 ; 
      RECT 33.084 168.076 33.156 169.16 ; 
      RECT 33.084 169.78 33.156 169.928 ; 
      RECT 33.084 172.9 33.156 176.828 ; 
      RECT 33.084 177.796 33.156 179.636 ; 
      RECT 33.084 181.036 33.156 183.992 ; 
      RECT 32.94 164.548 33.012 168.836 ; 
      RECT 32.94 175.204 33.012 176.072 ; 
      RECT 32.94 180.748 33.012 181.94 ; 
      RECT 32.796 167.14 32.868 168.98 ; 
      RECT 32.796 173.476 32.868 174.236 ; 
      RECT 32.796 174.4 32.868 174.548 ; 
      RECT 32.796 175.492 32.868 176.828 ; 
      RECT 32.796 177.364 32.868 182.732 ; 
      RECT 32.796 183.16 32.868 187.628 ; 
      RECT 32.652 164.836 32.724 165.596 ; 
      RECT 32.652 166.42 32.724 166.964 ; 
      RECT 32.652 168.076 32.724 180.716 ; 
      RECT 32.652 181.036 32.724 182.876 ; 
      RECT 32.652 185.356 32.724 187.196 ; 
      RECT 32.652 190.612 32.724 191.516 ; 
      RECT 32.508 160.788 32.58 161.404 ; 
      RECT 32.508 192.768 32.58 193.432 ; 
      RECT 32.364 160.788 32.436 160.988 ; 
      RECT 32.076 160.788 32.148 161.074 ; 
      RECT 32.076 193.046 32.148 193.51 ; 
      RECT 31.5 166.852 31.572 167.612 ; 
      RECT 31.5 169.804 31.572 171.284 ; 
      RECT 31.5 177.652 31.572 178.556 ; 
      RECT 31.5 179.812 31.572 184.388 ; 
      RECT 31.5 187.516 31.572 189.356 ; 
      RECT 31.5 191.668 31.572 191.816 ; 
      RECT 31.356 162.676 31.428 164.66 ; 
      RECT 31.356 178.996 31.428 179.144 ; 
      RECT 31.356 183.304 31.428 186.548 ; 
      RECT 31.212 164.548 31.284 165.596 ; 
      RECT 31.212 166.708 31.284 168.044 ; 
      RECT 31.212 168.868 31.284 169.268 ; 
      RECT 31.212 172.396 31.284 183.452 ; 
      RECT 31.212 183.988 31.284 184.892 ; 
      RECT 31.068 163.18 31.14 167.756 ; 
      RECT 31.068 182.116 31.14 182.876 ; 
      RECT 31.068 185.332 31.14 185.48 ; 
      RECT 31.068 186.436 31.14 189.644 ; 
      RECT 30.924 166.996 30.996 170.996 ; 
      RECT 30.924 184.756 30.996 184.904 ; 
      RECT 29.484 165.34 29.556 166.964 ; 
      RECT 29.196 165.484 29.268 167.9 ; 
      RECT 29.052 164.836 29.124 165.092 ; 
      RECT 28.908 161 28.98 161.204 ; 
      RECT 28.908 173.476 28.98 174.236 ; 
      RECT 28.836 175.96 28.908 193.354 ; 
      RECT 28.548 175.96 28.62 193.358 ; 
      RECT 28.476 162.676 28.548 163.436 ; 
      RECT 28.476 165.772 28.548 174.812 ; 
      RECT 28.404 177.932 28.476 179.79 ; 
      RECT 28.26 160.682 28.332 193.51 ; 
      RECT 28.116 175.76 28.188 178.85 ; 
      RECT 28.116 179.0548 28.188 181.02 ; 
      RECT 28.116 181.2 28.188 182.684 ; 
      RECT 28.116 182.988 28.188 185.628 ; 
      RECT 28.044 162.676 28.116 164.66 ; 
      RECT 28.044 167.788 28.116 170.06 ; 
      RECT 28.044 171.316 28.116 174.236 ; 
      RECT 27.972 176.102 28.044 178.67 ; 
      RECT 27.972 181.38 28.044 183.508 ; 
      RECT 27.828 160.682 27.9 175.068 ; 
      RECT 27.396 160.682 27.468 175.068 ; 
      RECT 26.964 160.682 27.036 175.068 ; 
      RECT 26.532 160.682 26.604 175.068 ; 
      RECT 26.1 160.682 26.172 175.068 ; 
      RECT 25.668 160.682 25.74 175.068 ; 
      RECT 25.236 160.682 25.308 175.068 ; 
      RECT 24.804 160.682 24.876 175.068 ; 
      RECT 24.372 160.682 24.444 175.068 ; 
      RECT 23.94 160.682 24.012 175.068 ; 
      RECT 23.508 160.682 23.58 175.068 ; 
      RECT 23.076 160.682 23.148 175.068 ; 
      RECT 22.644 160.682 22.716 175.068 ; 
      RECT 22.212 160.682 22.284 175.068 ; 
      RECT 21.78 160.682 21.852 175.068 ; 
      RECT 21.348 160.682 21.42 175.068 ; 
      RECT 20.916 160.682 20.988 175.068 ; 
      RECT 20.484 160.682 20.556 175.068 ; 
      RECT 20.052 160.682 20.124 175.068 ; 
      RECT 19.62 160.682 19.692 175.068 ; 
      RECT 19.188 160.682 19.26 175.068 ; 
      RECT 18.756 160.682 18.828 175.068 ; 
      RECT 18.324 160.682 18.396 175.068 ; 
      RECT 17.892 160.682 17.964 175.068 ; 
      RECT 17.46 160.682 17.532 175.068 ; 
      RECT 17.028 160.682 17.1 175.068 ; 
      RECT 16.596 160.682 16.668 175.068 ; 
      RECT 16.164 160.682 16.236 175.068 ; 
      RECT 15.732 160.682 15.804 175.068 ; 
      RECT 15.3 160.682 15.372 175.068 ; 
      RECT 14.868 160.682 14.94 175.068 ; 
      RECT 14.436 160.682 14.508 175.068 ; 
      RECT 14.004 160.682 14.076 175.068 ; 
      RECT 13.572 160.682 13.644 175.068 ; 
      RECT 13.14 160.682 13.212 175.068 ; 
      RECT 12.708 160.682 12.78 175.068 ; 
      RECT 12.276 160.682 12.348 175.068 ; 
      RECT 11.844 160.682 11.916 175.068 ; 
      RECT 11.412 160.682 11.484 175.068 ; 
      RECT 10.98 160.682 11.052 175.068 ; 
      RECT 10.548 160.682 10.62 175.068 ; 
      RECT 10.116 160.682 10.188 175.068 ; 
      RECT 9.684 160.682 9.756 175.068 ; 
      RECT 9.252 160.682 9.324 175.068 ; 
      RECT 8.82 160.682 8.892 175.068 ; 
      RECT 8.388 160.682 8.46 175.068 ; 
      RECT 7.956 160.682 8.028 175.068 ; 
      RECT 7.524 160.682 7.596 175.068 ; 
      RECT 7.092 160.682 7.164 175.068 ; 
      RECT 6.66 160.682 6.732 175.068 ; 
      RECT 6.228 160.682 6.3 175.068 ; 
      RECT 5.796 160.682 5.868 175.068 ; 
      RECT 5.364 160.682 5.436 175.068 ; 
      RECT 4.932 160.682 5.004 175.068 ; 
      RECT 4.5 160.682 4.572 175.068 ; 
      RECT 4.068 160.682 4.14 175.068 ; 
      RECT 3.636 160.682 3.708 175.068 ; 
      RECT 3.204 160.682 3.276 175.068 ; 
      RECT 2.772 160.682 2.844 175.068 ; 
      RECT 2.34 160.682 2.412 175.068 ; 
      RECT 1.908 160.682 1.98 175.068 ; 
      RECT 1.476 160.682 1.548 175.068 ; 
      RECT 1.332 175.836 1.404 178.6548 ; 
      RECT 1.332 181.668 1.404 186.348 ; 
      RECT 1.188 176.09 1.26 178.85 ; 
      RECT 1.188 179.054 1.26 183 ; 
      RECT 1.188 183.16 1.26 185.628 ; 
      RECT 1.044 160.682 1.116 193.51 ; 
      RECT 0.9 170.7 0.972 170.976 ; 
      RECT 0.9 177.18 0.972 177.512 ; 
      RECT 0.756 175.96 0.828 193.376 ; 
        RECT 34.796 193.728 34.868 197.47 ; 
        RECT 34.652 193.728 34.724 197.47 ; 
        RECT 34.508 196.036 34.58 197.326 ; 
        RECT 34.04 196.824 34.112 197.262 ; 
        RECT 34.004 193.858 34.076 194.816 ; 
        RECT 33.86 196.182 33.932 196.796 ; 
        RECT 33.536 196.284 33.608 197.316 ; 
        RECT 31.376 193.728 31.448 197.47 ; 
        RECT 31.232 193.728 31.304 197.47 ; 
        RECT 31.088 194.452 31.16 196.724 ; 
        RECT 34.796 198.048 34.868 201.79 ; 
        RECT 34.652 198.048 34.724 201.79 ; 
        RECT 34.508 200.356 34.58 201.646 ; 
        RECT 34.04 201.144 34.112 201.582 ; 
        RECT 34.004 198.178 34.076 199.136 ; 
        RECT 33.86 200.502 33.932 201.116 ; 
        RECT 33.536 200.604 33.608 201.636 ; 
        RECT 31.376 198.048 31.448 201.79 ; 
        RECT 31.232 198.048 31.304 201.79 ; 
        RECT 31.088 198.772 31.16 201.044 ; 
        RECT 34.796 202.368 34.868 206.11 ; 
        RECT 34.652 202.368 34.724 206.11 ; 
        RECT 34.508 204.676 34.58 205.966 ; 
        RECT 34.04 205.464 34.112 205.902 ; 
        RECT 34.004 202.498 34.076 203.456 ; 
        RECT 33.86 204.822 33.932 205.436 ; 
        RECT 33.536 204.924 33.608 205.956 ; 
        RECT 31.376 202.368 31.448 206.11 ; 
        RECT 31.232 202.368 31.304 206.11 ; 
        RECT 31.088 203.092 31.16 205.364 ; 
        RECT 34.796 206.688 34.868 210.43 ; 
        RECT 34.652 206.688 34.724 210.43 ; 
        RECT 34.508 208.996 34.58 210.286 ; 
        RECT 34.04 209.784 34.112 210.222 ; 
        RECT 34.004 206.818 34.076 207.776 ; 
        RECT 33.86 209.142 33.932 209.756 ; 
        RECT 33.536 209.244 33.608 210.276 ; 
        RECT 31.376 206.688 31.448 210.43 ; 
        RECT 31.232 206.688 31.304 210.43 ; 
        RECT 31.088 207.412 31.16 209.684 ; 
        RECT 34.796 211.008 34.868 214.75 ; 
        RECT 34.652 211.008 34.724 214.75 ; 
        RECT 34.508 213.316 34.58 214.606 ; 
        RECT 34.04 214.104 34.112 214.542 ; 
        RECT 34.004 211.138 34.076 212.096 ; 
        RECT 33.86 213.462 33.932 214.076 ; 
        RECT 33.536 213.564 33.608 214.596 ; 
        RECT 31.376 211.008 31.448 214.75 ; 
        RECT 31.232 211.008 31.304 214.75 ; 
        RECT 31.088 211.732 31.16 214.004 ; 
        RECT 34.796 215.328 34.868 219.07 ; 
        RECT 34.652 215.328 34.724 219.07 ; 
        RECT 34.508 217.636 34.58 218.926 ; 
        RECT 34.04 218.424 34.112 218.862 ; 
        RECT 34.004 215.458 34.076 216.416 ; 
        RECT 33.86 217.782 33.932 218.396 ; 
        RECT 33.536 217.884 33.608 218.916 ; 
        RECT 31.376 215.328 31.448 219.07 ; 
        RECT 31.232 215.328 31.304 219.07 ; 
        RECT 31.088 216.052 31.16 218.324 ; 
        RECT 34.796 219.648 34.868 223.39 ; 
        RECT 34.652 219.648 34.724 223.39 ; 
        RECT 34.508 221.956 34.58 223.246 ; 
        RECT 34.04 222.744 34.112 223.182 ; 
        RECT 34.004 219.778 34.076 220.736 ; 
        RECT 33.86 222.102 33.932 222.716 ; 
        RECT 33.536 222.204 33.608 223.236 ; 
        RECT 31.376 219.648 31.448 223.39 ; 
        RECT 31.232 219.648 31.304 223.39 ; 
        RECT 31.088 220.372 31.16 222.644 ; 
        RECT 34.796 223.968 34.868 227.71 ; 
        RECT 34.652 223.968 34.724 227.71 ; 
        RECT 34.508 226.276 34.58 227.566 ; 
        RECT 34.04 227.064 34.112 227.502 ; 
        RECT 34.004 224.098 34.076 225.056 ; 
        RECT 33.86 226.422 33.932 227.036 ; 
        RECT 33.536 226.524 33.608 227.556 ; 
        RECT 31.376 223.968 31.448 227.71 ; 
        RECT 31.232 223.968 31.304 227.71 ; 
        RECT 31.088 224.692 31.16 226.964 ; 
        RECT 34.796 228.288 34.868 232.03 ; 
        RECT 34.652 228.288 34.724 232.03 ; 
        RECT 34.508 230.596 34.58 231.886 ; 
        RECT 34.04 231.384 34.112 231.822 ; 
        RECT 34.004 228.418 34.076 229.376 ; 
        RECT 33.86 230.742 33.932 231.356 ; 
        RECT 33.536 230.844 33.608 231.876 ; 
        RECT 31.376 228.288 31.448 232.03 ; 
        RECT 31.232 228.288 31.304 232.03 ; 
        RECT 31.088 229.012 31.16 231.284 ; 
        RECT 34.796 232.608 34.868 236.35 ; 
        RECT 34.652 232.608 34.724 236.35 ; 
        RECT 34.508 234.916 34.58 236.206 ; 
        RECT 34.04 235.704 34.112 236.142 ; 
        RECT 34.004 232.738 34.076 233.696 ; 
        RECT 33.86 235.062 33.932 235.676 ; 
        RECT 33.536 235.164 33.608 236.196 ; 
        RECT 31.376 232.608 31.448 236.35 ; 
        RECT 31.232 232.608 31.304 236.35 ; 
        RECT 31.088 233.332 31.16 235.604 ; 
        RECT 34.796 236.928 34.868 240.67 ; 
        RECT 34.652 236.928 34.724 240.67 ; 
        RECT 34.508 239.236 34.58 240.526 ; 
        RECT 34.04 240.024 34.112 240.462 ; 
        RECT 34.004 237.058 34.076 238.016 ; 
        RECT 33.86 239.382 33.932 239.996 ; 
        RECT 33.536 239.484 33.608 240.516 ; 
        RECT 31.376 236.928 31.448 240.67 ; 
        RECT 31.232 236.928 31.304 240.67 ; 
        RECT 31.088 237.652 31.16 239.924 ; 
        RECT 34.796 241.248 34.868 244.99 ; 
        RECT 34.652 241.248 34.724 244.99 ; 
        RECT 34.508 243.556 34.58 244.846 ; 
        RECT 34.04 244.344 34.112 244.782 ; 
        RECT 34.004 241.378 34.076 242.336 ; 
        RECT 33.86 243.702 33.932 244.316 ; 
        RECT 33.536 243.804 33.608 244.836 ; 
        RECT 31.376 241.248 31.448 244.99 ; 
        RECT 31.232 241.248 31.304 244.99 ; 
        RECT 31.088 241.972 31.16 244.244 ; 
        RECT 34.796 245.568 34.868 249.31 ; 
        RECT 34.652 245.568 34.724 249.31 ; 
        RECT 34.508 247.876 34.58 249.166 ; 
        RECT 34.04 248.664 34.112 249.102 ; 
        RECT 34.004 245.698 34.076 246.656 ; 
        RECT 33.86 248.022 33.932 248.636 ; 
        RECT 33.536 248.124 33.608 249.156 ; 
        RECT 31.376 245.568 31.448 249.31 ; 
        RECT 31.232 245.568 31.304 249.31 ; 
        RECT 31.088 246.292 31.16 248.564 ; 
        RECT 34.796 249.888 34.868 253.63 ; 
        RECT 34.652 249.888 34.724 253.63 ; 
        RECT 34.508 252.196 34.58 253.486 ; 
        RECT 34.04 252.984 34.112 253.422 ; 
        RECT 34.004 250.018 34.076 250.976 ; 
        RECT 33.86 252.342 33.932 252.956 ; 
        RECT 33.536 252.444 33.608 253.476 ; 
        RECT 31.376 249.888 31.448 253.63 ; 
        RECT 31.232 249.888 31.304 253.63 ; 
        RECT 31.088 250.612 31.16 252.884 ; 
        RECT 34.796 254.208 34.868 257.95 ; 
        RECT 34.652 254.208 34.724 257.95 ; 
        RECT 34.508 256.516 34.58 257.806 ; 
        RECT 34.04 257.304 34.112 257.742 ; 
        RECT 34.004 254.338 34.076 255.296 ; 
        RECT 33.86 256.662 33.932 257.276 ; 
        RECT 33.536 256.764 33.608 257.796 ; 
        RECT 31.376 254.208 31.448 257.95 ; 
        RECT 31.232 254.208 31.304 257.95 ; 
        RECT 31.088 254.932 31.16 257.204 ; 
        RECT 34.796 258.528 34.868 262.27 ; 
        RECT 34.652 258.528 34.724 262.27 ; 
        RECT 34.508 260.836 34.58 262.126 ; 
        RECT 34.04 261.624 34.112 262.062 ; 
        RECT 34.004 258.658 34.076 259.616 ; 
        RECT 33.86 260.982 33.932 261.596 ; 
        RECT 33.536 261.084 33.608 262.116 ; 
        RECT 31.376 258.528 31.448 262.27 ; 
        RECT 31.232 258.528 31.304 262.27 ; 
        RECT 31.088 259.252 31.16 261.524 ; 
        RECT 34.796 262.848 34.868 266.59 ; 
        RECT 34.652 262.848 34.724 266.59 ; 
        RECT 34.508 265.156 34.58 266.446 ; 
        RECT 34.04 265.944 34.112 266.382 ; 
        RECT 34.004 262.978 34.076 263.936 ; 
        RECT 33.86 265.302 33.932 265.916 ; 
        RECT 33.536 265.404 33.608 266.436 ; 
        RECT 31.376 262.848 31.448 266.59 ; 
        RECT 31.232 262.848 31.304 266.59 ; 
        RECT 31.088 263.572 31.16 265.844 ; 
        RECT 34.796 267.168 34.868 270.91 ; 
        RECT 34.652 267.168 34.724 270.91 ; 
        RECT 34.508 269.476 34.58 270.766 ; 
        RECT 34.04 270.264 34.112 270.702 ; 
        RECT 34.004 267.298 34.076 268.256 ; 
        RECT 33.86 269.622 33.932 270.236 ; 
        RECT 33.536 269.724 33.608 270.756 ; 
        RECT 31.376 267.168 31.448 270.91 ; 
        RECT 31.232 267.168 31.304 270.91 ; 
        RECT 31.088 267.892 31.16 270.164 ; 
        RECT 34.796 271.488 34.868 275.23 ; 
        RECT 34.652 271.488 34.724 275.23 ; 
        RECT 34.508 273.796 34.58 275.086 ; 
        RECT 34.04 274.584 34.112 275.022 ; 
        RECT 34.004 271.618 34.076 272.576 ; 
        RECT 33.86 273.942 33.932 274.556 ; 
        RECT 33.536 274.044 33.608 275.076 ; 
        RECT 31.376 271.488 31.448 275.23 ; 
        RECT 31.232 271.488 31.304 275.23 ; 
        RECT 31.088 272.212 31.16 274.484 ; 
        RECT 34.796 275.808 34.868 279.55 ; 
        RECT 34.652 275.808 34.724 279.55 ; 
        RECT 34.508 278.116 34.58 279.406 ; 
        RECT 34.04 278.904 34.112 279.342 ; 
        RECT 34.004 275.938 34.076 276.896 ; 
        RECT 33.86 278.262 33.932 278.876 ; 
        RECT 33.536 278.364 33.608 279.396 ; 
        RECT 31.376 275.808 31.448 279.55 ; 
        RECT 31.232 275.808 31.304 279.55 ; 
        RECT 31.088 276.532 31.16 278.804 ; 
        RECT 34.796 280.128 34.868 283.87 ; 
        RECT 34.652 280.128 34.724 283.87 ; 
        RECT 34.508 282.436 34.58 283.726 ; 
        RECT 34.04 283.224 34.112 283.662 ; 
        RECT 34.004 280.258 34.076 281.216 ; 
        RECT 33.86 282.582 33.932 283.196 ; 
        RECT 33.536 282.684 33.608 283.716 ; 
        RECT 31.376 280.128 31.448 283.87 ; 
        RECT 31.232 280.128 31.304 283.87 ; 
        RECT 31.088 280.852 31.16 283.124 ; 
        RECT 34.796 284.448 34.868 288.19 ; 
        RECT 34.652 284.448 34.724 288.19 ; 
        RECT 34.508 286.756 34.58 288.046 ; 
        RECT 34.04 287.544 34.112 287.982 ; 
        RECT 34.004 284.578 34.076 285.536 ; 
        RECT 33.86 286.902 33.932 287.516 ; 
        RECT 33.536 287.004 33.608 288.036 ; 
        RECT 31.376 284.448 31.448 288.19 ; 
        RECT 31.232 284.448 31.304 288.19 ; 
        RECT 31.088 285.172 31.16 287.444 ; 
        RECT 34.796 288.768 34.868 292.51 ; 
        RECT 34.652 288.768 34.724 292.51 ; 
        RECT 34.508 291.076 34.58 292.366 ; 
        RECT 34.04 291.864 34.112 292.302 ; 
        RECT 34.004 288.898 34.076 289.856 ; 
        RECT 33.86 291.222 33.932 291.836 ; 
        RECT 33.536 291.324 33.608 292.356 ; 
        RECT 31.376 288.768 31.448 292.51 ; 
        RECT 31.232 288.768 31.304 292.51 ; 
        RECT 31.088 289.492 31.16 291.764 ; 
        RECT 34.796 293.088 34.868 296.83 ; 
        RECT 34.652 293.088 34.724 296.83 ; 
        RECT 34.508 295.396 34.58 296.686 ; 
        RECT 34.04 296.184 34.112 296.622 ; 
        RECT 34.004 293.218 34.076 294.176 ; 
        RECT 33.86 295.542 33.932 296.156 ; 
        RECT 33.536 295.644 33.608 296.676 ; 
        RECT 31.376 293.088 31.448 296.83 ; 
        RECT 31.232 293.088 31.304 296.83 ; 
        RECT 31.088 293.812 31.16 296.084 ; 
        RECT 34.796 297.408 34.868 301.15 ; 
        RECT 34.652 297.408 34.724 301.15 ; 
        RECT 34.508 299.716 34.58 301.006 ; 
        RECT 34.04 300.504 34.112 300.942 ; 
        RECT 34.004 297.538 34.076 298.496 ; 
        RECT 33.86 299.862 33.932 300.476 ; 
        RECT 33.536 299.964 33.608 300.996 ; 
        RECT 31.376 297.408 31.448 301.15 ; 
        RECT 31.232 297.408 31.304 301.15 ; 
        RECT 31.088 298.132 31.16 300.404 ; 
        RECT 34.796 301.728 34.868 305.47 ; 
        RECT 34.652 301.728 34.724 305.47 ; 
        RECT 34.508 304.036 34.58 305.326 ; 
        RECT 34.04 304.824 34.112 305.262 ; 
        RECT 34.004 301.858 34.076 302.816 ; 
        RECT 33.86 304.182 33.932 304.796 ; 
        RECT 33.536 304.284 33.608 305.316 ; 
        RECT 31.376 301.728 31.448 305.47 ; 
        RECT 31.232 301.728 31.304 305.47 ; 
        RECT 31.088 302.452 31.16 304.724 ; 
        RECT 34.796 306.048 34.868 309.79 ; 
        RECT 34.652 306.048 34.724 309.79 ; 
        RECT 34.508 308.356 34.58 309.646 ; 
        RECT 34.04 309.144 34.112 309.582 ; 
        RECT 34.004 306.178 34.076 307.136 ; 
        RECT 33.86 308.502 33.932 309.116 ; 
        RECT 33.536 308.604 33.608 309.636 ; 
        RECT 31.376 306.048 31.448 309.79 ; 
        RECT 31.232 306.048 31.304 309.79 ; 
        RECT 31.088 306.772 31.16 309.044 ; 
        RECT 34.796 310.368 34.868 314.11 ; 
        RECT 34.652 310.368 34.724 314.11 ; 
        RECT 34.508 312.676 34.58 313.966 ; 
        RECT 34.04 313.464 34.112 313.902 ; 
        RECT 34.004 310.498 34.076 311.456 ; 
        RECT 33.86 312.822 33.932 313.436 ; 
        RECT 33.536 312.924 33.608 313.956 ; 
        RECT 31.376 310.368 31.448 314.11 ; 
        RECT 31.232 310.368 31.304 314.11 ; 
        RECT 31.088 311.092 31.16 313.364 ; 
        RECT 34.796 314.688 34.868 318.43 ; 
        RECT 34.652 314.688 34.724 318.43 ; 
        RECT 34.508 316.996 34.58 318.286 ; 
        RECT 34.04 317.784 34.112 318.222 ; 
        RECT 34.004 314.818 34.076 315.776 ; 
        RECT 33.86 317.142 33.932 317.756 ; 
        RECT 33.536 317.244 33.608 318.276 ; 
        RECT 31.376 314.688 31.448 318.43 ; 
        RECT 31.232 314.688 31.304 318.43 ; 
        RECT 31.088 315.412 31.16 317.684 ; 
        RECT 34.796 319.008 34.868 322.75 ; 
        RECT 34.652 319.008 34.724 322.75 ; 
        RECT 34.508 321.316 34.58 322.606 ; 
        RECT 34.04 322.104 34.112 322.542 ; 
        RECT 34.004 319.138 34.076 320.096 ; 
        RECT 33.86 321.462 33.932 322.076 ; 
        RECT 33.536 321.564 33.608 322.596 ; 
        RECT 31.376 319.008 31.448 322.75 ; 
        RECT 31.232 319.008 31.304 322.75 ; 
        RECT 31.088 319.732 31.16 322.004 ; 
        RECT 34.796 323.328 34.868 327.07 ; 
        RECT 34.652 323.328 34.724 327.07 ; 
        RECT 34.508 325.636 34.58 326.926 ; 
        RECT 34.04 326.424 34.112 326.862 ; 
        RECT 34.004 323.458 34.076 324.416 ; 
        RECT 33.86 325.782 33.932 326.396 ; 
        RECT 33.536 325.884 33.608 326.916 ; 
        RECT 31.376 323.328 31.448 327.07 ; 
        RECT 31.232 323.328 31.304 327.07 ; 
        RECT 31.088 324.052 31.16 326.324 ; 
        RECT 34.796 327.648 34.868 331.39 ; 
        RECT 34.652 327.648 34.724 331.39 ; 
        RECT 34.508 329.956 34.58 331.246 ; 
        RECT 34.04 330.744 34.112 331.182 ; 
        RECT 34.004 327.778 34.076 328.736 ; 
        RECT 33.86 330.102 33.932 330.716 ; 
        RECT 33.536 330.204 33.608 331.236 ; 
        RECT 31.376 327.648 31.448 331.39 ; 
        RECT 31.232 327.648 31.304 331.39 ; 
        RECT 31.088 328.372 31.16 330.644 ; 
        RECT 34.796 331.968 34.868 335.71 ; 
        RECT 34.652 331.968 34.724 335.71 ; 
        RECT 34.508 334.276 34.58 335.566 ; 
        RECT 34.04 335.064 34.112 335.502 ; 
        RECT 34.004 332.098 34.076 333.056 ; 
        RECT 33.86 334.422 33.932 335.036 ; 
        RECT 33.536 334.524 33.608 335.556 ; 
        RECT 31.376 331.968 31.448 335.71 ; 
        RECT 31.232 331.968 31.304 335.71 ; 
        RECT 31.088 332.692 31.16 334.964 ; 
        RECT 34.796 336.288 34.868 340.03 ; 
        RECT 34.652 336.288 34.724 340.03 ; 
        RECT 34.508 338.596 34.58 339.886 ; 
        RECT 34.04 339.384 34.112 339.822 ; 
        RECT 34.004 336.418 34.076 337.376 ; 
        RECT 33.86 338.742 33.932 339.356 ; 
        RECT 33.536 338.844 33.608 339.876 ; 
        RECT 31.376 336.288 31.448 340.03 ; 
        RECT 31.232 336.288 31.304 340.03 ; 
        RECT 31.088 337.012 31.16 339.284 ; 
        RECT 34.796 340.608 34.868 344.35 ; 
        RECT 34.652 340.608 34.724 344.35 ; 
        RECT 34.508 342.916 34.58 344.206 ; 
        RECT 34.04 343.704 34.112 344.142 ; 
        RECT 34.004 340.738 34.076 341.696 ; 
        RECT 33.86 343.062 33.932 343.676 ; 
        RECT 33.536 343.164 33.608 344.196 ; 
        RECT 31.376 340.608 31.448 344.35 ; 
        RECT 31.232 340.608 31.304 344.35 ; 
        RECT 31.088 341.332 31.16 343.604 ; 
        RECT 34.796 344.928 34.868 348.67 ; 
        RECT 34.652 344.928 34.724 348.67 ; 
        RECT 34.508 347.236 34.58 348.526 ; 
        RECT 34.04 348.024 34.112 348.462 ; 
        RECT 34.004 345.058 34.076 346.016 ; 
        RECT 33.86 347.382 33.932 347.996 ; 
        RECT 33.536 347.484 33.608 348.516 ; 
        RECT 31.376 344.928 31.448 348.67 ; 
        RECT 31.232 344.928 31.304 348.67 ; 
        RECT 31.088 345.652 31.16 347.924 ; 
        RECT 34.796 349.248 34.868 352.99 ; 
        RECT 34.652 349.248 34.724 352.99 ; 
        RECT 34.508 351.556 34.58 352.846 ; 
        RECT 34.04 352.344 34.112 352.782 ; 
        RECT 34.004 349.378 34.076 350.336 ; 
        RECT 33.86 351.702 33.932 352.316 ; 
        RECT 33.536 351.804 33.608 352.836 ; 
        RECT 31.376 349.248 31.448 352.99 ; 
        RECT 31.232 349.248 31.304 352.99 ; 
        RECT 31.088 349.972 31.16 352.244 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 34.564 1.026 35.076 5.4 ; 
      RECT 34.508 3.688 35.076 4.978 ; 
      RECT 33.916 2.596 34.164 5.4 ; 
      RECT 33.86 3.834 34.164 4.448 ; 
      RECT 33.916 1.026 34.02 5.4 ; 
      RECT 33.916 1.51 34.076 2.468 ; 
      RECT 33.916 1.026 34.164 1.382 ; 
      RECT 32.728 2.828 33.552 5.4 ; 
      RECT 33.448 1.026 33.552 5.4 ; 
      RECT 32.728 3.936 33.608 4.968 ; 
      RECT 32.728 1.026 33.12 5.4 ; 
      RECT 31.06 1.026 31.392 5.4 ; 
      RECT 31.06 1.38 31.448 5.122 ; 
      RECT 65.776 1.026 66.116 5.4 ; 
      RECT 65.2 1.026 65.304 5.4 ; 
      RECT 64.768 1.026 64.872 5.4 ; 
      RECT 64.336 1.026 64.44 5.4 ; 
      RECT 63.904 1.026 64.008 5.4 ; 
      RECT 63.472 1.026 63.576 5.4 ; 
      RECT 63.04 1.026 63.144 5.4 ; 
      RECT 62.608 1.026 62.712 5.4 ; 
      RECT 62.176 1.026 62.28 5.4 ; 
      RECT 61.744 1.026 61.848 5.4 ; 
      RECT 61.312 1.026 61.416 5.4 ; 
      RECT 60.88 1.026 60.984 5.4 ; 
      RECT 60.448 1.026 60.552 5.4 ; 
      RECT 60.016 1.026 60.12 5.4 ; 
      RECT 59.584 1.026 59.688 5.4 ; 
      RECT 59.152 1.026 59.256 5.4 ; 
      RECT 58.72 1.026 58.824 5.4 ; 
      RECT 58.288 1.026 58.392 5.4 ; 
      RECT 57.856 1.026 57.96 5.4 ; 
      RECT 57.424 1.026 57.528 5.4 ; 
      RECT 56.992 1.026 57.096 5.4 ; 
      RECT 56.56 1.026 56.664 5.4 ; 
      RECT 56.128 1.026 56.232 5.4 ; 
      RECT 55.696 1.026 55.8 5.4 ; 
      RECT 55.264 1.026 55.368 5.4 ; 
      RECT 54.832 1.026 54.936 5.4 ; 
      RECT 54.4 1.026 54.504 5.4 ; 
      RECT 53.968 1.026 54.072 5.4 ; 
      RECT 53.536 1.026 53.64 5.4 ; 
      RECT 53.104 1.026 53.208 5.4 ; 
      RECT 52.672 1.026 52.776 5.4 ; 
      RECT 52.24 1.026 52.344 5.4 ; 
      RECT 51.808 1.026 51.912 5.4 ; 
      RECT 51.376 1.026 51.48 5.4 ; 
      RECT 50.944 1.026 51.048 5.4 ; 
      RECT 50.512 1.026 50.616 5.4 ; 
      RECT 50.08 1.026 50.184 5.4 ; 
      RECT 49.648 1.026 49.752 5.4 ; 
      RECT 49.216 1.026 49.32 5.4 ; 
      RECT 48.784 1.026 48.888 5.4 ; 
      RECT 48.352 1.026 48.456 5.4 ; 
      RECT 47.92 1.026 48.024 5.4 ; 
      RECT 47.488 1.026 47.592 5.4 ; 
      RECT 47.056 1.026 47.16 5.4 ; 
      RECT 46.624 1.026 46.728 5.4 ; 
      RECT 46.192 1.026 46.296 5.4 ; 
      RECT 45.76 1.026 45.864 5.4 ; 
      RECT 45.328 1.026 45.432 5.4 ; 
      RECT 44.896 1.026 45 5.4 ; 
      RECT 44.464 1.026 44.568 5.4 ; 
      RECT 44.032 1.026 44.136 5.4 ; 
      RECT 43.6 1.026 43.704 5.4 ; 
      RECT 43.168 1.026 43.272 5.4 ; 
      RECT 42.736 1.026 42.84 5.4 ; 
      RECT 42.304 1.026 42.408 5.4 ; 
      RECT 41.872 1.026 41.976 5.4 ; 
      RECT 41.44 1.026 41.544 5.4 ; 
      RECT 41.008 1.026 41.112 5.4 ; 
      RECT 40.576 1.026 40.68 5.4 ; 
      RECT 40.144 1.026 40.248 5.4 ; 
      RECT 39.712 1.026 39.816 5.4 ; 
      RECT 39.28 1.026 39.384 5.4 ; 
      RECT 38.848 1.026 38.952 5.4 ; 
      RECT 38.416 1.026 38.52 5.4 ; 
      RECT 37.984 1.026 38.088 5.4 ; 
      RECT 37.552 1.026 37.656 5.4 ; 
      RECT 36.7 1.026 37.008 5.4 ; 
      RECT 29.128 1.026 29.436 5.4 ; 
      RECT 28.48 1.026 28.584 5.4 ; 
      RECT 28.048 1.026 28.152 5.4 ; 
      RECT 27.616 1.026 27.72 5.4 ; 
      RECT 27.184 1.026 27.288 5.4 ; 
      RECT 26.752 1.026 26.856 5.4 ; 
      RECT 26.32 1.026 26.424 5.4 ; 
      RECT 25.888 1.026 25.992 5.4 ; 
      RECT 25.456 1.026 25.56 5.4 ; 
      RECT 25.024 1.026 25.128 5.4 ; 
      RECT 24.592 1.026 24.696 5.4 ; 
      RECT 24.16 1.026 24.264 5.4 ; 
      RECT 23.728 1.026 23.832 5.4 ; 
      RECT 23.296 1.026 23.4 5.4 ; 
      RECT 22.864 1.026 22.968 5.4 ; 
      RECT 22.432 1.026 22.536 5.4 ; 
      RECT 22 1.026 22.104 5.4 ; 
      RECT 21.568 1.026 21.672 5.4 ; 
      RECT 21.136 1.026 21.24 5.4 ; 
      RECT 20.704 1.026 20.808 5.4 ; 
      RECT 20.272 1.026 20.376 5.4 ; 
      RECT 19.84 1.026 19.944 5.4 ; 
      RECT 19.408 1.026 19.512 5.4 ; 
      RECT 18.976 1.026 19.08 5.4 ; 
      RECT 18.544 1.026 18.648 5.4 ; 
      RECT 18.112 1.026 18.216 5.4 ; 
      RECT 17.68 1.026 17.784 5.4 ; 
      RECT 17.248 1.026 17.352 5.4 ; 
      RECT 16.816 1.026 16.92 5.4 ; 
      RECT 16.384 1.026 16.488 5.4 ; 
      RECT 15.952 1.026 16.056 5.4 ; 
      RECT 15.52 1.026 15.624 5.4 ; 
      RECT 15.088 1.026 15.192 5.4 ; 
      RECT 14.656 1.026 14.76 5.4 ; 
      RECT 14.224 1.026 14.328 5.4 ; 
      RECT 13.792 1.026 13.896 5.4 ; 
      RECT 13.36 1.026 13.464 5.4 ; 
      RECT 12.928 1.026 13.032 5.4 ; 
      RECT 12.496 1.026 12.6 5.4 ; 
      RECT 12.064 1.026 12.168 5.4 ; 
      RECT 11.632 1.026 11.736 5.4 ; 
      RECT 11.2 1.026 11.304 5.4 ; 
      RECT 10.768 1.026 10.872 5.4 ; 
      RECT 10.336 1.026 10.44 5.4 ; 
      RECT 9.904 1.026 10.008 5.4 ; 
      RECT 9.472 1.026 9.576 5.4 ; 
      RECT 9.04 1.026 9.144 5.4 ; 
      RECT 8.608 1.026 8.712 5.4 ; 
      RECT 8.176 1.026 8.28 5.4 ; 
      RECT 7.744 1.026 7.848 5.4 ; 
      RECT 7.312 1.026 7.416 5.4 ; 
      RECT 6.88 1.026 6.984 5.4 ; 
      RECT 6.448 1.026 6.552 5.4 ; 
      RECT 6.016 1.026 6.12 5.4 ; 
      RECT 5.584 1.026 5.688 5.4 ; 
      RECT 5.152 1.026 5.256 5.4 ; 
      RECT 4.72 1.026 4.824 5.4 ; 
      RECT 4.288 1.026 4.392 5.4 ; 
      RECT 3.856 1.026 3.96 5.4 ; 
      RECT 3.424 1.026 3.528 5.4 ; 
      RECT 2.992 1.026 3.096 5.4 ; 
      RECT 2.56 1.026 2.664 5.4 ; 
      RECT 2.128 1.026 2.232 5.4 ; 
      RECT 1.696 1.026 1.8 5.4 ; 
      RECT 1.264 1.026 1.368 5.4 ; 
      RECT 0.832 1.026 0.936 5.4 ; 
      RECT 0.02 1.026 0.36 5.4 ; 
      RECT 34.564 5.346 35.076 9.72 ; 
      RECT 34.508 8.008 35.076 9.298 ; 
      RECT 33.916 6.916 34.164 9.72 ; 
      RECT 33.86 8.154 34.164 8.768 ; 
      RECT 33.916 5.346 34.02 9.72 ; 
      RECT 33.916 5.83 34.076 6.788 ; 
      RECT 33.916 5.346 34.164 5.702 ; 
      RECT 32.728 7.148 33.552 9.72 ; 
      RECT 33.448 5.346 33.552 9.72 ; 
      RECT 32.728 8.256 33.608 9.288 ; 
      RECT 32.728 5.346 33.12 9.72 ; 
      RECT 31.06 5.346 31.392 9.72 ; 
      RECT 31.06 5.7 31.448 9.442 ; 
      RECT 65.776 5.346 66.116 9.72 ; 
      RECT 65.2 5.346 65.304 9.72 ; 
      RECT 64.768 5.346 64.872 9.72 ; 
      RECT 64.336 5.346 64.44 9.72 ; 
      RECT 63.904 5.346 64.008 9.72 ; 
      RECT 63.472 5.346 63.576 9.72 ; 
      RECT 63.04 5.346 63.144 9.72 ; 
      RECT 62.608 5.346 62.712 9.72 ; 
      RECT 62.176 5.346 62.28 9.72 ; 
      RECT 61.744 5.346 61.848 9.72 ; 
      RECT 61.312 5.346 61.416 9.72 ; 
      RECT 60.88 5.346 60.984 9.72 ; 
      RECT 60.448 5.346 60.552 9.72 ; 
      RECT 60.016 5.346 60.12 9.72 ; 
      RECT 59.584 5.346 59.688 9.72 ; 
      RECT 59.152 5.346 59.256 9.72 ; 
      RECT 58.72 5.346 58.824 9.72 ; 
      RECT 58.288 5.346 58.392 9.72 ; 
      RECT 57.856 5.346 57.96 9.72 ; 
      RECT 57.424 5.346 57.528 9.72 ; 
      RECT 56.992 5.346 57.096 9.72 ; 
      RECT 56.56 5.346 56.664 9.72 ; 
      RECT 56.128 5.346 56.232 9.72 ; 
      RECT 55.696 5.346 55.8 9.72 ; 
      RECT 55.264 5.346 55.368 9.72 ; 
      RECT 54.832 5.346 54.936 9.72 ; 
      RECT 54.4 5.346 54.504 9.72 ; 
      RECT 53.968 5.346 54.072 9.72 ; 
      RECT 53.536 5.346 53.64 9.72 ; 
      RECT 53.104 5.346 53.208 9.72 ; 
      RECT 52.672 5.346 52.776 9.72 ; 
      RECT 52.24 5.346 52.344 9.72 ; 
      RECT 51.808 5.346 51.912 9.72 ; 
      RECT 51.376 5.346 51.48 9.72 ; 
      RECT 50.944 5.346 51.048 9.72 ; 
      RECT 50.512 5.346 50.616 9.72 ; 
      RECT 50.08 5.346 50.184 9.72 ; 
      RECT 49.648 5.346 49.752 9.72 ; 
      RECT 49.216 5.346 49.32 9.72 ; 
      RECT 48.784 5.346 48.888 9.72 ; 
      RECT 48.352 5.346 48.456 9.72 ; 
      RECT 47.92 5.346 48.024 9.72 ; 
      RECT 47.488 5.346 47.592 9.72 ; 
      RECT 47.056 5.346 47.16 9.72 ; 
      RECT 46.624 5.346 46.728 9.72 ; 
      RECT 46.192 5.346 46.296 9.72 ; 
      RECT 45.76 5.346 45.864 9.72 ; 
      RECT 45.328 5.346 45.432 9.72 ; 
      RECT 44.896 5.346 45 9.72 ; 
      RECT 44.464 5.346 44.568 9.72 ; 
      RECT 44.032 5.346 44.136 9.72 ; 
      RECT 43.6 5.346 43.704 9.72 ; 
      RECT 43.168 5.346 43.272 9.72 ; 
      RECT 42.736 5.346 42.84 9.72 ; 
      RECT 42.304 5.346 42.408 9.72 ; 
      RECT 41.872 5.346 41.976 9.72 ; 
      RECT 41.44 5.346 41.544 9.72 ; 
      RECT 41.008 5.346 41.112 9.72 ; 
      RECT 40.576 5.346 40.68 9.72 ; 
      RECT 40.144 5.346 40.248 9.72 ; 
      RECT 39.712 5.346 39.816 9.72 ; 
      RECT 39.28 5.346 39.384 9.72 ; 
      RECT 38.848 5.346 38.952 9.72 ; 
      RECT 38.416 5.346 38.52 9.72 ; 
      RECT 37.984 5.346 38.088 9.72 ; 
      RECT 37.552 5.346 37.656 9.72 ; 
      RECT 36.7 5.346 37.008 9.72 ; 
      RECT 29.128 5.346 29.436 9.72 ; 
      RECT 28.48 5.346 28.584 9.72 ; 
      RECT 28.048 5.346 28.152 9.72 ; 
      RECT 27.616 5.346 27.72 9.72 ; 
      RECT 27.184 5.346 27.288 9.72 ; 
      RECT 26.752 5.346 26.856 9.72 ; 
      RECT 26.32 5.346 26.424 9.72 ; 
      RECT 25.888 5.346 25.992 9.72 ; 
      RECT 25.456 5.346 25.56 9.72 ; 
      RECT 25.024 5.346 25.128 9.72 ; 
      RECT 24.592 5.346 24.696 9.72 ; 
      RECT 24.16 5.346 24.264 9.72 ; 
      RECT 23.728 5.346 23.832 9.72 ; 
      RECT 23.296 5.346 23.4 9.72 ; 
      RECT 22.864 5.346 22.968 9.72 ; 
      RECT 22.432 5.346 22.536 9.72 ; 
      RECT 22 5.346 22.104 9.72 ; 
      RECT 21.568 5.346 21.672 9.72 ; 
      RECT 21.136 5.346 21.24 9.72 ; 
      RECT 20.704 5.346 20.808 9.72 ; 
      RECT 20.272 5.346 20.376 9.72 ; 
      RECT 19.84 5.346 19.944 9.72 ; 
      RECT 19.408 5.346 19.512 9.72 ; 
      RECT 18.976 5.346 19.08 9.72 ; 
      RECT 18.544 5.346 18.648 9.72 ; 
      RECT 18.112 5.346 18.216 9.72 ; 
      RECT 17.68 5.346 17.784 9.72 ; 
      RECT 17.248 5.346 17.352 9.72 ; 
      RECT 16.816 5.346 16.92 9.72 ; 
      RECT 16.384 5.346 16.488 9.72 ; 
      RECT 15.952 5.346 16.056 9.72 ; 
      RECT 15.52 5.346 15.624 9.72 ; 
      RECT 15.088 5.346 15.192 9.72 ; 
      RECT 14.656 5.346 14.76 9.72 ; 
      RECT 14.224 5.346 14.328 9.72 ; 
      RECT 13.792 5.346 13.896 9.72 ; 
      RECT 13.36 5.346 13.464 9.72 ; 
      RECT 12.928 5.346 13.032 9.72 ; 
      RECT 12.496 5.346 12.6 9.72 ; 
      RECT 12.064 5.346 12.168 9.72 ; 
      RECT 11.632 5.346 11.736 9.72 ; 
      RECT 11.2 5.346 11.304 9.72 ; 
      RECT 10.768 5.346 10.872 9.72 ; 
      RECT 10.336 5.346 10.44 9.72 ; 
      RECT 9.904 5.346 10.008 9.72 ; 
      RECT 9.472 5.346 9.576 9.72 ; 
      RECT 9.04 5.346 9.144 9.72 ; 
      RECT 8.608 5.346 8.712 9.72 ; 
      RECT 8.176 5.346 8.28 9.72 ; 
      RECT 7.744 5.346 7.848 9.72 ; 
      RECT 7.312 5.346 7.416 9.72 ; 
      RECT 6.88 5.346 6.984 9.72 ; 
      RECT 6.448 5.346 6.552 9.72 ; 
      RECT 6.016 5.346 6.12 9.72 ; 
      RECT 5.584 5.346 5.688 9.72 ; 
      RECT 5.152 5.346 5.256 9.72 ; 
      RECT 4.72 5.346 4.824 9.72 ; 
      RECT 4.288 5.346 4.392 9.72 ; 
      RECT 3.856 5.346 3.96 9.72 ; 
      RECT 3.424 5.346 3.528 9.72 ; 
      RECT 2.992 5.346 3.096 9.72 ; 
      RECT 2.56 5.346 2.664 9.72 ; 
      RECT 2.128 5.346 2.232 9.72 ; 
      RECT 1.696 5.346 1.8 9.72 ; 
      RECT 1.264 5.346 1.368 9.72 ; 
      RECT 0.832 5.346 0.936 9.72 ; 
      RECT 0.02 5.346 0.36 9.72 ; 
      RECT 34.564 9.666 35.076 14.04 ; 
      RECT 34.508 12.328 35.076 13.618 ; 
      RECT 33.916 11.236 34.164 14.04 ; 
      RECT 33.86 12.474 34.164 13.088 ; 
      RECT 33.916 9.666 34.02 14.04 ; 
      RECT 33.916 10.15 34.076 11.108 ; 
      RECT 33.916 9.666 34.164 10.022 ; 
      RECT 32.728 11.468 33.552 14.04 ; 
      RECT 33.448 9.666 33.552 14.04 ; 
      RECT 32.728 12.576 33.608 13.608 ; 
      RECT 32.728 9.666 33.12 14.04 ; 
      RECT 31.06 9.666 31.392 14.04 ; 
      RECT 31.06 10.02 31.448 13.762 ; 
      RECT 65.776 9.666 66.116 14.04 ; 
      RECT 65.2 9.666 65.304 14.04 ; 
      RECT 64.768 9.666 64.872 14.04 ; 
      RECT 64.336 9.666 64.44 14.04 ; 
      RECT 63.904 9.666 64.008 14.04 ; 
      RECT 63.472 9.666 63.576 14.04 ; 
      RECT 63.04 9.666 63.144 14.04 ; 
      RECT 62.608 9.666 62.712 14.04 ; 
      RECT 62.176 9.666 62.28 14.04 ; 
      RECT 61.744 9.666 61.848 14.04 ; 
      RECT 61.312 9.666 61.416 14.04 ; 
      RECT 60.88 9.666 60.984 14.04 ; 
      RECT 60.448 9.666 60.552 14.04 ; 
      RECT 60.016 9.666 60.12 14.04 ; 
      RECT 59.584 9.666 59.688 14.04 ; 
      RECT 59.152 9.666 59.256 14.04 ; 
      RECT 58.72 9.666 58.824 14.04 ; 
      RECT 58.288 9.666 58.392 14.04 ; 
      RECT 57.856 9.666 57.96 14.04 ; 
      RECT 57.424 9.666 57.528 14.04 ; 
      RECT 56.992 9.666 57.096 14.04 ; 
      RECT 56.56 9.666 56.664 14.04 ; 
      RECT 56.128 9.666 56.232 14.04 ; 
      RECT 55.696 9.666 55.8 14.04 ; 
      RECT 55.264 9.666 55.368 14.04 ; 
      RECT 54.832 9.666 54.936 14.04 ; 
      RECT 54.4 9.666 54.504 14.04 ; 
      RECT 53.968 9.666 54.072 14.04 ; 
      RECT 53.536 9.666 53.64 14.04 ; 
      RECT 53.104 9.666 53.208 14.04 ; 
      RECT 52.672 9.666 52.776 14.04 ; 
      RECT 52.24 9.666 52.344 14.04 ; 
      RECT 51.808 9.666 51.912 14.04 ; 
      RECT 51.376 9.666 51.48 14.04 ; 
      RECT 50.944 9.666 51.048 14.04 ; 
      RECT 50.512 9.666 50.616 14.04 ; 
      RECT 50.08 9.666 50.184 14.04 ; 
      RECT 49.648 9.666 49.752 14.04 ; 
      RECT 49.216 9.666 49.32 14.04 ; 
      RECT 48.784 9.666 48.888 14.04 ; 
      RECT 48.352 9.666 48.456 14.04 ; 
      RECT 47.92 9.666 48.024 14.04 ; 
      RECT 47.488 9.666 47.592 14.04 ; 
      RECT 47.056 9.666 47.16 14.04 ; 
      RECT 46.624 9.666 46.728 14.04 ; 
      RECT 46.192 9.666 46.296 14.04 ; 
      RECT 45.76 9.666 45.864 14.04 ; 
      RECT 45.328 9.666 45.432 14.04 ; 
      RECT 44.896 9.666 45 14.04 ; 
      RECT 44.464 9.666 44.568 14.04 ; 
      RECT 44.032 9.666 44.136 14.04 ; 
      RECT 43.6 9.666 43.704 14.04 ; 
      RECT 43.168 9.666 43.272 14.04 ; 
      RECT 42.736 9.666 42.84 14.04 ; 
      RECT 42.304 9.666 42.408 14.04 ; 
      RECT 41.872 9.666 41.976 14.04 ; 
      RECT 41.44 9.666 41.544 14.04 ; 
      RECT 41.008 9.666 41.112 14.04 ; 
      RECT 40.576 9.666 40.68 14.04 ; 
      RECT 40.144 9.666 40.248 14.04 ; 
      RECT 39.712 9.666 39.816 14.04 ; 
      RECT 39.28 9.666 39.384 14.04 ; 
      RECT 38.848 9.666 38.952 14.04 ; 
      RECT 38.416 9.666 38.52 14.04 ; 
      RECT 37.984 9.666 38.088 14.04 ; 
      RECT 37.552 9.666 37.656 14.04 ; 
      RECT 36.7 9.666 37.008 14.04 ; 
      RECT 29.128 9.666 29.436 14.04 ; 
      RECT 28.48 9.666 28.584 14.04 ; 
      RECT 28.048 9.666 28.152 14.04 ; 
      RECT 27.616 9.666 27.72 14.04 ; 
      RECT 27.184 9.666 27.288 14.04 ; 
      RECT 26.752 9.666 26.856 14.04 ; 
      RECT 26.32 9.666 26.424 14.04 ; 
      RECT 25.888 9.666 25.992 14.04 ; 
      RECT 25.456 9.666 25.56 14.04 ; 
      RECT 25.024 9.666 25.128 14.04 ; 
      RECT 24.592 9.666 24.696 14.04 ; 
      RECT 24.16 9.666 24.264 14.04 ; 
      RECT 23.728 9.666 23.832 14.04 ; 
      RECT 23.296 9.666 23.4 14.04 ; 
      RECT 22.864 9.666 22.968 14.04 ; 
      RECT 22.432 9.666 22.536 14.04 ; 
      RECT 22 9.666 22.104 14.04 ; 
      RECT 21.568 9.666 21.672 14.04 ; 
      RECT 21.136 9.666 21.24 14.04 ; 
      RECT 20.704 9.666 20.808 14.04 ; 
      RECT 20.272 9.666 20.376 14.04 ; 
      RECT 19.84 9.666 19.944 14.04 ; 
      RECT 19.408 9.666 19.512 14.04 ; 
      RECT 18.976 9.666 19.08 14.04 ; 
      RECT 18.544 9.666 18.648 14.04 ; 
      RECT 18.112 9.666 18.216 14.04 ; 
      RECT 17.68 9.666 17.784 14.04 ; 
      RECT 17.248 9.666 17.352 14.04 ; 
      RECT 16.816 9.666 16.92 14.04 ; 
      RECT 16.384 9.666 16.488 14.04 ; 
      RECT 15.952 9.666 16.056 14.04 ; 
      RECT 15.52 9.666 15.624 14.04 ; 
      RECT 15.088 9.666 15.192 14.04 ; 
      RECT 14.656 9.666 14.76 14.04 ; 
      RECT 14.224 9.666 14.328 14.04 ; 
      RECT 13.792 9.666 13.896 14.04 ; 
      RECT 13.36 9.666 13.464 14.04 ; 
      RECT 12.928 9.666 13.032 14.04 ; 
      RECT 12.496 9.666 12.6 14.04 ; 
      RECT 12.064 9.666 12.168 14.04 ; 
      RECT 11.632 9.666 11.736 14.04 ; 
      RECT 11.2 9.666 11.304 14.04 ; 
      RECT 10.768 9.666 10.872 14.04 ; 
      RECT 10.336 9.666 10.44 14.04 ; 
      RECT 9.904 9.666 10.008 14.04 ; 
      RECT 9.472 9.666 9.576 14.04 ; 
      RECT 9.04 9.666 9.144 14.04 ; 
      RECT 8.608 9.666 8.712 14.04 ; 
      RECT 8.176 9.666 8.28 14.04 ; 
      RECT 7.744 9.666 7.848 14.04 ; 
      RECT 7.312 9.666 7.416 14.04 ; 
      RECT 6.88 9.666 6.984 14.04 ; 
      RECT 6.448 9.666 6.552 14.04 ; 
      RECT 6.016 9.666 6.12 14.04 ; 
      RECT 5.584 9.666 5.688 14.04 ; 
      RECT 5.152 9.666 5.256 14.04 ; 
      RECT 4.72 9.666 4.824 14.04 ; 
      RECT 4.288 9.666 4.392 14.04 ; 
      RECT 3.856 9.666 3.96 14.04 ; 
      RECT 3.424 9.666 3.528 14.04 ; 
      RECT 2.992 9.666 3.096 14.04 ; 
      RECT 2.56 9.666 2.664 14.04 ; 
      RECT 2.128 9.666 2.232 14.04 ; 
      RECT 1.696 9.666 1.8 14.04 ; 
      RECT 1.264 9.666 1.368 14.04 ; 
      RECT 0.832 9.666 0.936 14.04 ; 
      RECT 0.02 9.666 0.36 14.04 ; 
      RECT 34.564 13.986 35.076 18.36 ; 
      RECT 34.508 16.648 35.076 17.938 ; 
      RECT 33.916 15.556 34.164 18.36 ; 
      RECT 33.86 16.794 34.164 17.408 ; 
      RECT 33.916 13.986 34.02 18.36 ; 
      RECT 33.916 14.47 34.076 15.428 ; 
      RECT 33.916 13.986 34.164 14.342 ; 
      RECT 32.728 15.788 33.552 18.36 ; 
      RECT 33.448 13.986 33.552 18.36 ; 
      RECT 32.728 16.896 33.608 17.928 ; 
      RECT 32.728 13.986 33.12 18.36 ; 
      RECT 31.06 13.986 31.392 18.36 ; 
      RECT 31.06 14.34 31.448 18.082 ; 
      RECT 65.776 13.986 66.116 18.36 ; 
      RECT 65.2 13.986 65.304 18.36 ; 
      RECT 64.768 13.986 64.872 18.36 ; 
      RECT 64.336 13.986 64.44 18.36 ; 
      RECT 63.904 13.986 64.008 18.36 ; 
      RECT 63.472 13.986 63.576 18.36 ; 
      RECT 63.04 13.986 63.144 18.36 ; 
      RECT 62.608 13.986 62.712 18.36 ; 
      RECT 62.176 13.986 62.28 18.36 ; 
      RECT 61.744 13.986 61.848 18.36 ; 
      RECT 61.312 13.986 61.416 18.36 ; 
      RECT 60.88 13.986 60.984 18.36 ; 
      RECT 60.448 13.986 60.552 18.36 ; 
      RECT 60.016 13.986 60.12 18.36 ; 
      RECT 59.584 13.986 59.688 18.36 ; 
      RECT 59.152 13.986 59.256 18.36 ; 
      RECT 58.72 13.986 58.824 18.36 ; 
      RECT 58.288 13.986 58.392 18.36 ; 
      RECT 57.856 13.986 57.96 18.36 ; 
      RECT 57.424 13.986 57.528 18.36 ; 
      RECT 56.992 13.986 57.096 18.36 ; 
      RECT 56.56 13.986 56.664 18.36 ; 
      RECT 56.128 13.986 56.232 18.36 ; 
      RECT 55.696 13.986 55.8 18.36 ; 
      RECT 55.264 13.986 55.368 18.36 ; 
      RECT 54.832 13.986 54.936 18.36 ; 
      RECT 54.4 13.986 54.504 18.36 ; 
      RECT 53.968 13.986 54.072 18.36 ; 
      RECT 53.536 13.986 53.64 18.36 ; 
      RECT 53.104 13.986 53.208 18.36 ; 
      RECT 52.672 13.986 52.776 18.36 ; 
      RECT 52.24 13.986 52.344 18.36 ; 
      RECT 51.808 13.986 51.912 18.36 ; 
      RECT 51.376 13.986 51.48 18.36 ; 
      RECT 50.944 13.986 51.048 18.36 ; 
      RECT 50.512 13.986 50.616 18.36 ; 
      RECT 50.08 13.986 50.184 18.36 ; 
      RECT 49.648 13.986 49.752 18.36 ; 
      RECT 49.216 13.986 49.32 18.36 ; 
      RECT 48.784 13.986 48.888 18.36 ; 
      RECT 48.352 13.986 48.456 18.36 ; 
      RECT 47.92 13.986 48.024 18.36 ; 
      RECT 47.488 13.986 47.592 18.36 ; 
      RECT 47.056 13.986 47.16 18.36 ; 
      RECT 46.624 13.986 46.728 18.36 ; 
      RECT 46.192 13.986 46.296 18.36 ; 
      RECT 45.76 13.986 45.864 18.36 ; 
      RECT 45.328 13.986 45.432 18.36 ; 
      RECT 44.896 13.986 45 18.36 ; 
      RECT 44.464 13.986 44.568 18.36 ; 
      RECT 44.032 13.986 44.136 18.36 ; 
      RECT 43.6 13.986 43.704 18.36 ; 
      RECT 43.168 13.986 43.272 18.36 ; 
      RECT 42.736 13.986 42.84 18.36 ; 
      RECT 42.304 13.986 42.408 18.36 ; 
      RECT 41.872 13.986 41.976 18.36 ; 
      RECT 41.44 13.986 41.544 18.36 ; 
      RECT 41.008 13.986 41.112 18.36 ; 
      RECT 40.576 13.986 40.68 18.36 ; 
      RECT 40.144 13.986 40.248 18.36 ; 
      RECT 39.712 13.986 39.816 18.36 ; 
      RECT 39.28 13.986 39.384 18.36 ; 
      RECT 38.848 13.986 38.952 18.36 ; 
      RECT 38.416 13.986 38.52 18.36 ; 
      RECT 37.984 13.986 38.088 18.36 ; 
      RECT 37.552 13.986 37.656 18.36 ; 
      RECT 36.7 13.986 37.008 18.36 ; 
      RECT 29.128 13.986 29.436 18.36 ; 
      RECT 28.48 13.986 28.584 18.36 ; 
      RECT 28.048 13.986 28.152 18.36 ; 
      RECT 27.616 13.986 27.72 18.36 ; 
      RECT 27.184 13.986 27.288 18.36 ; 
      RECT 26.752 13.986 26.856 18.36 ; 
      RECT 26.32 13.986 26.424 18.36 ; 
      RECT 25.888 13.986 25.992 18.36 ; 
      RECT 25.456 13.986 25.56 18.36 ; 
      RECT 25.024 13.986 25.128 18.36 ; 
      RECT 24.592 13.986 24.696 18.36 ; 
      RECT 24.16 13.986 24.264 18.36 ; 
      RECT 23.728 13.986 23.832 18.36 ; 
      RECT 23.296 13.986 23.4 18.36 ; 
      RECT 22.864 13.986 22.968 18.36 ; 
      RECT 22.432 13.986 22.536 18.36 ; 
      RECT 22 13.986 22.104 18.36 ; 
      RECT 21.568 13.986 21.672 18.36 ; 
      RECT 21.136 13.986 21.24 18.36 ; 
      RECT 20.704 13.986 20.808 18.36 ; 
      RECT 20.272 13.986 20.376 18.36 ; 
      RECT 19.84 13.986 19.944 18.36 ; 
      RECT 19.408 13.986 19.512 18.36 ; 
      RECT 18.976 13.986 19.08 18.36 ; 
      RECT 18.544 13.986 18.648 18.36 ; 
      RECT 18.112 13.986 18.216 18.36 ; 
      RECT 17.68 13.986 17.784 18.36 ; 
      RECT 17.248 13.986 17.352 18.36 ; 
      RECT 16.816 13.986 16.92 18.36 ; 
      RECT 16.384 13.986 16.488 18.36 ; 
      RECT 15.952 13.986 16.056 18.36 ; 
      RECT 15.52 13.986 15.624 18.36 ; 
      RECT 15.088 13.986 15.192 18.36 ; 
      RECT 14.656 13.986 14.76 18.36 ; 
      RECT 14.224 13.986 14.328 18.36 ; 
      RECT 13.792 13.986 13.896 18.36 ; 
      RECT 13.36 13.986 13.464 18.36 ; 
      RECT 12.928 13.986 13.032 18.36 ; 
      RECT 12.496 13.986 12.6 18.36 ; 
      RECT 12.064 13.986 12.168 18.36 ; 
      RECT 11.632 13.986 11.736 18.36 ; 
      RECT 11.2 13.986 11.304 18.36 ; 
      RECT 10.768 13.986 10.872 18.36 ; 
      RECT 10.336 13.986 10.44 18.36 ; 
      RECT 9.904 13.986 10.008 18.36 ; 
      RECT 9.472 13.986 9.576 18.36 ; 
      RECT 9.04 13.986 9.144 18.36 ; 
      RECT 8.608 13.986 8.712 18.36 ; 
      RECT 8.176 13.986 8.28 18.36 ; 
      RECT 7.744 13.986 7.848 18.36 ; 
      RECT 7.312 13.986 7.416 18.36 ; 
      RECT 6.88 13.986 6.984 18.36 ; 
      RECT 6.448 13.986 6.552 18.36 ; 
      RECT 6.016 13.986 6.12 18.36 ; 
      RECT 5.584 13.986 5.688 18.36 ; 
      RECT 5.152 13.986 5.256 18.36 ; 
      RECT 4.72 13.986 4.824 18.36 ; 
      RECT 4.288 13.986 4.392 18.36 ; 
      RECT 3.856 13.986 3.96 18.36 ; 
      RECT 3.424 13.986 3.528 18.36 ; 
      RECT 2.992 13.986 3.096 18.36 ; 
      RECT 2.56 13.986 2.664 18.36 ; 
      RECT 2.128 13.986 2.232 18.36 ; 
      RECT 1.696 13.986 1.8 18.36 ; 
      RECT 1.264 13.986 1.368 18.36 ; 
      RECT 0.832 13.986 0.936 18.36 ; 
      RECT 0.02 13.986 0.36 18.36 ; 
      RECT 34.564 18.306 35.076 22.68 ; 
      RECT 34.508 20.968 35.076 22.258 ; 
      RECT 33.916 19.876 34.164 22.68 ; 
      RECT 33.86 21.114 34.164 21.728 ; 
      RECT 33.916 18.306 34.02 22.68 ; 
      RECT 33.916 18.79 34.076 19.748 ; 
      RECT 33.916 18.306 34.164 18.662 ; 
      RECT 32.728 20.108 33.552 22.68 ; 
      RECT 33.448 18.306 33.552 22.68 ; 
      RECT 32.728 21.216 33.608 22.248 ; 
      RECT 32.728 18.306 33.12 22.68 ; 
      RECT 31.06 18.306 31.392 22.68 ; 
      RECT 31.06 18.66 31.448 22.402 ; 
      RECT 65.776 18.306 66.116 22.68 ; 
      RECT 65.2 18.306 65.304 22.68 ; 
      RECT 64.768 18.306 64.872 22.68 ; 
      RECT 64.336 18.306 64.44 22.68 ; 
      RECT 63.904 18.306 64.008 22.68 ; 
      RECT 63.472 18.306 63.576 22.68 ; 
      RECT 63.04 18.306 63.144 22.68 ; 
      RECT 62.608 18.306 62.712 22.68 ; 
      RECT 62.176 18.306 62.28 22.68 ; 
      RECT 61.744 18.306 61.848 22.68 ; 
      RECT 61.312 18.306 61.416 22.68 ; 
      RECT 60.88 18.306 60.984 22.68 ; 
      RECT 60.448 18.306 60.552 22.68 ; 
      RECT 60.016 18.306 60.12 22.68 ; 
      RECT 59.584 18.306 59.688 22.68 ; 
      RECT 59.152 18.306 59.256 22.68 ; 
      RECT 58.72 18.306 58.824 22.68 ; 
      RECT 58.288 18.306 58.392 22.68 ; 
      RECT 57.856 18.306 57.96 22.68 ; 
      RECT 57.424 18.306 57.528 22.68 ; 
      RECT 56.992 18.306 57.096 22.68 ; 
      RECT 56.56 18.306 56.664 22.68 ; 
      RECT 56.128 18.306 56.232 22.68 ; 
      RECT 55.696 18.306 55.8 22.68 ; 
      RECT 55.264 18.306 55.368 22.68 ; 
      RECT 54.832 18.306 54.936 22.68 ; 
      RECT 54.4 18.306 54.504 22.68 ; 
      RECT 53.968 18.306 54.072 22.68 ; 
      RECT 53.536 18.306 53.64 22.68 ; 
      RECT 53.104 18.306 53.208 22.68 ; 
      RECT 52.672 18.306 52.776 22.68 ; 
      RECT 52.24 18.306 52.344 22.68 ; 
      RECT 51.808 18.306 51.912 22.68 ; 
      RECT 51.376 18.306 51.48 22.68 ; 
      RECT 50.944 18.306 51.048 22.68 ; 
      RECT 50.512 18.306 50.616 22.68 ; 
      RECT 50.08 18.306 50.184 22.68 ; 
      RECT 49.648 18.306 49.752 22.68 ; 
      RECT 49.216 18.306 49.32 22.68 ; 
      RECT 48.784 18.306 48.888 22.68 ; 
      RECT 48.352 18.306 48.456 22.68 ; 
      RECT 47.92 18.306 48.024 22.68 ; 
      RECT 47.488 18.306 47.592 22.68 ; 
      RECT 47.056 18.306 47.16 22.68 ; 
      RECT 46.624 18.306 46.728 22.68 ; 
      RECT 46.192 18.306 46.296 22.68 ; 
      RECT 45.76 18.306 45.864 22.68 ; 
      RECT 45.328 18.306 45.432 22.68 ; 
      RECT 44.896 18.306 45 22.68 ; 
      RECT 44.464 18.306 44.568 22.68 ; 
      RECT 44.032 18.306 44.136 22.68 ; 
      RECT 43.6 18.306 43.704 22.68 ; 
      RECT 43.168 18.306 43.272 22.68 ; 
      RECT 42.736 18.306 42.84 22.68 ; 
      RECT 42.304 18.306 42.408 22.68 ; 
      RECT 41.872 18.306 41.976 22.68 ; 
      RECT 41.44 18.306 41.544 22.68 ; 
      RECT 41.008 18.306 41.112 22.68 ; 
      RECT 40.576 18.306 40.68 22.68 ; 
      RECT 40.144 18.306 40.248 22.68 ; 
      RECT 39.712 18.306 39.816 22.68 ; 
      RECT 39.28 18.306 39.384 22.68 ; 
      RECT 38.848 18.306 38.952 22.68 ; 
      RECT 38.416 18.306 38.52 22.68 ; 
      RECT 37.984 18.306 38.088 22.68 ; 
      RECT 37.552 18.306 37.656 22.68 ; 
      RECT 36.7 18.306 37.008 22.68 ; 
      RECT 29.128 18.306 29.436 22.68 ; 
      RECT 28.48 18.306 28.584 22.68 ; 
      RECT 28.048 18.306 28.152 22.68 ; 
      RECT 27.616 18.306 27.72 22.68 ; 
      RECT 27.184 18.306 27.288 22.68 ; 
      RECT 26.752 18.306 26.856 22.68 ; 
      RECT 26.32 18.306 26.424 22.68 ; 
      RECT 25.888 18.306 25.992 22.68 ; 
      RECT 25.456 18.306 25.56 22.68 ; 
      RECT 25.024 18.306 25.128 22.68 ; 
      RECT 24.592 18.306 24.696 22.68 ; 
      RECT 24.16 18.306 24.264 22.68 ; 
      RECT 23.728 18.306 23.832 22.68 ; 
      RECT 23.296 18.306 23.4 22.68 ; 
      RECT 22.864 18.306 22.968 22.68 ; 
      RECT 22.432 18.306 22.536 22.68 ; 
      RECT 22 18.306 22.104 22.68 ; 
      RECT 21.568 18.306 21.672 22.68 ; 
      RECT 21.136 18.306 21.24 22.68 ; 
      RECT 20.704 18.306 20.808 22.68 ; 
      RECT 20.272 18.306 20.376 22.68 ; 
      RECT 19.84 18.306 19.944 22.68 ; 
      RECT 19.408 18.306 19.512 22.68 ; 
      RECT 18.976 18.306 19.08 22.68 ; 
      RECT 18.544 18.306 18.648 22.68 ; 
      RECT 18.112 18.306 18.216 22.68 ; 
      RECT 17.68 18.306 17.784 22.68 ; 
      RECT 17.248 18.306 17.352 22.68 ; 
      RECT 16.816 18.306 16.92 22.68 ; 
      RECT 16.384 18.306 16.488 22.68 ; 
      RECT 15.952 18.306 16.056 22.68 ; 
      RECT 15.52 18.306 15.624 22.68 ; 
      RECT 15.088 18.306 15.192 22.68 ; 
      RECT 14.656 18.306 14.76 22.68 ; 
      RECT 14.224 18.306 14.328 22.68 ; 
      RECT 13.792 18.306 13.896 22.68 ; 
      RECT 13.36 18.306 13.464 22.68 ; 
      RECT 12.928 18.306 13.032 22.68 ; 
      RECT 12.496 18.306 12.6 22.68 ; 
      RECT 12.064 18.306 12.168 22.68 ; 
      RECT 11.632 18.306 11.736 22.68 ; 
      RECT 11.2 18.306 11.304 22.68 ; 
      RECT 10.768 18.306 10.872 22.68 ; 
      RECT 10.336 18.306 10.44 22.68 ; 
      RECT 9.904 18.306 10.008 22.68 ; 
      RECT 9.472 18.306 9.576 22.68 ; 
      RECT 9.04 18.306 9.144 22.68 ; 
      RECT 8.608 18.306 8.712 22.68 ; 
      RECT 8.176 18.306 8.28 22.68 ; 
      RECT 7.744 18.306 7.848 22.68 ; 
      RECT 7.312 18.306 7.416 22.68 ; 
      RECT 6.88 18.306 6.984 22.68 ; 
      RECT 6.448 18.306 6.552 22.68 ; 
      RECT 6.016 18.306 6.12 22.68 ; 
      RECT 5.584 18.306 5.688 22.68 ; 
      RECT 5.152 18.306 5.256 22.68 ; 
      RECT 4.72 18.306 4.824 22.68 ; 
      RECT 4.288 18.306 4.392 22.68 ; 
      RECT 3.856 18.306 3.96 22.68 ; 
      RECT 3.424 18.306 3.528 22.68 ; 
      RECT 2.992 18.306 3.096 22.68 ; 
      RECT 2.56 18.306 2.664 22.68 ; 
      RECT 2.128 18.306 2.232 22.68 ; 
      RECT 1.696 18.306 1.8 22.68 ; 
      RECT 1.264 18.306 1.368 22.68 ; 
      RECT 0.832 18.306 0.936 22.68 ; 
      RECT 0.02 18.306 0.36 22.68 ; 
      RECT 34.564 22.626 35.076 27 ; 
      RECT 34.508 25.288 35.076 26.578 ; 
      RECT 33.916 24.196 34.164 27 ; 
      RECT 33.86 25.434 34.164 26.048 ; 
      RECT 33.916 22.626 34.02 27 ; 
      RECT 33.916 23.11 34.076 24.068 ; 
      RECT 33.916 22.626 34.164 22.982 ; 
      RECT 32.728 24.428 33.552 27 ; 
      RECT 33.448 22.626 33.552 27 ; 
      RECT 32.728 25.536 33.608 26.568 ; 
      RECT 32.728 22.626 33.12 27 ; 
      RECT 31.06 22.626 31.392 27 ; 
      RECT 31.06 22.98 31.448 26.722 ; 
      RECT 65.776 22.626 66.116 27 ; 
      RECT 65.2 22.626 65.304 27 ; 
      RECT 64.768 22.626 64.872 27 ; 
      RECT 64.336 22.626 64.44 27 ; 
      RECT 63.904 22.626 64.008 27 ; 
      RECT 63.472 22.626 63.576 27 ; 
      RECT 63.04 22.626 63.144 27 ; 
      RECT 62.608 22.626 62.712 27 ; 
      RECT 62.176 22.626 62.28 27 ; 
      RECT 61.744 22.626 61.848 27 ; 
      RECT 61.312 22.626 61.416 27 ; 
      RECT 60.88 22.626 60.984 27 ; 
      RECT 60.448 22.626 60.552 27 ; 
      RECT 60.016 22.626 60.12 27 ; 
      RECT 59.584 22.626 59.688 27 ; 
      RECT 59.152 22.626 59.256 27 ; 
      RECT 58.72 22.626 58.824 27 ; 
      RECT 58.288 22.626 58.392 27 ; 
      RECT 57.856 22.626 57.96 27 ; 
      RECT 57.424 22.626 57.528 27 ; 
      RECT 56.992 22.626 57.096 27 ; 
      RECT 56.56 22.626 56.664 27 ; 
      RECT 56.128 22.626 56.232 27 ; 
      RECT 55.696 22.626 55.8 27 ; 
      RECT 55.264 22.626 55.368 27 ; 
      RECT 54.832 22.626 54.936 27 ; 
      RECT 54.4 22.626 54.504 27 ; 
      RECT 53.968 22.626 54.072 27 ; 
      RECT 53.536 22.626 53.64 27 ; 
      RECT 53.104 22.626 53.208 27 ; 
      RECT 52.672 22.626 52.776 27 ; 
      RECT 52.24 22.626 52.344 27 ; 
      RECT 51.808 22.626 51.912 27 ; 
      RECT 51.376 22.626 51.48 27 ; 
      RECT 50.944 22.626 51.048 27 ; 
      RECT 50.512 22.626 50.616 27 ; 
      RECT 50.08 22.626 50.184 27 ; 
      RECT 49.648 22.626 49.752 27 ; 
      RECT 49.216 22.626 49.32 27 ; 
      RECT 48.784 22.626 48.888 27 ; 
      RECT 48.352 22.626 48.456 27 ; 
      RECT 47.92 22.626 48.024 27 ; 
      RECT 47.488 22.626 47.592 27 ; 
      RECT 47.056 22.626 47.16 27 ; 
      RECT 46.624 22.626 46.728 27 ; 
      RECT 46.192 22.626 46.296 27 ; 
      RECT 45.76 22.626 45.864 27 ; 
      RECT 45.328 22.626 45.432 27 ; 
      RECT 44.896 22.626 45 27 ; 
      RECT 44.464 22.626 44.568 27 ; 
      RECT 44.032 22.626 44.136 27 ; 
      RECT 43.6 22.626 43.704 27 ; 
      RECT 43.168 22.626 43.272 27 ; 
      RECT 42.736 22.626 42.84 27 ; 
      RECT 42.304 22.626 42.408 27 ; 
      RECT 41.872 22.626 41.976 27 ; 
      RECT 41.44 22.626 41.544 27 ; 
      RECT 41.008 22.626 41.112 27 ; 
      RECT 40.576 22.626 40.68 27 ; 
      RECT 40.144 22.626 40.248 27 ; 
      RECT 39.712 22.626 39.816 27 ; 
      RECT 39.28 22.626 39.384 27 ; 
      RECT 38.848 22.626 38.952 27 ; 
      RECT 38.416 22.626 38.52 27 ; 
      RECT 37.984 22.626 38.088 27 ; 
      RECT 37.552 22.626 37.656 27 ; 
      RECT 36.7 22.626 37.008 27 ; 
      RECT 29.128 22.626 29.436 27 ; 
      RECT 28.48 22.626 28.584 27 ; 
      RECT 28.048 22.626 28.152 27 ; 
      RECT 27.616 22.626 27.72 27 ; 
      RECT 27.184 22.626 27.288 27 ; 
      RECT 26.752 22.626 26.856 27 ; 
      RECT 26.32 22.626 26.424 27 ; 
      RECT 25.888 22.626 25.992 27 ; 
      RECT 25.456 22.626 25.56 27 ; 
      RECT 25.024 22.626 25.128 27 ; 
      RECT 24.592 22.626 24.696 27 ; 
      RECT 24.16 22.626 24.264 27 ; 
      RECT 23.728 22.626 23.832 27 ; 
      RECT 23.296 22.626 23.4 27 ; 
      RECT 22.864 22.626 22.968 27 ; 
      RECT 22.432 22.626 22.536 27 ; 
      RECT 22 22.626 22.104 27 ; 
      RECT 21.568 22.626 21.672 27 ; 
      RECT 21.136 22.626 21.24 27 ; 
      RECT 20.704 22.626 20.808 27 ; 
      RECT 20.272 22.626 20.376 27 ; 
      RECT 19.84 22.626 19.944 27 ; 
      RECT 19.408 22.626 19.512 27 ; 
      RECT 18.976 22.626 19.08 27 ; 
      RECT 18.544 22.626 18.648 27 ; 
      RECT 18.112 22.626 18.216 27 ; 
      RECT 17.68 22.626 17.784 27 ; 
      RECT 17.248 22.626 17.352 27 ; 
      RECT 16.816 22.626 16.92 27 ; 
      RECT 16.384 22.626 16.488 27 ; 
      RECT 15.952 22.626 16.056 27 ; 
      RECT 15.52 22.626 15.624 27 ; 
      RECT 15.088 22.626 15.192 27 ; 
      RECT 14.656 22.626 14.76 27 ; 
      RECT 14.224 22.626 14.328 27 ; 
      RECT 13.792 22.626 13.896 27 ; 
      RECT 13.36 22.626 13.464 27 ; 
      RECT 12.928 22.626 13.032 27 ; 
      RECT 12.496 22.626 12.6 27 ; 
      RECT 12.064 22.626 12.168 27 ; 
      RECT 11.632 22.626 11.736 27 ; 
      RECT 11.2 22.626 11.304 27 ; 
      RECT 10.768 22.626 10.872 27 ; 
      RECT 10.336 22.626 10.44 27 ; 
      RECT 9.904 22.626 10.008 27 ; 
      RECT 9.472 22.626 9.576 27 ; 
      RECT 9.04 22.626 9.144 27 ; 
      RECT 8.608 22.626 8.712 27 ; 
      RECT 8.176 22.626 8.28 27 ; 
      RECT 7.744 22.626 7.848 27 ; 
      RECT 7.312 22.626 7.416 27 ; 
      RECT 6.88 22.626 6.984 27 ; 
      RECT 6.448 22.626 6.552 27 ; 
      RECT 6.016 22.626 6.12 27 ; 
      RECT 5.584 22.626 5.688 27 ; 
      RECT 5.152 22.626 5.256 27 ; 
      RECT 4.72 22.626 4.824 27 ; 
      RECT 4.288 22.626 4.392 27 ; 
      RECT 3.856 22.626 3.96 27 ; 
      RECT 3.424 22.626 3.528 27 ; 
      RECT 2.992 22.626 3.096 27 ; 
      RECT 2.56 22.626 2.664 27 ; 
      RECT 2.128 22.626 2.232 27 ; 
      RECT 1.696 22.626 1.8 27 ; 
      RECT 1.264 22.626 1.368 27 ; 
      RECT 0.832 22.626 0.936 27 ; 
      RECT 0.02 22.626 0.36 27 ; 
      RECT 34.564 26.946 35.076 31.32 ; 
      RECT 34.508 29.608 35.076 30.898 ; 
      RECT 33.916 28.516 34.164 31.32 ; 
      RECT 33.86 29.754 34.164 30.368 ; 
      RECT 33.916 26.946 34.02 31.32 ; 
      RECT 33.916 27.43 34.076 28.388 ; 
      RECT 33.916 26.946 34.164 27.302 ; 
      RECT 32.728 28.748 33.552 31.32 ; 
      RECT 33.448 26.946 33.552 31.32 ; 
      RECT 32.728 29.856 33.608 30.888 ; 
      RECT 32.728 26.946 33.12 31.32 ; 
      RECT 31.06 26.946 31.392 31.32 ; 
      RECT 31.06 27.3 31.448 31.042 ; 
      RECT 65.776 26.946 66.116 31.32 ; 
      RECT 65.2 26.946 65.304 31.32 ; 
      RECT 64.768 26.946 64.872 31.32 ; 
      RECT 64.336 26.946 64.44 31.32 ; 
      RECT 63.904 26.946 64.008 31.32 ; 
      RECT 63.472 26.946 63.576 31.32 ; 
      RECT 63.04 26.946 63.144 31.32 ; 
      RECT 62.608 26.946 62.712 31.32 ; 
      RECT 62.176 26.946 62.28 31.32 ; 
      RECT 61.744 26.946 61.848 31.32 ; 
      RECT 61.312 26.946 61.416 31.32 ; 
      RECT 60.88 26.946 60.984 31.32 ; 
      RECT 60.448 26.946 60.552 31.32 ; 
      RECT 60.016 26.946 60.12 31.32 ; 
      RECT 59.584 26.946 59.688 31.32 ; 
      RECT 59.152 26.946 59.256 31.32 ; 
      RECT 58.72 26.946 58.824 31.32 ; 
      RECT 58.288 26.946 58.392 31.32 ; 
      RECT 57.856 26.946 57.96 31.32 ; 
      RECT 57.424 26.946 57.528 31.32 ; 
      RECT 56.992 26.946 57.096 31.32 ; 
      RECT 56.56 26.946 56.664 31.32 ; 
      RECT 56.128 26.946 56.232 31.32 ; 
      RECT 55.696 26.946 55.8 31.32 ; 
      RECT 55.264 26.946 55.368 31.32 ; 
      RECT 54.832 26.946 54.936 31.32 ; 
      RECT 54.4 26.946 54.504 31.32 ; 
      RECT 53.968 26.946 54.072 31.32 ; 
      RECT 53.536 26.946 53.64 31.32 ; 
      RECT 53.104 26.946 53.208 31.32 ; 
      RECT 52.672 26.946 52.776 31.32 ; 
      RECT 52.24 26.946 52.344 31.32 ; 
      RECT 51.808 26.946 51.912 31.32 ; 
      RECT 51.376 26.946 51.48 31.32 ; 
      RECT 50.944 26.946 51.048 31.32 ; 
      RECT 50.512 26.946 50.616 31.32 ; 
      RECT 50.08 26.946 50.184 31.32 ; 
      RECT 49.648 26.946 49.752 31.32 ; 
      RECT 49.216 26.946 49.32 31.32 ; 
      RECT 48.784 26.946 48.888 31.32 ; 
      RECT 48.352 26.946 48.456 31.32 ; 
      RECT 47.92 26.946 48.024 31.32 ; 
      RECT 47.488 26.946 47.592 31.32 ; 
      RECT 47.056 26.946 47.16 31.32 ; 
      RECT 46.624 26.946 46.728 31.32 ; 
      RECT 46.192 26.946 46.296 31.32 ; 
      RECT 45.76 26.946 45.864 31.32 ; 
      RECT 45.328 26.946 45.432 31.32 ; 
      RECT 44.896 26.946 45 31.32 ; 
      RECT 44.464 26.946 44.568 31.32 ; 
      RECT 44.032 26.946 44.136 31.32 ; 
      RECT 43.6 26.946 43.704 31.32 ; 
      RECT 43.168 26.946 43.272 31.32 ; 
      RECT 42.736 26.946 42.84 31.32 ; 
      RECT 42.304 26.946 42.408 31.32 ; 
      RECT 41.872 26.946 41.976 31.32 ; 
      RECT 41.44 26.946 41.544 31.32 ; 
      RECT 41.008 26.946 41.112 31.32 ; 
      RECT 40.576 26.946 40.68 31.32 ; 
      RECT 40.144 26.946 40.248 31.32 ; 
      RECT 39.712 26.946 39.816 31.32 ; 
      RECT 39.28 26.946 39.384 31.32 ; 
      RECT 38.848 26.946 38.952 31.32 ; 
      RECT 38.416 26.946 38.52 31.32 ; 
      RECT 37.984 26.946 38.088 31.32 ; 
      RECT 37.552 26.946 37.656 31.32 ; 
      RECT 36.7 26.946 37.008 31.32 ; 
      RECT 29.128 26.946 29.436 31.32 ; 
      RECT 28.48 26.946 28.584 31.32 ; 
      RECT 28.048 26.946 28.152 31.32 ; 
      RECT 27.616 26.946 27.72 31.32 ; 
      RECT 27.184 26.946 27.288 31.32 ; 
      RECT 26.752 26.946 26.856 31.32 ; 
      RECT 26.32 26.946 26.424 31.32 ; 
      RECT 25.888 26.946 25.992 31.32 ; 
      RECT 25.456 26.946 25.56 31.32 ; 
      RECT 25.024 26.946 25.128 31.32 ; 
      RECT 24.592 26.946 24.696 31.32 ; 
      RECT 24.16 26.946 24.264 31.32 ; 
      RECT 23.728 26.946 23.832 31.32 ; 
      RECT 23.296 26.946 23.4 31.32 ; 
      RECT 22.864 26.946 22.968 31.32 ; 
      RECT 22.432 26.946 22.536 31.32 ; 
      RECT 22 26.946 22.104 31.32 ; 
      RECT 21.568 26.946 21.672 31.32 ; 
      RECT 21.136 26.946 21.24 31.32 ; 
      RECT 20.704 26.946 20.808 31.32 ; 
      RECT 20.272 26.946 20.376 31.32 ; 
      RECT 19.84 26.946 19.944 31.32 ; 
      RECT 19.408 26.946 19.512 31.32 ; 
      RECT 18.976 26.946 19.08 31.32 ; 
      RECT 18.544 26.946 18.648 31.32 ; 
      RECT 18.112 26.946 18.216 31.32 ; 
      RECT 17.68 26.946 17.784 31.32 ; 
      RECT 17.248 26.946 17.352 31.32 ; 
      RECT 16.816 26.946 16.92 31.32 ; 
      RECT 16.384 26.946 16.488 31.32 ; 
      RECT 15.952 26.946 16.056 31.32 ; 
      RECT 15.52 26.946 15.624 31.32 ; 
      RECT 15.088 26.946 15.192 31.32 ; 
      RECT 14.656 26.946 14.76 31.32 ; 
      RECT 14.224 26.946 14.328 31.32 ; 
      RECT 13.792 26.946 13.896 31.32 ; 
      RECT 13.36 26.946 13.464 31.32 ; 
      RECT 12.928 26.946 13.032 31.32 ; 
      RECT 12.496 26.946 12.6 31.32 ; 
      RECT 12.064 26.946 12.168 31.32 ; 
      RECT 11.632 26.946 11.736 31.32 ; 
      RECT 11.2 26.946 11.304 31.32 ; 
      RECT 10.768 26.946 10.872 31.32 ; 
      RECT 10.336 26.946 10.44 31.32 ; 
      RECT 9.904 26.946 10.008 31.32 ; 
      RECT 9.472 26.946 9.576 31.32 ; 
      RECT 9.04 26.946 9.144 31.32 ; 
      RECT 8.608 26.946 8.712 31.32 ; 
      RECT 8.176 26.946 8.28 31.32 ; 
      RECT 7.744 26.946 7.848 31.32 ; 
      RECT 7.312 26.946 7.416 31.32 ; 
      RECT 6.88 26.946 6.984 31.32 ; 
      RECT 6.448 26.946 6.552 31.32 ; 
      RECT 6.016 26.946 6.12 31.32 ; 
      RECT 5.584 26.946 5.688 31.32 ; 
      RECT 5.152 26.946 5.256 31.32 ; 
      RECT 4.72 26.946 4.824 31.32 ; 
      RECT 4.288 26.946 4.392 31.32 ; 
      RECT 3.856 26.946 3.96 31.32 ; 
      RECT 3.424 26.946 3.528 31.32 ; 
      RECT 2.992 26.946 3.096 31.32 ; 
      RECT 2.56 26.946 2.664 31.32 ; 
      RECT 2.128 26.946 2.232 31.32 ; 
      RECT 1.696 26.946 1.8 31.32 ; 
      RECT 1.264 26.946 1.368 31.32 ; 
      RECT 0.832 26.946 0.936 31.32 ; 
      RECT 0.02 26.946 0.36 31.32 ; 
      RECT 34.564 31.266 35.076 35.64 ; 
      RECT 34.508 33.928 35.076 35.218 ; 
      RECT 33.916 32.836 34.164 35.64 ; 
      RECT 33.86 34.074 34.164 34.688 ; 
      RECT 33.916 31.266 34.02 35.64 ; 
      RECT 33.916 31.75 34.076 32.708 ; 
      RECT 33.916 31.266 34.164 31.622 ; 
      RECT 32.728 33.068 33.552 35.64 ; 
      RECT 33.448 31.266 33.552 35.64 ; 
      RECT 32.728 34.176 33.608 35.208 ; 
      RECT 32.728 31.266 33.12 35.64 ; 
      RECT 31.06 31.266 31.392 35.64 ; 
      RECT 31.06 31.62 31.448 35.362 ; 
      RECT 65.776 31.266 66.116 35.64 ; 
      RECT 65.2 31.266 65.304 35.64 ; 
      RECT 64.768 31.266 64.872 35.64 ; 
      RECT 64.336 31.266 64.44 35.64 ; 
      RECT 63.904 31.266 64.008 35.64 ; 
      RECT 63.472 31.266 63.576 35.64 ; 
      RECT 63.04 31.266 63.144 35.64 ; 
      RECT 62.608 31.266 62.712 35.64 ; 
      RECT 62.176 31.266 62.28 35.64 ; 
      RECT 61.744 31.266 61.848 35.64 ; 
      RECT 61.312 31.266 61.416 35.64 ; 
      RECT 60.88 31.266 60.984 35.64 ; 
      RECT 60.448 31.266 60.552 35.64 ; 
      RECT 60.016 31.266 60.12 35.64 ; 
      RECT 59.584 31.266 59.688 35.64 ; 
      RECT 59.152 31.266 59.256 35.64 ; 
      RECT 58.72 31.266 58.824 35.64 ; 
      RECT 58.288 31.266 58.392 35.64 ; 
      RECT 57.856 31.266 57.96 35.64 ; 
      RECT 57.424 31.266 57.528 35.64 ; 
      RECT 56.992 31.266 57.096 35.64 ; 
      RECT 56.56 31.266 56.664 35.64 ; 
      RECT 56.128 31.266 56.232 35.64 ; 
      RECT 55.696 31.266 55.8 35.64 ; 
      RECT 55.264 31.266 55.368 35.64 ; 
      RECT 54.832 31.266 54.936 35.64 ; 
      RECT 54.4 31.266 54.504 35.64 ; 
      RECT 53.968 31.266 54.072 35.64 ; 
      RECT 53.536 31.266 53.64 35.64 ; 
      RECT 53.104 31.266 53.208 35.64 ; 
      RECT 52.672 31.266 52.776 35.64 ; 
      RECT 52.24 31.266 52.344 35.64 ; 
      RECT 51.808 31.266 51.912 35.64 ; 
      RECT 51.376 31.266 51.48 35.64 ; 
      RECT 50.944 31.266 51.048 35.64 ; 
      RECT 50.512 31.266 50.616 35.64 ; 
      RECT 50.08 31.266 50.184 35.64 ; 
      RECT 49.648 31.266 49.752 35.64 ; 
      RECT 49.216 31.266 49.32 35.64 ; 
      RECT 48.784 31.266 48.888 35.64 ; 
      RECT 48.352 31.266 48.456 35.64 ; 
      RECT 47.92 31.266 48.024 35.64 ; 
      RECT 47.488 31.266 47.592 35.64 ; 
      RECT 47.056 31.266 47.16 35.64 ; 
      RECT 46.624 31.266 46.728 35.64 ; 
      RECT 46.192 31.266 46.296 35.64 ; 
      RECT 45.76 31.266 45.864 35.64 ; 
      RECT 45.328 31.266 45.432 35.64 ; 
      RECT 44.896 31.266 45 35.64 ; 
      RECT 44.464 31.266 44.568 35.64 ; 
      RECT 44.032 31.266 44.136 35.64 ; 
      RECT 43.6 31.266 43.704 35.64 ; 
      RECT 43.168 31.266 43.272 35.64 ; 
      RECT 42.736 31.266 42.84 35.64 ; 
      RECT 42.304 31.266 42.408 35.64 ; 
      RECT 41.872 31.266 41.976 35.64 ; 
      RECT 41.44 31.266 41.544 35.64 ; 
      RECT 41.008 31.266 41.112 35.64 ; 
      RECT 40.576 31.266 40.68 35.64 ; 
      RECT 40.144 31.266 40.248 35.64 ; 
      RECT 39.712 31.266 39.816 35.64 ; 
      RECT 39.28 31.266 39.384 35.64 ; 
      RECT 38.848 31.266 38.952 35.64 ; 
      RECT 38.416 31.266 38.52 35.64 ; 
      RECT 37.984 31.266 38.088 35.64 ; 
      RECT 37.552 31.266 37.656 35.64 ; 
      RECT 36.7 31.266 37.008 35.64 ; 
      RECT 29.128 31.266 29.436 35.64 ; 
      RECT 28.48 31.266 28.584 35.64 ; 
      RECT 28.048 31.266 28.152 35.64 ; 
      RECT 27.616 31.266 27.72 35.64 ; 
      RECT 27.184 31.266 27.288 35.64 ; 
      RECT 26.752 31.266 26.856 35.64 ; 
      RECT 26.32 31.266 26.424 35.64 ; 
      RECT 25.888 31.266 25.992 35.64 ; 
      RECT 25.456 31.266 25.56 35.64 ; 
      RECT 25.024 31.266 25.128 35.64 ; 
      RECT 24.592 31.266 24.696 35.64 ; 
      RECT 24.16 31.266 24.264 35.64 ; 
      RECT 23.728 31.266 23.832 35.64 ; 
      RECT 23.296 31.266 23.4 35.64 ; 
      RECT 22.864 31.266 22.968 35.64 ; 
      RECT 22.432 31.266 22.536 35.64 ; 
      RECT 22 31.266 22.104 35.64 ; 
      RECT 21.568 31.266 21.672 35.64 ; 
      RECT 21.136 31.266 21.24 35.64 ; 
      RECT 20.704 31.266 20.808 35.64 ; 
      RECT 20.272 31.266 20.376 35.64 ; 
      RECT 19.84 31.266 19.944 35.64 ; 
      RECT 19.408 31.266 19.512 35.64 ; 
      RECT 18.976 31.266 19.08 35.64 ; 
      RECT 18.544 31.266 18.648 35.64 ; 
      RECT 18.112 31.266 18.216 35.64 ; 
      RECT 17.68 31.266 17.784 35.64 ; 
      RECT 17.248 31.266 17.352 35.64 ; 
      RECT 16.816 31.266 16.92 35.64 ; 
      RECT 16.384 31.266 16.488 35.64 ; 
      RECT 15.952 31.266 16.056 35.64 ; 
      RECT 15.52 31.266 15.624 35.64 ; 
      RECT 15.088 31.266 15.192 35.64 ; 
      RECT 14.656 31.266 14.76 35.64 ; 
      RECT 14.224 31.266 14.328 35.64 ; 
      RECT 13.792 31.266 13.896 35.64 ; 
      RECT 13.36 31.266 13.464 35.64 ; 
      RECT 12.928 31.266 13.032 35.64 ; 
      RECT 12.496 31.266 12.6 35.64 ; 
      RECT 12.064 31.266 12.168 35.64 ; 
      RECT 11.632 31.266 11.736 35.64 ; 
      RECT 11.2 31.266 11.304 35.64 ; 
      RECT 10.768 31.266 10.872 35.64 ; 
      RECT 10.336 31.266 10.44 35.64 ; 
      RECT 9.904 31.266 10.008 35.64 ; 
      RECT 9.472 31.266 9.576 35.64 ; 
      RECT 9.04 31.266 9.144 35.64 ; 
      RECT 8.608 31.266 8.712 35.64 ; 
      RECT 8.176 31.266 8.28 35.64 ; 
      RECT 7.744 31.266 7.848 35.64 ; 
      RECT 7.312 31.266 7.416 35.64 ; 
      RECT 6.88 31.266 6.984 35.64 ; 
      RECT 6.448 31.266 6.552 35.64 ; 
      RECT 6.016 31.266 6.12 35.64 ; 
      RECT 5.584 31.266 5.688 35.64 ; 
      RECT 5.152 31.266 5.256 35.64 ; 
      RECT 4.72 31.266 4.824 35.64 ; 
      RECT 4.288 31.266 4.392 35.64 ; 
      RECT 3.856 31.266 3.96 35.64 ; 
      RECT 3.424 31.266 3.528 35.64 ; 
      RECT 2.992 31.266 3.096 35.64 ; 
      RECT 2.56 31.266 2.664 35.64 ; 
      RECT 2.128 31.266 2.232 35.64 ; 
      RECT 1.696 31.266 1.8 35.64 ; 
      RECT 1.264 31.266 1.368 35.64 ; 
      RECT 0.832 31.266 0.936 35.64 ; 
      RECT 0.02 31.266 0.36 35.64 ; 
      RECT 34.564 35.586 35.076 39.96 ; 
      RECT 34.508 38.248 35.076 39.538 ; 
      RECT 33.916 37.156 34.164 39.96 ; 
      RECT 33.86 38.394 34.164 39.008 ; 
      RECT 33.916 35.586 34.02 39.96 ; 
      RECT 33.916 36.07 34.076 37.028 ; 
      RECT 33.916 35.586 34.164 35.942 ; 
      RECT 32.728 37.388 33.552 39.96 ; 
      RECT 33.448 35.586 33.552 39.96 ; 
      RECT 32.728 38.496 33.608 39.528 ; 
      RECT 32.728 35.586 33.12 39.96 ; 
      RECT 31.06 35.586 31.392 39.96 ; 
      RECT 31.06 35.94 31.448 39.682 ; 
      RECT 65.776 35.586 66.116 39.96 ; 
      RECT 65.2 35.586 65.304 39.96 ; 
      RECT 64.768 35.586 64.872 39.96 ; 
      RECT 64.336 35.586 64.44 39.96 ; 
      RECT 63.904 35.586 64.008 39.96 ; 
      RECT 63.472 35.586 63.576 39.96 ; 
      RECT 63.04 35.586 63.144 39.96 ; 
      RECT 62.608 35.586 62.712 39.96 ; 
      RECT 62.176 35.586 62.28 39.96 ; 
      RECT 61.744 35.586 61.848 39.96 ; 
      RECT 61.312 35.586 61.416 39.96 ; 
      RECT 60.88 35.586 60.984 39.96 ; 
      RECT 60.448 35.586 60.552 39.96 ; 
      RECT 60.016 35.586 60.12 39.96 ; 
      RECT 59.584 35.586 59.688 39.96 ; 
      RECT 59.152 35.586 59.256 39.96 ; 
      RECT 58.72 35.586 58.824 39.96 ; 
      RECT 58.288 35.586 58.392 39.96 ; 
      RECT 57.856 35.586 57.96 39.96 ; 
      RECT 57.424 35.586 57.528 39.96 ; 
      RECT 56.992 35.586 57.096 39.96 ; 
      RECT 56.56 35.586 56.664 39.96 ; 
      RECT 56.128 35.586 56.232 39.96 ; 
      RECT 55.696 35.586 55.8 39.96 ; 
      RECT 55.264 35.586 55.368 39.96 ; 
      RECT 54.832 35.586 54.936 39.96 ; 
      RECT 54.4 35.586 54.504 39.96 ; 
      RECT 53.968 35.586 54.072 39.96 ; 
      RECT 53.536 35.586 53.64 39.96 ; 
      RECT 53.104 35.586 53.208 39.96 ; 
      RECT 52.672 35.586 52.776 39.96 ; 
      RECT 52.24 35.586 52.344 39.96 ; 
      RECT 51.808 35.586 51.912 39.96 ; 
      RECT 51.376 35.586 51.48 39.96 ; 
      RECT 50.944 35.586 51.048 39.96 ; 
      RECT 50.512 35.586 50.616 39.96 ; 
      RECT 50.08 35.586 50.184 39.96 ; 
      RECT 49.648 35.586 49.752 39.96 ; 
      RECT 49.216 35.586 49.32 39.96 ; 
      RECT 48.784 35.586 48.888 39.96 ; 
      RECT 48.352 35.586 48.456 39.96 ; 
      RECT 47.92 35.586 48.024 39.96 ; 
      RECT 47.488 35.586 47.592 39.96 ; 
      RECT 47.056 35.586 47.16 39.96 ; 
      RECT 46.624 35.586 46.728 39.96 ; 
      RECT 46.192 35.586 46.296 39.96 ; 
      RECT 45.76 35.586 45.864 39.96 ; 
      RECT 45.328 35.586 45.432 39.96 ; 
      RECT 44.896 35.586 45 39.96 ; 
      RECT 44.464 35.586 44.568 39.96 ; 
      RECT 44.032 35.586 44.136 39.96 ; 
      RECT 43.6 35.586 43.704 39.96 ; 
      RECT 43.168 35.586 43.272 39.96 ; 
      RECT 42.736 35.586 42.84 39.96 ; 
      RECT 42.304 35.586 42.408 39.96 ; 
      RECT 41.872 35.586 41.976 39.96 ; 
      RECT 41.44 35.586 41.544 39.96 ; 
      RECT 41.008 35.586 41.112 39.96 ; 
      RECT 40.576 35.586 40.68 39.96 ; 
      RECT 40.144 35.586 40.248 39.96 ; 
      RECT 39.712 35.586 39.816 39.96 ; 
      RECT 39.28 35.586 39.384 39.96 ; 
      RECT 38.848 35.586 38.952 39.96 ; 
      RECT 38.416 35.586 38.52 39.96 ; 
      RECT 37.984 35.586 38.088 39.96 ; 
      RECT 37.552 35.586 37.656 39.96 ; 
      RECT 36.7 35.586 37.008 39.96 ; 
      RECT 29.128 35.586 29.436 39.96 ; 
      RECT 28.48 35.586 28.584 39.96 ; 
      RECT 28.048 35.586 28.152 39.96 ; 
      RECT 27.616 35.586 27.72 39.96 ; 
      RECT 27.184 35.586 27.288 39.96 ; 
      RECT 26.752 35.586 26.856 39.96 ; 
      RECT 26.32 35.586 26.424 39.96 ; 
      RECT 25.888 35.586 25.992 39.96 ; 
      RECT 25.456 35.586 25.56 39.96 ; 
      RECT 25.024 35.586 25.128 39.96 ; 
      RECT 24.592 35.586 24.696 39.96 ; 
      RECT 24.16 35.586 24.264 39.96 ; 
      RECT 23.728 35.586 23.832 39.96 ; 
      RECT 23.296 35.586 23.4 39.96 ; 
      RECT 22.864 35.586 22.968 39.96 ; 
      RECT 22.432 35.586 22.536 39.96 ; 
      RECT 22 35.586 22.104 39.96 ; 
      RECT 21.568 35.586 21.672 39.96 ; 
      RECT 21.136 35.586 21.24 39.96 ; 
      RECT 20.704 35.586 20.808 39.96 ; 
      RECT 20.272 35.586 20.376 39.96 ; 
      RECT 19.84 35.586 19.944 39.96 ; 
      RECT 19.408 35.586 19.512 39.96 ; 
      RECT 18.976 35.586 19.08 39.96 ; 
      RECT 18.544 35.586 18.648 39.96 ; 
      RECT 18.112 35.586 18.216 39.96 ; 
      RECT 17.68 35.586 17.784 39.96 ; 
      RECT 17.248 35.586 17.352 39.96 ; 
      RECT 16.816 35.586 16.92 39.96 ; 
      RECT 16.384 35.586 16.488 39.96 ; 
      RECT 15.952 35.586 16.056 39.96 ; 
      RECT 15.52 35.586 15.624 39.96 ; 
      RECT 15.088 35.586 15.192 39.96 ; 
      RECT 14.656 35.586 14.76 39.96 ; 
      RECT 14.224 35.586 14.328 39.96 ; 
      RECT 13.792 35.586 13.896 39.96 ; 
      RECT 13.36 35.586 13.464 39.96 ; 
      RECT 12.928 35.586 13.032 39.96 ; 
      RECT 12.496 35.586 12.6 39.96 ; 
      RECT 12.064 35.586 12.168 39.96 ; 
      RECT 11.632 35.586 11.736 39.96 ; 
      RECT 11.2 35.586 11.304 39.96 ; 
      RECT 10.768 35.586 10.872 39.96 ; 
      RECT 10.336 35.586 10.44 39.96 ; 
      RECT 9.904 35.586 10.008 39.96 ; 
      RECT 9.472 35.586 9.576 39.96 ; 
      RECT 9.04 35.586 9.144 39.96 ; 
      RECT 8.608 35.586 8.712 39.96 ; 
      RECT 8.176 35.586 8.28 39.96 ; 
      RECT 7.744 35.586 7.848 39.96 ; 
      RECT 7.312 35.586 7.416 39.96 ; 
      RECT 6.88 35.586 6.984 39.96 ; 
      RECT 6.448 35.586 6.552 39.96 ; 
      RECT 6.016 35.586 6.12 39.96 ; 
      RECT 5.584 35.586 5.688 39.96 ; 
      RECT 5.152 35.586 5.256 39.96 ; 
      RECT 4.72 35.586 4.824 39.96 ; 
      RECT 4.288 35.586 4.392 39.96 ; 
      RECT 3.856 35.586 3.96 39.96 ; 
      RECT 3.424 35.586 3.528 39.96 ; 
      RECT 2.992 35.586 3.096 39.96 ; 
      RECT 2.56 35.586 2.664 39.96 ; 
      RECT 2.128 35.586 2.232 39.96 ; 
      RECT 1.696 35.586 1.8 39.96 ; 
      RECT 1.264 35.586 1.368 39.96 ; 
      RECT 0.832 35.586 0.936 39.96 ; 
      RECT 0.02 35.586 0.36 39.96 ; 
      RECT 34.564 39.906 35.076 44.28 ; 
      RECT 34.508 42.568 35.076 43.858 ; 
      RECT 33.916 41.476 34.164 44.28 ; 
      RECT 33.86 42.714 34.164 43.328 ; 
      RECT 33.916 39.906 34.02 44.28 ; 
      RECT 33.916 40.39 34.076 41.348 ; 
      RECT 33.916 39.906 34.164 40.262 ; 
      RECT 32.728 41.708 33.552 44.28 ; 
      RECT 33.448 39.906 33.552 44.28 ; 
      RECT 32.728 42.816 33.608 43.848 ; 
      RECT 32.728 39.906 33.12 44.28 ; 
      RECT 31.06 39.906 31.392 44.28 ; 
      RECT 31.06 40.26 31.448 44.002 ; 
      RECT 65.776 39.906 66.116 44.28 ; 
      RECT 65.2 39.906 65.304 44.28 ; 
      RECT 64.768 39.906 64.872 44.28 ; 
      RECT 64.336 39.906 64.44 44.28 ; 
      RECT 63.904 39.906 64.008 44.28 ; 
      RECT 63.472 39.906 63.576 44.28 ; 
      RECT 63.04 39.906 63.144 44.28 ; 
      RECT 62.608 39.906 62.712 44.28 ; 
      RECT 62.176 39.906 62.28 44.28 ; 
      RECT 61.744 39.906 61.848 44.28 ; 
      RECT 61.312 39.906 61.416 44.28 ; 
      RECT 60.88 39.906 60.984 44.28 ; 
      RECT 60.448 39.906 60.552 44.28 ; 
      RECT 60.016 39.906 60.12 44.28 ; 
      RECT 59.584 39.906 59.688 44.28 ; 
      RECT 59.152 39.906 59.256 44.28 ; 
      RECT 58.72 39.906 58.824 44.28 ; 
      RECT 58.288 39.906 58.392 44.28 ; 
      RECT 57.856 39.906 57.96 44.28 ; 
      RECT 57.424 39.906 57.528 44.28 ; 
      RECT 56.992 39.906 57.096 44.28 ; 
      RECT 56.56 39.906 56.664 44.28 ; 
      RECT 56.128 39.906 56.232 44.28 ; 
      RECT 55.696 39.906 55.8 44.28 ; 
      RECT 55.264 39.906 55.368 44.28 ; 
      RECT 54.832 39.906 54.936 44.28 ; 
      RECT 54.4 39.906 54.504 44.28 ; 
      RECT 53.968 39.906 54.072 44.28 ; 
      RECT 53.536 39.906 53.64 44.28 ; 
      RECT 53.104 39.906 53.208 44.28 ; 
      RECT 52.672 39.906 52.776 44.28 ; 
      RECT 52.24 39.906 52.344 44.28 ; 
      RECT 51.808 39.906 51.912 44.28 ; 
      RECT 51.376 39.906 51.48 44.28 ; 
      RECT 50.944 39.906 51.048 44.28 ; 
      RECT 50.512 39.906 50.616 44.28 ; 
      RECT 50.08 39.906 50.184 44.28 ; 
      RECT 49.648 39.906 49.752 44.28 ; 
      RECT 49.216 39.906 49.32 44.28 ; 
      RECT 48.784 39.906 48.888 44.28 ; 
      RECT 48.352 39.906 48.456 44.28 ; 
      RECT 47.92 39.906 48.024 44.28 ; 
      RECT 47.488 39.906 47.592 44.28 ; 
      RECT 47.056 39.906 47.16 44.28 ; 
      RECT 46.624 39.906 46.728 44.28 ; 
      RECT 46.192 39.906 46.296 44.28 ; 
      RECT 45.76 39.906 45.864 44.28 ; 
      RECT 45.328 39.906 45.432 44.28 ; 
      RECT 44.896 39.906 45 44.28 ; 
      RECT 44.464 39.906 44.568 44.28 ; 
      RECT 44.032 39.906 44.136 44.28 ; 
      RECT 43.6 39.906 43.704 44.28 ; 
      RECT 43.168 39.906 43.272 44.28 ; 
      RECT 42.736 39.906 42.84 44.28 ; 
      RECT 42.304 39.906 42.408 44.28 ; 
      RECT 41.872 39.906 41.976 44.28 ; 
      RECT 41.44 39.906 41.544 44.28 ; 
      RECT 41.008 39.906 41.112 44.28 ; 
      RECT 40.576 39.906 40.68 44.28 ; 
      RECT 40.144 39.906 40.248 44.28 ; 
      RECT 39.712 39.906 39.816 44.28 ; 
      RECT 39.28 39.906 39.384 44.28 ; 
      RECT 38.848 39.906 38.952 44.28 ; 
      RECT 38.416 39.906 38.52 44.28 ; 
      RECT 37.984 39.906 38.088 44.28 ; 
      RECT 37.552 39.906 37.656 44.28 ; 
      RECT 36.7 39.906 37.008 44.28 ; 
      RECT 29.128 39.906 29.436 44.28 ; 
      RECT 28.48 39.906 28.584 44.28 ; 
      RECT 28.048 39.906 28.152 44.28 ; 
      RECT 27.616 39.906 27.72 44.28 ; 
      RECT 27.184 39.906 27.288 44.28 ; 
      RECT 26.752 39.906 26.856 44.28 ; 
      RECT 26.32 39.906 26.424 44.28 ; 
      RECT 25.888 39.906 25.992 44.28 ; 
      RECT 25.456 39.906 25.56 44.28 ; 
      RECT 25.024 39.906 25.128 44.28 ; 
      RECT 24.592 39.906 24.696 44.28 ; 
      RECT 24.16 39.906 24.264 44.28 ; 
      RECT 23.728 39.906 23.832 44.28 ; 
      RECT 23.296 39.906 23.4 44.28 ; 
      RECT 22.864 39.906 22.968 44.28 ; 
      RECT 22.432 39.906 22.536 44.28 ; 
      RECT 22 39.906 22.104 44.28 ; 
      RECT 21.568 39.906 21.672 44.28 ; 
      RECT 21.136 39.906 21.24 44.28 ; 
      RECT 20.704 39.906 20.808 44.28 ; 
      RECT 20.272 39.906 20.376 44.28 ; 
      RECT 19.84 39.906 19.944 44.28 ; 
      RECT 19.408 39.906 19.512 44.28 ; 
      RECT 18.976 39.906 19.08 44.28 ; 
      RECT 18.544 39.906 18.648 44.28 ; 
      RECT 18.112 39.906 18.216 44.28 ; 
      RECT 17.68 39.906 17.784 44.28 ; 
      RECT 17.248 39.906 17.352 44.28 ; 
      RECT 16.816 39.906 16.92 44.28 ; 
      RECT 16.384 39.906 16.488 44.28 ; 
      RECT 15.952 39.906 16.056 44.28 ; 
      RECT 15.52 39.906 15.624 44.28 ; 
      RECT 15.088 39.906 15.192 44.28 ; 
      RECT 14.656 39.906 14.76 44.28 ; 
      RECT 14.224 39.906 14.328 44.28 ; 
      RECT 13.792 39.906 13.896 44.28 ; 
      RECT 13.36 39.906 13.464 44.28 ; 
      RECT 12.928 39.906 13.032 44.28 ; 
      RECT 12.496 39.906 12.6 44.28 ; 
      RECT 12.064 39.906 12.168 44.28 ; 
      RECT 11.632 39.906 11.736 44.28 ; 
      RECT 11.2 39.906 11.304 44.28 ; 
      RECT 10.768 39.906 10.872 44.28 ; 
      RECT 10.336 39.906 10.44 44.28 ; 
      RECT 9.904 39.906 10.008 44.28 ; 
      RECT 9.472 39.906 9.576 44.28 ; 
      RECT 9.04 39.906 9.144 44.28 ; 
      RECT 8.608 39.906 8.712 44.28 ; 
      RECT 8.176 39.906 8.28 44.28 ; 
      RECT 7.744 39.906 7.848 44.28 ; 
      RECT 7.312 39.906 7.416 44.28 ; 
      RECT 6.88 39.906 6.984 44.28 ; 
      RECT 6.448 39.906 6.552 44.28 ; 
      RECT 6.016 39.906 6.12 44.28 ; 
      RECT 5.584 39.906 5.688 44.28 ; 
      RECT 5.152 39.906 5.256 44.28 ; 
      RECT 4.72 39.906 4.824 44.28 ; 
      RECT 4.288 39.906 4.392 44.28 ; 
      RECT 3.856 39.906 3.96 44.28 ; 
      RECT 3.424 39.906 3.528 44.28 ; 
      RECT 2.992 39.906 3.096 44.28 ; 
      RECT 2.56 39.906 2.664 44.28 ; 
      RECT 2.128 39.906 2.232 44.28 ; 
      RECT 1.696 39.906 1.8 44.28 ; 
      RECT 1.264 39.906 1.368 44.28 ; 
      RECT 0.832 39.906 0.936 44.28 ; 
      RECT 0.02 39.906 0.36 44.28 ; 
      RECT 34.564 44.226 35.076 48.6 ; 
      RECT 34.508 46.888 35.076 48.178 ; 
      RECT 33.916 45.796 34.164 48.6 ; 
      RECT 33.86 47.034 34.164 47.648 ; 
      RECT 33.916 44.226 34.02 48.6 ; 
      RECT 33.916 44.71 34.076 45.668 ; 
      RECT 33.916 44.226 34.164 44.582 ; 
      RECT 32.728 46.028 33.552 48.6 ; 
      RECT 33.448 44.226 33.552 48.6 ; 
      RECT 32.728 47.136 33.608 48.168 ; 
      RECT 32.728 44.226 33.12 48.6 ; 
      RECT 31.06 44.226 31.392 48.6 ; 
      RECT 31.06 44.58 31.448 48.322 ; 
      RECT 65.776 44.226 66.116 48.6 ; 
      RECT 65.2 44.226 65.304 48.6 ; 
      RECT 64.768 44.226 64.872 48.6 ; 
      RECT 64.336 44.226 64.44 48.6 ; 
      RECT 63.904 44.226 64.008 48.6 ; 
      RECT 63.472 44.226 63.576 48.6 ; 
      RECT 63.04 44.226 63.144 48.6 ; 
      RECT 62.608 44.226 62.712 48.6 ; 
      RECT 62.176 44.226 62.28 48.6 ; 
      RECT 61.744 44.226 61.848 48.6 ; 
      RECT 61.312 44.226 61.416 48.6 ; 
      RECT 60.88 44.226 60.984 48.6 ; 
      RECT 60.448 44.226 60.552 48.6 ; 
      RECT 60.016 44.226 60.12 48.6 ; 
      RECT 59.584 44.226 59.688 48.6 ; 
      RECT 59.152 44.226 59.256 48.6 ; 
      RECT 58.72 44.226 58.824 48.6 ; 
      RECT 58.288 44.226 58.392 48.6 ; 
      RECT 57.856 44.226 57.96 48.6 ; 
      RECT 57.424 44.226 57.528 48.6 ; 
      RECT 56.992 44.226 57.096 48.6 ; 
      RECT 56.56 44.226 56.664 48.6 ; 
      RECT 56.128 44.226 56.232 48.6 ; 
      RECT 55.696 44.226 55.8 48.6 ; 
      RECT 55.264 44.226 55.368 48.6 ; 
      RECT 54.832 44.226 54.936 48.6 ; 
      RECT 54.4 44.226 54.504 48.6 ; 
      RECT 53.968 44.226 54.072 48.6 ; 
      RECT 53.536 44.226 53.64 48.6 ; 
      RECT 53.104 44.226 53.208 48.6 ; 
      RECT 52.672 44.226 52.776 48.6 ; 
      RECT 52.24 44.226 52.344 48.6 ; 
      RECT 51.808 44.226 51.912 48.6 ; 
      RECT 51.376 44.226 51.48 48.6 ; 
      RECT 50.944 44.226 51.048 48.6 ; 
      RECT 50.512 44.226 50.616 48.6 ; 
      RECT 50.08 44.226 50.184 48.6 ; 
      RECT 49.648 44.226 49.752 48.6 ; 
      RECT 49.216 44.226 49.32 48.6 ; 
      RECT 48.784 44.226 48.888 48.6 ; 
      RECT 48.352 44.226 48.456 48.6 ; 
      RECT 47.92 44.226 48.024 48.6 ; 
      RECT 47.488 44.226 47.592 48.6 ; 
      RECT 47.056 44.226 47.16 48.6 ; 
      RECT 46.624 44.226 46.728 48.6 ; 
      RECT 46.192 44.226 46.296 48.6 ; 
      RECT 45.76 44.226 45.864 48.6 ; 
      RECT 45.328 44.226 45.432 48.6 ; 
      RECT 44.896 44.226 45 48.6 ; 
      RECT 44.464 44.226 44.568 48.6 ; 
      RECT 44.032 44.226 44.136 48.6 ; 
      RECT 43.6 44.226 43.704 48.6 ; 
      RECT 43.168 44.226 43.272 48.6 ; 
      RECT 42.736 44.226 42.84 48.6 ; 
      RECT 42.304 44.226 42.408 48.6 ; 
      RECT 41.872 44.226 41.976 48.6 ; 
      RECT 41.44 44.226 41.544 48.6 ; 
      RECT 41.008 44.226 41.112 48.6 ; 
      RECT 40.576 44.226 40.68 48.6 ; 
      RECT 40.144 44.226 40.248 48.6 ; 
      RECT 39.712 44.226 39.816 48.6 ; 
      RECT 39.28 44.226 39.384 48.6 ; 
      RECT 38.848 44.226 38.952 48.6 ; 
      RECT 38.416 44.226 38.52 48.6 ; 
      RECT 37.984 44.226 38.088 48.6 ; 
      RECT 37.552 44.226 37.656 48.6 ; 
      RECT 36.7 44.226 37.008 48.6 ; 
      RECT 29.128 44.226 29.436 48.6 ; 
      RECT 28.48 44.226 28.584 48.6 ; 
      RECT 28.048 44.226 28.152 48.6 ; 
      RECT 27.616 44.226 27.72 48.6 ; 
      RECT 27.184 44.226 27.288 48.6 ; 
      RECT 26.752 44.226 26.856 48.6 ; 
      RECT 26.32 44.226 26.424 48.6 ; 
      RECT 25.888 44.226 25.992 48.6 ; 
      RECT 25.456 44.226 25.56 48.6 ; 
      RECT 25.024 44.226 25.128 48.6 ; 
      RECT 24.592 44.226 24.696 48.6 ; 
      RECT 24.16 44.226 24.264 48.6 ; 
      RECT 23.728 44.226 23.832 48.6 ; 
      RECT 23.296 44.226 23.4 48.6 ; 
      RECT 22.864 44.226 22.968 48.6 ; 
      RECT 22.432 44.226 22.536 48.6 ; 
      RECT 22 44.226 22.104 48.6 ; 
      RECT 21.568 44.226 21.672 48.6 ; 
      RECT 21.136 44.226 21.24 48.6 ; 
      RECT 20.704 44.226 20.808 48.6 ; 
      RECT 20.272 44.226 20.376 48.6 ; 
      RECT 19.84 44.226 19.944 48.6 ; 
      RECT 19.408 44.226 19.512 48.6 ; 
      RECT 18.976 44.226 19.08 48.6 ; 
      RECT 18.544 44.226 18.648 48.6 ; 
      RECT 18.112 44.226 18.216 48.6 ; 
      RECT 17.68 44.226 17.784 48.6 ; 
      RECT 17.248 44.226 17.352 48.6 ; 
      RECT 16.816 44.226 16.92 48.6 ; 
      RECT 16.384 44.226 16.488 48.6 ; 
      RECT 15.952 44.226 16.056 48.6 ; 
      RECT 15.52 44.226 15.624 48.6 ; 
      RECT 15.088 44.226 15.192 48.6 ; 
      RECT 14.656 44.226 14.76 48.6 ; 
      RECT 14.224 44.226 14.328 48.6 ; 
      RECT 13.792 44.226 13.896 48.6 ; 
      RECT 13.36 44.226 13.464 48.6 ; 
      RECT 12.928 44.226 13.032 48.6 ; 
      RECT 12.496 44.226 12.6 48.6 ; 
      RECT 12.064 44.226 12.168 48.6 ; 
      RECT 11.632 44.226 11.736 48.6 ; 
      RECT 11.2 44.226 11.304 48.6 ; 
      RECT 10.768 44.226 10.872 48.6 ; 
      RECT 10.336 44.226 10.44 48.6 ; 
      RECT 9.904 44.226 10.008 48.6 ; 
      RECT 9.472 44.226 9.576 48.6 ; 
      RECT 9.04 44.226 9.144 48.6 ; 
      RECT 8.608 44.226 8.712 48.6 ; 
      RECT 8.176 44.226 8.28 48.6 ; 
      RECT 7.744 44.226 7.848 48.6 ; 
      RECT 7.312 44.226 7.416 48.6 ; 
      RECT 6.88 44.226 6.984 48.6 ; 
      RECT 6.448 44.226 6.552 48.6 ; 
      RECT 6.016 44.226 6.12 48.6 ; 
      RECT 5.584 44.226 5.688 48.6 ; 
      RECT 5.152 44.226 5.256 48.6 ; 
      RECT 4.72 44.226 4.824 48.6 ; 
      RECT 4.288 44.226 4.392 48.6 ; 
      RECT 3.856 44.226 3.96 48.6 ; 
      RECT 3.424 44.226 3.528 48.6 ; 
      RECT 2.992 44.226 3.096 48.6 ; 
      RECT 2.56 44.226 2.664 48.6 ; 
      RECT 2.128 44.226 2.232 48.6 ; 
      RECT 1.696 44.226 1.8 48.6 ; 
      RECT 1.264 44.226 1.368 48.6 ; 
      RECT 0.832 44.226 0.936 48.6 ; 
      RECT 0.02 44.226 0.36 48.6 ; 
      RECT 34.564 48.546 35.076 52.92 ; 
      RECT 34.508 51.208 35.076 52.498 ; 
      RECT 33.916 50.116 34.164 52.92 ; 
      RECT 33.86 51.354 34.164 51.968 ; 
      RECT 33.916 48.546 34.02 52.92 ; 
      RECT 33.916 49.03 34.076 49.988 ; 
      RECT 33.916 48.546 34.164 48.902 ; 
      RECT 32.728 50.348 33.552 52.92 ; 
      RECT 33.448 48.546 33.552 52.92 ; 
      RECT 32.728 51.456 33.608 52.488 ; 
      RECT 32.728 48.546 33.12 52.92 ; 
      RECT 31.06 48.546 31.392 52.92 ; 
      RECT 31.06 48.9 31.448 52.642 ; 
      RECT 65.776 48.546 66.116 52.92 ; 
      RECT 65.2 48.546 65.304 52.92 ; 
      RECT 64.768 48.546 64.872 52.92 ; 
      RECT 64.336 48.546 64.44 52.92 ; 
      RECT 63.904 48.546 64.008 52.92 ; 
      RECT 63.472 48.546 63.576 52.92 ; 
      RECT 63.04 48.546 63.144 52.92 ; 
      RECT 62.608 48.546 62.712 52.92 ; 
      RECT 62.176 48.546 62.28 52.92 ; 
      RECT 61.744 48.546 61.848 52.92 ; 
      RECT 61.312 48.546 61.416 52.92 ; 
      RECT 60.88 48.546 60.984 52.92 ; 
      RECT 60.448 48.546 60.552 52.92 ; 
      RECT 60.016 48.546 60.12 52.92 ; 
      RECT 59.584 48.546 59.688 52.92 ; 
      RECT 59.152 48.546 59.256 52.92 ; 
      RECT 58.72 48.546 58.824 52.92 ; 
      RECT 58.288 48.546 58.392 52.92 ; 
      RECT 57.856 48.546 57.96 52.92 ; 
      RECT 57.424 48.546 57.528 52.92 ; 
      RECT 56.992 48.546 57.096 52.92 ; 
      RECT 56.56 48.546 56.664 52.92 ; 
      RECT 56.128 48.546 56.232 52.92 ; 
      RECT 55.696 48.546 55.8 52.92 ; 
      RECT 55.264 48.546 55.368 52.92 ; 
      RECT 54.832 48.546 54.936 52.92 ; 
      RECT 54.4 48.546 54.504 52.92 ; 
      RECT 53.968 48.546 54.072 52.92 ; 
      RECT 53.536 48.546 53.64 52.92 ; 
      RECT 53.104 48.546 53.208 52.92 ; 
      RECT 52.672 48.546 52.776 52.92 ; 
      RECT 52.24 48.546 52.344 52.92 ; 
      RECT 51.808 48.546 51.912 52.92 ; 
      RECT 51.376 48.546 51.48 52.92 ; 
      RECT 50.944 48.546 51.048 52.92 ; 
      RECT 50.512 48.546 50.616 52.92 ; 
      RECT 50.08 48.546 50.184 52.92 ; 
      RECT 49.648 48.546 49.752 52.92 ; 
      RECT 49.216 48.546 49.32 52.92 ; 
      RECT 48.784 48.546 48.888 52.92 ; 
      RECT 48.352 48.546 48.456 52.92 ; 
      RECT 47.92 48.546 48.024 52.92 ; 
      RECT 47.488 48.546 47.592 52.92 ; 
      RECT 47.056 48.546 47.16 52.92 ; 
      RECT 46.624 48.546 46.728 52.92 ; 
      RECT 46.192 48.546 46.296 52.92 ; 
      RECT 45.76 48.546 45.864 52.92 ; 
      RECT 45.328 48.546 45.432 52.92 ; 
      RECT 44.896 48.546 45 52.92 ; 
      RECT 44.464 48.546 44.568 52.92 ; 
      RECT 44.032 48.546 44.136 52.92 ; 
      RECT 43.6 48.546 43.704 52.92 ; 
      RECT 43.168 48.546 43.272 52.92 ; 
      RECT 42.736 48.546 42.84 52.92 ; 
      RECT 42.304 48.546 42.408 52.92 ; 
      RECT 41.872 48.546 41.976 52.92 ; 
      RECT 41.44 48.546 41.544 52.92 ; 
      RECT 41.008 48.546 41.112 52.92 ; 
      RECT 40.576 48.546 40.68 52.92 ; 
      RECT 40.144 48.546 40.248 52.92 ; 
      RECT 39.712 48.546 39.816 52.92 ; 
      RECT 39.28 48.546 39.384 52.92 ; 
      RECT 38.848 48.546 38.952 52.92 ; 
      RECT 38.416 48.546 38.52 52.92 ; 
      RECT 37.984 48.546 38.088 52.92 ; 
      RECT 37.552 48.546 37.656 52.92 ; 
      RECT 36.7 48.546 37.008 52.92 ; 
      RECT 29.128 48.546 29.436 52.92 ; 
      RECT 28.48 48.546 28.584 52.92 ; 
      RECT 28.048 48.546 28.152 52.92 ; 
      RECT 27.616 48.546 27.72 52.92 ; 
      RECT 27.184 48.546 27.288 52.92 ; 
      RECT 26.752 48.546 26.856 52.92 ; 
      RECT 26.32 48.546 26.424 52.92 ; 
      RECT 25.888 48.546 25.992 52.92 ; 
      RECT 25.456 48.546 25.56 52.92 ; 
      RECT 25.024 48.546 25.128 52.92 ; 
      RECT 24.592 48.546 24.696 52.92 ; 
      RECT 24.16 48.546 24.264 52.92 ; 
      RECT 23.728 48.546 23.832 52.92 ; 
      RECT 23.296 48.546 23.4 52.92 ; 
      RECT 22.864 48.546 22.968 52.92 ; 
      RECT 22.432 48.546 22.536 52.92 ; 
      RECT 22 48.546 22.104 52.92 ; 
      RECT 21.568 48.546 21.672 52.92 ; 
      RECT 21.136 48.546 21.24 52.92 ; 
      RECT 20.704 48.546 20.808 52.92 ; 
      RECT 20.272 48.546 20.376 52.92 ; 
      RECT 19.84 48.546 19.944 52.92 ; 
      RECT 19.408 48.546 19.512 52.92 ; 
      RECT 18.976 48.546 19.08 52.92 ; 
      RECT 18.544 48.546 18.648 52.92 ; 
      RECT 18.112 48.546 18.216 52.92 ; 
      RECT 17.68 48.546 17.784 52.92 ; 
      RECT 17.248 48.546 17.352 52.92 ; 
      RECT 16.816 48.546 16.92 52.92 ; 
      RECT 16.384 48.546 16.488 52.92 ; 
      RECT 15.952 48.546 16.056 52.92 ; 
      RECT 15.52 48.546 15.624 52.92 ; 
      RECT 15.088 48.546 15.192 52.92 ; 
      RECT 14.656 48.546 14.76 52.92 ; 
      RECT 14.224 48.546 14.328 52.92 ; 
      RECT 13.792 48.546 13.896 52.92 ; 
      RECT 13.36 48.546 13.464 52.92 ; 
      RECT 12.928 48.546 13.032 52.92 ; 
      RECT 12.496 48.546 12.6 52.92 ; 
      RECT 12.064 48.546 12.168 52.92 ; 
      RECT 11.632 48.546 11.736 52.92 ; 
      RECT 11.2 48.546 11.304 52.92 ; 
      RECT 10.768 48.546 10.872 52.92 ; 
      RECT 10.336 48.546 10.44 52.92 ; 
      RECT 9.904 48.546 10.008 52.92 ; 
      RECT 9.472 48.546 9.576 52.92 ; 
      RECT 9.04 48.546 9.144 52.92 ; 
      RECT 8.608 48.546 8.712 52.92 ; 
      RECT 8.176 48.546 8.28 52.92 ; 
      RECT 7.744 48.546 7.848 52.92 ; 
      RECT 7.312 48.546 7.416 52.92 ; 
      RECT 6.88 48.546 6.984 52.92 ; 
      RECT 6.448 48.546 6.552 52.92 ; 
      RECT 6.016 48.546 6.12 52.92 ; 
      RECT 5.584 48.546 5.688 52.92 ; 
      RECT 5.152 48.546 5.256 52.92 ; 
      RECT 4.72 48.546 4.824 52.92 ; 
      RECT 4.288 48.546 4.392 52.92 ; 
      RECT 3.856 48.546 3.96 52.92 ; 
      RECT 3.424 48.546 3.528 52.92 ; 
      RECT 2.992 48.546 3.096 52.92 ; 
      RECT 2.56 48.546 2.664 52.92 ; 
      RECT 2.128 48.546 2.232 52.92 ; 
      RECT 1.696 48.546 1.8 52.92 ; 
      RECT 1.264 48.546 1.368 52.92 ; 
      RECT 0.832 48.546 0.936 52.92 ; 
      RECT 0.02 48.546 0.36 52.92 ; 
      RECT 34.564 52.866 35.076 57.24 ; 
      RECT 34.508 55.528 35.076 56.818 ; 
      RECT 33.916 54.436 34.164 57.24 ; 
      RECT 33.86 55.674 34.164 56.288 ; 
      RECT 33.916 52.866 34.02 57.24 ; 
      RECT 33.916 53.35 34.076 54.308 ; 
      RECT 33.916 52.866 34.164 53.222 ; 
      RECT 32.728 54.668 33.552 57.24 ; 
      RECT 33.448 52.866 33.552 57.24 ; 
      RECT 32.728 55.776 33.608 56.808 ; 
      RECT 32.728 52.866 33.12 57.24 ; 
      RECT 31.06 52.866 31.392 57.24 ; 
      RECT 31.06 53.22 31.448 56.962 ; 
      RECT 65.776 52.866 66.116 57.24 ; 
      RECT 65.2 52.866 65.304 57.24 ; 
      RECT 64.768 52.866 64.872 57.24 ; 
      RECT 64.336 52.866 64.44 57.24 ; 
      RECT 63.904 52.866 64.008 57.24 ; 
      RECT 63.472 52.866 63.576 57.24 ; 
      RECT 63.04 52.866 63.144 57.24 ; 
      RECT 62.608 52.866 62.712 57.24 ; 
      RECT 62.176 52.866 62.28 57.24 ; 
      RECT 61.744 52.866 61.848 57.24 ; 
      RECT 61.312 52.866 61.416 57.24 ; 
      RECT 60.88 52.866 60.984 57.24 ; 
      RECT 60.448 52.866 60.552 57.24 ; 
      RECT 60.016 52.866 60.12 57.24 ; 
      RECT 59.584 52.866 59.688 57.24 ; 
      RECT 59.152 52.866 59.256 57.24 ; 
      RECT 58.72 52.866 58.824 57.24 ; 
      RECT 58.288 52.866 58.392 57.24 ; 
      RECT 57.856 52.866 57.96 57.24 ; 
      RECT 57.424 52.866 57.528 57.24 ; 
      RECT 56.992 52.866 57.096 57.24 ; 
      RECT 56.56 52.866 56.664 57.24 ; 
      RECT 56.128 52.866 56.232 57.24 ; 
      RECT 55.696 52.866 55.8 57.24 ; 
      RECT 55.264 52.866 55.368 57.24 ; 
      RECT 54.832 52.866 54.936 57.24 ; 
      RECT 54.4 52.866 54.504 57.24 ; 
      RECT 53.968 52.866 54.072 57.24 ; 
      RECT 53.536 52.866 53.64 57.24 ; 
      RECT 53.104 52.866 53.208 57.24 ; 
      RECT 52.672 52.866 52.776 57.24 ; 
      RECT 52.24 52.866 52.344 57.24 ; 
      RECT 51.808 52.866 51.912 57.24 ; 
      RECT 51.376 52.866 51.48 57.24 ; 
      RECT 50.944 52.866 51.048 57.24 ; 
      RECT 50.512 52.866 50.616 57.24 ; 
      RECT 50.08 52.866 50.184 57.24 ; 
      RECT 49.648 52.866 49.752 57.24 ; 
      RECT 49.216 52.866 49.32 57.24 ; 
      RECT 48.784 52.866 48.888 57.24 ; 
      RECT 48.352 52.866 48.456 57.24 ; 
      RECT 47.92 52.866 48.024 57.24 ; 
      RECT 47.488 52.866 47.592 57.24 ; 
      RECT 47.056 52.866 47.16 57.24 ; 
      RECT 46.624 52.866 46.728 57.24 ; 
      RECT 46.192 52.866 46.296 57.24 ; 
      RECT 45.76 52.866 45.864 57.24 ; 
      RECT 45.328 52.866 45.432 57.24 ; 
      RECT 44.896 52.866 45 57.24 ; 
      RECT 44.464 52.866 44.568 57.24 ; 
      RECT 44.032 52.866 44.136 57.24 ; 
      RECT 43.6 52.866 43.704 57.24 ; 
      RECT 43.168 52.866 43.272 57.24 ; 
      RECT 42.736 52.866 42.84 57.24 ; 
      RECT 42.304 52.866 42.408 57.24 ; 
      RECT 41.872 52.866 41.976 57.24 ; 
      RECT 41.44 52.866 41.544 57.24 ; 
      RECT 41.008 52.866 41.112 57.24 ; 
      RECT 40.576 52.866 40.68 57.24 ; 
      RECT 40.144 52.866 40.248 57.24 ; 
      RECT 39.712 52.866 39.816 57.24 ; 
      RECT 39.28 52.866 39.384 57.24 ; 
      RECT 38.848 52.866 38.952 57.24 ; 
      RECT 38.416 52.866 38.52 57.24 ; 
      RECT 37.984 52.866 38.088 57.24 ; 
      RECT 37.552 52.866 37.656 57.24 ; 
      RECT 36.7 52.866 37.008 57.24 ; 
      RECT 29.128 52.866 29.436 57.24 ; 
      RECT 28.48 52.866 28.584 57.24 ; 
      RECT 28.048 52.866 28.152 57.24 ; 
      RECT 27.616 52.866 27.72 57.24 ; 
      RECT 27.184 52.866 27.288 57.24 ; 
      RECT 26.752 52.866 26.856 57.24 ; 
      RECT 26.32 52.866 26.424 57.24 ; 
      RECT 25.888 52.866 25.992 57.24 ; 
      RECT 25.456 52.866 25.56 57.24 ; 
      RECT 25.024 52.866 25.128 57.24 ; 
      RECT 24.592 52.866 24.696 57.24 ; 
      RECT 24.16 52.866 24.264 57.24 ; 
      RECT 23.728 52.866 23.832 57.24 ; 
      RECT 23.296 52.866 23.4 57.24 ; 
      RECT 22.864 52.866 22.968 57.24 ; 
      RECT 22.432 52.866 22.536 57.24 ; 
      RECT 22 52.866 22.104 57.24 ; 
      RECT 21.568 52.866 21.672 57.24 ; 
      RECT 21.136 52.866 21.24 57.24 ; 
      RECT 20.704 52.866 20.808 57.24 ; 
      RECT 20.272 52.866 20.376 57.24 ; 
      RECT 19.84 52.866 19.944 57.24 ; 
      RECT 19.408 52.866 19.512 57.24 ; 
      RECT 18.976 52.866 19.08 57.24 ; 
      RECT 18.544 52.866 18.648 57.24 ; 
      RECT 18.112 52.866 18.216 57.24 ; 
      RECT 17.68 52.866 17.784 57.24 ; 
      RECT 17.248 52.866 17.352 57.24 ; 
      RECT 16.816 52.866 16.92 57.24 ; 
      RECT 16.384 52.866 16.488 57.24 ; 
      RECT 15.952 52.866 16.056 57.24 ; 
      RECT 15.52 52.866 15.624 57.24 ; 
      RECT 15.088 52.866 15.192 57.24 ; 
      RECT 14.656 52.866 14.76 57.24 ; 
      RECT 14.224 52.866 14.328 57.24 ; 
      RECT 13.792 52.866 13.896 57.24 ; 
      RECT 13.36 52.866 13.464 57.24 ; 
      RECT 12.928 52.866 13.032 57.24 ; 
      RECT 12.496 52.866 12.6 57.24 ; 
      RECT 12.064 52.866 12.168 57.24 ; 
      RECT 11.632 52.866 11.736 57.24 ; 
      RECT 11.2 52.866 11.304 57.24 ; 
      RECT 10.768 52.866 10.872 57.24 ; 
      RECT 10.336 52.866 10.44 57.24 ; 
      RECT 9.904 52.866 10.008 57.24 ; 
      RECT 9.472 52.866 9.576 57.24 ; 
      RECT 9.04 52.866 9.144 57.24 ; 
      RECT 8.608 52.866 8.712 57.24 ; 
      RECT 8.176 52.866 8.28 57.24 ; 
      RECT 7.744 52.866 7.848 57.24 ; 
      RECT 7.312 52.866 7.416 57.24 ; 
      RECT 6.88 52.866 6.984 57.24 ; 
      RECT 6.448 52.866 6.552 57.24 ; 
      RECT 6.016 52.866 6.12 57.24 ; 
      RECT 5.584 52.866 5.688 57.24 ; 
      RECT 5.152 52.866 5.256 57.24 ; 
      RECT 4.72 52.866 4.824 57.24 ; 
      RECT 4.288 52.866 4.392 57.24 ; 
      RECT 3.856 52.866 3.96 57.24 ; 
      RECT 3.424 52.866 3.528 57.24 ; 
      RECT 2.992 52.866 3.096 57.24 ; 
      RECT 2.56 52.866 2.664 57.24 ; 
      RECT 2.128 52.866 2.232 57.24 ; 
      RECT 1.696 52.866 1.8 57.24 ; 
      RECT 1.264 52.866 1.368 57.24 ; 
      RECT 0.832 52.866 0.936 57.24 ; 
      RECT 0.02 52.866 0.36 57.24 ; 
      RECT 34.564 57.186 35.076 61.56 ; 
      RECT 34.508 59.848 35.076 61.138 ; 
      RECT 33.916 58.756 34.164 61.56 ; 
      RECT 33.86 59.994 34.164 60.608 ; 
      RECT 33.916 57.186 34.02 61.56 ; 
      RECT 33.916 57.67 34.076 58.628 ; 
      RECT 33.916 57.186 34.164 57.542 ; 
      RECT 32.728 58.988 33.552 61.56 ; 
      RECT 33.448 57.186 33.552 61.56 ; 
      RECT 32.728 60.096 33.608 61.128 ; 
      RECT 32.728 57.186 33.12 61.56 ; 
      RECT 31.06 57.186 31.392 61.56 ; 
      RECT 31.06 57.54 31.448 61.282 ; 
      RECT 65.776 57.186 66.116 61.56 ; 
      RECT 65.2 57.186 65.304 61.56 ; 
      RECT 64.768 57.186 64.872 61.56 ; 
      RECT 64.336 57.186 64.44 61.56 ; 
      RECT 63.904 57.186 64.008 61.56 ; 
      RECT 63.472 57.186 63.576 61.56 ; 
      RECT 63.04 57.186 63.144 61.56 ; 
      RECT 62.608 57.186 62.712 61.56 ; 
      RECT 62.176 57.186 62.28 61.56 ; 
      RECT 61.744 57.186 61.848 61.56 ; 
      RECT 61.312 57.186 61.416 61.56 ; 
      RECT 60.88 57.186 60.984 61.56 ; 
      RECT 60.448 57.186 60.552 61.56 ; 
      RECT 60.016 57.186 60.12 61.56 ; 
      RECT 59.584 57.186 59.688 61.56 ; 
      RECT 59.152 57.186 59.256 61.56 ; 
      RECT 58.72 57.186 58.824 61.56 ; 
      RECT 58.288 57.186 58.392 61.56 ; 
      RECT 57.856 57.186 57.96 61.56 ; 
      RECT 57.424 57.186 57.528 61.56 ; 
      RECT 56.992 57.186 57.096 61.56 ; 
      RECT 56.56 57.186 56.664 61.56 ; 
      RECT 56.128 57.186 56.232 61.56 ; 
      RECT 55.696 57.186 55.8 61.56 ; 
      RECT 55.264 57.186 55.368 61.56 ; 
      RECT 54.832 57.186 54.936 61.56 ; 
      RECT 54.4 57.186 54.504 61.56 ; 
      RECT 53.968 57.186 54.072 61.56 ; 
      RECT 53.536 57.186 53.64 61.56 ; 
      RECT 53.104 57.186 53.208 61.56 ; 
      RECT 52.672 57.186 52.776 61.56 ; 
      RECT 52.24 57.186 52.344 61.56 ; 
      RECT 51.808 57.186 51.912 61.56 ; 
      RECT 51.376 57.186 51.48 61.56 ; 
      RECT 50.944 57.186 51.048 61.56 ; 
      RECT 50.512 57.186 50.616 61.56 ; 
      RECT 50.08 57.186 50.184 61.56 ; 
      RECT 49.648 57.186 49.752 61.56 ; 
      RECT 49.216 57.186 49.32 61.56 ; 
      RECT 48.784 57.186 48.888 61.56 ; 
      RECT 48.352 57.186 48.456 61.56 ; 
      RECT 47.92 57.186 48.024 61.56 ; 
      RECT 47.488 57.186 47.592 61.56 ; 
      RECT 47.056 57.186 47.16 61.56 ; 
      RECT 46.624 57.186 46.728 61.56 ; 
      RECT 46.192 57.186 46.296 61.56 ; 
      RECT 45.76 57.186 45.864 61.56 ; 
      RECT 45.328 57.186 45.432 61.56 ; 
      RECT 44.896 57.186 45 61.56 ; 
      RECT 44.464 57.186 44.568 61.56 ; 
      RECT 44.032 57.186 44.136 61.56 ; 
      RECT 43.6 57.186 43.704 61.56 ; 
      RECT 43.168 57.186 43.272 61.56 ; 
      RECT 42.736 57.186 42.84 61.56 ; 
      RECT 42.304 57.186 42.408 61.56 ; 
      RECT 41.872 57.186 41.976 61.56 ; 
      RECT 41.44 57.186 41.544 61.56 ; 
      RECT 41.008 57.186 41.112 61.56 ; 
      RECT 40.576 57.186 40.68 61.56 ; 
      RECT 40.144 57.186 40.248 61.56 ; 
      RECT 39.712 57.186 39.816 61.56 ; 
      RECT 39.28 57.186 39.384 61.56 ; 
      RECT 38.848 57.186 38.952 61.56 ; 
      RECT 38.416 57.186 38.52 61.56 ; 
      RECT 37.984 57.186 38.088 61.56 ; 
      RECT 37.552 57.186 37.656 61.56 ; 
      RECT 36.7 57.186 37.008 61.56 ; 
      RECT 29.128 57.186 29.436 61.56 ; 
      RECT 28.48 57.186 28.584 61.56 ; 
      RECT 28.048 57.186 28.152 61.56 ; 
      RECT 27.616 57.186 27.72 61.56 ; 
      RECT 27.184 57.186 27.288 61.56 ; 
      RECT 26.752 57.186 26.856 61.56 ; 
      RECT 26.32 57.186 26.424 61.56 ; 
      RECT 25.888 57.186 25.992 61.56 ; 
      RECT 25.456 57.186 25.56 61.56 ; 
      RECT 25.024 57.186 25.128 61.56 ; 
      RECT 24.592 57.186 24.696 61.56 ; 
      RECT 24.16 57.186 24.264 61.56 ; 
      RECT 23.728 57.186 23.832 61.56 ; 
      RECT 23.296 57.186 23.4 61.56 ; 
      RECT 22.864 57.186 22.968 61.56 ; 
      RECT 22.432 57.186 22.536 61.56 ; 
      RECT 22 57.186 22.104 61.56 ; 
      RECT 21.568 57.186 21.672 61.56 ; 
      RECT 21.136 57.186 21.24 61.56 ; 
      RECT 20.704 57.186 20.808 61.56 ; 
      RECT 20.272 57.186 20.376 61.56 ; 
      RECT 19.84 57.186 19.944 61.56 ; 
      RECT 19.408 57.186 19.512 61.56 ; 
      RECT 18.976 57.186 19.08 61.56 ; 
      RECT 18.544 57.186 18.648 61.56 ; 
      RECT 18.112 57.186 18.216 61.56 ; 
      RECT 17.68 57.186 17.784 61.56 ; 
      RECT 17.248 57.186 17.352 61.56 ; 
      RECT 16.816 57.186 16.92 61.56 ; 
      RECT 16.384 57.186 16.488 61.56 ; 
      RECT 15.952 57.186 16.056 61.56 ; 
      RECT 15.52 57.186 15.624 61.56 ; 
      RECT 15.088 57.186 15.192 61.56 ; 
      RECT 14.656 57.186 14.76 61.56 ; 
      RECT 14.224 57.186 14.328 61.56 ; 
      RECT 13.792 57.186 13.896 61.56 ; 
      RECT 13.36 57.186 13.464 61.56 ; 
      RECT 12.928 57.186 13.032 61.56 ; 
      RECT 12.496 57.186 12.6 61.56 ; 
      RECT 12.064 57.186 12.168 61.56 ; 
      RECT 11.632 57.186 11.736 61.56 ; 
      RECT 11.2 57.186 11.304 61.56 ; 
      RECT 10.768 57.186 10.872 61.56 ; 
      RECT 10.336 57.186 10.44 61.56 ; 
      RECT 9.904 57.186 10.008 61.56 ; 
      RECT 9.472 57.186 9.576 61.56 ; 
      RECT 9.04 57.186 9.144 61.56 ; 
      RECT 8.608 57.186 8.712 61.56 ; 
      RECT 8.176 57.186 8.28 61.56 ; 
      RECT 7.744 57.186 7.848 61.56 ; 
      RECT 7.312 57.186 7.416 61.56 ; 
      RECT 6.88 57.186 6.984 61.56 ; 
      RECT 6.448 57.186 6.552 61.56 ; 
      RECT 6.016 57.186 6.12 61.56 ; 
      RECT 5.584 57.186 5.688 61.56 ; 
      RECT 5.152 57.186 5.256 61.56 ; 
      RECT 4.72 57.186 4.824 61.56 ; 
      RECT 4.288 57.186 4.392 61.56 ; 
      RECT 3.856 57.186 3.96 61.56 ; 
      RECT 3.424 57.186 3.528 61.56 ; 
      RECT 2.992 57.186 3.096 61.56 ; 
      RECT 2.56 57.186 2.664 61.56 ; 
      RECT 2.128 57.186 2.232 61.56 ; 
      RECT 1.696 57.186 1.8 61.56 ; 
      RECT 1.264 57.186 1.368 61.56 ; 
      RECT 0.832 57.186 0.936 61.56 ; 
      RECT 0.02 57.186 0.36 61.56 ; 
      RECT 34.564 61.506 35.076 65.88 ; 
      RECT 34.508 64.168 35.076 65.458 ; 
      RECT 33.916 63.076 34.164 65.88 ; 
      RECT 33.86 64.314 34.164 64.928 ; 
      RECT 33.916 61.506 34.02 65.88 ; 
      RECT 33.916 61.99 34.076 62.948 ; 
      RECT 33.916 61.506 34.164 61.862 ; 
      RECT 32.728 63.308 33.552 65.88 ; 
      RECT 33.448 61.506 33.552 65.88 ; 
      RECT 32.728 64.416 33.608 65.448 ; 
      RECT 32.728 61.506 33.12 65.88 ; 
      RECT 31.06 61.506 31.392 65.88 ; 
      RECT 31.06 61.86 31.448 65.602 ; 
      RECT 65.776 61.506 66.116 65.88 ; 
      RECT 65.2 61.506 65.304 65.88 ; 
      RECT 64.768 61.506 64.872 65.88 ; 
      RECT 64.336 61.506 64.44 65.88 ; 
      RECT 63.904 61.506 64.008 65.88 ; 
      RECT 63.472 61.506 63.576 65.88 ; 
      RECT 63.04 61.506 63.144 65.88 ; 
      RECT 62.608 61.506 62.712 65.88 ; 
      RECT 62.176 61.506 62.28 65.88 ; 
      RECT 61.744 61.506 61.848 65.88 ; 
      RECT 61.312 61.506 61.416 65.88 ; 
      RECT 60.88 61.506 60.984 65.88 ; 
      RECT 60.448 61.506 60.552 65.88 ; 
      RECT 60.016 61.506 60.12 65.88 ; 
      RECT 59.584 61.506 59.688 65.88 ; 
      RECT 59.152 61.506 59.256 65.88 ; 
      RECT 58.72 61.506 58.824 65.88 ; 
      RECT 58.288 61.506 58.392 65.88 ; 
      RECT 57.856 61.506 57.96 65.88 ; 
      RECT 57.424 61.506 57.528 65.88 ; 
      RECT 56.992 61.506 57.096 65.88 ; 
      RECT 56.56 61.506 56.664 65.88 ; 
      RECT 56.128 61.506 56.232 65.88 ; 
      RECT 55.696 61.506 55.8 65.88 ; 
      RECT 55.264 61.506 55.368 65.88 ; 
      RECT 54.832 61.506 54.936 65.88 ; 
      RECT 54.4 61.506 54.504 65.88 ; 
      RECT 53.968 61.506 54.072 65.88 ; 
      RECT 53.536 61.506 53.64 65.88 ; 
      RECT 53.104 61.506 53.208 65.88 ; 
      RECT 52.672 61.506 52.776 65.88 ; 
      RECT 52.24 61.506 52.344 65.88 ; 
      RECT 51.808 61.506 51.912 65.88 ; 
      RECT 51.376 61.506 51.48 65.88 ; 
      RECT 50.944 61.506 51.048 65.88 ; 
      RECT 50.512 61.506 50.616 65.88 ; 
      RECT 50.08 61.506 50.184 65.88 ; 
      RECT 49.648 61.506 49.752 65.88 ; 
      RECT 49.216 61.506 49.32 65.88 ; 
      RECT 48.784 61.506 48.888 65.88 ; 
      RECT 48.352 61.506 48.456 65.88 ; 
      RECT 47.92 61.506 48.024 65.88 ; 
      RECT 47.488 61.506 47.592 65.88 ; 
      RECT 47.056 61.506 47.16 65.88 ; 
      RECT 46.624 61.506 46.728 65.88 ; 
      RECT 46.192 61.506 46.296 65.88 ; 
      RECT 45.76 61.506 45.864 65.88 ; 
      RECT 45.328 61.506 45.432 65.88 ; 
      RECT 44.896 61.506 45 65.88 ; 
      RECT 44.464 61.506 44.568 65.88 ; 
      RECT 44.032 61.506 44.136 65.88 ; 
      RECT 43.6 61.506 43.704 65.88 ; 
      RECT 43.168 61.506 43.272 65.88 ; 
      RECT 42.736 61.506 42.84 65.88 ; 
      RECT 42.304 61.506 42.408 65.88 ; 
      RECT 41.872 61.506 41.976 65.88 ; 
      RECT 41.44 61.506 41.544 65.88 ; 
      RECT 41.008 61.506 41.112 65.88 ; 
      RECT 40.576 61.506 40.68 65.88 ; 
      RECT 40.144 61.506 40.248 65.88 ; 
      RECT 39.712 61.506 39.816 65.88 ; 
      RECT 39.28 61.506 39.384 65.88 ; 
      RECT 38.848 61.506 38.952 65.88 ; 
      RECT 38.416 61.506 38.52 65.88 ; 
      RECT 37.984 61.506 38.088 65.88 ; 
      RECT 37.552 61.506 37.656 65.88 ; 
      RECT 36.7 61.506 37.008 65.88 ; 
      RECT 29.128 61.506 29.436 65.88 ; 
      RECT 28.48 61.506 28.584 65.88 ; 
      RECT 28.048 61.506 28.152 65.88 ; 
      RECT 27.616 61.506 27.72 65.88 ; 
      RECT 27.184 61.506 27.288 65.88 ; 
      RECT 26.752 61.506 26.856 65.88 ; 
      RECT 26.32 61.506 26.424 65.88 ; 
      RECT 25.888 61.506 25.992 65.88 ; 
      RECT 25.456 61.506 25.56 65.88 ; 
      RECT 25.024 61.506 25.128 65.88 ; 
      RECT 24.592 61.506 24.696 65.88 ; 
      RECT 24.16 61.506 24.264 65.88 ; 
      RECT 23.728 61.506 23.832 65.88 ; 
      RECT 23.296 61.506 23.4 65.88 ; 
      RECT 22.864 61.506 22.968 65.88 ; 
      RECT 22.432 61.506 22.536 65.88 ; 
      RECT 22 61.506 22.104 65.88 ; 
      RECT 21.568 61.506 21.672 65.88 ; 
      RECT 21.136 61.506 21.24 65.88 ; 
      RECT 20.704 61.506 20.808 65.88 ; 
      RECT 20.272 61.506 20.376 65.88 ; 
      RECT 19.84 61.506 19.944 65.88 ; 
      RECT 19.408 61.506 19.512 65.88 ; 
      RECT 18.976 61.506 19.08 65.88 ; 
      RECT 18.544 61.506 18.648 65.88 ; 
      RECT 18.112 61.506 18.216 65.88 ; 
      RECT 17.68 61.506 17.784 65.88 ; 
      RECT 17.248 61.506 17.352 65.88 ; 
      RECT 16.816 61.506 16.92 65.88 ; 
      RECT 16.384 61.506 16.488 65.88 ; 
      RECT 15.952 61.506 16.056 65.88 ; 
      RECT 15.52 61.506 15.624 65.88 ; 
      RECT 15.088 61.506 15.192 65.88 ; 
      RECT 14.656 61.506 14.76 65.88 ; 
      RECT 14.224 61.506 14.328 65.88 ; 
      RECT 13.792 61.506 13.896 65.88 ; 
      RECT 13.36 61.506 13.464 65.88 ; 
      RECT 12.928 61.506 13.032 65.88 ; 
      RECT 12.496 61.506 12.6 65.88 ; 
      RECT 12.064 61.506 12.168 65.88 ; 
      RECT 11.632 61.506 11.736 65.88 ; 
      RECT 11.2 61.506 11.304 65.88 ; 
      RECT 10.768 61.506 10.872 65.88 ; 
      RECT 10.336 61.506 10.44 65.88 ; 
      RECT 9.904 61.506 10.008 65.88 ; 
      RECT 9.472 61.506 9.576 65.88 ; 
      RECT 9.04 61.506 9.144 65.88 ; 
      RECT 8.608 61.506 8.712 65.88 ; 
      RECT 8.176 61.506 8.28 65.88 ; 
      RECT 7.744 61.506 7.848 65.88 ; 
      RECT 7.312 61.506 7.416 65.88 ; 
      RECT 6.88 61.506 6.984 65.88 ; 
      RECT 6.448 61.506 6.552 65.88 ; 
      RECT 6.016 61.506 6.12 65.88 ; 
      RECT 5.584 61.506 5.688 65.88 ; 
      RECT 5.152 61.506 5.256 65.88 ; 
      RECT 4.72 61.506 4.824 65.88 ; 
      RECT 4.288 61.506 4.392 65.88 ; 
      RECT 3.856 61.506 3.96 65.88 ; 
      RECT 3.424 61.506 3.528 65.88 ; 
      RECT 2.992 61.506 3.096 65.88 ; 
      RECT 2.56 61.506 2.664 65.88 ; 
      RECT 2.128 61.506 2.232 65.88 ; 
      RECT 1.696 61.506 1.8 65.88 ; 
      RECT 1.264 61.506 1.368 65.88 ; 
      RECT 0.832 61.506 0.936 65.88 ; 
      RECT 0.02 61.506 0.36 65.88 ; 
      RECT 34.564 65.826 35.076 70.2 ; 
      RECT 34.508 68.488 35.076 69.778 ; 
      RECT 33.916 67.396 34.164 70.2 ; 
      RECT 33.86 68.634 34.164 69.248 ; 
      RECT 33.916 65.826 34.02 70.2 ; 
      RECT 33.916 66.31 34.076 67.268 ; 
      RECT 33.916 65.826 34.164 66.182 ; 
      RECT 32.728 67.628 33.552 70.2 ; 
      RECT 33.448 65.826 33.552 70.2 ; 
      RECT 32.728 68.736 33.608 69.768 ; 
      RECT 32.728 65.826 33.12 70.2 ; 
      RECT 31.06 65.826 31.392 70.2 ; 
      RECT 31.06 66.18 31.448 69.922 ; 
      RECT 65.776 65.826 66.116 70.2 ; 
      RECT 65.2 65.826 65.304 70.2 ; 
      RECT 64.768 65.826 64.872 70.2 ; 
      RECT 64.336 65.826 64.44 70.2 ; 
      RECT 63.904 65.826 64.008 70.2 ; 
      RECT 63.472 65.826 63.576 70.2 ; 
      RECT 63.04 65.826 63.144 70.2 ; 
      RECT 62.608 65.826 62.712 70.2 ; 
      RECT 62.176 65.826 62.28 70.2 ; 
      RECT 61.744 65.826 61.848 70.2 ; 
      RECT 61.312 65.826 61.416 70.2 ; 
      RECT 60.88 65.826 60.984 70.2 ; 
      RECT 60.448 65.826 60.552 70.2 ; 
      RECT 60.016 65.826 60.12 70.2 ; 
      RECT 59.584 65.826 59.688 70.2 ; 
      RECT 59.152 65.826 59.256 70.2 ; 
      RECT 58.72 65.826 58.824 70.2 ; 
      RECT 58.288 65.826 58.392 70.2 ; 
      RECT 57.856 65.826 57.96 70.2 ; 
      RECT 57.424 65.826 57.528 70.2 ; 
      RECT 56.992 65.826 57.096 70.2 ; 
      RECT 56.56 65.826 56.664 70.2 ; 
      RECT 56.128 65.826 56.232 70.2 ; 
      RECT 55.696 65.826 55.8 70.2 ; 
      RECT 55.264 65.826 55.368 70.2 ; 
      RECT 54.832 65.826 54.936 70.2 ; 
      RECT 54.4 65.826 54.504 70.2 ; 
      RECT 53.968 65.826 54.072 70.2 ; 
      RECT 53.536 65.826 53.64 70.2 ; 
      RECT 53.104 65.826 53.208 70.2 ; 
      RECT 52.672 65.826 52.776 70.2 ; 
      RECT 52.24 65.826 52.344 70.2 ; 
      RECT 51.808 65.826 51.912 70.2 ; 
      RECT 51.376 65.826 51.48 70.2 ; 
      RECT 50.944 65.826 51.048 70.2 ; 
      RECT 50.512 65.826 50.616 70.2 ; 
      RECT 50.08 65.826 50.184 70.2 ; 
      RECT 49.648 65.826 49.752 70.2 ; 
      RECT 49.216 65.826 49.32 70.2 ; 
      RECT 48.784 65.826 48.888 70.2 ; 
      RECT 48.352 65.826 48.456 70.2 ; 
      RECT 47.92 65.826 48.024 70.2 ; 
      RECT 47.488 65.826 47.592 70.2 ; 
      RECT 47.056 65.826 47.16 70.2 ; 
      RECT 46.624 65.826 46.728 70.2 ; 
      RECT 46.192 65.826 46.296 70.2 ; 
      RECT 45.76 65.826 45.864 70.2 ; 
      RECT 45.328 65.826 45.432 70.2 ; 
      RECT 44.896 65.826 45 70.2 ; 
      RECT 44.464 65.826 44.568 70.2 ; 
      RECT 44.032 65.826 44.136 70.2 ; 
      RECT 43.6 65.826 43.704 70.2 ; 
      RECT 43.168 65.826 43.272 70.2 ; 
      RECT 42.736 65.826 42.84 70.2 ; 
      RECT 42.304 65.826 42.408 70.2 ; 
      RECT 41.872 65.826 41.976 70.2 ; 
      RECT 41.44 65.826 41.544 70.2 ; 
      RECT 41.008 65.826 41.112 70.2 ; 
      RECT 40.576 65.826 40.68 70.2 ; 
      RECT 40.144 65.826 40.248 70.2 ; 
      RECT 39.712 65.826 39.816 70.2 ; 
      RECT 39.28 65.826 39.384 70.2 ; 
      RECT 38.848 65.826 38.952 70.2 ; 
      RECT 38.416 65.826 38.52 70.2 ; 
      RECT 37.984 65.826 38.088 70.2 ; 
      RECT 37.552 65.826 37.656 70.2 ; 
      RECT 36.7 65.826 37.008 70.2 ; 
      RECT 29.128 65.826 29.436 70.2 ; 
      RECT 28.48 65.826 28.584 70.2 ; 
      RECT 28.048 65.826 28.152 70.2 ; 
      RECT 27.616 65.826 27.72 70.2 ; 
      RECT 27.184 65.826 27.288 70.2 ; 
      RECT 26.752 65.826 26.856 70.2 ; 
      RECT 26.32 65.826 26.424 70.2 ; 
      RECT 25.888 65.826 25.992 70.2 ; 
      RECT 25.456 65.826 25.56 70.2 ; 
      RECT 25.024 65.826 25.128 70.2 ; 
      RECT 24.592 65.826 24.696 70.2 ; 
      RECT 24.16 65.826 24.264 70.2 ; 
      RECT 23.728 65.826 23.832 70.2 ; 
      RECT 23.296 65.826 23.4 70.2 ; 
      RECT 22.864 65.826 22.968 70.2 ; 
      RECT 22.432 65.826 22.536 70.2 ; 
      RECT 22 65.826 22.104 70.2 ; 
      RECT 21.568 65.826 21.672 70.2 ; 
      RECT 21.136 65.826 21.24 70.2 ; 
      RECT 20.704 65.826 20.808 70.2 ; 
      RECT 20.272 65.826 20.376 70.2 ; 
      RECT 19.84 65.826 19.944 70.2 ; 
      RECT 19.408 65.826 19.512 70.2 ; 
      RECT 18.976 65.826 19.08 70.2 ; 
      RECT 18.544 65.826 18.648 70.2 ; 
      RECT 18.112 65.826 18.216 70.2 ; 
      RECT 17.68 65.826 17.784 70.2 ; 
      RECT 17.248 65.826 17.352 70.2 ; 
      RECT 16.816 65.826 16.92 70.2 ; 
      RECT 16.384 65.826 16.488 70.2 ; 
      RECT 15.952 65.826 16.056 70.2 ; 
      RECT 15.52 65.826 15.624 70.2 ; 
      RECT 15.088 65.826 15.192 70.2 ; 
      RECT 14.656 65.826 14.76 70.2 ; 
      RECT 14.224 65.826 14.328 70.2 ; 
      RECT 13.792 65.826 13.896 70.2 ; 
      RECT 13.36 65.826 13.464 70.2 ; 
      RECT 12.928 65.826 13.032 70.2 ; 
      RECT 12.496 65.826 12.6 70.2 ; 
      RECT 12.064 65.826 12.168 70.2 ; 
      RECT 11.632 65.826 11.736 70.2 ; 
      RECT 11.2 65.826 11.304 70.2 ; 
      RECT 10.768 65.826 10.872 70.2 ; 
      RECT 10.336 65.826 10.44 70.2 ; 
      RECT 9.904 65.826 10.008 70.2 ; 
      RECT 9.472 65.826 9.576 70.2 ; 
      RECT 9.04 65.826 9.144 70.2 ; 
      RECT 8.608 65.826 8.712 70.2 ; 
      RECT 8.176 65.826 8.28 70.2 ; 
      RECT 7.744 65.826 7.848 70.2 ; 
      RECT 7.312 65.826 7.416 70.2 ; 
      RECT 6.88 65.826 6.984 70.2 ; 
      RECT 6.448 65.826 6.552 70.2 ; 
      RECT 6.016 65.826 6.12 70.2 ; 
      RECT 5.584 65.826 5.688 70.2 ; 
      RECT 5.152 65.826 5.256 70.2 ; 
      RECT 4.72 65.826 4.824 70.2 ; 
      RECT 4.288 65.826 4.392 70.2 ; 
      RECT 3.856 65.826 3.96 70.2 ; 
      RECT 3.424 65.826 3.528 70.2 ; 
      RECT 2.992 65.826 3.096 70.2 ; 
      RECT 2.56 65.826 2.664 70.2 ; 
      RECT 2.128 65.826 2.232 70.2 ; 
      RECT 1.696 65.826 1.8 70.2 ; 
      RECT 1.264 65.826 1.368 70.2 ; 
      RECT 0.832 65.826 0.936 70.2 ; 
      RECT 0.02 65.826 0.36 70.2 ; 
      RECT 34.564 70.146 35.076 74.52 ; 
      RECT 34.508 72.808 35.076 74.098 ; 
      RECT 33.916 71.716 34.164 74.52 ; 
      RECT 33.86 72.954 34.164 73.568 ; 
      RECT 33.916 70.146 34.02 74.52 ; 
      RECT 33.916 70.63 34.076 71.588 ; 
      RECT 33.916 70.146 34.164 70.502 ; 
      RECT 32.728 71.948 33.552 74.52 ; 
      RECT 33.448 70.146 33.552 74.52 ; 
      RECT 32.728 73.056 33.608 74.088 ; 
      RECT 32.728 70.146 33.12 74.52 ; 
      RECT 31.06 70.146 31.392 74.52 ; 
      RECT 31.06 70.5 31.448 74.242 ; 
      RECT 65.776 70.146 66.116 74.52 ; 
      RECT 65.2 70.146 65.304 74.52 ; 
      RECT 64.768 70.146 64.872 74.52 ; 
      RECT 64.336 70.146 64.44 74.52 ; 
      RECT 63.904 70.146 64.008 74.52 ; 
      RECT 63.472 70.146 63.576 74.52 ; 
      RECT 63.04 70.146 63.144 74.52 ; 
      RECT 62.608 70.146 62.712 74.52 ; 
      RECT 62.176 70.146 62.28 74.52 ; 
      RECT 61.744 70.146 61.848 74.52 ; 
      RECT 61.312 70.146 61.416 74.52 ; 
      RECT 60.88 70.146 60.984 74.52 ; 
      RECT 60.448 70.146 60.552 74.52 ; 
      RECT 60.016 70.146 60.12 74.52 ; 
      RECT 59.584 70.146 59.688 74.52 ; 
      RECT 59.152 70.146 59.256 74.52 ; 
      RECT 58.72 70.146 58.824 74.52 ; 
      RECT 58.288 70.146 58.392 74.52 ; 
      RECT 57.856 70.146 57.96 74.52 ; 
      RECT 57.424 70.146 57.528 74.52 ; 
      RECT 56.992 70.146 57.096 74.52 ; 
      RECT 56.56 70.146 56.664 74.52 ; 
      RECT 56.128 70.146 56.232 74.52 ; 
      RECT 55.696 70.146 55.8 74.52 ; 
      RECT 55.264 70.146 55.368 74.52 ; 
      RECT 54.832 70.146 54.936 74.52 ; 
      RECT 54.4 70.146 54.504 74.52 ; 
      RECT 53.968 70.146 54.072 74.52 ; 
      RECT 53.536 70.146 53.64 74.52 ; 
      RECT 53.104 70.146 53.208 74.52 ; 
      RECT 52.672 70.146 52.776 74.52 ; 
      RECT 52.24 70.146 52.344 74.52 ; 
      RECT 51.808 70.146 51.912 74.52 ; 
      RECT 51.376 70.146 51.48 74.52 ; 
      RECT 50.944 70.146 51.048 74.52 ; 
      RECT 50.512 70.146 50.616 74.52 ; 
      RECT 50.08 70.146 50.184 74.52 ; 
      RECT 49.648 70.146 49.752 74.52 ; 
      RECT 49.216 70.146 49.32 74.52 ; 
      RECT 48.784 70.146 48.888 74.52 ; 
      RECT 48.352 70.146 48.456 74.52 ; 
      RECT 47.92 70.146 48.024 74.52 ; 
      RECT 47.488 70.146 47.592 74.52 ; 
      RECT 47.056 70.146 47.16 74.52 ; 
      RECT 46.624 70.146 46.728 74.52 ; 
      RECT 46.192 70.146 46.296 74.52 ; 
      RECT 45.76 70.146 45.864 74.52 ; 
      RECT 45.328 70.146 45.432 74.52 ; 
      RECT 44.896 70.146 45 74.52 ; 
      RECT 44.464 70.146 44.568 74.52 ; 
      RECT 44.032 70.146 44.136 74.52 ; 
      RECT 43.6 70.146 43.704 74.52 ; 
      RECT 43.168 70.146 43.272 74.52 ; 
      RECT 42.736 70.146 42.84 74.52 ; 
      RECT 42.304 70.146 42.408 74.52 ; 
      RECT 41.872 70.146 41.976 74.52 ; 
      RECT 41.44 70.146 41.544 74.52 ; 
      RECT 41.008 70.146 41.112 74.52 ; 
      RECT 40.576 70.146 40.68 74.52 ; 
      RECT 40.144 70.146 40.248 74.52 ; 
      RECT 39.712 70.146 39.816 74.52 ; 
      RECT 39.28 70.146 39.384 74.52 ; 
      RECT 38.848 70.146 38.952 74.52 ; 
      RECT 38.416 70.146 38.52 74.52 ; 
      RECT 37.984 70.146 38.088 74.52 ; 
      RECT 37.552 70.146 37.656 74.52 ; 
      RECT 36.7 70.146 37.008 74.52 ; 
      RECT 29.128 70.146 29.436 74.52 ; 
      RECT 28.48 70.146 28.584 74.52 ; 
      RECT 28.048 70.146 28.152 74.52 ; 
      RECT 27.616 70.146 27.72 74.52 ; 
      RECT 27.184 70.146 27.288 74.52 ; 
      RECT 26.752 70.146 26.856 74.52 ; 
      RECT 26.32 70.146 26.424 74.52 ; 
      RECT 25.888 70.146 25.992 74.52 ; 
      RECT 25.456 70.146 25.56 74.52 ; 
      RECT 25.024 70.146 25.128 74.52 ; 
      RECT 24.592 70.146 24.696 74.52 ; 
      RECT 24.16 70.146 24.264 74.52 ; 
      RECT 23.728 70.146 23.832 74.52 ; 
      RECT 23.296 70.146 23.4 74.52 ; 
      RECT 22.864 70.146 22.968 74.52 ; 
      RECT 22.432 70.146 22.536 74.52 ; 
      RECT 22 70.146 22.104 74.52 ; 
      RECT 21.568 70.146 21.672 74.52 ; 
      RECT 21.136 70.146 21.24 74.52 ; 
      RECT 20.704 70.146 20.808 74.52 ; 
      RECT 20.272 70.146 20.376 74.52 ; 
      RECT 19.84 70.146 19.944 74.52 ; 
      RECT 19.408 70.146 19.512 74.52 ; 
      RECT 18.976 70.146 19.08 74.52 ; 
      RECT 18.544 70.146 18.648 74.52 ; 
      RECT 18.112 70.146 18.216 74.52 ; 
      RECT 17.68 70.146 17.784 74.52 ; 
      RECT 17.248 70.146 17.352 74.52 ; 
      RECT 16.816 70.146 16.92 74.52 ; 
      RECT 16.384 70.146 16.488 74.52 ; 
      RECT 15.952 70.146 16.056 74.52 ; 
      RECT 15.52 70.146 15.624 74.52 ; 
      RECT 15.088 70.146 15.192 74.52 ; 
      RECT 14.656 70.146 14.76 74.52 ; 
      RECT 14.224 70.146 14.328 74.52 ; 
      RECT 13.792 70.146 13.896 74.52 ; 
      RECT 13.36 70.146 13.464 74.52 ; 
      RECT 12.928 70.146 13.032 74.52 ; 
      RECT 12.496 70.146 12.6 74.52 ; 
      RECT 12.064 70.146 12.168 74.52 ; 
      RECT 11.632 70.146 11.736 74.52 ; 
      RECT 11.2 70.146 11.304 74.52 ; 
      RECT 10.768 70.146 10.872 74.52 ; 
      RECT 10.336 70.146 10.44 74.52 ; 
      RECT 9.904 70.146 10.008 74.52 ; 
      RECT 9.472 70.146 9.576 74.52 ; 
      RECT 9.04 70.146 9.144 74.52 ; 
      RECT 8.608 70.146 8.712 74.52 ; 
      RECT 8.176 70.146 8.28 74.52 ; 
      RECT 7.744 70.146 7.848 74.52 ; 
      RECT 7.312 70.146 7.416 74.52 ; 
      RECT 6.88 70.146 6.984 74.52 ; 
      RECT 6.448 70.146 6.552 74.52 ; 
      RECT 6.016 70.146 6.12 74.52 ; 
      RECT 5.584 70.146 5.688 74.52 ; 
      RECT 5.152 70.146 5.256 74.52 ; 
      RECT 4.72 70.146 4.824 74.52 ; 
      RECT 4.288 70.146 4.392 74.52 ; 
      RECT 3.856 70.146 3.96 74.52 ; 
      RECT 3.424 70.146 3.528 74.52 ; 
      RECT 2.992 70.146 3.096 74.52 ; 
      RECT 2.56 70.146 2.664 74.52 ; 
      RECT 2.128 70.146 2.232 74.52 ; 
      RECT 1.696 70.146 1.8 74.52 ; 
      RECT 1.264 70.146 1.368 74.52 ; 
      RECT 0.832 70.146 0.936 74.52 ; 
      RECT 0.02 70.146 0.36 74.52 ; 
      RECT 34.564 74.466 35.076 78.84 ; 
      RECT 34.508 77.128 35.076 78.418 ; 
      RECT 33.916 76.036 34.164 78.84 ; 
      RECT 33.86 77.274 34.164 77.888 ; 
      RECT 33.916 74.466 34.02 78.84 ; 
      RECT 33.916 74.95 34.076 75.908 ; 
      RECT 33.916 74.466 34.164 74.822 ; 
      RECT 32.728 76.268 33.552 78.84 ; 
      RECT 33.448 74.466 33.552 78.84 ; 
      RECT 32.728 77.376 33.608 78.408 ; 
      RECT 32.728 74.466 33.12 78.84 ; 
      RECT 31.06 74.466 31.392 78.84 ; 
      RECT 31.06 74.82 31.448 78.562 ; 
      RECT 65.776 74.466 66.116 78.84 ; 
      RECT 65.2 74.466 65.304 78.84 ; 
      RECT 64.768 74.466 64.872 78.84 ; 
      RECT 64.336 74.466 64.44 78.84 ; 
      RECT 63.904 74.466 64.008 78.84 ; 
      RECT 63.472 74.466 63.576 78.84 ; 
      RECT 63.04 74.466 63.144 78.84 ; 
      RECT 62.608 74.466 62.712 78.84 ; 
      RECT 62.176 74.466 62.28 78.84 ; 
      RECT 61.744 74.466 61.848 78.84 ; 
      RECT 61.312 74.466 61.416 78.84 ; 
      RECT 60.88 74.466 60.984 78.84 ; 
      RECT 60.448 74.466 60.552 78.84 ; 
      RECT 60.016 74.466 60.12 78.84 ; 
      RECT 59.584 74.466 59.688 78.84 ; 
      RECT 59.152 74.466 59.256 78.84 ; 
      RECT 58.72 74.466 58.824 78.84 ; 
      RECT 58.288 74.466 58.392 78.84 ; 
      RECT 57.856 74.466 57.96 78.84 ; 
      RECT 57.424 74.466 57.528 78.84 ; 
      RECT 56.992 74.466 57.096 78.84 ; 
      RECT 56.56 74.466 56.664 78.84 ; 
      RECT 56.128 74.466 56.232 78.84 ; 
      RECT 55.696 74.466 55.8 78.84 ; 
      RECT 55.264 74.466 55.368 78.84 ; 
      RECT 54.832 74.466 54.936 78.84 ; 
      RECT 54.4 74.466 54.504 78.84 ; 
      RECT 53.968 74.466 54.072 78.84 ; 
      RECT 53.536 74.466 53.64 78.84 ; 
      RECT 53.104 74.466 53.208 78.84 ; 
      RECT 52.672 74.466 52.776 78.84 ; 
      RECT 52.24 74.466 52.344 78.84 ; 
      RECT 51.808 74.466 51.912 78.84 ; 
      RECT 51.376 74.466 51.48 78.84 ; 
      RECT 50.944 74.466 51.048 78.84 ; 
      RECT 50.512 74.466 50.616 78.84 ; 
      RECT 50.08 74.466 50.184 78.84 ; 
      RECT 49.648 74.466 49.752 78.84 ; 
      RECT 49.216 74.466 49.32 78.84 ; 
      RECT 48.784 74.466 48.888 78.84 ; 
      RECT 48.352 74.466 48.456 78.84 ; 
      RECT 47.92 74.466 48.024 78.84 ; 
      RECT 47.488 74.466 47.592 78.84 ; 
      RECT 47.056 74.466 47.16 78.84 ; 
      RECT 46.624 74.466 46.728 78.84 ; 
      RECT 46.192 74.466 46.296 78.84 ; 
      RECT 45.76 74.466 45.864 78.84 ; 
      RECT 45.328 74.466 45.432 78.84 ; 
      RECT 44.896 74.466 45 78.84 ; 
      RECT 44.464 74.466 44.568 78.84 ; 
      RECT 44.032 74.466 44.136 78.84 ; 
      RECT 43.6 74.466 43.704 78.84 ; 
      RECT 43.168 74.466 43.272 78.84 ; 
      RECT 42.736 74.466 42.84 78.84 ; 
      RECT 42.304 74.466 42.408 78.84 ; 
      RECT 41.872 74.466 41.976 78.84 ; 
      RECT 41.44 74.466 41.544 78.84 ; 
      RECT 41.008 74.466 41.112 78.84 ; 
      RECT 40.576 74.466 40.68 78.84 ; 
      RECT 40.144 74.466 40.248 78.84 ; 
      RECT 39.712 74.466 39.816 78.84 ; 
      RECT 39.28 74.466 39.384 78.84 ; 
      RECT 38.848 74.466 38.952 78.84 ; 
      RECT 38.416 74.466 38.52 78.84 ; 
      RECT 37.984 74.466 38.088 78.84 ; 
      RECT 37.552 74.466 37.656 78.84 ; 
      RECT 36.7 74.466 37.008 78.84 ; 
      RECT 29.128 74.466 29.436 78.84 ; 
      RECT 28.48 74.466 28.584 78.84 ; 
      RECT 28.048 74.466 28.152 78.84 ; 
      RECT 27.616 74.466 27.72 78.84 ; 
      RECT 27.184 74.466 27.288 78.84 ; 
      RECT 26.752 74.466 26.856 78.84 ; 
      RECT 26.32 74.466 26.424 78.84 ; 
      RECT 25.888 74.466 25.992 78.84 ; 
      RECT 25.456 74.466 25.56 78.84 ; 
      RECT 25.024 74.466 25.128 78.84 ; 
      RECT 24.592 74.466 24.696 78.84 ; 
      RECT 24.16 74.466 24.264 78.84 ; 
      RECT 23.728 74.466 23.832 78.84 ; 
      RECT 23.296 74.466 23.4 78.84 ; 
      RECT 22.864 74.466 22.968 78.84 ; 
      RECT 22.432 74.466 22.536 78.84 ; 
      RECT 22 74.466 22.104 78.84 ; 
      RECT 21.568 74.466 21.672 78.84 ; 
      RECT 21.136 74.466 21.24 78.84 ; 
      RECT 20.704 74.466 20.808 78.84 ; 
      RECT 20.272 74.466 20.376 78.84 ; 
      RECT 19.84 74.466 19.944 78.84 ; 
      RECT 19.408 74.466 19.512 78.84 ; 
      RECT 18.976 74.466 19.08 78.84 ; 
      RECT 18.544 74.466 18.648 78.84 ; 
      RECT 18.112 74.466 18.216 78.84 ; 
      RECT 17.68 74.466 17.784 78.84 ; 
      RECT 17.248 74.466 17.352 78.84 ; 
      RECT 16.816 74.466 16.92 78.84 ; 
      RECT 16.384 74.466 16.488 78.84 ; 
      RECT 15.952 74.466 16.056 78.84 ; 
      RECT 15.52 74.466 15.624 78.84 ; 
      RECT 15.088 74.466 15.192 78.84 ; 
      RECT 14.656 74.466 14.76 78.84 ; 
      RECT 14.224 74.466 14.328 78.84 ; 
      RECT 13.792 74.466 13.896 78.84 ; 
      RECT 13.36 74.466 13.464 78.84 ; 
      RECT 12.928 74.466 13.032 78.84 ; 
      RECT 12.496 74.466 12.6 78.84 ; 
      RECT 12.064 74.466 12.168 78.84 ; 
      RECT 11.632 74.466 11.736 78.84 ; 
      RECT 11.2 74.466 11.304 78.84 ; 
      RECT 10.768 74.466 10.872 78.84 ; 
      RECT 10.336 74.466 10.44 78.84 ; 
      RECT 9.904 74.466 10.008 78.84 ; 
      RECT 9.472 74.466 9.576 78.84 ; 
      RECT 9.04 74.466 9.144 78.84 ; 
      RECT 8.608 74.466 8.712 78.84 ; 
      RECT 8.176 74.466 8.28 78.84 ; 
      RECT 7.744 74.466 7.848 78.84 ; 
      RECT 7.312 74.466 7.416 78.84 ; 
      RECT 6.88 74.466 6.984 78.84 ; 
      RECT 6.448 74.466 6.552 78.84 ; 
      RECT 6.016 74.466 6.12 78.84 ; 
      RECT 5.584 74.466 5.688 78.84 ; 
      RECT 5.152 74.466 5.256 78.84 ; 
      RECT 4.72 74.466 4.824 78.84 ; 
      RECT 4.288 74.466 4.392 78.84 ; 
      RECT 3.856 74.466 3.96 78.84 ; 
      RECT 3.424 74.466 3.528 78.84 ; 
      RECT 2.992 74.466 3.096 78.84 ; 
      RECT 2.56 74.466 2.664 78.84 ; 
      RECT 2.128 74.466 2.232 78.84 ; 
      RECT 1.696 74.466 1.8 78.84 ; 
      RECT 1.264 74.466 1.368 78.84 ; 
      RECT 0.832 74.466 0.936 78.84 ; 
      RECT 0.02 74.466 0.36 78.84 ; 
      RECT 34.564 78.786 35.076 83.16 ; 
      RECT 34.508 81.448 35.076 82.738 ; 
      RECT 33.916 80.356 34.164 83.16 ; 
      RECT 33.86 81.594 34.164 82.208 ; 
      RECT 33.916 78.786 34.02 83.16 ; 
      RECT 33.916 79.27 34.076 80.228 ; 
      RECT 33.916 78.786 34.164 79.142 ; 
      RECT 32.728 80.588 33.552 83.16 ; 
      RECT 33.448 78.786 33.552 83.16 ; 
      RECT 32.728 81.696 33.608 82.728 ; 
      RECT 32.728 78.786 33.12 83.16 ; 
      RECT 31.06 78.786 31.392 83.16 ; 
      RECT 31.06 79.14 31.448 82.882 ; 
      RECT 65.776 78.786 66.116 83.16 ; 
      RECT 65.2 78.786 65.304 83.16 ; 
      RECT 64.768 78.786 64.872 83.16 ; 
      RECT 64.336 78.786 64.44 83.16 ; 
      RECT 63.904 78.786 64.008 83.16 ; 
      RECT 63.472 78.786 63.576 83.16 ; 
      RECT 63.04 78.786 63.144 83.16 ; 
      RECT 62.608 78.786 62.712 83.16 ; 
      RECT 62.176 78.786 62.28 83.16 ; 
      RECT 61.744 78.786 61.848 83.16 ; 
      RECT 61.312 78.786 61.416 83.16 ; 
      RECT 60.88 78.786 60.984 83.16 ; 
      RECT 60.448 78.786 60.552 83.16 ; 
      RECT 60.016 78.786 60.12 83.16 ; 
      RECT 59.584 78.786 59.688 83.16 ; 
      RECT 59.152 78.786 59.256 83.16 ; 
      RECT 58.72 78.786 58.824 83.16 ; 
      RECT 58.288 78.786 58.392 83.16 ; 
      RECT 57.856 78.786 57.96 83.16 ; 
      RECT 57.424 78.786 57.528 83.16 ; 
      RECT 56.992 78.786 57.096 83.16 ; 
      RECT 56.56 78.786 56.664 83.16 ; 
      RECT 56.128 78.786 56.232 83.16 ; 
      RECT 55.696 78.786 55.8 83.16 ; 
      RECT 55.264 78.786 55.368 83.16 ; 
      RECT 54.832 78.786 54.936 83.16 ; 
      RECT 54.4 78.786 54.504 83.16 ; 
      RECT 53.968 78.786 54.072 83.16 ; 
      RECT 53.536 78.786 53.64 83.16 ; 
      RECT 53.104 78.786 53.208 83.16 ; 
      RECT 52.672 78.786 52.776 83.16 ; 
      RECT 52.24 78.786 52.344 83.16 ; 
      RECT 51.808 78.786 51.912 83.16 ; 
      RECT 51.376 78.786 51.48 83.16 ; 
      RECT 50.944 78.786 51.048 83.16 ; 
      RECT 50.512 78.786 50.616 83.16 ; 
      RECT 50.08 78.786 50.184 83.16 ; 
      RECT 49.648 78.786 49.752 83.16 ; 
      RECT 49.216 78.786 49.32 83.16 ; 
      RECT 48.784 78.786 48.888 83.16 ; 
      RECT 48.352 78.786 48.456 83.16 ; 
      RECT 47.92 78.786 48.024 83.16 ; 
      RECT 47.488 78.786 47.592 83.16 ; 
      RECT 47.056 78.786 47.16 83.16 ; 
      RECT 46.624 78.786 46.728 83.16 ; 
      RECT 46.192 78.786 46.296 83.16 ; 
      RECT 45.76 78.786 45.864 83.16 ; 
      RECT 45.328 78.786 45.432 83.16 ; 
      RECT 44.896 78.786 45 83.16 ; 
      RECT 44.464 78.786 44.568 83.16 ; 
      RECT 44.032 78.786 44.136 83.16 ; 
      RECT 43.6 78.786 43.704 83.16 ; 
      RECT 43.168 78.786 43.272 83.16 ; 
      RECT 42.736 78.786 42.84 83.16 ; 
      RECT 42.304 78.786 42.408 83.16 ; 
      RECT 41.872 78.786 41.976 83.16 ; 
      RECT 41.44 78.786 41.544 83.16 ; 
      RECT 41.008 78.786 41.112 83.16 ; 
      RECT 40.576 78.786 40.68 83.16 ; 
      RECT 40.144 78.786 40.248 83.16 ; 
      RECT 39.712 78.786 39.816 83.16 ; 
      RECT 39.28 78.786 39.384 83.16 ; 
      RECT 38.848 78.786 38.952 83.16 ; 
      RECT 38.416 78.786 38.52 83.16 ; 
      RECT 37.984 78.786 38.088 83.16 ; 
      RECT 37.552 78.786 37.656 83.16 ; 
      RECT 36.7 78.786 37.008 83.16 ; 
      RECT 29.128 78.786 29.436 83.16 ; 
      RECT 28.48 78.786 28.584 83.16 ; 
      RECT 28.048 78.786 28.152 83.16 ; 
      RECT 27.616 78.786 27.72 83.16 ; 
      RECT 27.184 78.786 27.288 83.16 ; 
      RECT 26.752 78.786 26.856 83.16 ; 
      RECT 26.32 78.786 26.424 83.16 ; 
      RECT 25.888 78.786 25.992 83.16 ; 
      RECT 25.456 78.786 25.56 83.16 ; 
      RECT 25.024 78.786 25.128 83.16 ; 
      RECT 24.592 78.786 24.696 83.16 ; 
      RECT 24.16 78.786 24.264 83.16 ; 
      RECT 23.728 78.786 23.832 83.16 ; 
      RECT 23.296 78.786 23.4 83.16 ; 
      RECT 22.864 78.786 22.968 83.16 ; 
      RECT 22.432 78.786 22.536 83.16 ; 
      RECT 22 78.786 22.104 83.16 ; 
      RECT 21.568 78.786 21.672 83.16 ; 
      RECT 21.136 78.786 21.24 83.16 ; 
      RECT 20.704 78.786 20.808 83.16 ; 
      RECT 20.272 78.786 20.376 83.16 ; 
      RECT 19.84 78.786 19.944 83.16 ; 
      RECT 19.408 78.786 19.512 83.16 ; 
      RECT 18.976 78.786 19.08 83.16 ; 
      RECT 18.544 78.786 18.648 83.16 ; 
      RECT 18.112 78.786 18.216 83.16 ; 
      RECT 17.68 78.786 17.784 83.16 ; 
      RECT 17.248 78.786 17.352 83.16 ; 
      RECT 16.816 78.786 16.92 83.16 ; 
      RECT 16.384 78.786 16.488 83.16 ; 
      RECT 15.952 78.786 16.056 83.16 ; 
      RECT 15.52 78.786 15.624 83.16 ; 
      RECT 15.088 78.786 15.192 83.16 ; 
      RECT 14.656 78.786 14.76 83.16 ; 
      RECT 14.224 78.786 14.328 83.16 ; 
      RECT 13.792 78.786 13.896 83.16 ; 
      RECT 13.36 78.786 13.464 83.16 ; 
      RECT 12.928 78.786 13.032 83.16 ; 
      RECT 12.496 78.786 12.6 83.16 ; 
      RECT 12.064 78.786 12.168 83.16 ; 
      RECT 11.632 78.786 11.736 83.16 ; 
      RECT 11.2 78.786 11.304 83.16 ; 
      RECT 10.768 78.786 10.872 83.16 ; 
      RECT 10.336 78.786 10.44 83.16 ; 
      RECT 9.904 78.786 10.008 83.16 ; 
      RECT 9.472 78.786 9.576 83.16 ; 
      RECT 9.04 78.786 9.144 83.16 ; 
      RECT 8.608 78.786 8.712 83.16 ; 
      RECT 8.176 78.786 8.28 83.16 ; 
      RECT 7.744 78.786 7.848 83.16 ; 
      RECT 7.312 78.786 7.416 83.16 ; 
      RECT 6.88 78.786 6.984 83.16 ; 
      RECT 6.448 78.786 6.552 83.16 ; 
      RECT 6.016 78.786 6.12 83.16 ; 
      RECT 5.584 78.786 5.688 83.16 ; 
      RECT 5.152 78.786 5.256 83.16 ; 
      RECT 4.72 78.786 4.824 83.16 ; 
      RECT 4.288 78.786 4.392 83.16 ; 
      RECT 3.856 78.786 3.96 83.16 ; 
      RECT 3.424 78.786 3.528 83.16 ; 
      RECT 2.992 78.786 3.096 83.16 ; 
      RECT 2.56 78.786 2.664 83.16 ; 
      RECT 2.128 78.786 2.232 83.16 ; 
      RECT 1.696 78.786 1.8 83.16 ; 
      RECT 1.264 78.786 1.368 83.16 ; 
      RECT 0.832 78.786 0.936 83.16 ; 
      RECT 0.02 78.786 0.36 83.16 ; 
      RECT 34.564 83.106 35.076 87.48 ; 
      RECT 34.508 85.768 35.076 87.058 ; 
      RECT 33.916 84.676 34.164 87.48 ; 
      RECT 33.86 85.914 34.164 86.528 ; 
      RECT 33.916 83.106 34.02 87.48 ; 
      RECT 33.916 83.59 34.076 84.548 ; 
      RECT 33.916 83.106 34.164 83.462 ; 
      RECT 32.728 84.908 33.552 87.48 ; 
      RECT 33.448 83.106 33.552 87.48 ; 
      RECT 32.728 86.016 33.608 87.048 ; 
      RECT 32.728 83.106 33.12 87.48 ; 
      RECT 31.06 83.106 31.392 87.48 ; 
      RECT 31.06 83.46 31.448 87.202 ; 
      RECT 65.776 83.106 66.116 87.48 ; 
      RECT 65.2 83.106 65.304 87.48 ; 
      RECT 64.768 83.106 64.872 87.48 ; 
      RECT 64.336 83.106 64.44 87.48 ; 
      RECT 63.904 83.106 64.008 87.48 ; 
      RECT 63.472 83.106 63.576 87.48 ; 
      RECT 63.04 83.106 63.144 87.48 ; 
      RECT 62.608 83.106 62.712 87.48 ; 
      RECT 62.176 83.106 62.28 87.48 ; 
      RECT 61.744 83.106 61.848 87.48 ; 
      RECT 61.312 83.106 61.416 87.48 ; 
      RECT 60.88 83.106 60.984 87.48 ; 
      RECT 60.448 83.106 60.552 87.48 ; 
      RECT 60.016 83.106 60.12 87.48 ; 
      RECT 59.584 83.106 59.688 87.48 ; 
      RECT 59.152 83.106 59.256 87.48 ; 
      RECT 58.72 83.106 58.824 87.48 ; 
      RECT 58.288 83.106 58.392 87.48 ; 
      RECT 57.856 83.106 57.96 87.48 ; 
      RECT 57.424 83.106 57.528 87.48 ; 
      RECT 56.992 83.106 57.096 87.48 ; 
      RECT 56.56 83.106 56.664 87.48 ; 
      RECT 56.128 83.106 56.232 87.48 ; 
      RECT 55.696 83.106 55.8 87.48 ; 
      RECT 55.264 83.106 55.368 87.48 ; 
      RECT 54.832 83.106 54.936 87.48 ; 
      RECT 54.4 83.106 54.504 87.48 ; 
      RECT 53.968 83.106 54.072 87.48 ; 
      RECT 53.536 83.106 53.64 87.48 ; 
      RECT 53.104 83.106 53.208 87.48 ; 
      RECT 52.672 83.106 52.776 87.48 ; 
      RECT 52.24 83.106 52.344 87.48 ; 
      RECT 51.808 83.106 51.912 87.48 ; 
      RECT 51.376 83.106 51.48 87.48 ; 
      RECT 50.944 83.106 51.048 87.48 ; 
      RECT 50.512 83.106 50.616 87.48 ; 
      RECT 50.08 83.106 50.184 87.48 ; 
      RECT 49.648 83.106 49.752 87.48 ; 
      RECT 49.216 83.106 49.32 87.48 ; 
      RECT 48.784 83.106 48.888 87.48 ; 
      RECT 48.352 83.106 48.456 87.48 ; 
      RECT 47.92 83.106 48.024 87.48 ; 
      RECT 47.488 83.106 47.592 87.48 ; 
      RECT 47.056 83.106 47.16 87.48 ; 
      RECT 46.624 83.106 46.728 87.48 ; 
      RECT 46.192 83.106 46.296 87.48 ; 
      RECT 45.76 83.106 45.864 87.48 ; 
      RECT 45.328 83.106 45.432 87.48 ; 
      RECT 44.896 83.106 45 87.48 ; 
      RECT 44.464 83.106 44.568 87.48 ; 
      RECT 44.032 83.106 44.136 87.48 ; 
      RECT 43.6 83.106 43.704 87.48 ; 
      RECT 43.168 83.106 43.272 87.48 ; 
      RECT 42.736 83.106 42.84 87.48 ; 
      RECT 42.304 83.106 42.408 87.48 ; 
      RECT 41.872 83.106 41.976 87.48 ; 
      RECT 41.44 83.106 41.544 87.48 ; 
      RECT 41.008 83.106 41.112 87.48 ; 
      RECT 40.576 83.106 40.68 87.48 ; 
      RECT 40.144 83.106 40.248 87.48 ; 
      RECT 39.712 83.106 39.816 87.48 ; 
      RECT 39.28 83.106 39.384 87.48 ; 
      RECT 38.848 83.106 38.952 87.48 ; 
      RECT 38.416 83.106 38.52 87.48 ; 
      RECT 37.984 83.106 38.088 87.48 ; 
      RECT 37.552 83.106 37.656 87.48 ; 
      RECT 36.7 83.106 37.008 87.48 ; 
      RECT 29.128 83.106 29.436 87.48 ; 
      RECT 28.48 83.106 28.584 87.48 ; 
      RECT 28.048 83.106 28.152 87.48 ; 
      RECT 27.616 83.106 27.72 87.48 ; 
      RECT 27.184 83.106 27.288 87.48 ; 
      RECT 26.752 83.106 26.856 87.48 ; 
      RECT 26.32 83.106 26.424 87.48 ; 
      RECT 25.888 83.106 25.992 87.48 ; 
      RECT 25.456 83.106 25.56 87.48 ; 
      RECT 25.024 83.106 25.128 87.48 ; 
      RECT 24.592 83.106 24.696 87.48 ; 
      RECT 24.16 83.106 24.264 87.48 ; 
      RECT 23.728 83.106 23.832 87.48 ; 
      RECT 23.296 83.106 23.4 87.48 ; 
      RECT 22.864 83.106 22.968 87.48 ; 
      RECT 22.432 83.106 22.536 87.48 ; 
      RECT 22 83.106 22.104 87.48 ; 
      RECT 21.568 83.106 21.672 87.48 ; 
      RECT 21.136 83.106 21.24 87.48 ; 
      RECT 20.704 83.106 20.808 87.48 ; 
      RECT 20.272 83.106 20.376 87.48 ; 
      RECT 19.84 83.106 19.944 87.48 ; 
      RECT 19.408 83.106 19.512 87.48 ; 
      RECT 18.976 83.106 19.08 87.48 ; 
      RECT 18.544 83.106 18.648 87.48 ; 
      RECT 18.112 83.106 18.216 87.48 ; 
      RECT 17.68 83.106 17.784 87.48 ; 
      RECT 17.248 83.106 17.352 87.48 ; 
      RECT 16.816 83.106 16.92 87.48 ; 
      RECT 16.384 83.106 16.488 87.48 ; 
      RECT 15.952 83.106 16.056 87.48 ; 
      RECT 15.52 83.106 15.624 87.48 ; 
      RECT 15.088 83.106 15.192 87.48 ; 
      RECT 14.656 83.106 14.76 87.48 ; 
      RECT 14.224 83.106 14.328 87.48 ; 
      RECT 13.792 83.106 13.896 87.48 ; 
      RECT 13.36 83.106 13.464 87.48 ; 
      RECT 12.928 83.106 13.032 87.48 ; 
      RECT 12.496 83.106 12.6 87.48 ; 
      RECT 12.064 83.106 12.168 87.48 ; 
      RECT 11.632 83.106 11.736 87.48 ; 
      RECT 11.2 83.106 11.304 87.48 ; 
      RECT 10.768 83.106 10.872 87.48 ; 
      RECT 10.336 83.106 10.44 87.48 ; 
      RECT 9.904 83.106 10.008 87.48 ; 
      RECT 9.472 83.106 9.576 87.48 ; 
      RECT 9.04 83.106 9.144 87.48 ; 
      RECT 8.608 83.106 8.712 87.48 ; 
      RECT 8.176 83.106 8.28 87.48 ; 
      RECT 7.744 83.106 7.848 87.48 ; 
      RECT 7.312 83.106 7.416 87.48 ; 
      RECT 6.88 83.106 6.984 87.48 ; 
      RECT 6.448 83.106 6.552 87.48 ; 
      RECT 6.016 83.106 6.12 87.48 ; 
      RECT 5.584 83.106 5.688 87.48 ; 
      RECT 5.152 83.106 5.256 87.48 ; 
      RECT 4.72 83.106 4.824 87.48 ; 
      RECT 4.288 83.106 4.392 87.48 ; 
      RECT 3.856 83.106 3.96 87.48 ; 
      RECT 3.424 83.106 3.528 87.48 ; 
      RECT 2.992 83.106 3.096 87.48 ; 
      RECT 2.56 83.106 2.664 87.48 ; 
      RECT 2.128 83.106 2.232 87.48 ; 
      RECT 1.696 83.106 1.8 87.48 ; 
      RECT 1.264 83.106 1.368 87.48 ; 
      RECT 0.832 83.106 0.936 87.48 ; 
      RECT 0.02 83.106 0.36 87.48 ; 
      RECT 34.564 87.426 35.076 91.8 ; 
      RECT 34.508 90.088 35.076 91.378 ; 
      RECT 33.916 88.996 34.164 91.8 ; 
      RECT 33.86 90.234 34.164 90.848 ; 
      RECT 33.916 87.426 34.02 91.8 ; 
      RECT 33.916 87.91 34.076 88.868 ; 
      RECT 33.916 87.426 34.164 87.782 ; 
      RECT 32.728 89.228 33.552 91.8 ; 
      RECT 33.448 87.426 33.552 91.8 ; 
      RECT 32.728 90.336 33.608 91.368 ; 
      RECT 32.728 87.426 33.12 91.8 ; 
      RECT 31.06 87.426 31.392 91.8 ; 
      RECT 31.06 87.78 31.448 91.522 ; 
      RECT 65.776 87.426 66.116 91.8 ; 
      RECT 65.2 87.426 65.304 91.8 ; 
      RECT 64.768 87.426 64.872 91.8 ; 
      RECT 64.336 87.426 64.44 91.8 ; 
      RECT 63.904 87.426 64.008 91.8 ; 
      RECT 63.472 87.426 63.576 91.8 ; 
      RECT 63.04 87.426 63.144 91.8 ; 
      RECT 62.608 87.426 62.712 91.8 ; 
      RECT 62.176 87.426 62.28 91.8 ; 
      RECT 61.744 87.426 61.848 91.8 ; 
      RECT 61.312 87.426 61.416 91.8 ; 
      RECT 60.88 87.426 60.984 91.8 ; 
      RECT 60.448 87.426 60.552 91.8 ; 
      RECT 60.016 87.426 60.12 91.8 ; 
      RECT 59.584 87.426 59.688 91.8 ; 
      RECT 59.152 87.426 59.256 91.8 ; 
      RECT 58.72 87.426 58.824 91.8 ; 
      RECT 58.288 87.426 58.392 91.8 ; 
      RECT 57.856 87.426 57.96 91.8 ; 
      RECT 57.424 87.426 57.528 91.8 ; 
      RECT 56.992 87.426 57.096 91.8 ; 
      RECT 56.56 87.426 56.664 91.8 ; 
      RECT 56.128 87.426 56.232 91.8 ; 
      RECT 55.696 87.426 55.8 91.8 ; 
      RECT 55.264 87.426 55.368 91.8 ; 
      RECT 54.832 87.426 54.936 91.8 ; 
      RECT 54.4 87.426 54.504 91.8 ; 
      RECT 53.968 87.426 54.072 91.8 ; 
      RECT 53.536 87.426 53.64 91.8 ; 
      RECT 53.104 87.426 53.208 91.8 ; 
      RECT 52.672 87.426 52.776 91.8 ; 
      RECT 52.24 87.426 52.344 91.8 ; 
      RECT 51.808 87.426 51.912 91.8 ; 
      RECT 51.376 87.426 51.48 91.8 ; 
      RECT 50.944 87.426 51.048 91.8 ; 
      RECT 50.512 87.426 50.616 91.8 ; 
      RECT 50.08 87.426 50.184 91.8 ; 
      RECT 49.648 87.426 49.752 91.8 ; 
      RECT 49.216 87.426 49.32 91.8 ; 
      RECT 48.784 87.426 48.888 91.8 ; 
      RECT 48.352 87.426 48.456 91.8 ; 
      RECT 47.92 87.426 48.024 91.8 ; 
      RECT 47.488 87.426 47.592 91.8 ; 
      RECT 47.056 87.426 47.16 91.8 ; 
      RECT 46.624 87.426 46.728 91.8 ; 
      RECT 46.192 87.426 46.296 91.8 ; 
      RECT 45.76 87.426 45.864 91.8 ; 
      RECT 45.328 87.426 45.432 91.8 ; 
      RECT 44.896 87.426 45 91.8 ; 
      RECT 44.464 87.426 44.568 91.8 ; 
      RECT 44.032 87.426 44.136 91.8 ; 
      RECT 43.6 87.426 43.704 91.8 ; 
      RECT 43.168 87.426 43.272 91.8 ; 
      RECT 42.736 87.426 42.84 91.8 ; 
      RECT 42.304 87.426 42.408 91.8 ; 
      RECT 41.872 87.426 41.976 91.8 ; 
      RECT 41.44 87.426 41.544 91.8 ; 
      RECT 41.008 87.426 41.112 91.8 ; 
      RECT 40.576 87.426 40.68 91.8 ; 
      RECT 40.144 87.426 40.248 91.8 ; 
      RECT 39.712 87.426 39.816 91.8 ; 
      RECT 39.28 87.426 39.384 91.8 ; 
      RECT 38.848 87.426 38.952 91.8 ; 
      RECT 38.416 87.426 38.52 91.8 ; 
      RECT 37.984 87.426 38.088 91.8 ; 
      RECT 37.552 87.426 37.656 91.8 ; 
      RECT 36.7 87.426 37.008 91.8 ; 
      RECT 29.128 87.426 29.436 91.8 ; 
      RECT 28.48 87.426 28.584 91.8 ; 
      RECT 28.048 87.426 28.152 91.8 ; 
      RECT 27.616 87.426 27.72 91.8 ; 
      RECT 27.184 87.426 27.288 91.8 ; 
      RECT 26.752 87.426 26.856 91.8 ; 
      RECT 26.32 87.426 26.424 91.8 ; 
      RECT 25.888 87.426 25.992 91.8 ; 
      RECT 25.456 87.426 25.56 91.8 ; 
      RECT 25.024 87.426 25.128 91.8 ; 
      RECT 24.592 87.426 24.696 91.8 ; 
      RECT 24.16 87.426 24.264 91.8 ; 
      RECT 23.728 87.426 23.832 91.8 ; 
      RECT 23.296 87.426 23.4 91.8 ; 
      RECT 22.864 87.426 22.968 91.8 ; 
      RECT 22.432 87.426 22.536 91.8 ; 
      RECT 22 87.426 22.104 91.8 ; 
      RECT 21.568 87.426 21.672 91.8 ; 
      RECT 21.136 87.426 21.24 91.8 ; 
      RECT 20.704 87.426 20.808 91.8 ; 
      RECT 20.272 87.426 20.376 91.8 ; 
      RECT 19.84 87.426 19.944 91.8 ; 
      RECT 19.408 87.426 19.512 91.8 ; 
      RECT 18.976 87.426 19.08 91.8 ; 
      RECT 18.544 87.426 18.648 91.8 ; 
      RECT 18.112 87.426 18.216 91.8 ; 
      RECT 17.68 87.426 17.784 91.8 ; 
      RECT 17.248 87.426 17.352 91.8 ; 
      RECT 16.816 87.426 16.92 91.8 ; 
      RECT 16.384 87.426 16.488 91.8 ; 
      RECT 15.952 87.426 16.056 91.8 ; 
      RECT 15.52 87.426 15.624 91.8 ; 
      RECT 15.088 87.426 15.192 91.8 ; 
      RECT 14.656 87.426 14.76 91.8 ; 
      RECT 14.224 87.426 14.328 91.8 ; 
      RECT 13.792 87.426 13.896 91.8 ; 
      RECT 13.36 87.426 13.464 91.8 ; 
      RECT 12.928 87.426 13.032 91.8 ; 
      RECT 12.496 87.426 12.6 91.8 ; 
      RECT 12.064 87.426 12.168 91.8 ; 
      RECT 11.632 87.426 11.736 91.8 ; 
      RECT 11.2 87.426 11.304 91.8 ; 
      RECT 10.768 87.426 10.872 91.8 ; 
      RECT 10.336 87.426 10.44 91.8 ; 
      RECT 9.904 87.426 10.008 91.8 ; 
      RECT 9.472 87.426 9.576 91.8 ; 
      RECT 9.04 87.426 9.144 91.8 ; 
      RECT 8.608 87.426 8.712 91.8 ; 
      RECT 8.176 87.426 8.28 91.8 ; 
      RECT 7.744 87.426 7.848 91.8 ; 
      RECT 7.312 87.426 7.416 91.8 ; 
      RECT 6.88 87.426 6.984 91.8 ; 
      RECT 6.448 87.426 6.552 91.8 ; 
      RECT 6.016 87.426 6.12 91.8 ; 
      RECT 5.584 87.426 5.688 91.8 ; 
      RECT 5.152 87.426 5.256 91.8 ; 
      RECT 4.72 87.426 4.824 91.8 ; 
      RECT 4.288 87.426 4.392 91.8 ; 
      RECT 3.856 87.426 3.96 91.8 ; 
      RECT 3.424 87.426 3.528 91.8 ; 
      RECT 2.992 87.426 3.096 91.8 ; 
      RECT 2.56 87.426 2.664 91.8 ; 
      RECT 2.128 87.426 2.232 91.8 ; 
      RECT 1.696 87.426 1.8 91.8 ; 
      RECT 1.264 87.426 1.368 91.8 ; 
      RECT 0.832 87.426 0.936 91.8 ; 
      RECT 0.02 87.426 0.36 91.8 ; 
      RECT 34.564 91.746 35.076 96.12 ; 
      RECT 34.508 94.408 35.076 95.698 ; 
      RECT 33.916 93.316 34.164 96.12 ; 
      RECT 33.86 94.554 34.164 95.168 ; 
      RECT 33.916 91.746 34.02 96.12 ; 
      RECT 33.916 92.23 34.076 93.188 ; 
      RECT 33.916 91.746 34.164 92.102 ; 
      RECT 32.728 93.548 33.552 96.12 ; 
      RECT 33.448 91.746 33.552 96.12 ; 
      RECT 32.728 94.656 33.608 95.688 ; 
      RECT 32.728 91.746 33.12 96.12 ; 
      RECT 31.06 91.746 31.392 96.12 ; 
      RECT 31.06 92.1 31.448 95.842 ; 
      RECT 65.776 91.746 66.116 96.12 ; 
      RECT 65.2 91.746 65.304 96.12 ; 
      RECT 64.768 91.746 64.872 96.12 ; 
      RECT 64.336 91.746 64.44 96.12 ; 
      RECT 63.904 91.746 64.008 96.12 ; 
      RECT 63.472 91.746 63.576 96.12 ; 
      RECT 63.04 91.746 63.144 96.12 ; 
      RECT 62.608 91.746 62.712 96.12 ; 
      RECT 62.176 91.746 62.28 96.12 ; 
      RECT 61.744 91.746 61.848 96.12 ; 
      RECT 61.312 91.746 61.416 96.12 ; 
      RECT 60.88 91.746 60.984 96.12 ; 
      RECT 60.448 91.746 60.552 96.12 ; 
      RECT 60.016 91.746 60.12 96.12 ; 
      RECT 59.584 91.746 59.688 96.12 ; 
      RECT 59.152 91.746 59.256 96.12 ; 
      RECT 58.72 91.746 58.824 96.12 ; 
      RECT 58.288 91.746 58.392 96.12 ; 
      RECT 57.856 91.746 57.96 96.12 ; 
      RECT 57.424 91.746 57.528 96.12 ; 
      RECT 56.992 91.746 57.096 96.12 ; 
      RECT 56.56 91.746 56.664 96.12 ; 
      RECT 56.128 91.746 56.232 96.12 ; 
      RECT 55.696 91.746 55.8 96.12 ; 
      RECT 55.264 91.746 55.368 96.12 ; 
      RECT 54.832 91.746 54.936 96.12 ; 
      RECT 54.4 91.746 54.504 96.12 ; 
      RECT 53.968 91.746 54.072 96.12 ; 
      RECT 53.536 91.746 53.64 96.12 ; 
      RECT 53.104 91.746 53.208 96.12 ; 
      RECT 52.672 91.746 52.776 96.12 ; 
      RECT 52.24 91.746 52.344 96.12 ; 
      RECT 51.808 91.746 51.912 96.12 ; 
      RECT 51.376 91.746 51.48 96.12 ; 
      RECT 50.944 91.746 51.048 96.12 ; 
      RECT 50.512 91.746 50.616 96.12 ; 
      RECT 50.08 91.746 50.184 96.12 ; 
      RECT 49.648 91.746 49.752 96.12 ; 
      RECT 49.216 91.746 49.32 96.12 ; 
      RECT 48.784 91.746 48.888 96.12 ; 
      RECT 48.352 91.746 48.456 96.12 ; 
      RECT 47.92 91.746 48.024 96.12 ; 
      RECT 47.488 91.746 47.592 96.12 ; 
      RECT 47.056 91.746 47.16 96.12 ; 
      RECT 46.624 91.746 46.728 96.12 ; 
      RECT 46.192 91.746 46.296 96.12 ; 
      RECT 45.76 91.746 45.864 96.12 ; 
      RECT 45.328 91.746 45.432 96.12 ; 
      RECT 44.896 91.746 45 96.12 ; 
      RECT 44.464 91.746 44.568 96.12 ; 
      RECT 44.032 91.746 44.136 96.12 ; 
      RECT 43.6 91.746 43.704 96.12 ; 
      RECT 43.168 91.746 43.272 96.12 ; 
      RECT 42.736 91.746 42.84 96.12 ; 
      RECT 42.304 91.746 42.408 96.12 ; 
      RECT 41.872 91.746 41.976 96.12 ; 
      RECT 41.44 91.746 41.544 96.12 ; 
      RECT 41.008 91.746 41.112 96.12 ; 
      RECT 40.576 91.746 40.68 96.12 ; 
      RECT 40.144 91.746 40.248 96.12 ; 
      RECT 39.712 91.746 39.816 96.12 ; 
      RECT 39.28 91.746 39.384 96.12 ; 
      RECT 38.848 91.746 38.952 96.12 ; 
      RECT 38.416 91.746 38.52 96.12 ; 
      RECT 37.984 91.746 38.088 96.12 ; 
      RECT 37.552 91.746 37.656 96.12 ; 
      RECT 36.7 91.746 37.008 96.12 ; 
      RECT 29.128 91.746 29.436 96.12 ; 
      RECT 28.48 91.746 28.584 96.12 ; 
      RECT 28.048 91.746 28.152 96.12 ; 
      RECT 27.616 91.746 27.72 96.12 ; 
      RECT 27.184 91.746 27.288 96.12 ; 
      RECT 26.752 91.746 26.856 96.12 ; 
      RECT 26.32 91.746 26.424 96.12 ; 
      RECT 25.888 91.746 25.992 96.12 ; 
      RECT 25.456 91.746 25.56 96.12 ; 
      RECT 25.024 91.746 25.128 96.12 ; 
      RECT 24.592 91.746 24.696 96.12 ; 
      RECT 24.16 91.746 24.264 96.12 ; 
      RECT 23.728 91.746 23.832 96.12 ; 
      RECT 23.296 91.746 23.4 96.12 ; 
      RECT 22.864 91.746 22.968 96.12 ; 
      RECT 22.432 91.746 22.536 96.12 ; 
      RECT 22 91.746 22.104 96.12 ; 
      RECT 21.568 91.746 21.672 96.12 ; 
      RECT 21.136 91.746 21.24 96.12 ; 
      RECT 20.704 91.746 20.808 96.12 ; 
      RECT 20.272 91.746 20.376 96.12 ; 
      RECT 19.84 91.746 19.944 96.12 ; 
      RECT 19.408 91.746 19.512 96.12 ; 
      RECT 18.976 91.746 19.08 96.12 ; 
      RECT 18.544 91.746 18.648 96.12 ; 
      RECT 18.112 91.746 18.216 96.12 ; 
      RECT 17.68 91.746 17.784 96.12 ; 
      RECT 17.248 91.746 17.352 96.12 ; 
      RECT 16.816 91.746 16.92 96.12 ; 
      RECT 16.384 91.746 16.488 96.12 ; 
      RECT 15.952 91.746 16.056 96.12 ; 
      RECT 15.52 91.746 15.624 96.12 ; 
      RECT 15.088 91.746 15.192 96.12 ; 
      RECT 14.656 91.746 14.76 96.12 ; 
      RECT 14.224 91.746 14.328 96.12 ; 
      RECT 13.792 91.746 13.896 96.12 ; 
      RECT 13.36 91.746 13.464 96.12 ; 
      RECT 12.928 91.746 13.032 96.12 ; 
      RECT 12.496 91.746 12.6 96.12 ; 
      RECT 12.064 91.746 12.168 96.12 ; 
      RECT 11.632 91.746 11.736 96.12 ; 
      RECT 11.2 91.746 11.304 96.12 ; 
      RECT 10.768 91.746 10.872 96.12 ; 
      RECT 10.336 91.746 10.44 96.12 ; 
      RECT 9.904 91.746 10.008 96.12 ; 
      RECT 9.472 91.746 9.576 96.12 ; 
      RECT 9.04 91.746 9.144 96.12 ; 
      RECT 8.608 91.746 8.712 96.12 ; 
      RECT 8.176 91.746 8.28 96.12 ; 
      RECT 7.744 91.746 7.848 96.12 ; 
      RECT 7.312 91.746 7.416 96.12 ; 
      RECT 6.88 91.746 6.984 96.12 ; 
      RECT 6.448 91.746 6.552 96.12 ; 
      RECT 6.016 91.746 6.12 96.12 ; 
      RECT 5.584 91.746 5.688 96.12 ; 
      RECT 5.152 91.746 5.256 96.12 ; 
      RECT 4.72 91.746 4.824 96.12 ; 
      RECT 4.288 91.746 4.392 96.12 ; 
      RECT 3.856 91.746 3.96 96.12 ; 
      RECT 3.424 91.746 3.528 96.12 ; 
      RECT 2.992 91.746 3.096 96.12 ; 
      RECT 2.56 91.746 2.664 96.12 ; 
      RECT 2.128 91.746 2.232 96.12 ; 
      RECT 1.696 91.746 1.8 96.12 ; 
      RECT 1.264 91.746 1.368 96.12 ; 
      RECT 0.832 91.746 0.936 96.12 ; 
      RECT 0.02 91.746 0.36 96.12 ; 
      RECT 34.564 96.066 35.076 100.44 ; 
      RECT 34.508 98.728 35.076 100.018 ; 
      RECT 33.916 97.636 34.164 100.44 ; 
      RECT 33.86 98.874 34.164 99.488 ; 
      RECT 33.916 96.066 34.02 100.44 ; 
      RECT 33.916 96.55 34.076 97.508 ; 
      RECT 33.916 96.066 34.164 96.422 ; 
      RECT 32.728 97.868 33.552 100.44 ; 
      RECT 33.448 96.066 33.552 100.44 ; 
      RECT 32.728 98.976 33.608 100.008 ; 
      RECT 32.728 96.066 33.12 100.44 ; 
      RECT 31.06 96.066 31.392 100.44 ; 
      RECT 31.06 96.42 31.448 100.162 ; 
      RECT 65.776 96.066 66.116 100.44 ; 
      RECT 65.2 96.066 65.304 100.44 ; 
      RECT 64.768 96.066 64.872 100.44 ; 
      RECT 64.336 96.066 64.44 100.44 ; 
      RECT 63.904 96.066 64.008 100.44 ; 
      RECT 63.472 96.066 63.576 100.44 ; 
      RECT 63.04 96.066 63.144 100.44 ; 
      RECT 62.608 96.066 62.712 100.44 ; 
      RECT 62.176 96.066 62.28 100.44 ; 
      RECT 61.744 96.066 61.848 100.44 ; 
      RECT 61.312 96.066 61.416 100.44 ; 
      RECT 60.88 96.066 60.984 100.44 ; 
      RECT 60.448 96.066 60.552 100.44 ; 
      RECT 60.016 96.066 60.12 100.44 ; 
      RECT 59.584 96.066 59.688 100.44 ; 
      RECT 59.152 96.066 59.256 100.44 ; 
      RECT 58.72 96.066 58.824 100.44 ; 
      RECT 58.288 96.066 58.392 100.44 ; 
      RECT 57.856 96.066 57.96 100.44 ; 
      RECT 57.424 96.066 57.528 100.44 ; 
      RECT 56.992 96.066 57.096 100.44 ; 
      RECT 56.56 96.066 56.664 100.44 ; 
      RECT 56.128 96.066 56.232 100.44 ; 
      RECT 55.696 96.066 55.8 100.44 ; 
      RECT 55.264 96.066 55.368 100.44 ; 
      RECT 54.832 96.066 54.936 100.44 ; 
      RECT 54.4 96.066 54.504 100.44 ; 
      RECT 53.968 96.066 54.072 100.44 ; 
      RECT 53.536 96.066 53.64 100.44 ; 
      RECT 53.104 96.066 53.208 100.44 ; 
      RECT 52.672 96.066 52.776 100.44 ; 
      RECT 52.24 96.066 52.344 100.44 ; 
      RECT 51.808 96.066 51.912 100.44 ; 
      RECT 51.376 96.066 51.48 100.44 ; 
      RECT 50.944 96.066 51.048 100.44 ; 
      RECT 50.512 96.066 50.616 100.44 ; 
      RECT 50.08 96.066 50.184 100.44 ; 
      RECT 49.648 96.066 49.752 100.44 ; 
      RECT 49.216 96.066 49.32 100.44 ; 
      RECT 48.784 96.066 48.888 100.44 ; 
      RECT 48.352 96.066 48.456 100.44 ; 
      RECT 47.92 96.066 48.024 100.44 ; 
      RECT 47.488 96.066 47.592 100.44 ; 
      RECT 47.056 96.066 47.16 100.44 ; 
      RECT 46.624 96.066 46.728 100.44 ; 
      RECT 46.192 96.066 46.296 100.44 ; 
      RECT 45.76 96.066 45.864 100.44 ; 
      RECT 45.328 96.066 45.432 100.44 ; 
      RECT 44.896 96.066 45 100.44 ; 
      RECT 44.464 96.066 44.568 100.44 ; 
      RECT 44.032 96.066 44.136 100.44 ; 
      RECT 43.6 96.066 43.704 100.44 ; 
      RECT 43.168 96.066 43.272 100.44 ; 
      RECT 42.736 96.066 42.84 100.44 ; 
      RECT 42.304 96.066 42.408 100.44 ; 
      RECT 41.872 96.066 41.976 100.44 ; 
      RECT 41.44 96.066 41.544 100.44 ; 
      RECT 41.008 96.066 41.112 100.44 ; 
      RECT 40.576 96.066 40.68 100.44 ; 
      RECT 40.144 96.066 40.248 100.44 ; 
      RECT 39.712 96.066 39.816 100.44 ; 
      RECT 39.28 96.066 39.384 100.44 ; 
      RECT 38.848 96.066 38.952 100.44 ; 
      RECT 38.416 96.066 38.52 100.44 ; 
      RECT 37.984 96.066 38.088 100.44 ; 
      RECT 37.552 96.066 37.656 100.44 ; 
      RECT 36.7 96.066 37.008 100.44 ; 
      RECT 29.128 96.066 29.436 100.44 ; 
      RECT 28.48 96.066 28.584 100.44 ; 
      RECT 28.048 96.066 28.152 100.44 ; 
      RECT 27.616 96.066 27.72 100.44 ; 
      RECT 27.184 96.066 27.288 100.44 ; 
      RECT 26.752 96.066 26.856 100.44 ; 
      RECT 26.32 96.066 26.424 100.44 ; 
      RECT 25.888 96.066 25.992 100.44 ; 
      RECT 25.456 96.066 25.56 100.44 ; 
      RECT 25.024 96.066 25.128 100.44 ; 
      RECT 24.592 96.066 24.696 100.44 ; 
      RECT 24.16 96.066 24.264 100.44 ; 
      RECT 23.728 96.066 23.832 100.44 ; 
      RECT 23.296 96.066 23.4 100.44 ; 
      RECT 22.864 96.066 22.968 100.44 ; 
      RECT 22.432 96.066 22.536 100.44 ; 
      RECT 22 96.066 22.104 100.44 ; 
      RECT 21.568 96.066 21.672 100.44 ; 
      RECT 21.136 96.066 21.24 100.44 ; 
      RECT 20.704 96.066 20.808 100.44 ; 
      RECT 20.272 96.066 20.376 100.44 ; 
      RECT 19.84 96.066 19.944 100.44 ; 
      RECT 19.408 96.066 19.512 100.44 ; 
      RECT 18.976 96.066 19.08 100.44 ; 
      RECT 18.544 96.066 18.648 100.44 ; 
      RECT 18.112 96.066 18.216 100.44 ; 
      RECT 17.68 96.066 17.784 100.44 ; 
      RECT 17.248 96.066 17.352 100.44 ; 
      RECT 16.816 96.066 16.92 100.44 ; 
      RECT 16.384 96.066 16.488 100.44 ; 
      RECT 15.952 96.066 16.056 100.44 ; 
      RECT 15.52 96.066 15.624 100.44 ; 
      RECT 15.088 96.066 15.192 100.44 ; 
      RECT 14.656 96.066 14.76 100.44 ; 
      RECT 14.224 96.066 14.328 100.44 ; 
      RECT 13.792 96.066 13.896 100.44 ; 
      RECT 13.36 96.066 13.464 100.44 ; 
      RECT 12.928 96.066 13.032 100.44 ; 
      RECT 12.496 96.066 12.6 100.44 ; 
      RECT 12.064 96.066 12.168 100.44 ; 
      RECT 11.632 96.066 11.736 100.44 ; 
      RECT 11.2 96.066 11.304 100.44 ; 
      RECT 10.768 96.066 10.872 100.44 ; 
      RECT 10.336 96.066 10.44 100.44 ; 
      RECT 9.904 96.066 10.008 100.44 ; 
      RECT 9.472 96.066 9.576 100.44 ; 
      RECT 9.04 96.066 9.144 100.44 ; 
      RECT 8.608 96.066 8.712 100.44 ; 
      RECT 8.176 96.066 8.28 100.44 ; 
      RECT 7.744 96.066 7.848 100.44 ; 
      RECT 7.312 96.066 7.416 100.44 ; 
      RECT 6.88 96.066 6.984 100.44 ; 
      RECT 6.448 96.066 6.552 100.44 ; 
      RECT 6.016 96.066 6.12 100.44 ; 
      RECT 5.584 96.066 5.688 100.44 ; 
      RECT 5.152 96.066 5.256 100.44 ; 
      RECT 4.72 96.066 4.824 100.44 ; 
      RECT 4.288 96.066 4.392 100.44 ; 
      RECT 3.856 96.066 3.96 100.44 ; 
      RECT 3.424 96.066 3.528 100.44 ; 
      RECT 2.992 96.066 3.096 100.44 ; 
      RECT 2.56 96.066 2.664 100.44 ; 
      RECT 2.128 96.066 2.232 100.44 ; 
      RECT 1.696 96.066 1.8 100.44 ; 
      RECT 1.264 96.066 1.368 100.44 ; 
      RECT 0.832 96.066 0.936 100.44 ; 
      RECT 0.02 96.066 0.36 100.44 ; 
      RECT 34.564 100.386 35.076 104.76 ; 
      RECT 34.508 103.048 35.076 104.338 ; 
      RECT 33.916 101.956 34.164 104.76 ; 
      RECT 33.86 103.194 34.164 103.808 ; 
      RECT 33.916 100.386 34.02 104.76 ; 
      RECT 33.916 100.87 34.076 101.828 ; 
      RECT 33.916 100.386 34.164 100.742 ; 
      RECT 32.728 102.188 33.552 104.76 ; 
      RECT 33.448 100.386 33.552 104.76 ; 
      RECT 32.728 103.296 33.608 104.328 ; 
      RECT 32.728 100.386 33.12 104.76 ; 
      RECT 31.06 100.386 31.392 104.76 ; 
      RECT 31.06 100.74 31.448 104.482 ; 
      RECT 65.776 100.386 66.116 104.76 ; 
      RECT 65.2 100.386 65.304 104.76 ; 
      RECT 64.768 100.386 64.872 104.76 ; 
      RECT 64.336 100.386 64.44 104.76 ; 
      RECT 63.904 100.386 64.008 104.76 ; 
      RECT 63.472 100.386 63.576 104.76 ; 
      RECT 63.04 100.386 63.144 104.76 ; 
      RECT 62.608 100.386 62.712 104.76 ; 
      RECT 62.176 100.386 62.28 104.76 ; 
      RECT 61.744 100.386 61.848 104.76 ; 
      RECT 61.312 100.386 61.416 104.76 ; 
      RECT 60.88 100.386 60.984 104.76 ; 
      RECT 60.448 100.386 60.552 104.76 ; 
      RECT 60.016 100.386 60.12 104.76 ; 
      RECT 59.584 100.386 59.688 104.76 ; 
      RECT 59.152 100.386 59.256 104.76 ; 
      RECT 58.72 100.386 58.824 104.76 ; 
      RECT 58.288 100.386 58.392 104.76 ; 
      RECT 57.856 100.386 57.96 104.76 ; 
      RECT 57.424 100.386 57.528 104.76 ; 
      RECT 56.992 100.386 57.096 104.76 ; 
      RECT 56.56 100.386 56.664 104.76 ; 
      RECT 56.128 100.386 56.232 104.76 ; 
      RECT 55.696 100.386 55.8 104.76 ; 
      RECT 55.264 100.386 55.368 104.76 ; 
      RECT 54.832 100.386 54.936 104.76 ; 
      RECT 54.4 100.386 54.504 104.76 ; 
      RECT 53.968 100.386 54.072 104.76 ; 
      RECT 53.536 100.386 53.64 104.76 ; 
      RECT 53.104 100.386 53.208 104.76 ; 
      RECT 52.672 100.386 52.776 104.76 ; 
      RECT 52.24 100.386 52.344 104.76 ; 
      RECT 51.808 100.386 51.912 104.76 ; 
      RECT 51.376 100.386 51.48 104.76 ; 
      RECT 50.944 100.386 51.048 104.76 ; 
      RECT 50.512 100.386 50.616 104.76 ; 
      RECT 50.08 100.386 50.184 104.76 ; 
      RECT 49.648 100.386 49.752 104.76 ; 
      RECT 49.216 100.386 49.32 104.76 ; 
      RECT 48.784 100.386 48.888 104.76 ; 
      RECT 48.352 100.386 48.456 104.76 ; 
      RECT 47.92 100.386 48.024 104.76 ; 
      RECT 47.488 100.386 47.592 104.76 ; 
      RECT 47.056 100.386 47.16 104.76 ; 
      RECT 46.624 100.386 46.728 104.76 ; 
      RECT 46.192 100.386 46.296 104.76 ; 
      RECT 45.76 100.386 45.864 104.76 ; 
      RECT 45.328 100.386 45.432 104.76 ; 
      RECT 44.896 100.386 45 104.76 ; 
      RECT 44.464 100.386 44.568 104.76 ; 
      RECT 44.032 100.386 44.136 104.76 ; 
      RECT 43.6 100.386 43.704 104.76 ; 
      RECT 43.168 100.386 43.272 104.76 ; 
      RECT 42.736 100.386 42.84 104.76 ; 
      RECT 42.304 100.386 42.408 104.76 ; 
      RECT 41.872 100.386 41.976 104.76 ; 
      RECT 41.44 100.386 41.544 104.76 ; 
      RECT 41.008 100.386 41.112 104.76 ; 
      RECT 40.576 100.386 40.68 104.76 ; 
      RECT 40.144 100.386 40.248 104.76 ; 
      RECT 39.712 100.386 39.816 104.76 ; 
      RECT 39.28 100.386 39.384 104.76 ; 
      RECT 38.848 100.386 38.952 104.76 ; 
      RECT 38.416 100.386 38.52 104.76 ; 
      RECT 37.984 100.386 38.088 104.76 ; 
      RECT 37.552 100.386 37.656 104.76 ; 
      RECT 36.7 100.386 37.008 104.76 ; 
      RECT 29.128 100.386 29.436 104.76 ; 
      RECT 28.48 100.386 28.584 104.76 ; 
      RECT 28.048 100.386 28.152 104.76 ; 
      RECT 27.616 100.386 27.72 104.76 ; 
      RECT 27.184 100.386 27.288 104.76 ; 
      RECT 26.752 100.386 26.856 104.76 ; 
      RECT 26.32 100.386 26.424 104.76 ; 
      RECT 25.888 100.386 25.992 104.76 ; 
      RECT 25.456 100.386 25.56 104.76 ; 
      RECT 25.024 100.386 25.128 104.76 ; 
      RECT 24.592 100.386 24.696 104.76 ; 
      RECT 24.16 100.386 24.264 104.76 ; 
      RECT 23.728 100.386 23.832 104.76 ; 
      RECT 23.296 100.386 23.4 104.76 ; 
      RECT 22.864 100.386 22.968 104.76 ; 
      RECT 22.432 100.386 22.536 104.76 ; 
      RECT 22 100.386 22.104 104.76 ; 
      RECT 21.568 100.386 21.672 104.76 ; 
      RECT 21.136 100.386 21.24 104.76 ; 
      RECT 20.704 100.386 20.808 104.76 ; 
      RECT 20.272 100.386 20.376 104.76 ; 
      RECT 19.84 100.386 19.944 104.76 ; 
      RECT 19.408 100.386 19.512 104.76 ; 
      RECT 18.976 100.386 19.08 104.76 ; 
      RECT 18.544 100.386 18.648 104.76 ; 
      RECT 18.112 100.386 18.216 104.76 ; 
      RECT 17.68 100.386 17.784 104.76 ; 
      RECT 17.248 100.386 17.352 104.76 ; 
      RECT 16.816 100.386 16.92 104.76 ; 
      RECT 16.384 100.386 16.488 104.76 ; 
      RECT 15.952 100.386 16.056 104.76 ; 
      RECT 15.52 100.386 15.624 104.76 ; 
      RECT 15.088 100.386 15.192 104.76 ; 
      RECT 14.656 100.386 14.76 104.76 ; 
      RECT 14.224 100.386 14.328 104.76 ; 
      RECT 13.792 100.386 13.896 104.76 ; 
      RECT 13.36 100.386 13.464 104.76 ; 
      RECT 12.928 100.386 13.032 104.76 ; 
      RECT 12.496 100.386 12.6 104.76 ; 
      RECT 12.064 100.386 12.168 104.76 ; 
      RECT 11.632 100.386 11.736 104.76 ; 
      RECT 11.2 100.386 11.304 104.76 ; 
      RECT 10.768 100.386 10.872 104.76 ; 
      RECT 10.336 100.386 10.44 104.76 ; 
      RECT 9.904 100.386 10.008 104.76 ; 
      RECT 9.472 100.386 9.576 104.76 ; 
      RECT 9.04 100.386 9.144 104.76 ; 
      RECT 8.608 100.386 8.712 104.76 ; 
      RECT 8.176 100.386 8.28 104.76 ; 
      RECT 7.744 100.386 7.848 104.76 ; 
      RECT 7.312 100.386 7.416 104.76 ; 
      RECT 6.88 100.386 6.984 104.76 ; 
      RECT 6.448 100.386 6.552 104.76 ; 
      RECT 6.016 100.386 6.12 104.76 ; 
      RECT 5.584 100.386 5.688 104.76 ; 
      RECT 5.152 100.386 5.256 104.76 ; 
      RECT 4.72 100.386 4.824 104.76 ; 
      RECT 4.288 100.386 4.392 104.76 ; 
      RECT 3.856 100.386 3.96 104.76 ; 
      RECT 3.424 100.386 3.528 104.76 ; 
      RECT 2.992 100.386 3.096 104.76 ; 
      RECT 2.56 100.386 2.664 104.76 ; 
      RECT 2.128 100.386 2.232 104.76 ; 
      RECT 1.696 100.386 1.8 104.76 ; 
      RECT 1.264 100.386 1.368 104.76 ; 
      RECT 0.832 100.386 0.936 104.76 ; 
      RECT 0.02 100.386 0.36 104.76 ; 
      RECT 34.564 104.706 35.076 109.08 ; 
      RECT 34.508 107.368 35.076 108.658 ; 
      RECT 33.916 106.276 34.164 109.08 ; 
      RECT 33.86 107.514 34.164 108.128 ; 
      RECT 33.916 104.706 34.02 109.08 ; 
      RECT 33.916 105.19 34.076 106.148 ; 
      RECT 33.916 104.706 34.164 105.062 ; 
      RECT 32.728 106.508 33.552 109.08 ; 
      RECT 33.448 104.706 33.552 109.08 ; 
      RECT 32.728 107.616 33.608 108.648 ; 
      RECT 32.728 104.706 33.12 109.08 ; 
      RECT 31.06 104.706 31.392 109.08 ; 
      RECT 31.06 105.06 31.448 108.802 ; 
      RECT 65.776 104.706 66.116 109.08 ; 
      RECT 65.2 104.706 65.304 109.08 ; 
      RECT 64.768 104.706 64.872 109.08 ; 
      RECT 64.336 104.706 64.44 109.08 ; 
      RECT 63.904 104.706 64.008 109.08 ; 
      RECT 63.472 104.706 63.576 109.08 ; 
      RECT 63.04 104.706 63.144 109.08 ; 
      RECT 62.608 104.706 62.712 109.08 ; 
      RECT 62.176 104.706 62.28 109.08 ; 
      RECT 61.744 104.706 61.848 109.08 ; 
      RECT 61.312 104.706 61.416 109.08 ; 
      RECT 60.88 104.706 60.984 109.08 ; 
      RECT 60.448 104.706 60.552 109.08 ; 
      RECT 60.016 104.706 60.12 109.08 ; 
      RECT 59.584 104.706 59.688 109.08 ; 
      RECT 59.152 104.706 59.256 109.08 ; 
      RECT 58.72 104.706 58.824 109.08 ; 
      RECT 58.288 104.706 58.392 109.08 ; 
      RECT 57.856 104.706 57.96 109.08 ; 
      RECT 57.424 104.706 57.528 109.08 ; 
      RECT 56.992 104.706 57.096 109.08 ; 
      RECT 56.56 104.706 56.664 109.08 ; 
      RECT 56.128 104.706 56.232 109.08 ; 
      RECT 55.696 104.706 55.8 109.08 ; 
      RECT 55.264 104.706 55.368 109.08 ; 
      RECT 54.832 104.706 54.936 109.08 ; 
      RECT 54.4 104.706 54.504 109.08 ; 
      RECT 53.968 104.706 54.072 109.08 ; 
      RECT 53.536 104.706 53.64 109.08 ; 
      RECT 53.104 104.706 53.208 109.08 ; 
      RECT 52.672 104.706 52.776 109.08 ; 
      RECT 52.24 104.706 52.344 109.08 ; 
      RECT 51.808 104.706 51.912 109.08 ; 
      RECT 51.376 104.706 51.48 109.08 ; 
      RECT 50.944 104.706 51.048 109.08 ; 
      RECT 50.512 104.706 50.616 109.08 ; 
      RECT 50.08 104.706 50.184 109.08 ; 
      RECT 49.648 104.706 49.752 109.08 ; 
      RECT 49.216 104.706 49.32 109.08 ; 
      RECT 48.784 104.706 48.888 109.08 ; 
      RECT 48.352 104.706 48.456 109.08 ; 
      RECT 47.92 104.706 48.024 109.08 ; 
      RECT 47.488 104.706 47.592 109.08 ; 
      RECT 47.056 104.706 47.16 109.08 ; 
      RECT 46.624 104.706 46.728 109.08 ; 
      RECT 46.192 104.706 46.296 109.08 ; 
      RECT 45.76 104.706 45.864 109.08 ; 
      RECT 45.328 104.706 45.432 109.08 ; 
      RECT 44.896 104.706 45 109.08 ; 
      RECT 44.464 104.706 44.568 109.08 ; 
      RECT 44.032 104.706 44.136 109.08 ; 
      RECT 43.6 104.706 43.704 109.08 ; 
      RECT 43.168 104.706 43.272 109.08 ; 
      RECT 42.736 104.706 42.84 109.08 ; 
      RECT 42.304 104.706 42.408 109.08 ; 
      RECT 41.872 104.706 41.976 109.08 ; 
      RECT 41.44 104.706 41.544 109.08 ; 
      RECT 41.008 104.706 41.112 109.08 ; 
      RECT 40.576 104.706 40.68 109.08 ; 
      RECT 40.144 104.706 40.248 109.08 ; 
      RECT 39.712 104.706 39.816 109.08 ; 
      RECT 39.28 104.706 39.384 109.08 ; 
      RECT 38.848 104.706 38.952 109.08 ; 
      RECT 38.416 104.706 38.52 109.08 ; 
      RECT 37.984 104.706 38.088 109.08 ; 
      RECT 37.552 104.706 37.656 109.08 ; 
      RECT 36.7 104.706 37.008 109.08 ; 
      RECT 29.128 104.706 29.436 109.08 ; 
      RECT 28.48 104.706 28.584 109.08 ; 
      RECT 28.048 104.706 28.152 109.08 ; 
      RECT 27.616 104.706 27.72 109.08 ; 
      RECT 27.184 104.706 27.288 109.08 ; 
      RECT 26.752 104.706 26.856 109.08 ; 
      RECT 26.32 104.706 26.424 109.08 ; 
      RECT 25.888 104.706 25.992 109.08 ; 
      RECT 25.456 104.706 25.56 109.08 ; 
      RECT 25.024 104.706 25.128 109.08 ; 
      RECT 24.592 104.706 24.696 109.08 ; 
      RECT 24.16 104.706 24.264 109.08 ; 
      RECT 23.728 104.706 23.832 109.08 ; 
      RECT 23.296 104.706 23.4 109.08 ; 
      RECT 22.864 104.706 22.968 109.08 ; 
      RECT 22.432 104.706 22.536 109.08 ; 
      RECT 22 104.706 22.104 109.08 ; 
      RECT 21.568 104.706 21.672 109.08 ; 
      RECT 21.136 104.706 21.24 109.08 ; 
      RECT 20.704 104.706 20.808 109.08 ; 
      RECT 20.272 104.706 20.376 109.08 ; 
      RECT 19.84 104.706 19.944 109.08 ; 
      RECT 19.408 104.706 19.512 109.08 ; 
      RECT 18.976 104.706 19.08 109.08 ; 
      RECT 18.544 104.706 18.648 109.08 ; 
      RECT 18.112 104.706 18.216 109.08 ; 
      RECT 17.68 104.706 17.784 109.08 ; 
      RECT 17.248 104.706 17.352 109.08 ; 
      RECT 16.816 104.706 16.92 109.08 ; 
      RECT 16.384 104.706 16.488 109.08 ; 
      RECT 15.952 104.706 16.056 109.08 ; 
      RECT 15.52 104.706 15.624 109.08 ; 
      RECT 15.088 104.706 15.192 109.08 ; 
      RECT 14.656 104.706 14.76 109.08 ; 
      RECT 14.224 104.706 14.328 109.08 ; 
      RECT 13.792 104.706 13.896 109.08 ; 
      RECT 13.36 104.706 13.464 109.08 ; 
      RECT 12.928 104.706 13.032 109.08 ; 
      RECT 12.496 104.706 12.6 109.08 ; 
      RECT 12.064 104.706 12.168 109.08 ; 
      RECT 11.632 104.706 11.736 109.08 ; 
      RECT 11.2 104.706 11.304 109.08 ; 
      RECT 10.768 104.706 10.872 109.08 ; 
      RECT 10.336 104.706 10.44 109.08 ; 
      RECT 9.904 104.706 10.008 109.08 ; 
      RECT 9.472 104.706 9.576 109.08 ; 
      RECT 9.04 104.706 9.144 109.08 ; 
      RECT 8.608 104.706 8.712 109.08 ; 
      RECT 8.176 104.706 8.28 109.08 ; 
      RECT 7.744 104.706 7.848 109.08 ; 
      RECT 7.312 104.706 7.416 109.08 ; 
      RECT 6.88 104.706 6.984 109.08 ; 
      RECT 6.448 104.706 6.552 109.08 ; 
      RECT 6.016 104.706 6.12 109.08 ; 
      RECT 5.584 104.706 5.688 109.08 ; 
      RECT 5.152 104.706 5.256 109.08 ; 
      RECT 4.72 104.706 4.824 109.08 ; 
      RECT 4.288 104.706 4.392 109.08 ; 
      RECT 3.856 104.706 3.96 109.08 ; 
      RECT 3.424 104.706 3.528 109.08 ; 
      RECT 2.992 104.706 3.096 109.08 ; 
      RECT 2.56 104.706 2.664 109.08 ; 
      RECT 2.128 104.706 2.232 109.08 ; 
      RECT 1.696 104.706 1.8 109.08 ; 
      RECT 1.264 104.706 1.368 109.08 ; 
      RECT 0.832 104.706 0.936 109.08 ; 
      RECT 0.02 104.706 0.36 109.08 ; 
      RECT 34.564 109.026 35.076 113.4 ; 
      RECT 34.508 111.688 35.076 112.978 ; 
      RECT 33.916 110.596 34.164 113.4 ; 
      RECT 33.86 111.834 34.164 112.448 ; 
      RECT 33.916 109.026 34.02 113.4 ; 
      RECT 33.916 109.51 34.076 110.468 ; 
      RECT 33.916 109.026 34.164 109.382 ; 
      RECT 32.728 110.828 33.552 113.4 ; 
      RECT 33.448 109.026 33.552 113.4 ; 
      RECT 32.728 111.936 33.608 112.968 ; 
      RECT 32.728 109.026 33.12 113.4 ; 
      RECT 31.06 109.026 31.392 113.4 ; 
      RECT 31.06 109.38 31.448 113.122 ; 
      RECT 65.776 109.026 66.116 113.4 ; 
      RECT 65.2 109.026 65.304 113.4 ; 
      RECT 64.768 109.026 64.872 113.4 ; 
      RECT 64.336 109.026 64.44 113.4 ; 
      RECT 63.904 109.026 64.008 113.4 ; 
      RECT 63.472 109.026 63.576 113.4 ; 
      RECT 63.04 109.026 63.144 113.4 ; 
      RECT 62.608 109.026 62.712 113.4 ; 
      RECT 62.176 109.026 62.28 113.4 ; 
      RECT 61.744 109.026 61.848 113.4 ; 
      RECT 61.312 109.026 61.416 113.4 ; 
      RECT 60.88 109.026 60.984 113.4 ; 
      RECT 60.448 109.026 60.552 113.4 ; 
      RECT 60.016 109.026 60.12 113.4 ; 
      RECT 59.584 109.026 59.688 113.4 ; 
      RECT 59.152 109.026 59.256 113.4 ; 
      RECT 58.72 109.026 58.824 113.4 ; 
      RECT 58.288 109.026 58.392 113.4 ; 
      RECT 57.856 109.026 57.96 113.4 ; 
      RECT 57.424 109.026 57.528 113.4 ; 
      RECT 56.992 109.026 57.096 113.4 ; 
      RECT 56.56 109.026 56.664 113.4 ; 
      RECT 56.128 109.026 56.232 113.4 ; 
      RECT 55.696 109.026 55.8 113.4 ; 
      RECT 55.264 109.026 55.368 113.4 ; 
      RECT 54.832 109.026 54.936 113.4 ; 
      RECT 54.4 109.026 54.504 113.4 ; 
      RECT 53.968 109.026 54.072 113.4 ; 
      RECT 53.536 109.026 53.64 113.4 ; 
      RECT 53.104 109.026 53.208 113.4 ; 
      RECT 52.672 109.026 52.776 113.4 ; 
      RECT 52.24 109.026 52.344 113.4 ; 
      RECT 51.808 109.026 51.912 113.4 ; 
      RECT 51.376 109.026 51.48 113.4 ; 
      RECT 50.944 109.026 51.048 113.4 ; 
      RECT 50.512 109.026 50.616 113.4 ; 
      RECT 50.08 109.026 50.184 113.4 ; 
      RECT 49.648 109.026 49.752 113.4 ; 
      RECT 49.216 109.026 49.32 113.4 ; 
      RECT 48.784 109.026 48.888 113.4 ; 
      RECT 48.352 109.026 48.456 113.4 ; 
      RECT 47.92 109.026 48.024 113.4 ; 
      RECT 47.488 109.026 47.592 113.4 ; 
      RECT 47.056 109.026 47.16 113.4 ; 
      RECT 46.624 109.026 46.728 113.4 ; 
      RECT 46.192 109.026 46.296 113.4 ; 
      RECT 45.76 109.026 45.864 113.4 ; 
      RECT 45.328 109.026 45.432 113.4 ; 
      RECT 44.896 109.026 45 113.4 ; 
      RECT 44.464 109.026 44.568 113.4 ; 
      RECT 44.032 109.026 44.136 113.4 ; 
      RECT 43.6 109.026 43.704 113.4 ; 
      RECT 43.168 109.026 43.272 113.4 ; 
      RECT 42.736 109.026 42.84 113.4 ; 
      RECT 42.304 109.026 42.408 113.4 ; 
      RECT 41.872 109.026 41.976 113.4 ; 
      RECT 41.44 109.026 41.544 113.4 ; 
      RECT 41.008 109.026 41.112 113.4 ; 
      RECT 40.576 109.026 40.68 113.4 ; 
      RECT 40.144 109.026 40.248 113.4 ; 
      RECT 39.712 109.026 39.816 113.4 ; 
      RECT 39.28 109.026 39.384 113.4 ; 
      RECT 38.848 109.026 38.952 113.4 ; 
      RECT 38.416 109.026 38.52 113.4 ; 
      RECT 37.984 109.026 38.088 113.4 ; 
      RECT 37.552 109.026 37.656 113.4 ; 
      RECT 36.7 109.026 37.008 113.4 ; 
      RECT 29.128 109.026 29.436 113.4 ; 
      RECT 28.48 109.026 28.584 113.4 ; 
      RECT 28.048 109.026 28.152 113.4 ; 
      RECT 27.616 109.026 27.72 113.4 ; 
      RECT 27.184 109.026 27.288 113.4 ; 
      RECT 26.752 109.026 26.856 113.4 ; 
      RECT 26.32 109.026 26.424 113.4 ; 
      RECT 25.888 109.026 25.992 113.4 ; 
      RECT 25.456 109.026 25.56 113.4 ; 
      RECT 25.024 109.026 25.128 113.4 ; 
      RECT 24.592 109.026 24.696 113.4 ; 
      RECT 24.16 109.026 24.264 113.4 ; 
      RECT 23.728 109.026 23.832 113.4 ; 
      RECT 23.296 109.026 23.4 113.4 ; 
      RECT 22.864 109.026 22.968 113.4 ; 
      RECT 22.432 109.026 22.536 113.4 ; 
      RECT 22 109.026 22.104 113.4 ; 
      RECT 21.568 109.026 21.672 113.4 ; 
      RECT 21.136 109.026 21.24 113.4 ; 
      RECT 20.704 109.026 20.808 113.4 ; 
      RECT 20.272 109.026 20.376 113.4 ; 
      RECT 19.84 109.026 19.944 113.4 ; 
      RECT 19.408 109.026 19.512 113.4 ; 
      RECT 18.976 109.026 19.08 113.4 ; 
      RECT 18.544 109.026 18.648 113.4 ; 
      RECT 18.112 109.026 18.216 113.4 ; 
      RECT 17.68 109.026 17.784 113.4 ; 
      RECT 17.248 109.026 17.352 113.4 ; 
      RECT 16.816 109.026 16.92 113.4 ; 
      RECT 16.384 109.026 16.488 113.4 ; 
      RECT 15.952 109.026 16.056 113.4 ; 
      RECT 15.52 109.026 15.624 113.4 ; 
      RECT 15.088 109.026 15.192 113.4 ; 
      RECT 14.656 109.026 14.76 113.4 ; 
      RECT 14.224 109.026 14.328 113.4 ; 
      RECT 13.792 109.026 13.896 113.4 ; 
      RECT 13.36 109.026 13.464 113.4 ; 
      RECT 12.928 109.026 13.032 113.4 ; 
      RECT 12.496 109.026 12.6 113.4 ; 
      RECT 12.064 109.026 12.168 113.4 ; 
      RECT 11.632 109.026 11.736 113.4 ; 
      RECT 11.2 109.026 11.304 113.4 ; 
      RECT 10.768 109.026 10.872 113.4 ; 
      RECT 10.336 109.026 10.44 113.4 ; 
      RECT 9.904 109.026 10.008 113.4 ; 
      RECT 9.472 109.026 9.576 113.4 ; 
      RECT 9.04 109.026 9.144 113.4 ; 
      RECT 8.608 109.026 8.712 113.4 ; 
      RECT 8.176 109.026 8.28 113.4 ; 
      RECT 7.744 109.026 7.848 113.4 ; 
      RECT 7.312 109.026 7.416 113.4 ; 
      RECT 6.88 109.026 6.984 113.4 ; 
      RECT 6.448 109.026 6.552 113.4 ; 
      RECT 6.016 109.026 6.12 113.4 ; 
      RECT 5.584 109.026 5.688 113.4 ; 
      RECT 5.152 109.026 5.256 113.4 ; 
      RECT 4.72 109.026 4.824 113.4 ; 
      RECT 4.288 109.026 4.392 113.4 ; 
      RECT 3.856 109.026 3.96 113.4 ; 
      RECT 3.424 109.026 3.528 113.4 ; 
      RECT 2.992 109.026 3.096 113.4 ; 
      RECT 2.56 109.026 2.664 113.4 ; 
      RECT 2.128 109.026 2.232 113.4 ; 
      RECT 1.696 109.026 1.8 113.4 ; 
      RECT 1.264 109.026 1.368 113.4 ; 
      RECT 0.832 109.026 0.936 113.4 ; 
      RECT 0.02 109.026 0.36 113.4 ; 
      RECT 34.564 113.346 35.076 117.72 ; 
      RECT 34.508 116.008 35.076 117.298 ; 
      RECT 33.916 114.916 34.164 117.72 ; 
      RECT 33.86 116.154 34.164 116.768 ; 
      RECT 33.916 113.346 34.02 117.72 ; 
      RECT 33.916 113.83 34.076 114.788 ; 
      RECT 33.916 113.346 34.164 113.702 ; 
      RECT 32.728 115.148 33.552 117.72 ; 
      RECT 33.448 113.346 33.552 117.72 ; 
      RECT 32.728 116.256 33.608 117.288 ; 
      RECT 32.728 113.346 33.12 117.72 ; 
      RECT 31.06 113.346 31.392 117.72 ; 
      RECT 31.06 113.7 31.448 117.442 ; 
      RECT 65.776 113.346 66.116 117.72 ; 
      RECT 65.2 113.346 65.304 117.72 ; 
      RECT 64.768 113.346 64.872 117.72 ; 
      RECT 64.336 113.346 64.44 117.72 ; 
      RECT 63.904 113.346 64.008 117.72 ; 
      RECT 63.472 113.346 63.576 117.72 ; 
      RECT 63.04 113.346 63.144 117.72 ; 
      RECT 62.608 113.346 62.712 117.72 ; 
      RECT 62.176 113.346 62.28 117.72 ; 
      RECT 61.744 113.346 61.848 117.72 ; 
      RECT 61.312 113.346 61.416 117.72 ; 
      RECT 60.88 113.346 60.984 117.72 ; 
      RECT 60.448 113.346 60.552 117.72 ; 
      RECT 60.016 113.346 60.12 117.72 ; 
      RECT 59.584 113.346 59.688 117.72 ; 
      RECT 59.152 113.346 59.256 117.72 ; 
      RECT 58.72 113.346 58.824 117.72 ; 
      RECT 58.288 113.346 58.392 117.72 ; 
      RECT 57.856 113.346 57.96 117.72 ; 
      RECT 57.424 113.346 57.528 117.72 ; 
      RECT 56.992 113.346 57.096 117.72 ; 
      RECT 56.56 113.346 56.664 117.72 ; 
      RECT 56.128 113.346 56.232 117.72 ; 
      RECT 55.696 113.346 55.8 117.72 ; 
      RECT 55.264 113.346 55.368 117.72 ; 
      RECT 54.832 113.346 54.936 117.72 ; 
      RECT 54.4 113.346 54.504 117.72 ; 
      RECT 53.968 113.346 54.072 117.72 ; 
      RECT 53.536 113.346 53.64 117.72 ; 
      RECT 53.104 113.346 53.208 117.72 ; 
      RECT 52.672 113.346 52.776 117.72 ; 
      RECT 52.24 113.346 52.344 117.72 ; 
      RECT 51.808 113.346 51.912 117.72 ; 
      RECT 51.376 113.346 51.48 117.72 ; 
      RECT 50.944 113.346 51.048 117.72 ; 
      RECT 50.512 113.346 50.616 117.72 ; 
      RECT 50.08 113.346 50.184 117.72 ; 
      RECT 49.648 113.346 49.752 117.72 ; 
      RECT 49.216 113.346 49.32 117.72 ; 
      RECT 48.784 113.346 48.888 117.72 ; 
      RECT 48.352 113.346 48.456 117.72 ; 
      RECT 47.92 113.346 48.024 117.72 ; 
      RECT 47.488 113.346 47.592 117.72 ; 
      RECT 47.056 113.346 47.16 117.72 ; 
      RECT 46.624 113.346 46.728 117.72 ; 
      RECT 46.192 113.346 46.296 117.72 ; 
      RECT 45.76 113.346 45.864 117.72 ; 
      RECT 45.328 113.346 45.432 117.72 ; 
      RECT 44.896 113.346 45 117.72 ; 
      RECT 44.464 113.346 44.568 117.72 ; 
      RECT 44.032 113.346 44.136 117.72 ; 
      RECT 43.6 113.346 43.704 117.72 ; 
      RECT 43.168 113.346 43.272 117.72 ; 
      RECT 42.736 113.346 42.84 117.72 ; 
      RECT 42.304 113.346 42.408 117.72 ; 
      RECT 41.872 113.346 41.976 117.72 ; 
      RECT 41.44 113.346 41.544 117.72 ; 
      RECT 41.008 113.346 41.112 117.72 ; 
      RECT 40.576 113.346 40.68 117.72 ; 
      RECT 40.144 113.346 40.248 117.72 ; 
      RECT 39.712 113.346 39.816 117.72 ; 
      RECT 39.28 113.346 39.384 117.72 ; 
      RECT 38.848 113.346 38.952 117.72 ; 
      RECT 38.416 113.346 38.52 117.72 ; 
      RECT 37.984 113.346 38.088 117.72 ; 
      RECT 37.552 113.346 37.656 117.72 ; 
      RECT 36.7 113.346 37.008 117.72 ; 
      RECT 29.128 113.346 29.436 117.72 ; 
      RECT 28.48 113.346 28.584 117.72 ; 
      RECT 28.048 113.346 28.152 117.72 ; 
      RECT 27.616 113.346 27.72 117.72 ; 
      RECT 27.184 113.346 27.288 117.72 ; 
      RECT 26.752 113.346 26.856 117.72 ; 
      RECT 26.32 113.346 26.424 117.72 ; 
      RECT 25.888 113.346 25.992 117.72 ; 
      RECT 25.456 113.346 25.56 117.72 ; 
      RECT 25.024 113.346 25.128 117.72 ; 
      RECT 24.592 113.346 24.696 117.72 ; 
      RECT 24.16 113.346 24.264 117.72 ; 
      RECT 23.728 113.346 23.832 117.72 ; 
      RECT 23.296 113.346 23.4 117.72 ; 
      RECT 22.864 113.346 22.968 117.72 ; 
      RECT 22.432 113.346 22.536 117.72 ; 
      RECT 22 113.346 22.104 117.72 ; 
      RECT 21.568 113.346 21.672 117.72 ; 
      RECT 21.136 113.346 21.24 117.72 ; 
      RECT 20.704 113.346 20.808 117.72 ; 
      RECT 20.272 113.346 20.376 117.72 ; 
      RECT 19.84 113.346 19.944 117.72 ; 
      RECT 19.408 113.346 19.512 117.72 ; 
      RECT 18.976 113.346 19.08 117.72 ; 
      RECT 18.544 113.346 18.648 117.72 ; 
      RECT 18.112 113.346 18.216 117.72 ; 
      RECT 17.68 113.346 17.784 117.72 ; 
      RECT 17.248 113.346 17.352 117.72 ; 
      RECT 16.816 113.346 16.92 117.72 ; 
      RECT 16.384 113.346 16.488 117.72 ; 
      RECT 15.952 113.346 16.056 117.72 ; 
      RECT 15.52 113.346 15.624 117.72 ; 
      RECT 15.088 113.346 15.192 117.72 ; 
      RECT 14.656 113.346 14.76 117.72 ; 
      RECT 14.224 113.346 14.328 117.72 ; 
      RECT 13.792 113.346 13.896 117.72 ; 
      RECT 13.36 113.346 13.464 117.72 ; 
      RECT 12.928 113.346 13.032 117.72 ; 
      RECT 12.496 113.346 12.6 117.72 ; 
      RECT 12.064 113.346 12.168 117.72 ; 
      RECT 11.632 113.346 11.736 117.72 ; 
      RECT 11.2 113.346 11.304 117.72 ; 
      RECT 10.768 113.346 10.872 117.72 ; 
      RECT 10.336 113.346 10.44 117.72 ; 
      RECT 9.904 113.346 10.008 117.72 ; 
      RECT 9.472 113.346 9.576 117.72 ; 
      RECT 9.04 113.346 9.144 117.72 ; 
      RECT 8.608 113.346 8.712 117.72 ; 
      RECT 8.176 113.346 8.28 117.72 ; 
      RECT 7.744 113.346 7.848 117.72 ; 
      RECT 7.312 113.346 7.416 117.72 ; 
      RECT 6.88 113.346 6.984 117.72 ; 
      RECT 6.448 113.346 6.552 117.72 ; 
      RECT 6.016 113.346 6.12 117.72 ; 
      RECT 5.584 113.346 5.688 117.72 ; 
      RECT 5.152 113.346 5.256 117.72 ; 
      RECT 4.72 113.346 4.824 117.72 ; 
      RECT 4.288 113.346 4.392 117.72 ; 
      RECT 3.856 113.346 3.96 117.72 ; 
      RECT 3.424 113.346 3.528 117.72 ; 
      RECT 2.992 113.346 3.096 117.72 ; 
      RECT 2.56 113.346 2.664 117.72 ; 
      RECT 2.128 113.346 2.232 117.72 ; 
      RECT 1.696 113.346 1.8 117.72 ; 
      RECT 1.264 113.346 1.368 117.72 ; 
      RECT 0.832 113.346 0.936 117.72 ; 
      RECT 0.02 113.346 0.36 117.72 ; 
      RECT 34.564 117.666 35.076 122.04 ; 
      RECT 34.508 120.328 35.076 121.618 ; 
      RECT 33.916 119.236 34.164 122.04 ; 
      RECT 33.86 120.474 34.164 121.088 ; 
      RECT 33.916 117.666 34.02 122.04 ; 
      RECT 33.916 118.15 34.076 119.108 ; 
      RECT 33.916 117.666 34.164 118.022 ; 
      RECT 32.728 119.468 33.552 122.04 ; 
      RECT 33.448 117.666 33.552 122.04 ; 
      RECT 32.728 120.576 33.608 121.608 ; 
      RECT 32.728 117.666 33.12 122.04 ; 
      RECT 31.06 117.666 31.392 122.04 ; 
      RECT 31.06 118.02 31.448 121.762 ; 
      RECT 65.776 117.666 66.116 122.04 ; 
      RECT 65.2 117.666 65.304 122.04 ; 
      RECT 64.768 117.666 64.872 122.04 ; 
      RECT 64.336 117.666 64.44 122.04 ; 
      RECT 63.904 117.666 64.008 122.04 ; 
      RECT 63.472 117.666 63.576 122.04 ; 
      RECT 63.04 117.666 63.144 122.04 ; 
      RECT 62.608 117.666 62.712 122.04 ; 
      RECT 62.176 117.666 62.28 122.04 ; 
      RECT 61.744 117.666 61.848 122.04 ; 
      RECT 61.312 117.666 61.416 122.04 ; 
      RECT 60.88 117.666 60.984 122.04 ; 
      RECT 60.448 117.666 60.552 122.04 ; 
      RECT 60.016 117.666 60.12 122.04 ; 
      RECT 59.584 117.666 59.688 122.04 ; 
      RECT 59.152 117.666 59.256 122.04 ; 
      RECT 58.72 117.666 58.824 122.04 ; 
      RECT 58.288 117.666 58.392 122.04 ; 
      RECT 57.856 117.666 57.96 122.04 ; 
      RECT 57.424 117.666 57.528 122.04 ; 
      RECT 56.992 117.666 57.096 122.04 ; 
      RECT 56.56 117.666 56.664 122.04 ; 
      RECT 56.128 117.666 56.232 122.04 ; 
      RECT 55.696 117.666 55.8 122.04 ; 
      RECT 55.264 117.666 55.368 122.04 ; 
      RECT 54.832 117.666 54.936 122.04 ; 
      RECT 54.4 117.666 54.504 122.04 ; 
      RECT 53.968 117.666 54.072 122.04 ; 
      RECT 53.536 117.666 53.64 122.04 ; 
      RECT 53.104 117.666 53.208 122.04 ; 
      RECT 52.672 117.666 52.776 122.04 ; 
      RECT 52.24 117.666 52.344 122.04 ; 
      RECT 51.808 117.666 51.912 122.04 ; 
      RECT 51.376 117.666 51.48 122.04 ; 
      RECT 50.944 117.666 51.048 122.04 ; 
      RECT 50.512 117.666 50.616 122.04 ; 
      RECT 50.08 117.666 50.184 122.04 ; 
      RECT 49.648 117.666 49.752 122.04 ; 
      RECT 49.216 117.666 49.32 122.04 ; 
      RECT 48.784 117.666 48.888 122.04 ; 
      RECT 48.352 117.666 48.456 122.04 ; 
      RECT 47.92 117.666 48.024 122.04 ; 
      RECT 47.488 117.666 47.592 122.04 ; 
      RECT 47.056 117.666 47.16 122.04 ; 
      RECT 46.624 117.666 46.728 122.04 ; 
      RECT 46.192 117.666 46.296 122.04 ; 
      RECT 45.76 117.666 45.864 122.04 ; 
      RECT 45.328 117.666 45.432 122.04 ; 
      RECT 44.896 117.666 45 122.04 ; 
      RECT 44.464 117.666 44.568 122.04 ; 
      RECT 44.032 117.666 44.136 122.04 ; 
      RECT 43.6 117.666 43.704 122.04 ; 
      RECT 43.168 117.666 43.272 122.04 ; 
      RECT 42.736 117.666 42.84 122.04 ; 
      RECT 42.304 117.666 42.408 122.04 ; 
      RECT 41.872 117.666 41.976 122.04 ; 
      RECT 41.44 117.666 41.544 122.04 ; 
      RECT 41.008 117.666 41.112 122.04 ; 
      RECT 40.576 117.666 40.68 122.04 ; 
      RECT 40.144 117.666 40.248 122.04 ; 
      RECT 39.712 117.666 39.816 122.04 ; 
      RECT 39.28 117.666 39.384 122.04 ; 
      RECT 38.848 117.666 38.952 122.04 ; 
      RECT 38.416 117.666 38.52 122.04 ; 
      RECT 37.984 117.666 38.088 122.04 ; 
      RECT 37.552 117.666 37.656 122.04 ; 
      RECT 36.7 117.666 37.008 122.04 ; 
      RECT 29.128 117.666 29.436 122.04 ; 
      RECT 28.48 117.666 28.584 122.04 ; 
      RECT 28.048 117.666 28.152 122.04 ; 
      RECT 27.616 117.666 27.72 122.04 ; 
      RECT 27.184 117.666 27.288 122.04 ; 
      RECT 26.752 117.666 26.856 122.04 ; 
      RECT 26.32 117.666 26.424 122.04 ; 
      RECT 25.888 117.666 25.992 122.04 ; 
      RECT 25.456 117.666 25.56 122.04 ; 
      RECT 25.024 117.666 25.128 122.04 ; 
      RECT 24.592 117.666 24.696 122.04 ; 
      RECT 24.16 117.666 24.264 122.04 ; 
      RECT 23.728 117.666 23.832 122.04 ; 
      RECT 23.296 117.666 23.4 122.04 ; 
      RECT 22.864 117.666 22.968 122.04 ; 
      RECT 22.432 117.666 22.536 122.04 ; 
      RECT 22 117.666 22.104 122.04 ; 
      RECT 21.568 117.666 21.672 122.04 ; 
      RECT 21.136 117.666 21.24 122.04 ; 
      RECT 20.704 117.666 20.808 122.04 ; 
      RECT 20.272 117.666 20.376 122.04 ; 
      RECT 19.84 117.666 19.944 122.04 ; 
      RECT 19.408 117.666 19.512 122.04 ; 
      RECT 18.976 117.666 19.08 122.04 ; 
      RECT 18.544 117.666 18.648 122.04 ; 
      RECT 18.112 117.666 18.216 122.04 ; 
      RECT 17.68 117.666 17.784 122.04 ; 
      RECT 17.248 117.666 17.352 122.04 ; 
      RECT 16.816 117.666 16.92 122.04 ; 
      RECT 16.384 117.666 16.488 122.04 ; 
      RECT 15.952 117.666 16.056 122.04 ; 
      RECT 15.52 117.666 15.624 122.04 ; 
      RECT 15.088 117.666 15.192 122.04 ; 
      RECT 14.656 117.666 14.76 122.04 ; 
      RECT 14.224 117.666 14.328 122.04 ; 
      RECT 13.792 117.666 13.896 122.04 ; 
      RECT 13.36 117.666 13.464 122.04 ; 
      RECT 12.928 117.666 13.032 122.04 ; 
      RECT 12.496 117.666 12.6 122.04 ; 
      RECT 12.064 117.666 12.168 122.04 ; 
      RECT 11.632 117.666 11.736 122.04 ; 
      RECT 11.2 117.666 11.304 122.04 ; 
      RECT 10.768 117.666 10.872 122.04 ; 
      RECT 10.336 117.666 10.44 122.04 ; 
      RECT 9.904 117.666 10.008 122.04 ; 
      RECT 9.472 117.666 9.576 122.04 ; 
      RECT 9.04 117.666 9.144 122.04 ; 
      RECT 8.608 117.666 8.712 122.04 ; 
      RECT 8.176 117.666 8.28 122.04 ; 
      RECT 7.744 117.666 7.848 122.04 ; 
      RECT 7.312 117.666 7.416 122.04 ; 
      RECT 6.88 117.666 6.984 122.04 ; 
      RECT 6.448 117.666 6.552 122.04 ; 
      RECT 6.016 117.666 6.12 122.04 ; 
      RECT 5.584 117.666 5.688 122.04 ; 
      RECT 5.152 117.666 5.256 122.04 ; 
      RECT 4.72 117.666 4.824 122.04 ; 
      RECT 4.288 117.666 4.392 122.04 ; 
      RECT 3.856 117.666 3.96 122.04 ; 
      RECT 3.424 117.666 3.528 122.04 ; 
      RECT 2.992 117.666 3.096 122.04 ; 
      RECT 2.56 117.666 2.664 122.04 ; 
      RECT 2.128 117.666 2.232 122.04 ; 
      RECT 1.696 117.666 1.8 122.04 ; 
      RECT 1.264 117.666 1.368 122.04 ; 
      RECT 0.832 117.666 0.936 122.04 ; 
      RECT 0.02 117.666 0.36 122.04 ; 
      RECT 34.564 121.986 35.076 126.36 ; 
      RECT 34.508 124.648 35.076 125.938 ; 
      RECT 33.916 123.556 34.164 126.36 ; 
      RECT 33.86 124.794 34.164 125.408 ; 
      RECT 33.916 121.986 34.02 126.36 ; 
      RECT 33.916 122.47 34.076 123.428 ; 
      RECT 33.916 121.986 34.164 122.342 ; 
      RECT 32.728 123.788 33.552 126.36 ; 
      RECT 33.448 121.986 33.552 126.36 ; 
      RECT 32.728 124.896 33.608 125.928 ; 
      RECT 32.728 121.986 33.12 126.36 ; 
      RECT 31.06 121.986 31.392 126.36 ; 
      RECT 31.06 122.34 31.448 126.082 ; 
      RECT 65.776 121.986 66.116 126.36 ; 
      RECT 65.2 121.986 65.304 126.36 ; 
      RECT 64.768 121.986 64.872 126.36 ; 
      RECT 64.336 121.986 64.44 126.36 ; 
      RECT 63.904 121.986 64.008 126.36 ; 
      RECT 63.472 121.986 63.576 126.36 ; 
      RECT 63.04 121.986 63.144 126.36 ; 
      RECT 62.608 121.986 62.712 126.36 ; 
      RECT 62.176 121.986 62.28 126.36 ; 
      RECT 61.744 121.986 61.848 126.36 ; 
      RECT 61.312 121.986 61.416 126.36 ; 
      RECT 60.88 121.986 60.984 126.36 ; 
      RECT 60.448 121.986 60.552 126.36 ; 
      RECT 60.016 121.986 60.12 126.36 ; 
      RECT 59.584 121.986 59.688 126.36 ; 
      RECT 59.152 121.986 59.256 126.36 ; 
      RECT 58.72 121.986 58.824 126.36 ; 
      RECT 58.288 121.986 58.392 126.36 ; 
      RECT 57.856 121.986 57.96 126.36 ; 
      RECT 57.424 121.986 57.528 126.36 ; 
      RECT 56.992 121.986 57.096 126.36 ; 
      RECT 56.56 121.986 56.664 126.36 ; 
      RECT 56.128 121.986 56.232 126.36 ; 
      RECT 55.696 121.986 55.8 126.36 ; 
      RECT 55.264 121.986 55.368 126.36 ; 
      RECT 54.832 121.986 54.936 126.36 ; 
      RECT 54.4 121.986 54.504 126.36 ; 
      RECT 53.968 121.986 54.072 126.36 ; 
      RECT 53.536 121.986 53.64 126.36 ; 
      RECT 53.104 121.986 53.208 126.36 ; 
      RECT 52.672 121.986 52.776 126.36 ; 
      RECT 52.24 121.986 52.344 126.36 ; 
      RECT 51.808 121.986 51.912 126.36 ; 
      RECT 51.376 121.986 51.48 126.36 ; 
      RECT 50.944 121.986 51.048 126.36 ; 
      RECT 50.512 121.986 50.616 126.36 ; 
      RECT 50.08 121.986 50.184 126.36 ; 
      RECT 49.648 121.986 49.752 126.36 ; 
      RECT 49.216 121.986 49.32 126.36 ; 
      RECT 48.784 121.986 48.888 126.36 ; 
      RECT 48.352 121.986 48.456 126.36 ; 
      RECT 47.92 121.986 48.024 126.36 ; 
      RECT 47.488 121.986 47.592 126.36 ; 
      RECT 47.056 121.986 47.16 126.36 ; 
      RECT 46.624 121.986 46.728 126.36 ; 
      RECT 46.192 121.986 46.296 126.36 ; 
      RECT 45.76 121.986 45.864 126.36 ; 
      RECT 45.328 121.986 45.432 126.36 ; 
      RECT 44.896 121.986 45 126.36 ; 
      RECT 44.464 121.986 44.568 126.36 ; 
      RECT 44.032 121.986 44.136 126.36 ; 
      RECT 43.6 121.986 43.704 126.36 ; 
      RECT 43.168 121.986 43.272 126.36 ; 
      RECT 42.736 121.986 42.84 126.36 ; 
      RECT 42.304 121.986 42.408 126.36 ; 
      RECT 41.872 121.986 41.976 126.36 ; 
      RECT 41.44 121.986 41.544 126.36 ; 
      RECT 41.008 121.986 41.112 126.36 ; 
      RECT 40.576 121.986 40.68 126.36 ; 
      RECT 40.144 121.986 40.248 126.36 ; 
      RECT 39.712 121.986 39.816 126.36 ; 
      RECT 39.28 121.986 39.384 126.36 ; 
      RECT 38.848 121.986 38.952 126.36 ; 
      RECT 38.416 121.986 38.52 126.36 ; 
      RECT 37.984 121.986 38.088 126.36 ; 
      RECT 37.552 121.986 37.656 126.36 ; 
      RECT 36.7 121.986 37.008 126.36 ; 
      RECT 29.128 121.986 29.436 126.36 ; 
      RECT 28.48 121.986 28.584 126.36 ; 
      RECT 28.048 121.986 28.152 126.36 ; 
      RECT 27.616 121.986 27.72 126.36 ; 
      RECT 27.184 121.986 27.288 126.36 ; 
      RECT 26.752 121.986 26.856 126.36 ; 
      RECT 26.32 121.986 26.424 126.36 ; 
      RECT 25.888 121.986 25.992 126.36 ; 
      RECT 25.456 121.986 25.56 126.36 ; 
      RECT 25.024 121.986 25.128 126.36 ; 
      RECT 24.592 121.986 24.696 126.36 ; 
      RECT 24.16 121.986 24.264 126.36 ; 
      RECT 23.728 121.986 23.832 126.36 ; 
      RECT 23.296 121.986 23.4 126.36 ; 
      RECT 22.864 121.986 22.968 126.36 ; 
      RECT 22.432 121.986 22.536 126.36 ; 
      RECT 22 121.986 22.104 126.36 ; 
      RECT 21.568 121.986 21.672 126.36 ; 
      RECT 21.136 121.986 21.24 126.36 ; 
      RECT 20.704 121.986 20.808 126.36 ; 
      RECT 20.272 121.986 20.376 126.36 ; 
      RECT 19.84 121.986 19.944 126.36 ; 
      RECT 19.408 121.986 19.512 126.36 ; 
      RECT 18.976 121.986 19.08 126.36 ; 
      RECT 18.544 121.986 18.648 126.36 ; 
      RECT 18.112 121.986 18.216 126.36 ; 
      RECT 17.68 121.986 17.784 126.36 ; 
      RECT 17.248 121.986 17.352 126.36 ; 
      RECT 16.816 121.986 16.92 126.36 ; 
      RECT 16.384 121.986 16.488 126.36 ; 
      RECT 15.952 121.986 16.056 126.36 ; 
      RECT 15.52 121.986 15.624 126.36 ; 
      RECT 15.088 121.986 15.192 126.36 ; 
      RECT 14.656 121.986 14.76 126.36 ; 
      RECT 14.224 121.986 14.328 126.36 ; 
      RECT 13.792 121.986 13.896 126.36 ; 
      RECT 13.36 121.986 13.464 126.36 ; 
      RECT 12.928 121.986 13.032 126.36 ; 
      RECT 12.496 121.986 12.6 126.36 ; 
      RECT 12.064 121.986 12.168 126.36 ; 
      RECT 11.632 121.986 11.736 126.36 ; 
      RECT 11.2 121.986 11.304 126.36 ; 
      RECT 10.768 121.986 10.872 126.36 ; 
      RECT 10.336 121.986 10.44 126.36 ; 
      RECT 9.904 121.986 10.008 126.36 ; 
      RECT 9.472 121.986 9.576 126.36 ; 
      RECT 9.04 121.986 9.144 126.36 ; 
      RECT 8.608 121.986 8.712 126.36 ; 
      RECT 8.176 121.986 8.28 126.36 ; 
      RECT 7.744 121.986 7.848 126.36 ; 
      RECT 7.312 121.986 7.416 126.36 ; 
      RECT 6.88 121.986 6.984 126.36 ; 
      RECT 6.448 121.986 6.552 126.36 ; 
      RECT 6.016 121.986 6.12 126.36 ; 
      RECT 5.584 121.986 5.688 126.36 ; 
      RECT 5.152 121.986 5.256 126.36 ; 
      RECT 4.72 121.986 4.824 126.36 ; 
      RECT 4.288 121.986 4.392 126.36 ; 
      RECT 3.856 121.986 3.96 126.36 ; 
      RECT 3.424 121.986 3.528 126.36 ; 
      RECT 2.992 121.986 3.096 126.36 ; 
      RECT 2.56 121.986 2.664 126.36 ; 
      RECT 2.128 121.986 2.232 126.36 ; 
      RECT 1.696 121.986 1.8 126.36 ; 
      RECT 1.264 121.986 1.368 126.36 ; 
      RECT 0.832 121.986 0.936 126.36 ; 
      RECT 0.02 121.986 0.36 126.36 ; 
      RECT 34.564 126.306 35.076 130.68 ; 
      RECT 34.508 128.968 35.076 130.258 ; 
      RECT 33.916 127.876 34.164 130.68 ; 
      RECT 33.86 129.114 34.164 129.728 ; 
      RECT 33.916 126.306 34.02 130.68 ; 
      RECT 33.916 126.79 34.076 127.748 ; 
      RECT 33.916 126.306 34.164 126.662 ; 
      RECT 32.728 128.108 33.552 130.68 ; 
      RECT 33.448 126.306 33.552 130.68 ; 
      RECT 32.728 129.216 33.608 130.248 ; 
      RECT 32.728 126.306 33.12 130.68 ; 
      RECT 31.06 126.306 31.392 130.68 ; 
      RECT 31.06 126.66 31.448 130.402 ; 
      RECT 65.776 126.306 66.116 130.68 ; 
      RECT 65.2 126.306 65.304 130.68 ; 
      RECT 64.768 126.306 64.872 130.68 ; 
      RECT 64.336 126.306 64.44 130.68 ; 
      RECT 63.904 126.306 64.008 130.68 ; 
      RECT 63.472 126.306 63.576 130.68 ; 
      RECT 63.04 126.306 63.144 130.68 ; 
      RECT 62.608 126.306 62.712 130.68 ; 
      RECT 62.176 126.306 62.28 130.68 ; 
      RECT 61.744 126.306 61.848 130.68 ; 
      RECT 61.312 126.306 61.416 130.68 ; 
      RECT 60.88 126.306 60.984 130.68 ; 
      RECT 60.448 126.306 60.552 130.68 ; 
      RECT 60.016 126.306 60.12 130.68 ; 
      RECT 59.584 126.306 59.688 130.68 ; 
      RECT 59.152 126.306 59.256 130.68 ; 
      RECT 58.72 126.306 58.824 130.68 ; 
      RECT 58.288 126.306 58.392 130.68 ; 
      RECT 57.856 126.306 57.96 130.68 ; 
      RECT 57.424 126.306 57.528 130.68 ; 
      RECT 56.992 126.306 57.096 130.68 ; 
      RECT 56.56 126.306 56.664 130.68 ; 
      RECT 56.128 126.306 56.232 130.68 ; 
      RECT 55.696 126.306 55.8 130.68 ; 
      RECT 55.264 126.306 55.368 130.68 ; 
      RECT 54.832 126.306 54.936 130.68 ; 
      RECT 54.4 126.306 54.504 130.68 ; 
      RECT 53.968 126.306 54.072 130.68 ; 
      RECT 53.536 126.306 53.64 130.68 ; 
      RECT 53.104 126.306 53.208 130.68 ; 
      RECT 52.672 126.306 52.776 130.68 ; 
      RECT 52.24 126.306 52.344 130.68 ; 
      RECT 51.808 126.306 51.912 130.68 ; 
      RECT 51.376 126.306 51.48 130.68 ; 
      RECT 50.944 126.306 51.048 130.68 ; 
      RECT 50.512 126.306 50.616 130.68 ; 
      RECT 50.08 126.306 50.184 130.68 ; 
      RECT 49.648 126.306 49.752 130.68 ; 
      RECT 49.216 126.306 49.32 130.68 ; 
      RECT 48.784 126.306 48.888 130.68 ; 
      RECT 48.352 126.306 48.456 130.68 ; 
      RECT 47.92 126.306 48.024 130.68 ; 
      RECT 47.488 126.306 47.592 130.68 ; 
      RECT 47.056 126.306 47.16 130.68 ; 
      RECT 46.624 126.306 46.728 130.68 ; 
      RECT 46.192 126.306 46.296 130.68 ; 
      RECT 45.76 126.306 45.864 130.68 ; 
      RECT 45.328 126.306 45.432 130.68 ; 
      RECT 44.896 126.306 45 130.68 ; 
      RECT 44.464 126.306 44.568 130.68 ; 
      RECT 44.032 126.306 44.136 130.68 ; 
      RECT 43.6 126.306 43.704 130.68 ; 
      RECT 43.168 126.306 43.272 130.68 ; 
      RECT 42.736 126.306 42.84 130.68 ; 
      RECT 42.304 126.306 42.408 130.68 ; 
      RECT 41.872 126.306 41.976 130.68 ; 
      RECT 41.44 126.306 41.544 130.68 ; 
      RECT 41.008 126.306 41.112 130.68 ; 
      RECT 40.576 126.306 40.68 130.68 ; 
      RECT 40.144 126.306 40.248 130.68 ; 
      RECT 39.712 126.306 39.816 130.68 ; 
      RECT 39.28 126.306 39.384 130.68 ; 
      RECT 38.848 126.306 38.952 130.68 ; 
      RECT 38.416 126.306 38.52 130.68 ; 
      RECT 37.984 126.306 38.088 130.68 ; 
      RECT 37.552 126.306 37.656 130.68 ; 
      RECT 36.7 126.306 37.008 130.68 ; 
      RECT 29.128 126.306 29.436 130.68 ; 
      RECT 28.48 126.306 28.584 130.68 ; 
      RECT 28.048 126.306 28.152 130.68 ; 
      RECT 27.616 126.306 27.72 130.68 ; 
      RECT 27.184 126.306 27.288 130.68 ; 
      RECT 26.752 126.306 26.856 130.68 ; 
      RECT 26.32 126.306 26.424 130.68 ; 
      RECT 25.888 126.306 25.992 130.68 ; 
      RECT 25.456 126.306 25.56 130.68 ; 
      RECT 25.024 126.306 25.128 130.68 ; 
      RECT 24.592 126.306 24.696 130.68 ; 
      RECT 24.16 126.306 24.264 130.68 ; 
      RECT 23.728 126.306 23.832 130.68 ; 
      RECT 23.296 126.306 23.4 130.68 ; 
      RECT 22.864 126.306 22.968 130.68 ; 
      RECT 22.432 126.306 22.536 130.68 ; 
      RECT 22 126.306 22.104 130.68 ; 
      RECT 21.568 126.306 21.672 130.68 ; 
      RECT 21.136 126.306 21.24 130.68 ; 
      RECT 20.704 126.306 20.808 130.68 ; 
      RECT 20.272 126.306 20.376 130.68 ; 
      RECT 19.84 126.306 19.944 130.68 ; 
      RECT 19.408 126.306 19.512 130.68 ; 
      RECT 18.976 126.306 19.08 130.68 ; 
      RECT 18.544 126.306 18.648 130.68 ; 
      RECT 18.112 126.306 18.216 130.68 ; 
      RECT 17.68 126.306 17.784 130.68 ; 
      RECT 17.248 126.306 17.352 130.68 ; 
      RECT 16.816 126.306 16.92 130.68 ; 
      RECT 16.384 126.306 16.488 130.68 ; 
      RECT 15.952 126.306 16.056 130.68 ; 
      RECT 15.52 126.306 15.624 130.68 ; 
      RECT 15.088 126.306 15.192 130.68 ; 
      RECT 14.656 126.306 14.76 130.68 ; 
      RECT 14.224 126.306 14.328 130.68 ; 
      RECT 13.792 126.306 13.896 130.68 ; 
      RECT 13.36 126.306 13.464 130.68 ; 
      RECT 12.928 126.306 13.032 130.68 ; 
      RECT 12.496 126.306 12.6 130.68 ; 
      RECT 12.064 126.306 12.168 130.68 ; 
      RECT 11.632 126.306 11.736 130.68 ; 
      RECT 11.2 126.306 11.304 130.68 ; 
      RECT 10.768 126.306 10.872 130.68 ; 
      RECT 10.336 126.306 10.44 130.68 ; 
      RECT 9.904 126.306 10.008 130.68 ; 
      RECT 9.472 126.306 9.576 130.68 ; 
      RECT 9.04 126.306 9.144 130.68 ; 
      RECT 8.608 126.306 8.712 130.68 ; 
      RECT 8.176 126.306 8.28 130.68 ; 
      RECT 7.744 126.306 7.848 130.68 ; 
      RECT 7.312 126.306 7.416 130.68 ; 
      RECT 6.88 126.306 6.984 130.68 ; 
      RECT 6.448 126.306 6.552 130.68 ; 
      RECT 6.016 126.306 6.12 130.68 ; 
      RECT 5.584 126.306 5.688 130.68 ; 
      RECT 5.152 126.306 5.256 130.68 ; 
      RECT 4.72 126.306 4.824 130.68 ; 
      RECT 4.288 126.306 4.392 130.68 ; 
      RECT 3.856 126.306 3.96 130.68 ; 
      RECT 3.424 126.306 3.528 130.68 ; 
      RECT 2.992 126.306 3.096 130.68 ; 
      RECT 2.56 126.306 2.664 130.68 ; 
      RECT 2.128 126.306 2.232 130.68 ; 
      RECT 1.696 126.306 1.8 130.68 ; 
      RECT 1.264 126.306 1.368 130.68 ; 
      RECT 0.832 126.306 0.936 130.68 ; 
      RECT 0.02 126.306 0.36 130.68 ; 
      RECT 34.564 130.626 35.076 135 ; 
      RECT 34.508 133.288 35.076 134.578 ; 
      RECT 33.916 132.196 34.164 135 ; 
      RECT 33.86 133.434 34.164 134.048 ; 
      RECT 33.916 130.626 34.02 135 ; 
      RECT 33.916 131.11 34.076 132.068 ; 
      RECT 33.916 130.626 34.164 130.982 ; 
      RECT 32.728 132.428 33.552 135 ; 
      RECT 33.448 130.626 33.552 135 ; 
      RECT 32.728 133.536 33.608 134.568 ; 
      RECT 32.728 130.626 33.12 135 ; 
      RECT 31.06 130.626 31.392 135 ; 
      RECT 31.06 130.98 31.448 134.722 ; 
      RECT 65.776 130.626 66.116 135 ; 
      RECT 65.2 130.626 65.304 135 ; 
      RECT 64.768 130.626 64.872 135 ; 
      RECT 64.336 130.626 64.44 135 ; 
      RECT 63.904 130.626 64.008 135 ; 
      RECT 63.472 130.626 63.576 135 ; 
      RECT 63.04 130.626 63.144 135 ; 
      RECT 62.608 130.626 62.712 135 ; 
      RECT 62.176 130.626 62.28 135 ; 
      RECT 61.744 130.626 61.848 135 ; 
      RECT 61.312 130.626 61.416 135 ; 
      RECT 60.88 130.626 60.984 135 ; 
      RECT 60.448 130.626 60.552 135 ; 
      RECT 60.016 130.626 60.12 135 ; 
      RECT 59.584 130.626 59.688 135 ; 
      RECT 59.152 130.626 59.256 135 ; 
      RECT 58.72 130.626 58.824 135 ; 
      RECT 58.288 130.626 58.392 135 ; 
      RECT 57.856 130.626 57.96 135 ; 
      RECT 57.424 130.626 57.528 135 ; 
      RECT 56.992 130.626 57.096 135 ; 
      RECT 56.56 130.626 56.664 135 ; 
      RECT 56.128 130.626 56.232 135 ; 
      RECT 55.696 130.626 55.8 135 ; 
      RECT 55.264 130.626 55.368 135 ; 
      RECT 54.832 130.626 54.936 135 ; 
      RECT 54.4 130.626 54.504 135 ; 
      RECT 53.968 130.626 54.072 135 ; 
      RECT 53.536 130.626 53.64 135 ; 
      RECT 53.104 130.626 53.208 135 ; 
      RECT 52.672 130.626 52.776 135 ; 
      RECT 52.24 130.626 52.344 135 ; 
      RECT 51.808 130.626 51.912 135 ; 
      RECT 51.376 130.626 51.48 135 ; 
      RECT 50.944 130.626 51.048 135 ; 
      RECT 50.512 130.626 50.616 135 ; 
      RECT 50.08 130.626 50.184 135 ; 
      RECT 49.648 130.626 49.752 135 ; 
      RECT 49.216 130.626 49.32 135 ; 
      RECT 48.784 130.626 48.888 135 ; 
      RECT 48.352 130.626 48.456 135 ; 
      RECT 47.92 130.626 48.024 135 ; 
      RECT 47.488 130.626 47.592 135 ; 
      RECT 47.056 130.626 47.16 135 ; 
      RECT 46.624 130.626 46.728 135 ; 
      RECT 46.192 130.626 46.296 135 ; 
      RECT 45.76 130.626 45.864 135 ; 
      RECT 45.328 130.626 45.432 135 ; 
      RECT 44.896 130.626 45 135 ; 
      RECT 44.464 130.626 44.568 135 ; 
      RECT 44.032 130.626 44.136 135 ; 
      RECT 43.6 130.626 43.704 135 ; 
      RECT 43.168 130.626 43.272 135 ; 
      RECT 42.736 130.626 42.84 135 ; 
      RECT 42.304 130.626 42.408 135 ; 
      RECT 41.872 130.626 41.976 135 ; 
      RECT 41.44 130.626 41.544 135 ; 
      RECT 41.008 130.626 41.112 135 ; 
      RECT 40.576 130.626 40.68 135 ; 
      RECT 40.144 130.626 40.248 135 ; 
      RECT 39.712 130.626 39.816 135 ; 
      RECT 39.28 130.626 39.384 135 ; 
      RECT 38.848 130.626 38.952 135 ; 
      RECT 38.416 130.626 38.52 135 ; 
      RECT 37.984 130.626 38.088 135 ; 
      RECT 37.552 130.626 37.656 135 ; 
      RECT 36.7 130.626 37.008 135 ; 
      RECT 29.128 130.626 29.436 135 ; 
      RECT 28.48 130.626 28.584 135 ; 
      RECT 28.048 130.626 28.152 135 ; 
      RECT 27.616 130.626 27.72 135 ; 
      RECT 27.184 130.626 27.288 135 ; 
      RECT 26.752 130.626 26.856 135 ; 
      RECT 26.32 130.626 26.424 135 ; 
      RECT 25.888 130.626 25.992 135 ; 
      RECT 25.456 130.626 25.56 135 ; 
      RECT 25.024 130.626 25.128 135 ; 
      RECT 24.592 130.626 24.696 135 ; 
      RECT 24.16 130.626 24.264 135 ; 
      RECT 23.728 130.626 23.832 135 ; 
      RECT 23.296 130.626 23.4 135 ; 
      RECT 22.864 130.626 22.968 135 ; 
      RECT 22.432 130.626 22.536 135 ; 
      RECT 22 130.626 22.104 135 ; 
      RECT 21.568 130.626 21.672 135 ; 
      RECT 21.136 130.626 21.24 135 ; 
      RECT 20.704 130.626 20.808 135 ; 
      RECT 20.272 130.626 20.376 135 ; 
      RECT 19.84 130.626 19.944 135 ; 
      RECT 19.408 130.626 19.512 135 ; 
      RECT 18.976 130.626 19.08 135 ; 
      RECT 18.544 130.626 18.648 135 ; 
      RECT 18.112 130.626 18.216 135 ; 
      RECT 17.68 130.626 17.784 135 ; 
      RECT 17.248 130.626 17.352 135 ; 
      RECT 16.816 130.626 16.92 135 ; 
      RECT 16.384 130.626 16.488 135 ; 
      RECT 15.952 130.626 16.056 135 ; 
      RECT 15.52 130.626 15.624 135 ; 
      RECT 15.088 130.626 15.192 135 ; 
      RECT 14.656 130.626 14.76 135 ; 
      RECT 14.224 130.626 14.328 135 ; 
      RECT 13.792 130.626 13.896 135 ; 
      RECT 13.36 130.626 13.464 135 ; 
      RECT 12.928 130.626 13.032 135 ; 
      RECT 12.496 130.626 12.6 135 ; 
      RECT 12.064 130.626 12.168 135 ; 
      RECT 11.632 130.626 11.736 135 ; 
      RECT 11.2 130.626 11.304 135 ; 
      RECT 10.768 130.626 10.872 135 ; 
      RECT 10.336 130.626 10.44 135 ; 
      RECT 9.904 130.626 10.008 135 ; 
      RECT 9.472 130.626 9.576 135 ; 
      RECT 9.04 130.626 9.144 135 ; 
      RECT 8.608 130.626 8.712 135 ; 
      RECT 8.176 130.626 8.28 135 ; 
      RECT 7.744 130.626 7.848 135 ; 
      RECT 7.312 130.626 7.416 135 ; 
      RECT 6.88 130.626 6.984 135 ; 
      RECT 6.448 130.626 6.552 135 ; 
      RECT 6.016 130.626 6.12 135 ; 
      RECT 5.584 130.626 5.688 135 ; 
      RECT 5.152 130.626 5.256 135 ; 
      RECT 4.72 130.626 4.824 135 ; 
      RECT 4.288 130.626 4.392 135 ; 
      RECT 3.856 130.626 3.96 135 ; 
      RECT 3.424 130.626 3.528 135 ; 
      RECT 2.992 130.626 3.096 135 ; 
      RECT 2.56 130.626 2.664 135 ; 
      RECT 2.128 130.626 2.232 135 ; 
      RECT 1.696 130.626 1.8 135 ; 
      RECT 1.264 130.626 1.368 135 ; 
      RECT 0.832 130.626 0.936 135 ; 
      RECT 0.02 130.626 0.36 135 ; 
      RECT 34.564 134.946 35.076 139.32 ; 
      RECT 34.508 137.608 35.076 138.898 ; 
      RECT 33.916 136.516 34.164 139.32 ; 
      RECT 33.86 137.754 34.164 138.368 ; 
      RECT 33.916 134.946 34.02 139.32 ; 
      RECT 33.916 135.43 34.076 136.388 ; 
      RECT 33.916 134.946 34.164 135.302 ; 
      RECT 32.728 136.748 33.552 139.32 ; 
      RECT 33.448 134.946 33.552 139.32 ; 
      RECT 32.728 137.856 33.608 138.888 ; 
      RECT 32.728 134.946 33.12 139.32 ; 
      RECT 31.06 134.946 31.392 139.32 ; 
      RECT 31.06 135.3 31.448 139.042 ; 
      RECT 65.776 134.946 66.116 139.32 ; 
      RECT 65.2 134.946 65.304 139.32 ; 
      RECT 64.768 134.946 64.872 139.32 ; 
      RECT 64.336 134.946 64.44 139.32 ; 
      RECT 63.904 134.946 64.008 139.32 ; 
      RECT 63.472 134.946 63.576 139.32 ; 
      RECT 63.04 134.946 63.144 139.32 ; 
      RECT 62.608 134.946 62.712 139.32 ; 
      RECT 62.176 134.946 62.28 139.32 ; 
      RECT 61.744 134.946 61.848 139.32 ; 
      RECT 61.312 134.946 61.416 139.32 ; 
      RECT 60.88 134.946 60.984 139.32 ; 
      RECT 60.448 134.946 60.552 139.32 ; 
      RECT 60.016 134.946 60.12 139.32 ; 
      RECT 59.584 134.946 59.688 139.32 ; 
      RECT 59.152 134.946 59.256 139.32 ; 
      RECT 58.72 134.946 58.824 139.32 ; 
      RECT 58.288 134.946 58.392 139.32 ; 
      RECT 57.856 134.946 57.96 139.32 ; 
      RECT 57.424 134.946 57.528 139.32 ; 
      RECT 56.992 134.946 57.096 139.32 ; 
      RECT 56.56 134.946 56.664 139.32 ; 
      RECT 56.128 134.946 56.232 139.32 ; 
      RECT 55.696 134.946 55.8 139.32 ; 
      RECT 55.264 134.946 55.368 139.32 ; 
      RECT 54.832 134.946 54.936 139.32 ; 
      RECT 54.4 134.946 54.504 139.32 ; 
      RECT 53.968 134.946 54.072 139.32 ; 
      RECT 53.536 134.946 53.64 139.32 ; 
      RECT 53.104 134.946 53.208 139.32 ; 
      RECT 52.672 134.946 52.776 139.32 ; 
      RECT 52.24 134.946 52.344 139.32 ; 
      RECT 51.808 134.946 51.912 139.32 ; 
      RECT 51.376 134.946 51.48 139.32 ; 
      RECT 50.944 134.946 51.048 139.32 ; 
      RECT 50.512 134.946 50.616 139.32 ; 
      RECT 50.08 134.946 50.184 139.32 ; 
      RECT 49.648 134.946 49.752 139.32 ; 
      RECT 49.216 134.946 49.32 139.32 ; 
      RECT 48.784 134.946 48.888 139.32 ; 
      RECT 48.352 134.946 48.456 139.32 ; 
      RECT 47.92 134.946 48.024 139.32 ; 
      RECT 47.488 134.946 47.592 139.32 ; 
      RECT 47.056 134.946 47.16 139.32 ; 
      RECT 46.624 134.946 46.728 139.32 ; 
      RECT 46.192 134.946 46.296 139.32 ; 
      RECT 45.76 134.946 45.864 139.32 ; 
      RECT 45.328 134.946 45.432 139.32 ; 
      RECT 44.896 134.946 45 139.32 ; 
      RECT 44.464 134.946 44.568 139.32 ; 
      RECT 44.032 134.946 44.136 139.32 ; 
      RECT 43.6 134.946 43.704 139.32 ; 
      RECT 43.168 134.946 43.272 139.32 ; 
      RECT 42.736 134.946 42.84 139.32 ; 
      RECT 42.304 134.946 42.408 139.32 ; 
      RECT 41.872 134.946 41.976 139.32 ; 
      RECT 41.44 134.946 41.544 139.32 ; 
      RECT 41.008 134.946 41.112 139.32 ; 
      RECT 40.576 134.946 40.68 139.32 ; 
      RECT 40.144 134.946 40.248 139.32 ; 
      RECT 39.712 134.946 39.816 139.32 ; 
      RECT 39.28 134.946 39.384 139.32 ; 
      RECT 38.848 134.946 38.952 139.32 ; 
      RECT 38.416 134.946 38.52 139.32 ; 
      RECT 37.984 134.946 38.088 139.32 ; 
      RECT 37.552 134.946 37.656 139.32 ; 
      RECT 36.7 134.946 37.008 139.32 ; 
      RECT 29.128 134.946 29.436 139.32 ; 
      RECT 28.48 134.946 28.584 139.32 ; 
      RECT 28.048 134.946 28.152 139.32 ; 
      RECT 27.616 134.946 27.72 139.32 ; 
      RECT 27.184 134.946 27.288 139.32 ; 
      RECT 26.752 134.946 26.856 139.32 ; 
      RECT 26.32 134.946 26.424 139.32 ; 
      RECT 25.888 134.946 25.992 139.32 ; 
      RECT 25.456 134.946 25.56 139.32 ; 
      RECT 25.024 134.946 25.128 139.32 ; 
      RECT 24.592 134.946 24.696 139.32 ; 
      RECT 24.16 134.946 24.264 139.32 ; 
      RECT 23.728 134.946 23.832 139.32 ; 
      RECT 23.296 134.946 23.4 139.32 ; 
      RECT 22.864 134.946 22.968 139.32 ; 
      RECT 22.432 134.946 22.536 139.32 ; 
      RECT 22 134.946 22.104 139.32 ; 
      RECT 21.568 134.946 21.672 139.32 ; 
      RECT 21.136 134.946 21.24 139.32 ; 
      RECT 20.704 134.946 20.808 139.32 ; 
      RECT 20.272 134.946 20.376 139.32 ; 
      RECT 19.84 134.946 19.944 139.32 ; 
      RECT 19.408 134.946 19.512 139.32 ; 
      RECT 18.976 134.946 19.08 139.32 ; 
      RECT 18.544 134.946 18.648 139.32 ; 
      RECT 18.112 134.946 18.216 139.32 ; 
      RECT 17.68 134.946 17.784 139.32 ; 
      RECT 17.248 134.946 17.352 139.32 ; 
      RECT 16.816 134.946 16.92 139.32 ; 
      RECT 16.384 134.946 16.488 139.32 ; 
      RECT 15.952 134.946 16.056 139.32 ; 
      RECT 15.52 134.946 15.624 139.32 ; 
      RECT 15.088 134.946 15.192 139.32 ; 
      RECT 14.656 134.946 14.76 139.32 ; 
      RECT 14.224 134.946 14.328 139.32 ; 
      RECT 13.792 134.946 13.896 139.32 ; 
      RECT 13.36 134.946 13.464 139.32 ; 
      RECT 12.928 134.946 13.032 139.32 ; 
      RECT 12.496 134.946 12.6 139.32 ; 
      RECT 12.064 134.946 12.168 139.32 ; 
      RECT 11.632 134.946 11.736 139.32 ; 
      RECT 11.2 134.946 11.304 139.32 ; 
      RECT 10.768 134.946 10.872 139.32 ; 
      RECT 10.336 134.946 10.44 139.32 ; 
      RECT 9.904 134.946 10.008 139.32 ; 
      RECT 9.472 134.946 9.576 139.32 ; 
      RECT 9.04 134.946 9.144 139.32 ; 
      RECT 8.608 134.946 8.712 139.32 ; 
      RECT 8.176 134.946 8.28 139.32 ; 
      RECT 7.744 134.946 7.848 139.32 ; 
      RECT 7.312 134.946 7.416 139.32 ; 
      RECT 6.88 134.946 6.984 139.32 ; 
      RECT 6.448 134.946 6.552 139.32 ; 
      RECT 6.016 134.946 6.12 139.32 ; 
      RECT 5.584 134.946 5.688 139.32 ; 
      RECT 5.152 134.946 5.256 139.32 ; 
      RECT 4.72 134.946 4.824 139.32 ; 
      RECT 4.288 134.946 4.392 139.32 ; 
      RECT 3.856 134.946 3.96 139.32 ; 
      RECT 3.424 134.946 3.528 139.32 ; 
      RECT 2.992 134.946 3.096 139.32 ; 
      RECT 2.56 134.946 2.664 139.32 ; 
      RECT 2.128 134.946 2.232 139.32 ; 
      RECT 1.696 134.946 1.8 139.32 ; 
      RECT 1.264 134.946 1.368 139.32 ; 
      RECT 0.832 134.946 0.936 139.32 ; 
      RECT 0.02 134.946 0.36 139.32 ; 
      RECT 34.564 139.266 35.076 143.64 ; 
      RECT 34.508 141.928 35.076 143.218 ; 
      RECT 33.916 140.836 34.164 143.64 ; 
      RECT 33.86 142.074 34.164 142.688 ; 
      RECT 33.916 139.266 34.02 143.64 ; 
      RECT 33.916 139.75 34.076 140.708 ; 
      RECT 33.916 139.266 34.164 139.622 ; 
      RECT 32.728 141.068 33.552 143.64 ; 
      RECT 33.448 139.266 33.552 143.64 ; 
      RECT 32.728 142.176 33.608 143.208 ; 
      RECT 32.728 139.266 33.12 143.64 ; 
      RECT 31.06 139.266 31.392 143.64 ; 
      RECT 31.06 139.62 31.448 143.362 ; 
      RECT 65.776 139.266 66.116 143.64 ; 
      RECT 65.2 139.266 65.304 143.64 ; 
      RECT 64.768 139.266 64.872 143.64 ; 
      RECT 64.336 139.266 64.44 143.64 ; 
      RECT 63.904 139.266 64.008 143.64 ; 
      RECT 63.472 139.266 63.576 143.64 ; 
      RECT 63.04 139.266 63.144 143.64 ; 
      RECT 62.608 139.266 62.712 143.64 ; 
      RECT 62.176 139.266 62.28 143.64 ; 
      RECT 61.744 139.266 61.848 143.64 ; 
      RECT 61.312 139.266 61.416 143.64 ; 
      RECT 60.88 139.266 60.984 143.64 ; 
      RECT 60.448 139.266 60.552 143.64 ; 
      RECT 60.016 139.266 60.12 143.64 ; 
      RECT 59.584 139.266 59.688 143.64 ; 
      RECT 59.152 139.266 59.256 143.64 ; 
      RECT 58.72 139.266 58.824 143.64 ; 
      RECT 58.288 139.266 58.392 143.64 ; 
      RECT 57.856 139.266 57.96 143.64 ; 
      RECT 57.424 139.266 57.528 143.64 ; 
      RECT 56.992 139.266 57.096 143.64 ; 
      RECT 56.56 139.266 56.664 143.64 ; 
      RECT 56.128 139.266 56.232 143.64 ; 
      RECT 55.696 139.266 55.8 143.64 ; 
      RECT 55.264 139.266 55.368 143.64 ; 
      RECT 54.832 139.266 54.936 143.64 ; 
      RECT 54.4 139.266 54.504 143.64 ; 
      RECT 53.968 139.266 54.072 143.64 ; 
      RECT 53.536 139.266 53.64 143.64 ; 
      RECT 53.104 139.266 53.208 143.64 ; 
      RECT 52.672 139.266 52.776 143.64 ; 
      RECT 52.24 139.266 52.344 143.64 ; 
      RECT 51.808 139.266 51.912 143.64 ; 
      RECT 51.376 139.266 51.48 143.64 ; 
      RECT 50.944 139.266 51.048 143.64 ; 
      RECT 50.512 139.266 50.616 143.64 ; 
      RECT 50.08 139.266 50.184 143.64 ; 
      RECT 49.648 139.266 49.752 143.64 ; 
      RECT 49.216 139.266 49.32 143.64 ; 
      RECT 48.784 139.266 48.888 143.64 ; 
      RECT 48.352 139.266 48.456 143.64 ; 
      RECT 47.92 139.266 48.024 143.64 ; 
      RECT 47.488 139.266 47.592 143.64 ; 
      RECT 47.056 139.266 47.16 143.64 ; 
      RECT 46.624 139.266 46.728 143.64 ; 
      RECT 46.192 139.266 46.296 143.64 ; 
      RECT 45.76 139.266 45.864 143.64 ; 
      RECT 45.328 139.266 45.432 143.64 ; 
      RECT 44.896 139.266 45 143.64 ; 
      RECT 44.464 139.266 44.568 143.64 ; 
      RECT 44.032 139.266 44.136 143.64 ; 
      RECT 43.6 139.266 43.704 143.64 ; 
      RECT 43.168 139.266 43.272 143.64 ; 
      RECT 42.736 139.266 42.84 143.64 ; 
      RECT 42.304 139.266 42.408 143.64 ; 
      RECT 41.872 139.266 41.976 143.64 ; 
      RECT 41.44 139.266 41.544 143.64 ; 
      RECT 41.008 139.266 41.112 143.64 ; 
      RECT 40.576 139.266 40.68 143.64 ; 
      RECT 40.144 139.266 40.248 143.64 ; 
      RECT 39.712 139.266 39.816 143.64 ; 
      RECT 39.28 139.266 39.384 143.64 ; 
      RECT 38.848 139.266 38.952 143.64 ; 
      RECT 38.416 139.266 38.52 143.64 ; 
      RECT 37.984 139.266 38.088 143.64 ; 
      RECT 37.552 139.266 37.656 143.64 ; 
      RECT 36.7 139.266 37.008 143.64 ; 
      RECT 29.128 139.266 29.436 143.64 ; 
      RECT 28.48 139.266 28.584 143.64 ; 
      RECT 28.048 139.266 28.152 143.64 ; 
      RECT 27.616 139.266 27.72 143.64 ; 
      RECT 27.184 139.266 27.288 143.64 ; 
      RECT 26.752 139.266 26.856 143.64 ; 
      RECT 26.32 139.266 26.424 143.64 ; 
      RECT 25.888 139.266 25.992 143.64 ; 
      RECT 25.456 139.266 25.56 143.64 ; 
      RECT 25.024 139.266 25.128 143.64 ; 
      RECT 24.592 139.266 24.696 143.64 ; 
      RECT 24.16 139.266 24.264 143.64 ; 
      RECT 23.728 139.266 23.832 143.64 ; 
      RECT 23.296 139.266 23.4 143.64 ; 
      RECT 22.864 139.266 22.968 143.64 ; 
      RECT 22.432 139.266 22.536 143.64 ; 
      RECT 22 139.266 22.104 143.64 ; 
      RECT 21.568 139.266 21.672 143.64 ; 
      RECT 21.136 139.266 21.24 143.64 ; 
      RECT 20.704 139.266 20.808 143.64 ; 
      RECT 20.272 139.266 20.376 143.64 ; 
      RECT 19.84 139.266 19.944 143.64 ; 
      RECT 19.408 139.266 19.512 143.64 ; 
      RECT 18.976 139.266 19.08 143.64 ; 
      RECT 18.544 139.266 18.648 143.64 ; 
      RECT 18.112 139.266 18.216 143.64 ; 
      RECT 17.68 139.266 17.784 143.64 ; 
      RECT 17.248 139.266 17.352 143.64 ; 
      RECT 16.816 139.266 16.92 143.64 ; 
      RECT 16.384 139.266 16.488 143.64 ; 
      RECT 15.952 139.266 16.056 143.64 ; 
      RECT 15.52 139.266 15.624 143.64 ; 
      RECT 15.088 139.266 15.192 143.64 ; 
      RECT 14.656 139.266 14.76 143.64 ; 
      RECT 14.224 139.266 14.328 143.64 ; 
      RECT 13.792 139.266 13.896 143.64 ; 
      RECT 13.36 139.266 13.464 143.64 ; 
      RECT 12.928 139.266 13.032 143.64 ; 
      RECT 12.496 139.266 12.6 143.64 ; 
      RECT 12.064 139.266 12.168 143.64 ; 
      RECT 11.632 139.266 11.736 143.64 ; 
      RECT 11.2 139.266 11.304 143.64 ; 
      RECT 10.768 139.266 10.872 143.64 ; 
      RECT 10.336 139.266 10.44 143.64 ; 
      RECT 9.904 139.266 10.008 143.64 ; 
      RECT 9.472 139.266 9.576 143.64 ; 
      RECT 9.04 139.266 9.144 143.64 ; 
      RECT 8.608 139.266 8.712 143.64 ; 
      RECT 8.176 139.266 8.28 143.64 ; 
      RECT 7.744 139.266 7.848 143.64 ; 
      RECT 7.312 139.266 7.416 143.64 ; 
      RECT 6.88 139.266 6.984 143.64 ; 
      RECT 6.448 139.266 6.552 143.64 ; 
      RECT 6.016 139.266 6.12 143.64 ; 
      RECT 5.584 139.266 5.688 143.64 ; 
      RECT 5.152 139.266 5.256 143.64 ; 
      RECT 4.72 139.266 4.824 143.64 ; 
      RECT 4.288 139.266 4.392 143.64 ; 
      RECT 3.856 139.266 3.96 143.64 ; 
      RECT 3.424 139.266 3.528 143.64 ; 
      RECT 2.992 139.266 3.096 143.64 ; 
      RECT 2.56 139.266 2.664 143.64 ; 
      RECT 2.128 139.266 2.232 143.64 ; 
      RECT 1.696 139.266 1.8 143.64 ; 
      RECT 1.264 139.266 1.368 143.64 ; 
      RECT 0.832 139.266 0.936 143.64 ; 
      RECT 0.02 139.266 0.36 143.64 ; 
      RECT 34.564 143.586 35.076 147.96 ; 
      RECT 34.508 146.248 35.076 147.538 ; 
      RECT 33.916 145.156 34.164 147.96 ; 
      RECT 33.86 146.394 34.164 147.008 ; 
      RECT 33.916 143.586 34.02 147.96 ; 
      RECT 33.916 144.07 34.076 145.028 ; 
      RECT 33.916 143.586 34.164 143.942 ; 
      RECT 32.728 145.388 33.552 147.96 ; 
      RECT 33.448 143.586 33.552 147.96 ; 
      RECT 32.728 146.496 33.608 147.528 ; 
      RECT 32.728 143.586 33.12 147.96 ; 
      RECT 31.06 143.586 31.392 147.96 ; 
      RECT 31.06 143.94 31.448 147.682 ; 
      RECT 65.776 143.586 66.116 147.96 ; 
      RECT 65.2 143.586 65.304 147.96 ; 
      RECT 64.768 143.586 64.872 147.96 ; 
      RECT 64.336 143.586 64.44 147.96 ; 
      RECT 63.904 143.586 64.008 147.96 ; 
      RECT 63.472 143.586 63.576 147.96 ; 
      RECT 63.04 143.586 63.144 147.96 ; 
      RECT 62.608 143.586 62.712 147.96 ; 
      RECT 62.176 143.586 62.28 147.96 ; 
      RECT 61.744 143.586 61.848 147.96 ; 
      RECT 61.312 143.586 61.416 147.96 ; 
      RECT 60.88 143.586 60.984 147.96 ; 
      RECT 60.448 143.586 60.552 147.96 ; 
      RECT 60.016 143.586 60.12 147.96 ; 
      RECT 59.584 143.586 59.688 147.96 ; 
      RECT 59.152 143.586 59.256 147.96 ; 
      RECT 58.72 143.586 58.824 147.96 ; 
      RECT 58.288 143.586 58.392 147.96 ; 
      RECT 57.856 143.586 57.96 147.96 ; 
      RECT 57.424 143.586 57.528 147.96 ; 
      RECT 56.992 143.586 57.096 147.96 ; 
      RECT 56.56 143.586 56.664 147.96 ; 
      RECT 56.128 143.586 56.232 147.96 ; 
      RECT 55.696 143.586 55.8 147.96 ; 
      RECT 55.264 143.586 55.368 147.96 ; 
      RECT 54.832 143.586 54.936 147.96 ; 
      RECT 54.4 143.586 54.504 147.96 ; 
      RECT 53.968 143.586 54.072 147.96 ; 
      RECT 53.536 143.586 53.64 147.96 ; 
      RECT 53.104 143.586 53.208 147.96 ; 
      RECT 52.672 143.586 52.776 147.96 ; 
      RECT 52.24 143.586 52.344 147.96 ; 
      RECT 51.808 143.586 51.912 147.96 ; 
      RECT 51.376 143.586 51.48 147.96 ; 
      RECT 50.944 143.586 51.048 147.96 ; 
      RECT 50.512 143.586 50.616 147.96 ; 
      RECT 50.08 143.586 50.184 147.96 ; 
      RECT 49.648 143.586 49.752 147.96 ; 
      RECT 49.216 143.586 49.32 147.96 ; 
      RECT 48.784 143.586 48.888 147.96 ; 
      RECT 48.352 143.586 48.456 147.96 ; 
      RECT 47.92 143.586 48.024 147.96 ; 
      RECT 47.488 143.586 47.592 147.96 ; 
      RECT 47.056 143.586 47.16 147.96 ; 
      RECT 46.624 143.586 46.728 147.96 ; 
      RECT 46.192 143.586 46.296 147.96 ; 
      RECT 45.76 143.586 45.864 147.96 ; 
      RECT 45.328 143.586 45.432 147.96 ; 
      RECT 44.896 143.586 45 147.96 ; 
      RECT 44.464 143.586 44.568 147.96 ; 
      RECT 44.032 143.586 44.136 147.96 ; 
      RECT 43.6 143.586 43.704 147.96 ; 
      RECT 43.168 143.586 43.272 147.96 ; 
      RECT 42.736 143.586 42.84 147.96 ; 
      RECT 42.304 143.586 42.408 147.96 ; 
      RECT 41.872 143.586 41.976 147.96 ; 
      RECT 41.44 143.586 41.544 147.96 ; 
      RECT 41.008 143.586 41.112 147.96 ; 
      RECT 40.576 143.586 40.68 147.96 ; 
      RECT 40.144 143.586 40.248 147.96 ; 
      RECT 39.712 143.586 39.816 147.96 ; 
      RECT 39.28 143.586 39.384 147.96 ; 
      RECT 38.848 143.586 38.952 147.96 ; 
      RECT 38.416 143.586 38.52 147.96 ; 
      RECT 37.984 143.586 38.088 147.96 ; 
      RECT 37.552 143.586 37.656 147.96 ; 
      RECT 36.7 143.586 37.008 147.96 ; 
      RECT 29.128 143.586 29.436 147.96 ; 
      RECT 28.48 143.586 28.584 147.96 ; 
      RECT 28.048 143.586 28.152 147.96 ; 
      RECT 27.616 143.586 27.72 147.96 ; 
      RECT 27.184 143.586 27.288 147.96 ; 
      RECT 26.752 143.586 26.856 147.96 ; 
      RECT 26.32 143.586 26.424 147.96 ; 
      RECT 25.888 143.586 25.992 147.96 ; 
      RECT 25.456 143.586 25.56 147.96 ; 
      RECT 25.024 143.586 25.128 147.96 ; 
      RECT 24.592 143.586 24.696 147.96 ; 
      RECT 24.16 143.586 24.264 147.96 ; 
      RECT 23.728 143.586 23.832 147.96 ; 
      RECT 23.296 143.586 23.4 147.96 ; 
      RECT 22.864 143.586 22.968 147.96 ; 
      RECT 22.432 143.586 22.536 147.96 ; 
      RECT 22 143.586 22.104 147.96 ; 
      RECT 21.568 143.586 21.672 147.96 ; 
      RECT 21.136 143.586 21.24 147.96 ; 
      RECT 20.704 143.586 20.808 147.96 ; 
      RECT 20.272 143.586 20.376 147.96 ; 
      RECT 19.84 143.586 19.944 147.96 ; 
      RECT 19.408 143.586 19.512 147.96 ; 
      RECT 18.976 143.586 19.08 147.96 ; 
      RECT 18.544 143.586 18.648 147.96 ; 
      RECT 18.112 143.586 18.216 147.96 ; 
      RECT 17.68 143.586 17.784 147.96 ; 
      RECT 17.248 143.586 17.352 147.96 ; 
      RECT 16.816 143.586 16.92 147.96 ; 
      RECT 16.384 143.586 16.488 147.96 ; 
      RECT 15.952 143.586 16.056 147.96 ; 
      RECT 15.52 143.586 15.624 147.96 ; 
      RECT 15.088 143.586 15.192 147.96 ; 
      RECT 14.656 143.586 14.76 147.96 ; 
      RECT 14.224 143.586 14.328 147.96 ; 
      RECT 13.792 143.586 13.896 147.96 ; 
      RECT 13.36 143.586 13.464 147.96 ; 
      RECT 12.928 143.586 13.032 147.96 ; 
      RECT 12.496 143.586 12.6 147.96 ; 
      RECT 12.064 143.586 12.168 147.96 ; 
      RECT 11.632 143.586 11.736 147.96 ; 
      RECT 11.2 143.586 11.304 147.96 ; 
      RECT 10.768 143.586 10.872 147.96 ; 
      RECT 10.336 143.586 10.44 147.96 ; 
      RECT 9.904 143.586 10.008 147.96 ; 
      RECT 9.472 143.586 9.576 147.96 ; 
      RECT 9.04 143.586 9.144 147.96 ; 
      RECT 8.608 143.586 8.712 147.96 ; 
      RECT 8.176 143.586 8.28 147.96 ; 
      RECT 7.744 143.586 7.848 147.96 ; 
      RECT 7.312 143.586 7.416 147.96 ; 
      RECT 6.88 143.586 6.984 147.96 ; 
      RECT 6.448 143.586 6.552 147.96 ; 
      RECT 6.016 143.586 6.12 147.96 ; 
      RECT 5.584 143.586 5.688 147.96 ; 
      RECT 5.152 143.586 5.256 147.96 ; 
      RECT 4.72 143.586 4.824 147.96 ; 
      RECT 4.288 143.586 4.392 147.96 ; 
      RECT 3.856 143.586 3.96 147.96 ; 
      RECT 3.424 143.586 3.528 147.96 ; 
      RECT 2.992 143.586 3.096 147.96 ; 
      RECT 2.56 143.586 2.664 147.96 ; 
      RECT 2.128 143.586 2.232 147.96 ; 
      RECT 1.696 143.586 1.8 147.96 ; 
      RECT 1.264 143.586 1.368 147.96 ; 
      RECT 0.832 143.586 0.936 147.96 ; 
      RECT 0.02 143.586 0.36 147.96 ; 
      RECT 34.564 147.906 35.076 152.28 ; 
      RECT 34.508 150.568 35.076 151.858 ; 
      RECT 33.916 149.476 34.164 152.28 ; 
      RECT 33.86 150.714 34.164 151.328 ; 
      RECT 33.916 147.906 34.02 152.28 ; 
      RECT 33.916 148.39 34.076 149.348 ; 
      RECT 33.916 147.906 34.164 148.262 ; 
      RECT 32.728 149.708 33.552 152.28 ; 
      RECT 33.448 147.906 33.552 152.28 ; 
      RECT 32.728 150.816 33.608 151.848 ; 
      RECT 32.728 147.906 33.12 152.28 ; 
      RECT 31.06 147.906 31.392 152.28 ; 
      RECT 31.06 148.26 31.448 152.002 ; 
      RECT 65.776 147.906 66.116 152.28 ; 
      RECT 65.2 147.906 65.304 152.28 ; 
      RECT 64.768 147.906 64.872 152.28 ; 
      RECT 64.336 147.906 64.44 152.28 ; 
      RECT 63.904 147.906 64.008 152.28 ; 
      RECT 63.472 147.906 63.576 152.28 ; 
      RECT 63.04 147.906 63.144 152.28 ; 
      RECT 62.608 147.906 62.712 152.28 ; 
      RECT 62.176 147.906 62.28 152.28 ; 
      RECT 61.744 147.906 61.848 152.28 ; 
      RECT 61.312 147.906 61.416 152.28 ; 
      RECT 60.88 147.906 60.984 152.28 ; 
      RECT 60.448 147.906 60.552 152.28 ; 
      RECT 60.016 147.906 60.12 152.28 ; 
      RECT 59.584 147.906 59.688 152.28 ; 
      RECT 59.152 147.906 59.256 152.28 ; 
      RECT 58.72 147.906 58.824 152.28 ; 
      RECT 58.288 147.906 58.392 152.28 ; 
      RECT 57.856 147.906 57.96 152.28 ; 
      RECT 57.424 147.906 57.528 152.28 ; 
      RECT 56.992 147.906 57.096 152.28 ; 
      RECT 56.56 147.906 56.664 152.28 ; 
      RECT 56.128 147.906 56.232 152.28 ; 
      RECT 55.696 147.906 55.8 152.28 ; 
      RECT 55.264 147.906 55.368 152.28 ; 
      RECT 54.832 147.906 54.936 152.28 ; 
      RECT 54.4 147.906 54.504 152.28 ; 
      RECT 53.968 147.906 54.072 152.28 ; 
      RECT 53.536 147.906 53.64 152.28 ; 
      RECT 53.104 147.906 53.208 152.28 ; 
      RECT 52.672 147.906 52.776 152.28 ; 
      RECT 52.24 147.906 52.344 152.28 ; 
      RECT 51.808 147.906 51.912 152.28 ; 
      RECT 51.376 147.906 51.48 152.28 ; 
      RECT 50.944 147.906 51.048 152.28 ; 
      RECT 50.512 147.906 50.616 152.28 ; 
      RECT 50.08 147.906 50.184 152.28 ; 
      RECT 49.648 147.906 49.752 152.28 ; 
      RECT 49.216 147.906 49.32 152.28 ; 
      RECT 48.784 147.906 48.888 152.28 ; 
      RECT 48.352 147.906 48.456 152.28 ; 
      RECT 47.92 147.906 48.024 152.28 ; 
      RECT 47.488 147.906 47.592 152.28 ; 
      RECT 47.056 147.906 47.16 152.28 ; 
      RECT 46.624 147.906 46.728 152.28 ; 
      RECT 46.192 147.906 46.296 152.28 ; 
      RECT 45.76 147.906 45.864 152.28 ; 
      RECT 45.328 147.906 45.432 152.28 ; 
      RECT 44.896 147.906 45 152.28 ; 
      RECT 44.464 147.906 44.568 152.28 ; 
      RECT 44.032 147.906 44.136 152.28 ; 
      RECT 43.6 147.906 43.704 152.28 ; 
      RECT 43.168 147.906 43.272 152.28 ; 
      RECT 42.736 147.906 42.84 152.28 ; 
      RECT 42.304 147.906 42.408 152.28 ; 
      RECT 41.872 147.906 41.976 152.28 ; 
      RECT 41.44 147.906 41.544 152.28 ; 
      RECT 41.008 147.906 41.112 152.28 ; 
      RECT 40.576 147.906 40.68 152.28 ; 
      RECT 40.144 147.906 40.248 152.28 ; 
      RECT 39.712 147.906 39.816 152.28 ; 
      RECT 39.28 147.906 39.384 152.28 ; 
      RECT 38.848 147.906 38.952 152.28 ; 
      RECT 38.416 147.906 38.52 152.28 ; 
      RECT 37.984 147.906 38.088 152.28 ; 
      RECT 37.552 147.906 37.656 152.28 ; 
      RECT 36.7 147.906 37.008 152.28 ; 
      RECT 29.128 147.906 29.436 152.28 ; 
      RECT 28.48 147.906 28.584 152.28 ; 
      RECT 28.048 147.906 28.152 152.28 ; 
      RECT 27.616 147.906 27.72 152.28 ; 
      RECT 27.184 147.906 27.288 152.28 ; 
      RECT 26.752 147.906 26.856 152.28 ; 
      RECT 26.32 147.906 26.424 152.28 ; 
      RECT 25.888 147.906 25.992 152.28 ; 
      RECT 25.456 147.906 25.56 152.28 ; 
      RECT 25.024 147.906 25.128 152.28 ; 
      RECT 24.592 147.906 24.696 152.28 ; 
      RECT 24.16 147.906 24.264 152.28 ; 
      RECT 23.728 147.906 23.832 152.28 ; 
      RECT 23.296 147.906 23.4 152.28 ; 
      RECT 22.864 147.906 22.968 152.28 ; 
      RECT 22.432 147.906 22.536 152.28 ; 
      RECT 22 147.906 22.104 152.28 ; 
      RECT 21.568 147.906 21.672 152.28 ; 
      RECT 21.136 147.906 21.24 152.28 ; 
      RECT 20.704 147.906 20.808 152.28 ; 
      RECT 20.272 147.906 20.376 152.28 ; 
      RECT 19.84 147.906 19.944 152.28 ; 
      RECT 19.408 147.906 19.512 152.28 ; 
      RECT 18.976 147.906 19.08 152.28 ; 
      RECT 18.544 147.906 18.648 152.28 ; 
      RECT 18.112 147.906 18.216 152.28 ; 
      RECT 17.68 147.906 17.784 152.28 ; 
      RECT 17.248 147.906 17.352 152.28 ; 
      RECT 16.816 147.906 16.92 152.28 ; 
      RECT 16.384 147.906 16.488 152.28 ; 
      RECT 15.952 147.906 16.056 152.28 ; 
      RECT 15.52 147.906 15.624 152.28 ; 
      RECT 15.088 147.906 15.192 152.28 ; 
      RECT 14.656 147.906 14.76 152.28 ; 
      RECT 14.224 147.906 14.328 152.28 ; 
      RECT 13.792 147.906 13.896 152.28 ; 
      RECT 13.36 147.906 13.464 152.28 ; 
      RECT 12.928 147.906 13.032 152.28 ; 
      RECT 12.496 147.906 12.6 152.28 ; 
      RECT 12.064 147.906 12.168 152.28 ; 
      RECT 11.632 147.906 11.736 152.28 ; 
      RECT 11.2 147.906 11.304 152.28 ; 
      RECT 10.768 147.906 10.872 152.28 ; 
      RECT 10.336 147.906 10.44 152.28 ; 
      RECT 9.904 147.906 10.008 152.28 ; 
      RECT 9.472 147.906 9.576 152.28 ; 
      RECT 9.04 147.906 9.144 152.28 ; 
      RECT 8.608 147.906 8.712 152.28 ; 
      RECT 8.176 147.906 8.28 152.28 ; 
      RECT 7.744 147.906 7.848 152.28 ; 
      RECT 7.312 147.906 7.416 152.28 ; 
      RECT 6.88 147.906 6.984 152.28 ; 
      RECT 6.448 147.906 6.552 152.28 ; 
      RECT 6.016 147.906 6.12 152.28 ; 
      RECT 5.584 147.906 5.688 152.28 ; 
      RECT 5.152 147.906 5.256 152.28 ; 
      RECT 4.72 147.906 4.824 152.28 ; 
      RECT 4.288 147.906 4.392 152.28 ; 
      RECT 3.856 147.906 3.96 152.28 ; 
      RECT 3.424 147.906 3.528 152.28 ; 
      RECT 2.992 147.906 3.096 152.28 ; 
      RECT 2.56 147.906 2.664 152.28 ; 
      RECT 2.128 147.906 2.232 152.28 ; 
      RECT 1.696 147.906 1.8 152.28 ; 
      RECT 1.264 147.906 1.368 152.28 ; 
      RECT 0.832 147.906 0.936 152.28 ; 
      RECT 0.02 147.906 0.36 152.28 ; 
      RECT 34.564 152.226 35.076 156.6 ; 
      RECT 34.508 154.888 35.076 156.178 ; 
      RECT 33.916 153.796 34.164 156.6 ; 
      RECT 33.86 155.034 34.164 155.648 ; 
      RECT 33.916 152.226 34.02 156.6 ; 
      RECT 33.916 152.71 34.076 153.668 ; 
      RECT 33.916 152.226 34.164 152.582 ; 
      RECT 32.728 154.028 33.552 156.6 ; 
      RECT 33.448 152.226 33.552 156.6 ; 
      RECT 32.728 155.136 33.608 156.168 ; 
      RECT 32.728 152.226 33.12 156.6 ; 
      RECT 31.06 152.226 31.392 156.6 ; 
      RECT 31.06 152.58 31.448 156.322 ; 
      RECT 65.776 152.226 66.116 156.6 ; 
      RECT 65.2 152.226 65.304 156.6 ; 
      RECT 64.768 152.226 64.872 156.6 ; 
      RECT 64.336 152.226 64.44 156.6 ; 
      RECT 63.904 152.226 64.008 156.6 ; 
      RECT 63.472 152.226 63.576 156.6 ; 
      RECT 63.04 152.226 63.144 156.6 ; 
      RECT 62.608 152.226 62.712 156.6 ; 
      RECT 62.176 152.226 62.28 156.6 ; 
      RECT 61.744 152.226 61.848 156.6 ; 
      RECT 61.312 152.226 61.416 156.6 ; 
      RECT 60.88 152.226 60.984 156.6 ; 
      RECT 60.448 152.226 60.552 156.6 ; 
      RECT 60.016 152.226 60.12 156.6 ; 
      RECT 59.584 152.226 59.688 156.6 ; 
      RECT 59.152 152.226 59.256 156.6 ; 
      RECT 58.72 152.226 58.824 156.6 ; 
      RECT 58.288 152.226 58.392 156.6 ; 
      RECT 57.856 152.226 57.96 156.6 ; 
      RECT 57.424 152.226 57.528 156.6 ; 
      RECT 56.992 152.226 57.096 156.6 ; 
      RECT 56.56 152.226 56.664 156.6 ; 
      RECT 56.128 152.226 56.232 156.6 ; 
      RECT 55.696 152.226 55.8 156.6 ; 
      RECT 55.264 152.226 55.368 156.6 ; 
      RECT 54.832 152.226 54.936 156.6 ; 
      RECT 54.4 152.226 54.504 156.6 ; 
      RECT 53.968 152.226 54.072 156.6 ; 
      RECT 53.536 152.226 53.64 156.6 ; 
      RECT 53.104 152.226 53.208 156.6 ; 
      RECT 52.672 152.226 52.776 156.6 ; 
      RECT 52.24 152.226 52.344 156.6 ; 
      RECT 51.808 152.226 51.912 156.6 ; 
      RECT 51.376 152.226 51.48 156.6 ; 
      RECT 50.944 152.226 51.048 156.6 ; 
      RECT 50.512 152.226 50.616 156.6 ; 
      RECT 50.08 152.226 50.184 156.6 ; 
      RECT 49.648 152.226 49.752 156.6 ; 
      RECT 49.216 152.226 49.32 156.6 ; 
      RECT 48.784 152.226 48.888 156.6 ; 
      RECT 48.352 152.226 48.456 156.6 ; 
      RECT 47.92 152.226 48.024 156.6 ; 
      RECT 47.488 152.226 47.592 156.6 ; 
      RECT 47.056 152.226 47.16 156.6 ; 
      RECT 46.624 152.226 46.728 156.6 ; 
      RECT 46.192 152.226 46.296 156.6 ; 
      RECT 45.76 152.226 45.864 156.6 ; 
      RECT 45.328 152.226 45.432 156.6 ; 
      RECT 44.896 152.226 45 156.6 ; 
      RECT 44.464 152.226 44.568 156.6 ; 
      RECT 44.032 152.226 44.136 156.6 ; 
      RECT 43.6 152.226 43.704 156.6 ; 
      RECT 43.168 152.226 43.272 156.6 ; 
      RECT 42.736 152.226 42.84 156.6 ; 
      RECT 42.304 152.226 42.408 156.6 ; 
      RECT 41.872 152.226 41.976 156.6 ; 
      RECT 41.44 152.226 41.544 156.6 ; 
      RECT 41.008 152.226 41.112 156.6 ; 
      RECT 40.576 152.226 40.68 156.6 ; 
      RECT 40.144 152.226 40.248 156.6 ; 
      RECT 39.712 152.226 39.816 156.6 ; 
      RECT 39.28 152.226 39.384 156.6 ; 
      RECT 38.848 152.226 38.952 156.6 ; 
      RECT 38.416 152.226 38.52 156.6 ; 
      RECT 37.984 152.226 38.088 156.6 ; 
      RECT 37.552 152.226 37.656 156.6 ; 
      RECT 36.7 152.226 37.008 156.6 ; 
      RECT 29.128 152.226 29.436 156.6 ; 
      RECT 28.48 152.226 28.584 156.6 ; 
      RECT 28.048 152.226 28.152 156.6 ; 
      RECT 27.616 152.226 27.72 156.6 ; 
      RECT 27.184 152.226 27.288 156.6 ; 
      RECT 26.752 152.226 26.856 156.6 ; 
      RECT 26.32 152.226 26.424 156.6 ; 
      RECT 25.888 152.226 25.992 156.6 ; 
      RECT 25.456 152.226 25.56 156.6 ; 
      RECT 25.024 152.226 25.128 156.6 ; 
      RECT 24.592 152.226 24.696 156.6 ; 
      RECT 24.16 152.226 24.264 156.6 ; 
      RECT 23.728 152.226 23.832 156.6 ; 
      RECT 23.296 152.226 23.4 156.6 ; 
      RECT 22.864 152.226 22.968 156.6 ; 
      RECT 22.432 152.226 22.536 156.6 ; 
      RECT 22 152.226 22.104 156.6 ; 
      RECT 21.568 152.226 21.672 156.6 ; 
      RECT 21.136 152.226 21.24 156.6 ; 
      RECT 20.704 152.226 20.808 156.6 ; 
      RECT 20.272 152.226 20.376 156.6 ; 
      RECT 19.84 152.226 19.944 156.6 ; 
      RECT 19.408 152.226 19.512 156.6 ; 
      RECT 18.976 152.226 19.08 156.6 ; 
      RECT 18.544 152.226 18.648 156.6 ; 
      RECT 18.112 152.226 18.216 156.6 ; 
      RECT 17.68 152.226 17.784 156.6 ; 
      RECT 17.248 152.226 17.352 156.6 ; 
      RECT 16.816 152.226 16.92 156.6 ; 
      RECT 16.384 152.226 16.488 156.6 ; 
      RECT 15.952 152.226 16.056 156.6 ; 
      RECT 15.52 152.226 15.624 156.6 ; 
      RECT 15.088 152.226 15.192 156.6 ; 
      RECT 14.656 152.226 14.76 156.6 ; 
      RECT 14.224 152.226 14.328 156.6 ; 
      RECT 13.792 152.226 13.896 156.6 ; 
      RECT 13.36 152.226 13.464 156.6 ; 
      RECT 12.928 152.226 13.032 156.6 ; 
      RECT 12.496 152.226 12.6 156.6 ; 
      RECT 12.064 152.226 12.168 156.6 ; 
      RECT 11.632 152.226 11.736 156.6 ; 
      RECT 11.2 152.226 11.304 156.6 ; 
      RECT 10.768 152.226 10.872 156.6 ; 
      RECT 10.336 152.226 10.44 156.6 ; 
      RECT 9.904 152.226 10.008 156.6 ; 
      RECT 9.472 152.226 9.576 156.6 ; 
      RECT 9.04 152.226 9.144 156.6 ; 
      RECT 8.608 152.226 8.712 156.6 ; 
      RECT 8.176 152.226 8.28 156.6 ; 
      RECT 7.744 152.226 7.848 156.6 ; 
      RECT 7.312 152.226 7.416 156.6 ; 
      RECT 6.88 152.226 6.984 156.6 ; 
      RECT 6.448 152.226 6.552 156.6 ; 
      RECT 6.016 152.226 6.12 156.6 ; 
      RECT 5.584 152.226 5.688 156.6 ; 
      RECT 5.152 152.226 5.256 156.6 ; 
      RECT 4.72 152.226 4.824 156.6 ; 
      RECT 4.288 152.226 4.392 156.6 ; 
      RECT 3.856 152.226 3.96 156.6 ; 
      RECT 3.424 152.226 3.528 156.6 ; 
      RECT 2.992 152.226 3.096 156.6 ; 
      RECT 2.56 152.226 2.664 156.6 ; 
      RECT 2.128 152.226 2.232 156.6 ; 
      RECT 1.696 152.226 1.8 156.6 ; 
      RECT 1.264 152.226 1.368 156.6 ; 
      RECT 0.832 152.226 0.936 156.6 ; 
      RECT 0.02 152.226 0.36 156.6 ; 
      RECT 34.564 156.546 35.076 160.92 ; 
      RECT 34.508 159.208 35.076 160.498 ; 
      RECT 33.916 158.116 34.164 160.92 ; 
      RECT 33.86 159.354 34.164 159.968 ; 
      RECT 33.916 156.546 34.02 160.92 ; 
      RECT 33.916 157.03 34.076 157.988 ; 
      RECT 33.916 156.546 34.164 156.902 ; 
      RECT 32.728 158.348 33.552 160.92 ; 
      RECT 33.448 156.546 33.552 160.92 ; 
      RECT 32.728 159.456 33.608 160.488 ; 
      RECT 32.728 156.546 33.12 160.92 ; 
      RECT 31.06 156.546 31.392 160.92 ; 
      RECT 31.06 156.9 31.448 160.642 ; 
      RECT 65.776 156.546 66.116 160.92 ; 
      RECT 65.2 156.546 65.304 160.92 ; 
      RECT 64.768 156.546 64.872 160.92 ; 
      RECT 64.336 156.546 64.44 160.92 ; 
      RECT 63.904 156.546 64.008 160.92 ; 
      RECT 63.472 156.546 63.576 160.92 ; 
      RECT 63.04 156.546 63.144 160.92 ; 
      RECT 62.608 156.546 62.712 160.92 ; 
      RECT 62.176 156.546 62.28 160.92 ; 
      RECT 61.744 156.546 61.848 160.92 ; 
      RECT 61.312 156.546 61.416 160.92 ; 
      RECT 60.88 156.546 60.984 160.92 ; 
      RECT 60.448 156.546 60.552 160.92 ; 
      RECT 60.016 156.546 60.12 160.92 ; 
      RECT 59.584 156.546 59.688 160.92 ; 
      RECT 59.152 156.546 59.256 160.92 ; 
      RECT 58.72 156.546 58.824 160.92 ; 
      RECT 58.288 156.546 58.392 160.92 ; 
      RECT 57.856 156.546 57.96 160.92 ; 
      RECT 57.424 156.546 57.528 160.92 ; 
      RECT 56.992 156.546 57.096 160.92 ; 
      RECT 56.56 156.546 56.664 160.92 ; 
      RECT 56.128 156.546 56.232 160.92 ; 
      RECT 55.696 156.546 55.8 160.92 ; 
      RECT 55.264 156.546 55.368 160.92 ; 
      RECT 54.832 156.546 54.936 160.92 ; 
      RECT 54.4 156.546 54.504 160.92 ; 
      RECT 53.968 156.546 54.072 160.92 ; 
      RECT 53.536 156.546 53.64 160.92 ; 
      RECT 53.104 156.546 53.208 160.92 ; 
      RECT 52.672 156.546 52.776 160.92 ; 
      RECT 52.24 156.546 52.344 160.92 ; 
      RECT 51.808 156.546 51.912 160.92 ; 
      RECT 51.376 156.546 51.48 160.92 ; 
      RECT 50.944 156.546 51.048 160.92 ; 
      RECT 50.512 156.546 50.616 160.92 ; 
      RECT 50.08 156.546 50.184 160.92 ; 
      RECT 49.648 156.546 49.752 160.92 ; 
      RECT 49.216 156.546 49.32 160.92 ; 
      RECT 48.784 156.546 48.888 160.92 ; 
      RECT 48.352 156.546 48.456 160.92 ; 
      RECT 47.92 156.546 48.024 160.92 ; 
      RECT 47.488 156.546 47.592 160.92 ; 
      RECT 47.056 156.546 47.16 160.92 ; 
      RECT 46.624 156.546 46.728 160.92 ; 
      RECT 46.192 156.546 46.296 160.92 ; 
      RECT 45.76 156.546 45.864 160.92 ; 
      RECT 45.328 156.546 45.432 160.92 ; 
      RECT 44.896 156.546 45 160.92 ; 
      RECT 44.464 156.546 44.568 160.92 ; 
      RECT 44.032 156.546 44.136 160.92 ; 
      RECT 43.6 156.546 43.704 160.92 ; 
      RECT 43.168 156.546 43.272 160.92 ; 
      RECT 42.736 156.546 42.84 160.92 ; 
      RECT 42.304 156.546 42.408 160.92 ; 
      RECT 41.872 156.546 41.976 160.92 ; 
      RECT 41.44 156.546 41.544 160.92 ; 
      RECT 41.008 156.546 41.112 160.92 ; 
      RECT 40.576 156.546 40.68 160.92 ; 
      RECT 40.144 156.546 40.248 160.92 ; 
      RECT 39.712 156.546 39.816 160.92 ; 
      RECT 39.28 156.546 39.384 160.92 ; 
      RECT 38.848 156.546 38.952 160.92 ; 
      RECT 38.416 156.546 38.52 160.92 ; 
      RECT 37.984 156.546 38.088 160.92 ; 
      RECT 37.552 156.546 37.656 160.92 ; 
      RECT 36.7 156.546 37.008 160.92 ; 
      RECT 29.128 156.546 29.436 160.92 ; 
      RECT 28.48 156.546 28.584 160.92 ; 
      RECT 28.048 156.546 28.152 160.92 ; 
      RECT 27.616 156.546 27.72 160.92 ; 
      RECT 27.184 156.546 27.288 160.92 ; 
      RECT 26.752 156.546 26.856 160.92 ; 
      RECT 26.32 156.546 26.424 160.92 ; 
      RECT 25.888 156.546 25.992 160.92 ; 
      RECT 25.456 156.546 25.56 160.92 ; 
      RECT 25.024 156.546 25.128 160.92 ; 
      RECT 24.592 156.546 24.696 160.92 ; 
      RECT 24.16 156.546 24.264 160.92 ; 
      RECT 23.728 156.546 23.832 160.92 ; 
      RECT 23.296 156.546 23.4 160.92 ; 
      RECT 22.864 156.546 22.968 160.92 ; 
      RECT 22.432 156.546 22.536 160.92 ; 
      RECT 22 156.546 22.104 160.92 ; 
      RECT 21.568 156.546 21.672 160.92 ; 
      RECT 21.136 156.546 21.24 160.92 ; 
      RECT 20.704 156.546 20.808 160.92 ; 
      RECT 20.272 156.546 20.376 160.92 ; 
      RECT 19.84 156.546 19.944 160.92 ; 
      RECT 19.408 156.546 19.512 160.92 ; 
      RECT 18.976 156.546 19.08 160.92 ; 
      RECT 18.544 156.546 18.648 160.92 ; 
      RECT 18.112 156.546 18.216 160.92 ; 
      RECT 17.68 156.546 17.784 160.92 ; 
      RECT 17.248 156.546 17.352 160.92 ; 
      RECT 16.816 156.546 16.92 160.92 ; 
      RECT 16.384 156.546 16.488 160.92 ; 
      RECT 15.952 156.546 16.056 160.92 ; 
      RECT 15.52 156.546 15.624 160.92 ; 
      RECT 15.088 156.546 15.192 160.92 ; 
      RECT 14.656 156.546 14.76 160.92 ; 
      RECT 14.224 156.546 14.328 160.92 ; 
      RECT 13.792 156.546 13.896 160.92 ; 
      RECT 13.36 156.546 13.464 160.92 ; 
      RECT 12.928 156.546 13.032 160.92 ; 
      RECT 12.496 156.546 12.6 160.92 ; 
      RECT 12.064 156.546 12.168 160.92 ; 
      RECT 11.632 156.546 11.736 160.92 ; 
      RECT 11.2 156.546 11.304 160.92 ; 
      RECT 10.768 156.546 10.872 160.92 ; 
      RECT 10.336 156.546 10.44 160.92 ; 
      RECT 9.904 156.546 10.008 160.92 ; 
      RECT 9.472 156.546 9.576 160.92 ; 
      RECT 9.04 156.546 9.144 160.92 ; 
      RECT 8.608 156.546 8.712 160.92 ; 
      RECT 8.176 156.546 8.28 160.92 ; 
      RECT 7.744 156.546 7.848 160.92 ; 
      RECT 7.312 156.546 7.416 160.92 ; 
      RECT 6.88 156.546 6.984 160.92 ; 
      RECT 6.448 156.546 6.552 160.92 ; 
      RECT 6.016 156.546 6.12 160.92 ; 
      RECT 5.584 156.546 5.688 160.92 ; 
      RECT 5.152 156.546 5.256 160.92 ; 
      RECT 4.72 156.546 4.824 160.92 ; 
      RECT 4.288 156.546 4.392 160.92 ; 
      RECT 3.856 156.546 3.96 160.92 ; 
      RECT 3.424 156.546 3.528 160.92 ; 
      RECT 2.992 156.546 3.096 160.92 ; 
      RECT 2.56 156.546 2.664 160.92 ; 
      RECT 2.128 156.546 2.232 160.92 ; 
      RECT 1.696 156.546 1.8 160.92 ; 
      RECT 1.264 156.546 1.368 160.92 ; 
      RECT 0.832 156.546 0.936 160.92 ; 
      RECT 0.02 156.546 0.36 160.92 ; 
      RECT 0 193.638 66.096 195.402 ; 
      RECT 65.756 160.788 66.096 195.402 ; 
      RECT 37.532 166.804 65.284 195.402 ; 
      RECT 43.364 160.788 65.284 195.402 ; 
      RECT 28.892 193.608 37.204 195.402 ; 
      RECT 31.988 193.482 37.204 195.402 ; 
      RECT 0.812 166.024 28.564 195.402 ; 
      RECT 27.38 160.788 28.564 195.402 ; 
      RECT 0 160.788 0.34 195.402 ; 
      RECT 28.892 167.236 31.372 195.402 ; 
      RECT 31.988 193.464 37.06 195.402 ; 
      RECT 34.58 166.408 37.06 195.402 ; 
      RECT 34.544 192.436 37.06 195.402 ; 
      RECT 33.896 192.436 34.144 195.402 ; 
      RECT 31.988 192.436 33.532 195.402 ; 
      RECT 37.532 175.96 65.34 193.376 ; 
      RECT 0.756 175.96 28.564 193.376 ; 
      RECT 37.476 175.96 65.34 193.358 ; 
      RECT 0.756 175.96 28.62 193.358 ; 
      RECT 28.836 175.96 31.372 193.354 ; 
      RECT 32.708 163.528 33.388 195.402 ; 
      RECT 33.14 160.788 33.388 195.402 ; 
      RECT 29.972 162.472 31.516 191.848 ; 
      RECT 28.836 191.668 31.572 191.816 ; 
      RECT 34.524 187.372 37.06 191.804 ; 
      RECT 32.652 190.612 33.388 191.516 ; 
      RECT 32.708 188.308 33.444 189.356 ; 
      RECT 28.836 187.516 31.572 189.356 ; 
      RECT 32.652 185.356 33.388 187.196 ; 
      RECT 34.524 177.22 37.06 186.548 ; 
      RECT 28.836 179.812 31.572 184.388 ; 
      RECT 32.708 178.732 33.444 183.956 ; 
      RECT 32.652 181.036 33.444 182.876 ; 
      RECT 32.652 168.076 33.388 180.716 ; 
      RECT 32.652 168.076 33.444 178.556 ; 
      RECT 28.836 177.652 31.572 178.556 ; 
      RECT 34.58 166.408 37.204 175.832 ; 
      RECT 34.524 165.916 36.988 173.06 ; 
      RECT 28.892 169.804 31.572 171.284 ; 
      RECT 32.708 166.996 33.444 167.756 ; 
      RECT 29.108 166.852 31.572 167.612 ; 
      RECT 32.652 166.42 33.388 166.964 ; 
      RECT 29.108 163.852 31.516 191.848 ; 
      RECT 32.708 165.916 33.444 166.82 ; 
      RECT 38.18 166.036 65.284 195.402 ; 
      RECT 42.5 166.024 65.284 195.402 ; 
      RECT 37.532 160.788 37.852 195.402 ; 
      RECT 28.892 163.528 29.644 166.784 ; 
      RECT 37.532 160.788 38.716 166.4 ; 
      RECT 37.532 165.256 42.172 166.4 ; 
      RECT 42.5 160.788 43.036 195.402 ; 
      RECT 23.924 164.5 27.052 195.402 ; 
      RECT 0.812 160.788 23.596 195.402 ; 
      RECT 34.58 163.852 36.988 195.402 ; 
      RECT 34.724 161.494 37.204 165.788 ; 
      RECT 37.532 165.256 43.036 165.632 ; 
      RECT 41.636 160.788 65.284 165.62 ; 
      RECT 26.516 160.788 28.564 165.62 ; 
      RECT 32.652 165.34 33.444 165.596 ; 
      RECT 32.652 164.836 33.388 165.596 ; 
      RECT 40.772 163.72 65.284 165.62 ; 
      RECT 37.532 163.852 40.444 166.4 ; 
      RECT 32.708 163.756 33.444 164.804 ; 
      RECT 0.812 163.72 26.188 165.62 ; 
      RECT 25.652 160.788 26.188 195.402 ; 
      RECT 39.908 160.788 41.308 164.276 ; 
      RECT 37.532 163.528 39.58 166.4 ; 
      RECT 39.044 160.788 39.58 195.402 ; 
      RECT 24.788 163.528 26.188 195.402 ; 
      RECT 0.812 160.788 24.46 165.62 ; 
      RECT 32.708 160.788 32.812 195.402 ; 
      RECT 29.252 160.788 29.644 195.402 ; 
      RECT 24.788 160.788 25.324 195.402 ; 
      RECT 39.044 160.788 41.308 163.328 ; 
      RECT 34.58 160.788 36.988 163.328 ; 
      RECT 29.252 160.788 31.372 163.328 ; 
      RECT 25.652 160.788 28.564 163.328 ; 
      RECT 39.044 160.788 65.284 163.316 ; 
      RECT 0.812 160.788 25.324 163.316 ; 
      RECT 34.524 162.676 37.204 163.292 ; 
      RECT 37.532 160.788 65.284 162.26 ; 
      RECT 32.708 160.788 33.388 162.26 ; 
      RECT 28.892 160.788 31.372 162.26 ; 
      RECT 0.812 160.788 28.564 162.26 ; 
      RECT 31.988 160.788 33.388 161.848 ; 
      RECT 34.544 160.788 36.988 161.448 ; 
      RECT 31.988 160.788 33.532 161.448 ; 
      RECT 39.06 160.682 39.132 195.402 ; 
      RECT 38.628 160.682 38.7 195.402 ; 
      RECT 27.396 160.732 27.468 195.402 ; 
      RECT 26.964 160.732 27.036 195.402 ; 
      RECT 26.532 160.732 26.604 195.402 ; 
      RECT 26.1 160.732 26.172 195.402 ; 
      RECT 25.668 160.682 25.74 195.402 ; 
      RECT 25.236 160.682 25.308 195.402 ; 
      RECT 24.804 160.732 24.876 195.402 ; 
      RECT 24.372 160.732 24.444 195.402 ; 
      RECT 23.94 160.732 24.012 195.402 ; 
      RECT 23.508 160.732 23.58 195.402 ; 
      RECT 33.896 160.788 34.144 161.448 ; 
        RECT 34.564 193.374 35.076 197.748 ; 
        RECT 34.508 196.036 35.076 197.326 ; 
        RECT 33.916 194.944 34.164 197.748 ; 
        RECT 33.86 196.182 34.164 196.796 ; 
        RECT 33.916 193.374 34.02 197.748 ; 
        RECT 33.916 193.858 34.076 194.816 ; 
        RECT 33.916 193.374 34.164 193.73 ; 
        RECT 32.728 195.176 33.552 197.748 ; 
        RECT 33.448 193.374 33.552 197.748 ; 
        RECT 32.728 196.284 33.608 197.316 ; 
        RECT 32.728 193.374 33.12 197.748 ; 
        RECT 31.06 193.374 31.392 197.748 ; 
        RECT 31.06 193.728 31.448 197.47 ; 
        RECT 65.776 193.374 66.116 197.748 ; 
        RECT 65.2 193.374 65.304 197.748 ; 
        RECT 64.768 193.374 64.872 197.748 ; 
        RECT 64.336 193.374 64.44 197.748 ; 
        RECT 63.904 193.374 64.008 197.748 ; 
        RECT 63.472 193.374 63.576 197.748 ; 
        RECT 63.04 193.374 63.144 197.748 ; 
        RECT 62.608 193.374 62.712 197.748 ; 
        RECT 62.176 193.374 62.28 197.748 ; 
        RECT 61.744 193.374 61.848 197.748 ; 
        RECT 61.312 193.374 61.416 197.748 ; 
        RECT 60.88 193.374 60.984 197.748 ; 
        RECT 60.448 193.374 60.552 197.748 ; 
        RECT 60.016 193.374 60.12 197.748 ; 
        RECT 59.584 193.374 59.688 197.748 ; 
        RECT 59.152 193.374 59.256 197.748 ; 
        RECT 58.72 193.374 58.824 197.748 ; 
        RECT 58.288 193.374 58.392 197.748 ; 
        RECT 57.856 193.374 57.96 197.748 ; 
        RECT 57.424 193.374 57.528 197.748 ; 
        RECT 56.992 193.374 57.096 197.748 ; 
        RECT 56.56 193.374 56.664 197.748 ; 
        RECT 56.128 193.374 56.232 197.748 ; 
        RECT 55.696 193.374 55.8 197.748 ; 
        RECT 55.264 193.374 55.368 197.748 ; 
        RECT 54.832 193.374 54.936 197.748 ; 
        RECT 54.4 193.374 54.504 197.748 ; 
        RECT 53.968 193.374 54.072 197.748 ; 
        RECT 53.536 193.374 53.64 197.748 ; 
        RECT 53.104 193.374 53.208 197.748 ; 
        RECT 52.672 193.374 52.776 197.748 ; 
        RECT 52.24 193.374 52.344 197.748 ; 
        RECT 51.808 193.374 51.912 197.748 ; 
        RECT 51.376 193.374 51.48 197.748 ; 
        RECT 50.944 193.374 51.048 197.748 ; 
        RECT 50.512 193.374 50.616 197.748 ; 
        RECT 50.08 193.374 50.184 197.748 ; 
        RECT 49.648 193.374 49.752 197.748 ; 
        RECT 49.216 193.374 49.32 197.748 ; 
        RECT 48.784 193.374 48.888 197.748 ; 
        RECT 48.352 193.374 48.456 197.748 ; 
        RECT 47.92 193.374 48.024 197.748 ; 
        RECT 47.488 193.374 47.592 197.748 ; 
        RECT 47.056 193.374 47.16 197.748 ; 
        RECT 46.624 193.374 46.728 197.748 ; 
        RECT 46.192 193.374 46.296 197.748 ; 
        RECT 45.76 193.374 45.864 197.748 ; 
        RECT 45.328 193.374 45.432 197.748 ; 
        RECT 44.896 193.374 45 197.748 ; 
        RECT 44.464 193.374 44.568 197.748 ; 
        RECT 44.032 193.374 44.136 197.748 ; 
        RECT 43.6 193.374 43.704 197.748 ; 
        RECT 43.168 193.374 43.272 197.748 ; 
        RECT 42.736 193.374 42.84 197.748 ; 
        RECT 42.304 193.374 42.408 197.748 ; 
        RECT 41.872 193.374 41.976 197.748 ; 
        RECT 41.44 193.374 41.544 197.748 ; 
        RECT 41.008 193.374 41.112 197.748 ; 
        RECT 40.576 193.374 40.68 197.748 ; 
        RECT 40.144 193.374 40.248 197.748 ; 
        RECT 39.712 193.374 39.816 197.748 ; 
        RECT 39.28 193.374 39.384 197.748 ; 
        RECT 38.848 193.374 38.952 197.748 ; 
        RECT 38.416 193.374 38.52 197.748 ; 
        RECT 37.984 193.374 38.088 197.748 ; 
        RECT 37.552 193.374 37.656 197.748 ; 
        RECT 36.7 193.374 37.008 197.748 ; 
        RECT 29.128 193.374 29.436 197.748 ; 
        RECT 28.48 193.374 28.584 197.748 ; 
        RECT 28.048 193.374 28.152 197.748 ; 
        RECT 27.616 193.374 27.72 197.748 ; 
        RECT 27.184 193.374 27.288 197.748 ; 
        RECT 26.752 193.374 26.856 197.748 ; 
        RECT 26.32 193.374 26.424 197.748 ; 
        RECT 25.888 193.374 25.992 197.748 ; 
        RECT 25.456 193.374 25.56 197.748 ; 
        RECT 25.024 193.374 25.128 197.748 ; 
        RECT 24.592 193.374 24.696 197.748 ; 
        RECT 24.16 193.374 24.264 197.748 ; 
        RECT 23.728 193.374 23.832 197.748 ; 
        RECT 23.296 193.374 23.4 197.748 ; 
        RECT 22.864 193.374 22.968 197.748 ; 
        RECT 22.432 193.374 22.536 197.748 ; 
        RECT 22 193.374 22.104 197.748 ; 
        RECT 21.568 193.374 21.672 197.748 ; 
        RECT 21.136 193.374 21.24 197.748 ; 
        RECT 20.704 193.374 20.808 197.748 ; 
        RECT 20.272 193.374 20.376 197.748 ; 
        RECT 19.84 193.374 19.944 197.748 ; 
        RECT 19.408 193.374 19.512 197.748 ; 
        RECT 18.976 193.374 19.08 197.748 ; 
        RECT 18.544 193.374 18.648 197.748 ; 
        RECT 18.112 193.374 18.216 197.748 ; 
        RECT 17.68 193.374 17.784 197.748 ; 
        RECT 17.248 193.374 17.352 197.748 ; 
        RECT 16.816 193.374 16.92 197.748 ; 
        RECT 16.384 193.374 16.488 197.748 ; 
        RECT 15.952 193.374 16.056 197.748 ; 
        RECT 15.52 193.374 15.624 197.748 ; 
        RECT 15.088 193.374 15.192 197.748 ; 
        RECT 14.656 193.374 14.76 197.748 ; 
        RECT 14.224 193.374 14.328 197.748 ; 
        RECT 13.792 193.374 13.896 197.748 ; 
        RECT 13.36 193.374 13.464 197.748 ; 
        RECT 12.928 193.374 13.032 197.748 ; 
        RECT 12.496 193.374 12.6 197.748 ; 
        RECT 12.064 193.374 12.168 197.748 ; 
        RECT 11.632 193.374 11.736 197.748 ; 
        RECT 11.2 193.374 11.304 197.748 ; 
        RECT 10.768 193.374 10.872 197.748 ; 
        RECT 10.336 193.374 10.44 197.748 ; 
        RECT 9.904 193.374 10.008 197.748 ; 
        RECT 9.472 193.374 9.576 197.748 ; 
        RECT 9.04 193.374 9.144 197.748 ; 
        RECT 8.608 193.374 8.712 197.748 ; 
        RECT 8.176 193.374 8.28 197.748 ; 
        RECT 7.744 193.374 7.848 197.748 ; 
        RECT 7.312 193.374 7.416 197.748 ; 
        RECT 6.88 193.374 6.984 197.748 ; 
        RECT 6.448 193.374 6.552 197.748 ; 
        RECT 6.016 193.374 6.12 197.748 ; 
        RECT 5.584 193.374 5.688 197.748 ; 
        RECT 5.152 193.374 5.256 197.748 ; 
        RECT 4.72 193.374 4.824 197.748 ; 
        RECT 4.288 193.374 4.392 197.748 ; 
        RECT 3.856 193.374 3.96 197.748 ; 
        RECT 3.424 193.374 3.528 197.748 ; 
        RECT 2.992 193.374 3.096 197.748 ; 
        RECT 2.56 193.374 2.664 197.748 ; 
        RECT 2.128 193.374 2.232 197.748 ; 
        RECT 1.696 193.374 1.8 197.748 ; 
        RECT 1.264 193.374 1.368 197.748 ; 
        RECT 0.832 193.374 0.936 197.748 ; 
        RECT 0.02 193.374 0.36 197.748 ; 
        RECT 34.564 197.694 35.076 202.068 ; 
        RECT 34.508 200.356 35.076 201.646 ; 
        RECT 33.916 199.264 34.164 202.068 ; 
        RECT 33.86 200.502 34.164 201.116 ; 
        RECT 33.916 197.694 34.02 202.068 ; 
        RECT 33.916 198.178 34.076 199.136 ; 
        RECT 33.916 197.694 34.164 198.05 ; 
        RECT 32.728 199.496 33.552 202.068 ; 
        RECT 33.448 197.694 33.552 202.068 ; 
        RECT 32.728 200.604 33.608 201.636 ; 
        RECT 32.728 197.694 33.12 202.068 ; 
        RECT 31.06 197.694 31.392 202.068 ; 
        RECT 31.06 198.048 31.448 201.79 ; 
        RECT 65.776 197.694 66.116 202.068 ; 
        RECT 65.2 197.694 65.304 202.068 ; 
        RECT 64.768 197.694 64.872 202.068 ; 
        RECT 64.336 197.694 64.44 202.068 ; 
        RECT 63.904 197.694 64.008 202.068 ; 
        RECT 63.472 197.694 63.576 202.068 ; 
        RECT 63.04 197.694 63.144 202.068 ; 
        RECT 62.608 197.694 62.712 202.068 ; 
        RECT 62.176 197.694 62.28 202.068 ; 
        RECT 61.744 197.694 61.848 202.068 ; 
        RECT 61.312 197.694 61.416 202.068 ; 
        RECT 60.88 197.694 60.984 202.068 ; 
        RECT 60.448 197.694 60.552 202.068 ; 
        RECT 60.016 197.694 60.12 202.068 ; 
        RECT 59.584 197.694 59.688 202.068 ; 
        RECT 59.152 197.694 59.256 202.068 ; 
        RECT 58.72 197.694 58.824 202.068 ; 
        RECT 58.288 197.694 58.392 202.068 ; 
        RECT 57.856 197.694 57.96 202.068 ; 
        RECT 57.424 197.694 57.528 202.068 ; 
        RECT 56.992 197.694 57.096 202.068 ; 
        RECT 56.56 197.694 56.664 202.068 ; 
        RECT 56.128 197.694 56.232 202.068 ; 
        RECT 55.696 197.694 55.8 202.068 ; 
        RECT 55.264 197.694 55.368 202.068 ; 
        RECT 54.832 197.694 54.936 202.068 ; 
        RECT 54.4 197.694 54.504 202.068 ; 
        RECT 53.968 197.694 54.072 202.068 ; 
        RECT 53.536 197.694 53.64 202.068 ; 
        RECT 53.104 197.694 53.208 202.068 ; 
        RECT 52.672 197.694 52.776 202.068 ; 
        RECT 52.24 197.694 52.344 202.068 ; 
        RECT 51.808 197.694 51.912 202.068 ; 
        RECT 51.376 197.694 51.48 202.068 ; 
        RECT 50.944 197.694 51.048 202.068 ; 
        RECT 50.512 197.694 50.616 202.068 ; 
        RECT 50.08 197.694 50.184 202.068 ; 
        RECT 49.648 197.694 49.752 202.068 ; 
        RECT 49.216 197.694 49.32 202.068 ; 
        RECT 48.784 197.694 48.888 202.068 ; 
        RECT 48.352 197.694 48.456 202.068 ; 
        RECT 47.92 197.694 48.024 202.068 ; 
        RECT 47.488 197.694 47.592 202.068 ; 
        RECT 47.056 197.694 47.16 202.068 ; 
        RECT 46.624 197.694 46.728 202.068 ; 
        RECT 46.192 197.694 46.296 202.068 ; 
        RECT 45.76 197.694 45.864 202.068 ; 
        RECT 45.328 197.694 45.432 202.068 ; 
        RECT 44.896 197.694 45 202.068 ; 
        RECT 44.464 197.694 44.568 202.068 ; 
        RECT 44.032 197.694 44.136 202.068 ; 
        RECT 43.6 197.694 43.704 202.068 ; 
        RECT 43.168 197.694 43.272 202.068 ; 
        RECT 42.736 197.694 42.84 202.068 ; 
        RECT 42.304 197.694 42.408 202.068 ; 
        RECT 41.872 197.694 41.976 202.068 ; 
        RECT 41.44 197.694 41.544 202.068 ; 
        RECT 41.008 197.694 41.112 202.068 ; 
        RECT 40.576 197.694 40.68 202.068 ; 
        RECT 40.144 197.694 40.248 202.068 ; 
        RECT 39.712 197.694 39.816 202.068 ; 
        RECT 39.28 197.694 39.384 202.068 ; 
        RECT 38.848 197.694 38.952 202.068 ; 
        RECT 38.416 197.694 38.52 202.068 ; 
        RECT 37.984 197.694 38.088 202.068 ; 
        RECT 37.552 197.694 37.656 202.068 ; 
        RECT 36.7 197.694 37.008 202.068 ; 
        RECT 29.128 197.694 29.436 202.068 ; 
        RECT 28.48 197.694 28.584 202.068 ; 
        RECT 28.048 197.694 28.152 202.068 ; 
        RECT 27.616 197.694 27.72 202.068 ; 
        RECT 27.184 197.694 27.288 202.068 ; 
        RECT 26.752 197.694 26.856 202.068 ; 
        RECT 26.32 197.694 26.424 202.068 ; 
        RECT 25.888 197.694 25.992 202.068 ; 
        RECT 25.456 197.694 25.56 202.068 ; 
        RECT 25.024 197.694 25.128 202.068 ; 
        RECT 24.592 197.694 24.696 202.068 ; 
        RECT 24.16 197.694 24.264 202.068 ; 
        RECT 23.728 197.694 23.832 202.068 ; 
        RECT 23.296 197.694 23.4 202.068 ; 
        RECT 22.864 197.694 22.968 202.068 ; 
        RECT 22.432 197.694 22.536 202.068 ; 
        RECT 22 197.694 22.104 202.068 ; 
        RECT 21.568 197.694 21.672 202.068 ; 
        RECT 21.136 197.694 21.24 202.068 ; 
        RECT 20.704 197.694 20.808 202.068 ; 
        RECT 20.272 197.694 20.376 202.068 ; 
        RECT 19.84 197.694 19.944 202.068 ; 
        RECT 19.408 197.694 19.512 202.068 ; 
        RECT 18.976 197.694 19.08 202.068 ; 
        RECT 18.544 197.694 18.648 202.068 ; 
        RECT 18.112 197.694 18.216 202.068 ; 
        RECT 17.68 197.694 17.784 202.068 ; 
        RECT 17.248 197.694 17.352 202.068 ; 
        RECT 16.816 197.694 16.92 202.068 ; 
        RECT 16.384 197.694 16.488 202.068 ; 
        RECT 15.952 197.694 16.056 202.068 ; 
        RECT 15.52 197.694 15.624 202.068 ; 
        RECT 15.088 197.694 15.192 202.068 ; 
        RECT 14.656 197.694 14.76 202.068 ; 
        RECT 14.224 197.694 14.328 202.068 ; 
        RECT 13.792 197.694 13.896 202.068 ; 
        RECT 13.36 197.694 13.464 202.068 ; 
        RECT 12.928 197.694 13.032 202.068 ; 
        RECT 12.496 197.694 12.6 202.068 ; 
        RECT 12.064 197.694 12.168 202.068 ; 
        RECT 11.632 197.694 11.736 202.068 ; 
        RECT 11.2 197.694 11.304 202.068 ; 
        RECT 10.768 197.694 10.872 202.068 ; 
        RECT 10.336 197.694 10.44 202.068 ; 
        RECT 9.904 197.694 10.008 202.068 ; 
        RECT 9.472 197.694 9.576 202.068 ; 
        RECT 9.04 197.694 9.144 202.068 ; 
        RECT 8.608 197.694 8.712 202.068 ; 
        RECT 8.176 197.694 8.28 202.068 ; 
        RECT 7.744 197.694 7.848 202.068 ; 
        RECT 7.312 197.694 7.416 202.068 ; 
        RECT 6.88 197.694 6.984 202.068 ; 
        RECT 6.448 197.694 6.552 202.068 ; 
        RECT 6.016 197.694 6.12 202.068 ; 
        RECT 5.584 197.694 5.688 202.068 ; 
        RECT 5.152 197.694 5.256 202.068 ; 
        RECT 4.72 197.694 4.824 202.068 ; 
        RECT 4.288 197.694 4.392 202.068 ; 
        RECT 3.856 197.694 3.96 202.068 ; 
        RECT 3.424 197.694 3.528 202.068 ; 
        RECT 2.992 197.694 3.096 202.068 ; 
        RECT 2.56 197.694 2.664 202.068 ; 
        RECT 2.128 197.694 2.232 202.068 ; 
        RECT 1.696 197.694 1.8 202.068 ; 
        RECT 1.264 197.694 1.368 202.068 ; 
        RECT 0.832 197.694 0.936 202.068 ; 
        RECT 0.02 197.694 0.36 202.068 ; 
        RECT 34.564 202.014 35.076 206.388 ; 
        RECT 34.508 204.676 35.076 205.966 ; 
        RECT 33.916 203.584 34.164 206.388 ; 
        RECT 33.86 204.822 34.164 205.436 ; 
        RECT 33.916 202.014 34.02 206.388 ; 
        RECT 33.916 202.498 34.076 203.456 ; 
        RECT 33.916 202.014 34.164 202.37 ; 
        RECT 32.728 203.816 33.552 206.388 ; 
        RECT 33.448 202.014 33.552 206.388 ; 
        RECT 32.728 204.924 33.608 205.956 ; 
        RECT 32.728 202.014 33.12 206.388 ; 
        RECT 31.06 202.014 31.392 206.388 ; 
        RECT 31.06 202.368 31.448 206.11 ; 
        RECT 65.776 202.014 66.116 206.388 ; 
        RECT 65.2 202.014 65.304 206.388 ; 
        RECT 64.768 202.014 64.872 206.388 ; 
        RECT 64.336 202.014 64.44 206.388 ; 
        RECT 63.904 202.014 64.008 206.388 ; 
        RECT 63.472 202.014 63.576 206.388 ; 
        RECT 63.04 202.014 63.144 206.388 ; 
        RECT 62.608 202.014 62.712 206.388 ; 
        RECT 62.176 202.014 62.28 206.388 ; 
        RECT 61.744 202.014 61.848 206.388 ; 
        RECT 61.312 202.014 61.416 206.388 ; 
        RECT 60.88 202.014 60.984 206.388 ; 
        RECT 60.448 202.014 60.552 206.388 ; 
        RECT 60.016 202.014 60.12 206.388 ; 
        RECT 59.584 202.014 59.688 206.388 ; 
        RECT 59.152 202.014 59.256 206.388 ; 
        RECT 58.72 202.014 58.824 206.388 ; 
        RECT 58.288 202.014 58.392 206.388 ; 
        RECT 57.856 202.014 57.96 206.388 ; 
        RECT 57.424 202.014 57.528 206.388 ; 
        RECT 56.992 202.014 57.096 206.388 ; 
        RECT 56.56 202.014 56.664 206.388 ; 
        RECT 56.128 202.014 56.232 206.388 ; 
        RECT 55.696 202.014 55.8 206.388 ; 
        RECT 55.264 202.014 55.368 206.388 ; 
        RECT 54.832 202.014 54.936 206.388 ; 
        RECT 54.4 202.014 54.504 206.388 ; 
        RECT 53.968 202.014 54.072 206.388 ; 
        RECT 53.536 202.014 53.64 206.388 ; 
        RECT 53.104 202.014 53.208 206.388 ; 
        RECT 52.672 202.014 52.776 206.388 ; 
        RECT 52.24 202.014 52.344 206.388 ; 
        RECT 51.808 202.014 51.912 206.388 ; 
        RECT 51.376 202.014 51.48 206.388 ; 
        RECT 50.944 202.014 51.048 206.388 ; 
        RECT 50.512 202.014 50.616 206.388 ; 
        RECT 50.08 202.014 50.184 206.388 ; 
        RECT 49.648 202.014 49.752 206.388 ; 
        RECT 49.216 202.014 49.32 206.388 ; 
        RECT 48.784 202.014 48.888 206.388 ; 
        RECT 48.352 202.014 48.456 206.388 ; 
        RECT 47.92 202.014 48.024 206.388 ; 
        RECT 47.488 202.014 47.592 206.388 ; 
        RECT 47.056 202.014 47.16 206.388 ; 
        RECT 46.624 202.014 46.728 206.388 ; 
        RECT 46.192 202.014 46.296 206.388 ; 
        RECT 45.76 202.014 45.864 206.388 ; 
        RECT 45.328 202.014 45.432 206.388 ; 
        RECT 44.896 202.014 45 206.388 ; 
        RECT 44.464 202.014 44.568 206.388 ; 
        RECT 44.032 202.014 44.136 206.388 ; 
        RECT 43.6 202.014 43.704 206.388 ; 
        RECT 43.168 202.014 43.272 206.388 ; 
        RECT 42.736 202.014 42.84 206.388 ; 
        RECT 42.304 202.014 42.408 206.388 ; 
        RECT 41.872 202.014 41.976 206.388 ; 
        RECT 41.44 202.014 41.544 206.388 ; 
        RECT 41.008 202.014 41.112 206.388 ; 
        RECT 40.576 202.014 40.68 206.388 ; 
        RECT 40.144 202.014 40.248 206.388 ; 
        RECT 39.712 202.014 39.816 206.388 ; 
        RECT 39.28 202.014 39.384 206.388 ; 
        RECT 38.848 202.014 38.952 206.388 ; 
        RECT 38.416 202.014 38.52 206.388 ; 
        RECT 37.984 202.014 38.088 206.388 ; 
        RECT 37.552 202.014 37.656 206.388 ; 
        RECT 36.7 202.014 37.008 206.388 ; 
        RECT 29.128 202.014 29.436 206.388 ; 
        RECT 28.48 202.014 28.584 206.388 ; 
        RECT 28.048 202.014 28.152 206.388 ; 
        RECT 27.616 202.014 27.72 206.388 ; 
        RECT 27.184 202.014 27.288 206.388 ; 
        RECT 26.752 202.014 26.856 206.388 ; 
        RECT 26.32 202.014 26.424 206.388 ; 
        RECT 25.888 202.014 25.992 206.388 ; 
        RECT 25.456 202.014 25.56 206.388 ; 
        RECT 25.024 202.014 25.128 206.388 ; 
        RECT 24.592 202.014 24.696 206.388 ; 
        RECT 24.16 202.014 24.264 206.388 ; 
        RECT 23.728 202.014 23.832 206.388 ; 
        RECT 23.296 202.014 23.4 206.388 ; 
        RECT 22.864 202.014 22.968 206.388 ; 
        RECT 22.432 202.014 22.536 206.388 ; 
        RECT 22 202.014 22.104 206.388 ; 
        RECT 21.568 202.014 21.672 206.388 ; 
        RECT 21.136 202.014 21.24 206.388 ; 
        RECT 20.704 202.014 20.808 206.388 ; 
        RECT 20.272 202.014 20.376 206.388 ; 
        RECT 19.84 202.014 19.944 206.388 ; 
        RECT 19.408 202.014 19.512 206.388 ; 
        RECT 18.976 202.014 19.08 206.388 ; 
        RECT 18.544 202.014 18.648 206.388 ; 
        RECT 18.112 202.014 18.216 206.388 ; 
        RECT 17.68 202.014 17.784 206.388 ; 
        RECT 17.248 202.014 17.352 206.388 ; 
        RECT 16.816 202.014 16.92 206.388 ; 
        RECT 16.384 202.014 16.488 206.388 ; 
        RECT 15.952 202.014 16.056 206.388 ; 
        RECT 15.52 202.014 15.624 206.388 ; 
        RECT 15.088 202.014 15.192 206.388 ; 
        RECT 14.656 202.014 14.76 206.388 ; 
        RECT 14.224 202.014 14.328 206.388 ; 
        RECT 13.792 202.014 13.896 206.388 ; 
        RECT 13.36 202.014 13.464 206.388 ; 
        RECT 12.928 202.014 13.032 206.388 ; 
        RECT 12.496 202.014 12.6 206.388 ; 
        RECT 12.064 202.014 12.168 206.388 ; 
        RECT 11.632 202.014 11.736 206.388 ; 
        RECT 11.2 202.014 11.304 206.388 ; 
        RECT 10.768 202.014 10.872 206.388 ; 
        RECT 10.336 202.014 10.44 206.388 ; 
        RECT 9.904 202.014 10.008 206.388 ; 
        RECT 9.472 202.014 9.576 206.388 ; 
        RECT 9.04 202.014 9.144 206.388 ; 
        RECT 8.608 202.014 8.712 206.388 ; 
        RECT 8.176 202.014 8.28 206.388 ; 
        RECT 7.744 202.014 7.848 206.388 ; 
        RECT 7.312 202.014 7.416 206.388 ; 
        RECT 6.88 202.014 6.984 206.388 ; 
        RECT 6.448 202.014 6.552 206.388 ; 
        RECT 6.016 202.014 6.12 206.388 ; 
        RECT 5.584 202.014 5.688 206.388 ; 
        RECT 5.152 202.014 5.256 206.388 ; 
        RECT 4.72 202.014 4.824 206.388 ; 
        RECT 4.288 202.014 4.392 206.388 ; 
        RECT 3.856 202.014 3.96 206.388 ; 
        RECT 3.424 202.014 3.528 206.388 ; 
        RECT 2.992 202.014 3.096 206.388 ; 
        RECT 2.56 202.014 2.664 206.388 ; 
        RECT 2.128 202.014 2.232 206.388 ; 
        RECT 1.696 202.014 1.8 206.388 ; 
        RECT 1.264 202.014 1.368 206.388 ; 
        RECT 0.832 202.014 0.936 206.388 ; 
        RECT 0.02 202.014 0.36 206.388 ; 
        RECT 34.564 206.334 35.076 210.708 ; 
        RECT 34.508 208.996 35.076 210.286 ; 
        RECT 33.916 207.904 34.164 210.708 ; 
        RECT 33.86 209.142 34.164 209.756 ; 
        RECT 33.916 206.334 34.02 210.708 ; 
        RECT 33.916 206.818 34.076 207.776 ; 
        RECT 33.916 206.334 34.164 206.69 ; 
        RECT 32.728 208.136 33.552 210.708 ; 
        RECT 33.448 206.334 33.552 210.708 ; 
        RECT 32.728 209.244 33.608 210.276 ; 
        RECT 32.728 206.334 33.12 210.708 ; 
        RECT 31.06 206.334 31.392 210.708 ; 
        RECT 31.06 206.688 31.448 210.43 ; 
        RECT 65.776 206.334 66.116 210.708 ; 
        RECT 65.2 206.334 65.304 210.708 ; 
        RECT 64.768 206.334 64.872 210.708 ; 
        RECT 64.336 206.334 64.44 210.708 ; 
        RECT 63.904 206.334 64.008 210.708 ; 
        RECT 63.472 206.334 63.576 210.708 ; 
        RECT 63.04 206.334 63.144 210.708 ; 
        RECT 62.608 206.334 62.712 210.708 ; 
        RECT 62.176 206.334 62.28 210.708 ; 
        RECT 61.744 206.334 61.848 210.708 ; 
        RECT 61.312 206.334 61.416 210.708 ; 
        RECT 60.88 206.334 60.984 210.708 ; 
        RECT 60.448 206.334 60.552 210.708 ; 
        RECT 60.016 206.334 60.12 210.708 ; 
        RECT 59.584 206.334 59.688 210.708 ; 
        RECT 59.152 206.334 59.256 210.708 ; 
        RECT 58.72 206.334 58.824 210.708 ; 
        RECT 58.288 206.334 58.392 210.708 ; 
        RECT 57.856 206.334 57.96 210.708 ; 
        RECT 57.424 206.334 57.528 210.708 ; 
        RECT 56.992 206.334 57.096 210.708 ; 
        RECT 56.56 206.334 56.664 210.708 ; 
        RECT 56.128 206.334 56.232 210.708 ; 
        RECT 55.696 206.334 55.8 210.708 ; 
        RECT 55.264 206.334 55.368 210.708 ; 
        RECT 54.832 206.334 54.936 210.708 ; 
        RECT 54.4 206.334 54.504 210.708 ; 
        RECT 53.968 206.334 54.072 210.708 ; 
        RECT 53.536 206.334 53.64 210.708 ; 
        RECT 53.104 206.334 53.208 210.708 ; 
        RECT 52.672 206.334 52.776 210.708 ; 
        RECT 52.24 206.334 52.344 210.708 ; 
        RECT 51.808 206.334 51.912 210.708 ; 
        RECT 51.376 206.334 51.48 210.708 ; 
        RECT 50.944 206.334 51.048 210.708 ; 
        RECT 50.512 206.334 50.616 210.708 ; 
        RECT 50.08 206.334 50.184 210.708 ; 
        RECT 49.648 206.334 49.752 210.708 ; 
        RECT 49.216 206.334 49.32 210.708 ; 
        RECT 48.784 206.334 48.888 210.708 ; 
        RECT 48.352 206.334 48.456 210.708 ; 
        RECT 47.92 206.334 48.024 210.708 ; 
        RECT 47.488 206.334 47.592 210.708 ; 
        RECT 47.056 206.334 47.16 210.708 ; 
        RECT 46.624 206.334 46.728 210.708 ; 
        RECT 46.192 206.334 46.296 210.708 ; 
        RECT 45.76 206.334 45.864 210.708 ; 
        RECT 45.328 206.334 45.432 210.708 ; 
        RECT 44.896 206.334 45 210.708 ; 
        RECT 44.464 206.334 44.568 210.708 ; 
        RECT 44.032 206.334 44.136 210.708 ; 
        RECT 43.6 206.334 43.704 210.708 ; 
        RECT 43.168 206.334 43.272 210.708 ; 
        RECT 42.736 206.334 42.84 210.708 ; 
        RECT 42.304 206.334 42.408 210.708 ; 
        RECT 41.872 206.334 41.976 210.708 ; 
        RECT 41.44 206.334 41.544 210.708 ; 
        RECT 41.008 206.334 41.112 210.708 ; 
        RECT 40.576 206.334 40.68 210.708 ; 
        RECT 40.144 206.334 40.248 210.708 ; 
        RECT 39.712 206.334 39.816 210.708 ; 
        RECT 39.28 206.334 39.384 210.708 ; 
        RECT 38.848 206.334 38.952 210.708 ; 
        RECT 38.416 206.334 38.52 210.708 ; 
        RECT 37.984 206.334 38.088 210.708 ; 
        RECT 37.552 206.334 37.656 210.708 ; 
        RECT 36.7 206.334 37.008 210.708 ; 
        RECT 29.128 206.334 29.436 210.708 ; 
        RECT 28.48 206.334 28.584 210.708 ; 
        RECT 28.048 206.334 28.152 210.708 ; 
        RECT 27.616 206.334 27.72 210.708 ; 
        RECT 27.184 206.334 27.288 210.708 ; 
        RECT 26.752 206.334 26.856 210.708 ; 
        RECT 26.32 206.334 26.424 210.708 ; 
        RECT 25.888 206.334 25.992 210.708 ; 
        RECT 25.456 206.334 25.56 210.708 ; 
        RECT 25.024 206.334 25.128 210.708 ; 
        RECT 24.592 206.334 24.696 210.708 ; 
        RECT 24.16 206.334 24.264 210.708 ; 
        RECT 23.728 206.334 23.832 210.708 ; 
        RECT 23.296 206.334 23.4 210.708 ; 
        RECT 22.864 206.334 22.968 210.708 ; 
        RECT 22.432 206.334 22.536 210.708 ; 
        RECT 22 206.334 22.104 210.708 ; 
        RECT 21.568 206.334 21.672 210.708 ; 
        RECT 21.136 206.334 21.24 210.708 ; 
        RECT 20.704 206.334 20.808 210.708 ; 
        RECT 20.272 206.334 20.376 210.708 ; 
        RECT 19.84 206.334 19.944 210.708 ; 
        RECT 19.408 206.334 19.512 210.708 ; 
        RECT 18.976 206.334 19.08 210.708 ; 
        RECT 18.544 206.334 18.648 210.708 ; 
        RECT 18.112 206.334 18.216 210.708 ; 
        RECT 17.68 206.334 17.784 210.708 ; 
        RECT 17.248 206.334 17.352 210.708 ; 
        RECT 16.816 206.334 16.92 210.708 ; 
        RECT 16.384 206.334 16.488 210.708 ; 
        RECT 15.952 206.334 16.056 210.708 ; 
        RECT 15.52 206.334 15.624 210.708 ; 
        RECT 15.088 206.334 15.192 210.708 ; 
        RECT 14.656 206.334 14.76 210.708 ; 
        RECT 14.224 206.334 14.328 210.708 ; 
        RECT 13.792 206.334 13.896 210.708 ; 
        RECT 13.36 206.334 13.464 210.708 ; 
        RECT 12.928 206.334 13.032 210.708 ; 
        RECT 12.496 206.334 12.6 210.708 ; 
        RECT 12.064 206.334 12.168 210.708 ; 
        RECT 11.632 206.334 11.736 210.708 ; 
        RECT 11.2 206.334 11.304 210.708 ; 
        RECT 10.768 206.334 10.872 210.708 ; 
        RECT 10.336 206.334 10.44 210.708 ; 
        RECT 9.904 206.334 10.008 210.708 ; 
        RECT 9.472 206.334 9.576 210.708 ; 
        RECT 9.04 206.334 9.144 210.708 ; 
        RECT 8.608 206.334 8.712 210.708 ; 
        RECT 8.176 206.334 8.28 210.708 ; 
        RECT 7.744 206.334 7.848 210.708 ; 
        RECT 7.312 206.334 7.416 210.708 ; 
        RECT 6.88 206.334 6.984 210.708 ; 
        RECT 6.448 206.334 6.552 210.708 ; 
        RECT 6.016 206.334 6.12 210.708 ; 
        RECT 5.584 206.334 5.688 210.708 ; 
        RECT 5.152 206.334 5.256 210.708 ; 
        RECT 4.72 206.334 4.824 210.708 ; 
        RECT 4.288 206.334 4.392 210.708 ; 
        RECT 3.856 206.334 3.96 210.708 ; 
        RECT 3.424 206.334 3.528 210.708 ; 
        RECT 2.992 206.334 3.096 210.708 ; 
        RECT 2.56 206.334 2.664 210.708 ; 
        RECT 2.128 206.334 2.232 210.708 ; 
        RECT 1.696 206.334 1.8 210.708 ; 
        RECT 1.264 206.334 1.368 210.708 ; 
        RECT 0.832 206.334 0.936 210.708 ; 
        RECT 0.02 206.334 0.36 210.708 ; 
        RECT 34.564 210.654 35.076 215.028 ; 
        RECT 34.508 213.316 35.076 214.606 ; 
        RECT 33.916 212.224 34.164 215.028 ; 
        RECT 33.86 213.462 34.164 214.076 ; 
        RECT 33.916 210.654 34.02 215.028 ; 
        RECT 33.916 211.138 34.076 212.096 ; 
        RECT 33.916 210.654 34.164 211.01 ; 
        RECT 32.728 212.456 33.552 215.028 ; 
        RECT 33.448 210.654 33.552 215.028 ; 
        RECT 32.728 213.564 33.608 214.596 ; 
        RECT 32.728 210.654 33.12 215.028 ; 
        RECT 31.06 210.654 31.392 215.028 ; 
        RECT 31.06 211.008 31.448 214.75 ; 
        RECT 65.776 210.654 66.116 215.028 ; 
        RECT 65.2 210.654 65.304 215.028 ; 
        RECT 64.768 210.654 64.872 215.028 ; 
        RECT 64.336 210.654 64.44 215.028 ; 
        RECT 63.904 210.654 64.008 215.028 ; 
        RECT 63.472 210.654 63.576 215.028 ; 
        RECT 63.04 210.654 63.144 215.028 ; 
        RECT 62.608 210.654 62.712 215.028 ; 
        RECT 62.176 210.654 62.28 215.028 ; 
        RECT 61.744 210.654 61.848 215.028 ; 
        RECT 61.312 210.654 61.416 215.028 ; 
        RECT 60.88 210.654 60.984 215.028 ; 
        RECT 60.448 210.654 60.552 215.028 ; 
        RECT 60.016 210.654 60.12 215.028 ; 
        RECT 59.584 210.654 59.688 215.028 ; 
        RECT 59.152 210.654 59.256 215.028 ; 
        RECT 58.72 210.654 58.824 215.028 ; 
        RECT 58.288 210.654 58.392 215.028 ; 
        RECT 57.856 210.654 57.96 215.028 ; 
        RECT 57.424 210.654 57.528 215.028 ; 
        RECT 56.992 210.654 57.096 215.028 ; 
        RECT 56.56 210.654 56.664 215.028 ; 
        RECT 56.128 210.654 56.232 215.028 ; 
        RECT 55.696 210.654 55.8 215.028 ; 
        RECT 55.264 210.654 55.368 215.028 ; 
        RECT 54.832 210.654 54.936 215.028 ; 
        RECT 54.4 210.654 54.504 215.028 ; 
        RECT 53.968 210.654 54.072 215.028 ; 
        RECT 53.536 210.654 53.64 215.028 ; 
        RECT 53.104 210.654 53.208 215.028 ; 
        RECT 52.672 210.654 52.776 215.028 ; 
        RECT 52.24 210.654 52.344 215.028 ; 
        RECT 51.808 210.654 51.912 215.028 ; 
        RECT 51.376 210.654 51.48 215.028 ; 
        RECT 50.944 210.654 51.048 215.028 ; 
        RECT 50.512 210.654 50.616 215.028 ; 
        RECT 50.08 210.654 50.184 215.028 ; 
        RECT 49.648 210.654 49.752 215.028 ; 
        RECT 49.216 210.654 49.32 215.028 ; 
        RECT 48.784 210.654 48.888 215.028 ; 
        RECT 48.352 210.654 48.456 215.028 ; 
        RECT 47.92 210.654 48.024 215.028 ; 
        RECT 47.488 210.654 47.592 215.028 ; 
        RECT 47.056 210.654 47.16 215.028 ; 
        RECT 46.624 210.654 46.728 215.028 ; 
        RECT 46.192 210.654 46.296 215.028 ; 
        RECT 45.76 210.654 45.864 215.028 ; 
        RECT 45.328 210.654 45.432 215.028 ; 
        RECT 44.896 210.654 45 215.028 ; 
        RECT 44.464 210.654 44.568 215.028 ; 
        RECT 44.032 210.654 44.136 215.028 ; 
        RECT 43.6 210.654 43.704 215.028 ; 
        RECT 43.168 210.654 43.272 215.028 ; 
        RECT 42.736 210.654 42.84 215.028 ; 
        RECT 42.304 210.654 42.408 215.028 ; 
        RECT 41.872 210.654 41.976 215.028 ; 
        RECT 41.44 210.654 41.544 215.028 ; 
        RECT 41.008 210.654 41.112 215.028 ; 
        RECT 40.576 210.654 40.68 215.028 ; 
        RECT 40.144 210.654 40.248 215.028 ; 
        RECT 39.712 210.654 39.816 215.028 ; 
        RECT 39.28 210.654 39.384 215.028 ; 
        RECT 38.848 210.654 38.952 215.028 ; 
        RECT 38.416 210.654 38.52 215.028 ; 
        RECT 37.984 210.654 38.088 215.028 ; 
        RECT 37.552 210.654 37.656 215.028 ; 
        RECT 36.7 210.654 37.008 215.028 ; 
        RECT 29.128 210.654 29.436 215.028 ; 
        RECT 28.48 210.654 28.584 215.028 ; 
        RECT 28.048 210.654 28.152 215.028 ; 
        RECT 27.616 210.654 27.72 215.028 ; 
        RECT 27.184 210.654 27.288 215.028 ; 
        RECT 26.752 210.654 26.856 215.028 ; 
        RECT 26.32 210.654 26.424 215.028 ; 
        RECT 25.888 210.654 25.992 215.028 ; 
        RECT 25.456 210.654 25.56 215.028 ; 
        RECT 25.024 210.654 25.128 215.028 ; 
        RECT 24.592 210.654 24.696 215.028 ; 
        RECT 24.16 210.654 24.264 215.028 ; 
        RECT 23.728 210.654 23.832 215.028 ; 
        RECT 23.296 210.654 23.4 215.028 ; 
        RECT 22.864 210.654 22.968 215.028 ; 
        RECT 22.432 210.654 22.536 215.028 ; 
        RECT 22 210.654 22.104 215.028 ; 
        RECT 21.568 210.654 21.672 215.028 ; 
        RECT 21.136 210.654 21.24 215.028 ; 
        RECT 20.704 210.654 20.808 215.028 ; 
        RECT 20.272 210.654 20.376 215.028 ; 
        RECT 19.84 210.654 19.944 215.028 ; 
        RECT 19.408 210.654 19.512 215.028 ; 
        RECT 18.976 210.654 19.08 215.028 ; 
        RECT 18.544 210.654 18.648 215.028 ; 
        RECT 18.112 210.654 18.216 215.028 ; 
        RECT 17.68 210.654 17.784 215.028 ; 
        RECT 17.248 210.654 17.352 215.028 ; 
        RECT 16.816 210.654 16.92 215.028 ; 
        RECT 16.384 210.654 16.488 215.028 ; 
        RECT 15.952 210.654 16.056 215.028 ; 
        RECT 15.52 210.654 15.624 215.028 ; 
        RECT 15.088 210.654 15.192 215.028 ; 
        RECT 14.656 210.654 14.76 215.028 ; 
        RECT 14.224 210.654 14.328 215.028 ; 
        RECT 13.792 210.654 13.896 215.028 ; 
        RECT 13.36 210.654 13.464 215.028 ; 
        RECT 12.928 210.654 13.032 215.028 ; 
        RECT 12.496 210.654 12.6 215.028 ; 
        RECT 12.064 210.654 12.168 215.028 ; 
        RECT 11.632 210.654 11.736 215.028 ; 
        RECT 11.2 210.654 11.304 215.028 ; 
        RECT 10.768 210.654 10.872 215.028 ; 
        RECT 10.336 210.654 10.44 215.028 ; 
        RECT 9.904 210.654 10.008 215.028 ; 
        RECT 9.472 210.654 9.576 215.028 ; 
        RECT 9.04 210.654 9.144 215.028 ; 
        RECT 8.608 210.654 8.712 215.028 ; 
        RECT 8.176 210.654 8.28 215.028 ; 
        RECT 7.744 210.654 7.848 215.028 ; 
        RECT 7.312 210.654 7.416 215.028 ; 
        RECT 6.88 210.654 6.984 215.028 ; 
        RECT 6.448 210.654 6.552 215.028 ; 
        RECT 6.016 210.654 6.12 215.028 ; 
        RECT 5.584 210.654 5.688 215.028 ; 
        RECT 5.152 210.654 5.256 215.028 ; 
        RECT 4.72 210.654 4.824 215.028 ; 
        RECT 4.288 210.654 4.392 215.028 ; 
        RECT 3.856 210.654 3.96 215.028 ; 
        RECT 3.424 210.654 3.528 215.028 ; 
        RECT 2.992 210.654 3.096 215.028 ; 
        RECT 2.56 210.654 2.664 215.028 ; 
        RECT 2.128 210.654 2.232 215.028 ; 
        RECT 1.696 210.654 1.8 215.028 ; 
        RECT 1.264 210.654 1.368 215.028 ; 
        RECT 0.832 210.654 0.936 215.028 ; 
        RECT 0.02 210.654 0.36 215.028 ; 
        RECT 34.564 214.974 35.076 219.348 ; 
        RECT 34.508 217.636 35.076 218.926 ; 
        RECT 33.916 216.544 34.164 219.348 ; 
        RECT 33.86 217.782 34.164 218.396 ; 
        RECT 33.916 214.974 34.02 219.348 ; 
        RECT 33.916 215.458 34.076 216.416 ; 
        RECT 33.916 214.974 34.164 215.33 ; 
        RECT 32.728 216.776 33.552 219.348 ; 
        RECT 33.448 214.974 33.552 219.348 ; 
        RECT 32.728 217.884 33.608 218.916 ; 
        RECT 32.728 214.974 33.12 219.348 ; 
        RECT 31.06 214.974 31.392 219.348 ; 
        RECT 31.06 215.328 31.448 219.07 ; 
        RECT 65.776 214.974 66.116 219.348 ; 
        RECT 65.2 214.974 65.304 219.348 ; 
        RECT 64.768 214.974 64.872 219.348 ; 
        RECT 64.336 214.974 64.44 219.348 ; 
        RECT 63.904 214.974 64.008 219.348 ; 
        RECT 63.472 214.974 63.576 219.348 ; 
        RECT 63.04 214.974 63.144 219.348 ; 
        RECT 62.608 214.974 62.712 219.348 ; 
        RECT 62.176 214.974 62.28 219.348 ; 
        RECT 61.744 214.974 61.848 219.348 ; 
        RECT 61.312 214.974 61.416 219.348 ; 
        RECT 60.88 214.974 60.984 219.348 ; 
        RECT 60.448 214.974 60.552 219.348 ; 
        RECT 60.016 214.974 60.12 219.348 ; 
        RECT 59.584 214.974 59.688 219.348 ; 
        RECT 59.152 214.974 59.256 219.348 ; 
        RECT 58.72 214.974 58.824 219.348 ; 
        RECT 58.288 214.974 58.392 219.348 ; 
        RECT 57.856 214.974 57.96 219.348 ; 
        RECT 57.424 214.974 57.528 219.348 ; 
        RECT 56.992 214.974 57.096 219.348 ; 
        RECT 56.56 214.974 56.664 219.348 ; 
        RECT 56.128 214.974 56.232 219.348 ; 
        RECT 55.696 214.974 55.8 219.348 ; 
        RECT 55.264 214.974 55.368 219.348 ; 
        RECT 54.832 214.974 54.936 219.348 ; 
        RECT 54.4 214.974 54.504 219.348 ; 
        RECT 53.968 214.974 54.072 219.348 ; 
        RECT 53.536 214.974 53.64 219.348 ; 
        RECT 53.104 214.974 53.208 219.348 ; 
        RECT 52.672 214.974 52.776 219.348 ; 
        RECT 52.24 214.974 52.344 219.348 ; 
        RECT 51.808 214.974 51.912 219.348 ; 
        RECT 51.376 214.974 51.48 219.348 ; 
        RECT 50.944 214.974 51.048 219.348 ; 
        RECT 50.512 214.974 50.616 219.348 ; 
        RECT 50.08 214.974 50.184 219.348 ; 
        RECT 49.648 214.974 49.752 219.348 ; 
        RECT 49.216 214.974 49.32 219.348 ; 
        RECT 48.784 214.974 48.888 219.348 ; 
        RECT 48.352 214.974 48.456 219.348 ; 
        RECT 47.92 214.974 48.024 219.348 ; 
        RECT 47.488 214.974 47.592 219.348 ; 
        RECT 47.056 214.974 47.16 219.348 ; 
        RECT 46.624 214.974 46.728 219.348 ; 
        RECT 46.192 214.974 46.296 219.348 ; 
        RECT 45.76 214.974 45.864 219.348 ; 
        RECT 45.328 214.974 45.432 219.348 ; 
        RECT 44.896 214.974 45 219.348 ; 
        RECT 44.464 214.974 44.568 219.348 ; 
        RECT 44.032 214.974 44.136 219.348 ; 
        RECT 43.6 214.974 43.704 219.348 ; 
        RECT 43.168 214.974 43.272 219.348 ; 
        RECT 42.736 214.974 42.84 219.348 ; 
        RECT 42.304 214.974 42.408 219.348 ; 
        RECT 41.872 214.974 41.976 219.348 ; 
        RECT 41.44 214.974 41.544 219.348 ; 
        RECT 41.008 214.974 41.112 219.348 ; 
        RECT 40.576 214.974 40.68 219.348 ; 
        RECT 40.144 214.974 40.248 219.348 ; 
        RECT 39.712 214.974 39.816 219.348 ; 
        RECT 39.28 214.974 39.384 219.348 ; 
        RECT 38.848 214.974 38.952 219.348 ; 
        RECT 38.416 214.974 38.52 219.348 ; 
        RECT 37.984 214.974 38.088 219.348 ; 
        RECT 37.552 214.974 37.656 219.348 ; 
        RECT 36.7 214.974 37.008 219.348 ; 
        RECT 29.128 214.974 29.436 219.348 ; 
        RECT 28.48 214.974 28.584 219.348 ; 
        RECT 28.048 214.974 28.152 219.348 ; 
        RECT 27.616 214.974 27.72 219.348 ; 
        RECT 27.184 214.974 27.288 219.348 ; 
        RECT 26.752 214.974 26.856 219.348 ; 
        RECT 26.32 214.974 26.424 219.348 ; 
        RECT 25.888 214.974 25.992 219.348 ; 
        RECT 25.456 214.974 25.56 219.348 ; 
        RECT 25.024 214.974 25.128 219.348 ; 
        RECT 24.592 214.974 24.696 219.348 ; 
        RECT 24.16 214.974 24.264 219.348 ; 
        RECT 23.728 214.974 23.832 219.348 ; 
        RECT 23.296 214.974 23.4 219.348 ; 
        RECT 22.864 214.974 22.968 219.348 ; 
        RECT 22.432 214.974 22.536 219.348 ; 
        RECT 22 214.974 22.104 219.348 ; 
        RECT 21.568 214.974 21.672 219.348 ; 
        RECT 21.136 214.974 21.24 219.348 ; 
        RECT 20.704 214.974 20.808 219.348 ; 
        RECT 20.272 214.974 20.376 219.348 ; 
        RECT 19.84 214.974 19.944 219.348 ; 
        RECT 19.408 214.974 19.512 219.348 ; 
        RECT 18.976 214.974 19.08 219.348 ; 
        RECT 18.544 214.974 18.648 219.348 ; 
        RECT 18.112 214.974 18.216 219.348 ; 
        RECT 17.68 214.974 17.784 219.348 ; 
        RECT 17.248 214.974 17.352 219.348 ; 
        RECT 16.816 214.974 16.92 219.348 ; 
        RECT 16.384 214.974 16.488 219.348 ; 
        RECT 15.952 214.974 16.056 219.348 ; 
        RECT 15.52 214.974 15.624 219.348 ; 
        RECT 15.088 214.974 15.192 219.348 ; 
        RECT 14.656 214.974 14.76 219.348 ; 
        RECT 14.224 214.974 14.328 219.348 ; 
        RECT 13.792 214.974 13.896 219.348 ; 
        RECT 13.36 214.974 13.464 219.348 ; 
        RECT 12.928 214.974 13.032 219.348 ; 
        RECT 12.496 214.974 12.6 219.348 ; 
        RECT 12.064 214.974 12.168 219.348 ; 
        RECT 11.632 214.974 11.736 219.348 ; 
        RECT 11.2 214.974 11.304 219.348 ; 
        RECT 10.768 214.974 10.872 219.348 ; 
        RECT 10.336 214.974 10.44 219.348 ; 
        RECT 9.904 214.974 10.008 219.348 ; 
        RECT 9.472 214.974 9.576 219.348 ; 
        RECT 9.04 214.974 9.144 219.348 ; 
        RECT 8.608 214.974 8.712 219.348 ; 
        RECT 8.176 214.974 8.28 219.348 ; 
        RECT 7.744 214.974 7.848 219.348 ; 
        RECT 7.312 214.974 7.416 219.348 ; 
        RECT 6.88 214.974 6.984 219.348 ; 
        RECT 6.448 214.974 6.552 219.348 ; 
        RECT 6.016 214.974 6.12 219.348 ; 
        RECT 5.584 214.974 5.688 219.348 ; 
        RECT 5.152 214.974 5.256 219.348 ; 
        RECT 4.72 214.974 4.824 219.348 ; 
        RECT 4.288 214.974 4.392 219.348 ; 
        RECT 3.856 214.974 3.96 219.348 ; 
        RECT 3.424 214.974 3.528 219.348 ; 
        RECT 2.992 214.974 3.096 219.348 ; 
        RECT 2.56 214.974 2.664 219.348 ; 
        RECT 2.128 214.974 2.232 219.348 ; 
        RECT 1.696 214.974 1.8 219.348 ; 
        RECT 1.264 214.974 1.368 219.348 ; 
        RECT 0.832 214.974 0.936 219.348 ; 
        RECT 0.02 214.974 0.36 219.348 ; 
        RECT 34.564 219.294 35.076 223.668 ; 
        RECT 34.508 221.956 35.076 223.246 ; 
        RECT 33.916 220.864 34.164 223.668 ; 
        RECT 33.86 222.102 34.164 222.716 ; 
        RECT 33.916 219.294 34.02 223.668 ; 
        RECT 33.916 219.778 34.076 220.736 ; 
        RECT 33.916 219.294 34.164 219.65 ; 
        RECT 32.728 221.096 33.552 223.668 ; 
        RECT 33.448 219.294 33.552 223.668 ; 
        RECT 32.728 222.204 33.608 223.236 ; 
        RECT 32.728 219.294 33.12 223.668 ; 
        RECT 31.06 219.294 31.392 223.668 ; 
        RECT 31.06 219.648 31.448 223.39 ; 
        RECT 65.776 219.294 66.116 223.668 ; 
        RECT 65.2 219.294 65.304 223.668 ; 
        RECT 64.768 219.294 64.872 223.668 ; 
        RECT 64.336 219.294 64.44 223.668 ; 
        RECT 63.904 219.294 64.008 223.668 ; 
        RECT 63.472 219.294 63.576 223.668 ; 
        RECT 63.04 219.294 63.144 223.668 ; 
        RECT 62.608 219.294 62.712 223.668 ; 
        RECT 62.176 219.294 62.28 223.668 ; 
        RECT 61.744 219.294 61.848 223.668 ; 
        RECT 61.312 219.294 61.416 223.668 ; 
        RECT 60.88 219.294 60.984 223.668 ; 
        RECT 60.448 219.294 60.552 223.668 ; 
        RECT 60.016 219.294 60.12 223.668 ; 
        RECT 59.584 219.294 59.688 223.668 ; 
        RECT 59.152 219.294 59.256 223.668 ; 
        RECT 58.72 219.294 58.824 223.668 ; 
        RECT 58.288 219.294 58.392 223.668 ; 
        RECT 57.856 219.294 57.96 223.668 ; 
        RECT 57.424 219.294 57.528 223.668 ; 
        RECT 56.992 219.294 57.096 223.668 ; 
        RECT 56.56 219.294 56.664 223.668 ; 
        RECT 56.128 219.294 56.232 223.668 ; 
        RECT 55.696 219.294 55.8 223.668 ; 
        RECT 55.264 219.294 55.368 223.668 ; 
        RECT 54.832 219.294 54.936 223.668 ; 
        RECT 54.4 219.294 54.504 223.668 ; 
        RECT 53.968 219.294 54.072 223.668 ; 
        RECT 53.536 219.294 53.64 223.668 ; 
        RECT 53.104 219.294 53.208 223.668 ; 
        RECT 52.672 219.294 52.776 223.668 ; 
        RECT 52.24 219.294 52.344 223.668 ; 
        RECT 51.808 219.294 51.912 223.668 ; 
        RECT 51.376 219.294 51.48 223.668 ; 
        RECT 50.944 219.294 51.048 223.668 ; 
        RECT 50.512 219.294 50.616 223.668 ; 
        RECT 50.08 219.294 50.184 223.668 ; 
        RECT 49.648 219.294 49.752 223.668 ; 
        RECT 49.216 219.294 49.32 223.668 ; 
        RECT 48.784 219.294 48.888 223.668 ; 
        RECT 48.352 219.294 48.456 223.668 ; 
        RECT 47.92 219.294 48.024 223.668 ; 
        RECT 47.488 219.294 47.592 223.668 ; 
        RECT 47.056 219.294 47.16 223.668 ; 
        RECT 46.624 219.294 46.728 223.668 ; 
        RECT 46.192 219.294 46.296 223.668 ; 
        RECT 45.76 219.294 45.864 223.668 ; 
        RECT 45.328 219.294 45.432 223.668 ; 
        RECT 44.896 219.294 45 223.668 ; 
        RECT 44.464 219.294 44.568 223.668 ; 
        RECT 44.032 219.294 44.136 223.668 ; 
        RECT 43.6 219.294 43.704 223.668 ; 
        RECT 43.168 219.294 43.272 223.668 ; 
        RECT 42.736 219.294 42.84 223.668 ; 
        RECT 42.304 219.294 42.408 223.668 ; 
        RECT 41.872 219.294 41.976 223.668 ; 
        RECT 41.44 219.294 41.544 223.668 ; 
        RECT 41.008 219.294 41.112 223.668 ; 
        RECT 40.576 219.294 40.68 223.668 ; 
        RECT 40.144 219.294 40.248 223.668 ; 
        RECT 39.712 219.294 39.816 223.668 ; 
        RECT 39.28 219.294 39.384 223.668 ; 
        RECT 38.848 219.294 38.952 223.668 ; 
        RECT 38.416 219.294 38.52 223.668 ; 
        RECT 37.984 219.294 38.088 223.668 ; 
        RECT 37.552 219.294 37.656 223.668 ; 
        RECT 36.7 219.294 37.008 223.668 ; 
        RECT 29.128 219.294 29.436 223.668 ; 
        RECT 28.48 219.294 28.584 223.668 ; 
        RECT 28.048 219.294 28.152 223.668 ; 
        RECT 27.616 219.294 27.72 223.668 ; 
        RECT 27.184 219.294 27.288 223.668 ; 
        RECT 26.752 219.294 26.856 223.668 ; 
        RECT 26.32 219.294 26.424 223.668 ; 
        RECT 25.888 219.294 25.992 223.668 ; 
        RECT 25.456 219.294 25.56 223.668 ; 
        RECT 25.024 219.294 25.128 223.668 ; 
        RECT 24.592 219.294 24.696 223.668 ; 
        RECT 24.16 219.294 24.264 223.668 ; 
        RECT 23.728 219.294 23.832 223.668 ; 
        RECT 23.296 219.294 23.4 223.668 ; 
        RECT 22.864 219.294 22.968 223.668 ; 
        RECT 22.432 219.294 22.536 223.668 ; 
        RECT 22 219.294 22.104 223.668 ; 
        RECT 21.568 219.294 21.672 223.668 ; 
        RECT 21.136 219.294 21.24 223.668 ; 
        RECT 20.704 219.294 20.808 223.668 ; 
        RECT 20.272 219.294 20.376 223.668 ; 
        RECT 19.84 219.294 19.944 223.668 ; 
        RECT 19.408 219.294 19.512 223.668 ; 
        RECT 18.976 219.294 19.08 223.668 ; 
        RECT 18.544 219.294 18.648 223.668 ; 
        RECT 18.112 219.294 18.216 223.668 ; 
        RECT 17.68 219.294 17.784 223.668 ; 
        RECT 17.248 219.294 17.352 223.668 ; 
        RECT 16.816 219.294 16.92 223.668 ; 
        RECT 16.384 219.294 16.488 223.668 ; 
        RECT 15.952 219.294 16.056 223.668 ; 
        RECT 15.52 219.294 15.624 223.668 ; 
        RECT 15.088 219.294 15.192 223.668 ; 
        RECT 14.656 219.294 14.76 223.668 ; 
        RECT 14.224 219.294 14.328 223.668 ; 
        RECT 13.792 219.294 13.896 223.668 ; 
        RECT 13.36 219.294 13.464 223.668 ; 
        RECT 12.928 219.294 13.032 223.668 ; 
        RECT 12.496 219.294 12.6 223.668 ; 
        RECT 12.064 219.294 12.168 223.668 ; 
        RECT 11.632 219.294 11.736 223.668 ; 
        RECT 11.2 219.294 11.304 223.668 ; 
        RECT 10.768 219.294 10.872 223.668 ; 
        RECT 10.336 219.294 10.44 223.668 ; 
        RECT 9.904 219.294 10.008 223.668 ; 
        RECT 9.472 219.294 9.576 223.668 ; 
        RECT 9.04 219.294 9.144 223.668 ; 
        RECT 8.608 219.294 8.712 223.668 ; 
        RECT 8.176 219.294 8.28 223.668 ; 
        RECT 7.744 219.294 7.848 223.668 ; 
        RECT 7.312 219.294 7.416 223.668 ; 
        RECT 6.88 219.294 6.984 223.668 ; 
        RECT 6.448 219.294 6.552 223.668 ; 
        RECT 6.016 219.294 6.12 223.668 ; 
        RECT 5.584 219.294 5.688 223.668 ; 
        RECT 5.152 219.294 5.256 223.668 ; 
        RECT 4.72 219.294 4.824 223.668 ; 
        RECT 4.288 219.294 4.392 223.668 ; 
        RECT 3.856 219.294 3.96 223.668 ; 
        RECT 3.424 219.294 3.528 223.668 ; 
        RECT 2.992 219.294 3.096 223.668 ; 
        RECT 2.56 219.294 2.664 223.668 ; 
        RECT 2.128 219.294 2.232 223.668 ; 
        RECT 1.696 219.294 1.8 223.668 ; 
        RECT 1.264 219.294 1.368 223.668 ; 
        RECT 0.832 219.294 0.936 223.668 ; 
        RECT 0.02 219.294 0.36 223.668 ; 
        RECT 34.564 223.614 35.076 227.988 ; 
        RECT 34.508 226.276 35.076 227.566 ; 
        RECT 33.916 225.184 34.164 227.988 ; 
        RECT 33.86 226.422 34.164 227.036 ; 
        RECT 33.916 223.614 34.02 227.988 ; 
        RECT 33.916 224.098 34.076 225.056 ; 
        RECT 33.916 223.614 34.164 223.97 ; 
        RECT 32.728 225.416 33.552 227.988 ; 
        RECT 33.448 223.614 33.552 227.988 ; 
        RECT 32.728 226.524 33.608 227.556 ; 
        RECT 32.728 223.614 33.12 227.988 ; 
        RECT 31.06 223.614 31.392 227.988 ; 
        RECT 31.06 223.968 31.448 227.71 ; 
        RECT 65.776 223.614 66.116 227.988 ; 
        RECT 65.2 223.614 65.304 227.988 ; 
        RECT 64.768 223.614 64.872 227.988 ; 
        RECT 64.336 223.614 64.44 227.988 ; 
        RECT 63.904 223.614 64.008 227.988 ; 
        RECT 63.472 223.614 63.576 227.988 ; 
        RECT 63.04 223.614 63.144 227.988 ; 
        RECT 62.608 223.614 62.712 227.988 ; 
        RECT 62.176 223.614 62.28 227.988 ; 
        RECT 61.744 223.614 61.848 227.988 ; 
        RECT 61.312 223.614 61.416 227.988 ; 
        RECT 60.88 223.614 60.984 227.988 ; 
        RECT 60.448 223.614 60.552 227.988 ; 
        RECT 60.016 223.614 60.12 227.988 ; 
        RECT 59.584 223.614 59.688 227.988 ; 
        RECT 59.152 223.614 59.256 227.988 ; 
        RECT 58.72 223.614 58.824 227.988 ; 
        RECT 58.288 223.614 58.392 227.988 ; 
        RECT 57.856 223.614 57.96 227.988 ; 
        RECT 57.424 223.614 57.528 227.988 ; 
        RECT 56.992 223.614 57.096 227.988 ; 
        RECT 56.56 223.614 56.664 227.988 ; 
        RECT 56.128 223.614 56.232 227.988 ; 
        RECT 55.696 223.614 55.8 227.988 ; 
        RECT 55.264 223.614 55.368 227.988 ; 
        RECT 54.832 223.614 54.936 227.988 ; 
        RECT 54.4 223.614 54.504 227.988 ; 
        RECT 53.968 223.614 54.072 227.988 ; 
        RECT 53.536 223.614 53.64 227.988 ; 
        RECT 53.104 223.614 53.208 227.988 ; 
        RECT 52.672 223.614 52.776 227.988 ; 
        RECT 52.24 223.614 52.344 227.988 ; 
        RECT 51.808 223.614 51.912 227.988 ; 
        RECT 51.376 223.614 51.48 227.988 ; 
        RECT 50.944 223.614 51.048 227.988 ; 
        RECT 50.512 223.614 50.616 227.988 ; 
        RECT 50.08 223.614 50.184 227.988 ; 
        RECT 49.648 223.614 49.752 227.988 ; 
        RECT 49.216 223.614 49.32 227.988 ; 
        RECT 48.784 223.614 48.888 227.988 ; 
        RECT 48.352 223.614 48.456 227.988 ; 
        RECT 47.92 223.614 48.024 227.988 ; 
        RECT 47.488 223.614 47.592 227.988 ; 
        RECT 47.056 223.614 47.16 227.988 ; 
        RECT 46.624 223.614 46.728 227.988 ; 
        RECT 46.192 223.614 46.296 227.988 ; 
        RECT 45.76 223.614 45.864 227.988 ; 
        RECT 45.328 223.614 45.432 227.988 ; 
        RECT 44.896 223.614 45 227.988 ; 
        RECT 44.464 223.614 44.568 227.988 ; 
        RECT 44.032 223.614 44.136 227.988 ; 
        RECT 43.6 223.614 43.704 227.988 ; 
        RECT 43.168 223.614 43.272 227.988 ; 
        RECT 42.736 223.614 42.84 227.988 ; 
        RECT 42.304 223.614 42.408 227.988 ; 
        RECT 41.872 223.614 41.976 227.988 ; 
        RECT 41.44 223.614 41.544 227.988 ; 
        RECT 41.008 223.614 41.112 227.988 ; 
        RECT 40.576 223.614 40.68 227.988 ; 
        RECT 40.144 223.614 40.248 227.988 ; 
        RECT 39.712 223.614 39.816 227.988 ; 
        RECT 39.28 223.614 39.384 227.988 ; 
        RECT 38.848 223.614 38.952 227.988 ; 
        RECT 38.416 223.614 38.52 227.988 ; 
        RECT 37.984 223.614 38.088 227.988 ; 
        RECT 37.552 223.614 37.656 227.988 ; 
        RECT 36.7 223.614 37.008 227.988 ; 
        RECT 29.128 223.614 29.436 227.988 ; 
        RECT 28.48 223.614 28.584 227.988 ; 
        RECT 28.048 223.614 28.152 227.988 ; 
        RECT 27.616 223.614 27.72 227.988 ; 
        RECT 27.184 223.614 27.288 227.988 ; 
        RECT 26.752 223.614 26.856 227.988 ; 
        RECT 26.32 223.614 26.424 227.988 ; 
        RECT 25.888 223.614 25.992 227.988 ; 
        RECT 25.456 223.614 25.56 227.988 ; 
        RECT 25.024 223.614 25.128 227.988 ; 
        RECT 24.592 223.614 24.696 227.988 ; 
        RECT 24.16 223.614 24.264 227.988 ; 
        RECT 23.728 223.614 23.832 227.988 ; 
        RECT 23.296 223.614 23.4 227.988 ; 
        RECT 22.864 223.614 22.968 227.988 ; 
        RECT 22.432 223.614 22.536 227.988 ; 
        RECT 22 223.614 22.104 227.988 ; 
        RECT 21.568 223.614 21.672 227.988 ; 
        RECT 21.136 223.614 21.24 227.988 ; 
        RECT 20.704 223.614 20.808 227.988 ; 
        RECT 20.272 223.614 20.376 227.988 ; 
        RECT 19.84 223.614 19.944 227.988 ; 
        RECT 19.408 223.614 19.512 227.988 ; 
        RECT 18.976 223.614 19.08 227.988 ; 
        RECT 18.544 223.614 18.648 227.988 ; 
        RECT 18.112 223.614 18.216 227.988 ; 
        RECT 17.68 223.614 17.784 227.988 ; 
        RECT 17.248 223.614 17.352 227.988 ; 
        RECT 16.816 223.614 16.92 227.988 ; 
        RECT 16.384 223.614 16.488 227.988 ; 
        RECT 15.952 223.614 16.056 227.988 ; 
        RECT 15.52 223.614 15.624 227.988 ; 
        RECT 15.088 223.614 15.192 227.988 ; 
        RECT 14.656 223.614 14.76 227.988 ; 
        RECT 14.224 223.614 14.328 227.988 ; 
        RECT 13.792 223.614 13.896 227.988 ; 
        RECT 13.36 223.614 13.464 227.988 ; 
        RECT 12.928 223.614 13.032 227.988 ; 
        RECT 12.496 223.614 12.6 227.988 ; 
        RECT 12.064 223.614 12.168 227.988 ; 
        RECT 11.632 223.614 11.736 227.988 ; 
        RECT 11.2 223.614 11.304 227.988 ; 
        RECT 10.768 223.614 10.872 227.988 ; 
        RECT 10.336 223.614 10.44 227.988 ; 
        RECT 9.904 223.614 10.008 227.988 ; 
        RECT 9.472 223.614 9.576 227.988 ; 
        RECT 9.04 223.614 9.144 227.988 ; 
        RECT 8.608 223.614 8.712 227.988 ; 
        RECT 8.176 223.614 8.28 227.988 ; 
        RECT 7.744 223.614 7.848 227.988 ; 
        RECT 7.312 223.614 7.416 227.988 ; 
        RECT 6.88 223.614 6.984 227.988 ; 
        RECT 6.448 223.614 6.552 227.988 ; 
        RECT 6.016 223.614 6.12 227.988 ; 
        RECT 5.584 223.614 5.688 227.988 ; 
        RECT 5.152 223.614 5.256 227.988 ; 
        RECT 4.72 223.614 4.824 227.988 ; 
        RECT 4.288 223.614 4.392 227.988 ; 
        RECT 3.856 223.614 3.96 227.988 ; 
        RECT 3.424 223.614 3.528 227.988 ; 
        RECT 2.992 223.614 3.096 227.988 ; 
        RECT 2.56 223.614 2.664 227.988 ; 
        RECT 2.128 223.614 2.232 227.988 ; 
        RECT 1.696 223.614 1.8 227.988 ; 
        RECT 1.264 223.614 1.368 227.988 ; 
        RECT 0.832 223.614 0.936 227.988 ; 
        RECT 0.02 223.614 0.36 227.988 ; 
        RECT 34.564 227.934 35.076 232.308 ; 
        RECT 34.508 230.596 35.076 231.886 ; 
        RECT 33.916 229.504 34.164 232.308 ; 
        RECT 33.86 230.742 34.164 231.356 ; 
        RECT 33.916 227.934 34.02 232.308 ; 
        RECT 33.916 228.418 34.076 229.376 ; 
        RECT 33.916 227.934 34.164 228.29 ; 
        RECT 32.728 229.736 33.552 232.308 ; 
        RECT 33.448 227.934 33.552 232.308 ; 
        RECT 32.728 230.844 33.608 231.876 ; 
        RECT 32.728 227.934 33.12 232.308 ; 
        RECT 31.06 227.934 31.392 232.308 ; 
        RECT 31.06 228.288 31.448 232.03 ; 
        RECT 65.776 227.934 66.116 232.308 ; 
        RECT 65.2 227.934 65.304 232.308 ; 
        RECT 64.768 227.934 64.872 232.308 ; 
        RECT 64.336 227.934 64.44 232.308 ; 
        RECT 63.904 227.934 64.008 232.308 ; 
        RECT 63.472 227.934 63.576 232.308 ; 
        RECT 63.04 227.934 63.144 232.308 ; 
        RECT 62.608 227.934 62.712 232.308 ; 
        RECT 62.176 227.934 62.28 232.308 ; 
        RECT 61.744 227.934 61.848 232.308 ; 
        RECT 61.312 227.934 61.416 232.308 ; 
        RECT 60.88 227.934 60.984 232.308 ; 
        RECT 60.448 227.934 60.552 232.308 ; 
        RECT 60.016 227.934 60.12 232.308 ; 
        RECT 59.584 227.934 59.688 232.308 ; 
        RECT 59.152 227.934 59.256 232.308 ; 
        RECT 58.72 227.934 58.824 232.308 ; 
        RECT 58.288 227.934 58.392 232.308 ; 
        RECT 57.856 227.934 57.96 232.308 ; 
        RECT 57.424 227.934 57.528 232.308 ; 
        RECT 56.992 227.934 57.096 232.308 ; 
        RECT 56.56 227.934 56.664 232.308 ; 
        RECT 56.128 227.934 56.232 232.308 ; 
        RECT 55.696 227.934 55.8 232.308 ; 
        RECT 55.264 227.934 55.368 232.308 ; 
        RECT 54.832 227.934 54.936 232.308 ; 
        RECT 54.4 227.934 54.504 232.308 ; 
        RECT 53.968 227.934 54.072 232.308 ; 
        RECT 53.536 227.934 53.64 232.308 ; 
        RECT 53.104 227.934 53.208 232.308 ; 
        RECT 52.672 227.934 52.776 232.308 ; 
        RECT 52.24 227.934 52.344 232.308 ; 
        RECT 51.808 227.934 51.912 232.308 ; 
        RECT 51.376 227.934 51.48 232.308 ; 
        RECT 50.944 227.934 51.048 232.308 ; 
        RECT 50.512 227.934 50.616 232.308 ; 
        RECT 50.08 227.934 50.184 232.308 ; 
        RECT 49.648 227.934 49.752 232.308 ; 
        RECT 49.216 227.934 49.32 232.308 ; 
        RECT 48.784 227.934 48.888 232.308 ; 
        RECT 48.352 227.934 48.456 232.308 ; 
        RECT 47.92 227.934 48.024 232.308 ; 
        RECT 47.488 227.934 47.592 232.308 ; 
        RECT 47.056 227.934 47.16 232.308 ; 
        RECT 46.624 227.934 46.728 232.308 ; 
        RECT 46.192 227.934 46.296 232.308 ; 
        RECT 45.76 227.934 45.864 232.308 ; 
        RECT 45.328 227.934 45.432 232.308 ; 
        RECT 44.896 227.934 45 232.308 ; 
        RECT 44.464 227.934 44.568 232.308 ; 
        RECT 44.032 227.934 44.136 232.308 ; 
        RECT 43.6 227.934 43.704 232.308 ; 
        RECT 43.168 227.934 43.272 232.308 ; 
        RECT 42.736 227.934 42.84 232.308 ; 
        RECT 42.304 227.934 42.408 232.308 ; 
        RECT 41.872 227.934 41.976 232.308 ; 
        RECT 41.44 227.934 41.544 232.308 ; 
        RECT 41.008 227.934 41.112 232.308 ; 
        RECT 40.576 227.934 40.68 232.308 ; 
        RECT 40.144 227.934 40.248 232.308 ; 
        RECT 39.712 227.934 39.816 232.308 ; 
        RECT 39.28 227.934 39.384 232.308 ; 
        RECT 38.848 227.934 38.952 232.308 ; 
        RECT 38.416 227.934 38.52 232.308 ; 
        RECT 37.984 227.934 38.088 232.308 ; 
        RECT 37.552 227.934 37.656 232.308 ; 
        RECT 36.7 227.934 37.008 232.308 ; 
        RECT 29.128 227.934 29.436 232.308 ; 
        RECT 28.48 227.934 28.584 232.308 ; 
        RECT 28.048 227.934 28.152 232.308 ; 
        RECT 27.616 227.934 27.72 232.308 ; 
        RECT 27.184 227.934 27.288 232.308 ; 
        RECT 26.752 227.934 26.856 232.308 ; 
        RECT 26.32 227.934 26.424 232.308 ; 
        RECT 25.888 227.934 25.992 232.308 ; 
        RECT 25.456 227.934 25.56 232.308 ; 
        RECT 25.024 227.934 25.128 232.308 ; 
        RECT 24.592 227.934 24.696 232.308 ; 
        RECT 24.16 227.934 24.264 232.308 ; 
        RECT 23.728 227.934 23.832 232.308 ; 
        RECT 23.296 227.934 23.4 232.308 ; 
        RECT 22.864 227.934 22.968 232.308 ; 
        RECT 22.432 227.934 22.536 232.308 ; 
        RECT 22 227.934 22.104 232.308 ; 
        RECT 21.568 227.934 21.672 232.308 ; 
        RECT 21.136 227.934 21.24 232.308 ; 
        RECT 20.704 227.934 20.808 232.308 ; 
        RECT 20.272 227.934 20.376 232.308 ; 
        RECT 19.84 227.934 19.944 232.308 ; 
        RECT 19.408 227.934 19.512 232.308 ; 
        RECT 18.976 227.934 19.08 232.308 ; 
        RECT 18.544 227.934 18.648 232.308 ; 
        RECT 18.112 227.934 18.216 232.308 ; 
        RECT 17.68 227.934 17.784 232.308 ; 
        RECT 17.248 227.934 17.352 232.308 ; 
        RECT 16.816 227.934 16.92 232.308 ; 
        RECT 16.384 227.934 16.488 232.308 ; 
        RECT 15.952 227.934 16.056 232.308 ; 
        RECT 15.52 227.934 15.624 232.308 ; 
        RECT 15.088 227.934 15.192 232.308 ; 
        RECT 14.656 227.934 14.76 232.308 ; 
        RECT 14.224 227.934 14.328 232.308 ; 
        RECT 13.792 227.934 13.896 232.308 ; 
        RECT 13.36 227.934 13.464 232.308 ; 
        RECT 12.928 227.934 13.032 232.308 ; 
        RECT 12.496 227.934 12.6 232.308 ; 
        RECT 12.064 227.934 12.168 232.308 ; 
        RECT 11.632 227.934 11.736 232.308 ; 
        RECT 11.2 227.934 11.304 232.308 ; 
        RECT 10.768 227.934 10.872 232.308 ; 
        RECT 10.336 227.934 10.44 232.308 ; 
        RECT 9.904 227.934 10.008 232.308 ; 
        RECT 9.472 227.934 9.576 232.308 ; 
        RECT 9.04 227.934 9.144 232.308 ; 
        RECT 8.608 227.934 8.712 232.308 ; 
        RECT 8.176 227.934 8.28 232.308 ; 
        RECT 7.744 227.934 7.848 232.308 ; 
        RECT 7.312 227.934 7.416 232.308 ; 
        RECT 6.88 227.934 6.984 232.308 ; 
        RECT 6.448 227.934 6.552 232.308 ; 
        RECT 6.016 227.934 6.12 232.308 ; 
        RECT 5.584 227.934 5.688 232.308 ; 
        RECT 5.152 227.934 5.256 232.308 ; 
        RECT 4.72 227.934 4.824 232.308 ; 
        RECT 4.288 227.934 4.392 232.308 ; 
        RECT 3.856 227.934 3.96 232.308 ; 
        RECT 3.424 227.934 3.528 232.308 ; 
        RECT 2.992 227.934 3.096 232.308 ; 
        RECT 2.56 227.934 2.664 232.308 ; 
        RECT 2.128 227.934 2.232 232.308 ; 
        RECT 1.696 227.934 1.8 232.308 ; 
        RECT 1.264 227.934 1.368 232.308 ; 
        RECT 0.832 227.934 0.936 232.308 ; 
        RECT 0.02 227.934 0.36 232.308 ; 
        RECT 34.564 232.254 35.076 236.628 ; 
        RECT 34.508 234.916 35.076 236.206 ; 
        RECT 33.916 233.824 34.164 236.628 ; 
        RECT 33.86 235.062 34.164 235.676 ; 
        RECT 33.916 232.254 34.02 236.628 ; 
        RECT 33.916 232.738 34.076 233.696 ; 
        RECT 33.916 232.254 34.164 232.61 ; 
        RECT 32.728 234.056 33.552 236.628 ; 
        RECT 33.448 232.254 33.552 236.628 ; 
        RECT 32.728 235.164 33.608 236.196 ; 
        RECT 32.728 232.254 33.12 236.628 ; 
        RECT 31.06 232.254 31.392 236.628 ; 
        RECT 31.06 232.608 31.448 236.35 ; 
        RECT 65.776 232.254 66.116 236.628 ; 
        RECT 65.2 232.254 65.304 236.628 ; 
        RECT 64.768 232.254 64.872 236.628 ; 
        RECT 64.336 232.254 64.44 236.628 ; 
        RECT 63.904 232.254 64.008 236.628 ; 
        RECT 63.472 232.254 63.576 236.628 ; 
        RECT 63.04 232.254 63.144 236.628 ; 
        RECT 62.608 232.254 62.712 236.628 ; 
        RECT 62.176 232.254 62.28 236.628 ; 
        RECT 61.744 232.254 61.848 236.628 ; 
        RECT 61.312 232.254 61.416 236.628 ; 
        RECT 60.88 232.254 60.984 236.628 ; 
        RECT 60.448 232.254 60.552 236.628 ; 
        RECT 60.016 232.254 60.12 236.628 ; 
        RECT 59.584 232.254 59.688 236.628 ; 
        RECT 59.152 232.254 59.256 236.628 ; 
        RECT 58.72 232.254 58.824 236.628 ; 
        RECT 58.288 232.254 58.392 236.628 ; 
        RECT 57.856 232.254 57.96 236.628 ; 
        RECT 57.424 232.254 57.528 236.628 ; 
        RECT 56.992 232.254 57.096 236.628 ; 
        RECT 56.56 232.254 56.664 236.628 ; 
        RECT 56.128 232.254 56.232 236.628 ; 
        RECT 55.696 232.254 55.8 236.628 ; 
        RECT 55.264 232.254 55.368 236.628 ; 
        RECT 54.832 232.254 54.936 236.628 ; 
        RECT 54.4 232.254 54.504 236.628 ; 
        RECT 53.968 232.254 54.072 236.628 ; 
        RECT 53.536 232.254 53.64 236.628 ; 
        RECT 53.104 232.254 53.208 236.628 ; 
        RECT 52.672 232.254 52.776 236.628 ; 
        RECT 52.24 232.254 52.344 236.628 ; 
        RECT 51.808 232.254 51.912 236.628 ; 
        RECT 51.376 232.254 51.48 236.628 ; 
        RECT 50.944 232.254 51.048 236.628 ; 
        RECT 50.512 232.254 50.616 236.628 ; 
        RECT 50.08 232.254 50.184 236.628 ; 
        RECT 49.648 232.254 49.752 236.628 ; 
        RECT 49.216 232.254 49.32 236.628 ; 
        RECT 48.784 232.254 48.888 236.628 ; 
        RECT 48.352 232.254 48.456 236.628 ; 
        RECT 47.92 232.254 48.024 236.628 ; 
        RECT 47.488 232.254 47.592 236.628 ; 
        RECT 47.056 232.254 47.16 236.628 ; 
        RECT 46.624 232.254 46.728 236.628 ; 
        RECT 46.192 232.254 46.296 236.628 ; 
        RECT 45.76 232.254 45.864 236.628 ; 
        RECT 45.328 232.254 45.432 236.628 ; 
        RECT 44.896 232.254 45 236.628 ; 
        RECT 44.464 232.254 44.568 236.628 ; 
        RECT 44.032 232.254 44.136 236.628 ; 
        RECT 43.6 232.254 43.704 236.628 ; 
        RECT 43.168 232.254 43.272 236.628 ; 
        RECT 42.736 232.254 42.84 236.628 ; 
        RECT 42.304 232.254 42.408 236.628 ; 
        RECT 41.872 232.254 41.976 236.628 ; 
        RECT 41.44 232.254 41.544 236.628 ; 
        RECT 41.008 232.254 41.112 236.628 ; 
        RECT 40.576 232.254 40.68 236.628 ; 
        RECT 40.144 232.254 40.248 236.628 ; 
        RECT 39.712 232.254 39.816 236.628 ; 
        RECT 39.28 232.254 39.384 236.628 ; 
        RECT 38.848 232.254 38.952 236.628 ; 
        RECT 38.416 232.254 38.52 236.628 ; 
        RECT 37.984 232.254 38.088 236.628 ; 
        RECT 37.552 232.254 37.656 236.628 ; 
        RECT 36.7 232.254 37.008 236.628 ; 
        RECT 29.128 232.254 29.436 236.628 ; 
        RECT 28.48 232.254 28.584 236.628 ; 
        RECT 28.048 232.254 28.152 236.628 ; 
        RECT 27.616 232.254 27.72 236.628 ; 
        RECT 27.184 232.254 27.288 236.628 ; 
        RECT 26.752 232.254 26.856 236.628 ; 
        RECT 26.32 232.254 26.424 236.628 ; 
        RECT 25.888 232.254 25.992 236.628 ; 
        RECT 25.456 232.254 25.56 236.628 ; 
        RECT 25.024 232.254 25.128 236.628 ; 
        RECT 24.592 232.254 24.696 236.628 ; 
        RECT 24.16 232.254 24.264 236.628 ; 
        RECT 23.728 232.254 23.832 236.628 ; 
        RECT 23.296 232.254 23.4 236.628 ; 
        RECT 22.864 232.254 22.968 236.628 ; 
        RECT 22.432 232.254 22.536 236.628 ; 
        RECT 22 232.254 22.104 236.628 ; 
        RECT 21.568 232.254 21.672 236.628 ; 
        RECT 21.136 232.254 21.24 236.628 ; 
        RECT 20.704 232.254 20.808 236.628 ; 
        RECT 20.272 232.254 20.376 236.628 ; 
        RECT 19.84 232.254 19.944 236.628 ; 
        RECT 19.408 232.254 19.512 236.628 ; 
        RECT 18.976 232.254 19.08 236.628 ; 
        RECT 18.544 232.254 18.648 236.628 ; 
        RECT 18.112 232.254 18.216 236.628 ; 
        RECT 17.68 232.254 17.784 236.628 ; 
        RECT 17.248 232.254 17.352 236.628 ; 
        RECT 16.816 232.254 16.92 236.628 ; 
        RECT 16.384 232.254 16.488 236.628 ; 
        RECT 15.952 232.254 16.056 236.628 ; 
        RECT 15.52 232.254 15.624 236.628 ; 
        RECT 15.088 232.254 15.192 236.628 ; 
        RECT 14.656 232.254 14.76 236.628 ; 
        RECT 14.224 232.254 14.328 236.628 ; 
        RECT 13.792 232.254 13.896 236.628 ; 
        RECT 13.36 232.254 13.464 236.628 ; 
        RECT 12.928 232.254 13.032 236.628 ; 
        RECT 12.496 232.254 12.6 236.628 ; 
        RECT 12.064 232.254 12.168 236.628 ; 
        RECT 11.632 232.254 11.736 236.628 ; 
        RECT 11.2 232.254 11.304 236.628 ; 
        RECT 10.768 232.254 10.872 236.628 ; 
        RECT 10.336 232.254 10.44 236.628 ; 
        RECT 9.904 232.254 10.008 236.628 ; 
        RECT 9.472 232.254 9.576 236.628 ; 
        RECT 9.04 232.254 9.144 236.628 ; 
        RECT 8.608 232.254 8.712 236.628 ; 
        RECT 8.176 232.254 8.28 236.628 ; 
        RECT 7.744 232.254 7.848 236.628 ; 
        RECT 7.312 232.254 7.416 236.628 ; 
        RECT 6.88 232.254 6.984 236.628 ; 
        RECT 6.448 232.254 6.552 236.628 ; 
        RECT 6.016 232.254 6.12 236.628 ; 
        RECT 5.584 232.254 5.688 236.628 ; 
        RECT 5.152 232.254 5.256 236.628 ; 
        RECT 4.72 232.254 4.824 236.628 ; 
        RECT 4.288 232.254 4.392 236.628 ; 
        RECT 3.856 232.254 3.96 236.628 ; 
        RECT 3.424 232.254 3.528 236.628 ; 
        RECT 2.992 232.254 3.096 236.628 ; 
        RECT 2.56 232.254 2.664 236.628 ; 
        RECT 2.128 232.254 2.232 236.628 ; 
        RECT 1.696 232.254 1.8 236.628 ; 
        RECT 1.264 232.254 1.368 236.628 ; 
        RECT 0.832 232.254 0.936 236.628 ; 
        RECT 0.02 232.254 0.36 236.628 ; 
        RECT 34.564 236.574 35.076 240.948 ; 
        RECT 34.508 239.236 35.076 240.526 ; 
        RECT 33.916 238.144 34.164 240.948 ; 
        RECT 33.86 239.382 34.164 239.996 ; 
        RECT 33.916 236.574 34.02 240.948 ; 
        RECT 33.916 237.058 34.076 238.016 ; 
        RECT 33.916 236.574 34.164 236.93 ; 
        RECT 32.728 238.376 33.552 240.948 ; 
        RECT 33.448 236.574 33.552 240.948 ; 
        RECT 32.728 239.484 33.608 240.516 ; 
        RECT 32.728 236.574 33.12 240.948 ; 
        RECT 31.06 236.574 31.392 240.948 ; 
        RECT 31.06 236.928 31.448 240.67 ; 
        RECT 65.776 236.574 66.116 240.948 ; 
        RECT 65.2 236.574 65.304 240.948 ; 
        RECT 64.768 236.574 64.872 240.948 ; 
        RECT 64.336 236.574 64.44 240.948 ; 
        RECT 63.904 236.574 64.008 240.948 ; 
        RECT 63.472 236.574 63.576 240.948 ; 
        RECT 63.04 236.574 63.144 240.948 ; 
        RECT 62.608 236.574 62.712 240.948 ; 
        RECT 62.176 236.574 62.28 240.948 ; 
        RECT 61.744 236.574 61.848 240.948 ; 
        RECT 61.312 236.574 61.416 240.948 ; 
        RECT 60.88 236.574 60.984 240.948 ; 
        RECT 60.448 236.574 60.552 240.948 ; 
        RECT 60.016 236.574 60.12 240.948 ; 
        RECT 59.584 236.574 59.688 240.948 ; 
        RECT 59.152 236.574 59.256 240.948 ; 
        RECT 58.72 236.574 58.824 240.948 ; 
        RECT 58.288 236.574 58.392 240.948 ; 
        RECT 57.856 236.574 57.96 240.948 ; 
        RECT 57.424 236.574 57.528 240.948 ; 
        RECT 56.992 236.574 57.096 240.948 ; 
        RECT 56.56 236.574 56.664 240.948 ; 
        RECT 56.128 236.574 56.232 240.948 ; 
        RECT 55.696 236.574 55.8 240.948 ; 
        RECT 55.264 236.574 55.368 240.948 ; 
        RECT 54.832 236.574 54.936 240.948 ; 
        RECT 54.4 236.574 54.504 240.948 ; 
        RECT 53.968 236.574 54.072 240.948 ; 
        RECT 53.536 236.574 53.64 240.948 ; 
        RECT 53.104 236.574 53.208 240.948 ; 
        RECT 52.672 236.574 52.776 240.948 ; 
        RECT 52.24 236.574 52.344 240.948 ; 
        RECT 51.808 236.574 51.912 240.948 ; 
        RECT 51.376 236.574 51.48 240.948 ; 
        RECT 50.944 236.574 51.048 240.948 ; 
        RECT 50.512 236.574 50.616 240.948 ; 
        RECT 50.08 236.574 50.184 240.948 ; 
        RECT 49.648 236.574 49.752 240.948 ; 
        RECT 49.216 236.574 49.32 240.948 ; 
        RECT 48.784 236.574 48.888 240.948 ; 
        RECT 48.352 236.574 48.456 240.948 ; 
        RECT 47.92 236.574 48.024 240.948 ; 
        RECT 47.488 236.574 47.592 240.948 ; 
        RECT 47.056 236.574 47.16 240.948 ; 
        RECT 46.624 236.574 46.728 240.948 ; 
        RECT 46.192 236.574 46.296 240.948 ; 
        RECT 45.76 236.574 45.864 240.948 ; 
        RECT 45.328 236.574 45.432 240.948 ; 
        RECT 44.896 236.574 45 240.948 ; 
        RECT 44.464 236.574 44.568 240.948 ; 
        RECT 44.032 236.574 44.136 240.948 ; 
        RECT 43.6 236.574 43.704 240.948 ; 
        RECT 43.168 236.574 43.272 240.948 ; 
        RECT 42.736 236.574 42.84 240.948 ; 
        RECT 42.304 236.574 42.408 240.948 ; 
        RECT 41.872 236.574 41.976 240.948 ; 
        RECT 41.44 236.574 41.544 240.948 ; 
        RECT 41.008 236.574 41.112 240.948 ; 
        RECT 40.576 236.574 40.68 240.948 ; 
        RECT 40.144 236.574 40.248 240.948 ; 
        RECT 39.712 236.574 39.816 240.948 ; 
        RECT 39.28 236.574 39.384 240.948 ; 
        RECT 38.848 236.574 38.952 240.948 ; 
        RECT 38.416 236.574 38.52 240.948 ; 
        RECT 37.984 236.574 38.088 240.948 ; 
        RECT 37.552 236.574 37.656 240.948 ; 
        RECT 36.7 236.574 37.008 240.948 ; 
        RECT 29.128 236.574 29.436 240.948 ; 
        RECT 28.48 236.574 28.584 240.948 ; 
        RECT 28.048 236.574 28.152 240.948 ; 
        RECT 27.616 236.574 27.72 240.948 ; 
        RECT 27.184 236.574 27.288 240.948 ; 
        RECT 26.752 236.574 26.856 240.948 ; 
        RECT 26.32 236.574 26.424 240.948 ; 
        RECT 25.888 236.574 25.992 240.948 ; 
        RECT 25.456 236.574 25.56 240.948 ; 
        RECT 25.024 236.574 25.128 240.948 ; 
        RECT 24.592 236.574 24.696 240.948 ; 
        RECT 24.16 236.574 24.264 240.948 ; 
        RECT 23.728 236.574 23.832 240.948 ; 
        RECT 23.296 236.574 23.4 240.948 ; 
        RECT 22.864 236.574 22.968 240.948 ; 
        RECT 22.432 236.574 22.536 240.948 ; 
        RECT 22 236.574 22.104 240.948 ; 
        RECT 21.568 236.574 21.672 240.948 ; 
        RECT 21.136 236.574 21.24 240.948 ; 
        RECT 20.704 236.574 20.808 240.948 ; 
        RECT 20.272 236.574 20.376 240.948 ; 
        RECT 19.84 236.574 19.944 240.948 ; 
        RECT 19.408 236.574 19.512 240.948 ; 
        RECT 18.976 236.574 19.08 240.948 ; 
        RECT 18.544 236.574 18.648 240.948 ; 
        RECT 18.112 236.574 18.216 240.948 ; 
        RECT 17.68 236.574 17.784 240.948 ; 
        RECT 17.248 236.574 17.352 240.948 ; 
        RECT 16.816 236.574 16.92 240.948 ; 
        RECT 16.384 236.574 16.488 240.948 ; 
        RECT 15.952 236.574 16.056 240.948 ; 
        RECT 15.52 236.574 15.624 240.948 ; 
        RECT 15.088 236.574 15.192 240.948 ; 
        RECT 14.656 236.574 14.76 240.948 ; 
        RECT 14.224 236.574 14.328 240.948 ; 
        RECT 13.792 236.574 13.896 240.948 ; 
        RECT 13.36 236.574 13.464 240.948 ; 
        RECT 12.928 236.574 13.032 240.948 ; 
        RECT 12.496 236.574 12.6 240.948 ; 
        RECT 12.064 236.574 12.168 240.948 ; 
        RECT 11.632 236.574 11.736 240.948 ; 
        RECT 11.2 236.574 11.304 240.948 ; 
        RECT 10.768 236.574 10.872 240.948 ; 
        RECT 10.336 236.574 10.44 240.948 ; 
        RECT 9.904 236.574 10.008 240.948 ; 
        RECT 9.472 236.574 9.576 240.948 ; 
        RECT 9.04 236.574 9.144 240.948 ; 
        RECT 8.608 236.574 8.712 240.948 ; 
        RECT 8.176 236.574 8.28 240.948 ; 
        RECT 7.744 236.574 7.848 240.948 ; 
        RECT 7.312 236.574 7.416 240.948 ; 
        RECT 6.88 236.574 6.984 240.948 ; 
        RECT 6.448 236.574 6.552 240.948 ; 
        RECT 6.016 236.574 6.12 240.948 ; 
        RECT 5.584 236.574 5.688 240.948 ; 
        RECT 5.152 236.574 5.256 240.948 ; 
        RECT 4.72 236.574 4.824 240.948 ; 
        RECT 4.288 236.574 4.392 240.948 ; 
        RECT 3.856 236.574 3.96 240.948 ; 
        RECT 3.424 236.574 3.528 240.948 ; 
        RECT 2.992 236.574 3.096 240.948 ; 
        RECT 2.56 236.574 2.664 240.948 ; 
        RECT 2.128 236.574 2.232 240.948 ; 
        RECT 1.696 236.574 1.8 240.948 ; 
        RECT 1.264 236.574 1.368 240.948 ; 
        RECT 0.832 236.574 0.936 240.948 ; 
        RECT 0.02 236.574 0.36 240.948 ; 
        RECT 34.564 240.894 35.076 245.268 ; 
        RECT 34.508 243.556 35.076 244.846 ; 
        RECT 33.916 242.464 34.164 245.268 ; 
        RECT 33.86 243.702 34.164 244.316 ; 
        RECT 33.916 240.894 34.02 245.268 ; 
        RECT 33.916 241.378 34.076 242.336 ; 
        RECT 33.916 240.894 34.164 241.25 ; 
        RECT 32.728 242.696 33.552 245.268 ; 
        RECT 33.448 240.894 33.552 245.268 ; 
        RECT 32.728 243.804 33.608 244.836 ; 
        RECT 32.728 240.894 33.12 245.268 ; 
        RECT 31.06 240.894 31.392 245.268 ; 
        RECT 31.06 241.248 31.448 244.99 ; 
        RECT 65.776 240.894 66.116 245.268 ; 
        RECT 65.2 240.894 65.304 245.268 ; 
        RECT 64.768 240.894 64.872 245.268 ; 
        RECT 64.336 240.894 64.44 245.268 ; 
        RECT 63.904 240.894 64.008 245.268 ; 
        RECT 63.472 240.894 63.576 245.268 ; 
        RECT 63.04 240.894 63.144 245.268 ; 
        RECT 62.608 240.894 62.712 245.268 ; 
        RECT 62.176 240.894 62.28 245.268 ; 
        RECT 61.744 240.894 61.848 245.268 ; 
        RECT 61.312 240.894 61.416 245.268 ; 
        RECT 60.88 240.894 60.984 245.268 ; 
        RECT 60.448 240.894 60.552 245.268 ; 
        RECT 60.016 240.894 60.12 245.268 ; 
        RECT 59.584 240.894 59.688 245.268 ; 
        RECT 59.152 240.894 59.256 245.268 ; 
        RECT 58.72 240.894 58.824 245.268 ; 
        RECT 58.288 240.894 58.392 245.268 ; 
        RECT 57.856 240.894 57.96 245.268 ; 
        RECT 57.424 240.894 57.528 245.268 ; 
        RECT 56.992 240.894 57.096 245.268 ; 
        RECT 56.56 240.894 56.664 245.268 ; 
        RECT 56.128 240.894 56.232 245.268 ; 
        RECT 55.696 240.894 55.8 245.268 ; 
        RECT 55.264 240.894 55.368 245.268 ; 
        RECT 54.832 240.894 54.936 245.268 ; 
        RECT 54.4 240.894 54.504 245.268 ; 
        RECT 53.968 240.894 54.072 245.268 ; 
        RECT 53.536 240.894 53.64 245.268 ; 
        RECT 53.104 240.894 53.208 245.268 ; 
        RECT 52.672 240.894 52.776 245.268 ; 
        RECT 52.24 240.894 52.344 245.268 ; 
        RECT 51.808 240.894 51.912 245.268 ; 
        RECT 51.376 240.894 51.48 245.268 ; 
        RECT 50.944 240.894 51.048 245.268 ; 
        RECT 50.512 240.894 50.616 245.268 ; 
        RECT 50.08 240.894 50.184 245.268 ; 
        RECT 49.648 240.894 49.752 245.268 ; 
        RECT 49.216 240.894 49.32 245.268 ; 
        RECT 48.784 240.894 48.888 245.268 ; 
        RECT 48.352 240.894 48.456 245.268 ; 
        RECT 47.92 240.894 48.024 245.268 ; 
        RECT 47.488 240.894 47.592 245.268 ; 
        RECT 47.056 240.894 47.16 245.268 ; 
        RECT 46.624 240.894 46.728 245.268 ; 
        RECT 46.192 240.894 46.296 245.268 ; 
        RECT 45.76 240.894 45.864 245.268 ; 
        RECT 45.328 240.894 45.432 245.268 ; 
        RECT 44.896 240.894 45 245.268 ; 
        RECT 44.464 240.894 44.568 245.268 ; 
        RECT 44.032 240.894 44.136 245.268 ; 
        RECT 43.6 240.894 43.704 245.268 ; 
        RECT 43.168 240.894 43.272 245.268 ; 
        RECT 42.736 240.894 42.84 245.268 ; 
        RECT 42.304 240.894 42.408 245.268 ; 
        RECT 41.872 240.894 41.976 245.268 ; 
        RECT 41.44 240.894 41.544 245.268 ; 
        RECT 41.008 240.894 41.112 245.268 ; 
        RECT 40.576 240.894 40.68 245.268 ; 
        RECT 40.144 240.894 40.248 245.268 ; 
        RECT 39.712 240.894 39.816 245.268 ; 
        RECT 39.28 240.894 39.384 245.268 ; 
        RECT 38.848 240.894 38.952 245.268 ; 
        RECT 38.416 240.894 38.52 245.268 ; 
        RECT 37.984 240.894 38.088 245.268 ; 
        RECT 37.552 240.894 37.656 245.268 ; 
        RECT 36.7 240.894 37.008 245.268 ; 
        RECT 29.128 240.894 29.436 245.268 ; 
        RECT 28.48 240.894 28.584 245.268 ; 
        RECT 28.048 240.894 28.152 245.268 ; 
        RECT 27.616 240.894 27.72 245.268 ; 
        RECT 27.184 240.894 27.288 245.268 ; 
        RECT 26.752 240.894 26.856 245.268 ; 
        RECT 26.32 240.894 26.424 245.268 ; 
        RECT 25.888 240.894 25.992 245.268 ; 
        RECT 25.456 240.894 25.56 245.268 ; 
        RECT 25.024 240.894 25.128 245.268 ; 
        RECT 24.592 240.894 24.696 245.268 ; 
        RECT 24.16 240.894 24.264 245.268 ; 
        RECT 23.728 240.894 23.832 245.268 ; 
        RECT 23.296 240.894 23.4 245.268 ; 
        RECT 22.864 240.894 22.968 245.268 ; 
        RECT 22.432 240.894 22.536 245.268 ; 
        RECT 22 240.894 22.104 245.268 ; 
        RECT 21.568 240.894 21.672 245.268 ; 
        RECT 21.136 240.894 21.24 245.268 ; 
        RECT 20.704 240.894 20.808 245.268 ; 
        RECT 20.272 240.894 20.376 245.268 ; 
        RECT 19.84 240.894 19.944 245.268 ; 
        RECT 19.408 240.894 19.512 245.268 ; 
        RECT 18.976 240.894 19.08 245.268 ; 
        RECT 18.544 240.894 18.648 245.268 ; 
        RECT 18.112 240.894 18.216 245.268 ; 
        RECT 17.68 240.894 17.784 245.268 ; 
        RECT 17.248 240.894 17.352 245.268 ; 
        RECT 16.816 240.894 16.92 245.268 ; 
        RECT 16.384 240.894 16.488 245.268 ; 
        RECT 15.952 240.894 16.056 245.268 ; 
        RECT 15.52 240.894 15.624 245.268 ; 
        RECT 15.088 240.894 15.192 245.268 ; 
        RECT 14.656 240.894 14.76 245.268 ; 
        RECT 14.224 240.894 14.328 245.268 ; 
        RECT 13.792 240.894 13.896 245.268 ; 
        RECT 13.36 240.894 13.464 245.268 ; 
        RECT 12.928 240.894 13.032 245.268 ; 
        RECT 12.496 240.894 12.6 245.268 ; 
        RECT 12.064 240.894 12.168 245.268 ; 
        RECT 11.632 240.894 11.736 245.268 ; 
        RECT 11.2 240.894 11.304 245.268 ; 
        RECT 10.768 240.894 10.872 245.268 ; 
        RECT 10.336 240.894 10.44 245.268 ; 
        RECT 9.904 240.894 10.008 245.268 ; 
        RECT 9.472 240.894 9.576 245.268 ; 
        RECT 9.04 240.894 9.144 245.268 ; 
        RECT 8.608 240.894 8.712 245.268 ; 
        RECT 8.176 240.894 8.28 245.268 ; 
        RECT 7.744 240.894 7.848 245.268 ; 
        RECT 7.312 240.894 7.416 245.268 ; 
        RECT 6.88 240.894 6.984 245.268 ; 
        RECT 6.448 240.894 6.552 245.268 ; 
        RECT 6.016 240.894 6.12 245.268 ; 
        RECT 5.584 240.894 5.688 245.268 ; 
        RECT 5.152 240.894 5.256 245.268 ; 
        RECT 4.72 240.894 4.824 245.268 ; 
        RECT 4.288 240.894 4.392 245.268 ; 
        RECT 3.856 240.894 3.96 245.268 ; 
        RECT 3.424 240.894 3.528 245.268 ; 
        RECT 2.992 240.894 3.096 245.268 ; 
        RECT 2.56 240.894 2.664 245.268 ; 
        RECT 2.128 240.894 2.232 245.268 ; 
        RECT 1.696 240.894 1.8 245.268 ; 
        RECT 1.264 240.894 1.368 245.268 ; 
        RECT 0.832 240.894 0.936 245.268 ; 
        RECT 0.02 240.894 0.36 245.268 ; 
        RECT 34.564 245.214 35.076 249.588 ; 
        RECT 34.508 247.876 35.076 249.166 ; 
        RECT 33.916 246.784 34.164 249.588 ; 
        RECT 33.86 248.022 34.164 248.636 ; 
        RECT 33.916 245.214 34.02 249.588 ; 
        RECT 33.916 245.698 34.076 246.656 ; 
        RECT 33.916 245.214 34.164 245.57 ; 
        RECT 32.728 247.016 33.552 249.588 ; 
        RECT 33.448 245.214 33.552 249.588 ; 
        RECT 32.728 248.124 33.608 249.156 ; 
        RECT 32.728 245.214 33.12 249.588 ; 
        RECT 31.06 245.214 31.392 249.588 ; 
        RECT 31.06 245.568 31.448 249.31 ; 
        RECT 65.776 245.214 66.116 249.588 ; 
        RECT 65.2 245.214 65.304 249.588 ; 
        RECT 64.768 245.214 64.872 249.588 ; 
        RECT 64.336 245.214 64.44 249.588 ; 
        RECT 63.904 245.214 64.008 249.588 ; 
        RECT 63.472 245.214 63.576 249.588 ; 
        RECT 63.04 245.214 63.144 249.588 ; 
        RECT 62.608 245.214 62.712 249.588 ; 
        RECT 62.176 245.214 62.28 249.588 ; 
        RECT 61.744 245.214 61.848 249.588 ; 
        RECT 61.312 245.214 61.416 249.588 ; 
        RECT 60.88 245.214 60.984 249.588 ; 
        RECT 60.448 245.214 60.552 249.588 ; 
        RECT 60.016 245.214 60.12 249.588 ; 
        RECT 59.584 245.214 59.688 249.588 ; 
        RECT 59.152 245.214 59.256 249.588 ; 
        RECT 58.72 245.214 58.824 249.588 ; 
        RECT 58.288 245.214 58.392 249.588 ; 
        RECT 57.856 245.214 57.96 249.588 ; 
        RECT 57.424 245.214 57.528 249.588 ; 
        RECT 56.992 245.214 57.096 249.588 ; 
        RECT 56.56 245.214 56.664 249.588 ; 
        RECT 56.128 245.214 56.232 249.588 ; 
        RECT 55.696 245.214 55.8 249.588 ; 
        RECT 55.264 245.214 55.368 249.588 ; 
        RECT 54.832 245.214 54.936 249.588 ; 
        RECT 54.4 245.214 54.504 249.588 ; 
        RECT 53.968 245.214 54.072 249.588 ; 
        RECT 53.536 245.214 53.64 249.588 ; 
        RECT 53.104 245.214 53.208 249.588 ; 
        RECT 52.672 245.214 52.776 249.588 ; 
        RECT 52.24 245.214 52.344 249.588 ; 
        RECT 51.808 245.214 51.912 249.588 ; 
        RECT 51.376 245.214 51.48 249.588 ; 
        RECT 50.944 245.214 51.048 249.588 ; 
        RECT 50.512 245.214 50.616 249.588 ; 
        RECT 50.08 245.214 50.184 249.588 ; 
        RECT 49.648 245.214 49.752 249.588 ; 
        RECT 49.216 245.214 49.32 249.588 ; 
        RECT 48.784 245.214 48.888 249.588 ; 
        RECT 48.352 245.214 48.456 249.588 ; 
        RECT 47.92 245.214 48.024 249.588 ; 
        RECT 47.488 245.214 47.592 249.588 ; 
        RECT 47.056 245.214 47.16 249.588 ; 
        RECT 46.624 245.214 46.728 249.588 ; 
        RECT 46.192 245.214 46.296 249.588 ; 
        RECT 45.76 245.214 45.864 249.588 ; 
        RECT 45.328 245.214 45.432 249.588 ; 
        RECT 44.896 245.214 45 249.588 ; 
        RECT 44.464 245.214 44.568 249.588 ; 
        RECT 44.032 245.214 44.136 249.588 ; 
        RECT 43.6 245.214 43.704 249.588 ; 
        RECT 43.168 245.214 43.272 249.588 ; 
        RECT 42.736 245.214 42.84 249.588 ; 
        RECT 42.304 245.214 42.408 249.588 ; 
        RECT 41.872 245.214 41.976 249.588 ; 
        RECT 41.44 245.214 41.544 249.588 ; 
        RECT 41.008 245.214 41.112 249.588 ; 
        RECT 40.576 245.214 40.68 249.588 ; 
        RECT 40.144 245.214 40.248 249.588 ; 
        RECT 39.712 245.214 39.816 249.588 ; 
        RECT 39.28 245.214 39.384 249.588 ; 
        RECT 38.848 245.214 38.952 249.588 ; 
        RECT 38.416 245.214 38.52 249.588 ; 
        RECT 37.984 245.214 38.088 249.588 ; 
        RECT 37.552 245.214 37.656 249.588 ; 
        RECT 36.7 245.214 37.008 249.588 ; 
        RECT 29.128 245.214 29.436 249.588 ; 
        RECT 28.48 245.214 28.584 249.588 ; 
        RECT 28.048 245.214 28.152 249.588 ; 
        RECT 27.616 245.214 27.72 249.588 ; 
        RECT 27.184 245.214 27.288 249.588 ; 
        RECT 26.752 245.214 26.856 249.588 ; 
        RECT 26.32 245.214 26.424 249.588 ; 
        RECT 25.888 245.214 25.992 249.588 ; 
        RECT 25.456 245.214 25.56 249.588 ; 
        RECT 25.024 245.214 25.128 249.588 ; 
        RECT 24.592 245.214 24.696 249.588 ; 
        RECT 24.16 245.214 24.264 249.588 ; 
        RECT 23.728 245.214 23.832 249.588 ; 
        RECT 23.296 245.214 23.4 249.588 ; 
        RECT 22.864 245.214 22.968 249.588 ; 
        RECT 22.432 245.214 22.536 249.588 ; 
        RECT 22 245.214 22.104 249.588 ; 
        RECT 21.568 245.214 21.672 249.588 ; 
        RECT 21.136 245.214 21.24 249.588 ; 
        RECT 20.704 245.214 20.808 249.588 ; 
        RECT 20.272 245.214 20.376 249.588 ; 
        RECT 19.84 245.214 19.944 249.588 ; 
        RECT 19.408 245.214 19.512 249.588 ; 
        RECT 18.976 245.214 19.08 249.588 ; 
        RECT 18.544 245.214 18.648 249.588 ; 
        RECT 18.112 245.214 18.216 249.588 ; 
        RECT 17.68 245.214 17.784 249.588 ; 
        RECT 17.248 245.214 17.352 249.588 ; 
        RECT 16.816 245.214 16.92 249.588 ; 
        RECT 16.384 245.214 16.488 249.588 ; 
        RECT 15.952 245.214 16.056 249.588 ; 
        RECT 15.52 245.214 15.624 249.588 ; 
        RECT 15.088 245.214 15.192 249.588 ; 
        RECT 14.656 245.214 14.76 249.588 ; 
        RECT 14.224 245.214 14.328 249.588 ; 
        RECT 13.792 245.214 13.896 249.588 ; 
        RECT 13.36 245.214 13.464 249.588 ; 
        RECT 12.928 245.214 13.032 249.588 ; 
        RECT 12.496 245.214 12.6 249.588 ; 
        RECT 12.064 245.214 12.168 249.588 ; 
        RECT 11.632 245.214 11.736 249.588 ; 
        RECT 11.2 245.214 11.304 249.588 ; 
        RECT 10.768 245.214 10.872 249.588 ; 
        RECT 10.336 245.214 10.44 249.588 ; 
        RECT 9.904 245.214 10.008 249.588 ; 
        RECT 9.472 245.214 9.576 249.588 ; 
        RECT 9.04 245.214 9.144 249.588 ; 
        RECT 8.608 245.214 8.712 249.588 ; 
        RECT 8.176 245.214 8.28 249.588 ; 
        RECT 7.744 245.214 7.848 249.588 ; 
        RECT 7.312 245.214 7.416 249.588 ; 
        RECT 6.88 245.214 6.984 249.588 ; 
        RECT 6.448 245.214 6.552 249.588 ; 
        RECT 6.016 245.214 6.12 249.588 ; 
        RECT 5.584 245.214 5.688 249.588 ; 
        RECT 5.152 245.214 5.256 249.588 ; 
        RECT 4.72 245.214 4.824 249.588 ; 
        RECT 4.288 245.214 4.392 249.588 ; 
        RECT 3.856 245.214 3.96 249.588 ; 
        RECT 3.424 245.214 3.528 249.588 ; 
        RECT 2.992 245.214 3.096 249.588 ; 
        RECT 2.56 245.214 2.664 249.588 ; 
        RECT 2.128 245.214 2.232 249.588 ; 
        RECT 1.696 245.214 1.8 249.588 ; 
        RECT 1.264 245.214 1.368 249.588 ; 
        RECT 0.832 245.214 0.936 249.588 ; 
        RECT 0.02 245.214 0.36 249.588 ; 
        RECT 34.564 249.534 35.076 253.908 ; 
        RECT 34.508 252.196 35.076 253.486 ; 
        RECT 33.916 251.104 34.164 253.908 ; 
        RECT 33.86 252.342 34.164 252.956 ; 
        RECT 33.916 249.534 34.02 253.908 ; 
        RECT 33.916 250.018 34.076 250.976 ; 
        RECT 33.916 249.534 34.164 249.89 ; 
        RECT 32.728 251.336 33.552 253.908 ; 
        RECT 33.448 249.534 33.552 253.908 ; 
        RECT 32.728 252.444 33.608 253.476 ; 
        RECT 32.728 249.534 33.12 253.908 ; 
        RECT 31.06 249.534 31.392 253.908 ; 
        RECT 31.06 249.888 31.448 253.63 ; 
        RECT 65.776 249.534 66.116 253.908 ; 
        RECT 65.2 249.534 65.304 253.908 ; 
        RECT 64.768 249.534 64.872 253.908 ; 
        RECT 64.336 249.534 64.44 253.908 ; 
        RECT 63.904 249.534 64.008 253.908 ; 
        RECT 63.472 249.534 63.576 253.908 ; 
        RECT 63.04 249.534 63.144 253.908 ; 
        RECT 62.608 249.534 62.712 253.908 ; 
        RECT 62.176 249.534 62.28 253.908 ; 
        RECT 61.744 249.534 61.848 253.908 ; 
        RECT 61.312 249.534 61.416 253.908 ; 
        RECT 60.88 249.534 60.984 253.908 ; 
        RECT 60.448 249.534 60.552 253.908 ; 
        RECT 60.016 249.534 60.12 253.908 ; 
        RECT 59.584 249.534 59.688 253.908 ; 
        RECT 59.152 249.534 59.256 253.908 ; 
        RECT 58.72 249.534 58.824 253.908 ; 
        RECT 58.288 249.534 58.392 253.908 ; 
        RECT 57.856 249.534 57.96 253.908 ; 
        RECT 57.424 249.534 57.528 253.908 ; 
        RECT 56.992 249.534 57.096 253.908 ; 
        RECT 56.56 249.534 56.664 253.908 ; 
        RECT 56.128 249.534 56.232 253.908 ; 
        RECT 55.696 249.534 55.8 253.908 ; 
        RECT 55.264 249.534 55.368 253.908 ; 
        RECT 54.832 249.534 54.936 253.908 ; 
        RECT 54.4 249.534 54.504 253.908 ; 
        RECT 53.968 249.534 54.072 253.908 ; 
        RECT 53.536 249.534 53.64 253.908 ; 
        RECT 53.104 249.534 53.208 253.908 ; 
        RECT 52.672 249.534 52.776 253.908 ; 
        RECT 52.24 249.534 52.344 253.908 ; 
        RECT 51.808 249.534 51.912 253.908 ; 
        RECT 51.376 249.534 51.48 253.908 ; 
        RECT 50.944 249.534 51.048 253.908 ; 
        RECT 50.512 249.534 50.616 253.908 ; 
        RECT 50.08 249.534 50.184 253.908 ; 
        RECT 49.648 249.534 49.752 253.908 ; 
        RECT 49.216 249.534 49.32 253.908 ; 
        RECT 48.784 249.534 48.888 253.908 ; 
        RECT 48.352 249.534 48.456 253.908 ; 
        RECT 47.92 249.534 48.024 253.908 ; 
        RECT 47.488 249.534 47.592 253.908 ; 
        RECT 47.056 249.534 47.16 253.908 ; 
        RECT 46.624 249.534 46.728 253.908 ; 
        RECT 46.192 249.534 46.296 253.908 ; 
        RECT 45.76 249.534 45.864 253.908 ; 
        RECT 45.328 249.534 45.432 253.908 ; 
        RECT 44.896 249.534 45 253.908 ; 
        RECT 44.464 249.534 44.568 253.908 ; 
        RECT 44.032 249.534 44.136 253.908 ; 
        RECT 43.6 249.534 43.704 253.908 ; 
        RECT 43.168 249.534 43.272 253.908 ; 
        RECT 42.736 249.534 42.84 253.908 ; 
        RECT 42.304 249.534 42.408 253.908 ; 
        RECT 41.872 249.534 41.976 253.908 ; 
        RECT 41.44 249.534 41.544 253.908 ; 
        RECT 41.008 249.534 41.112 253.908 ; 
        RECT 40.576 249.534 40.68 253.908 ; 
        RECT 40.144 249.534 40.248 253.908 ; 
        RECT 39.712 249.534 39.816 253.908 ; 
        RECT 39.28 249.534 39.384 253.908 ; 
        RECT 38.848 249.534 38.952 253.908 ; 
        RECT 38.416 249.534 38.52 253.908 ; 
        RECT 37.984 249.534 38.088 253.908 ; 
        RECT 37.552 249.534 37.656 253.908 ; 
        RECT 36.7 249.534 37.008 253.908 ; 
        RECT 29.128 249.534 29.436 253.908 ; 
        RECT 28.48 249.534 28.584 253.908 ; 
        RECT 28.048 249.534 28.152 253.908 ; 
        RECT 27.616 249.534 27.72 253.908 ; 
        RECT 27.184 249.534 27.288 253.908 ; 
        RECT 26.752 249.534 26.856 253.908 ; 
        RECT 26.32 249.534 26.424 253.908 ; 
        RECT 25.888 249.534 25.992 253.908 ; 
        RECT 25.456 249.534 25.56 253.908 ; 
        RECT 25.024 249.534 25.128 253.908 ; 
        RECT 24.592 249.534 24.696 253.908 ; 
        RECT 24.16 249.534 24.264 253.908 ; 
        RECT 23.728 249.534 23.832 253.908 ; 
        RECT 23.296 249.534 23.4 253.908 ; 
        RECT 22.864 249.534 22.968 253.908 ; 
        RECT 22.432 249.534 22.536 253.908 ; 
        RECT 22 249.534 22.104 253.908 ; 
        RECT 21.568 249.534 21.672 253.908 ; 
        RECT 21.136 249.534 21.24 253.908 ; 
        RECT 20.704 249.534 20.808 253.908 ; 
        RECT 20.272 249.534 20.376 253.908 ; 
        RECT 19.84 249.534 19.944 253.908 ; 
        RECT 19.408 249.534 19.512 253.908 ; 
        RECT 18.976 249.534 19.08 253.908 ; 
        RECT 18.544 249.534 18.648 253.908 ; 
        RECT 18.112 249.534 18.216 253.908 ; 
        RECT 17.68 249.534 17.784 253.908 ; 
        RECT 17.248 249.534 17.352 253.908 ; 
        RECT 16.816 249.534 16.92 253.908 ; 
        RECT 16.384 249.534 16.488 253.908 ; 
        RECT 15.952 249.534 16.056 253.908 ; 
        RECT 15.52 249.534 15.624 253.908 ; 
        RECT 15.088 249.534 15.192 253.908 ; 
        RECT 14.656 249.534 14.76 253.908 ; 
        RECT 14.224 249.534 14.328 253.908 ; 
        RECT 13.792 249.534 13.896 253.908 ; 
        RECT 13.36 249.534 13.464 253.908 ; 
        RECT 12.928 249.534 13.032 253.908 ; 
        RECT 12.496 249.534 12.6 253.908 ; 
        RECT 12.064 249.534 12.168 253.908 ; 
        RECT 11.632 249.534 11.736 253.908 ; 
        RECT 11.2 249.534 11.304 253.908 ; 
        RECT 10.768 249.534 10.872 253.908 ; 
        RECT 10.336 249.534 10.44 253.908 ; 
        RECT 9.904 249.534 10.008 253.908 ; 
        RECT 9.472 249.534 9.576 253.908 ; 
        RECT 9.04 249.534 9.144 253.908 ; 
        RECT 8.608 249.534 8.712 253.908 ; 
        RECT 8.176 249.534 8.28 253.908 ; 
        RECT 7.744 249.534 7.848 253.908 ; 
        RECT 7.312 249.534 7.416 253.908 ; 
        RECT 6.88 249.534 6.984 253.908 ; 
        RECT 6.448 249.534 6.552 253.908 ; 
        RECT 6.016 249.534 6.12 253.908 ; 
        RECT 5.584 249.534 5.688 253.908 ; 
        RECT 5.152 249.534 5.256 253.908 ; 
        RECT 4.72 249.534 4.824 253.908 ; 
        RECT 4.288 249.534 4.392 253.908 ; 
        RECT 3.856 249.534 3.96 253.908 ; 
        RECT 3.424 249.534 3.528 253.908 ; 
        RECT 2.992 249.534 3.096 253.908 ; 
        RECT 2.56 249.534 2.664 253.908 ; 
        RECT 2.128 249.534 2.232 253.908 ; 
        RECT 1.696 249.534 1.8 253.908 ; 
        RECT 1.264 249.534 1.368 253.908 ; 
        RECT 0.832 249.534 0.936 253.908 ; 
        RECT 0.02 249.534 0.36 253.908 ; 
        RECT 34.564 253.854 35.076 258.228 ; 
        RECT 34.508 256.516 35.076 257.806 ; 
        RECT 33.916 255.424 34.164 258.228 ; 
        RECT 33.86 256.662 34.164 257.276 ; 
        RECT 33.916 253.854 34.02 258.228 ; 
        RECT 33.916 254.338 34.076 255.296 ; 
        RECT 33.916 253.854 34.164 254.21 ; 
        RECT 32.728 255.656 33.552 258.228 ; 
        RECT 33.448 253.854 33.552 258.228 ; 
        RECT 32.728 256.764 33.608 257.796 ; 
        RECT 32.728 253.854 33.12 258.228 ; 
        RECT 31.06 253.854 31.392 258.228 ; 
        RECT 31.06 254.208 31.448 257.95 ; 
        RECT 65.776 253.854 66.116 258.228 ; 
        RECT 65.2 253.854 65.304 258.228 ; 
        RECT 64.768 253.854 64.872 258.228 ; 
        RECT 64.336 253.854 64.44 258.228 ; 
        RECT 63.904 253.854 64.008 258.228 ; 
        RECT 63.472 253.854 63.576 258.228 ; 
        RECT 63.04 253.854 63.144 258.228 ; 
        RECT 62.608 253.854 62.712 258.228 ; 
        RECT 62.176 253.854 62.28 258.228 ; 
        RECT 61.744 253.854 61.848 258.228 ; 
        RECT 61.312 253.854 61.416 258.228 ; 
        RECT 60.88 253.854 60.984 258.228 ; 
        RECT 60.448 253.854 60.552 258.228 ; 
        RECT 60.016 253.854 60.12 258.228 ; 
        RECT 59.584 253.854 59.688 258.228 ; 
        RECT 59.152 253.854 59.256 258.228 ; 
        RECT 58.72 253.854 58.824 258.228 ; 
        RECT 58.288 253.854 58.392 258.228 ; 
        RECT 57.856 253.854 57.96 258.228 ; 
        RECT 57.424 253.854 57.528 258.228 ; 
        RECT 56.992 253.854 57.096 258.228 ; 
        RECT 56.56 253.854 56.664 258.228 ; 
        RECT 56.128 253.854 56.232 258.228 ; 
        RECT 55.696 253.854 55.8 258.228 ; 
        RECT 55.264 253.854 55.368 258.228 ; 
        RECT 54.832 253.854 54.936 258.228 ; 
        RECT 54.4 253.854 54.504 258.228 ; 
        RECT 53.968 253.854 54.072 258.228 ; 
        RECT 53.536 253.854 53.64 258.228 ; 
        RECT 53.104 253.854 53.208 258.228 ; 
        RECT 52.672 253.854 52.776 258.228 ; 
        RECT 52.24 253.854 52.344 258.228 ; 
        RECT 51.808 253.854 51.912 258.228 ; 
        RECT 51.376 253.854 51.48 258.228 ; 
        RECT 50.944 253.854 51.048 258.228 ; 
        RECT 50.512 253.854 50.616 258.228 ; 
        RECT 50.08 253.854 50.184 258.228 ; 
        RECT 49.648 253.854 49.752 258.228 ; 
        RECT 49.216 253.854 49.32 258.228 ; 
        RECT 48.784 253.854 48.888 258.228 ; 
        RECT 48.352 253.854 48.456 258.228 ; 
        RECT 47.92 253.854 48.024 258.228 ; 
        RECT 47.488 253.854 47.592 258.228 ; 
        RECT 47.056 253.854 47.16 258.228 ; 
        RECT 46.624 253.854 46.728 258.228 ; 
        RECT 46.192 253.854 46.296 258.228 ; 
        RECT 45.76 253.854 45.864 258.228 ; 
        RECT 45.328 253.854 45.432 258.228 ; 
        RECT 44.896 253.854 45 258.228 ; 
        RECT 44.464 253.854 44.568 258.228 ; 
        RECT 44.032 253.854 44.136 258.228 ; 
        RECT 43.6 253.854 43.704 258.228 ; 
        RECT 43.168 253.854 43.272 258.228 ; 
        RECT 42.736 253.854 42.84 258.228 ; 
        RECT 42.304 253.854 42.408 258.228 ; 
        RECT 41.872 253.854 41.976 258.228 ; 
        RECT 41.44 253.854 41.544 258.228 ; 
        RECT 41.008 253.854 41.112 258.228 ; 
        RECT 40.576 253.854 40.68 258.228 ; 
        RECT 40.144 253.854 40.248 258.228 ; 
        RECT 39.712 253.854 39.816 258.228 ; 
        RECT 39.28 253.854 39.384 258.228 ; 
        RECT 38.848 253.854 38.952 258.228 ; 
        RECT 38.416 253.854 38.52 258.228 ; 
        RECT 37.984 253.854 38.088 258.228 ; 
        RECT 37.552 253.854 37.656 258.228 ; 
        RECT 36.7 253.854 37.008 258.228 ; 
        RECT 29.128 253.854 29.436 258.228 ; 
        RECT 28.48 253.854 28.584 258.228 ; 
        RECT 28.048 253.854 28.152 258.228 ; 
        RECT 27.616 253.854 27.72 258.228 ; 
        RECT 27.184 253.854 27.288 258.228 ; 
        RECT 26.752 253.854 26.856 258.228 ; 
        RECT 26.32 253.854 26.424 258.228 ; 
        RECT 25.888 253.854 25.992 258.228 ; 
        RECT 25.456 253.854 25.56 258.228 ; 
        RECT 25.024 253.854 25.128 258.228 ; 
        RECT 24.592 253.854 24.696 258.228 ; 
        RECT 24.16 253.854 24.264 258.228 ; 
        RECT 23.728 253.854 23.832 258.228 ; 
        RECT 23.296 253.854 23.4 258.228 ; 
        RECT 22.864 253.854 22.968 258.228 ; 
        RECT 22.432 253.854 22.536 258.228 ; 
        RECT 22 253.854 22.104 258.228 ; 
        RECT 21.568 253.854 21.672 258.228 ; 
        RECT 21.136 253.854 21.24 258.228 ; 
        RECT 20.704 253.854 20.808 258.228 ; 
        RECT 20.272 253.854 20.376 258.228 ; 
        RECT 19.84 253.854 19.944 258.228 ; 
        RECT 19.408 253.854 19.512 258.228 ; 
        RECT 18.976 253.854 19.08 258.228 ; 
        RECT 18.544 253.854 18.648 258.228 ; 
        RECT 18.112 253.854 18.216 258.228 ; 
        RECT 17.68 253.854 17.784 258.228 ; 
        RECT 17.248 253.854 17.352 258.228 ; 
        RECT 16.816 253.854 16.92 258.228 ; 
        RECT 16.384 253.854 16.488 258.228 ; 
        RECT 15.952 253.854 16.056 258.228 ; 
        RECT 15.52 253.854 15.624 258.228 ; 
        RECT 15.088 253.854 15.192 258.228 ; 
        RECT 14.656 253.854 14.76 258.228 ; 
        RECT 14.224 253.854 14.328 258.228 ; 
        RECT 13.792 253.854 13.896 258.228 ; 
        RECT 13.36 253.854 13.464 258.228 ; 
        RECT 12.928 253.854 13.032 258.228 ; 
        RECT 12.496 253.854 12.6 258.228 ; 
        RECT 12.064 253.854 12.168 258.228 ; 
        RECT 11.632 253.854 11.736 258.228 ; 
        RECT 11.2 253.854 11.304 258.228 ; 
        RECT 10.768 253.854 10.872 258.228 ; 
        RECT 10.336 253.854 10.44 258.228 ; 
        RECT 9.904 253.854 10.008 258.228 ; 
        RECT 9.472 253.854 9.576 258.228 ; 
        RECT 9.04 253.854 9.144 258.228 ; 
        RECT 8.608 253.854 8.712 258.228 ; 
        RECT 8.176 253.854 8.28 258.228 ; 
        RECT 7.744 253.854 7.848 258.228 ; 
        RECT 7.312 253.854 7.416 258.228 ; 
        RECT 6.88 253.854 6.984 258.228 ; 
        RECT 6.448 253.854 6.552 258.228 ; 
        RECT 6.016 253.854 6.12 258.228 ; 
        RECT 5.584 253.854 5.688 258.228 ; 
        RECT 5.152 253.854 5.256 258.228 ; 
        RECT 4.72 253.854 4.824 258.228 ; 
        RECT 4.288 253.854 4.392 258.228 ; 
        RECT 3.856 253.854 3.96 258.228 ; 
        RECT 3.424 253.854 3.528 258.228 ; 
        RECT 2.992 253.854 3.096 258.228 ; 
        RECT 2.56 253.854 2.664 258.228 ; 
        RECT 2.128 253.854 2.232 258.228 ; 
        RECT 1.696 253.854 1.8 258.228 ; 
        RECT 1.264 253.854 1.368 258.228 ; 
        RECT 0.832 253.854 0.936 258.228 ; 
        RECT 0.02 253.854 0.36 258.228 ; 
        RECT 34.564 258.174 35.076 262.548 ; 
        RECT 34.508 260.836 35.076 262.126 ; 
        RECT 33.916 259.744 34.164 262.548 ; 
        RECT 33.86 260.982 34.164 261.596 ; 
        RECT 33.916 258.174 34.02 262.548 ; 
        RECT 33.916 258.658 34.076 259.616 ; 
        RECT 33.916 258.174 34.164 258.53 ; 
        RECT 32.728 259.976 33.552 262.548 ; 
        RECT 33.448 258.174 33.552 262.548 ; 
        RECT 32.728 261.084 33.608 262.116 ; 
        RECT 32.728 258.174 33.12 262.548 ; 
        RECT 31.06 258.174 31.392 262.548 ; 
        RECT 31.06 258.528 31.448 262.27 ; 
        RECT 65.776 258.174 66.116 262.548 ; 
        RECT 65.2 258.174 65.304 262.548 ; 
        RECT 64.768 258.174 64.872 262.548 ; 
        RECT 64.336 258.174 64.44 262.548 ; 
        RECT 63.904 258.174 64.008 262.548 ; 
        RECT 63.472 258.174 63.576 262.548 ; 
        RECT 63.04 258.174 63.144 262.548 ; 
        RECT 62.608 258.174 62.712 262.548 ; 
        RECT 62.176 258.174 62.28 262.548 ; 
        RECT 61.744 258.174 61.848 262.548 ; 
        RECT 61.312 258.174 61.416 262.548 ; 
        RECT 60.88 258.174 60.984 262.548 ; 
        RECT 60.448 258.174 60.552 262.548 ; 
        RECT 60.016 258.174 60.12 262.548 ; 
        RECT 59.584 258.174 59.688 262.548 ; 
        RECT 59.152 258.174 59.256 262.548 ; 
        RECT 58.72 258.174 58.824 262.548 ; 
        RECT 58.288 258.174 58.392 262.548 ; 
        RECT 57.856 258.174 57.96 262.548 ; 
        RECT 57.424 258.174 57.528 262.548 ; 
        RECT 56.992 258.174 57.096 262.548 ; 
        RECT 56.56 258.174 56.664 262.548 ; 
        RECT 56.128 258.174 56.232 262.548 ; 
        RECT 55.696 258.174 55.8 262.548 ; 
        RECT 55.264 258.174 55.368 262.548 ; 
        RECT 54.832 258.174 54.936 262.548 ; 
        RECT 54.4 258.174 54.504 262.548 ; 
        RECT 53.968 258.174 54.072 262.548 ; 
        RECT 53.536 258.174 53.64 262.548 ; 
        RECT 53.104 258.174 53.208 262.548 ; 
        RECT 52.672 258.174 52.776 262.548 ; 
        RECT 52.24 258.174 52.344 262.548 ; 
        RECT 51.808 258.174 51.912 262.548 ; 
        RECT 51.376 258.174 51.48 262.548 ; 
        RECT 50.944 258.174 51.048 262.548 ; 
        RECT 50.512 258.174 50.616 262.548 ; 
        RECT 50.08 258.174 50.184 262.548 ; 
        RECT 49.648 258.174 49.752 262.548 ; 
        RECT 49.216 258.174 49.32 262.548 ; 
        RECT 48.784 258.174 48.888 262.548 ; 
        RECT 48.352 258.174 48.456 262.548 ; 
        RECT 47.92 258.174 48.024 262.548 ; 
        RECT 47.488 258.174 47.592 262.548 ; 
        RECT 47.056 258.174 47.16 262.548 ; 
        RECT 46.624 258.174 46.728 262.548 ; 
        RECT 46.192 258.174 46.296 262.548 ; 
        RECT 45.76 258.174 45.864 262.548 ; 
        RECT 45.328 258.174 45.432 262.548 ; 
        RECT 44.896 258.174 45 262.548 ; 
        RECT 44.464 258.174 44.568 262.548 ; 
        RECT 44.032 258.174 44.136 262.548 ; 
        RECT 43.6 258.174 43.704 262.548 ; 
        RECT 43.168 258.174 43.272 262.548 ; 
        RECT 42.736 258.174 42.84 262.548 ; 
        RECT 42.304 258.174 42.408 262.548 ; 
        RECT 41.872 258.174 41.976 262.548 ; 
        RECT 41.44 258.174 41.544 262.548 ; 
        RECT 41.008 258.174 41.112 262.548 ; 
        RECT 40.576 258.174 40.68 262.548 ; 
        RECT 40.144 258.174 40.248 262.548 ; 
        RECT 39.712 258.174 39.816 262.548 ; 
        RECT 39.28 258.174 39.384 262.548 ; 
        RECT 38.848 258.174 38.952 262.548 ; 
        RECT 38.416 258.174 38.52 262.548 ; 
        RECT 37.984 258.174 38.088 262.548 ; 
        RECT 37.552 258.174 37.656 262.548 ; 
        RECT 36.7 258.174 37.008 262.548 ; 
        RECT 29.128 258.174 29.436 262.548 ; 
        RECT 28.48 258.174 28.584 262.548 ; 
        RECT 28.048 258.174 28.152 262.548 ; 
        RECT 27.616 258.174 27.72 262.548 ; 
        RECT 27.184 258.174 27.288 262.548 ; 
        RECT 26.752 258.174 26.856 262.548 ; 
        RECT 26.32 258.174 26.424 262.548 ; 
        RECT 25.888 258.174 25.992 262.548 ; 
        RECT 25.456 258.174 25.56 262.548 ; 
        RECT 25.024 258.174 25.128 262.548 ; 
        RECT 24.592 258.174 24.696 262.548 ; 
        RECT 24.16 258.174 24.264 262.548 ; 
        RECT 23.728 258.174 23.832 262.548 ; 
        RECT 23.296 258.174 23.4 262.548 ; 
        RECT 22.864 258.174 22.968 262.548 ; 
        RECT 22.432 258.174 22.536 262.548 ; 
        RECT 22 258.174 22.104 262.548 ; 
        RECT 21.568 258.174 21.672 262.548 ; 
        RECT 21.136 258.174 21.24 262.548 ; 
        RECT 20.704 258.174 20.808 262.548 ; 
        RECT 20.272 258.174 20.376 262.548 ; 
        RECT 19.84 258.174 19.944 262.548 ; 
        RECT 19.408 258.174 19.512 262.548 ; 
        RECT 18.976 258.174 19.08 262.548 ; 
        RECT 18.544 258.174 18.648 262.548 ; 
        RECT 18.112 258.174 18.216 262.548 ; 
        RECT 17.68 258.174 17.784 262.548 ; 
        RECT 17.248 258.174 17.352 262.548 ; 
        RECT 16.816 258.174 16.92 262.548 ; 
        RECT 16.384 258.174 16.488 262.548 ; 
        RECT 15.952 258.174 16.056 262.548 ; 
        RECT 15.52 258.174 15.624 262.548 ; 
        RECT 15.088 258.174 15.192 262.548 ; 
        RECT 14.656 258.174 14.76 262.548 ; 
        RECT 14.224 258.174 14.328 262.548 ; 
        RECT 13.792 258.174 13.896 262.548 ; 
        RECT 13.36 258.174 13.464 262.548 ; 
        RECT 12.928 258.174 13.032 262.548 ; 
        RECT 12.496 258.174 12.6 262.548 ; 
        RECT 12.064 258.174 12.168 262.548 ; 
        RECT 11.632 258.174 11.736 262.548 ; 
        RECT 11.2 258.174 11.304 262.548 ; 
        RECT 10.768 258.174 10.872 262.548 ; 
        RECT 10.336 258.174 10.44 262.548 ; 
        RECT 9.904 258.174 10.008 262.548 ; 
        RECT 9.472 258.174 9.576 262.548 ; 
        RECT 9.04 258.174 9.144 262.548 ; 
        RECT 8.608 258.174 8.712 262.548 ; 
        RECT 8.176 258.174 8.28 262.548 ; 
        RECT 7.744 258.174 7.848 262.548 ; 
        RECT 7.312 258.174 7.416 262.548 ; 
        RECT 6.88 258.174 6.984 262.548 ; 
        RECT 6.448 258.174 6.552 262.548 ; 
        RECT 6.016 258.174 6.12 262.548 ; 
        RECT 5.584 258.174 5.688 262.548 ; 
        RECT 5.152 258.174 5.256 262.548 ; 
        RECT 4.72 258.174 4.824 262.548 ; 
        RECT 4.288 258.174 4.392 262.548 ; 
        RECT 3.856 258.174 3.96 262.548 ; 
        RECT 3.424 258.174 3.528 262.548 ; 
        RECT 2.992 258.174 3.096 262.548 ; 
        RECT 2.56 258.174 2.664 262.548 ; 
        RECT 2.128 258.174 2.232 262.548 ; 
        RECT 1.696 258.174 1.8 262.548 ; 
        RECT 1.264 258.174 1.368 262.548 ; 
        RECT 0.832 258.174 0.936 262.548 ; 
        RECT 0.02 258.174 0.36 262.548 ; 
        RECT 34.564 262.494 35.076 266.868 ; 
        RECT 34.508 265.156 35.076 266.446 ; 
        RECT 33.916 264.064 34.164 266.868 ; 
        RECT 33.86 265.302 34.164 265.916 ; 
        RECT 33.916 262.494 34.02 266.868 ; 
        RECT 33.916 262.978 34.076 263.936 ; 
        RECT 33.916 262.494 34.164 262.85 ; 
        RECT 32.728 264.296 33.552 266.868 ; 
        RECT 33.448 262.494 33.552 266.868 ; 
        RECT 32.728 265.404 33.608 266.436 ; 
        RECT 32.728 262.494 33.12 266.868 ; 
        RECT 31.06 262.494 31.392 266.868 ; 
        RECT 31.06 262.848 31.448 266.59 ; 
        RECT 65.776 262.494 66.116 266.868 ; 
        RECT 65.2 262.494 65.304 266.868 ; 
        RECT 64.768 262.494 64.872 266.868 ; 
        RECT 64.336 262.494 64.44 266.868 ; 
        RECT 63.904 262.494 64.008 266.868 ; 
        RECT 63.472 262.494 63.576 266.868 ; 
        RECT 63.04 262.494 63.144 266.868 ; 
        RECT 62.608 262.494 62.712 266.868 ; 
        RECT 62.176 262.494 62.28 266.868 ; 
        RECT 61.744 262.494 61.848 266.868 ; 
        RECT 61.312 262.494 61.416 266.868 ; 
        RECT 60.88 262.494 60.984 266.868 ; 
        RECT 60.448 262.494 60.552 266.868 ; 
        RECT 60.016 262.494 60.12 266.868 ; 
        RECT 59.584 262.494 59.688 266.868 ; 
        RECT 59.152 262.494 59.256 266.868 ; 
        RECT 58.72 262.494 58.824 266.868 ; 
        RECT 58.288 262.494 58.392 266.868 ; 
        RECT 57.856 262.494 57.96 266.868 ; 
        RECT 57.424 262.494 57.528 266.868 ; 
        RECT 56.992 262.494 57.096 266.868 ; 
        RECT 56.56 262.494 56.664 266.868 ; 
        RECT 56.128 262.494 56.232 266.868 ; 
        RECT 55.696 262.494 55.8 266.868 ; 
        RECT 55.264 262.494 55.368 266.868 ; 
        RECT 54.832 262.494 54.936 266.868 ; 
        RECT 54.4 262.494 54.504 266.868 ; 
        RECT 53.968 262.494 54.072 266.868 ; 
        RECT 53.536 262.494 53.64 266.868 ; 
        RECT 53.104 262.494 53.208 266.868 ; 
        RECT 52.672 262.494 52.776 266.868 ; 
        RECT 52.24 262.494 52.344 266.868 ; 
        RECT 51.808 262.494 51.912 266.868 ; 
        RECT 51.376 262.494 51.48 266.868 ; 
        RECT 50.944 262.494 51.048 266.868 ; 
        RECT 50.512 262.494 50.616 266.868 ; 
        RECT 50.08 262.494 50.184 266.868 ; 
        RECT 49.648 262.494 49.752 266.868 ; 
        RECT 49.216 262.494 49.32 266.868 ; 
        RECT 48.784 262.494 48.888 266.868 ; 
        RECT 48.352 262.494 48.456 266.868 ; 
        RECT 47.92 262.494 48.024 266.868 ; 
        RECT 47.488 262.494 47.592 266.868 ; 
        RECT 47.056 262.494 47.16 266.868 ; 
        RECT 46.624 262.494 46.728 266.868 ; 
        RECT 46.192 262.494 46.296 266.868 ; 
        RECT 45.76 262.494 45.864 266.868 ; 
        RECT 45.328 262.494 45.432 266.868 ; 
        RECT 44.896 262.494 45 266.868 ; 
        RECT 44.464 262.494 44.568 266.868 ; 
        RECT 44.032 262.494 44.136 266.868 ; 
        RECT 43.6 262.494 43.704 266.868 ; 
        RECT 43.168 262.494 43.272 266.868 ; 
        RECT 42.736 262.494 42.84 266.868 ; 
        RECT 42.304 262.494 42.408 266.868 ; 
        RECT 41.872 262.494 41.976 266.868 ; 
        RECT 41.44 262.494 41.544 266.868 ; 
        RECT 41.008 262.494 41.112 266.868 ; 
        RECT 40.576 262.494 40.68 266.868 ; 
        RECT 40.144 262.494 40.248 266.868 ; 
        RECT 39.712 262.494 39.816 266.868 ; 
        RECT 39.28 262.494 39.384 266.868 ; 
        RECT 38.848 262.494 38.952 266.868 ; 
        RECT 38.416 262.494 38.52 266.868 ; 
        RECT 37.984 262.494 38.088 266.868 ; 
        RECT 37.552 262.494 37.656 266.868 ; 
        RECT 36.7 262.494 37.008 266.868 ; 
        RECT 29.128 262.494 29.436 266.868 ; 
        RECT 28.48 262.494 28.584 266.868 ; 
        RECT 28.048 262.494 28.152 266.868 ; 
        RECT 27.616 262.494 27.72 266.868 ; 
        RECT 27.184 262.494 27.288 266.868 ; 
        RECT 26.752 262.494 26.856 266.868 ; 
        RECT 26.32 262.494 26.424 266.868 ; 
        RECT 25.888 262.494 25.992 266.868 ; 
        RECT 25.456 262.494 25.56 266.868 ; 
        RECT 25.024 262.494 25.128 266.868 ; 
        RECT 24.592 262.494 24.696 266.868 ; 
        RECT 24.16 262.494 24.264 266.868 ; 
        RECT 23.728 262.494 23.832 266.868 ; 
        RECT 23.296 262.494 23.4 266.868 ; 
        RECT 22.864 262.494 22.968 266.868 ; 
        RECT 22.432 262.494 22.536 266.868 ; 
        RECT 22 262.494 22.104 266.868 ; 
        RECT 21.568 262.494 21.672 266.868 ; 
        RECT 21.136 262.494 21.24 266.868 ; 
        RECT 20.704 262.494 20.808 266.868 ; 
        RECT 20.272 262.494 20.376 266.868 ; 
        RECT 19.84 262.494 19.944 266.868 ; 
        RECT 19.408 262.494 19.512 266.868 ; 
        RECT 18.976 262.494 19.08 266.868 ; 
        RECT 18.544 262.494 18.648 266.868 ; 
        RECT 18.112 262.494 18.216 266.868 ; 
        RECT 17.68 262.494 17.784 266.868 ; 
        RECT 17.248 262.494 17.352 266.868 ; 
        RECT 16.816 262.494 16.92 266.868 ; 
        RECT 16.384 262.494 16.488 266.868 ; 
        RECT 15.952 262.494 16.056 266.868 ; 
        RECT 15.52 262.494 15.624 266.868 ; 
        RECT 15.088 262.494 15.192 266.868 ; 
        RECT 14.656 262.494 14.76 266.868 ; 
        RECT 14.224 262.494 14.328 266.868 ; 
        RECT 13.792 262.494 13.896 266.868 ; 
        RECT 13.36 262.494 13.464 266.868 ; 
        RECT 12.928 262.494 13.032 266.868 ; 
        RECT 12.496 262.494 12.6 266.868 ; 
        RECT 12.064 262.494 12.168 266.868 ; 
        RECT 11.632 262.494 11.736 266.868 ; 
        RECT 11.2 262.494 11.304 266.868 ; 
        RECT 10.768 262.494 10.872 266.868 ; 
        RECT 10.336 262.494 10.44 266.868 ; 
        RECT 9.904 262.494 10.008 266.868 ; 
        RECT 9.472 262.494 9.576 266.868 ; 
        RECT 9.04 262.494 9.144 266.868 ; 
        RECT 8.608 262.494 8.712 266.868 ; 
        RECT 8.176 262.494 8.28 266.868 ; 
        RECT 7.744 262.494 7.848 266.868 ; 
        RECT 7.312 262.494 7.416 266.868 ; 
        RECT 6.88 262.494 6.984 266.868 ; 
        RECT 6.448 262.494 6.552 266.868 ; 
        RECT 6.016 262.494 6.12 266.868 ; 
        RECT 5.584 262.494 5.688 266.868 ; 
        RECT 5.152 262.494 5.256 266.868 ; 
        RECT 4.72 262.494 4.824 266.868 ; 
        RECT 4.288 262.494 4.392 266.868 ; 
        RECT 3.856 262.494 3.96 266.868 ; 
        RECT 3.424 262.494 3.528 266.868 ; 
        RECT 2.992 262.494 3.096 266.868 ; 
        RECT 2.56 262.494 2.664 266.868 ; 
        RECT 2.128 262.494 2.232 266.868 ; 
        RECT 1.696 262.494 1.8 266.868 ; 
        RECT 1.264 262.494 1.368 266.868 ; 
        RECT 0.832 262.494 0.936 266.868 ; 
        RECT 0.02 262.494 0.36 266.868 ; 
        RECT 34.564 266.814 35.076 271.188 ; 
        RECT 34.508 269.476 35.076 270.766 ; 
        RECT 33.916 268.384 34.164 271.188 ; 
        RECT 33.86 269.622 34.164 270.236 ; 
        RECT 33.916 266.814 34.02 271.188 ; 
        RECT 33.916 267.298 34.076 268.256 ; 
        RECT 33.916 266.814 34.164 267.17 ; 
        RECT 32.728 268.616 33.552 271.188 ; 
        RECT 33.448 266.814 33.552 271.188 ; 
        RECT 32.728 269.724 33.608 270.756 ; 
        RECT 32.728 266.814 33.12 271.188 ; 
        RECT 31.06 266.814 31.392 271.188 ; 
        RECT 31.06 267.168 31.448 270.91 ; 
        RECT 65.776 266.814 66.116 271.188 ; 
        RECT 65.2 266.814 65.304 271.188 ; 
        RECT 64.768 266.814 64.872 271.188 ; 
        RECT 64.336 266.814 64.44 271.188 ; 
        RECT 63.904 266.814 64.008 271.188 ; 
        RECT 63.472 266.814 63.576 271.188 ; 
        RECT 63.04 266.814 63.144 271.188 ; 
        RECT 62.608 266.814 62.712 271.188 ; 
        RECT 62.176 266.814 62.28 271.188 ; 
        RECT 61.744 266.814 61.848 271.188 ; 
        RECT 61.312 266.814 61.416 271.188 ; 
        RECT 60.88 266.814 60.984 271.188 ; 
        RECT 60.448 266.814 60.552 271.188 ; 
        RECT 60.016 266.814 60.12 271.188 ; 
        RECT 59.584 266.814 59.688 271.188 ; 
        RECT 59.152 266.814 59.256 271.188 ; 
        RECT 58.72 266.814 58.824 271.188 ; 
        RECT 58.288 266.814 58.392 271.188 ; 
        RECT 57.856 266.814 57.96 271.188 ; 
        RECT 57.424 266.814 57.528 271.188 ; 
        RECT 56.992 266.814 57.096 271.188 ; 
        RECT 56.56 266.814 56.664 271.188 ; 
        RECT 56.128 266.814 56.232 271.188 ; 
        RECT 55.696 266.814 55.8 271.188 ; 
        RECT 55.264 266.814 55.368 271.188 ; 
        RECT 54.832 266.814 54.936 271.188 ; 
        RECT 54.4 266.814 54.504 271.188 ; 
        RECT 53.968 266.814 54.072 271.188 ; 
        RECT 53.536 266.814 53.64 271.188 ; 
        RECT 53.104 266.814 53.208 271.188 ; 
        RECT 52.672 266.814 52.776 271.188 ; 
        RECT 52.24 266.814 52.344 271.188 ; 
        RECT 51.808 266.814 51.912 271.188 ; 
        RECT 51.376 266.814 51.48 271.188 ; 
        RECT 50.944 266.814 51.048 271.188 ; 
        RECT 50.512 266.814 50.616 271.188 ; 
        RECT 50.08 266.814 50.184 271.188 ; 
        RECT 49.648 266.814 49.752 271.188 ; 
        RECT 49.216 266.814 49.32 271.188 ; 
        RECT 48.784 266.814 48.888 271.188 ; 
        RECT 48.352 266.814 48.456 271.188 ; 
        RECT 47.92 266.814 48.024 271.188 ; 
        RECT 47.488 266.814 47.592 271.188 ; 
        RECT 47.056 266.814 47.16 271.188 ; 
        RECT 46.624 266.814 46.728 271.188 ; 
        RECT 46.192 266.814 46.296 271.188 ; 
        RECT 45.76 266.814 45.864 271.188 ; 
        RECT 45.328 266.814 45.432 271.188 ; 
        RECT 44.896 266.814 45 271.188 ; 
        RECT 44.464 266.814 44.568 271.188 ; 
        RECT 44.032 266.814 44.136 271.188 ; 
        RECT 43.6 266.814 43.704 271.188 ; 
        RECT 43.168 266.814 43.272 271.188 ; 
        RECT 42.736 266.814 42.84 271.188 ; 
        RECT 42.304 266.814 42.408 271.188 ; 
        RECT 41.872 266.814 41.976 271.188 ; 
        RECT 41.44 266.814 41.544 271.188 ; 
        RECT 41.008 266.814 41.112 271.188 ; 
        RECT 40.576 266.814 40.68 271.188 ; 
        RECT 40.144 266.814 40.248 271.188 ; 
        RECT 39.712 266.814 39.816 271.188 ; 
        RECT 39.28 266.814 39.384 271.188 ; 
        RECT 38.848 266.814 38.952 271.188 ; 
        RECT 38.416 266.814 38.52 271.188 ; 
        RECT 37.984 266.814 38.088 271.188 ; 
        RECT 37.552 266.814 37.656 271.188 ; 
        RECT 36.7 266.814 37.008 271.188 ; 
        RECT 29.128 266.814 29.436 271.188 ; 
        RECT 28.48 266.814 28.584 271.188 ; 
        RECT 28.048 266.814 28.152 271.188 ; 
        RECT 27.616 266.814 27.72 271.188 ; 
        RECT 27.184 266.814 27.288 271.188 ; 
        RECT 26.752 266.814 26.856 271.188 ; 
        RECT 26.32 266.814 26.424 271.188 ; 
        RECT 25.888 266.814 25.992 271.188 ; 
        RECT 25.456 266.814 25.56 271.188 ; 
        RECT 25.024 266.814 25.128 271.188 ; 
        RECT 24.592 266.814 24.696 271.188 ; 
        RECT 24.16 266.814 24.264 271.188 ; 
        RECT 23.728 266.814 23.832 271.188 ; 
        RECT 23.296 266.814 23.4 271.188 ; 
        RECT 22.864 266.814 22.968 271.188 ; 
        RECT 22.432 266.814 22.536 271.188 ; 
        RECT 22 266.814 22.104 271.188 ; 
        RECT 21.568 266.814 21.672 271.188 ; 
        RECT 21.136 266.814 21.24 271.188 ; 
        RECT 20.704 266.814 20.808 271.188 ; 
        RECT 20.272 266.814 20.376 271.188 ; 
        RECT 19.84 266.814 19.944 271.188 ; 
        RECT 19.408 266.814 19.512 271.188 ; 
        RECT 18.976 266.814 19.08 271.188 ; 
        RECT 18.544 266.814 18.648 271.188 ; 
        RECT 18.112 266.814 18.216 271.188 ; 
        RECT 17.68 266.814 17.784 271.188 ; 
        RECT 17.248 266.814 17.352 271.188 ; 
        RECT 16.816 266.814 16.92 271.188 ; 
        RECT 16.384 266.814 16.488 271.188 ; 
        RECT 15.952 266.814 16.056 271.188 ; 
        RECT 15.52 266.814 15.624 271.188 ; 
        RECT 15.088 266.814 15.192 271.188 ; 
        RECT 14.656 266.814 14.76 271.188 ; 
        RECT 14.224 266.814 14.328 271.188 ; 
        RECT 13.792 266.814 13.896 271.188 ; 
        RECT 13.36 266.814 13.464 271.188 ; 
        RECT 12.928 266.814 13.032 271.188 ; 
        RECT 12.496 266.814 12.6 271.188 ; 
        RECT 12.064 266.814 12.168 271.188 ; 
        RECT 11.632 266.814 11.736 271.188 ; 
        RECT 11.2 266.814 11.304 271.188 ; 
        RECT 10.768 266.814 10.872 271.188 ; 
        RECT 10.336 266.814 10.44 271.188 ; 
        RECT 9.904 266.814 10.008 271.188 ; 
        RECT 9.472 266.814 9.576 271.188 ; 
        RECT 9.04 266.814 9.144 271.188 ; 
        RECT 8.608 266.814 8.712 271.188 ; 
        RECT 8.176 266.814 8.28 271.188 ; 
        RECT 7.744 266.814 7.848 271.188 ; 
        RECT 7.312 266.814 7.416 271.188 ; 
        RECT 6.88 266.814 6.984 271.188 ; 
        RECT 6.448 266.814 6.552 271.188 ; 
        RECT 6.016 266.814 6.12 271.188 ; 
        RECT 5.584 266.814 5.688 271.188 ; 
        RECT 5.152 266.814 5.256 271.188 ; 
        RECT 4.72 266.814 4.824 271.188 ; 
        RECT 4.288 266.814 4.392 271.188 ; 
        RECT 3.856 266.814 3.96 271.188 ; 
        RECT 3.424 266.814 3.528 271.188 ; 
        RECT 2.992 266.814 3.096 271.188 ; 
        RECT 2.56 266.814 2.664 271.188 ; 
        RECT 2.128 266.814 2.232 271.188 ; 
        RECT 1.696 266.814 1.8 271.188 ; 
        RECT 1.264 266.814 1.368 271.188 ; 
        RECT 0.832 266.814 0.936 271.188 ; 
        RECT 0.02 266.814 0.36 271.188 ; 
        RECT 34.564 271.134 35.076 275.508 ; 
        RECT 34.508 273.796 35.076 275.086 ; 
        RECT 33.916 272.704 34.164 275.508 ; 
        RECT 33.86 273.942 34.164 274.556 ; 
        RECT 33.916 271.134 34.02 275.508 ; 
        RECT 33.916 271.618 34.076 272.576 ; 
        RECT 33.916 271.134 34.164 271.49 ; 
        RECT 32.728 272.936 33.552 275.508 ; 
        RECT 33.448 271.134 33.552 275.508 ; 
        RECT 32.728 274.044 33.608 275.076 ; 
        RECT 32.728 271.134 33.12 275.508 ; 
        RECT 31.06 271.134 31.392 275.508 ; 
        RECT 31.06 271.488 31.448 275.23 ; 
        RECT 65.776 271.134 66.116 275.508 ; 
        RECT 65.2 271.134 65.304 275.508 ; 
        RECT 64.768 271.134 64.872 275.508 ; 
        RECT 64.336 271.134 64.44 275.508 ; 
        RECT 63.904 271.134 64.008 275.508 ; 
        RECT 63.472 271.134 63.576 275.508 ; 
        RECT 63.04 271.134 63.144 275.508 ; 
        RECT 62.608 271.134 62.712 275.508 ; 
        RECT 62.176 271.134 62.28 275.508 ; 
        RECT 61.744 271.134 61.848 275.508 ; 
        RECT 61.312 271.134 61.416 275.508 ; 
        RECT 60.88 271.134 60.984 275.508 ; 
        RECT 60.448 271.134 60.552 275.508 ; 
        RECT 60.016 271.134 60.12 275.508 ; 
        RECT 59.584 271.134 59.688 275.508 ; 
        RECT 59.152 271.134 59.256 275.508 ; 
        RECT 58.72 271.134 58.824 275.508 ; 
        RECT 58.288 271.134 58.392 275.508 ; 
        RECT 57.856 271.134 57.96 275.508 ; 
        RECT 57.424 271.134 57.528 275.508 ; 
        RECT 56.992 271.134 57.096 275.508 ; 
        RECT 56.56 271.134 56.664 275.508 ; 
        RECT 56.128 271.134 56.232 275.508 ; 
        RECT 55.696 271.134 55.8 275.508 ; 
        RECT 55.264 271.134 55.368 275.508 ; 
        RECT 54.832 271.134 54.936 275.508 ; 
        RECT 54.4 271.134 54.504 275.508 ; 
        RECT 53.968 271.134 54.072 275.508 ; 
        RECT 53.536 271.134 53.64 275.508 ; 
        RECT 53.104 271.134 53.208 275.508 ; 
        RECT 52.672 271.134 52.776 275.508 ; 
        RECT 52.24 271.134 52.344 275.508 ; 
        RECT 51.808 271.134 51.912 275.508 ; 
        RECT 51.376 271.134 51.48 275.508 ; 
        RECT 50.944 271.134 51.048 275.508 ; 
        RECT 50.512 271.134 50.616 275.508 ; 
        RECT 50.08 271.134 50.184 275.508 ; 
        RECT 49.648 271.134 49.752 275.508 ; 
        RECT 49.216 271.134 49.32 275.508 ; 
        RECT 48.784 271.134 48.888 275.508 ; 
        RECT 48.352 271.134 48.456 275.508 ; 
        RECT 47.92 271.134 48.024 275.508 ; 
        RECT 47.488 271.134 47.592 275.508 ; 
        RECT 47.056 271.134 47.16 275.508 ; 
        RECT 46.624 271.134 46.728 275.508 ; 
        RECT 46.192 271.134 46.296 275.508 ; 
        RECT 45.76 271.134 45.864 275.508 ; 
        RECT 45.328 271.134 45.432 275.508 ; 
        RECT 44.896 271.134 45 275.508 ; 
        RECT 44.464 271.134 44.568 275.508 ; 
        RECT 44.032 271.134 44.136 275.508 ; 
        RECT 43.6 271.134 43.704 275.508 ; 
        RECT 43.168 271.134 43.272 275.508 ; 
        RECT 42.736 271.134 42.84 275.508 ; 
        RECT 42.304 271.134 42.408 275.508 ; 
        RECT 41.872 271.134 41.976 275.508 ; 
        RECT 41.44 271.134 41.544 275.508 ; 
        RECT 41.008 271.134 41.112 275.508 ; 
        RECT 40.576 271.134 40.68 275.508 ; 
        RECT 40.144 271.134 40.248 275.508 ; 
        RECT 39.712 271.134 39.816 275.508 ; 
        RECT 39.28 271.134 39.384 275.508 ; 
        RECT 38.848 271.134 38.952 275.508 ; 
        RECT 38.416 271.134 38.52 275.508 ; 
        RECT 37.984 271.134 38.088 275.508 ; 
        RECT 37.552 271.134 37.656 275.508 ; 
        RECT 36.7 271.134 37.008 275.508 ; 
        RECT 29.128 271.134 29.436 275.508 ; 
        RECT 28.48 271.134 28.584 275.508 ; 
        RECT 28.048 271.134 28.152 275.508 ; 
        RECT 27.616 271.134 27.72 275.508 ; 
        RECT 27.184 271.134 27.288 275.508 ; 
        RECT 26.752 271.134 26.856 275.508 ; 
        RECT 26.32 271.134 26.424 275.508 ; 
        RECT 25.888 271.134 25.992 275.508 ; 
        RECT 25.456 271.134 25.56 275.508 ; 
        RECT 25.024 271.134 25.128 275.508 ; 
        RECT 24.592 271.134 24.696 275.508 ; 
        RECT 24.16 271.134 24.264 275.508 ; 
        RECT 23.728 271.134 23.832 275.508 ; 
        RECT 23.296 271.134 23.4 275.508 ; 
        RECT 22.864 271.134 22.968 275.508 ; 
        RECT 22.432 271.134 22.536 275.508 ; 
        RECT 22 271.134 22.104 275.508 ; 
        RECT 21.568 271.134 21.672 275.508 ; 
        RECT 21.136 271.134 21.24 275.508 ; 
        RECT 20.704 271.134 20.808 275.508 ; 
        RECT 20.272 271.134 20.376 275.508 ; 
        RECT 19.84 271.134 19.944 275.508 ; 
        RECT 19.408 271.134 19.512 275.508 ; 
        RECT 18.976 271.134 19.08 275.508 ; 
        RECT 18.544 271.134 18.648 275.508 ; 
        RECT 18.112 271.134 18.216 275.508 ; 
        RECT 17.68 271.134 17.784 275.508 ; 
        RECT 17.248 271.134 17.352 275.508 ; 
        RECT 16.816 271.134 16.92 275.508 ; 
        RECT 16.384 271.134 16.488 275.508 ; 
        RECT 15.952 271.134 16.056 275.508 ; 
        RECT 15.52 271.134 15.624 275.508 ; 
        RECT 15.088 271.134 15.192 275.508 ; 
        RECT 14.656 271.134 14.76 275.508 ; 
        RECT 14.224 271.134 14.328 275.508 ; 
        RECT 13.792 271.134 13.896 275.508 ; 
        RECT 13.36 271.134 13.464 275.508 ; 
        RECT 12.928 271.134 13.032 275.508 ; 
        RECT 12.496 271.134 12.6 275.508 ; 
        RECT 12.064 271.134 12.168 275.508 ; 
        RECT 11.632 271.134 11.736 275.508 ; 
        RECT 11.2 271.134 11.304 275.508 ; 
        RECT 10.768 271.134 10.872 275.508 ; 
        RECT 10.336 271.134 10.44 275.508 ; 
        RECT 9.904 271.134 10.008 275.508 ; 
        RECT 9.472 271.134 9.576 275.508 ; 
        RECT 9.04 271.134 9.144 275.508 ; 
        RECT 8.608 271.134 8.712 275.508 ; 
        RECT 8.176 271.134 8.28 275.508 ; 
        RECT 7.744 271.134 7.848 275.508 ; 
        RECT 7.312 271.134 7.416 275.508 ; 
        RECT 6.88 271.134 6.984 275.508 ; 
        RECT 6.448 271.134 6.552 275.508 ; 
        RECT 6.016 271.134 6.12 275.508 ; 
        RECT 5.584 271.134 5.688 275.508 ; 
        RECT 5.152 271.134 5.256 275.508 ; 
        RECT 4.72 271.134 4.824 275.508 ; 
        RECT 4.288 271.134 4.392 275.508 ; 
        RECT 3.856 271.134 3.96 275.508 ; 
        RECT 3.424 271.134 3.528 275.508 ; 
        RECT 2.992 271.134 3.096 275.508 ; 
        RECT 2.56 271.134 2.664 275.508 ; 
        RECT 2.128 271.134 2.232 275.508 ; 
        RECT 1.696 271.134 1.8 275.508 ; 
        RECT 1.264 271.134 1.368 275.508 ; 
        RECT 0.832 271.134 0.936 275.508 ; 
        RECT 0.02 271.134 0.36 275.508 ; 
        RECT 34.564 275.454 35.076 279.828 ; 
        RECT 34.508 278.116 35.076 279.406 ; 
        RECT 33.916 277.024 34.164 279.828 ; 
        RECT 33.86 278.262 34.164 278.876 ; 
        RECT 33.916 275.454 34.02 279.828 ; 
        RECT 33.916 275.938 34.076 276.896 ; 
        RECT 33.916 275.454 34.164 275.81 ; 
        RECT 32.728 277.256 33.552 279.828 ; 
        RECT 33.448 275.454 33.552 279.828 ; 
        RECT 32.728 278.364 33.608 279.396 ; 
        RECT 32.728 275.454 33.12 279.828 ; 
        RECT 31.06 275.454 31.392 279.828 ; 
        RECT 31.06 275.808 31.448 279.55 ; 
        RECT 65.776 275.454 66.116 279.828 ; 
        RECT 65.2 275.454 65.304 279.828 ; 
        RECT 64.768 275.454 64.872 279.828 ; 
        RECT 64.336 275.454 64.44 279.828 ; 
        RECT 63.904 275.454 64.008 279.828 ; 
        RECT 63.472 275.454 63.576 279.828 ; 
        RECT 63.04 275.454 63.144 279.828 ; 
        RECT 62.608 275.454 62.712 279.828 ; 
        RECT 62.176 275.454 62.28 279.828 ; 
        RECT 61.744 275.454 61.848 279.828 ; 
        RECT 61.312 275.454 61.416 279.828 ; 
        RECT 60.88 275.454 60.984 279.828 ; 
        RECT 60.448 275.454 60.552 279.828 ; 
        RECT 60.016 275.454 60.12 279.828 ; 
        RECT 59.584 275.454 59.688 279.828 ; 
        RECT 59.152 275.454 59.256 279.828 ; 
        RECT 58.72 275.454 58.824 279.828 ; 
        RECT 58.288 275.454 58.392 279.828 ; 
        RECT 57.856 275.454 57.96 279.828 ; 
        RECT 57.424 275.454 57.528 279.828 ; 
        RECT 56.992 275.454 57.096 279.828 ; 
        RECT 56.56 275.454 56.664 279.828 ; 
        RECT 56.128 275.454 56.232 279.828 ; 
        RECT 55.696 275.454 55.8 279.828 ; 
        RECT 55.264 275.454 55.368 279.828 ; 
        RECT 54.832 275.454 54.936 279.828 ; 
        RECT 54.4 275.454 54.504 279.828 ; 
        RECT 53.968 275.454 54.072 279.828 ; 
        RECT 53.536 275.454 53.64 279.828 ; 
        RECT 53.104 275.454 53.208 279.828 ; 
        RECT 52.672 275.454 52.776 279.828 ; 
        RECT 52.24 275.454 52.344 279.828 ; 
        RECT 51.808 275.454 51.912 279.828 ; 
        RECT 51.376 275.454 51.48 279.828 ; 
        RECT 50.944 275.454 51.048 279.828 ; 
        RECT 50.512 275.454 50.616 279.828 ; 
        RECT 50.08 275.454 50.184 279.828 ; 
        RECT 49.648 275.454 49.752 279.828 ; 
        RECT 49.216 275.454 49.32 279.828 ; 
        RECT 48.784 275.454 48.888 279.828 ; 
        RECT 48.352 275.454 48.456 279.828 ; 
        RECT 47.92 275.454 48.024 279.828 ; 
        RECT 47.488 275.454 47.592 279.828 ; 
        RECT 47.056 275.454 47.16 279.828 ; 
        RECT 46.624 275.454 46.728 279.828 ; 
        RECT 46.192 275.454 46.296 279.828 ; 
        RECT 45.76 275.454 45.864 279.828 ; 
        RECT 45.328 275.454 45.432 279.828 ; 
        RECT 44.896 275.454 45 279.828 ; 
        RECT 44.464 275.454 44.568 279.828 ; 
        RECT 44.032 275.454 44.136 279.828 ; 
        RECT 43.6 275.454 43.704 279.828 ; 
        RECT 43.168 275.454 43.272 279.828 ; 
        RECT 42.736 275.454 42.84 279.828 ; 
        RECT 42.304 275.454 42.408 279.828 ; 
        RECT 41.872 275.454 41.976 279.828 ; 
        RECT 41.44 275.454 41.544 279.828 ; 
        RECT 41.008 275.454 41.112 279.828 ; 
        RECT 40.576 275.454 40.68 279.828 ; 
        RECT 40.144 275.454 40.248 279.828 ; 
        RECT 39.712 275.454 39.816 279.828 ; 
        RECT 39.28 275.454 39.384 279.828 ; 
        RECT 38.848 275.454 38.952 279.828 ; 
        RECT 38.416 275.454 38.52 279.828 ; 
        RECT 37.984 275.454 38.088 279.828 ; 
        RECT 37.552 275.454 37.656 279.828 ; 
        RECT 36.7 275.454 37.008 279.828 ; 
        RECT 29.128 275.454 29.436 279.828 ; 
        RECT 28.48 275.454 28.584 279.828 ; 
        RECT 28.048 275.454 28.152 279.828 ; 
        RECT 27.616 275.454 27.72 279.828 ; 
        RECT 27.184 275.454 27.288 279.828 ; 
        RECT 26.752 275.454 26.856 279.828 ; 
        RECT 26.32 275.454 26.424 279.828 ; 
        RECT 25.888 275.454 25.992 279.828 ; 
        RECT 25.456 275.454 25.56 279.828 ; 
        RECT 25.024 275.454 25.128 279.828 ; 
        RECT 24.592 275.454 24.696 279.828 ; 
        RECT 24.16 275.454 24.264 279.828 ; 
        RECT 23.728 275.454 23.832 279.828 ; 
        RECT 23.296 275.454 23.4 279.828 ; 
        RECT 22.864 275.454 22.968 279.828 ; 
        RECT 22.432 275.454 22.536 279.828 ; 
        RECT 22 275.454 22.104 279.828 ; 
        RECT 21.568 275.454 21.672 279.828 ; 
        RECT 21.136 275.454 21.24 279.828 ; 
        RECT 20.704 275.454 20.808 279.828 ; 
        RECT 20.272 275.454 20.376 279.828 ; 
        RECT 19.84 275.454 19.944 279.828 ; 
        RECT 19.408 275.454 19.512 279.828 ; 
        RECT 18.976 275.454 19.08 279.828 ; 
        RECT 18.544 275.454 18.648 279.828 ; 
        RECT 18.112 275.454 18.216 279.828 ; 
        RECT 17.68 275.454 17.784 279.828 ; 
        RECT 17.248 275.454 17.352 279.828 ; 
        RECT 16.816 275.454 16.92 279.828 ; 
        RECT 16.384 275.454 16.488 279.828 ; 
        RECT 15.952 275.454 16.056 279.828 ; 
        RECT 15.52 275.454 15.624 279.828 ; 
        RECT 15.088 275.454 15.192 279.828 ; 
        RECT 14.656 275.454 14.76 279.828 ; 
        RECT 14.224 275.454 14.328 279.828 ; 
        RECT 13.792 275.454 13.896 279.828 ; 
        RECT 13.36 275.454 13.464 279.828 ; 
        RECT 12.928 275.454 13.032 279.828 ; 
        RECT 12.496 275.454 12.6 279.828 ; 
        RECT 12.064 275.454 12.168 279.828 ; 
        RECT 11.632 275.454 11.736 279.828 ; 
        RECT 11.2 275.454 11.304 279.828 ; 
        RECT 10.768 275.454 10.872 279.828 ; 
        RECT 10.336 275.454 10.44 279.828 ; 
        RECT 9.904 275.454 10.008 279.828 ; 
        RECT 9.472 275.454 9.576 279.828 ; 
        RECT 9.04 275.454 9.144 279.828 ; 
        RECT 8.608 275.454 8.712 279.828 ; 
        RECT 8.176 275.454 8.28 279.828 ; 
        RECT 7.744 275.454 7.848 279.828 ; 
        RECT 7.312 275.454 7.416 279.828 ; 
        RECT 6.88 275.454 6.984 279.828 ; 
        RECT 6.448 275.454 6.552 279.828 ; 
        RECT 6.016 275.454 6.12 279.828 ; 
        RECT 5.584 275.454 5.688 279.828 ; 
        RECT 5.152 275.454 5.256 279.828 ; 
        RECT 4.72 275.454 4.824 279.828 ; 
        RECT 4.288 275.454 4.392 279.828 ; 
        RECT 3.856 275.454 3.96 279.828 ; 
        RECT 3.424 275.454 3.528 279.828 ; 
        RECT 2.992 275.454 3.096 279.828 ; 
        RECT 2.56 275.454 2.664 279.828 ; 
        RECT 2.128 275.454 2.232 279.828 ; 
        RECT 1.696 275.454 1.8 279.828 ; 
        RECT 1.264 275.454 1.368 279.828 ; 
        RECT 0.832 275.454 0.936 279.828 ; 
        RECT 0.02 275.454 0.36 279.828 ; 
        RECT 34.564 279.774 35.076 284.148 ; 
        RECT 34.508 282.436 35.076 283.726 ; 
        RECT 33.916 281.344 34.164 284.148 ; 
        RECT 33.86 282.582 34.164 283.196 ; 
        RECT 33.916 279.774 34.02 284.148 ; 
        RECT 33.916 280.258 34.076 281.216 ; 
        RECT 33.916 279.774 34.164 280.13 ; 
        RECT 32.728 281.576 33.552 284.148 ; 
        RECT 33.448 279.774 33.552 284.148 ; 
        RECT 32.728 282.684 33.608 283.716 ; 
        RECT 32.728 279.774 33.12 284.148 ; 
        RECT 31.06 279.774 31.392 284.148 ; 
        RECT 31.06 280.128 31.448 283.87 ; 
        RECT 65.776 279.774 66.116 284.148 ; 
        RECT 65.2 279.774 65.304 284.148 ; 
        RECT 64.768 279.774 64.872 284.148 ; 
        RECT 64.336 279.774 64.44 284.148 ; 
        RECT 63.904 279.774 64.008 284.148 ; 
        RECT 63.472 279.774 63.576 284.148 ; 
        RECT 63.04 279.774 63.144 284.148 ; 
        RECT 62.608 279.774 62.712 284.148 ; 
        RECT 62.176 279.774 62.28 284.148 ; 
        RECT 61.744 279.774 61.848 284.148 ; 
        RECT 61.312 279.774 61.416 284.148 ; 
        RECT 60.88 279.774 60.984 284.148 ; 
        RECT 60.448 279.774 60.552 284.148 ; 
        RECT 60.016 279.774 60.12 284.148 ; 
        RECT 59.584 279.774 59.688 284.148 ; 
        RECT 59.152 279.774 59.256 284.148 ; 
        RECT 58.72 279.774 58.824 284.148 ; 
        RECT 58.288 279.774 58.392 284.148 ; 
        RECT 57.856 279.774 57.96 284.148 ; 
        RECT 57.424 279.774 57.528 284.148 ; 
        RECT 56.992 279.774 57.096 284.148 ; 
        RECT 56.56 279.774 56.664 284.148 ; 
        RECT 56.128 279.774 56.232 284.148 ; 
        RECT 55.696 279.774 55.8 284.148 ; 
        RECT 55.264 279.774 55.368 284.148 ; 
        RECT 54.832 279.774 54.936 284.148 ; 
        RECT 54.4 279.774 54.504 284.148 ; 
        RECT 53.968 279.774 54.072 284.148 ; 
        RECT 53.536 279.774 53.64 284.148 ; 
        RECT 53.104 279.774 53.208 284.148 ; 
        RECT 52.672 279.774 52.776 284.148 ; 
        RECT 52.24 279.774 52.344 284.148 ; 
        RECT 51.808 279.774 51.912 284.148 ; 
        RECT 51.376 279.774 51.48 284.148 ; 
        RECT 50.944 279.774 51.048 284.148 ; 
        RECT 50.512 279.774 50.616 284.148 ; 
        RECT 50.08 279.774 50.184 284.148 ; 
        RECT 49.648 279.774 49.752 284.148 ; 
        RECT 49.216 279.774 49.32 284.148 ; 
        RECT 48.784 279.774 48.888 284.148 ; 
        RECT 48.352 279.774 48.456 284.148 ; 
        RECT 47.92 279.774 48.024 284.148 ; 
        RECT 47.488 279.774 47.592 284.148 ; 
        RECT 47.056 279.774 47.16 284.148 ; 
        RECT 46.624 279.774 46.728 284.148 ; 
        RECT 46.192 279.774 46.296 284.148 ; 
        RECT 45.76 279.774 45.864 284.148 ; 
        RECT 45.328 279.774 45.432 284.148 ; 
        RECT 44.896 279.774 45 284.148 ; 
        RECT 44.464 279.774 44.568 284.148 ; 
        RECT 44.032 279.774 44.136 284.148 ; 
        RECT 43.6 279.774 43.704 284.148 ; 
        RECT 43.168 279.774 43.272 284.148 ; 
        RECT 42.736 279.774 42.84 284.148 ; 
        RECT 42.304 279.774 42.408 284.148 ; 
        RECT 41.872 279.774 41.976 284.148 ; 
        RECT 41.44 279.774 41.544 284.148 ; 
        RECT 41.008 279.774 41.112 284.148 ; 
        RECT 40.576 279.774 40.68 284.148 ; 
        RECT 40.144 279.774 40.248 284.148 ; 
        RECT 39.712 279.774 39.816 284.148 ; 
        RECT 39.28 279.774 39.384 284.148 ; 
        RECT 38.848 279.774 38.952 284.148 ; 
        RECT 38.416 279.774 38.52 284.148 ; 
        RECT 37.984 279.774 38.088 284.148 ; 
        RECT 37.552 279.774 37.656 284.148 ; 
        RECT 36.7 279.774 37.008 284.148 ; 
        RECT 29.128 279.774 29.436 284.148 ; 
        RECT 28.48 279.774 28.584 284.148 ; 
        RECT 28.048 279.774 28.152 284.148 ; 
        RECT 27.616 279.774 27.72 284.148 ; 
        RECT 27.184 279.774 27.288 284.148 ; 
        RECT 26.752 279.774 26.856 284.148 ; 
        RECT 26.32 279.774 26.424 284.148 ; 
        RECT 25.888 279.774 25.992 284.148 ; 
        RECT 25.456 279.774 25.56 284.148 ; 
        RECT 25.024 279.774 25.128 284.148 ; 
        RECT 24.592 279.774 24.696 284.148 ; 
        RECT 24.16 279.774 24.264 284.148 ; 
        RECT 23.728 279.774 23.832 284.148 ; 
        RECT 23.296 279.774 23.4 284.148 ; 
        RECT 22.864 279.774 22.968 284.148 ; 
        RECT 22.432 279.774 22.536 284.148 ; 
        RECT 22 279.774 22.104 284.148 ; 
        RECT 21.568 279.774 21.672 284.148 ; 
        RECT 21.136 279.774 21.24 284.148 ; 
        RECT 20.704 279.774 20.808 284.148 ; 
        RECT 20.272 279.774 20.376 284.148 ; 
        RECT 19.84 279.774 19.944 284.148 ; 
        RECT 19.408 279.774 19.512 284.148 ; 
        RECT 18.976 279.774 19.08 284.148 ; 
        RECT 18.544 279.774 18.648 284.148 ; 
        RECT 18.112 279.774 18.216 284.148 ; 
        RECT 17.68 279.774 17.784 284.148 ; 
        RECT 17.248 279.774 17.352 284.148 ; 
        RECT 16.816 279.774 16.92 284.148 ; 
        RECT 16.384 279.774 16.488 284.148 ; 
        RECT 15.952 279.774 16.056 284.148 ; 
        RECT 15.52 279.774 15.624 284.148 ; 
        RECT 15.088 279.774 15.192 284.148 ; 
        RECT 14.656 279.774 14.76 284.148 ; 
        RECT 14.224 279.774 14.328 284.148 ; 
        RECT 13.792 279.774 13.896 284.148 ; 
        RECT 13.36 279.774 13.464 284.148 ; 
        RECT 12.928 279.774 13.032 284.148 ; 
        RECT 12.496 279.774 12.6 284.148 ; 
        RECT 12.064 279.774 12.168 284.148 ; 
        RECT 11.632 279.774 11.736 284.148 ; 
        RECT 11.2 279.774 11.304 284.148 ; 
        RECT 10.768 279.774 10.872 284.148 ; 
        RECT 10.336 279.774 10.44 284.148 ; 
        RECT 9.904 279.774 10.008 284.148 ; 
        RECT 9.472 279.774 9.576 284.148 ; 
        RECT 9.04 279.774 9.144 284.148 ; 
        RECT 8.608 279.774 8.712 284.148 ; 
        RECT 8.176 279.774 8.28 284.148 ; 
        RECT 7.744 279.774 7.848 284.148 ; 
        RECT 7.312 279.774 7.416 284.148 ; 
        RECT 6.88 279.774 6.984 284.148 ; 
        RECT 6.448 279.774 6.552 284.148 ; 
        RECT 6.016 279.774 6.12 284.148 ; 
        RECT 5.584 279.774 5.688 284.148 ; 
        RECT 5.152 279.774 5.256 284.148 ; 
        RECT 4.72 279.774 4.824 284.148 ; 
        RECT 4.288 279.774 4.392 284.148 ; 
        RECT 3.856 279.774 3.96 284.148 ; 
        RECT 3.424 279.774 3.528 284.148 ; 
        RECT 2.992 279.774 3.096 284.148 ; 
        RECT 2.56 279.774 2.664 284.148 ; 
        RECT 2.128 279.774 2.232 284.148 ; 
        RECT 1.696 279.774 1.8 284.148 ; 
        RECT 1.264 279.774 1.368 284.148 ; 
        RECT 0.832 279.774 0.936 284.148 ; 
        RECT 0.02 279.774 0.36 284.148 ; 
        RECT 34.564 284.094 35.076 288.468 ; 
        RECT 34.508 286.756 35.076 288.046 ; 
        RECT 33.916 285.664 34.164 288.468 ; 
        RECT 33.86 286.902 34.164 287.516 ; 
        RECT 33.916 284.094 34.02 288.468 ; 
        RECT 33.916 284.578 34.076 285.536 ; 
        RECT 33.916 284.094 34.164 284.45 ; 
        RECT 32.728 285.896 33.552 288.468 ; 
        RECT 33.448 284.094 33.552 288.468 ; 
        RECT 32.728 287.004 33.608 288.036 ; 
        RECT 32.728 284.094 33.12 288.468 ; 
        RECT 31.06 284.094 31.392 288.468 ; 
        RECT 31.06 284.448 31.448 288.19 ; 
        RECT 65.776 284.094 66.116 288.468 ; 
        RECT 65.2 284.094 65.304 288.468 ; 
        RECT 64.768 284.094 64.872 288.468 ; 
        RECT 64.336 284.094 64.44 288.468 ; 
        RECT 63.904 284.094 64.008 288.468 ; 
        RECT 63.472 284.094 63.576 288.468 ; 
        RECT 63.04 284.094 63.144 288.468 ; 
        RECT 62.608 284.094 62.712 288.468 ; 
        RECT 62.176 284.094 62.28 288.468 ; 
        RECT 61.744 284.094 61.848 288.468 ; 
        RECT 61.312 284.094 61.416 288.468 ; 
        RECT 60.88 284.094 60.984 288.468 ; 
        RECT 60.448 284.094 60.552 288.468 ; 
        RECT 60.016 284.094 60.12 288.468 ; 
        RECT 59.584 284.094 59.688 288.468 ; 
        RECT 59.152 284.094 59.256 288.468 ; 
        RECT 58.72 284.094 58.824 288.468 ; 
        RECT 58.288 284.094 58.392 288.468 ; 
        RECT 57.856 284.094 57.96 288.468 ; 
        RECT 57.424 284.094 57.528 288.468 ; 
        RECT 56.992 284.094 57.096 288.468 ; 
        RECT 56.56 284.094 56.664 288.468 ; 
        RECT 56.128 284.094 56.232 288.468 ; 
        RECT 55.696 284.094 55.8 288.468 ; 
        RECT 55.264 284.094 55.368 288.468 ; 
        RECT 54.832 284.094 54.936 288.468 ; 
        RECT 54.4 284.094 54.504 288.468 ; 
        RECT 53.968 284.094 54.072 288.468 ; 
        RECT 53.536 284.094 53.64 288.468 ; 
        RECT 53.104 284.094 53.208 288.468 ; 
        RECT 52.672 284.094 52.776 288.468 ; 
        RECT 52.24 284.094 52.344 288.468 ; 
        RECT 51.808 284.094 51.912 288.468 ; 
        RECT 51.376 284.094 51.48 288.468 ; 
        RECT 50.944 284.094 51.048 288.468 ; 
        RECT 50.512 284.094 50.616 288.468 ; 
        RECT 50.08 284.094 50.184 288.468 ; 
        RECT 49.648 284.094 49.752 288.468 ; 
        RECT 49.216 284.094 49.32 288.468 ; 
        RECT 48.784 284.094 48.888 288.468 ; 
        RECT 48.352 284.094 48.456 288.468 ; 
        RECT 47.92 284.094 48.024 288.468 ; 
        RECT 47.488 284.094 47.592 288.468 ; 
        RECT 47.056 284.094 47.16 288.468 ; 
        RECT 46.624 284.094 46.728 288.468 ; 
        RECT 46.192 284.094 46.296 288.468 ; 
        RECT 45.76 284.094 45.864 288.468 ; 
        RECT 45.328 284.094 45.432 288.468 ; 
        RECT 44.896 284.094 45 288.468 ; 
        RECT 44.464 284.094 44.568 288.468 ; 
        RECT 44.032 284.094 44.136 288.468 ; 
        RECT 43.6 284.094 43.704 288.468 ; 
        RECT 43.168 284.094 43.272 288.468 ; 
        RECT 42.736 284.094 42.84 288.468 ; 
        RECT 42.304 284.094 42.408 288.468 ; 
        RECT 41.872 284.094 41.976 288.468 ; 
        RECT 41.44 284.094 41.544 288.468 ; 
        RECT 41.008 284.094 41.112 288.468 ; 
        RECT 40.576 284.094 40.68 288.468 ; 
        RECT 40.144 284.094 40.248 288.468 ; 
        RECT 39.712 284.094 39.816 288.468 ; 
        RECT 39.28 284.094 39.384 288.468 ; 
        RECT 38.848 284.094 38.952 288.468 ; 
        RECT 38.416 284.094 38.52 288.468 ; 
        RECT 37.984 284.094 38.088 288.468 ; 
        RECT 37.552 284.094 37.656 288.468 ; 
        RECT 36.7 284.094 37.008 288.468 ; 
        RECT 29.128 284.094 29.436 288.468 ; 
        RECT 28.48 284.094 28.584 288.468 ; 
        RECT 28.048 284.094 28.152 288.468 ; 
        RECT 27.616 284.094 27.72 288.468 ; 
        RECT 27.184 284.094 27.288 288.468 ; 
        RECT 26.752 284.094 26.856 288.468 ; 
        RECT 26.32 284.094 26.424 288.468 ; 
        RECT 25.888 284.094 25.992 288.468 ; 
        RECT 25.456 284.094 25.56 288.468 ; 
        RECT 25.024 284.094 25.128 288.468 ; 
        RECT 24.592 284.094 24.696 288.468 ; 
        RECT 24.16 284.094 24.264 288.468 ; 
        RECT 23.728 284.094 23.832 288.468 ; 
        RECT 23.296 284.094 23.4 288.468 ; 
        RECT 22.864 284.094 22.968 288.468 ; 
        RECT 22.432 284.094 22.536 288.468 ; 
        RECT 22 284.094 22.104 288.468 ; 
        RECT 21.568 284.094 21.672 288.468 ; 
        RECT 21.136 284.094 21.24 288.468 ; 
        RECT 20.704 284.094 20.808 288.468 ; 
        RECT 20.272 284.094 20.376 288.468 ; 
        RECT 19.84 284.094 19.944 288.468 ; 
        RECT 19.408 284.094 19.512 288.468 ; 
        RECT 18.976 284.094 19.08 288.468 ; 
        RECT 18.544 284.094 18.648 288.468 ; 
        RECT 18.112 284.094 18.216 288.468 ; 
        RECT 17.68 284.094 17.784 288.468 ; 
        RECT 17.248 284.094 17.352 288.468 ; 
        RECT 16.816 284.094 16.92 288.468 ; 
        RECT 16.384 284.094 16.488 288.468 ; 
        RECT 15.952 284.094 16.056 288.468 ; 
        RECT 15.52 284.094 15.624 288.468 ; 
        RECT 15.088 284.094 15.192 288.468 ; 
        RECT 14.656 284.094 14.76 288.468 ; 
        RECT 14.224 284.094 14.328 288.468 ; 
        RECT 13.792 284.094 13.896 288.468 ; 
        RECT 13.36 284.094 13.464 288.468 ; 
        RECT 12.928 284.094 13.032 288.468 ; 
        RECT 12.496 284.094 12.6 288.468 ; 
        RECT 12.064 284.094 12.168 288.468 ; 
        RECT 11.632 284.094 11.736 288.468 ; 
        RECT 11.2 284.094 11.304 288.468 ; 
        RECT 10.768 284.094 10.872 288.468 ; 
        RECT 10.336 284.094 10.44 288.468 ; 
        RECT 9.904 284.094 10.008 288.468 ; 
        RECT 9.472 284.094 9.576 288.468 ; 
        RECT 9.04 284.094 9.144 288.468 ; 
        RECT 8.608 284.094 8.712 288.468 ; 
        RECT 8.176 284.094 8.28 288.468 ; 
        RECT 7.744 284.094 7.848 288.468 ; 
        RECT 7.312 284.094 7.416 288.468 ; 
        RECT 6.88 284.094 6.984 288.468 ; 
        RECT 6.448 284.094 6.552 288.468 ; 
        RECT 6.016 284.094 6.12 288.468 ; 
        RECT 5.584 284.094 5.688 288.468 ; 
        RECT 5.152 284.094 5.256 288.468 ; 
        RECT 4.72 284.094 4.824 288.468 ; 
        RECT 4.288 284.094 4.392 288.468 ; 
        RECT 3.856 284.094 3.96 288.468 ; 
        RECT 3.424 284.094 3.528 288.468 ; 
        RECT 2.992 284.094 3.096 288.468 ; 
        RECT 2.56 284.094 2.664 288.468 ; 
        RECT 2.128 284.094 2.232 288.468 ; 
        RECT 1.696 284.094 1.8 288.468 ; 
        RECT 1.264 284.094 1.368 288.468 ; 
        RECT 0.832 284.094 0.936 288.468 ; 
        RECT 0.02 284.094 0.36 288.468 ; 
        RECT 34.564 288.414 35.076 292.788 ; 
        RECT 34.508 291.076 35.076 292.366 ; 
        RECT 33.916 289.984 34.164 292.788 ; 
        RECT 33.86 291.222 34.164 291.836 ; 
        RECT 33.916 288.414 34.02 292.788 ; 
        RECT 33.916 288.898 34.076 289.856 ; 
        RECT 33.916 288.414 34.164 288.77 ; 
        RECT 32.728 290.216 33.552 292.788 ; 
        RECT 33.448 288.414 33.552 292.788 ; 
        RECT 32.728 291.324 33.608 292.356 ; 
        RECT 32.728 288.414 33.12 292.788 ; 
        RECT 31.06 288.414 31.392 292.788 ; 
        RECT 31.06 288.768 31.448 292.51 ; 
        RECT 65.776 288.414 66.116 292.788 ; 
        RECT 65.2 288.414 65.304 292.788 ; 
        RECT 64.768 288.414 64.872 292.788 ; 
        RECT 64.336 288.414 64.44 292.788 ; 
        RECT 63.904 288.414 64.008 292.788 ; 
        RECT 63.472 288.414 63.576 292.788 ; 
        RECT 63.04 288.414 63.144 292.788 ; 
        RECT 62.608 288.414 62.712 292.788 ; 
        RECT 62.176 288.414 62.28 292.788 ; 
        RECT 61.744 288.414 61.848 292.788 ; 
        RECT 61.312 288.414 61.416 292.788 ; 
        RECT 60.88 288.414 60.984 292.788 ; 
        RECT 60.448 288.414 60.552 292.788 ; 
        RECT 60.016 288.414 60.12 292.788 ; 
        RECT 59.584 288.414 59.688 292.788 ; 
        RECT 59.152 288.414 59.256 292.788 ; 
        RECT 58.72 288.414 58.824 292.788 ; 
        RECT 58.288 288.414 58.392 292.788 ; 
        RECT 57.856 288.414 57.96 292.788 ; 
        RECT 57.424 288.414 57.528 292.788 ; 
        RECT 56.992 288.414 57.096 292.788 ; 
        RECT 56.56 288.414 56.664 292.788 ; 
        RECT 56.128 288.414 56.232 292.788 ; 
        RECT 55.696 288.414 55.8 292.788 ; 
        RECT 55.264 288.414 55.368 292.788 ; 
        RECT 54.832 288.414 54.936 292.788 ; 
        RECT 54.4 288.414 54.504 292.788 ; 
        RECT 53.968 288.414 54.072 292.788 ; 
        RECT 53.536 288.414 53.64 292.788 ; 
        RECT 53.104 288.414 53.208 292.788 ; 
        RECT 52.672 288.414 52.776 292.788 ; 
        RECT 52.24 288.414 52.344 292.788 ; 
        RECT 51.808 288.414 51.912 292.788 ; 
        RECT 51.376 288.414 51.48 292.788 ; 
        RECT 50.944 288.414 51.048 292.788 ; 
        RECT 50.512 288.414 50.616 292.788 ; 
        RECT 50.08 288.414 50.184 292.788 ; 
        RECT 49.648 288.414 49.752 292.788 ; 
        RECT 49.216 288.414 49.32 292.788 ; 
        RECT 48.784 288.414 48.888 292.788 ; 
        RECT 48.352 288.414 48.456 292.788 ; 
        RECT 47.92 288.414 48.024 292.788 ; 
        RECT 47.488 288.414 47.592 292.788 ; 
        RECT 47.056 288.414 47.16 292.788 ; 
        RECT 46.624 288.414 46.728 292.788 ; 
        RECT 46.192 288.414 46.296 292.788 ; 
        RECT 45.76 288.414 45.864 292.788 ; 
        RECT 45.328 288.414 45.432 292.788 ; 
        RECT 44.896 288.414 45 292.788 ; 
        RECT 44.464 288.414 44.568 292.788 ; 
        RECT 44.032 288.414 44.136 292.788 ; 
        RECT 43.6 288.414 43.704 292.788 ; 
        RECT 43.168 288.414 43.272 292.788 ; 
        RECT 42.736 288.414 42.84 292.788 ; 
        RECT 42.304 288.414 42.408 292.788 ; 
        RECT 41.872 288.414 41.976 292.788 ; 
        RECT 41.44 288.414 41.544 292.788 ; 
        RECT 41.008 288.414 41.112 292.788 ; 
        RECT 40.576 288.414 40.68 292.788 ; 
        RECT 40.144 288.414 40.248 292.788 ; 
        RECT 39.712 288.414 39.816 292.788 ; 
        RECT 39.28 288.414 39.384 292.788 ; 
        RECT 38.848 288.414 38.952 292.788 ; 
        RECT 38.416 288.414 38.52 292.788 ; 
        RECT 37.984 288.414 38.088 292.788 ; 
        RECT 37.552 288.414 37.656 292.788 ; 
        RECT 36.7 288.414 37.008 292.788 ; 
        RECT 29.128 288.414 29.436 292.788 ; 
        RECT 28.48 288.414 28.584 292.788 ; 
        RECT 28.048 288.414 28.152 292.788 ; 
        RECT 27.616 288.414 27.72 292.788 ; 
        RECT 27.184 288.414 27.288 292.788 ; 
        RECT 26.752 288.414 26.856 292.788 ; 
        RECT 26.32 288.414 26.424 292.788 ; 
        RECT 25.888 288.414 25.992 292.788 ; 
        RECT 25.456 288.414 25.56 292.788 ; 
        RECT 25.024 288.414 25.128 292.788 ; 
        RECT 24.592 288.414 24.696 292.788 ; 
        RECT 24.16 288.414 24.264 292.788 ; 
        RECT 23.728 288.414 23.832 292.788 ; 
        RECT 23.296 288.414 23.4 292.788 ; 
        RECT 22.864 288.414 22.968 292.788 ; 
        RECT 22.432 288.414 22.536 292.788 ; 
        RECT 22 288.414 22.104 292.788 ; 
        RECT 21.568 288.414 21.672 292.788 ; 
        RECT 21.136 288.414 21.24 292.788 ; 
        RECT 20.704 288.414 20.808 292.788 ; 
        RECT 20.272 288.414 20.376 292.788 ; 
        RECT 19.84 288.414 19.944 292.788 ; 
        RECT 19.408 288.414 19.512 292.788 ; 
        RECT 18.976 288.414 19.08 292.788 ; 
        RECT 18.544 288.414 18.648 292.788 ; 
        RECT 18.112 288.414 18.216 292.788 ; 
        RECT 17.68 288.414 17.784 292.788 ; 
        RECT 17.248 288.414 17.352 292.788 ; 
        RECT 16.816 288.414 16.92 292.788 ; 
        RECT 16.384 288.414 16.488 292.788 ; 
        RECT 15.952 288.414 16.056 292.788 ; 
        RECT 15.52 288.414 15.624 292.788 ; 
        RECT 15.088 288.414 15.192 292.788 ; 
        RECT 14.656 288.414 14.76 292.788 ; 
        RECT 14.224 288.414 14.328 292.788 ; 
        RECT 13.792 288.414 13.896 292.788 ; 
        RECT 13.36 288.414 13.464 292.788 ; 
        RECT 12.928 288.414 13.032 292.788 ; 
        RECT 12.496 288.414 12.6 292.788 ; 
        RECT 12.064 288.414 12.168 292.788 ; 
        RECT 11.632 288.414 11.736 292.788 ; 
        RECT 11.2 288.414 11.304 292.788 ; 
        RECT 10.768 288.414 10.872 292.788 ; 
        RECT 10.336 288.414 10.44 292.788 ; 
        RECT 9.904 288.414 10.008 292.788 ; 
        RECT 9.472 288.414 9.576 292.788 ; 
        RECT 9.04 288.414 9.144 292.788 ; 
        RECT 8.608 288.414 8.712 292.788 ; 
        RECT 8.176 288.414 8.28 292.788 ; 
        RECT 7.744 288.414 7.848 292.788 ; 
        RECT 7.312 288.414 7.416 292.788 ; 
        RECT 6.88 288.414 6.984 292.788 ; 
        RECT 6.448 288.414 6.552 292.788 ; 
        RECT 6.016 288.414 6.12 292.788 ; 
        RECT 5.584 288.414 5.688 292.788 ; 
        RECT 5.152 288.414 5.256 292.788 ; 
        RECT 4.72 288.414 4.824 292.788 ; 
        RECT 4.288 288.414 4.392 292.788 ; 
        RECT 3.856 288.414 3.96 292.788 ; 
        RECT 3.424 288.414 3.528 292.788 ; 
        RECT 2.992 288.414 3.096 292.788 ; 
        RECT 2.56 288.414 2.664 292.788 ; 
        RECT 2.128 288.414 2.232 292.788 ; 
        RECT 1.696 288.414 1.8 292.788 ; 
        RECT 1.264 288.414 1.368 292.788 ; 
        RECT 0.832 288.414 0.936 292.788 ; 
        RECT 0.02 288.414 0.36 292.788 ; 
        RECT 34.564 292.734 35.076 297.108 ; 
        RECT 34.508 295.396 35.076 296.686 ; 
        RECT 33.916 294.304 34.164 297.108 ; 
        RECT 33.86 295.542 34.164 296.156 ; 
        RECT 33.916 292.734 34.02 297.108 ; 
        RECT 33.916 293.218 34.076 294.176 ; 
        RECT 33.916 292.734 34.164 293.09 ; 
        RECT 32.728 294.536 33.552 297.108 ; 
        RECT 33.448 292.734 33.552 297.108 ; 
        RECT 32.728 295.644 33.608 296.676 ; 
        RECT 32.728 292.734 33.12 297.108 ; 
        RECT 31.06 292.734 31.392 297.108 ; 
        RECT 31.06 293.088 31.448 296.83 ; 
        RECT 65.776 292.734 66.116 297.108 ; 
        RECT 65.2 292.734 65.304 297.108 ; 
        RECT 64.768 292.734 64.872 297.108 ; 
        RECT 64.336 292.734 64.44 297.108 ; 
        RECT 63.904 292.734 64.008 297.108 ; 
        RECT 63.472 292.734 63.576 297.108 ; 
        RECT 63.04 292.734 63.144 297.108 ; 
        RECT 62.608 292.734 62.712 297.108 ; 
        RECT 62.176 292.734 62.28 297.108 ; 
        RECT 61.744 292.734 61.848 297.108 ; 
        RECT 61.312 292.734 61.416 297.108 ; 
        RECT 60.88 292.734 60.984 297.108 ; 
        RECT 60.448 292.734 60.552 297.108 ; 
        RECT 60.016 292.734 60.12 297.108 ; 
        RECT 59.584 292.734 59.688 297.108 ; 
        RECT 59.152 292.734 59.256 297.108 ; 
        RECT 58.72 292.734 58.824 297.108 ; 
        RECT 58.288 292.734 58.392 297.108 ; 
        RECT 57.856 292.734 57.96 297.108 ; 
        RECT 57.424 292.734 57.528 297.108 ; 
        RECT 56.992 292.734 57.096 297.108 ; 
        RECT 56.56 292.734 56.664 297.108 ; 
        RECT 56.128 292.734 56.232 297.108 ; 
        RECT 55.696 292.734 55.8 297.108 ; 
        RECT 55.264 292.734 55.368 297.108 ; 
        RECT 54.832 292.734 54.936 297.108 ; 
        RECT 54.4 292.734 54.504 297.108 ; 
        RECT 53.968 292.734 54.072 297.108 ; 
        RECT 53.536 292.734 53.64 297.108 ; 
        RECT 53.104 292.734 53.208 297.108 ; 
        RECT 52.672 292.734 52.776 297.108 ; 
        RECT 52.24 292.734 52.344 297.108 ; 
        RECT 51.808 292.734 51.912 297.108 ; 
        RECT 51.376 292.734 51.48 297.108 ; 
        RECT 50.944 292.734 51.048 297.108 ; 
        RECT 50.512 292.734 50.616 297.108 ; 
        RECT 50.08 292.734 50.184 297.108 ; 
        RECT 49.648 292.734 49.752 297.108 ; 
        RECT 49.216 292.734 49.32 297.108 ; 
        RECT 48.784 292.734 48.888 297.108 ; 
        RECT 48.352 292.734 48.456 297.108 ; 
        RECT 47.92 292.734 48.024 297.108 ; 
        RECT 47.488 292.734 47.592 297.108 ; 
        RECT 47.056 292.734 47.16 297.108 ; 
        RECT 46.624 292.734 46.728 297.108 ; 
        RECT 46.192 292.734 46.296 297.108 ; 
        RECT 45.76 292.734 45.864 297.108 ; 
        RECT 45.328 292.734 45.432 297.108 ; 
        RECT 44.896 292.734 45 297.108 ; 
        RECT 44.464 292.734 44.568 297.108 ; 
        RECT 44.032 292.734 44.136 297.108 ; 
        RECT 43.6 292.734 43.704 297.108 ; 
        RECT 43.168 292.734 43.272 297.108 ; 
        RECT 42.736 292.734 42.84 297.108 ; 
        RECT 42.304 292.734 42.408 297.108 ; 
        RECT 41.872 292.734 41.976 297.108 ; 
        RECT 41.44 292.734 41.544 297.108 ; 
        RECT 41.008 292.734 41.112 297.108 ; 
        RECT 40.576 292.734 40.68 297.108 ; 
        RECT 40.144 292.734 40.248 297.108 ; 
        RECT 39.712 292.734 39.816 297.108 ; 
        RECT 39.28 292.734 39.384 297.108 ; 
        RECT 38.848 292.734 38.952 297.108 ; 
        RECT 38.416 292.734 38.52 297.108 ; 
        RECT 37.984 292.734 38.088 297.108 ; 
        RECT 37.552 292.734 37.656 297.108 ; 
        RECT 36.7 292.734 37.008 297.108 ; 
        RECT 29.128 292.734 29.436 297.108 ; 
        RECT 28.48 292.734 28.584 297.108 ; 
        RECT 28.048 292.734 28.152 297.108 ; 
        RECT 27.616 292.734 27.72 297.108 ; 
        RECT 27.184 292.734 27.288 297.108 ; 
        RECT 26.752 292.734 26.856 297.108 ; 
        RECT 26.32 292.734 26.424 297.108 ; 
        RECT 25.888 292.734 25.992 297.108 ; 
        RECT 25.456 292.734 25.56 297.108 ; 
        RECT 25.024 292.734 25.128 297.108 ; 
        RECT 24.592 292.734 24.696 297.108 ; 
        RECT 24.16 292.734 24.264 297.108 ; 
        RECT 23.728 292.734 23.832 297.108 ; 
        RECT 23.296 292.734 23.4 297.108 ; 
        RECT 22.864 292.734 22.968 297.108 ; 
        RECT 22.432 292.734 22.536 297.108 ; 
        RECT 22 292.734 22.104 297.108 ; 
        RECT 21.568 292.734 21.672 297.108 ; 
        RECT 21.136 292.734 21.24 297.108 ; 
        RECT 20.704 292.734 20.808 297.108 ; 
        RECT 20.272 292.734 20.376 297.108 ; 
        RECT 19.84 292.734 19.944 297.108 ; 
        RECT 19.408 292.734 19.512 297.108 ; 
        RECT 18.976 292.734 19.08 297.108 ; 
        RECT 18.544 292.734 18.648 297.108 ; 
        RECT 18.112 292.734 18.216 297.108 ; 
        RECT 17.68 292.734 17.784 297.108 ; 
        RECT 17.248 292.734 17.352 297.108 ; 
        RECT 16.816 292.734 16.92 297.108 ; 
        RECT 16.384 292.734 16.488 297.108 ; 
        RECT 15.952 292.734 16.056 297.108 ; 
        RECT 15.52 292.734 15.624 297.108 ; 
        RECT 15.088 292.734 15.192 297.108 ; 
        RECT 14.656 292.734 14.76 297.108 ; 
        RECT 14.224 292.734 14.328 297.108 ; 
        RECT 13.792 292.734 13.896 297.108 ; 
        RECT 13.36 292.734 13.464 297.108 ; 
        RECT 12.928 292.734 13.032 297.108 ; 
        RECT 12.496 292.734 12.6 297.108 ; 
        RECT 12.064 292.734 12.168 297.108 ; 
        RECT 11.632 292.734 11.736 297.108 ; 
        RECT 11.2 292.734 11.304 297.108 ; 
        RECT 10.768 292.734 10.872 297.108 ; 
        RECT 10.336 292.734 10.44 297.108 ; 
        RECT 9.904 292.734 10.008 297.108 ; 
        RECT 9.472 292.734 9.576 297.108 ; 
        RECT 9.04 292.734 9.144 297.108 ; 
        RECT 8.608 292.734 8.712 297.108 ; 
        RECT 8.176 292.734 8.28 297.108 ; 
        RECT 7.744 292.734 7.848 297.108 ; 
        RECT 7.312 292.734 7.416 297.108 ; 
        RECT 6.88 292.734 6.984 297.108 ; 
        RECT 6.448 292.734 6.552 297.108 ; 
        RECT 6.016 292.734 6.12 297.108 ; 
        RECT 5.584 292.734 5.688 297.108 ; 
        RECT 5.152 292.734 5.256 297.108 ; 
        RECT 4.72 292.734 4.824 297.108 ; 
        RECT 4.288 292.734 4.392 297.108 ; 
        RECT 3.856 292.734 3.96 297.108 ; 
        RECT 3.424 292.734 3.528 297.108 ; 
        RECT 2.992 292.734 3.096 297.108 ; 
        RECT 2.56 292.734 2.664 297.108 ; 
        RECT 2.128 292.734 2.232 297.108 ; 
        RECT 1.696 292.734 1.8 297.108 ; 
        RECT 1.264 292.734 1.368 297.108 ; 
        RECT 0.832 292.734 0.936 297.108 ; 
        RECT 0.02 292.734 0.36 297.108 ; 
        RECT 34.564 297.054 35.076 301.428 ; 
        RECT 34.508 299.716 35.076 301.006 ; 
        RECT 33.916 298.624 34.164 301.428 ; 
        RECT 33.86 299.862 34.164 300.476 ; 
        RECT 33.916 297.054 34.02 301.428 ; 
        RECT 33.916 297.538 34.076 298.496 ; 
        RECT 33.916 297.054 34.164 297.41 ; 
        RECT 32.728 298.856 33.552 301.428 ; 
        RECT 33.448 297.054 33.552 301.428 ; 
        RECT 32.728 299.964 33.608 300.996 ; 
        RECT 32.728 297.054 33.12 301.428 ; 
        RECT 31.06 297.054 31.392 301.428 ; 
        RECT 31.06 297.408 31.448 301.15 ; 
        RECT 65.776 297.054 66.116 301.428 ; 
        RECT 65.2 297.054 65.304 301.428 ; 
        RECT 64.768 297.054 64.872 301.428 ; 
        RECT 64.336 297.054 64.44 301.428 ; 
        RECT 63.904 297.054 64.008 301.428 ; 
        RECT 63.472 297.054 63.576 301.428 ; 
        RECT 63.04 297.054 63.144 301.428 ; 
        RECT 62.608 297.054 62.712 301.428 ; 
        RECT 62.176 297.054 62.28 301.428 ; 
        RECT 61.744 297.054 61.848 301.428 ; 
        RECT 61.312 297.054 61.416 301.428 ; 
        RECT 60.88 297.054 60.984 301.428 ; 
        RECT 60.448 297.054 60.552 301.428 ; 
        RECT 60.016 297.054 60.12 301.428 ; 
        RECT 59.584 297.054 59.688 301.428 ; 
        RECT 59.152 297.054 59.256 301.428 ; 
        RECT 58.72 297.054 58.824 301.428 ; 
        RECT 58.288 297.054 58.392 301.428 ; 
        RECT 57.856 297.054 57.96 301.428 ; 
        RECT 57.424 297.054 57.528 301.428 ; 
        RECT 56.992 297.054 57.096 301.428 ; 
        RECT 56.56 297.054 56.664 301.428 ; 
        RECT 56.128 297.054 56.232 301.428 ; 
        RECT 55.696 297.054 55.8 301.428 ; 
        RECT 55.264 297.054 55.368 301.428 ; 
        RECT 54.832 297.054 54.936 301.428 ; 
        RECT 54.4 297.054 54.504 301.428 ; 
        RECT 53.968 297.054 54.072 301.428 ; 
        RECT 53.536 297.054 53.64 301.428 ; 
        RECT 53.104 297.054 53.208 301.428 ; 
        RECT 52.672 297.054 52.776 301.428 ; 
        RECT 52.24 297.054 52.344 301.428 ; 
        RECT 51.808 297.054 51.912 301.428 ; 
        RECT 51.376 297.054 51.48 301.428 ; 
        RECT 50.944 297.054 51.048 301.428 ; 
        RECT 50.512 297.054 50.616 301.428 ; 
        RECT 50.08 297.054 50.184 301.428 ; 
        RECT 49.648 297.054 49.752 301.428 ; 
        RECT 49.216 297.054 49.32 301.428 ; 
        RECT 48.784 297.054 48.888 301.428 ; 
        RECT 48.352 297.054 48.456 301.428 ; 
        RECT 47.92 297.054 48.024 301.428 ; 
        RECT 47.488 297.054 47.592 301.428 ; 
        RECT 47.056 297.054 47.16 301.428 ; 
        RECT 46.624 297.054 46.728 301.428 ; 
        RECT 46.192 297.054 46.296 301.428 ; 
        RECT 45.76 297.054 45.864 301.428 ; 
        RECT 45.328 297.054 45.432 301.428 ; 
        RECT 44.896 297.054 45 301.428 ; 
        RECT 44.464 297.054 44.568 301.428 ; 
        RECT 44.032 297.054 44.136 301.428 ; 
        RECT 43.6 297.054 43.704 301.428 ; 
        RECT 43.168 297.054 43.272 301.428 ; 
        RECT 42.736 297.054 42.84 301.428 ; 
        RECT 42.304 297.054 42.408 301.428 ; 
        RECT 41.872 297.054 41.976 301.428 ; 
        RECT 41.44 297.054 41.544 301.428 ; 
        RECT 41.008 297.054 41.112 301.428 ; 
        RECT 40.576 297.054 40.68 301.428 ; 
        RECT 40.144 297.054 40.248 301.428 ; 
        RECT 39.712 297.054 39.816 301.428 ; 
        RECT 39.28 297.054 39.384 301.428 ; 
        RECT 38.848 297.054 38.952 301.428 ; 
        RECT 38.416 297.054 38.52 301.428 ; 
        RECT 37.984 297.054 38.088 301.428 ; 
        RECT 37.552 297.054 37.656 301.428 ; 
        RECT 36.7 297.054 37.008 301.428 ; 
        RECT 29.128 297.054 29.436 301.428 ; 
        RECT 28.48 297.054 28.584 301.428 ; 
        RECT 28.048 297.054 28.152 301.428 ; 
        RECT 27.616 297.054 27.72 301.428 ; 
        RECT 27.184 297.054 27.288 301.428 ; 
        RECT 26.752 297.054 26.856 301.428 ; 
        RECT 26.32 297.054 26.424 301.428 ; 
        RECT 25.888 297.054 25.992 301.428 ; 
        RECT 25.456 297.054 25.56 301.428 ; 
        RECT 25.024 297.054 25.128 301.428 ; 
        RECT 24.592 297.054 24.696 301.428 ; 
        RECT 24.16 297.054 24.264 301.428 ; 
        RECT 23.728 297.054 23.832 301.428 ; 
        RECT 23.296 297.054 23.4 301.428 ; 
        RECT 22.864 297.054 22.968 301.428 ; 
        RECT 22.432 297.054 22.536 301.428 ; 
        RECT 22 297.054 22.104 301.428 ; 
        RECT 21.568 297.054 21.672 301.428 ; 
        RECT 21.136 297.054 21.24 301.428 ; 
        RECT 20.704 297.054 20.808 301.428 ; 
        RECT 20.272 297.054 20.376 301.428 ; 
        RECT 19.84 297.054 19.944 301.428 ; 
        RECT 19.408 297.054 19.512 301.428 ; 
        RECT 18.976 297.054 19.08 301.428 ; 
        RECT 18.544 297.054 18.648 301.428 ; 
        RECT 18.112 297.054 18.216 301.428 ; 
        RECT 17.68 297.054 17.784 301.428 ; 
        RECT 17.248 297.054 17.352 301.428 ; 
        RECT 16.816 297.054 16.92 301.428 ; 
        RECT 16.384 297.054 16.488 301.428 ; 
        RECT 15.952 297.054 16.056 301.428 ; 
        RECT 15.52 297.054 15.624 301.428 ; 
        RECT 15.088 297.054 15.192 301.428 ; 
        RECT 14.656 297.054 14.76 301.428 ; 
        RECT 14.224 297.054 14.328 301.428 ; 
        RECT 13.792 297.054 13.896 301.428 ; 
        RECT 13.36 297.054 13.464 301.428 ; 
        RECT 12.928 297.054 13.032 301.428 ; 
        RECT 12.496 297.054 12.6 301.428 ; 
        RECT 12.064 297.054 12.168 301.428 ; 
        RECT 11.632 297.054 11.736 301.428 ; 
        RECT 11.2 297.054 11.304 301.428 ; 
        RECT 10.768 297.054 10.872 301.428 ; 
        RECT 10.336 297.054 10.44 301.428 ; 
        RECT 9.904 297.054 10.008 301.428 ; 
        RECT 9.472 297.054 9.576 301.428 ; 
        RECT 9.04 297.054 9.144 301.428 ; 
        RECT 8.608 297.054 8.712 301.428 ; 
        RECT 8.176 297.054 8.28 301.428 ; 
        RECT 7.744 297.054 7.848 301.428 ; 
        RECT 7.312 297.054 7.416 301.428 ; 
        RECT 6.88 297.054 6.984 301.428 ; 
        RECT 6.448 297.054 6.552 301.428 ; 
        RECT 6.016 297.054 6.12 301.428 ; 
        RECT 5.584 297.054 5.688 301.428 ; 
        RECT 5.152 297.054 5.256 301.428 ; 
        RECT 4.72 297.054 4.824 301.428 ; 
        RECT 4.288 297.054 4.392 301.428 ; 
        RECT 3.856 297.054 3.96 301.428 ; 
        RECT 3.424 297.054 3.528 301.428 ; 
        RECT 2.992 297.054 3.096 301.428 ; 
        RECT 2.56 297.054 2.664 301.428 ; 
        RECT 2.128 297.054 2.232 301.428 ; 
        RECT 1.696 297.054 1.8 301.428 ; 
        RECT 1.264 297.054 1.368 301.428 ; 
        RECT 0.832 297.054 0.936 301.428 ; 
        RECT 0.02 297.054 0.36 301.428 ; 
        RECT 34.564 301.374 35.076 305.748 ; 
        RECT 34.508 304.036 35.076 305.326 ; 
        RECT 33.916 302.944 34.164 305.748 ; 
        RECT 33.86 304.182 34.164 304.796 ; 
        RECT 33.916 301.374 34.02 305.748 ; 
        RECT 33.916 301.858 34.076 302.816 ; 
        RECT 33.916 301.374 34.164 301.73 ; 
        RECT 32.728 303.176 33.552 305.748 ; 
        RECT 33.448 301.374 33.552 305.748 ; 
        RECT 32.728 304.284 33.608 305.316 ; 
        RECT 32.728 301.374 33.12 305.748 ; 
        RECT 31.06 301.374 31.392 305.748 ; 
        RECT 31.06 301.728 31.448 305.47 ; 
        RECT 65.776 301.374 66.116 305.748 ; 
        RECT 65.2 301.374 65.304 305.748 ; 
        RECT 64.768 301.374 64.872 305.748 ; 
        RECT 64.336 301.374 64.44 305.748 ; 
        RECT 63.904 301.374 64.008 305.748 ; 
        RECT 63.472 301.374 63.576 305.748 ; 
        RECT 63.04 301.374 63.144 305.748 ; 
        RECT 62.608 301.374 62.712 305.748 ; 
        RECT 62.176 301.374 62.28 305.748 ; 
        RECT 61.744 301.374 61.848 305.748 ; 
        RECT 61.312 301.374 61.416 305.748 ; 
        RECT 60.88 301.374 60.984 305.748 ; 
        RECT 60.448 301.374 60.552 305.748 ; 
        RECT 60.016 301.374 60.12 305.748 ; 
        RECT 59.584 301.374 59.688 305.748 ; 
        RECT 59.152 301.374 59.256 305.748 ; 
        RECT 58.72 301.374 58.824 305.748 ; 
        RECT 58.288 301.374 58.392 305.748 ; 
        RECT 57.856 301.374 57.96 305.748 ; 
        RECT 57.424 301.374 57.528 305.748 ; 
        RECT 56.992 301.374 57.096 305.748 ; 
        RECT 56.56 301.374 56.664 305.748 ; 
        RECT 56.128 301.374 56.232 305.748 ; 
        RECT 55.696 301.374 55.8 305.748 ; 
        RECT 55.264 301.374 55.368 305.748 ; 
        RECT 54.832 301.374 54.936 305.748 ; 
        RECT 54.4 301.374 54.504 305.748 ; 
        RECT 53.968 301.374 54.072 305.748 ; 
        RECT 53.536 301.374 53.64 305.748 ; 
        RECT 53.104 301.374 53.208 305.748 ; 
        RECT 52.672 301.374 52.776 305.748 ; 
        RECT 52.24 301.374 52.344 305.748 ; 
        RECT 51.808 301.374 51.912 305.748 ; 
        RECT 51.376 301.374 51.48 305.748 ; 
        RECT 50.944 301.374 51.048 305.748 ; 
        RECT 50.512 301.374 50.616 305.748 ; 
        RECT 50.08 301.374 50.184 305.748 ; 
        RECT 49.648 301.374 49.752 305.748 ; 
        RECT 49.216 301.374 49.32 305.748 ; 
        RECT 48.784 301.374 48.888 305.748 ; 
        RECT 48.352 301.374 48.456 305.748 ; 
        RECT 47.92 301.374 48.024 305.748 ; 
        RECT 47.488 301.374 47.592 305.748 ; 
        RECT 47.056 301.374 47.16 305.748 ; 
        RECT 46.624 301.374 46.728 305.748 ; 
        RECT 46.192 301.374 46.296 305.748 ; 
        RECT 45.76 301.374 45.864 305.748 ; 
        RECT 45.328 301.374 45.432 305.748 ; 
        RECT 44.896 301.374 45 305.748 ; 
        RECT 44.464 301.374 44.568 305.748 ; 
        RECT 44.032 301.374 44.136 305.748 ; 
        RECT 43.6 301.374 43.704 305.748 ; 
        RECT 43.168 301.374 43.272 305.748 ; 
        RECT 42.736 301.374 42.84 305.748 ; 
        RECT 42.304 301.374 42.408 305.748 ; 
        RECT 41.872 301.374 41.976 305.748 ; 
        RECT 41.44 301.374 41.544 305.748 ; 
        RECT 41.008 301.374 41.112 305.748 ; 
        RECT 40.576 301.374 40.68 305.748 ; 
        RECT 40.144 301.374 40.248 305.748 ; 
        RECT 39.712 301.374 39.816 305.748 ; 
        RECT 39.28 301.374 39.384 305.748 ; 
        RECT 38.848 301.374 38.952 305.748 ; 
        RECT 38.416 301.374 38.52 305.748 ; 
        RECT 37.984 301.374 38.088 305.748 ; 
        RECT 37.552 301.374 37.656 305.748 ; 
        RECT 36.7 301.374 37.008 305.748 ; 
        RECT 29.128 301.374 29.436 305.748 ; 
        RECT 28.48 301.374 28.584 305.748 ; 
        RECT 28.048 301.374 28.152 305.748 ; 
        RECT 27.616 301.374 27.72 305.748 ; 
        RECT 27.184 301.374 27.288 305.748 ; 
        RECT 26.752 301.374 26.856 305.748 ; 
        RECT 26.32 301.374 26.424 305.748 ; 
        RECT 25.888 301.374 25.992 305.748 ; 
        RECT 25.456 301.374 25.56 305.748 ; 
        RECT 25.024 301.374 25.128 305.748 ; 
        RECT 24.592 301.374 24.696 305.748 ; 
        RECT 24.16 301.374 24.264 305.748 ; 
        RECT 23.728 301.374 23.832 305.748 ; 
        RECT 23.296 301.374 23.4 305.748 ; 
        RECT 22.864 301.374 22.968 305.748 ; 
        RECT 22.432 301.374 22.536 305.748 ; 
        RECT 22 301.374 22.104 305.748 ; 
        RECT 21.568 301.374 21.672 305.748 ; 
        RECT 21.136 301.374 21.24 305.748 ; 
        RECT 20.704 301.374 20.808 305.748 ; 
        RECT 20.272 301.374 20.376 305.748 ; 
        RECT 19.84 301.374 19.944 305.748 ; 
        RECT 19.408 301.374 19.512 305.748 ; 
        RECT 18.976 301.374 19.08 305.748 ; 
        RECT 18.544 301.374 18.648 305.748 ; 
        RECT 18.112 301.374 18.216 305.748 ; 
        RECT 17.68 301.374 17.784 305.748 ; 
        RECT 17.248 301.374 17.352 305.748 ; 
        RECT 16.816 301.374 16.92 305.748 ; 
        RECT 16.384 301.374 16.488 305.748 ; 
        RECT 15.952 301.374 16.056 305.748 ; 
        RECT 15.52 301.374 15.624 305.748 ; 
        RECT 15.088 301.374 15.192 305.748 ; 
        RECT 14.656 301.374 14.76 305.748 ; 
        RECT 14.224 301.374 14.328 305.748 ; 
        RECT 13.792 301.374 13.896 305.748 ; 
        RECT 13.36 301.374 13.464 305.748 ; 
        RECT 12.928 301.374 13.032 305.748 ; 
        RECT 12.496 301.374 12.6 305.748 ; 
        RECT 12.064 301.374 12.168 305.748 ; 
        RECT 11.632 301.374 11.736 305.748 ; 
        RECT 11.2 301.374 11.304 305.748 ; 
        RECT 10.768 301.374 10.872 305.748 ; 
        RECT 10.336 301.374 10.44 305.748 ; 
        RECT 9.904 301.374 10.008 305.748 ; 
        RECT 9.472 301.374 9.576 305.748 ; 
        RECT 9.04 301.374 9.144 305.748 ; 
        RECT 8.608 301.374 8.712 305.748 ; 
        RECT 8.176 301.374 8.28 305.748 ; 
        RECT 7.744 301.374 7.848 305.748 ; 
        RECT 7.312 301.374 7.416 305.748 ; 
        RECT 6.88 301.374 6.984 305.748 ; 
        RECT 6.448 301.374 6.552 305.748 ; 
        RECT 6.016 301.374 6.12 305.748 ; 
        RECT 5.584 301.374 5.688 305.748 ; 
        RECT 5.152 301.374 5.256 305.748 ; 
        RECT 4.72 301.374 4.824 305.748 ; 
        RECT 4.288 301.374 4.392 305.748 ; 
        RECT 3.856 301.374 3.96 305.748 ; 
        RECT 3.424 301.374 3.528 305.748 ; 
        RECT 2.992 301.374 3.096 305.748 ; 
        RECT 2.56 301.374 2.664 305.748 ; 
        RECT 2.128 301.374 2.232 305.748 ; 
        RECT 1.696 301.374 1.8 305.748 ; 
        RECT 1.264 301.374 1.368 305.748 ; 
        RECT 0.832 301.374 0.936 305.748 ; 
        RECT 0.02 301.374 0.36 305.748 ; 
        RECT 34.564 305.694 35.076 310.068 ; 
        RECT 34.508 308.356 35.076 309.646 ; 
        RECT 33.916 307.264 34.164 310.068 ; 
        RECT 33.86 308.502 34.164 309.116 ; 
        RECT 33.916 305.694 34.02 310.068 ; 
        RECT 33.916 306.178 34.076 307.136 ; 
        RECT 33.916 305.694 34.164 306.05 ; 
        RECT 32.728 307.496 33.552 310.068 ; 
        RECT 33.448 305.694 33.552 310.068 ; 
        RECT 32.728 308.604 33.608 309.636 ; 
        RECT 32.728 305.694 33.12 310.068 ; 
        RECT 31.06 305.694 31.392 310.068 ; 
        RECT 31.06 306.048 31.448 309.79 ; 
        RECT 65.776 305.694 66.116 310.068 ; 
        RECT 65.2 305.694 65.304 310.068 ; 
        RECT 64.768 305.694 64.872 310.068 ; 
        RECT 64.336 305.694 64.44 310.068 ; 
        RECT 63.904 305.694 64.008 310.068 ; 
        RECT 63.472 305.694 63.576 310.068 ; 
        RECT 63.04 305.694 63.144 310.068 ; 
        RECT 62.608 305.694 62.712 310.068 ; 
        RECT 62.176 305.694 62.28 310.068 ; 
        RECT 61.744 305.694 61.848 310.068 ; 
        RECT 61.312 305.694 61.416 310.068 ; 
        RECT 60.88 305.694 60.984 310.068 ; 
        RECT 60.448 305.694 60.552 310.068 ; 
        RECT 60.016 305.694 60.12 310.068 ; 
        RECT 59.584 305.694 59.688 310.068 ; 
        RECT 59.152 305.694 59.256 310.068 ; 
        RECT 58.72 305.694 58.824 310.068 ; 
        RECT 58.288 305.694 58.392 310.068 ; 
        RECT 57.856 305.694 57.96 310.068 ; 
        RECT 57.424 305.694 57.528 310.068 ; 
        RECT 56.992 305.694 57.096 310.068 ; 
        RECT 56.56 305.694 56.664 310.068 ; 
        RECT 56.128 305.694 56.232 310.068 ; 
        RECT 55.696 305.694 55.8 310.068 ; 
        RECT 55.264 305.694 55.368 310.068 ; 
        RECT 54.832 305.694 54.936 310.068 ; 
        RECT 54.4 305.694 54.504 310.068 ; 
        RECT 53.968 305.694 54.072 310.068 ; 
        RECT 53.536 305.694 53.64 310.068 ; 
        RECT 53.104 305.694 53.208 310.068 ; 
        RECT 52.672 305.694 52.776 310.068 ; 
        RECT 52.24 305.694 52.344 310.068 ; 
        RECT 51.808 305.694 51.912 310.068 ; 
        RECT 51.376 305.694 51.48 310.068 ; 
        RECT 50.944 305.694 51.048 310.068 ; 
        RECT 50.512 305.694 50.616 310.068 ; 
        RECT 50.08 305.694 50.184 310.068 ; 
        RECT 49.648 305.694 49.752 310.068 ; 
        RECT 49.216 305.694 49.32 310.068 ; 
        RECT 48.784 305.694 48.888 310.068 ; 
        RECT 48.352 305.694 48.456 310.068 ; 
        RECT 47.92 305.694 48.024 310.068 ; 
        RECT 47.488 305.694 47.592 310.068 ; 
        RECT 47.056 305.694 47.16 310.068 ; 
        RECT 46.624 305.694 46.728 310.068 ; 
        RECT 46.192 305.694 46.296 310.068 ; 
        RECT 45.76 305.694 45.864 310.068 ; 
        RECT 45.328 305.694 45.432 310.068 ; 
        RECT 44.896 305.694 45 310.068 ; 
        RECT 44.464 305.694 44.568 310.068 ; 
        RECT 44.032 305.694 44.136 310.068 ; 
        RECT 43.6 305.694 43.704 310.068 ; 
        RECT 43.168 305.694 43.272 310.068 ; 
        RECT 42.736 305.694 42.84 310.068 ; 
        RECT 42.304 305.694 42.408 310.068 ; 
        RECT 41.872 305.694 41.976 310.068 ; 
        RECT 41.44 305.694 41.544 310.068 ; 
        RECT 41.008 305.694 41.112 310.068 ; 
        RECT 40.576 305.694 40.68 310.068 ; 
        RECT 40.144 305.694 40.248 310.068 ; 
        RECT 39.712 305.694 39.816 310.068 ; 
        RECT 39.28 305.694 39.384 310.068 ; 
        RECT 38.848 305.694 38.952 310.068 ; 
        RECT 38.416 305.694 38.52 310.068 ; 
        RECT 37.984 305.694 38.088 310.068 ; 
        RECT 37.552 305.694 37.656 310.068 ; 
        RECT 36.7 305.694 37.008 310.068 ; 
        RECT 29.128 305.694 29.436 310.068 ; 
        RECT 28.48 305.694 28.584 310.068 ; 
        RECT 28.048 305.694 28.152 310.068 ; 
        RECT 27.616 305.694 27.72 310.068 ; 
        RECT 27.184 305.694 27.288 310.068 ; 
        RECT 26.752 305.694 26.856 310.068 ; 
        RECT 26.32 305.694 26.424 310.068 ; 
        RECT 25.888 305.694 25.992 310.068 ; 
        RECT 25.456 305.694 25.56 310.068 ; 
        RECT 25.024 305.694 25.128 310.068 ; 
        RECT 24.592 305.694 24.696 310.068 ; 
        RECT 24.16 305.694 24.264 310.068 ; 
        RECT 23.728 305.694 23.832 310.068 ; 
        RECT 23.296 305.694 23.4 310.068 ; 
        RECT 22.864 305.694 22.968 310.068 ; 
        RECT 22.432 305.694 22.536 310.068 ; 
        RECT 22 305.694 22.104 310.068 ; 
        RECT 21.568 305.694 21.672 310.068 ; 
        RECT 21.136 305.694 21.24 310.068 ; 
        RECT 20.704 305.694 20.808 310.068 ; 
        RECT 20.272 305.694 20.376 310.068 ; 
        RECT 19.84 305.694 19.944 310.068 ; 
        RECT 19.408 305.694 19.512 310.068 ; 
        RECT 18.976 305.694 19.08 310.068 ; 
        RECT 18.544 305.694 18.648 310.068 ; 
        RECT 18.112 305.694 18.216 310.068 ; 
        RECT 17.68 305.694 17.784 310.068 ; 
        RECT 17.248 305.694 17.352 310.068 ; 
        RECT 16.816 305.694 16.92 310.068 ; 
        RECT 16.384 305.694 16.488 310.068 ; 
        RECT 15.952 305.694 16.056 310.068 ; 
        RECT 15.52 305.694 15.624 310.068 ; 
        RECT 15.088 305.694 15.192 310.068 ; 
        RECT 14.656 305.694 14.76 310.068 ; 
        RECT 14.224 305.694 14.328 310.068 ; 
        RECT 13.792 305.694 13.896 310.068 ; 
        RECT 13.36 305.694 13.464 310.068 ; 
        RECT 12.928 305.694 13.032 310.068 ; 
        RECT 12.496 305.694 12.6 310.068 ; 
        RECT 12.064 305.694 12.168 310.068 ; 
        RECT 11.632 305.694 11.736 310.068 ; 
        RECT 11.2 305.694 11.304 310.068 ; 
        RECT 10.768 305.694 10.872 310.068 ; 
        RECT 10.336 305.694 10.44 310.068 ; 
        RECT 9.904 305.694 10.008 310.068 ; 
        RECT 9.472 305.694 9.576 310.068 ; 
        RECT 9.04 305.694 9.144 310.068 ; 
        RECT 8.608 305.694 8.712 310.068 ; 
        RECT 8.176 305.694 8.28 310.068 ; 
        RECT 7.744 305.694 7.848 310.068 ; 
        RECT 7.312 305.694 7.416 310.068 ; 
        RECT 6.88 305.694 6.984 310.068 ; 
        RECT 6.448 305.694 6.552 310.068 ; 
        RECT 6.016 305.694 6.12 310.068 ; 
        RECT 5.584 305.694 5.688 310.068 ; 
        RECT 5.152 305.694 5.256 310.068 ; 
        RECT 4.72 305.694 4.824 310.068 ; 
        RECT 4.288 305.694 4.392 310.068 ; 
        RECT 3.856 305.694 3.96 310.068 ; 
        RECT 3.424 305.694 3.528 310.068 ; 
        RECT 2.992 305.694 3.096 310.068 ; 
        RECT 2.56 305.694 2.664 310.068 ; 
        RECT 2.128 305.694 2.232 310.068 ; 
        RECT 1.696 305.694 1.8 310.068 ; 
        RECT 1.264 305.694 1.368 310.068 ; 
        RECT 0.832 305.694 0.936 310.068 ; 
        RECT 0.02 305.694 0.36 310.068 ; 
        RECT 34.564 310.014 35.076 314.388 ; 
        RECT 34.508 312.676 35.076 313.966 ; 
        RECT 33.916 311.584 34.164 314.388 ; 
        RECT 33.86 312.822 34.164 313.436 ; 
        RECT 33.916 310.014 34.02 314.388 ; 
        RECT 33.916 310.498 34.076 311.456 ; 
        RECT 33.916 310.014 34.164 310.37 ; 
        RECT 32.728 311.816 33.552 314.388 ; 
        RECT 33.448 310.014 33.552 314.388 ; 
        RECT 32.728 312.924 33.608 313.956 ; 
        RECT 32.728 310.014 33.12 314.388 ; 
        RECT 31.06 310.014 31.392 314.388 ; 
        RECT 31.06 310.368 31.448 314.11 ; 
        RECT 65.776 310.014 66.116 314.388 ; 
        RECT 65.2 310.014 65.304 314.388 ; 
        RECT 64.768 310.014 64.872 314.388 ; 
        RECT 64.336 310.014 64.44 314.388 ; 
        RECT 63.904 310.014 64.008 314.388 ; 
        RECT 63.472 310.014 63.576 314.388 ; 
        RECT 63.04 310.014 63.144 314.388 ; 
        RECT 62.608 310.014 62.712 314.388 ; 
        RECT 62.176 310.014 62.28 314.388 ; 
        RECT 61.744 310.014 61.848 314.388 ; 
        RECT 61.312 310.014 61.416 314.388 ; 
        RECT 60.88 310.014 60.984 314.388 ; 
        RECT 60.448 310.014 60.552 314.388 ; 
        RECT 60.016 310.014 60.12 314.388 ; 
        RECT 59.584 310.014 59.688 314.388 ; 
        RECT 59.152 310.014 59.256 314.388 ; 
        RECT 58.72 310.014 58.824 314.388 ; 
        RECT 58.288 310.014 58.392 314.388 ; 
        RECT 57.856 310.014 57.96 314.388 ; 
        RECT 57.424 310.014 57.528 314.388 ; 
        RECT 56.992 310.014 57.096 314.388 ; 
        RECT 56.56 310.014 56.664 314.388 ; 
        RECT 56.128 310.014 56.232 314.388 ; 
        RECT 55.696 310.014 55.8 314.388 ; 
        RECT 55.264 310.014 55.368 314.388 ; 
        RECT 54.832 310.014 54.936 314.388 ; 
        RECT 54.4 310.014 54.504 314.388 ; 
        RECT 53.968 310.014 54.072 314.388 ; 
        RECT 53.536 310.014 53.64 314.388 ; 
        RECT 53.104 310.014 53.208 314.388 ; 
        RECT 52.672 310.014 52.776 314.388 ; 
        RECT 52.24 310.014 52.344 314.388 ; 
        RECT 51.808 310.014 51.912 314.388 ; 
        RECT 51.376 310.014 51.48 314.388 ; 
        RECT 50.944 310.014 51.048 314.388 ; 
        RECT 50.512 310.014 50.616 314.388 ; 
        RECT 50.08 310.014 50.184 314.388 ; 
        RECT 49.648 310.014 49.752 314.388 ; 
        RECT 49.216 310.014 49.32 314.388 ; 
        RECT 48.784 310.014 48.888 314.388 ; 
        RECT 48.352 310.014 48.456 314.388 ; 
        RECT 47.92 310.014 48.024 314.388 ; 
        RECT 47.488 310.014 47.592 314.388 ; 
        RECT 47.056 310.014 47.16 314.388 ; 
        RECT 46.624 310.014 46.728 314.388 ; 
        RECT 46.192 310.014 46.296 314.388 ; 
        RECT 45.76 310.014 45.864 314.388 ; 
        RECT 45.328 310.014 45.432 314.388 ; 
        RECT 44.896 310.014 45 314.388 ; 
        RECT 44.464 310.014 44.568 314.388 ; 
        RECT 44.032 310.014 44.136 314.388 ; 
        RECT 43.6 310.014 43.704 314.388 ; 
        RECT 43.168 310.014 43.272 314.388 ; 
        RECT 42.736 310.014 42.84 314.388 ; 
        RECT 42.304 310.014 42.408 314.388 ; 
        RECT 41.872 310.014 41.976 314.388 ; 
        RECT 41.44 310.014 41.544 314.388 ; 
        RECT 41.008 310.014 41.112 314.388 ; 
        RECT 40.576 310.014 40.68 314.388 ; 
        RECT 40.144 310.014 40.248 314.388 ; 
        RECT 39.712 310.014 39.816 314.388 ; 
        RECT 39.28 310.014 39.384 314.388 ; 
        RECT 38.848 310.014 38.952 314.388 ; 
        RECT 38.416 310.014 38.52 314.388 ; 
        RECT 37.984 310.014 38.088 314.388 ; 
        RECT 37.552 310.014 37.656 314.388 ; 
        RECT 36.7 310.014 37.008 314.388 ; 
        RECT 29.128 310.014 29.436 314.388 ; 
        RECT 28.48 310.014 28.584 314.388 ; 
        RECT 28.048 310.014 28.152 314.388 ; 
        RECT 27.616 310.014 27.72 314.388 ; 
        RECT 27.184 310.014 27.288 314.388 ; 
        RECT 26.752 310.014 26.856 314.388 ; 
        RECT 26.32 310.014 26.424 314.388 ; 
        RECT 25.888 310.014 25.992 314.388 ; 
        RECT 25.456 310.014 25.56 314.388 ; 
        RECT 25.024 310.014 25.128 314.388 ; 
        RECT 24.592 310.014 24.696 314.388 ; 
        RECT 24.16 310.014 24.264 314.388 ; 
        RECT 23.728 310.014 23.832 314.388 ; 
        RECT 23.296 310.014 23.4 314.388 ; 
        RECT 22.864 310.014 22.968 314.388 ; 
        RECT 22.432 310.014 22.536 314.388 ; 
        RECT 22 310.014 22.104 314.388 ; 
        RECT 21.568 310.014 21.672 314.388 ; 
        RECT 21.136 310.014 21.24 314.388 ; 
        RECT 20.704 310.014 20.808 314.388 ; 
        RECT 20.272 310.014 20.376 314.388 ; 
        RECT 19.84 310.014 19.944 314.388 ; 
        RECT 19.408 310.014 19.512 314.388 ; 
        RECT 18.976 310.014 19.08 314.388 ; 
        RECT 18.544 310.014 18.648 314.388 ; 
        RECT 18.112 310.014 18.216 314.388 ; 
        RECT 17.68 310.014 17.784 314.388 ; 
        RECT 17.248 310.014 17.352 314.388 ; 
        RECT 16.816 310.014 16.92 314.388 ; 
        RECT 16.384 310.014 16.488 314.388 ; 
        RECT 15.952 310.014 16.056 314.388 ; 
        RECT 15.52 310.014 15.624 314.388 ; 
        RECT 15.088 310.014 15.192 314.388 ; 
        RECT 14.656 310.014 14.76 314.388 ; 
        RECT 14.224 310.014 14.328 314.388 ; 
        RECT 13.792 310.014 13.896 314.388 ; 
        RECT 13.36 310.014 13.464 314.388 ; 
        RECT 12.928 310.014 13.032 314.388 ; 
        RECT 12.496 310.014 12.6 314.388 ; 
        RECT 12.064 310.014 12.168 314.388 ; 
        RECT 11.632 310.014 11.736 314.388 ; 
        RECT 11.2 310.014 11.304 314.388 ; 
        RECT 10.768 310.014 10.872 314.388 ; 
        RECT 10.336 310.014 10.44 314.388 ; 
        RECT 9.904 310.014 10.008 314.388 ; 
        RECT 9.472 310.014 9.576 314.388 ; 
        RECT 9.04 310.014 9.144 314.388 ; 
        RECT 8.608 310.014 8.712 314.388 ; 
        RECT 8.176 310.014 8.28 314.388 ; 
        RECT 7.744 310.014 7.848 314.388 ; 
        RECT 7.312 310.014 7.416 314.388 ; 
        RECT 6.88 310.014 6.984 314.388 ; 
        RECT 6.448 310.014 6.552 314.388 ; 
        RECT 6.016 310.014 6.12 314.388 ; 
        RECT 5.584 310.014 5.688 314.388 ; 
        RECT 5.152 310.014 5.256 314.388 ; 
        RECT 4.72 310.014 4.824 314.388 ; 
        RECT 4.288 310.014 4.392 314.388 ; 
        RECT 3.856 310.014 3.96 314.388 ; 
        RECT 3.424 310.014 3.528 314.388 ; 
        RECT 2.992 310.014 3.096 314.388 ; 
        RECT 2.56 310.014 2.664 314.388 ; 
        RECT 2.128 310.014 2.232 314.388 ; 
        RECT 1.696 310.014 1.8 314.388 ; 
        RECT 1.264 310.014 1.368 314.388 ; 
        RECT 0.832 310.014 0.936 314.388 ; 
        RECT 0.02 310.014 0.36 314.388 ; 
        RECT 34.564 314.334 35.076 318.708 ; 
        RECT 34.508 316.996 35.076 318.286 ; 
        RECT 33.916 315.904 34.164 318.708 ; 
        RECT 33.86 317.142 34.164 317.756 ; 
        RECT 33.916 314.334 34.02 318.708 ; 
        RECT 33.916 314.818 34.076 315.776 ; 
        RECT 33.916 314.334 34.164 314.69 ; 
        RECT 32.728 316.136 33.552 318.708 ; 
        RECT 33.448 314.334 33.552 318.708 ; 
        RECT 32.728 317.244 33.608 318.276 ; 
        RECT 32.728 314.334 33.12 318.708 ; 
        RECT 31.06 314.334 31.392 318.708 ; 
        RECT 31.06 314.688 31.448 318.43 ; 
        RECT 65.776 314.334 66.116 318.708 ; 
        RECT 65.2 314.334 65.304 318.708 ; 
        RECT 64.768 314.334 64.872 318.708 ; 
        RECT 64.336 314.334 64.44 318.708 ; 
        RECT 63.904 314.334 64.008 318.708 ; 
        RECT 63.472 314.334 63.576 318.708 ; 
        RECT 63.04 314.334 63.144 318.708 ; 
        RECT 62.608 314.334 62.712 318.708 ; 
        RECT 62.176 314.334 62.28 318.708 ; 
        RECT 61.744 314.334 61.848 318.708 ; 
        RECT 61.312 314.334 61.416 318.708 ; 
        RECT 60.88 314.334 60.984 318.708 ; 
        RECT 60.448 314.334 60.552 318.708 ; 
        RECT 60.016 314.334 60.12 318.708 ; 
        RECT 59.584 314.334 59.688 318.708 ; 
        RECT 59.152 314.334 59.256 318.708 ; 
        RECT 58.72 314.334 58.824 318.708 ; 
        RECT 58.288 314.334 58.392 318.708 ; 
        RECT 57.856 314.334 57.96 318.708 ; 
        RECT 57.424 314.334 57.528 318.708 ; 
        RECT 56.992 314.334 57.096 318.708 ; 
        RECT 56.56 314.334 56.664 318.708 ; 
        RECT 56.128 314.334 56.232 318.708 ; 
        RECT 55.696 314.334 55.8 318.708 ; 
        RECT 55.264 314.334 55.368 318.708 ; 
        RECT 54.832 314.334 54.936 318.708 ; 
        RECT 54.4 314.334 54.504 318.708 ; 
        RECT 53.968 314.334 54.072 318.708 ; 
        RECT 53.536 314.334 53.64 318.708 ; 
        RECT 53.104 314.334 53.208 318.708 ; 
        RECT 52.672 314.334 52.776 318.708 ; 
        RECT 52.24 314.334 52.344 318.708 ; 
        RECT 51.808 314.334 51.912 318.708 ; 
        RECT 51.376 314.334 51.48 318.708 ; 
        RECT 50.944 314.334 51.048 318.708 ; 
        RECT 50.512 314.334 50.616 318.708 ; 
        RECT 50.08 314.334 50.184 318.708 ; 
        RECT 49.648 314.334 49.752 318.708 ; 
        RECT 49.216 314.334 49.32 318.708 ; 
        RECT 48.784 314.334 48.888 318.708 ; 
        RECT 48.352 314.334 48.456 318.708 ; 
        RECT 47.92 314.334 48.024 318.708 ; 
        RECT 47.488 314.334 47.592 318.708 ; 
        RECT 47.056 314.334 47.16 318.708 ; 
        RECT 46.624 314.334 46.728 318.708 ; 
        RECT 46.192 314.334 46.296 318.708 ; 
        RECT 45.76 314.334 45.864 318.708 ; 
        RECT 45.328 314.334 45.432 318.708 ; 
        RECT 44.896 314.334 45 318.708 ; 
        RECT 44.464 314.334 44.568 318.708 ; 
        RECT 44.032 314.334 44.136 318.708 ; 
        RECT 43.6 314.334 43.704 318.708 ; 
        RECT 43.168 314.334 43.272 318.708 ; 
        RECT 42.736 314.334 42.84 318.708 ; 
        RECT 42.304 314.334 42.408 318.708 ; 
        RECT 41.872 314.334 41.976 318.708 ; 
        RECT 41.44 314.334 41.544 318.708 ; 
        RECT 41.008 314.334 41.112 318.708 ; 
        RECT 40.576 314.334 40.68 318.708 ; 
        RECT 40.144 314.334 40.248 318.708 ; 
        RECT 39.712 314.334 39.816 318.708 ; 
        RECT 39.28 314.334 39.384 318.708 ; 
        RECT 38.848 314.334 38.952 318.708 ; 
        RECT 38.416 314.334 38.52 318.708 ; 
        RECT 37.984 314.334 38.088 318.708 ; 
        RECT 37.552 314.334 37.656 318.708 ; 
        RECT 36.7 314.334 37.008 318.708 ; 
        RECT 29.128 314.334 29.436 318.708 ; 
        RECT 28.48 314.334 28.584 318.708 ; 
        RECT 28.048 314.334 28.152 318.708 ; 
        RECT 27.616 314.334 27.72 318.708 ; 
        RECT 27.184 314.334 27.288 318.708 ; 
        RECT 26.752 314.334 26.856 318.708 ; 
        RECT 26.32 314.334 26.424 318.708 ; 
        RECT 25.888 314.334 25.992 318.708 ; 
        RECT 25.456 314.334 25.56 318.708 ; 
        RECT 25.024 314.334 25.128 318.708 ; 
        RECT 24.592 314.334 24.696 318.708 ; 
        RECT 24.16 314.334 24.264 318.708 ; 
        RECT 23.728 314.334 23.832 318.708 ; 
        RECT 23.296 314.334 23.4 318.708 ; 
        RECT 22.864 314.334 22.968 318.708 ; 
        RECT 22.432 314.334 22.536 318.708 ; 
        RECT 22 314.334 22.104 318.708 ; 
        RECT 21.568 314.334 21.672 318.708 ; 
        RECT 21.136 314.334 21.24 318.708 ; 
        RECT 20.704 314.334 20.808 318.708 ; 
        RECT 20.272 314.334 20.376 318.708 ; 
        RECT 19.84 314.334 19.944 318.708 ; 
        RECT 19.408 314.334 19.512 318.708 ; 
        RECT 18.976 314.334 19.08 318.708 ; 
        RECT 18.544 314.334 18.648 318.708 ; 
        RECT 18.112 314.334 18.216 318.708 ; 
        RECT 17.68 314.334 17.784 318.708 ; 
        RECT 17.248 314.334 17.352 318.708 ; 
        RECT 16.816 314.334 16.92 318.708 ; 
        RECT 16.384 314.334 16.488 318.708 ; 
        RECT 15.952 314.334 16.056 318.708 ; 
        RECT 15.52 314.334 15.624 318.708 ; 
        RECT 15.088 314.334 15.192 318.708 ; 
        RECT 14.656 314.334 14.76 318.708 ; 
        RECT 14.224 314.334 14.328 318.708 ; 
        RECT 13.792 314.334 13.896 318.708 ; 
        RECT 13.36 314.334 13.464 318.708 ; 
        RECT 12.928 314.334 13.032 318.708 ; 
        RECT 12.496 314.334 12.6 318.708 ; 
        RECT 12.064 314.334 12.168 318.708 ; 
        RECT 11.632 314.334 11.736 318.708 ; 
        RECT 11.2 314.334 11.304 318.708 ; 
        RECT 10.768 314.334 10.872 318.708 ; 
        RECT 10.336 314.334 10.44 318.708 ; 
        RECT 9.904 314.334 10.008 318.708 ; 
        RECT 9.472 314.334 9.576 318.708 ; 
        RECT 9.04 314.334 9.144 318.708 ; 
        RECT 8.608 314.334 8.712 318.708 ; 
        RECT 8.176 314.334 8.28 318.708 ; 
        RECT 7.744 314.334 7.848 318.708 ; 
        RECT 7.312 314.334 7.416 318.708 ; 
        RECT 6.88 314.334 6.984 318.708 ; 
        RECT 6.448 314.334 6.552 318.708 ; 
        RECT 6.016 314.334 6.12 318.708 ; 
        RECT 5.584 314.334 5.688 318.708 ; 
        RECT 5.152 314.334 5.256 318.708 ; 
        RECT 4.72 314.334 4.824 318.708 ; 
        RECT 4.288 314.334 4.392 318.708 ; 
        RECT 3.856 314.334 3.96 318.708 ; 
        RECT 3.424 314.334 3.528 318.708 ; 
        RECT 2.992 314.334 3.096 318.708 ; 
        RECT 2.56 314.334 2.664 318.708 ; 
        RECT 2.128 314.334 2.232 318.708 ; 
        RECT 1.696 314.334 1.8 318.708 ; 
        RECT 1.264 314.334 1.368 318.708 ; 
        RECT 0.832 314.334 0.936 318.708 ; 
        RECT 0.02 314.334 0.36 318.708 ; 
        RECT 34.564 318.654 35.076 323.028 ; 
        RECT 34.508 321.316 35.076 322.606 ; 
        RECT 33.916 320.224 34.164 323.028 ; 
        RECT 33.86 321.462 34.164 322.076 ; 
        RECT 33.916 318.654 34.02 323.028 ; 
        RECT 33.916 319.138 34.076 320.096 ; 
        RECT 33.916 318.654 34.164 319.01 ; 
        RECT 32.728 320.456 33.552 323.028 ; 
        RECT 33.448 318.654 33.552 323.028 ; 
        RECT 32.728 321.564 33.608 322.596 ; 
        RECT 32.728 318.654 33.12 323.028 ; 
        RECT 31.06 318.654 31.392 323.028 ; 
        RECT 31.06 319.008 31.448 322.75 ; 
        RECT 65.776 318.654 66.116 323.028 ; 
        RECT 65.2 318.654 65.304 323.028 ; 
        RECT 64.768 318.654 64.872 323.028 ; 
        RECT 64.336 318.654 64.44 323.028 ; 
        RECT 63.904 318.654 64.008 323.028 ; 
        RECT 63.472 318.654 63.576 323.028 ; 
        RECT 63.04 318.654 63.144 323.028 ; 
        RECT 62.608 318.654 62.712 323.028 ; 
        RECT 62.176 318.654 62.28 323.028 ; 
        RECT 61.744 318.654 61.848 323.028 ; 
        RECT 61.312 318.654 61.416 323.028 ; 
        RECT 60.88 318.654 60.984 323.028 ; 
        RECT 60.448 318.654 60.552 323.028 ; 
        RECT 60.016 318.654 60.12 323.028 ; 
        RECT 59.584 318.654 59.688 323.028 ; 
        RECT 59.152 318.654 59.256 323.028 ; 
        RECT 58.72 318.654 58.824 323.028 ; 
        RECT 58.288 318.654 58.392 323.028 ; 
        RECT 57.856 318.654 57.96 323.028 ; 
        RECT 57.424 318.654 57.528 323.028 ; 
        RECT 56.992 318.654 57.096 323.028 ; 
        RECT 56.56 318.654 56.664 323.028 ; 
        RECT 56.128 318.654 56.232 323.028 ; 
        RECT 55.696 318.654 55.8 323.028 ; 
        RECT 55.264 318.654 55.368 323.028 ; 
        RECT 54.832 318.654 54.936 323.028 ; 
        RECT 54.4 318.654 54.504 323.028 ; 
        RECT 53.968 318.654 54.072 323.028 ; 
        RECT 53.536 318.654 53.64 323.028 ; 
        RECT 53.104 318.654 53.208 323.028 ; 
        RECT 52.672 318.654 52.776 323.028 ; 
        RECT 52.24 318.654 52.344 323.028 ; 
        RECT 51.808 318.654 51.912 323.028 ; 
        RECT 51.376 318.654 51.48 323.028 ; 
        RECT 50.944 318.654 51.048 323.028 ; 
        RECT 50.512 318.654 50.616 323.028 ; 
        RECT 50.08 318.654 50.184 323.028 ; 
        RECT 49.648 318.654 49.752 323.028 ; 
        RECT 49.216 318.654 49.32 323.028 ; 
        RECT 48.784 318.654 48.888 323.028 ; 
        RECT 48.352 318.654 48.456 323.028 ; 
        RECT 47.92 318.654 48.024 323.028 ; 
        RECT 47.488 318.654 47.592 323.028 ; 
        RECT 47.056 318.654 47.16 323.028 ; 
        RECT 46.624 318.654 46.728 323.028 ; 
        RECT 46.192 318.654 46.296 323.028 ; 
        RECT 45.76 318.654 45.864 323.028 ; 
        RECT 45.328 318.654 45.432 323.028 ; 
        RECT 44.896 318.654 45 323.028 ; 
        RECT 44.464 318.654 44.568 323.028 ; 
        RECT 44.032 318.654 44.136 323.028 ; 
        RECT 43.6 318.654 43.704 323.028 ; 
        RECT 43.168 318.654 43.272 323.028 ; 
        RECT 42.736 318.654 42.84 323.028 ; 
        RECT 42.304 318.654 42.408 323.028 ; 
        RECT 41.872 318.654 41.976 323.028 ; 
        RECT 41.44 318.654 41.544 323.028 ; 
        RECT 41.008 318.654 41.112 323.028 ; 
        RECT 40.576 318.654 40.68 323.028 ; 
        RECT 40.144 318.654 40.248 323.028 ; 
        RECT 39.712 318.654 39.816 323.028 ; 
        RECT 39.28 318.654 39.384 323.028 ; 
        RECT 38.848 318.654 38.952 323.028 ; 
        RECT 38.416 318.654 38.52 323.028 ; 
        RECT 37.984 318.654 38.088 323.028 ; 
        RECT 37.552 318.654 37.656 323.028 ; 
        RECT 36.7 318.654 37.008 323.028 ; 
        RECT 29.128 318.654 29.436 323.028 ; 
        RECT 28.48 318.654 28.584 323.028 ; 
        RECT 28.048 318.654 28.152 323.028 ; 
        RECT 27.616 318.654 27.72 323.028 ; 
        RECT 27.184 318.654 27.288 323.028 ; 
        RECT 26.752 318.654 26.856 323.028 ; 
        RECT 26.32 318.654 26.424 323.028 ; 
        RECT 25.888 318.654 25.992 323.028 ; 
        RECT 25.456 318.654 25.56 323.028 ; 
        RECT 25.024 318.654 25.128 323.028 ; 
        RECT 24.592 318.654 24.696 323.028 ; 
        RECT 24.16 318.654 24.264 323.028 ; 
        RECT 23.728 318.654 23.832 323.028 ; 
        RECT 23.296 318.654 23.4 323.028 ; 
        RECT 22.864 318.654 22.968 323.028 ; 
        RECT 22.432 318.654 22.536 323.028 ; 
        RECT 22 318.654 22.104 323.028 ; 
        RECT 21.568 318.654 21.672 323.028 ; 
        RECT 21.136 318.654 21.24 323.028 ; 
        RECT 20.704 318.654 20.808 323.028 ; 
        RECT 20.272 318.654 20.376 323.028 ; 
        RECT 19.84 318.654 19.944 323.028 ; 
        RECT 19.408 318.654 19.512 323.028 ; 
        RECT 18.976 318.654 19.08 323.028 ; 
        RECT 18.544 318.654 18.648 323.028 ; 
        RECT 18.112 318.654 18.216 323.028 ; 
        RECT 17.68 318.654 17.784 323.028 ; 
        RECT 17.248 318.654 17.352 323.028 ; 
        RECT 16.816 318.654 16.92 323.028 ; 
        RECT 16.384 318.654 16.488 323.028 ; 
        RECT 15.952 318.654 16.056 323.028 ; 
        RECT 15.52 318.654 15.624 323.028 ; 
        RECT 15.088 318.654 15.192 323.028 ; 
        RECT 14.656 318.654 14.76 323.028 ; 
        RECT 14.224 318.654 14.328 323.028 ; 
        RECT 13.792 318.654 13.896 323.028 ; 
        RECT 13.36 318.654 13.464 323.028 ; 
        RECT 12.928 318.654 13.032 323.028 ; 
        RECT 12.496 318.654 12.6 323.028 ; 
        RECT 12.064 318.654 12.168 323.028 ; 
        RECT 11.632 318.654 11.736 323.028 ; 
        RECT 11.2 318.654 11.304 323.028 ; 
        RECT 10.768 318.654 10.872 323.028 ; 
        RECT 10.336 318.654 10.44 323.028 ; 
        RECT 9.904 318.654 10.008 323.028 ; 
        RECT 9.472 318.654 9.576 323.028 ; 
        RECT 9.04 318.654 9.144 323.028 ; 
        RECT 8.608 318.654 8.712 323.028 ; 
        RECT 8.176 318.654 8.28 323.028 ; 
        RECT 7.744 318.654 7.848 323.028 ; 
        RECT 7.312 318.654 7.416 323.028 ; 
        RECT 6.88 318.654 6.984 323.028 ; 
        RECT 6.448 318.654 6.552 323.028 ; 
        RECT 6.016 318.654 6.12 323.028 ; 
        RECT 5.584 318.654 5.688 323.028 ; 
        RECT 5.152 318.654 5.256 323.028 ; 
        RECT 4.72 318.654 4.824 323.028 ; 
        RECT 4.288 318.654 4.392 323.028 ; 
        RECT 3.856 318.654 3.96 323.028 ; 
        RECT 3.424 318.654 3.528 323.028 ; 
        RECT 2.992 318.654 3.096 323.028 ; 
        RECT 2.56 318.654 2.664 323.028 ; 
        RECT 2.128 318.654 2.232 323.028 ; 
        RECT 1.696 318.654 1.8 323.028 ; 
        RECT 1.264 318.654 1.368 323.028 ; 
        RECT 0.832 318.654 0.936 323.028 ; 
        RECT 0.02 318.654 0.36 323.028 ; 
        RECT 34.564 322.974 35.076 327.348 ; 
        RECT 34.508 325.636 35.076 326.926 ; 
        RECT 33.916 324.544 34.164 327.348 ; 
        RECT 33.86 325.782 34.164 326.396 ; 
        RECT 33.916 322.974 34.02 327.348 ; 
        RECT 33.916 323.458 34.076 324.416 ; 
        RECT 33.916 322.974 34.164 323.33 ; 
        RECT 32.728 324.776 33.552 327.348 ; 
        RECT 33.448 322.974 33.552 327.348 ; 
        RECT 32.728 325.884 33.608 326.916 ; 
        RECT 32.728 322.974 33.12 327.348 ; 
        RECT 31.06 322.974 31.392 327.348 ; 
        RECT 31.06 323.328 31.448 327.07 ; 
        RECT 65.776 322.974 66.116 327.348 ; 
        RECT 65.2 322.974 65.304 327.348 ; 
        RECT 64.768 322.974 64.872 327.348 ; 
        RECT 64.336 322.974 64.44 327.348 ; 
        RECT 63.904 322.974 64.008 327.348 ; 
        RECT 63.472 322.974 63.576 327.348 ; 
        RECT 63.04 322.974 63.144 327.348 ; 
        RECT 62.608 322.974 62.712 327.348 ; 
        RECT 62.176 322.974 62.28 327.348 ; 
        RECT 61.744 322.974 61.848 327.348 ; 
        RECT 61.312 322.974 61.416 327.348 ; 
        RECT 60.88 322.974 60.984 327.348 ; 
        RECT 60.448 322.974 60.552 327.348 ; 
        RECT 60.016 322.974 60.12 327.348 ; 
        RECT 59.584 322.974 59.688 327.348 ; 
        RECT 59.152 322.974 59.256 327.348 ; 
        RECT 58.72 322.974 58.824 327.348 ; 
        RECT 58.288 322.974 58.392 327.348 ; 
        RECT 57.856 322.974 57.96 327.348 ; 
        RECT 57.424 322.974 57.528 327.348 ; 
        RECT 56.992 322.974 57.096 327.348 ; 
        RECT 56.56 322.974 56.664 327.348 ; 
        RECT 56.128 322.974 56.232 327.348 ; 
        RECT 55.696 322.974 55.8 327.348 ; 
        RECT 55.264 322.974 55.368 327.348 ; 
        RECT 54.832 322.974 54.936 327.348 ; 
        RECT 54.4 322.974 54.504 327.348 ; 
        RECT 53.968 322.974 54.072 327.348 ; 
        RECT 53.536 322.974 53.64 327.348 ; 
        RECT 53.104 322.974 53.208 327.348 ; 
        RECT 52.672 322.974 52.776 327.348 ; 
        RECT 52.24 322.974 52.344 327.348 ; 
        RECT 51.808 322.974 51.912 327.348 ; 
        RECT 51.376 322.974 51.48 327.348 ; 
        RECT 50.944 322.974 51.048 327.348 ; 
        RECT 50.512 322.974 50.616 327.348 ; 
        RECT 50.08 322.974 50.184 327.348 ; 
        RECT 49.648 322.974 49.752 327.348 ; 
        RECT 49.216 322.974 49.32 327.348 ; 
        RECT 48.784 322.974 48.888 327.348 ; 
        RECT 48.352 322.974 48.456 327.348 ; 
        RECT 47.92 322.974 48.024 327.348 ; 
        RECT 47.488 322.974 47.592 327.348 ; 
        RECT 47.056 322.974 47.16 327.348 ; 
        RECT 46.624 322.974 46.728 327.348 ; 
        RECT 46.192 322.974 46.296 327.348 ; 
        RECT 45.76 322.974 45.864 327.348 ; 
        RECT 45.328 322.974 45.432 327.348 ; 
        RECT 44.896 322.974 45 327.348 ; 
        RECT 44.464 322.974 44.568 327.348 ; 
        RECT 44.032 322.974 44.136 327.348 ; 
        RECT 43.6 322.974 43.704 327.348 ; 
        RECT 43.168 322.974 43.272 327.348 ; 
        RECT 42.736 322.974 42.84 327.348 ; 
        RECT 42.304 322.974 42.408 327.348 ; 
        RECT 41.872 322.974 41.976 327.348 ; 
        RECT 41.44 322.974 41.544 327.348 ; 
        RECT 41.008 322.974 41.112 327.348 ; 
        RECT 40.576 322.974 40.68 327.348 ; 
        RECT 40.144 322.974 40.248 327.348 ; 
        RECT 39.712 322.974 39.816 327.348 ; 
        RECT 39.28 322.974 39.384 327.348 ; 
        RECT 38.848 322.974 38.952 327.348 ; 
        RECT 38.416 322.974 38.52 327.348 ; 
        RECT 37.984 322.974 38.088 327.348 ; 
        RECT 37.552 322.974 37.656 327.348 ; 
        RECT 36.7 322.974 37.008 327.348 ; 
        RECT 29.128 322.974 29.436 327.348 ; 
        RECT 28.48 322.974 28.584 327.348 ; 
        RECT 28.048 322.974 28.152 327.348 ; 
        RECT 27.616 322.974 27.72 327.348 ; 
        RECT 27.184 322.974 27.288 327.348 ; 
        RECT 26.752 322.974 26.856 327.348 ; 
        RECT 26.32 322.974 26.424 327.348 ; 
        RECT 25.888 322.974 25.992 327.348 ; 
        RECT 25.456 322.974 25.56 327.348 ; 
        RECT 25.024 322.974 25.128 327.348 ; 
        RECT 24.592 322.974 24.696 327.348 ; 
        RECT 24.16 322.974 24.264 327.348 ; 
        RECT 23.728 322.974 23.832 327.348 ; 
        RECT 23.296 322.974 23.4 327.348 ; 
        RECT 22.864 322.974 22.968 327.348 ; 
        RECT 22.432 322.974 22.536 327.348 ; 
        RECT 22 322.974 22.104 327.348 ; 
        RECT 21.568 322.974 21.672 327.348 ; 
        RECT 21.136 322.974 21.24 327.348 ; 
        RECT 20.704 322.974 20.808 327.348 ; 
        RECT 20.272 322.974 20.376 327.348 ; 
        RECT 19.84 322.974 19.944 327.348 ; 
        RECT 19.408 322.974 19.512 327.348 ; 
        RECT 18.976 322.974 19.08 327.348 ; 
        RECT 18.544 322.974 18.648 327.348 ; 
        RECT 18.112 322.974 18.216 327.348 ; 
        RECT 17.68 322.974 17.784 327.348 ; 
        RECT 17.248 322.974 17.352 327.348 ; 
        RECT 16.816 322.974 16.92 327.348 ; 
        RECT 16.384 322.974 16.488 327.348 ; 
        RECT 15.952 322.974 16.056 327.348 ; 
        RECT 15.52 322.974 15.624 327.348 ; 
        RECT 15.088 322.974 15.192 327.348 ; 
        RECT 14.656 322.974 14.76 327.348 ; 
        RECT 14.224 322.974 14.328 327.348 ; 
        RECT 13.792 322.974 13.896 327.348 ; 
        RECT 13.36 322.974 13.464 327.348 ; 
        RECT 12.928 322.974 13.032 327.348 ; 
        RECT 12.496 322.974 12.6 327.348 ; 
        RECT 12.064 322.974 12.168 327.348 ; 
        RECT 11.632 322.974 11.736 327.348 ; 
        RECT 11.2 322.974 11.304 327.348 ; 
        RECT 10.768 322.974 10.872 327.348 ; 
        RECT 10.336 322.974 10.44 327.348 ; 
        RECT 9.904 322.974 10.008 327.348 ; 
        RECT 9.472 322.974 9.576 327.348 ; 
        RECT 9.04 322.974 9.144 327.348 ; 
        RECT 8.608 322.974 8.712 327.348 ; 
        RECT 8.176 322.974 8.28 327.348 ; 
        RECT 7.744 322.974 7.848 327.348 ; 
        RECT 7.312 322.974 7.416 327.348 ; 
        RECT 6.88 322.974 6.984 327.348 ; 
        RECT 6.448 322.974 6.552 327.348 ; 
        RECT 6.016 322.974 6.12 327.348 ; 
        RECT 5.584 322.974 5.688 327.348 ; 
        RECT 5.152 322.974 5.256 327.348 ; 
        RECT 4.72 322.974 4.824 327.348 ; 
        RECT 4.288 322.974 4.392 327.348 ; 
        RECT 3.856 322.974 3.96 327.348 ; 
        RECT 3.424 322.974 3.528 327.348 ; 
        RECT 2.992 322.974 3.096 327.348 ; 
        RECT 2.56 322.974 2.664 327.348 ; 
        RECT 2.128 322.974 2.232 327.348 ; 
        RECT 1.696 322.974 1.8 327.348 ; 
        RECT 1.264 322.974 1.368 327.348 ; 
        RECT 0.832 322.974 0.936 327.348 ; 
        RECT 0.02 322.974 0.36 327.348 ; 
        RECT 34.564 327.294 35.076 331.668 ; 
        RECT 34.508 329.956 35.076 331.246 ; 
        RECT 33.916 328.864 34.164 331.668 ; 
        RECT 33.86 330.102 34.164 330.716 ; 
        RECT 33.916 327.294 34.02 331.668 ; 
        RECT 33.916 327.778 34.076 328.736 ; 
        RECT 33.916 327.294 34.164 327.65 ; 
        RECT 32.728 329.096 33.552 331.668 ; 
        RECT 33.448 327.294 33.552 331.668 ; 
        RECT 32.728 330.204 33.608 331.236 ; 
        RECT 32.728 327.294 33.12 331.668 ; 
        RECT 31.06 327.294 31.392 331.668 ; 
        RECT 31.06 327.648 31.448 331.39 ; 
        RECT 65.776 327.294 66.116 331.668 ; 
        RECT 65.2 327.294 65.304 331.668 ; 
        RECT 64.768 327.294 64.872 331.668 ; 
        RECT 64.336 327.294 64.44 331.668 ; 
        RECT 63.904 327.294 64.008 331.668 ; 
        RECT 63.472 327.294 63.576 331.668 ; 
        RECT 63.04 327.294 63.144 331.668 ; 
        RECT 62.608 327.294 62.712 331.668 ; 
        RECT 62.176 327.294 62.28 331.668 ; 
        RECT 61.744 327.294 61.848 331.668 ; 
        RECT 61.312 327.294 61.416 331.668 ; 
        RECT 60.88 327.294 60.984 331.668 ; 
        RECT 60.448 327.294 60.552 331.668 ; 
        RECT 60.016 327.294 60.12 331.668 ; 
        RECT 59.584 327.294 59.688 331.668 ; 
        RECT 59.152 327.294 59.256 331.668 ; 
        RECT 58.72 327.294 58.824 331.668 ; 
        RECT 58.288 327.294 58.392 331.668 ; 
        RECT 57.856 327.294 57.96 331.668 ; 
        RECT 57.424 327.294 57.528 331.668 ; 
        RECT 56.992 327.294 57.096 331.668 ; 
        RECT 56.56 327.294 56.664 331.668 ; 
        RECT 56.128 327.294 56.232 331.668 ; 
        RECT 55.696 327.294 55.8 331.668 ; 
        RECT 55.264 327.294 55.368 331.668 ; 
        RECT 54.832 327.294 54.936 331.668 ; 
        RECT 54.4 327.294 54.504 331.668 ; 
        RECT 53.968 327.294 54.072 331.668 ; 
        RECT 53.536 327.294 53.64 331.668 ; 
        RECT 53.104 327.294 53.208 331.668 ; 
        RECT 52.672 327.294 52.776 331.668 ; 
        RECT 52.24 327.294 52.344 331.668 ; 
        RECT 51.808 327.294 51.912 331.668 ; 
        RECT 51.376 327.294 51.48 331.668 ; 
        RECT 50.944 327.294 51.048 331.668 ; 
        RECT 50.512 327.294 50.616 331.668 ; 
        RECT 50.08 327.294 50.184 331.668 ; 
        RECT 49.648 327.294 49.752 331.668 ; 
        RECT 49.216 327.294 49.32 331.668 ; 
        RECT 48.784 327.294 48.888 331.668 ; 
        RECT 48.352 327.294 48.456 331.668 ; 
        RECT 47.92 327.294 48.024 331.668 ; 
        RECT 47.488 327.294 47.592 331.668 ; 
        RECT 47.056 327.294 47.16 331.668 ; 
        RECT 46.624 327.294 46.728 331.668 ; 
        RECT 46.192 327.294 46.296 331.668 ; 
        RECT 45.76 327.294 45.864 331.668 ; 
        RECT 45.328 327.294 45.432 331.668 ; 
        RECT 44.896 327.294 45 331.668 ; 
        RECT 44.464 327.294 44.568 331.668 ; 
        RECT 44.032 327.294 44.136 331.668 ; 
        RECT 43.6 327.294 43.704 331.668 ; 
        RECT 43.168 327.294 43.272 331.668 ; 
        RECT 42.736 327.294 42.84 331.668 ; 
        RECT 42.304 327.294 42.408 331.668 ; 
        RECT 41.872 327.294 41.976 331.668 ; 
        RECT 41.44 327.294 41.544 331.668 ; 
        RECT 41.008 327.294 41.112 331.668 ; 
        RECT 40.576 327.294 40.68 331.668 ; 
        RECT 40.144 327.294 40.248 331.668 ; 
        RECT 39.712 327.294 39.816 331.668 ; 
        RECT 39.28 327.294 39.384 331.668 ; 
        RECT 38.848 327.294 38.952 331.668 ; 
        RECT 38.416 327.294 38.52 331.668 ; 
        RECT 37.984 327.294 38.088 331.668 ; 
        RECT 37.552 327.294 37.656 331.668 ; 
        RECT 36.7 327.294 37.008 331.668 ; 
        RECT 29.128 327.294 29.436 331.668 ; 
        RECT 28.48 327.294 28.584 331.668 ; 
        RECT 28.048 327.294 28.152 331.668 ; 
        RECT 27.616 327.294 27.72 331.668 ; 
        RECT 27.184 327.294 27.288 331.668 ; 
        RECT 26.752 327.294 26.856 331.668 ; 
        RECT 26.32 327.294 26.424 331.668 ; 
        RECT 25.888 327.294 25.992 331.668 ; 
        RECT 25.456 327.294 25.56 331.668 ; 
        RECT 25.024 327.294 25.128 331.668 ; 
        RECT 24.592 327.294 24.696 331.668 ; 
        RECT 24.16 327.294 24.264 331.668 ; 
        RECT 23.728 327.294 23.832 331.668 ; 
        RECT 23.296 327.294 23.4 331.668 ; 
        RECT 22.864 327.294 22.968 331.668 ; 
        RECT 22.432 327.294 22.536 331.668 ; 
        RECT 22 327.294 22.104 331.668 ; 
        RECT 21.568 327.294 21.672 331.668 ; 
        RECT 21.136 327.294 21.24 331.668 ; 
        RECT 20.704 327.294 20.808 331.668 ; 
        RECT 20.272 327.294 20.376 331.668 ; 
        RECT 19.84 327.294 19.944 331.668 ; 
        RECT 19.408 327.294 19.512 331.668 ; 
        RECT 18.976 327.294 19.08 331.668 ; 
        RECT 18.544 327.294 18.648 331.668 ; 
        RECT 18.112 327.294 18.216 331.668 ; 
        RECT 17.68 327.294 17.784 331.668 ; 
        RECT 17.248 327.294 17.352 331.668 ; 
        RECT 16.816 327.294 16.92 331.668 ; 
        RECT 16.384 327.294 16.488 331.668 ; 
        RECT 15.952 327.294 16.056 331.668 ; 
        RECT 15.52 327.294 15.624 331.668 ; 
        RECT 15.088 327.294 15.192 331.668 ; 
        RECT 14.656 327.294 14.76 331.668 ; 
        RECT 14.224 327.294 14.328 331.668 ; 
        RECT 13.792 327.294 13.896 331.668 ; 
        RECT 13.36 327.294 13.464 331.668 ; 
        RECT 12.928 327.294 13.032 331.668 ; 
        RECT 12.496 327.294 12.6 331.668 ; 
        RECT 12.064 327.294 12.168 331.668 ; 
        RECT 11.632 327.294 11.736 331.668 ; 
        RECT 11.2 327.294 11.304 331.668 ; 
        RECT 10.768 327.294 10.872 331.668 ; 
        RECT 10.336 327.294 10.44 331.668 ; 
        RECT 9.904 327.294 10.008 331.668 ; 
        RECT 9.472 327.294 9.576 331.668 ; 
        RECT 9.04 327.294 9.144 331.668 ; 
        RECT 8.608 327.294 8.712 331.668 ; 
        RECT 8.176 327.294 8.28 331.668 ; 
        RECT 7.744 327.294 7.848 331.668 ; 
        RECT 7.312 327.294 7.416 331.668 ; 
        RECT 6.88 327.294 6.984 331.668 ; 
        RECT 6.448 327.294 6.552 331.668 ; 
        RECT 6.016 327.294 6.12 331.668 ; 
        RECT 5.584 327.294 5.688 331.668 ; 
        RECT 5.152 327.294 5.256 331.668 ; 
        RECT 4.72 327.294 4.824 331.668 ; 
        RECT 4.288 327.294 4.392 331.668 ; 
        RECT 3.856 327.294 3.96 331.668 ; 
        RECT 3.424 327.294 3.528 331.668 ; 
        RECT 2.992 327.294 3.096 331.668 ; 
        RECT 2.56 327.294 2.664 331.668 ; 
        RECT 2.128 327.294 2.232 331.668 ; 
        RECT 1.696 327.294 1.8 331.668 ; 
        RECT 1.264 327.294 1.368 331.668 ; 
        RECT 0.832 327.294 0.936 331.668 ; 
        RECT 0.02 327.294 0.36 331.668 ; 
        RECT 34.564 331.614 35.076 335.988 ; 
        RECT 34.508 334.276 35.076 335.566 ; 
        RECT 33.916 333.184 34.164 335.988 ; 
        RECT 33.86 334.422 34.164 335.036 ; 
        RECT 33.916 331.614 34.02 335.988 ; 
        RECT 33.916 332.098 34.076 333.056 ; 
        RECT 33.916 331.614 34.164 331.97 ; 
        RECT 32.728 333.416 33.552 335.988 ; 
        RECT 33.448 331.614 33.552 335.988 ; 
        RECT 32.728 334.524 33.608 335.556 ; 
        RECT 32.728 331.614 33.12 335.988 ; 
        RECT 31.06 331.614 31.392 335.988 ; 
        RECT 31.06 331.968 31.448 335.71 ; 
        RECT 65.776 331.614 66.116 335.988 ; 
        RECT 65.2 331.614 65.304 335.988 ; 
        RECT 64.768 331.614 64.872 335.988 ; 
        RECT 64.336 331.614 64.44 335.988 ; 
        RECT 63.904 331.614 64.008 335.988 ; 
        RECT 63.472 331.614 63.576 335.988 ; 
        RECT 63.04 331.614 63.144 335.988 ; 
        RECT 62.608 331.614 62.712 335.988 ; 
        RECT 62.176 331.614 62.28 335.988 ; 
        RECT 61.744 331.614 61.848 335.988 ; 
        RECT 61.312 331.614 61.416 335.988 ; 
        RECT 60.88 331.614 60.984 335.988 ; 
        RECT 60.448 331.614 60.552 335.988 ; 
        RECT 60.016 331.614 60.12 335.988 ; 
        RECT 59.584 331.614 59.688 335.988 ; 
        RECT 59.152 331.614 59.256 335.988 ; 
        RECT 58.72 331.614 58.824 335.988 ; 
        RECT 58.288 331.614 58.392 335.988 ; 
        RECT 57.856 331.614 57.96 335.988 ; 
        RECT 57.424 331.614 57.528 335.988 ; 
        RECT 56.992 331.614 57.096 335.988 ; 
        RECT 56.56 331.614 56.664 335.988 ; 
        RECT 56.128 331.614 56.232 335.988 ; 
        RECT 55.696 331.614 55.8 335.988 ; 
        RECT 55.264 331.614 55.368 335.988 ; 
        RECT 54.832 331.614 54.936 335.988 ; 
        RECT 54.4 331.614 54.504 335.988 ; 
        RECT 53.968 331.614 54.072 335.988 ; 
        RECT 53.536 331.614 53.64 335.988 ; 
        RECT 53.104 331.614 53.208 335.988 ; 
        RECT 52.672 331.614 52.776 335.988 ; 
        RECT 52.24 331.614 52.344 335.988 ; 
        RECT 51.808 331.614 51.912 335.988 ; 
        RECT 51.376 331.614 51.48 335.988 ; 
        RECT 50.944 331.614 51.048 335.988 ; 
        RECT 50.512 331.614 50.616 335.988 ; 
        RECT 50.08 331.614 50.184 335.988 ; 
        RECT 49.648 331.614 49.752 335.988 ; 
        RECT 49.216 331.614 49.32 335.988 ; 
        RECT 48.784 331.614 48.888 335.988 ; 
        RECT 48.352 331.614 48.456 335.988 ; 
        RECT 47.92 331.614 48.024 335.988 ; 
        RECT 47.488 331.614 47.592 335.988 ; 
        RECT 47.056 331.614 47.16 335.988 ; 
        RECT 46.624 331.614 46.728 335.988 ; 
        RECT 46.192 331.614 46.296 335.988 ; 
        RECT 45.76 331.614 45.864 335.988 ; 
        RECT 45.328 331.614 45.432 335.988 ; 
        RECT 44.896 331.614 45 335.988 ; 
        RECT 44.464 331.614 44.568 335.988 ; 
        RECT 44.032 331.614 44.136 335.988 ; 
        RECT 43.6 331.614 43.704 335.988 ; 
        RECT 43.168 331.614 43.272 335.988 ; 
        RECT 42.736 331.614 42.84 335.988 ; 
        RECT 42.304 331.614 42.408 335.988 ; 
        RECT 41.872 331.614 41.976 335.988 ; 
        RECT 41.44 331.614 41.544 335.988 ; 
        RECT 41.008 331.614 41.112 335.988 ; 
        RECT 40.576 331.614 40.68 335.988 ; 
        RECT 40.144 331.614 40.248 335.988 ; 
        RECT 39.712 331.614 39.816 335.988 ; 
        RECT 39.28 331.614 39.384 335.988 ; 
        RECT 38.848 331.614 38.952 335.988 ; 
        RECT 38.416 331.614 38.52 335.988 ; 
        RECT 37.984 331.614 38.088 335.988 ; 
        RECT 37.552 331.614 37.656 335.988 ; 
        RECT 36.7 331.614 37.008 335.988 ; 
        RECT 29.128 331.614 29.436 335.988 ; 
        RECT 28.48 331.614 28.584 335.988 ; 
        RECT 28.048 331.614 28.152 335.988 ; 
        RECT 27.616 331.614 27.72 335.988 ; 
        RECT 27.184 331.614 27.288 335.988 ; 
        RECT 26.752 331.614 26.856 335.988 ; 
        RECT 26.32 331.614 26.424 335.988 ; 
        RECT 25.888 331.614 25.992 335.988 ; 
        RECT 25.456 331.614 25.56 335.988 ; 
        RECT 25.024 331.614 25.128 335.988 ; 
        RECT 24.592 331.614 24.696 335.988 ; 
        RECT 24.16 331.614 24.264 335.988 ; 
        RECT 23.728 331.614 23.832 335.988 ; 
        RECT 23.296 331.614 23.4 335.988 ; 
        RECT 22.864 331.614 22.968 335.988 ; 
        RECT 22.432 331.614 22.536 335.988 ; 
        RECT 22 331.614 22.104 335.988 ; 
        RECT 21.568 331.614 21.672 335.988 ; 
        RECT 21.136 331.614 21.24 335.988 ; 
        RECT 20.704 331.614 20.808 335.988 ; 
        RECT 20.272 331.614 20.376 335.988 ; 
        RECT 19.84 331.614 19.944 335.988 ; 
        RECT 19.408 331.614 19.512 335.988 ; 
        RECT 18.976 331.614 19.08 335.988 ; 
        RECT 18.544 331.614 18.648 335.988 ; 
        RECT 18.112 331.614 18.216 335.988 ; 
        RECT 17.68 331.614 17.784 335.988 ; 
        RECT 17.248 331.614 17.352 335.988 ; 
        RECT 16.816 331.614 16.92 335.988 ; 
        RECT 16.384 331.614 16.488 335.988 ; 
        RECT 15.952 331.614 16.056 335.988 ; 
        RECT 15.52 331.614 15.624 335.988 ; 
        RECT 15.088 331.614 15.192 335.988 ; 
        RECT 14.656 331.614 14.76 335.988 ; 
        RECT 14.224 331.614 14.328 335.988 ; 
        RECT 13.792 331.614 13.896 335.988 ; 
        RECT 13.36 331.614 13.464 335.988 ; 
        RECT 12.928 331.614 13.032 335.988 ; 
        RECT 12.496 331.614 12.6 335.988 ; 
        RECT 12.064 331.614 12.168 335.988 ; 
        RECT 11.632 331.614 11.736 335.988 ; 
        RECT 11.2 331.614 11.304 335.988 ; 
        RECT 10.768 331.614 10.872 335.988 ; 
        RECT 10.336 331.614 10.44 335.988 ; 
        RECT 9.904 331.614 10.008 335.988 ; 
        RECT 9.472 331.614 9.576 335.988 ; 
        RECT 9.04 331.614 9.144 335.988 ; 
        RECT 8.608 331.614 8.712 335.988 ; 
        RECT 8.176 331.614 8.28 335.988 ; 
        RECT 7.744 331.614 7.848 335.988 ; 
        RECT 7.312 331.614 7.416 335.988 ; 
        RECT 6.88 331.614 6.984 335.988 ; 
        RECT 6.448 331.614 6.552 335.988 ; 
        RECT 6.016 331.614 6.12 335.988 ; 
        RECT 5.584 331.614 5.688 335.988 ; 
        RECT 5.152 331.614 5.256 335.988 ; 
        RECT 4.72 331.614 4.824 335.988 ; 
        RECT 4.288 331.614 4.392 335.988 ; 
        RECT 3.856 331.614 3.96 335.988 ; 
        RECT 3.424 331.614 3.528 335.988 ; 
        RECT 2.992 331.614 3.096 335.988 ; 
        RECT 2.56 331.614 2.664 335.988 ; 
        RECT 2.128 331.614 2.232 335.988 ; 
        RECT 1.696 331.614 1.8 335.988 ; 
        RECT 1.264 331.614 1.368 335.988 ; 
        RECT 0.832 331.614 0.936 335.988 ; 
        RECT 0.02 331.614 0.36 335.988 ; 
        RECT 34.564 335.934 35.076 340.308 ; 
        RECT 34.508 338.596 35.076 339.886 ; 
        RECT 33.916 337.504 34.164 340.308 ; 
        RECT 33.86 338.742 34.164 339.356 ; 
        RECT 33.916 335.934 34.02 340.308 ; 
        RECT 33.916 336.418 34.076 337.376 ; 
        RECT 33.916 335.934 34.164 336.29 ; 
        RECT 32.728 337.736 33.552 340.308 ; 
        RECT 33.448 335.934 33.552 340.308 ; 
        RECT 32.728 338.844 33.608 339.876 ; 
        RECT 32.728 335.934 33.12 340.308 ; 
        RECT 31.06 335.934 31.392 340.308 ; 
        RECT 31.06 336.288 31.448 340.03 ; 
        RECT 65.776 335.934 66.116 340.308 ; 
        RECT 65.2 335.934 65.304 340.308 ; 
        RECT 64.768 335.934 64.872 340.308 ; 
        RECT 64.336 335.934 64.44 340.308 ; 
        RECT 63.904 335.934 64.008 340.308 ; 
        RECT 63.472 335.934 63.576 340.308 ; 
        RECT 63.04 335.934 63.144 340.308 ; 
        RECT 62.608 335.934 62.712 340.308 ; 
        RECT 62.176 335.934 62.28 340.308 ; 
        RECT 61.744 335.934 61.848 340.308 ; 
        RECT 61.312 335.934 61.416 340.308 ; 
        RECT 60.88 335.934 60.984 340.308 ; 
        RECT 60.448 335.934 60.552 340.308 ; 
        RECT 60.016 335.934 60.12 340.308 ; 
        RECT 59.584 335.934 59.688 340.308 ; 
        RECT 59.152 335.934 59.256 340.308 ; 
        RECT 58.72 335.934 58.824 340.308 ; 
        RECT 58.288 335.934 58.392 340.308 ; 
        RECT 57.856 335.934 57.96 340.308 ; 
        RECT 57.424 335.934 57.528 340.308 ; 
        RECT 56.992 335.934 57.096 340.308 ; 
        RECT 56.56 335.934 56.664 340.308 ; 
        RECT 56.128 335.934 56.232 340.308 ; 
        RECT 55.696 335.934 55.8 340.308 ; 
        RECT 55.264 335.934 55.368 340.308 ; 
        RECT 54.832 335.934 54.936 340.308 ; 
        RECT 54.4 335.934 54.504 340.308 ; 
        RECT 53.968 335.934 54.072 340.308 ; 
        RECT 53.536 335.934 53.64 340.308 ; 
        RECT 53.104 335.934 53.208 340.308 ; 
        RECT 52.672 335.934 52.776 340.308 ; 
        RECT 52.24 335.934 52.344 340.308 ; 
        RECT 51.808 335.934 51.912 340.308 ; 
        RECT 51.376 335.934 51.48 340.308 ; 
        RECT 50.944 335.934 51.048 340.308 ; 
        RECT 50.512 335.934 50.616 340.308 ; 
        RECT 50.08 335.934 50.184 340.308 ; 
        RECT 49.648 335.934 49.752 340.308 ; 
        RECT 49.216 335.934 49.32 340.308 ; 
        RECT 48.784 335.934 48.888 340.308 ; 
        RECT 48.352 335.934 48.456 340.308 ; 
        RECT 47.92 335.934 48.024 340.308 ; 
        RECT 47.488 335.934 47.592 340.308 ; 
        RECT 47.056 335.934 47.16 340.308 ; 
        RECT 46.624 335.934 46.728 340.308 ; 
        RECT 46.192 335.934 46.296 340.308 ; 
        RECT 45.76 335.934 45.864 340.308 ; 
        RECT 45.328 335.934 45.432 340.308 ; 
        RECT 44.896 335.934 45 340.308 ; 
        RECT 44.464 335.934 44.568 340.308 ; 
        RECT 44.032 335.934 44.136 340.308 ; 
        RECT 43.6 335.934 43.704 340.308 ; 
        RECT 43.168 335.934 43.272 340.308 ; 
        RECT 42.736 335.934 42.84 340.308 ; 
        RECT 42.304 335.934 42.408 340.308 ; 
        RECT 41.872 335.934 41.976 340.308 ; 
        RECT 41.44 335.934 41.544 340.308 ; 
        RECT 41.008 335.934 41.112 340.308 ; 
        RECT 40.576 335.934 40.68 340.308 ; 
        RECT 40.144 335.934 40.248 340.308 ; 
        RECT 39.712 335.934 39.816 340.308 ; 
        RECT 39.28 335.934 39.384 340.308 ; 
        RECT 38.848 335.934 38.952 340.308 ; 
        RECT 38.416 335.934 38.52 340.308 ; 
        RECT 37.984 335.934 38.088 340.308 ; 
        RECT 37.552 335.934 37.656 340.308 ; 
        RECT 36.7 335.934 37.008 340.308 ; 
        RECT 29.128 335.934 29.436 340.308 ; 
        RECT 28.48 335.934 28.584 340.308 ; 
        RECT 28.048 335.934 28.152 340.308 ; 
        RECT 27.616 335.934 27.72 340.308 ; 
        RECT 27.184 335.934 27.288 340.308 ; 
        RECT 26.752 335.934 26.856 340.308 ; 
        RECT 26.32 335.934 26.424 340.308 ; 
        RECT 25.888 335.934 25.992 340.308 ; 
        RECT 25.456 335.934 25.56 340.308 ; 
        RECT 25.024 335.934 25.128 340.308 ; 
        RECT 24.592 335.934 24.696 340.308 ; 
        RECT 24.16 335.934 24.264 340.308 ; 
        RECT 23.728 335.934 23.832 340.308 ; 
        RECT 23.296 335.934 23.4 340.308 ; 
        RECT 22.864 335.934 22.968 340.308 ; 
        RECT 22.432 335.934 22.536 340.308 ; 
        RECT 22 335.934 22.104 340.308 ; 
        RECT 21.568 335.934 21.672 340.308 ; 
        RECT 21.136 335.934 21.24 340.308 ; 
        RECT 20.704 335.934 20.808 340.308 ; 
        RECT 20.272 335.934 20.376 340.308 ; 
        RECT 19.84 335.934 19.944 340.308 ; 
        RECT 19.408 335.934 19.512 340.308 ; 
        RECT 18.976 335.934 19.08 340.308 ; 
        RECT 18.544 335.934 18.648 340.308 ; 
        RECT 18.112 335.934 18.216 340.308 ; 
        RECT 17.68 335.934 17.784 340.308 ; 
        RECT 17.248 335.934 17.352 340.308 ; 
        RECT 16.816 335.934 16.92 340.308 ; 
        RECT 16.384 335.934 16.488 340.308 ; 
        RECT 15.952 335.934 16.056 340.308 ; 
        RECT 15.52 335.934 15.624 340.308 ; 
        RECT 15.088 335.934 15.192 340.308 ; 
        RECT 14.656 335.934 14.76 340.308 ; 
        RECT 14.224 335.934 14.328 340.308 ; 
        RECT 13.792 335.934 13.896 340.308 ; 
        RECT 13.36 335.934 13.464 340.308 ; 
        RECT 12.928 335.934 13.032 340.308 ; 
        RECT 12.496 335.934 12.6 340.308 ; 
        RECT 12.064 335.934 12.168 340.308 ; 
        RECT 11.632 335.934 11.736 340.308 ; 
        RECT 11.2 335.934 11.304 340.308 ; 
        RECT 10.768 335.934 10.872 340.308 ; 
        RECT 10.336 335.934 10.44 340.308 ; 
        RECT 9.904 335.934 10.008 340.308 ; 
        RECT 9.472 335.934 9.576 340.308 ; 
        RECT 9.04 335.934 9.144 340.308 ; 
        RECT 8.608 335.934 8.712 340.308 ; 
        RECT 8.176 335.934 8.28 340.308 ; 
        RECT 7.744 335.934 7.848 340.308 ; 
        RECT 7.312 335.934 7.416 340.308 ; 
        RECT 6.88 335.934 6.984 340.308 ; 
        RECT 6.448 335.934 6.552 340.308 ; 
        RECT 6.016 335.934 6.12 340.308 ; 
        RECT 5.584 335.934 5.688 340.308 ; 
        RECT 5.152 335.934 5.256 340.308 ; 
        RECT 4.72 335.934 4.824 340.308 ; 
        RECT 4.288 335.934 4.392 340.308 ; 
        RECT 3.856 335.934 3.96 340.308 ; 
        RECT 3.424 335.934 3.528 340.308 ; 
        RECT 2.992 335.934 3.096 340.308 ; 
        RECT 2.56 335.934 2.664 340.308 ; 
        RECT 2.128 335.934 2.232 340.308 ; 
        RECT 1.696 335.934 1.8 340.308 ; 
        RECT 1.264 335.934 1.368 340.308 ; 
        RECT 0.832 335.934 0.936 340.308 ; 
        RECT 0.02 335.934 0.36 340.308 ; 
        RECT 34.564 340.254 35.076 344.628 ; 
        RECT 34.508 342.916 35.076 344.206 ; 
        RECT 33.916 341.824 34.164 344.628 ; 
        RECT 33.86 343.062 34.164 343.676 ; 
        RECT 33.916 340.254 34.02 344.628 ; 
        RECT 33.916 340.738 34.076 341.696 ; 
        RECT 33.916 340.254 34.164 340.61 ; 
        RECT 32.728 342.056 33.552 344.628 ; 
        RECT 33.448 340.254 33.552 344.628 ; 
        RECT 32.728 343.164 33.608 344.196 ; 
        RECT 32.728 340.254 33.12 344.628 ; 
        RECT 31.06 340.254 31.392 344.628 ; 
        RECT 31.06 340.608 31.448 344.35 ; 
        RECT 65.776 340.254 66.116 344.628 ; 
        RECT 65.2 340.254 65.304 344.628 ; 
        RECT 64.768 340.254 64.872 344.628 ; 
        RECT 64.336 340.254 64.44 344.628 ; 
        RECT 63.904 340.254 64.008 344.628 ; 
        RECT 63.472 340.254 63.576 344.628 ; 
        RECT 63.04 340.254 63.144 344.628 ; 
        RECT 62.608 340.254 62.712 344.628 ; 
        RECT 62.176 340.254 62.28 344.628 ; 
        RECT 61.744 340.254 61.848 344.628 ; 
        RECT 61.312 340.254 61.416 344.628 ; 
        RECT 60.88 340.254 60.984 344.628 ; 
        RECT 60.448 340.254 60.552 344.628 ; 
        RECT 60.016 340.254 60.12 344.628 ; 
        RECT 59.584 340.254 59.688 344.628 ; 
        RECT 59.152 340.254 59.256 344.628 ; 
        RECT 58.72 340.254 58.824 344.628 ; 
        RECT 58.288 340.254 58.392 344.628 ; 
        RECT 57.856 340.254 57.96 344.628 ; 
        RECT 57.424 340.254 57.528 344.628 ; 
        RECT 56.992 340.254 57.096 344.628 ; 
        RECT 56.56 340.254 56.664 344.628 ; 
        RECT 56.128 340.254 56.232 344.628 ; 
        RECT 55.696 340.254 55.8 344.628 ; 
        RECT 55.264 340.254 55.368 344.628 ; 
        RECT 54.832 340.254 54.936 344.628 ; 
        RECT 54.4 340.254 54.504 344.628 ; 
        RECT 53.968 340.254 54.072 344.628 ; 
        RECT 53.536 340.254 53.64 344.628 ; 
        RECT 53.104 340.254 53.208 344.628 ; 
        RECT 52.672 340.254 52.776 344.628 ; 
        RECT 52.24 340.254 52.344 344.628 ; 
        RECT 51.808 340.254 51.912 344.628 ; 
        RECT 51.376 340.254 51.48 344.628 ; 
        RECT 50.944 340.254 51.048 344.628 ; 
        RECT 50.512 340.254 50.616 344.628 ; 
        RECT 50.08 340.254 50.184 344.628 ; 
        RECT 49.648 340.254 49.752 344.628 ; 
        RECT 49.216 340.254 49.32 344.628 ; 
        RECT 48.784 340.254 48.888 344.628 ; 
        RECT 48.352 340.254 48.456 344.628 ; 
        RECT 47.92 340.254 48.024 344.628 ; 
        RECT 47.488 340.254 47.592 344.628 ; 
        RECT 47.056 340.254 47.16 344.628 ; 
        RECT 46.624 340.254 46.728 344.628 ; 
        RECT 46.192 340.254 46.296 344.628 ; 
        RECT 45.76 340.254 45.864 344.628 ; 
        RECT 45.328 340.254 45.432 344.628 ; 
        RECT 44.896 340.254 45 344.628 ; 
        RECT 44.464 340.254 44.568 344.628 ; 
        RECT 44.032 340.254 44.136 344.628 ; 
        RECT 43.6 340.254 43.704 344.628 ; 
        RECT 43.168 340.254 43.272 344.628 ; 
        RECT 42.736 340.254 42.84 344.628 ; 
        RECT 42.304 340.254 42.408 344.628 ; 
        RECT 41.872 340.254 41.976 344.628 ; 
        RECT 41.44 340.254 41.544 344.628 ; 
        RECT 41.008 340.254 41.112 344.628 ; 
        RECT 40.576 340.254 40.68 344.628 ; 
        RECT 40.144 340.254 40.248 344.628 ; 
        RECT 39.712 340.254 39.816 344.628 ; 
        RECT 39.28 340.254 39.384 344.628 ; 
        RECT 38.848 340.254 38.952 344.628 ; 
        RECT 38.416 340.254 38.52 344.628 ; 
        RECT 37.984 340.254 38.088 344.628 ; 
        RECT 37.552 340.254 37.656 344.628 ; 
        RECT 36.7 340.254 37.008 344.628 ; 
        RECT 29.128 340.254 29.436 344.628 ; 
        RECT 28.48 340.254 28.584 344.628 ; 
        RECT 28.048 340.254 28.152 344.628 ; 
        RECT 27.616 340.254 27.72 344.628 ; 
        RECT 27.184 340.254 27.288 344.628 ; 
        RECT 26.752 340.254 26.856 344.628 ; 
        RECT 26.32 340.254 26.424 344.628 ; 
        RECT 25.888 340.254 25.992 344.628 ; 
        RECT 25.456 340.254 25.56 344.628 ; 
        RECT 25.024 340.254 25.128 344.628 ; 
        RECT 24.592 340.254 24.696 344.628 ; 
        RECT 24.16 340.254 24.264 344.628 ; 
        RECT 23.728 340.254 23.832 344.628 ; 
        RECT 23.296 340.254 23.4 344.628 ; 
        RECT 22.864 340.254 22.968 344.628 ; 
        RECT 22.432 340.254 22.536 344.628 ; 
        RECT 22 340.254 22.104 344.628 ; 
        RECT 21.568 340.254 21.672 344.628 ; 
        RECT 21.136 340.254 21.24 344.628 ; 
        RECT 20.704 340.254 20.808 344.628 ; 
        RECT 20.272 340.254 20.376 344.628 ; 
        RECT 19.84 340.254 19.944 344.628 ; 
        RECT 19.408 340.254 19.512 344.628 ; 
        RECT 18.976 340.254 19.08 344.628 ; 
        RECT 18.544 340.254 18.648 344.628 ; 
        RECT 18.112 340.254 18.216 344.628 ; 
        RECT 17.68 340.254 17.784 344.628 ; 
        RECT 17.248 340.254 17.352 344.628 ; 
        RECT 16.816 340.254 16.92 344.628 ; 
        RECT 16.384 340.254 16.488 344.628 ; 
        RECT 15.952 340.254 16.056 344.628 ; 
        RECT 15.52 340.254 15.624 344.628 ; 
        RECT 15.088 340.254 15.192 344.628 ; 
        RECT 14.656 340.254 14.76 344.628 ; 
        RECT 14.224 340.254 14.328 344.628 ; 
        RECT 13.792 340.254 13.896 344.628 ; 
        RECT 13.36 340.254 13.464 344.628 ; 
        RECT 12.928 340.254 13.032 344.628 ; 
        RECT 12.496 340.254 12.6 344.628 ; 
        RECT 12.064 340.254 12.168 344.628 ; 
        RECT 11.632 340.254 11.736 344.628 ; 
        RECT 11.2 340.254 11.304 344.628 ; 
        RECT 10.768 340.254 10.872 344.628 ; 
        RECT 10.336 340.254 10.44 344.628 ; 
        RECT 9.904 340.254 10.008 344.628 ; 
        RECT 9.472 340.254 9.576 344.628 ; 
        RECT 9.04 340.254 9.144 344.628 ; 
        RECT 8.608 340.254 8.712 344.628 ; 
        RECT 8.176 340.254 8.28 344.628 ; 
        RECT 7.744 340.254 7.848 344.628 ; 
        RECT 7.312 340.254 7.416 344.628 ; 
        RECT 6.88 340.254 6.984 344.628 ; 
        RECT 6.448 340.254 6.552 344.628 ; 
        RECT 6.016 340.254 6.12 344.628 ; 
        RECT 5.584 340.254 5.688 344.628 ; 
        RECT 5.152 340.254 5.256 344.628 ; 
        RECT 4.72 340.254 4.824 344.628 ; 
        RECT 4.288 340.254 4.392 344.628 ; 
        RECT 3.856 340.254 3.96 344.628 ; 
        RECT 3.424 340.254 3.528 344.628 ; 
        RECT 2.992 340.254 3.096 344.628 ; 
        RECT 2.56 340.254 2.664 344.628 ; 
        RECT 2.128 340.254 2.232 344.628 ; 
        RECT 1.696 340.254 1.8 344.628 ; 
        RECT 1.264 340.254 1.368 344.628 ; 
        RECT 0.832 340.254 0.936 344.628 ; 
        RECT 0.02 340.254 0.36 344.628 ; 
        RECT 34.564 344.574 35.076 348.948 ; 
        RECT 34.508 347.236 35.076 348.526 ; 
        RECT 33.916 346.144 34.164 348.948 ; 
        RECT 33.86 347.382 34.164 347.996 ; 
        RECT 33.916 344.574 34.02 348.948 ; 
        RECT 33.916 345.058 34.076 346.016 ; 
        RECT 33.916 344.574 34.164 344.93 ; 
        RECT 32.728 346.376 33.552 348.948 ; 
        RECT 33.448 344.574 33.552 348.948 ; 
        RECT 32.728 347.484 33.608 348.516 ; 
        RECT 32.728 344.574 33.12 348.948 ; 
        RECT 31.06 344.574 31.392 348.948 ; 
        RECT 31.06 344.928 31.448 348.67 ; 
        RECT 65.776 344.574 66.116 348.948 ; 
        RECT 65.2 344.574 65.304 348.948 ; 
        RECT 64.768 344.574 64.872 348.948 ; 
        RECT 64.336 344.574 64.44 348.948 ; 
        RECT 63.904 344.574 64.008 348.948 ; 
        RECT 63.472 344.574 63.576 348.948 ; 
        RECT 63.04 344.574 63.144 348.948 ; 
        RECT 62.608 344.574 62.712 348.948 ; 
        RECT 62.176 344.574 62.28 348.948 ; 
        RECT 61.744 344.574 61.848 348.948 ; 
        RECT 61.312 344.574 61.416 348.948 ; 
        RECT 60.88 344.574 60.984 348.948 ; 
        RECT 60.448 344.574 60.552 348.948 ; 
        RECT 60.016 344.574 60.12 348.948 ; 
        RECT 59.584 344.574 59.688 348.948 ; 
        RECT 59.152 344.574 59.256 348.948 ; 
        RECT 58.72 344.574 58.824 348.948 ; 
        RECT 58.288 344.574 58.392 348.948 ; 
        RECT 57.856 344.574 57.96 348.948 ; 
        RECT 57.424 344.574 57.528 348.948 ; 
        RECT 56.992 344.574 57.096 348.948 ; 
        RECT 56.56 344.574 56.664 348.948 ; 
        RECT 56.128 344.574 56.232 348.948 ; 
        RECT 55.696 344.574 55.8 348.948 ; 
        RECT 55.264 344.574 55.368 348.948 ; 
        RECT 54.832 344.574 54.936 348.948 ; 
        RECT 54.4 344.574 54.504 348.948 ; 
        RECT 53.968 344.574 54.072 348.948 ; 
        RECT 53.536 344.574 53.64 348.948 ; 
        RECT 53.104 344.574 53.208 348.948 ; 
        RECT 52.672 344.574 52.776 348.948 ; 
        RECT 52.24 344.574 52.344 348.948 ; 
        RECT 51.808 344.574 51.912 348.948 ; 
        RECT 51.376 344.574 51.48 348.948 ; 
        RECT 50.944 344.574 51.048 348.948 ; 
        RECT 50.512 344.574 50.616 348.948 ; 
        RECT 50.08 344.574 50.184 348.948 ; 
        RECT 49.648 344.574 49.752 348.948 ; 
        RECT 49.216 344.574 49.32 348.948 ; 
        RECT 48.784 344.574 48.888 348.948 ; 
        RECT 48.352 344.574 48.456 348.948 ; 
        RECT 47.92 344.574 48.024 348.948 ; 
        RECT 47.488 344.574 47.592 348.948 ; 
        RECT 47.056 344.574 47.16 348.948 ; 
        RECT 46.624 344.574 46.728 348.948 ; 
        RECT 46.192 344.574 46.296 348.948 ; 
        RECT 45.76 344.574 45.864 348.948 ; 
        RECT 45.328 344.574 45.432 348.948 ; 
        RECT 44.896 344.574 45 348.948 ; 
        RECT 44.464 344.574 44.568 348.948 ; 
        RECT 44.032 344.574 44.136 348.948 ; 
        RECT 43.6 344.574 43.704 348.948 ; 
        RECT 43.168 344.574 43.272 348.948 ; 
        RECT 42.736 344.574 42.84 348.948 ; 
        RECT 42.304 344.574 42.408 348.948 ; 
        RECT 41.872 344.574 41.976 348.948 ; 
        RECT 41.44 344.574 41.544 348.948 ; 
        RECT 41.008 344.574 41.112 348.948 ; 
        RECT 40.576 344.574 40.68 348.948 ; 
        RECT 40.144 344.574 40.248 348.948 ; 
        RECT 39.712 344.574 39.816 348.948 ; 
        RECT 39.28 344.574 39.384 348.948 ; 
        RECT 38.848 344.574 38.952 348.948 ; 
        RECT 38.416 344.574 38.52 348.948 ; 
        RECT 37.984 344.574 38.088 348.948 ; 
        RECT 37.552 344.574 37.656 348.948 ; 
        RECT 36.7 344.574 37.008 348.948 ; 
        RECT 29.128 344.574 29.436 348.948 ; 
        RECT 28.48 344.574 28.584 348.948 ; 
        RECT 28.048 344.574 28.152 348.948 ; 
        RECT 27.616 344.574 27.72 348.948 ; 
        RECT 27.184 344.574 27.288 348.948 ; 
        RECT 26.752 344.574 26.856 348.948 ; 
        RECT 26.32 344.574 26.424 348.948 ; 
        RECT 25.888 344.574 25.992 348.948 ; 
        RECT 25.456 344.574 25.56 348.948 ; 
        RECT 25.024 344.574 25.128 348.948 ; 
        RECT 24.592 344.574 24.696 348.948 ; 
        RECT 24.16 344.574 24.264 348.948 ; 
        RECT 23.728 344.574 23.832 348.948 ; 
        RECT 23.296 344.574 23.4 348.948 ; 
        RECT 22.864 344.574 22.968 348.948 ; 
        RECT 22.432 344.574 22.536 348.948 ; 
        RECT 22 344.574 22.104 348.948 ; 
        RECT 21.568 344.574 21.672 348.948 ; 
        RECT 21.136 344.574 21.24 348.948 ; 
        RECT 20.704 344.574 20.808 348.948 ; 
        RECT 20.272 344.574 20.376 348.948 ; 
        RECT 19.84 344.574 19.944 348.948 ; 
        RECT 19.408 344.574 19.512 348.948 ; 
        RECT 18.976 344.574 19.08 348.948 ; 
        RECT 18.544 344.574 18.648 348.948 ; 
        RECT 18.112 344.574 18.216 348.948 ; 
        RECT 17.68 344.574 17.784 348.948 ; 
        RECT 17.248 344.574 17.352 348.948 ; 
        RECT 16.816 344.574 16.92 348.948 ; 
        RECT 16.384 344.574 16.488 348.948 ; 
        RECT 15.952 344.574 16.056 348.948 ; 
        RECT 15.52 344.574 15.624 348.948 ; 
        RECT 15.088 344.574 15.192 348.948 ; 
        RECT 14.656 344.574 14.76 348.948 ; 
        RECT 14.224 344.574 14.328 348.948 ; 
        RECT 13.792 344.574 13.896 348.948 ; 
        RECT 13.36 344.574 13.464 348.948 ; 
        RECT 12.928 344.574 13.032 348.948 ; 
        RECT 12.496 344.574 12.6 348.948 ; 
        RECT 12.064 344.574 12.168 348.948 ; 
        RECT 11.632 344.574 11.736 348.948 ; 
        RECT 11.2 344.574 11.304 348.948 ; 
        RECT 10.768 344.574 10.872 348.948 ; 
        RECT 10.336 344.574 10.44 348.948 ; 
        RECT 9.904 344.574 10.008 348.948 ; 
        RECT 9.472 344.574 9.576 348.948 ; 
        RECT 9.04 344.574 9.144 348.948 ; 
        RECT 8.608 344.574 8.712 348.948 ; 
        RECT 8.176 344.574 8.28 348.948 ; 
        RECT 7.744 344.574 7.848 348.948 ; 
        RECT 7.312 344.574 7.416 348.948 ; 
        RECT 6.88 344.574 6.984 348.948 ; 
        RECT 6.448 344.574 6.552 348.948 ; 
        RECT 6.016 344.574 6.12 348.948 ; 
        RECT 5.584 344.574 5.688 348.948 ; 
        RECT 5.152 344.574 5.256 348.948 ; 
        RECT 4.72 344.574 4.824 348.948 ; 
        RECT 4.288 344.574 4.392 348.948 ; 
        RECT 3.856 344.574 3.96 348.948 ; 
        RECT 3.424 344.574 3.528 348.948 ; 
        RECT 2.992 344.574 3.096 348.948 ; 
        RECT 2.56 344.574 2.664 348.948 ; 
        RECT 2.128 344.574 2.232 348.948 ; 
        RECT 1.696 344.574 1.8 348.948 ; 
        RECT 1.264 344.574 1.368 348.948 ; 
        RECT 0.832 344.574 0.936 348.948 ; 
        RECT 0.02 344.574 0.36 348.948 ; 
        RECT 34.564 348.894 35.076 353.268 ; 
        RECT 34.508 351.556 35.076 352.846 ; 
        RECT 33.916 350.464 34.164 353.268 ; 
        RECT 33.86 351.702 34.164 352.316 ; 
        RECT 33.916 348.894 34.02 353.268 ; 
        RECT 33.916 349.378 34.076 350.336 ; 
        RECT 33.916 348.894 34.164 349.25 ; 
        RECT 32.728 350.696 33.552 353.268 ; 
        RECT 33.448 348.894 33.552 353.268 ; 
        RECT 32.728 351.804 33.608 352.836 ; 
        RECT 32.728 348.894 33.12 353.268 ; 
        RECT 31.06 348.894 31.392 353.268 ; 
        RECT 31.06 349.248 31.448 352.99 ; 
        RECT 65.776 348.894 66.116 353.268 ; 
        RECT 65.2 348.894 65.304 353.268 ; 
        RECT 64.768 348.894 64.872 353.268 ; 
        RECT 64.336 348.894 64.44 353.268 ; 
        RECT 63.904 348.894 64.008 353.268 ; 
        RECT 63.472 348.894 63.576 353.268 ; 
        RECT 63.04 348.894 63.144 353.268 ; 
        RECT 62.608 348.894 62.712 353.268 ; 
        RECT 62.176 348.894 62.28 353.268 ; 
        RECT 61.744 348.894 61.848 353.268 ; 
        RECT 61.312 348.894 61.416 353.268 ; 
        RECT 60.88 348.894 60.984 353.268 ; 
        RECT 60.448 348.894 60.552 353.268 ; 
        RECT 60.016 348.894 60.12 353.268 ; 
        RECT 59.584 348.894 59.688 353.268 ; 
        RECT 59.152 348.894 59.256 353.268 ; 
        RECT 58.72 348.894 58.824 353.268 ; 
        RECT 58.288 348.894 58.392 353.268 ; 
        RECT 57.856 348.894 57.96 353.268 ; 
        RECT 57.424 348.894 57.528 353.268 ; 
        RECT 56.992 348.894 57.096 353.268 ; 
        RECT 56.56 348.894 56.664 353.268 ; 
        RECT 56.128 348.894 56.232 353.268 ; 
        RECT 55.696 348.894 55.8 353.268 ; 
        RECT 55.264 348.894 55.368 353.268 ; 
        RECT 54.832 348.894 54.936 353.268 ; 
        RECT 54.4 348.894 54.504 353.268 ; 
        RECT 53.968 348.894 54.072 353.268 ; 
        RECT 53.536 348.894 53.64 353.268 ; 
        RECT 53.104 348.894 53.208 353.268 ; 
        RECT 52.672 348.894 52.776 353.268 ; 
        RECT 52.24 348.894 52.344 353.268 ; 
        RECT 51.808 348.894 51.912 353.268 ; 
        RECT 51.376 348.894 51.48 353.268 ; 
        RECT 50.944 348.894 51.048 353.268 ; 
        RECT 50.512 348.894 50.616 353.268 ; 
        RECT 50.08 348.894 50.184 353.268 ; 
        RECT 49.648 348.894 49.752 353.268 ; 
        RECT 49.216 348.894 49.32 353.268 ; 
        RECT 48.784 348.894 48.888 353.268 ; 
        RECT 48.352 348.894 48.456 353.268 ; 
        RECT 47.92 348.894 48.024 353.268 ; 
        RECT 47.488 348.894 47.592 353.268 ; 
        RECT 47.056 348.894 47.16 353.268 ; 
        RECT 46.624 348.894 46.728 353.268 ; 
        RECT 46.192 348.894 46.296 353.268 ; 
        RECT 45.76 348.894 45.864 353.268 ; 
        RECT 45.328 348.894 45.432 353.268 ; 
        RECT 44.896 348.894 45 353.268 ; 
        RECT 44.464 348.894 44.568 353.268 ; 
        RECT 44.032 348.894 44.136 353.268 ; 
        RECT 43.6 348.894 43.704 353.268 ; 
        RECT 43.168 348.894 43.272 353.268 ; 
        RECT 42.736 348.894 42.84 353.268 ; 
        RECT 42.304 348.894 42.408 353.268 ; 
        RECT 41.872 348.894 41.976 353.268 ; 
        RECT 41.44 348.894 41.544 353.268 ; 
        RECT 41.008 348.894 41.112 353.268 ; 
        RECT 40.576 348.894 40.68 353.268 ; 
        RECT 40.144 348.894 40.248 353.268 ; 
        RECT 39.712 348.894 39.816 353.268 ; 
        RECT 39.28 348.894 39.384 353.268 ; 
        RECT 38.848 348.894 38.952 353.268 ; 
        RECT 38.416 348.894 38.52 353.268 ; 
        RECT 37.984 348.894 38.088 353.268 ; 
        RECT 37.552 348.894 37.656 353.268 ; 
        RECT 36.7 348.894 37.008 353.268 ; 
        RECT 29.128 348.894 29.436 353.268 ; 
        RECT 28.48 348.894 28.584 353.268 ; 
        RECT 28.048 348.894 28.152 353.268 ; 
        RECT 27.616 348.894 27.72 353.268 ; 
        RECT 27.184 348.894 27.288 353.268 ; 
        RECT 26.752 348.894 26.856 353.268 ; 
        RECT 26.32 348.894 26.424 353.268 ; 
        RECT 25.888 348.894 25.992 353.268 ; 
        RECT 25.456 348.894 25.56 353.268 ; 
        RECT 25.024 348.894 25.128 353.268 ; 
        RECT 24.592 348.894 24.696 353.268 ; 
        RECT 24.16 348.894 24.264 353.268 ; 
        RECT 23.728 348.894 23.832 353.268 ; 
        RECT 23.296 348.894 23.4 353.268 ; 
        RECT 22.864 348.894 22.968 353.268 ; 
        RECT 22.432 348.894 22.536 353.268 ; 
        RECT 22 348.894 22.104 353.268 ; 
        RECT 21.568 348.894 21.672 353.268 ; 
        RECT 21.136 348.894 21.24 353.268 ; 
        RECT 20.704 348.894 20.808 353.268 ; 
        RECT 20.272 348.894 20.376 353.268 ; 
        RECT 19.84 348.894 19.944 353.268 ; 
        RECT 19.408 348.894 19.512 353.268 ; 
        RECT 18.976 348.894 19.08 353.268 ; 
        RECT 18.544 348.894 18.648 353.268 ; 
        RECT 18.112 348.894 18.216 353.268 ; 
        RECT 17.68 348.894 17.784 353.268 ; 
        RECT 17.248 348.894 17.352 353.268 ; 
        RECT 16.816 348.894 16.92 353.268 ; 
        RECT 16.384 348.894 16.488 353.268 ; 
        RECT 15.952 348.894 16.056 353.268 ; 
        RECT 15.52 348.894 15.624 353.268 ; 
        RECT 15.088 348.894 15.192 353.268 ; 
        RECT 14.656 348.894 14.76 353.268 ; 
        RECT 14.224 348.894 14.328 353.268 ; 
        RECT 13.792 348.894 13.896 353.268 ; 
        RECT 13.36 348.894 13.464 353.268 ; 
        RECT 12.928 348.894 13.032 353.268 ; 
        RECT 12.496 348.894 12.6 353.268 ; 
        RECT 12.064 348.894 12.168 353.268 ; 
        RECT 11.632 348.894 11.736 353.268 ; 
        RECT 11.2 348.894 11.304 353.268 ; 
        RECT 10.768 348.894 10.872 353.268 ; 
        RECT 10.336 348.894 10.44 353.268 ; 
        RECT 9.904 348.894 10.008 353.268 ; 
        RECT 9.472 348.894 9.576 353.268 ; 
        RECT 9.04 348.894 9.144 353.268 ; 
        RECT 8.608 348.894 8.712 353.268 ; 
        RECT 8.176 348.894 8.28 353.268 ; 
        RECT 7.744 348.894 7.848 353.268 ; 
        RECT 7.312 348.894 7.416 353.268 ; 
        RECT 6.88 348.894 6.984 353.268 ; 
        RECT 6.448 348.894 6.552 353.268 ; 
        RECT 6.016 348.894 6.12 353.268 ; 
        RECT 5.584 348.894 5.688 353.268 ; 
        RECT 5.152 348.894 5.256 353.268 ; 
        RECT 4.72 348.894 4.824 353.268 ; 
        RECT 4.288 348.894 4.392 353.268 ; 
        RECT 3.856 348.894 3.96 353.268 ; 
        RECT 3.424 348.894 3.528 353.268 ; 
        RECT 2.992 348.894 3.096 353.268 ; 
        RECT 2.56 348.894 2.664 353.268 ; 
        RECT 2.128 348.894 2.232 353.268 ; 
        RECT 1.696 348.894 1.8 353.268 ; 
        RECT 1.264 348.894 1.368 353.268 ; 
        RECT 0.832 348.894 0.936 353.268 ; 
        RECT 0.02 348.894 0.36 353.268 ; 
  LAYER V3 SPACING 0.072 ; 
      RECT 0.02 4.88 66.116 5.4 ; 
      RECT 65.648 1.026 66.116 5.4 ; 
      RECT 37.208 4.496 65.576 5.4 ; 
      RECT 31.88 4.496 37.136 5.4 ; 
      RECT 29 1.026 31.52 5.4 ; 
      RECT 0.56 4.496 28.928 5.4 ; 
      RECT 0.02 1.026 0.488 5.4 ; 
      RECT 65.504 1.026 66.116 4.688 ; 
      RECT 37.424 1.026 65.432 5.4 ; 
      RECT 34.436 1.026 37.352 4.688 ; 
      RECT 33.788 1.808 34.292 5.4 ; 
      RECT 28.784 1.424 33.68 4.688 ; 
      RECT 0.704 1.026 28.712 5.4 ; 
      RECT 0.02 1.026 0.632 4.688 ; 
      RECT 34.22 1.026 66.116 4.304 ; 
      RECT 0.02 1.424 34.148 4.304 ; 
      RECT 33.32 1.026 66.116 1.712 ; 
      RECT 0.02 1.026 33.248 4.304 ; 
      RECT 0.02 1.026 66.116 1.328 ; 
      RECT 0.02 9.2 66.116 9.72 ; 
      RECT 65.648 5.346 66.116 9.72 ; 
      RECT 37.208 8.816 65.576 9.72 ; 
      RECT 31.88 8.816 37.136 9.72 ; 
      RECT 29 5.346 31.52 9.72 ; 
      RECT 0.56 8.816 28.928 9.72 ; 
      RECT 0.02 5.346 0.488 9.72 ; 
      RECT 65.504 5.346 66.116 9.008 ; 
      RECT 37.424 5.346 65.432 9.72 ; 
      RECT 34.436 5.346 37.352 9.008 ; 
      RECT 33.788 6.128 34.292 9.72 ; 
      RECT 28.784 5.744 33.68 9.008 ; 
      RECT 0.704 5.346 28.712 9.72 ; 
      RECT 0.02 5.346 0.632 9.008 ; 
      RECT 34.22 5.346 66.116 8.624 ; 
      RECT 0.02 5.744 34.148 8.624 ; 
      RECT 33.32 5.346 66.116 6.032 ; 
      RECT 0.02 5.346 33.248 8.624 ; 
      RECT 0.02 5.346 66.116 5.648 ; 
      RECT 0.02 13.52 66.116 14.04 ; 
      RECT 65.648 9.666 66.116 14.04 ; 
      RECT 37.208 13.136 65.576 14.04 ; 
      RECT 31.88 13.136 37.136 14.04 ; 
      RECT 29 9.666 31.52 14.04 ; 
      RECT 0.56 13.136 28.928 14.04 ; 
      RECT 0.02 9.666 0.488 14.04 ; 
      RECT 65.504 9.666 66.116 13.328 ; 
      RECT 37.424 9.666 65.432 14.04 ; 
      RECT 34.436 9.666 37.352 13.328 ; 
      RECT 33.788 10.448 34.292 14.04 ; 
      RECT 28.784 10.064 33.68 13.328 ; 
      RECT 0.704 9.666 28.712 14.04 ; 
      RECT 0.02 9.666 0.632 13.328 ; 
      RECT 34.22 9.666 66.116 12.944 ; 
      RECT 0.02 10.064 34.148 12.944 ; 
      RECT 33.32 9.666 66.116 10.352 ; 
      RECT 0.02 9.666 33.248 12.944 ; 
      RECT 0.02 9.666 66.116 9.968 ; 
      RECT 0.02 17.84 66.116 18.36 ; 
      RECT 65.648 13.986 66.116 18.36 ; 
      RECT 37.208 17.456 65.576 18.36 ; 
      RECT 31.88 17.456 37.136 18.36 ; 
      RECT 29 13.986 31.52 18.36 ; 
      RECT 0.56 17.456 28.928 18.36 ; 
      RECT 0.02 13.986 0.488 18.36 ; 
      RECT 65.504 13.986 66.116 17.648 ; 
      RECT 37.424 13.986 65.432 18.36 ; 
      RECT 34.436 13.986 37.352 17.648 ; 
      RECT 33.788 14.768 34.292 18.36 ; 
      RECT 28.784 14.384 33.68 17.648 ; 
      RECT 0.704 13.986 28.712 18.36 ; 
      RECT 0.02 13.986 0.632 17.648 ; 
      RECT 34.22 13.986 66.116 17.264 ; 
      RECT 0.02 14.384 34.148 17.264 ; 
      RECT 33.32 13.986 66.116 14.672 ; 
      RECT 0.02 13.986 33.248 17.264 ; 
      RECT 0.02 13.986 66.116 14.288 ; 
      RECT 0.02 22.16 66.116 22.68 ; 
      RECT 65.648 18.306 66.116 22.68 ; 
      RECT 37.208 21.776 65.576 22.68 ; 
      RECT 31.88 21.776 37.136 22.68 ; 
      RECT 29 18.306 31.52 22.68 ; 
      RECT 0.56 21.776 28.928 22.68 ; 
      RECT 0.02 18.306 0.488 22.68 ; 
      RECT 65.504 18.306 66.116 21.968 ; 
      RECT 37.424 18.306 65.432 22.68 ; 
      RECT 34.436 18.306 37.352 21.968 ; 
      RECT 33.788 19.088 34.292 22.68 ; 
      RECT 28.784 18.704 33.68 21.968 ; 
      RECT 0.704 18.306 28.712 22.68 ; 
      RECT 0.02 18.306 0.632 21.968 ; 
      RECT 34.22 18.306 66.116 21.584 ; 
      RECT 0.02 18.704 34.148 21.584 ; 
      RECT 33.32 18.306 66.116 18.992 ; 
      RECT 0.02 18.306 33.248 21.584 ; 
      RECT 0.02 18.306 66.116 18.608 ; 
      RECT 0.02 26.48 66.116 27 ; 
      RECT 65.648 22.626 66.116 27 ; 
      RECT 37.208 26.096 65.576 27 ; 
      RECT 31.88 26.096 37.136 27 ; 
      RECT 29 22.626 31.52 27 ; 
      RECT 0.56 26.096 28.928 27 ; 
      RECT 0.02 22.626 0.488 27 ; 
      RECT 65.504 22.626 66.116 26.288 ; 
      RECT 37.424 22.626 65.432 27 ; 
      RECT 34.436 22.626 37.352 26.288 ; 
      RECT 33.788 23.408 34.292 27 ; 
      RECT 28.784 23.024 33.68 26.288 ; 
      RECT 0.704 22.626 28.712 27 ; 
      RECT 0.02 22.626 0.632 26.288 ; 
      RECT 34.22 22.626 66.116 25.904 ; 
      RECT 0.02 23.024 34.148 25.904 ; 
      RECT 33.32 22.626 66.116 23.312 ; 
      RECT 0.02 22.626 33.248 25.904 ; 
      RECT 0.02 22.626 66.116 22.928 ; 
      RECT 0.02 30.8 66.116 31.32 ; 
      RECT 65.648 26.946 66.116 31.32 ; 
      RECT 37.208 30.416 65.576 31.32 ; 
      RECT 31.88 30.416 37.136 31.32 ; 
      RECT 29 26.946 31.52 31.32 ; 
      RECT 0.56 30.416 28.928 31.32 ; 
      RECT 0.02 26.946 0.488 31.32 ; 
      RECT 65.504 26.946 66.116 30.608 ; 
      RECT 37.424 26.946 65.432 31.32 ; 
      RECT 34.436 26.946 37.352 30.608 ; 
      RECT 33.788 27.728 34.292 31.32 ; 
      RECT 28.784 27.344 33.68 30.608 ; 
      RECT 0.704 26.946 28.712 31.32 ; 
      RECT 0.02 26.946 0.632 30.608 ; 
      RECT 34.22 26.946 66.116 30.224 ; 
      RECT 0.02 27.344 34.148 30.224 ; 
      RECT 33.32 26.946 66.116 27.632 ; 
      RECT 0.02 26.946 33.248 30.224 ; 
      RECT 0.02 26.946 66.116 27.248 ; 
      RECT 0.02 35.12 66.116 35.64 ; 
      RECT 65.648 31.266 66.116 35.64 ; 
      RECT 37.208 34.736 65.576 35.64 ; 
      RECT 31.88 34.736 37.136 35.64 ; 
      RECT 29 31.266 31.52 35.64 ; 
      RECT 0.56 34.736 28.928 35.64 ; 
      RECT 0.02 31.266 0.488 35.64 ; 
      RECT 65.504 31.266 66.116 34.928 ; 
      RECT 37.424 31.266 65.432 35.64 ; 
      RECT 34.436 31.266 37.352 34.928 ; 
      RECT 33.788 32.048 34.292 35.64 ; 
      RECT 28.784 31.664 33.68 34.928 ; 
      RECT 0.704 31.266 28.712 35.64 ; 
      RECT 0.02 31.266 0.632 34.928 ; 
      RECT 34.22 31.266 66.116 34.544 ; 
      RECT 0.02 31.664 34.148 34.544 ; 
      RECT 33.32 31.266 66.116 31.952 ; 
      RECT 0.02 31.266 33.248 34.544 ; 
      RECT 0.02 31.266 66.116 31.568 ; 
      RECT 0.02 39.44 66.116 39.96 ; 
      RECT 65.648 35.586 66.116 39.96 ; 
      RECT 37.208 39.056 65.576 39.96 ; 
      RECT 31.88 39.056 37.136 39.96 ; 
      RECT 29 35.586 31.52 39.96 ; 
      RECT 0.56 39.056 28.928 39.96 ; 
      RECT 0.02 35.586 0.488 39.96 ; 
      RECT 65.504 35.586 66.116 39.248 ; 
      RECT 37.424 35.586 65.432 39.96 ; 
      RECT 34.436 35.586 37.352 39.248 ; 
      RECT 33.788 36.368 34.292 39.96 ; 
      RECT 28.784 35.984 33.68 39.248 ; 
      RECT 0.704 35.586 28.712 39.96 ; 
      RECT 0.02 35.586 0.632 39.248 ; 
      RECT 34.22 35.586 66.116 38.864 ; 
      RECT 0.02 35.984 34.148 38.864 ; 
      RECT 33.32 35.586 66.116 36.272 ; 
      RECT 0.02 35.586 33.248 38.864 ; 
      RECT 0.02 35.586 66.116 35.888 ; 
      RECT 0.02 43.76 66.116 44.28 ; 
      RECT 65.648 39.906 66.116 44.28 ; 
      RECT 37.208 43.376 65.576 44.28 ; 
      RECT 31.88 43.376 37.136 44.28 ; 
      RECT 29 39.906 31.52 44.28 ; 
      RECT 0.56 43.376 28.928 44.28 ; 
      RECT 0.02 39.906 0.488 44.28 ; 
      RECT 65.504 39.906 66.116 43.568 ; 
      RECT 37.424 39.906 65.432 44.28 ; 
      RECT 34.436 39.906 37.352 43.568 ; 
      RECT 33.788 40.688 34.292 44.28 ; 
      RECT 28.784 40.304 33.68 43.568 ; 
      RECT 0.704 39.906 28.712 44.28 ; 
      RECT 0.02 39.906 0.632 43.568 ; 
      RECT 34.22 39.906 66.116 43.184 ; 
      RECT 0.02 40.304 34.148 43.184 ; 
      RECT 33.32 39.906 66.116 40.592 ; 
      RECT 0.02 39.906 33.248 43.184 ; 
      RECT 0.02 39.906 66.116 40.208 ; 
      RECT 0.02 48.08 66.116 48.6 ; 
      RECT 65.648 44.226 66.116 48.6 ; 
      RECT 37.208 47.696 65.576 48.6 ; 
      RECT 31.88 47.696 37.136 48.6 ; 
      RECT 29 44.226 31.52 48.6 ; 
      RECT 0.56 47.696 28.928 48.6 ; 
      RECT 0.02 44.226 0.488 48.6 ; 
      RECT 65.504 44.226 66.116 47.888 ; 
      RECT 37.424 44.226 65.432 48.6 ; 
      RECT 34.436 44.226 37.352 47.888 ; 
      RECT 33.788 45.008 34.292 48.6 ; 
      RECT 28.784 44.624 33.68 47.888 ; 
      RECT 0.704 44.226 28.712 48.6 ; 
      RECT 0.02 44.226 0.632 47.888 ; 
      RECT 34.22 44.226 66.116 47.504 ; 
      RECT 0.02 44.624 34.148 47.504 ; 
      RECT 33.32 44.226 66.116 44.912 ; 
      RECT 0.02 44.226 33.248 47.504 ; 
      RECT 0.02 44.226 66.116 44.528 ; 
      RECT 0.02 52.4 66.116 52.92 ; 
      RECT 65.648 48.546 66.116 52.92 ; 
      RECT 37.208 52.016 65.576 52.92 ; 
      RECT 31.88 52.016 37.136 52.92 ; 
      RECT 29 48.546 31.52 52.92 ; 
      RECT 0.56 52.016 28.928 52.92 ; 
      RECT 0.02 48.546 0.488 52.92 ; 
      RECT 65.504 48.546 66.116 52.208 ; 
      RECT 37.424 48.546 65.432 52.92 ; 
      RECT 34.436 48.546 37.352 52.208 ; 
      RECT 33.788 49.328 34.292 52.92 ; 
      RECT 28.784 48.944 33.68 52.208 ; 
      RECT 0.704 48.546 28.712 52.92 ; 
      RECT 0.02 48.546 0.632 52.208 ; 
      RECT 34.22 48.546 66.116 51.824 ; 
      RECT 0.02 48.944 34.148 51.824 ; 
      RECT 33.32 48.546 66.116 49.232 ; 
      RECT 0.02 48.546 33.248 51.824 ; 
      RECT 0.02 48.546 66.116 48.848 ; 
      RECT 0.02 56.72 66.116 57.24 ; 
      RECT 65.648 52.866 66.116 57.24 ; 
      RECT 37.208 56.336 65.576 57.24 ; 
      RECT 31.88 56.336 37.136 57.24 ; 
      RECT 29 52.866 31.52 57.24 ; 
      RECT 0.56 56.336 28.928 57.24 ; 
      RECT 0.02 52.866 0.488 57.24 ; 
      RECT 65.504 52.866 66.116 56.528 ; 
      RECT 37.424 52.866 65.432 57.24 ; 
      RECT 34.436 52.866 37.352 56.528 ; 
      RECT 33.788 53.648 34.292 57.24 ; 
      RECT 28.784 53.264 33.68 56.528 ; 
      RECT 0.704 52.866 28.712 57.24 ; 
      RECT 0.02 52.866 0.632 56.528 ; 
      RECT 34.22 52.866 66.116 56.144 ; 
      RECT 0.02 53.264 34.148 56.144 ; 
      RECT 33.32 52.866 66.116 53.552 ; 
      RECT 0.02 52.866 33.248 56.144 ; 
      RECT 0.02 52.866 66.116 53.168 ; 
      RECT 0.02 61.04 66.116 61.56 ; 
      RECT 65.648 57.186 66.116 61.56 ; 
      RECT 37.208 60.656 65.576 61.56 ; 
      RECT 31.88 60.656 37.136 61.56 ; 
      RECT 29 57.186 31.52 61.56 ; 
      RECT 0.56 60.656 28.928 61.56 ; 
      RECT 0.02 57.186 0.488 61.56 ; 
      RECT 65.504 57.186 66.116 60.848 ; 
      RECT 37.424 57.186 65.432 61.56 ; 
      RECT 34.436 57.186 37.352 60.848 ; 
      RECT 33.788 57.968 34.292 61.56 ; 
      RECT 28.784 57.584 33.68 60.848 ; 
      RECT 0.704 57.186 28.712 61.56 ; 
      RECT 0.02 57.186 0.632 60.848 ; 
      RECT 34.22 57.186 66.116 60.464 ; 
      RECT 0.02 57.584 34.148 60.464 ; 
      RECT 33.32 57.186 66.116 57.872 ; 
      RECT 0.02 57.186 33.248 60.464 ; 
      RECT 0.02 57.186 66.116 57.488 ; 
      RECT 0.02 65.36 66.116 65.88 ; 
      RECT 65.648 61.506 66.116 65.88 ; 
      RECT 37.208 64.976 65.576 65.88 ; 
      RECT 31.88 64.976 37.136 65.88 ; 
      RECT 29 61.506 31.52 65.88 ; 
      RECT 0.56 64.976 28.928 65.88 ; 
      RECT 0.02 61.506 0.488 65.88 ; 
      RECT 65.504 61.506 66.116 65.168 ; 
      RECT 37.424 61.506 65.432 65.88 ; 
      RECT 34.436 61.506 37.352 65.168 ; 
      RECT 33.788 62.288 34.292 65.88 ; 
      RECT 28.784 61.904 33.68 65.168 ; 
      RECT 0.704 61.506 28.712 65.88 ; 
      RECT 0.02 61.506 0.632 65.168 ; 
      RECT 34.22 61.506 66.116 64.784 ; 
      RECT 0.02 61.904 34.148 64.784 ; 
      RECT 33.32 61.506 66.116 62.192 ; 
      RECT 0.02 61.506 33.248 64.784 ; 
      RECT 0.02 61.506 66.116 61.808 ; 
      RECT 0.02 69.68 66.116 70.2 ; 
      RECT 65.648 65.826 66.116 70.2 ; 
      RECT 37.208 69.296 65.576 70.2 ; 
      RECT 31.88 69.296 37.136 70.2 ; 
      RECT 29 65.826 31.52 70.2 ; 
      RECT 0.56 69.296 28.928 70.2 ; 
      RECT 0.02 65.826 0.488 70.2 ; 
      RECT 65.504 65.826 66.116 69.488 ; 
      RECT 37.424 65.826 65.432 70.2 ; 
      RECT 34.436 65.826 37.352 69.488 ; 
      RECT 33.788 66.608 34.292 70.2 ; 
      RECT 28.784 66.224 33.68 69.488 ; 
      RECT 0.704 65.826 28.712 70.2 ; 
      RECT 0.02 65.826 0.632 69.488 ; 
      RECT 34.22 65.826 66.116 69.104 ; 
      RECT 0.02 66.224 34.148 69.104 ; 
      RECT 33.32 65.826 66.116 66.512 ; 
      RECT 0.02 65.826 33.248 69.104 ; 
      RECT 0.02 65.826 66.116 66.128 ; 
      RECT 0.02 74 66.116 74.52 ; 
      RECT 65.648 70.146 66.116 74.52 ; 
      RECT 37.208 73.616 65.576 74.52 ; 
      RECT 31.88 73.616 37.136 74.52 ; 
      RECT 29 70.146 31.52 74.52 ; 
      RECT 0.56 73.616 28.928 74.52 ; 
      RECT 0.02 70.146 0.488 74.52 ; 
      RECT 65.504 70.146 66.116 73.808 ; 
      RECT 37.424 70.146 65.432 74.52 ; 
      RECT 34.436 70.146 37.352 73.808 ; 
      RECT 33.788 70.928 34.292 74.52 ; 
      RECT 28.784 70.544 33.68 73.808 ; 
      RECT 0.704 70.146 28.712 74.52 ; 
      RECT 0.02 70.146 0.632 73.808 ; 
      RECT 34.22 70.146 66.116 73.424 ; 
      RECT 0.02 70.544 34.148 73.424 ; 
      RECT 33.32 70.146 66.116 70.832 ; 
      RECT 0.02 70.146 33.248 73.424 ; 
      RECT 0.02 70.146 66.116 70.448 ; 
      RECT 0.02 78.32 66.116 78.84 ; 
      RECT 65.648 74.466 66.116 78.84 ; 
      RECT 37.208 77.936 65.576 78.84 ; 
      RECT 31.88 77.936 37.136 78.84 ; 
      RECT 29 74.466 31.52 78.84 ; 
      RECT 0.56 77.936 28.928 78.84 ; 
      RECT 0.02 74.466 0.488 78.84 ; 
      RECT 65.504 74.466 66.116 78.128 ; 
      RECT 37.424 74.466 65.432 78.84 ; 
      RECT 34.436 74.466 37.352 78.128 ; 
      RECT 33.788 75.248 34.292 78.84 ; 
      RECT 28.784 74.864 33.68 78.128 ; 
      RECT 0.704 74.466 28.712 78.84 ; 
      RECT 0.02 74.466 0.632 78.128 ; 
      RECT 34.22 74.466 66.116 77.744 ; 
      RECT 0.02 74.864 34.148 77.744 ; 
      RECT 33.32 74.466 66.116 75.152 ; 
      RECT 0.02 74.466 33.248 77.744 ; 
      RECT 0.02 74.466 66.116 74.768 ; 
      RECT 0.02 82.64 66.116 83.16 ; 
      RECT 65.648 78.786 66.116 83.16 ; 
      RECT 37.208 82.256 65.576 83.16 ; 
      RECT 31.88 82.256 37.136 83.16 ; 
      RECT 29 78.786 31.52 83.16 ; 
      RECT 0.56 82.256 28.928 83.16 ; 
      RECT 0.02 78.786 0.488 83.16 ; 
      RECT 65.504 78.786 66.116 82.448 ; 
      RECT 37.424 78.786 65.432 83.16 ; 
      RECT 34.436 78.786 37.352 82.448 ; 
      RECT 33.788 79.568 34.292 83.16 ; 
      RECT 28.784 79.184 33.68 82.448 ; 
      RECT 0.704 78.786 28.712 83.16 ; 
      RECT 0.02 78.786 0.632 82.448 ; 
      RECT 34.22 78.786 66.116 82.064 ; 
      RECT 0.02 79.184 34.148 82.064 ; 
      RECT 33.32 78.786 66.116 79.472 ; 
      RECT 0.02 78.786 33.248 82.064 ; 
      RECT 0.02 78.786 66.116 79.088 ; 
      RECT 0.02 86.96 66.116 87.48 ; 
      RECT 65.648 83.106 66.116 87.48 ; 
      RECT 37.208 86.576 65.576 87.48 ; 
      RECT 31.88 86.576 37.136 87.48 ; 
      RECT 29 83.106 31.52 87.48 ; 
      RECT 0.56 86.576 28.928 87.48 ; 
      RECT 0.02 83.106 0.488 87.48 ; 
      RECT 65.504 83.106 66.116 86.768 ; 
      RECT 37.424 83.106 65.432 87.48 ; 
      RECT 34.436 83.106 37.352 86.768 ; 
      RECT 33.788 83.888 34.292 87.48 ; 
      RECT 28.784 83.504 33.68 86.768 ; 
      RECT 0.704 83.106 28.712 87.48 ; 
      RECT 0.02 83.106 0.632 86.768 ; 
      RECT 34.22 83.106 66.116 86.384 ; 
      RECT 0.02 83.504 34.148 86.384 ; 
      RECT 33.32 83.106 66.116 83.792 ; 
      RECT 0.02 83.106 33.248 86.384 ; 
      RECT 0.02 83.106 66.116 83.408 ; 
      RECT 0.02 91.28 66.116 91.8 ; 
      RECT 65.648 87.426 66.116 91.8 ; 
      RECT 37.208 90.896 65.576 91.8 ; 
      RECT 31.88 90.896 37.136 91.8 ; 
      RECT 29 87.426 31.52 91.8 ; 
      RECT 0.56 90.896 28.928 91.8 ; 
      RECT 0.02 87.426 0.488 91.8 ; 
      RECT 65.504 87.426 66.116 91.088 ; 
      RECT 37.424 87.426 65.432 91.8 ; 
      RECT 34.436 87.426 37.352 91.088 ; 
      RECT 33.788 88.208 34.292 91.8 ; 
      RECT 28.784 87.824 33.68 91.088 ; 
      RECT 0.704 87.426 28.712 91.8 ; 
      RECT 0.02 87.426 0.632 91.088 ; 
      RECT 34.22 87.426 66.116 90.704 ; 
      RECT 0.02 87.824 34.148 90.704 ; 
      RECT 33.32 87.426 66.116 88.112 ; 
      RECT 0.02 87.426 33.248 90.704 ; 
      RECT 0.02 87.426 66.116 87.728 ; 
      RECT 0.02 95.6 66.116 96.12 ; 
      RECT 65.648 91.746 66.116 96.12 ; 
      RECT 37.208 95.216 65.576 96.12 ; 
      RECT 31.88 95.216 37.136 96.12 ; 
      RECT 29 91.746 31.52 96.12 ; 
      RECT 0.56 95.216 28.928 96.12 ; 
      RECT 0.02 91.746 0.488 96.12 ; 
      RECT 65.504 91.746 66.116 95.408 ; 
      RECT 37.424 91.746 65.432 96.12 ; 
      RECT 34.436 91.746 37.352 95.408 ; 
      RECT 33.788 92.528 34.292 96.12 ; 
      RECT 28.784 92.144 33.68 95.408 ; 
      RECT 0.704 91.746 28.712 96.12 ; 
      RECT 0.02 91.746 0.632 95.408 ; 
      RECT 34.22 91.746 66.116 95.024 ; 
      RECT 0.02 92.144 34.148 95.024 ; 
      RECT 33.32 91.746 66.116 92.432 ; 
      RECT 0.02 91.746 33.248 95.024 ; 
      RECT 0.02 91.746 66.116 92.048 ; 
      RECT 0.02 99.92 66.116 100.44 ; 
      RECT 65.648 96.066 66.116 100.44 ; 
      RECT 37.208 99.536 65.576 100.44 ; 
      RECT 31.88 99.536 37.136 100.44 ; 
      RECT 29 96.066 31.52 100.44 ; 
      RECT 0.56 99.536 28.928 100.44 ; 
      RECT 0.02 96.066 0.488 100.44 ; 
      RECT 65.504 96.066 66.116 99.728 ; 
      RECT 37.424 96.066 65.432 100.44 ; 
      RECT 34.436 96.066 37.352 99.728 ; 
      RECT 33.788 96.848 34.292 100.44 ; 
      RECT 28.784 96.464 33.68 99.728 ; 
      RECT 0.704 96.066 28.712 100.44 ; 
      RECT 0.02 96.066 0.632 99.728 ; 
      RECT 34.22 96.066 66.116 99.344 ; 
      RECT 0.02 96.464 34.148 99.344 ; 
      RECT 33.32 96.066 66.116 96.752 ; 
      RECT 0.02 96.066 33.248 99.344 ; 
      RECT 0.02 96.066 66.116 96.368 ; 
      RECT 0.02 104.24 66.116 104.76 ; 
      RECT 65.648 100.386 66.116 104.76 ; 
      RECT 37.208 103.856 65.576 104.76 ; 
      RECT 31.88 103.856 37.136 104.76 ; 
      RECT 29 100.386 31.52 104.76 ; 
      RECT 0.56 103.856 28.928 104.76 ; 
      RECT 0.02 100.386 0.488 104.76 ; 
      RECT 65.504 100.386 66.116 104.048 ; 
      RECT 37.424 100.386 65.432 104.76 ; 
      RECT 34.436 100.386 37.352 104.048 ; 
      RECT 33.788 101.168 34.292 104.76 ; 
      RECT 28.784 100.784 33.68 104.048 ; 
      RECT 0.704 100.386 28.712 104.76 ; 
      RECT 0.02 100.386 0.632 104.048 ; 
      RECT 34.22 100.386 66.116 103.664 ; 
      RECT 0.02 100.784 34.148 103.664 ; 
      RECT 33.32 100.386 66.116 101.072 ; 
      RECT 0.02 100.386 33.248 103.664 ; 
      RECT 0.02 100.386 66.116 100.688 ; 
      RECT 0.02 108.56 66.116 109.08 ; 
      RECT 65.648 104.706 66.116 109.08 ; 
      RECT 37.208 108.176 65.576 109.08 ; 
      RECT 31.88 108.176 37.136 109.08 ; 
      RECT 29 104.706 31.52 109.08 ; 
      RECT 0.56 108.176 28.928 109.08 ; 
      RECT 0.02 104.706 0.488 109.08 ; 
      RECT 65.504 104.706 66.116 108.368 ; 
      RECT 37.424 104.706 65.432 109.08 ; 
      RECT 34.436 104.706 37.352 108.368 ; 
      RECT 33.788 105.488 34.292 109.08 ; 
      RECT 28.784 105.104 33.68 108.368 ; 
      RECT 0.704 104.706 28.712 109.08 ; 
      RECT 0.02 104.706 0.632 108.368 ; 
      RECT 34.22 104.706 66.116 107.984 ; 
      RECT 0.02 105.104 34.148 107.984 ; 
      RECT 33.32 104.706 66.116 105.392 ; 
      RECT 0.02 104.706 33.248 107.984 ; 
      RECT 0.02 104.706 66.116 105.008 ; 
      RECT 0.02 112.88 66.116 113.4 ; 
      RECT 65.648 109.026 66.116 113.4 ; 
      RECT 37.208 112.496 65.576 113.4 ; 
      RECT 31.88 112.496 37.136 113.4 ; 
      RECT 29 109.026 31.52 113.4 ; 
      RECT 0.56 112.496 28.928 113.4 ; 
      RECT 0.02 109.026 0.488 113.4 ; 
      RECT 65.504 109.026 66.116 112.688 ; 
      RECT 37.424 109.026 65.432 113.4 ; 
      RECT 34.436 109.026 37.352 112.688 ; 
      RECT 33.788 109.808 34.292 113.4 ; 
      RECT 28.784 109.424 33.68 112.688 ; 
      RECT 0.704 109.026 28.712 113.4 ; 
      RECT 0.02 109.026 0.632 112.688 ; 
      RECT 34.22 109.026 66.116 112.304 ; 
      RECT 0.02 109.424 34.148 112.304 ; 
      RECT 33.32 109.026 66.116 109.712 ; 
      RECT 0.02 109.026 33.248 112.304 ; 
      RECT 0.02 109.026 66.116 109.328 ; 
      RECT 0.02 117.2 66.116 117.72 ; 
      RECT 65.648 113.346 66.116 117.72 ; 
      RECT 37.208 116.816 65.576 117.72 ; 
      RECT 31.88 116.816 37.136 117.72 ; 
      RECT 29 113.346 31.52 117.72 ; 
      RECT 0.56 116.816 28.928 117.72 ; 
      RECT 0.02 113.346 0.488 117.72 ; 
      RECT 65.504 113.346 66.116 117.008 ; 
      RECT 37.424 113.346 65.432 117.72 ; 
      RECT 34.436 113.346 37.352 117.008 ; 
      RECT 33.788 114.128 34.292 117.72 ; 
      RECT 28.784 113.744 33.68 117.008 ; 
      RECT 0.704 113.346 28.712 117.72 ; 
      RECT 0.02 113.346 0.632 117.008 ; 
      RECT 34.22 113.346 66.116 116.624 ; 
      RECT 0.02 113.744 34.148 116.624 ; 
      RECT 33.32 113.346 66.116 114.032 ; 
      RECT 0.02 113.346 33.248 116.624 ; 
      RECT 0.02 113.346 66.116 113.648 ; 
      RECT 0.02 121.52 66.116 122.04 ; 
      RECT 65.648 117.666 66.116 122.04 ; 
      RECT 37.208 121.136 65.576 122.04 ; 
      RECT 31.88 121.136 37.136 122.04 ; 
      RECT 29 117.666 31.52 122.04 ; 
      RECT 0.56 121.136 28.928 122.04 ; 
      RECT 0.02 117.666 0.488 122.04 ; 
      RECT 65.504 117.666 66.116 121.328 ; 
      RECT 37.424 117.666 65.432 122.04 ; 
      RECT 34.436 117.666 37.352 121.328 ; 
      RECT 33.788 118.448 34.292 122.04 ; 
      RECT 28.784 118.064 33.68 121.328 ; 
      RECT 0.704 117.666 28.712 122.04 ; 
      RECT 0.02 117.666 0.632 121.328 ; 
      RECT 34.22 117.666 66.116 120.944 ; 
      RECT 0.02 118.064 34.148 120.944 ; 
      RECT 33.32 117.666 66.116 118.352 ; 
      RECT 0.02 117.666 33.248 120.944 ; 
      RECT 0.02 117.666 66.116 117.968 ; 
      RECT 0.02 125.84 66.116 126.36 ; 
      RECT 65.648 121.986 66.116 126.36 ; 
      RECT 37.208 125.456 65.576 126.36 ; 
      RECT 31.88 125.456 37.136 126.36 ; 
      RECT 29 121.986 31.52 126.36 ; 
      RECT 0.56 125.456 28.928 126.36 ; 
      RECT 0.02 121.986 0.488 126.36 ; 
      RECT 65.504 121.986 66.116 125.648 ; 
      RECT 37.424 121.986 65.432 126.36 ; 
      RECT 34.436 121.986 37.352 125.648 ; 
      RECT 33.788 122.768 34.292 126.36 ; 
      RECT 28.784 122.384 33.68 125.648 ; 
      RECT 0.704 121.986 28.712 126.36 ; 
      RECT 0.02 121.986 0.632 125.648 ; 
      RECT 34.22 121.986 66.116 125.264 ; 
      RECT 0.02 122.384 34.148 125.264 ; 
      RECT 33.32 121.986 66.116 122.672 ; 
      RECT 0.02 121.986 33.248 125.264 ; 
      RECT 0.02 121.986 66.116 122.288 ; 
      RECT 0.02 130.16 66.116 130.68 ; 
      RECT 65.648 126.306 66.116 130.68 ; 
      RECT 37.208 129.776 65.576 130.68 ; 
      RECT 31.88 129.776 37.136 130.68 ; 
      RECT 29 126.306 31.52 130.68 ; 
      RECT 0.56 129.776 28.928 130.68 ; 
      RECT 0.02 126.306 0.488 130.68 ; 
      RECT 65.504 126.306 66.116 129.968 ; 
      RECT 37.424 126.306 65.432 130.68 ; 
      RECT 34.436 126.306 37.352 129.968 ; 
      RECT 33.788 127.088 34.292 130.68 ; 
      RECT 28.784 126.704 33.68 129.968 ; 
      RECT 0.704 126.306 28.712 130.68 ; 
      RECT 0.02 126.306 0.632 129.968 ; 
      RECT 34.22 126.306 66.116 129.584 ; 
      RECT 0.02 126.704 34.148 129.584 ; 
      RECT 33.32 126.306 66.116 126.992 ; 
      RECT 0.02 126.306 33.248 129.584 ; 
      RECT 0.02 126.306 66.116 126.608 ; 
      RECT 0.02 134.48 66.116 135 ; 
      RECT 65.648 130.626 66.116 135 ; 
      RECT 37.208 134.096 65.576 135 ; 
      RECT 31.88 134.096 37.136 135 ; 
      RECT 29 130.626 31.52 135 ; 
      RECT 0.56 134.096 28.928 135 ; 
      RECT 0.02 130.626 0.488 135 ; 
      RECT 65.504 130.626 66.116 134.288 ; 
      RECT 37.424 130.626 65.432 135 ; 
      RECT 34.436 130.626 37.352 134.288 ; 
      RECT 33.788 131.408 34.292 135 ; 
      RECT 28.784 131.024 33.68 134.288 ; 
      RECT 0.704 130.626 28.712 135 ; 
      RECT 0.02 130.626 0.632 134.288 ; 
      RECT 34.22 130.626 66.116 133.904 ; 
      RECT 0.02 131.024 34.148 133.904 ; 
      RECT 33.32 130.626 66.116 131.312 ; 
      RECT 0.02 130.626 33.248 133.904 ; 
      RECT 0.02 130.626 66.116 130.928 ; 
      RECT 0.02 138.8 66.116 139.32 ; 
      RECT 65.648 134.946 66.116 139.32 ; 
      RECT 37.208 138.416 65.576 139.32 ; 
      RECT 31.88 138.416 37.136 139.32 ; 
      RECT 29 134.946 31.52 139.32 ; 
      RECT 0.56 138.416 28.928 139.32 ; 
      RECT 0.02 134.946 0.488 139.32 ; 
      RECT 65.504 134.946 66.116 138.608 ; 
      RECT 37.424 134.946 65.432 139.32 ; 
      RECT 34.436 134.946 37.352 138.608 ; 
      RECT 33.788 135.728 34.292 139.32 ; 
      RECT 28.784 135.344 33.68 138.608 ; 
      RECT 0.704 134.946 28.712 139.32 ; 
      RECT 0.02 134.946 0.632 138.608 ; 
      RECT 34.22 134.946 66.116 138.224 ; 
      RECT 0.02 135.344 34.148 138.224 ; 
      RECT 33.32 134.946 66.116 135.632 ; 
      RECT 0.02 134.946 33.248 138.224 ; 
      RECT 0.02 134.946 66.116 135.248 ; 
      RECT 0.02 143.12 66.116 143.64 ; 
      RECT 65.648 139.266 66.116 143.64 ; 
      RECT 37.208 142.736 65.576 143.64 ; 
      RECT 31.88 142.736 37.136 143.64 ; 
      RECT 29 139.266 31.52 143.64 ; 
      RECT 0.56 142.736 28.928 143.64 ; 
      RECT 0.02 139.266 0.488 143.64 ; 
      RECT 65.504 139.266 66.116 142.928 ; 
      RECT 37.424 139.266 65.432 143.64 ; 
      RECT 34.436 139.266 37.352 142.928 ; 
      RECT 33.788 140.048 34.292 143.64 ; 
      RECT 28.784 139.664 33.68 142.928 ; 
      RECT 0.704 139.266 28.712 143.64 ; 
      RECT 0.02 139.266 0.632 142.928 ; 
      RECT 34.22 139.266 66.116 142.544 ; 
      RECT 0.02 139.664 34.148 142.544 ; 
      RECT 33.32 139.266 66.116 139.952 ; 
      RECT 0.02 139.266 33.248 142.544 ; 
      RECT 0.02 139.266 66.116 139.568 ; 
      RECT 0.02 147.44 66.116 147.96 ; 
      RECT 65.648 143.586 66.116 147.96 ; 
      RECT 37.208 147.056 65.576 147.96 ; 
      RECT 31.88 147.056 37.136 147.96 ; 
      RECT 29 143.586 31.52 147.96 ; 
      RECT 0.56 147.056 28.928 147.96 ; 
      RECT 0.02 143.586 0.488 147.96 ; 
      RECT 65.504 143.586 66.116 147.248 ; 
      RECT 37.424 143.586 65.432 147.96 ; 
      RECT 34.436 143.586 37.352 147.248 ; 
      RECT 33.788 144.368 34.292 147.96 ; 
      RECT 28.784 143.984 33.68 147.248 ; 
      RECT 0.704 143.586 28.712 147.96 ; 
      RECT 0.02 143.586 0.632 147.248 ; 
      RECT 34.22 143.586 66.116 146.864 ; 
      RECT 0.02 143.984 34.148 146.864 ; 
      RECT 33.32 143.586 66.116 144.272 ; 
      RECT 0.02 143.586 33.248 146.864 ; 
      RECT 0.02 143.586 66.116 143.888 ; 
      RECT 0.02 151.76 66.116 152.28 ; 
      RECT 65.648 147.906 66.116 152.28 ; 
      RECT 37.208 151.376 65.576 152.28 ; 
      RECT 31.88 151.376 37.136 152.28 ; 
      RECT 29 147.906 31.52 152.28 ; 
      RECT 0.56 151.376 28.928 152.28 ; 
      RECT 0.02 147.906 0.488 152.28 ; 
      RECT 65.504 147.906 66.116 151.568 ; 
      RECT 37.424 147.906 65.432 152.28 ; 
      RECT 34.436 147.906 37.352 151.568 ; 
      RECT 33.788 148.688 34.292 152.28 ; 
      RECT 28.784 148.304 33.68 151.568 ; 
      RECT 0.704 147.906 28.712 152.28 ; 
      RECT 0.02 147.906 0.632 151.568 ; 
      RECT 34.22 147.906 66.116 151.184 ; 
      RECT 0.02 148.304 34.148 151.184 ; 
      RECT 33.32 147.906 66.116 148.592 ; 
      RECT 0.02 147.906 33.248 151.184 ; 
      RECT 0.02 147.906 66.116 148.208 ; 
      RECT 0.02 156.08 66.116 156.6 ; 
      RECT 65.648 152.226 66.116 156.6 ; 
      RECT 37.208 155.696 65.576 156.6 ; 
      RECT 31.88 155.696 37.136 156.6 ; 
      RECT 29 152.226 31.52 156.6 ; 
      RECT 0.56 155.696 28.928 156.6 ; 
      RECT 0.02 152.226 0.488 156.6 ; 
      RECT 65.504 152.226 66.116 155.888 ; 
      RECT 37.424 152.226 65.432 156.6 ; 
      RECT 34.436 152.226 37.352 155.888 ; 
      RECT 33.788 153.008 34.292 156.6 ; 
      RECT 28.784 152.624 33.68 155.888 ; 
      RECT 0.704 152.226 28.712 156.6 ; 
      RECT 0.02 152.226 0.632 155.888 ; 
      RECT 34.22 152.226 66.116 155.504 ; 
      RECT 0.02 152.624 34.148 155.504 ; 
      RECT 33.32 152.226 66.116 152.912 ; 
      RECT 0.02 152.226 33.248 155.504 ; 
      RECT 0.02 152.226 66.116 152.528 ; 
      RECT 0.02 160.4 66.116 160.92 ; 
      RECT 65.648 156.546 66.116 160.92 ; 
      RECT 37.208 160.016 65.576 160.92 ; 
      RECT 31.88 160.016 37.136 160.92 ; 
      RECT 29 156.546 31.52 160.92 ; 
      RECT 0.56 160.016 28.928 160.92 ; 
      RECT 0.02 156.546 0.488 160.92 ; 
      RECT 65.504 156.546 66.116 160.208 ; 
      RECT 37.424 156.546 65.432 160.92 ; 
      RECT 34.436 156.546 37.352 160.208 ; 
      RECT 33.788 157.328 34.292 160.92 ; 
      RECT 28.784 156.944 33.68 160.208 ; 
      RECT 0.704 156.546 28.712 160.92 ; 
      RECT 0.02 156.546 0.632 160.208 ; 
      RECT 34.22 156.546 66.116 159.824 ; 
      RECT 0.02 156.944 34.148 159.824 ; 
      RECT 33.32 156.546 66.116 157.232 ; 
      RECT 0.02 156.546 33.248 159.824 ; 
      RECT 0.02 156.546 66.116 156.848 ; 
      RECT 0 190.068 66.096 195.402 ; 
      RECT 43.236 160.788 66.096 195.402 ; 
      RECT 34.436 176.244 66.096 195.402 ; 
      RECT 38.052 165.876 66.096 195.402 ; 
      RECT 34.228 160.788 34.364 195.402 ; 
      RECT 34.02 160.788 34.156 195.402 ; 
      RECT 33.812 160.788 33.948 195.402 ; 
      RECT 33.604 160.788 33.74 195.402 ; 
      RECT 0 188.34 33.532 195.402 ; 
      RECT 32.564 177.396 66.096 189.204 ; 
      RECT 32.356 160.788 32.492 195.402 ; 
      RECT 32.148 160.788 32.284 195.402 ; 
      RECT 31.94 160.788 32.076 195.402 ; 
      RECT 31.732 160.788 31.868 195.402 ; 
      RECT 0 167.028 31.66 195.402 ; 
      RECT 0 175.668 33.532 187.476 ; 
      RECT 32.564 164.724 37.116 176.532 ; 
      RECT 37.26 166.644 66.096 195.402 ; 
      RECT 0 175.668 37.188 176.532 ; 
      RECT 32.564 166.644 66.096 176.148 ; 
      RECT 29.844 162.996 32.94 174.804 ; 
      RECT 28.98 163.572 31.66 195.402 ; 
      RECT 0 165.876 28.908 195.402 ; 
      RECT 27.252 160.788 29.052 166.932 ; 
      RECT 0 166.26 37.98 166.932 ; 
      RECT 37.188 165.876 66.096 166.548 ; 
      RECT 42.372 160.788 43.164 195.402 ; 
      RECT 27.252 165.108 42.3 166.164 ; 
      RECT 23.796 163.572 27.18 195.402 ; 
      RECT 0 160.788 23.724 195.402 ; 
      RECT 41.508 160.788 66.096 165.78 ; 
      RECT 40.644 163.572 66.096 165.78 ; 
      RECT 0 164.726 40.572 165.78 ; 
      RECT 39.78 160.788 41.436 165.012 ; 
      RECT 37.404 163.572 66.096 165.012 ; 
      RECT 34.436 163.572 37.332 166.164 ; 
      RECT 32.564 163.38 33.532 195.402 ; 
      RECT 33.012 160.788 34.524 163.86 ; 
      RECT 34.596 163.38 39.708 163.862 ; 
      RECT 26.388 163.38 29.772 165.78 ; 
      RECT 24.66 163.38 26.316 195.402 ; 
      RECT 0 160.788 24.588 165.78 ; 
      RECT 38.916 160.788 66.096 163.476 ; 
      RECT 33.012 161.108 38.844 163.476 ; 
      RECT 29.124 162.996 32.94 163.476 ; 
      RECT 25.524 160.788 29.052 163.476 ; 
      RECT 0 160.788 25.452 163.476 ; 
      RECT 37.188 160.788 66.096 163.284 ; 
      RECT 32.564 161.108 66.096 163.284 ; 
      RECT 0 160.788 31.66 163.284 ; 
      RECT 0 160.788 37.116 162.132 ; 
      RECT 0 160.788 66.096 161.012 ; 
        RECT 0.02 197.228 66.116 197.748 ; 
        RECT 65.648 193.374 66.116 197.748 ; 
        RECT 37.208 196.844 65.576 197.748 ; 
        RECT 31.88 196.844 37.136 197.748 ; 
        RECT 29 193.374 31.52 197.748 ; 
        RECT 0.56 196.844 28.928 197.748 ; 
        RECT 0.02 193.374 0.488 197.748 ; 
        RECT 65.504 193.374 66.116 197.036 ; 
        RECT 37.424 193.374 65.432 197.748 ; 
        RECT 34.436 193.374 37.352 197.036 ; 
        RECT 33.788 194.156 34.292 197.748 ; 
        RECT 28.784 193.772 33.68 197.036 ; 
        RECT 0.704 193.374 28.712 197.748 ; 
        RECT 0.02 193.374 0.632 197.036 ; 
        RECT 34.22 193.374 66.116 196.652 ; 
        RECT 0.02 193.772 34.148 196.652 ; 
        RECT 33.32 193.374 66.116 194.06 ; 
        RECT 0.02 193.374 33.248 196.652 ; 
        RECT 0.02 193.374 66.116 193.676 ; 
        RECT 0.02 201.548 66.116 202.068 ; 
        RECT 65.648 197.694 66.116 202.068 ; 
        RECT 37.208 201.164 65.576 202.068 ; 
        RECT 31.88 201.164 37.136 202.068 ; 
        RECT 29 197.694 31.52 202.068 ; 
        RECT 0.56 201.164 28.928 202.068 ; 
        RECT 0.02 197.694 0.488 202.068 ; 
        RECT 65.504 197.694 66.116 201.356 ; 
        RECT 37.424 197.694 65.432 202.068 ; 
        RECT 34.436 197.694 37.352 201.356 ; 
        RECT 33.788 198.476 34.292 202.068 ; 
        RECT 28.784 198.092 33.68 201.356 ; 
        RECT 0.704 197.694 28.712 202.068 ; 
        RECT 0.02 197.694 0.632 201.356 ; 
        RECT 34.22 197.694 66.116 200.972 ; 
        RECT 0.02 198.092 34.148 200.972 ; 
        RECT 33.32 197.694 66.116 198.38 ; 
        RECT 0.02 197.694 33.248 200.972 ; 
        RECT 0.02 197.694 66.116 197.996 ; 
        RECT 0.02 205.868 66.116 206.388 ; 
        RECT 65.648 202.014 66.116 206.388 ; 
        RECT 37.208 205.484 65.576 206.388 ; 
        RECT 31.88 205.484 37.136 206.388 ; 
        RECT 29 202.014 31.52 206.388 ; 
        RECT 0.56 205.484 28.928 206.388 ; 
        RECT 0.02 202.014 0.488 206.388 ; 
        RECT 65.504 202.014 66.116 205.676 ; 
        RECT 37.424 202.014 65.432 206.388 ; 
        RECT 34.436 202.014 37.352 205.676 ; 
        RECT 33.788 202.796 34.292 206.388 ; 
        RECT 28.784 202.412 33.68 205.676 ; 
        RECT 0.704 202.014 28.712 206.388 ; 
        RECT 0.02 202.014 0.632 205.676 ; 
        RECT 34.22 202.014 66.116 205.292 ; 
        RECT 0.02 202.412 34.148 205.292 ; 
        RECT 33.32 202.014 66.116 202.7 ; 
        RECT 0.02 202.014 33.248 205.292 ; 
        RECT 0.02 202.014 66.116 202.316 ; 
        RECT 0.02 210.188 66.116 210.708 ; 
        RECT 65.648 206.334 66.116 210.708 ; 
        RECT 37.208 209.804 65.576 210.708 ; 
        RECT 31.88 209.804 37.136 210.708 ; 
        RECT 29 206.334 31.52 210.708 ; 
        RECT 0.56 209.804 28.928 210.708 ; 
        RECT 0.02 206.334 0.488 210.708 ; 
        RECT 65.504 206.334 66.116 209.996 ; 
        RECT 37.424 206.334 65.432 210.708 ; 
        RECT 34.436 206.334 37.352 209.996 ; 
        RECT 33.788 207.116 34.292 210.708 ; 
        RECT 28.784 206.732 33.68 209.996 ; 
        RECT 0.704 206.334 28.712 210.708 ; 
        RECT 0.02 206.334 0.632 209.996 ; 
        RECT 34.22 206.334 66.116 209.612 ; 
        RECT 0.02 206.732 34.148 209.612 ; 
        RECT 33.32 206.334 66.116 207.02 ; 
        RECT 0.02 206.334 33.248 209.612 ; 
        RECT 0.02 206.334 66.116 206.636 ; 
        RECT 0.02 214.508 66.116 215.028 ; 
        RECT 65.648 210.654 66.116 215.028 ; 
        RECT 37.208 214.124 65.576 215.028 ; 
        RECT 31.88 214.124 37.136 215.028 ; 
        RECT 29 210.654 31.52 215.028 ; 
        RECT 0.56 214.124 28.928 215.028 ; 
        RECT 0.02 210.654 0.488 215.028 ; 
        RECT 65.504 210.654 66.116 214.316 ; 
        RECT 37.424 210.654 65.432 215.028 ; 
        RECT 34.436 210.654 37.352 214.316 ; 
        RECT 33.788 211.436 34.292 215.028 ; 
        RECT 28.784 211.052 33.68 214.316 ; 
        RECT 0.704 210.654 28.712 215.028 ; 
        RECT 0.02 210.654 0.632 214.316 ; 
        RECT 34.22 210.654 66.116 213.932 ; 
        RECT 0.02 211.052 34.148 213.932 ; 
        RECT 33.32 210.654 66.116 211.34 ; 
        RECT 0.02 210.654 33.248 213.932 ; 
        RECT 0.02 210.654 66.116 210.956 ; 
        RECT 0.02 218.828 66.116 219.348 ; 
        RECT 65.648 214.974 66.116 219.348 ; 
        RECT 37.208 218.444 65.576 219.348 ; 
        RECT 31.88 218.444 37.136 219.348 ; 
        RECT 29 214.974 31.52 219.348 ; 
        RECT 0.56 218.444 28.928 219.348 ; 
        RECT 0.02 214.974 0.488 219.348 ; 
        RECT 65.504 214.974 66.116 218.636 ; 
        RECT 37.424 214.974 65.432 219.348 ; 
        RECT 34.436 214.974 37.352 218.636 ; 
        RECT 33.788 215.756 34.292 219.348 ; 
        RECT 28.784 215.372 33.68 218.636 ; 
        RECT 0.704 214.974 28.712 219.348 ; 
        RECT 0.02 214.974 0.632 218.636 ; 
        RECT 34.22 214.974 66.116 218.252 ; 
        RECT 0.02 215.372 34.148 218.252 ; 
        RECT 33.32 214.974 66.116 215.66 ; 
        RECT 0.02 214.974 33.248 218.252 ; 
        RECT 0.02 214.974 66.116 215.276 ; 
        RECT 0.02 223.148 66.116 223.668 ; 
        RECT 65.648 219.294 66.116 223.668 ; 
        RECT 37.208 222.764 65.576 223.668 ; 
        RECT 31.88 222.764 37.136 223.668 ; 
        RECT 29 219.294 31.52 223.668 ; 
        RECT 0.56 222.764 28.928 223.668 ; 
        RECT 0.02 219.294 0.488 223.668 ; 
        RECT 65.504 219.294 66.116 222.956 ; 
        RECT 37.424 219.294 65.432 223.668 ; 
        RECT 34.436 219.294 37.352 222.956 ; 
        RECT 33.788 220.076 34.292 223.668 ; 
        RECT 28.784 219.692 33.68 222.956 ; 
        RECT 0.704 219.294 28.712 223.668 ; 
        RECT 0.02 219.294 0.632 222.956 ; 
        RECT 34.22 219.294 66.116 222.572 ; 
        RECT 0.02 219.692 34.148 222.572 ; 
        RECT 33.32 219.294 66.116 219.98 ; 
        RECT 0.02 219.294 33.248 222.572 ; 
        RECT 0.02 219.294 66.116 219.596 ; 
        RECT 0.02 227.468 66.116 227.988 ; 
        RECT 65.648 223.614 66.116 227.988 ; 
        RECT 37.208 227.084 65.576 227.988 ; 
        RECT 31.88 227.084 37.136 227.988 ; 
        RECT 29 223.614 31.52 227.988 ; 
        RECT 0.56 227.084 28.928 227.988 ; 
        RECT 0.02 223.614 0.488 227.988 ; 
        RECT 65.504 223.614 66.116 227.276 ; 
        RECT 37.424 223.614 65.432 227.988 ; 
        RECT 34.436 223.614 37.352 227.276 ; 
        RECT 33.788 224.396 34.292 227.988 ; 
        RECT 28.784 224.012 33.68 227.276 ; 
        RECT 0.704 223.614 28.712 227.988 ; 
        RECT 0.02 223.614 0.632 227.276 ; 
        RECT 34.22 223.614 66.116 226.892 ; 
        RECT 0.02 224.012 34.148 226.892 ; 
        RECT 33.32 223.614 66.116 224.3 ; 
        RECT 0.02 223.614 33.248 226.892 ; 
        RECT 0.02 223.614 66.116 223.916 ; 
        RECT 0.02 231.788 66.116 232.308 ; 
        RECT 65.648 227.934 66.116 232.308 ; 
        RECT 37.208 231.404 65.576 232.308 ; 
        RECT 31.88 231.404 37.136 232.308 ; 
        RECT 29 227.934 31.52 232.308 ; 
        RECT 0.56 231.404 28.928 232.308 ; 
        RECT 0.02 227.934 0.488 232.308 ; 
        RECT 65.504 227.934 66.116 231.596 ; 
        RECT 37.424 227.934 65.432 232.308 ; 
        RECT 34.436 227.934 37.352 231.596 ; 
        RECT 33.788 228.716 34.292 232.308 ; 
        RECT 28.784 228.332 33.68 231.596 ; 
        RECT 0.704 227.934 28.712 232.308 ; 
        RECT 0.02 227.934 0.632 231.596 ; 
        RECT 34.22 227.934 66.116 231.212 ; 
        RECT 0.02 228.332 34.148 231.212 ; 
        RECT 33.32 227.934 66.116 228.62 ; 
        RECT 0.02 227.934 33.248 231.212 ; 
        RECT 0.02 227.934 66.116 228.236 ; 
        RECT 0.02 236.108 66.116 236.628 ; 
        RECT 65.648 232.254 66.116 236.628 ; 
        RECT 37.208 235.724 65.576 236.628 ; 
        RECT 31.88 235.724 37.136 236.628 ; 
        RECT 29 232.254 31.52 236.628 ; 
        RECT 0.56 235.724 28.928 236.628 ; 
        RECT 0.02 232.254 0.488 236.628 ; 
        RECT 65.504 232.254 66.116 235.916 ; 
        RECT 37.424 232.254 65.432 236.628 ; 
        RECT 34.436 232.254 37.352 235.916 ; 
        RECT 33.788 233.036 34.292 236.628 ; 
        RECT 28.784 232.652 33.68 235.916 ; 
        RECT 0.704 232.254 28.712 236.628 ; 
        RECT 0.02 232.254 0.632 235.916 ; 
        RECT 34.22 232.254 66.116 235.532 ; 
        RECT 0.02 232.652 34.148 235.532 ; 
        RECT 33.32 232.254 66.116 232.94 ; 
        RECT 0.02 232.254 33.248 235.532 ; 
        RECT 0.02 232.254 66.116 232.556 ; 
        RECT 0.02 240.428 66.116 240.948 ; 
        RECT 65.648 236.574 66.116 240.948 ; 
        RECT 37.208 240.044 65.576 240.948 ; 
        RECT 31.88 240.044 37.136 240.948 ; 
        RECT 29 236.574 31.52 240.948 ; 
        RECT 0.56 240.044 28.928 240.948 ; 
        RECT 0.02 236.574 0.488 240.948 ; 
        RECT 65.504 236.574 66.116 240.236 ; 
        RECT 37.424 236.574 65.432 240.948 ; 
        RECT 34.436 236.574 37.352 240.236 ; 
        RECT 33.788 237.356 34.292 240.948 ; 
        RECT 28.784 236.972 33.68 240.236 ; 
        RECT 0.704 236.574 28.712 240.948 ; 
        RECT 0.02 236.574 0.632 240.236 ; 
        RECT 34.22 236.574 66.116 239.852 ; 
        RECT 0.02 236.972 34.148 239.852 ; 
        RECT 33.32 236.574 66.116 237.26 ; 
        RECT 0.02 236.574 33.248 239.852 ; 
        RECT 0.02 236.574 66.116 236.876 ; 
        RECT 0.02 244.748 66.116 245.268 ; 
        RECT 65.648 240.894 66.116 245.268 ; 
        RECT 37.208 244.364 65.576 245.268 ; 
        RECT 31.88 244.364 37.136 245.268 ; 
        RECT 29 240.894 31.52 245.268 ; 
        RECT 0.56 244.364 28.928 245.268 ; 
        RECT 0.02 240.894 0.488 245.268 ; 
        RECT 65.504 240.894 66.116 244.556 ; 
        RECT 37.424 240.894 65.432 245.268 ; 
        RECT 34.436 240.894 37.352 244.556 ; 
        RECT 33.788 241.676 34.292 245.268 ; 
        RECT 28.784 241.292 33.68 244.556 ; 
        RECT 0.704 240.894 28.712 245.268 ; 
        RECT 0.02 240.894 0.632 244.556 ; 
        RECT 34.22 240.894 66.116 244.172 ; 
        RECT 0.02 241.292 34.148 244.172 ; 
        RECT 33.32 240.894 66.116 241.58 ; 
        RECT 0.02 240.894 33.248 244.172 ; 
        RECT 0.02 240.894 66.116 241.196 ; 
        RECT 0.02 249.068 66.116 249.588 ; 
        RECT 65.648 245.214 66.116 249.588 ; 
        RECT 37.208 248.684 65.576 249.588 ; 
        RECT 31.88 248.684 37.136 249.588 ; 
        RECT 29 245.214 31.52 249.588 ; 
        RECT 0.56 248.684 28.928 249.588 ; 
        RECT 0.02 245.214 0.488 249.588 ; 
        RECT 65.504 245.214 66.116 248.876 ; 
        RECT 37.424 245.214 65.432 249.588 ; 
        RECT 34.436 245.214 37.352 248.876 ; 
        RECT 33.788 245.996 34.292 249.588 ; 
        RECT 28.784 245.612 33.68 248.876 ; 
        RECT 0.704 245.214 28.712 249.588 ; 
        RECT 0.02 245.214 0.632 248.876 ; 
        RECT 34.22 245.214 66.116 248.492 ; 
        RECT 0.02 245.612 34.148 248.492 ; 
        RECT 33.32 245.214 66.116 245.9 ; 
        RECT 0.02 245.214 33.248 248.492 ; 
        RECT 0.02 245.214 66.116 245.516 ; 
        RECT 0.02 253.388 66.116 253.908 ; 
        RECT 65.648 249.534 66.116 253.908 ; 
        RECT 37.208 253.004 65.576 253.908 ; 
        RECT 31.88 253.004 37.136 253.908 ; 
        RECT 29 249.534 31.52 253.908 ; 
        RECT 0.56 253.004 28.928 253.908 ; 
        RECT 0.02 249.534 0.488 253.908 ; 
        RECT 65.504 249.534 66.116 253.196 ; 
        RECT 37.424 249.534 65.432 253.908 ; 
        RECT 34.436 249.534 37.352 253.196 ; 
        RECT 33.788 250.316 34.292 253.908 ; 
        RECT 28.784 249.932 33.68 253.196 ; 
        RECT 0.704 249.534 28.712 253.908 ; 
        RECT 0.02 249.534 0.632 253.196 ; 
        RECT 34.22 249.534 66.116 252.812 ; 
        RECT 0.02 249.932 34.148 252.812 ; 
        RECT 33.32 249.534 66.116 250.22 ; 
        RECT 0.02 249.534 33.248 252.812 ; 
        RECT 0.02 249.534 66.116 249.836 ; 
        RECT 0.02 257.708 66.116 258.228 ; 
        RECT 65.648 253.854 66.116 258.228 ; 
        RECT 37.208 257.324 65.576 258.228 ; 
        RECT 31.88 257.324 37.136 258.228 ; 
        RECT 29 253.854 31.52 258.228 ; 
        RECT 0.56 257.324 28.928 258.228 ; 
        RECT 0.02 253.854 0.488 258.228 ; 
        RECT 65.504 253.854 66.116 257.516 ; 
        RECT 37.424 253.854 65.432 258.228 ; 
        RECT 34.436 253.854 37.352 257.516 ; 
        RECT 33.788 254.636 34.292 258.228 ; 
        RECT 28.784 254.252 33.68 257.516 ; 
        RECT 0.704 253.854 28.712 258.228 ; 
        RECT 0.02 253.854 0.632 257.516 ; 
        RECT 34.22 253.854 66.116 257.132 ; 
        RECT 0.02 254.252 34.148 257.132 ; 
        RECT 33.32 253.854 66.116 254.54 ; 
        RECT 0.02 253.854 33.248 257.132 ; 
        RECT 0.02 253.854 66.116 254.156 ; 
        RECT 0.02 262.028 66.116 262.548 ; 
        RECT 65.648 258.174 66.116 262.548 ; 
        RECT 37.208 261.644 65.576 262.548 ; 
        RECT 31.88 261.644 37.136 262.548 ; 
        RECT 29 258.174 31.52 262.548 ; 
        RECT 0.56 261.644 28.928 262.548 ; 
        RECT 0.02 258.174 0.488 262.548 ; 
        RECT 65.504 258.174 66.116 261.836 ; 
        RECT 37.424 258.174 65.432 262.548 ; 
        RECT 34.436 258.174 37.352 261.836 ; 
        RECT 33.788 258.956 34.292 262.548 ; 
        RECT 28.784 258.572 33.68 261.836 ; 
        RECT 0.704 258.174 28.712 262.548 ; 
        RECT 0.02 258.174 0.632 261.836 ; 
        RECT 34.22 258.174 66.116 261.452 ; 
        RECT 0.02 258.572 34.148 261.452 ; 
        RECT 33.32 258.174 66.116 258.86 ; 
        RECT 0.02 258.174 33.248 261.452 ; 
        RECT 0.02 258.174 66.116 258.476 ; 
        RECT 0.02 266.348 66.116 266.868 ; 
        RECT 65.648 262.494 66.116 266.868 ; 
        RECT 37.208 265.964 65.576 266.868 ; 
        RECT 31.88 265.964 37.136 266.868 ; 
        RECT 29 262.494 31.52 266.868 ; 
        RECT 0.56 265.964 28.928 266.868 ; 
        RECT 0.02 262.494 0.488 266.868 ; 
        RECT 65.504 262.494 66.116 266.156 ; 
        RECT 37.424 262.494 65.432 266.868 ; 
        RECT 34.436 262.494 37.352 266.156 ; 
        RECT 33.788 263.276 34.292 266.868 ; 
        RECT 28.784 262.892 33.68 266.156 ; 
        RECT 0.704 262.494 28.712 266.868 ; 
        RECT 0.02 262.494 0.632 266.156 ; 
        RECT 34.22 262.494 66.116 265.772 ; 
        RECT 0.02 262.892 34.148 265.772 ; 
        RECT 33.32 262.494 66.116 263.18 ; 
        RECT 0.02 262.494 33.248 265.772 ; 
        RECT 0.02 262.494 66.116 262.796 ; 
        RECT 0.02 270.668 66.116 271.188 ; 
        RECT 65.648 266.814 66.116 271.188 ; 
        RECT 37.208 270.284 65.576 271.188 ; 
        RECT 31.88 270.284 37.136 271.188 ; 
        RECT 29 266.814 31.52 271.188 ; 
        RECT 0.56 270.284 28.928 271.188 ; 
        RECT 0.02 266.814 0.488 271.188 ; 
        RECT 65.504 266.814 66.116 270.476 ; 
        RECT 37.424 266.814 65.432 271.188 ; 
        RECT 34.436 266.814 37.352 270.476 ; 
        RECT 33.788 267.596 34.292 271.188 ; 
        RECT 28.784 267.212 33.68 270.476 ; 
        RECT 0.704 266.814 28.712 271.188 ; 
        RECT 0.02 266.814 0.632 270.476 ; 
        RECT 34.22 266.814 66.116 270.092 ; 
        RECT 0.02 267.212 34.148 270.092 ; 
        RECT 33.32 266.814 66.116 267.5 ; 
        RECT 0.02 266.814 33.248 270.092 ; 
        RECT 0.02 266.814 66.116 267.116 ; 
        RECT 0.02 274.988 66.116 275.508 ; 
        RECT 65.648 271.134 66.116 275.508 ; 
        RECT 37.208 274.604 65.576 275.508 ; 
        RECT 31.88 274.604 37.136 275.508 ; 
        RECT 29 271.134 31.52 275.508 ; 
        RECT 0.56 274.604 28.928 275.508 ; 
        RECT 0.02 271.134 0.488 275.508 ; 
        RECT 65.504 271.134 66.116 274.796 ; 
        RECT 37.424 271.134 65.432 275.508 ; 
        RECT 34.436 271.134 37.352 274.796 ; 
        RECT 33.788 271.916 34.292 275.508 ; 
        RECT 28.784 271.532 33.68 274.796 ; 
        RECT 0.704 271.134 28.712 275.508 ; 
        RECT 0.02 271.134 0.632 274.796 ; 
        RECT 34.22 271.134 66.116 274.412 ; 
        RECT 0.02 271.532 34.148 274.412 ; 
        RECT 33.32 271.134 66.116 271.82 ; 
        RECT 0.02 271.134 33.248 274.412 ; 
        RECT 0.02 271.134 66.116 271.436 ; 
        RECT 0.02 279.308 66.116 279.828 ; 
        RECT 65.648 275.454 66.116 279.828 ; 
        RECT 37.208 278.924 65.576 279.828 ; 
        RECT 31.88 278.924 37.136 279.828 ; 
        RECT 29 275.454 31.52 279.828 ; 
        RECT 0.56 278.924 28.928 279.828 ; 
        RECT 0.02 275.454 0.488 279.828 ; 
        RECT 65.504 275.454 66.116 279.116 ; 
        RECT 37.424 275.454 65.432 279.828 ; 
        RECT 34.436 275.454 37.352 279.116 ; 
        RECT 33.788 276.236 34.292 279.828 ; 
        RECT 28.784 275.852 33.68 279.116 ; 
        RECT 0.704 275.454 28.712 279.828 ; 
        RECT 0.02 275.454 0.632 279.116 ; 
        RECT 34.22 275.454 66.116 278.732 ; 
        RECT 0.02 275.852 34.148 278.732 ; 
        RECT 33.32 275.454 66.116 276.14 ; 
        RECT 0.02 275.454 33.248 278.732 ; 
        RECT 0.02 275.454 66.116 275.756 ; 
        RECT 0.02 283.628 66.116 284.148 ; 
        RECT 65.648 279.774 66.116 284.148 ; 
        RECT 37.208 283.244 65.576 284.148 ; 
        RECT 31.88 283.244 37.136 284.148 ; 
        RECT 29 279.774 31.52 284.148 ; 
        RECT 0.56 283.244 28.928 284.148 ; 
        RECT 0.02 279.774 0.488 284.148 ; 
        RECT 65.504 279.774 66.116 283.436 ; 
        RECT 37.424 279.774 65.432 284.148 ; 
        RECT 34.436 279.774 37.352 283.436 ; 
        RECT 33.788 280.556 34.292 284.148 ; 
        RECT 28.784 280.172 33.68 283.436 ; 
        RECT 0.704 279.774 28.712 284.148 ; 
        RECT 0.02 279.774 0.632 283.436 ; 
        RECT 34.22 279.774 66.116 283.052 ; 
        RECT 0.02 280.172 34.148 283.052 ; 
        RECT 33.32 279.774 66.116 280.46 ; 
        RECT 0.02 279.774 33.248 283.052 ; 
        RECT 0.02 279.774 66.116 280.076 ; 
        RECT 0.02 287.948 66.116 288.468 ; 
        RECT 65.648 284.094 66.116 288.468 ; 
        RECT 37.208 287.564 65.576 288.468 ; 
        RECT 31.88 287.564 37.136 288.468 ; 
        RECT 29 284.094 31.52 288.468 ; 
        RECT 0.56 287.564 28.928 288.468 ; 
        RECT 0.02 284.094 0.488 288.468 ; 
        RECT 65.504 284.094 66.116 287.756 ; 
        RECT 37.424 284.094 65.432 288.468 ; 
        RECT 34.436 284.094 37.352 287.756 ; 
        RECT 33.788 284.876 34.292 288.468 ; 
        RECT 28.784 284.492 33.68 287.756 ; 
        RECT 0.704 284.094 28.712 288.468 ; 
        RECT 0.02 284.094 0.632 287.756 ; 
        RECT 34.22 284.094 66.116 287.372 ; 
        RECT 0.02 284.492 34.148 287.372 ; 
        RECT 33.32 284.094 66.116 284.78 ; 
        RECT 0.02 284.094 33.248 287.372 ; 
        RECT 0.02 284.094 66.116 284.396 ; 
        RECT 0.02 292.268 66.116 292.788 ; 
        RECT 65.648 288.414 66.116 292.788 ; 
        RECT 37.208 291.884 65.576 292.788 ; 
        RECT 31.88 291.884 37.136 292.788 ; 
        RECT 29 288.414 31.52 292.788 ; 
        RECT 0.56 291.884 28.928 292.788 ; 
        RECT 0.02 288.414 0.488 292.788 ; 
        RECT 65.504 288.414 66.116 292.076 ; 
        RECT 37.424 288.414 65.432 292.788 ; 
        RECT 34.436 288.414 37.352 292.076 ; 
        RECT 33.788 289.196 34.292 292.788 ; 
        RECT 28.784 288.812 33.68 292.076 ; 
        RECT 0.704 288.414 28.712 292.788 ; 
        RECT 0.02 288.414 0.632 292.076 ; 
        RECT 34.22 288.414 66.116 291.692 ; 
        RECT 0.02 288.812 34.148 291.692 ; 
        RECT 33.32 288.414 66.116 289.1 ; 
        RECT 0.02 288.414 33.248 291.692 ; 
        RECT 0.02 288.414 66.116 288.716 ; 
        RECT 0.02 296.588 66.116 297.108 ; 
        RECT 65.648 292.734 66.116 297.108 ; 
        RECT 37.208 296.204 65.576 297.108 ; 
        RECT 31.88 296.204 37.136 297.108 ; 
        RECT 29 292.734 31.52 297.108 ; 
        RECT 0.56 296.204 28.928 297.108 ; 
        RECT 0.02 292.734 0.488 297.108 ; 
        RECT 65.504 292.734 66.116 296.396 ; 
        RECT 37.424 292.734 65.432 297.108 ; 
        RECT 34.436 292.734 37.352 296.396 ; 
        RECT 33.788 293.516 34.292 297.108 ; 
        RECT 28.784 293.132 33.68 296.396 ; 
        RECT 0.704 292.734 28.712 297.108 ; 
        RECT 0.02 292.734 0.632 296.396 ; 
        RECT 34.22 292.734 66.116 296.012 ; 
        RECT 0.02 293.132 34.148 296.012 ; 
        RECT 33.32 292.734 66.116 293.42 ; 
        RECT 0.02 292.734 33.248 296.012 ; 
        RECT 0.02 292.734 66.116 293.036 ; 
        RECT 0.02 300.908 66.116 301.428 ; 
        RECT 65.648 297.054 66.116 301.428 ; 
        RECT 37.208 300.524 65.576 301.428 ; 
        RECT 31.88 300.524 37.136 301.428 ; 
        RECT 29 297.054 31.52 301.428 ; 
        RECT 0.56 300.524 28.928 301.428 ; 
        RECT 0.02 297.054 0.488 301.428 ; 
        RECT 65.504 297.054 66.116 300.716 ; 
        RECT 37.424 297.054 65.432 301.428 ; 
        RECT 34.436 297.054 37.352 300.716 ; 
        RECT 33.788 297.836 34.292 301.428 ; 
        RECT 28.784 297.452 33.68 300.716 ; 
        RECT 0.704 297.054 28.712 301.428 ; 
        RECT 0.02 297.054 0.632 300.716 ; 
        RECT 34.22 297.054 66.116 300.332 ; 
        RECT 0.02 297.452 34.148 300.332 ; 
        RECT 33.32 297.054 66.116 297.74 ; 
        RECT 0.02 297.054 33.248 300.332 ; 
        RECT 0.02 297.054 66.116 297.356 ; 
        RECT 0.02 305.228 66.116 305.748 ; 
        RECT 65.648 301.374 66.116 305.748 ; 
        RECT 37.208 304.844 65.576 305.748 ; 
        RECT 31.88 304.844 37.136 305.748 ; 
        RECT 29 301.374 31.52 305.748 ; 
        RECT 0.56 304.844 28.928 305.748 ; 
        RECT 0.02 301.374 0.488 305.748 ; 
        RECT 65.504 301.374 66.116 305.036 ; 
        RECT 37.424 301.374 65.432 305.748 ; 
        RECT 34.436 301.374 37.352 305.036 ; 
        RECT 33.788 302.156 34.292 305.748 ; 
        RECT 28.784 301.772 33.68 305.036 ; 
        RECT 0.704 301.374 28.712 305.748 ; 
        RECT 0.02 301.374 0.632 305.036 ; 
        RECT 34.22 301.374 66.116 304.652 ; 
        RECT 0.02 301.772 34.148 304.652 ; 
        RECT 33.32 301.374 66.116 302.06 ; 
        RECT 0.02 301.374 33.248 304.652 ; 
        RECT 0.02 301.374 66.116 301.676 ; 
        RECT 0.02 309.548 66.116 310.068 ; 
        RECT 65.648 305.694 66.116 310.068 ; 
        RECT 37.208 309.164 65.576 310.068 ; 
        RECT 31.88 309.164 37.136 310.068 ; 
        RECT 29 305.694 31.52 310.068 ; 
        RECT 0.56 309.164 28.928 310.068 ; 
        RECT 0.02 305.694 0.488 310.068 ; 
        RECT 65.504 305.694 66.116 309.356 ; 
        RECT 37.424 305.694 65.432 310.068 ; 
        RECT 34.436 305.694 37.352 309.356 ; 
        RECT 33.788 306.476 34.292 310.068 ; 
        RECT 28.784 306.092 33.68 309.356 ; 
        RECT 0.704 305.694 28.712 310.068 ; 
        RECT 0.02 305.694 0.632 309.356 ; 
        RECT 34.22 305.694 66.116 308.972 ; 
        RECT 0.02 306.092 34.148 308.972 ; 
        RECT 33.32 305.694 66.116 306.38 ; 
        RECT 0.02 305.694 33.248 308.972 ; 
        RECT 0.02 305.694 66.116 305.996 ; 
        RECT 0.02 313.868 66.116 314.388 ; 
        RECT 65.648 310.014 66.116 314.388 ; 
        RECT 37.208 313.484 65.576 314.388 ; 
        RECT 31.88 313.484 37.136 314.388 ; 
        RECT 29 310.014 31.52 314.388 ; 
        RECT 0.56 313.484 28.928 314.388 ; 
        RECT 0.02 310.014 0.488 314.388 ; 
        RECT 65.504 310.014 66.116 313.676 ; 
        RECT 37.424 310.014 65.432 314.388 ; 
        RECT 34.436 310.014 37.352 313.676 ; 
        RECT 33.788 310.796 34.292 314.388 ; 
        RECT 28.784 310.412 33.68 313.676 ; 
        RECT 0.704 310.014 28.712 314.388 ; 
        RECT 0.02 310.014 0.632 313.676 ; 
        RECT 34.22 310.014 66.116 313.292 ; 
        RECT 0.02 310.412 34.148 313.292 ; 
        RECT 33.32 310.014 66.116 310.7 ; 
        RECT 0.02 310.014 33.248 313.292 ; 
        RECT 0.02 310.014 66.116 310.316 ; 
        RECT 0.02 318.188 66.116 318.708 ; 
        RECT 65.648 314.334 66.116 318.708 ; 
        RECT 37.208 317.804 65.576 318.708 ; 
        RECT 31.88 317.804 37.136 318.708 ; 
        RECT 29 314.334 31.52 318.708 ; 
        RECT 0.56 317.804 28.928 318.708 ; 
        RECT 0.02 314.334 0.488 318.708 ; 
        RECT 65.504 314.334 66.116 317.996 ; 
        RECT 37.424 314.334 65.432 318.708 ; 
        RECT 34.436 314.334 37.352 317.996 ; 
        RECT 33.788 315.116 34.292 318.708 ; 
        RECT 28.784 314.732 33.68 317.996 ; 
        RECT 0.704 314.334 28.712 318.708 ; 
        RECT 0.02 314.334 0.632 317.996 ; 
        RECT 34.22 314.334 66.116 317.612 ; 
        RECT 0.02 314.732 34.148 317.612 ; 
        RECT 33.32 314.334 66.116 315.02 ; 
        RECT 0.02 314.334 33.248 317.612 ; 
        RECT 0.02 314.334 66.116 314.636 ; 
        RECT 0.02 322.508 66.116 323.028 ; 
        RECT 65.648 318.654 66.116 323.028 ; 
        RECT 37.208 322.124 65.576 323.028 ; 
        RECT 31.88 322.124 37.136 323.028 ; 
        RECT 29 318.654 31.52 323.028 ; 
        RECT 0.56 322.124 28.928 323.028 ; 
        RECT 0.02 318.654 0.488 323.028 ; 
        RECT 65.504 318.654 66.116 322.316 ; 
        RECT 37.424 318.654 65.432 323.028 ; 
        RECT 34.436 318.654 37.352 322.316 ; 
        RECT 33.788 319.436 34.292 323.028 ; 
        RECT 28.784 319.052 33.68 322.316 ; 
        RECT 0.704 318.654 28.712 323.028 ; 
        RECT 0.02 318.654 0.632 322.316 ; 
        RECT 34.22 318.654 66.116 321.932 ; 
        RECT 0.02 319.052 34.148 321.932 ; 
        RECT 33.32 318.654 66.116 319.34 ; 
        RECT 0.02 318.654 33.248 321.932 ; 
        RECT 0.02 318.654 66.116 318.956 ; 
        RECT 0.02 326.828 66.116 327.348 ; 
        RECT 65.648 322.974 66.116 327.348 ; 
        RECT 37.208 326.444 65.576 327.348 ; 
        RECT 31.88 326.444 37.136 327.348 ; 
        RECT 29 322.974 31.52 327.348 ; 
        RECT 0.56 326.444 28.928 327.348 ; 
        RECT 0.02 322.974 0.488 327.348 ; 
        RECT 65.504 322.974 66.116 326.636 ; 
        RECT 37.424 322.974 65.432 327.348 ; 
        RECT 34.436 322.974 37.352 326.636 ; 
        RECT 33.788 323.756 34.292 327.348 ; 
        RECT 28.784 323.372 33.68 326.636 ; 
        RECT 0.704 322.974 28.712 327.348 ; 
        RECT 0.02 322.974 0.632 326.636 ; 
        RECT 34.22 322.974 66.116 326.252 ; 
        RECT 0.02 323.372 34.148 326.252 ; 
        RECT 33.32 322.974 66.116 323.66 ; 
        RECT 0.02 322.974 33.248 326.252 ; 
        RECT 0.02 322.974 66.116 323.276 ; 
        RECT 0.02 331.148 66.116 331.668 ; 
        RECT 65.648 327.294 66.116 331.668 ; 
        RECT 37.208 330.764 65.576 331.668 ; 
        RECT 31.88 330.764 37.136 331.668 ; 
        RECT 29 327.294 31.52 331.668 ; 
        RECT 0.56 330.764 28.928 331.668 ; 
        RECT 0.02 327.294 0.488 331.668 ; 
        RECT 65.504 327.294 66.116 330.956 ; 
        RECT 37.424 327.294 65.432 331.668 ; 
        RECT 34.436 327.294 37.352 330.956 ; 
        RECT 33.788 328.076 34.292 331.668 ; 
        RECT 28.784 327.692 33.68 330.956 ; 
        RECT 0.704 327.294 28.712 331.668 ; 
        RECT 0.02 327.294 0.632 330.956 ; 
        RECT 34.22 327.294 66.116 330.572 ; 
        RECT 0.02 327.692 34.148 330.572 ; 
        RECT 33.32 327.294 66.116 327.98 ; 
        RECT 0.02 327.294 33.248 330.572 ; 
        RECT 0.02 327.294 66.116 327.596 ; 
        RECT 0.02 335.468 66.116 335.988 ; 
        RECT 65.648 331.614 66.116 335.988 ; 
        RECT 37.208 335.084 65.576 335.988 ; 
        RECT 31.88 335.084 37.136 335.988 ; 
        RECT 29 331.614 31.52 335.988 ; 
        RECT 0.56 335.084 28.928 335.988 ; 
        RECT 0.02 331.614 0.488 335.988 ; 
        RECT 65.504 331.614 66.116 335.276 ; 
        RECT 37.424 331.614 65.432 335.988 ; 
        RECT 34.436 331.614 37.352 335.276 ; 
        RECT 33.788 332.396 34.292 335.988 ; 
        RECT 28.784 332.012 33.68 335.276 ; 
        RECT 0.704 331.614 28.712 335.988 ; 
        RECT 0.02 331.614 0.632 335.276 ; 
        RECT 34.22 331.614 66.116 334.892 ; 
        RECT 0.02 332.012 34.148 334.892 ; 
        RECT 33.32 331.614 66.116 332.3 ; 
        RECT 0.02 331.614 33.248 334.892 ; 
        RECT 0.02 331.614 66.116 331.916 ; 
        RECT 0.02 339.788 66.116 340.308 ; 
        RECT 65.648 335.934 66.116 340.308 ; 
        RECT 37.208 339.404 65.576 340.308 ; 
        RECT 31.88 339.404 37.136 340.308 ; 
        RECT 29 335.934 31.52 340.308 ; 
        RECT 0.56 339.404 28.928 340.308 ; 
        RECT 0.02 335.934 0.488 340.308 ; 
        RECT 65.504 335.934 66.116 339.596 ; 
        RECT 37.424 335.934 65.432 340.308 ; 
        RECT 34.436 335.934 37.352 339.596 ; 
        RECT 33.788 336.716 34.292 340.308 ; 
        RECT 28.784 336.332 33.68 339.596 ; 
        RECT 0.704 335.934 28.712 340.308 ; 
        RECT 0.02 335.934 0.632 339.596 ; 
        RECT 34.22 335.934 66.116 339.212 ; 
        RECT 0.02 336.332 34.148 339.212 ; 
        RECT 33.32 335.934 66.116 336.62 ; 
        RECT 0.02 335.934 33.248 339.212 ; 
        RECT 0.02 335.934 66.116 336.236 ; 
        RECT 0.02 344.108 66.116 344.628 ; 
        RECT 65.648 340.254 66.116 344.628 ; 
        RECT 37.208 343.724 65.576 344.628 ; 
        RECT 31.88 343.724 37.136 344.628 ; 
        RECT 29 340.254 31.52 344.628 ; 
        RECT 0.56 343.724 28.928 344.628 ; 
        RECT 0.02 340.254 0.488 344.628 ; 
        RECT 65.504 340.254 66.116 343.916 ; 
        RECT 37.424 340.254 65.432 344.628 ; 
        RECT 34.436 340.254 37.352 343.916 ; 
        RECT 33.788 341.036 34.292 344.628 ; 
        RECT 28.784 340.652 33.68 343.916 ; 
        RECT 0.704 340.254 28.712 344.628 ; 
        RECT 0.02 340.254 0.632 343.916 ; 
        RECT 34.22 340.254 66.116 343.532 ; 
        RECT 0.02 340.652 34.148 343.532 ; 
        RECT 33.32 340.254 66.116 340.94 ; 
        RECT 0.02 340.254 33.248 343.532 ; 
        RECT 0.02 340.254 66.116 340.556 ; 
        RECT 0.02 348.428 66.116 348.948 ; 
        RECT 65.648 344.574 66.116 348.948 ; 
        RECT 37.208 348.044 65.576 348.948 ; 
        RECT 31.88 348.044 37.136 348.948 ; 
        RECT 29 344.574 31.52 348.948 ; 
        RECT 0.56 348.044 28.928 348.948 ; 
        RECT 0.02 344.574 0.488 348.948 ; 
        RECT 65.504 344.574 66.116 348.236 ; 
        RECT 37.424 344.574 65.432 348.948 ; 
        RECT 34.436 344.574 37.352 348.236 ; 
        RECT 33.788 345.356 34.292 348.948 ; 
        RECT 28.784 344.972 33.68 348.236 ; 
        RECT 0.704 344.574 28.712 348.948 ; 
        RECT 0.02 344.574 0.632 348.236 ; 
        RECT 34.22 344.574 66.116 347.852 ; 
        RECT 0.02 344.972 34.148 347.852 ; 
        RECT 33.32 344.574 66.116 345.26 ; 
        RECT 0.02 344.574 33.248 347.852 ; 
        RECT 0.02 344.574 66.116 344.876 ; 
        RECT 0.02 352.748 66.116 353.268 ; 
        RECT 65.648 348.894 66.116 353.268 ; 
        RECT 37.208 352.364 65.576 353.268 ; 
        RECT 31.88 352.364 37.136 353.268 ; 
        RECT 29 348.894 31.52 353.268 ; 
        RECT 0.56 352.364 28.928 353.268 ; 
        RECT 0.02 348.894 0.488 353.268 ; 
        RECT 65.504 348.894 66.116 352.556 ; 
        RECT 37.424 348.894 65.432 353.268 ; 
        RECT 34.436 348.894 37.352 352.556 ; 
        RECT 33.788 349.676 34.292 353.268 ; 
        RECT 28.784 349.292 33.68 352.556 ; 
        RECT 0.704 348.894 28.712 353.268 ; 
        RECT 0.02 348.894 0.632 352.556 ; 
        RECT 34.22 348.894 66.116 352.172 ; 
        RECT 0.02 349.292 34.148 352.172 ; 
        RECT 33.32 348.894 66.116 349.58 ; 
        RECT 0.02 348.894 33.248 352.172 ; 
        RECT 0.02 348.894 66.116 349.196 ; 
  LAYER M4 ; 
      RECT 6.276 167.64 60.038 167.736 ; 
      RECT 6.276 168.792 60.038 168.888 ; 
      RECT 6.276 170.328 60.038 170.424 ; 
      RECT 6.276 170.712 60.038 170.808 ; 
      RECT 6.276 172.056 60.038 172.152 ; 
      RECT 6.276 173.592 60.038 173.688 ; 
      RECT 43.82 163.476 44.156 163.572 ; 
      RECT 43.068 165.204 43.588 165.3 ; 
      RECT 43.1 167.834 43.568 167.93 ; 
      RECT 43.1 168.984 43.568 169.08 ; 
      RECT 40.544 165.204 42.828 165.3 ; 
      RECT 40.784 168.312 41.216 168.408 ; 
      RECT 35.452 169.812 39.824 169.908 ; 
      RECT 38.204 168.084 38.54 168.18 ; 
      RECT 35.068 172.884 38.54 172.98 ; 
      RECT 38.204 173.268 38.54 173.364 ; 
      RECT 37.492 166.164 37.828 166.26 ; 
      RECT 37.34 171.54 37.676 171.636 ; 
      RECT 37.34 174.42 37.676 174.516 ; 
      RECT 36.628 165.78 36.964 165.876 ; 
      RECT 35.772 160.628 36.824 160.724 ; 
      RECT 35.772 195.124 36.824 195.22 ; 
      RECT 35.836 171.732 36.812 171.828 ; 
      RECT 36.476 172.308 36.812 172.404 ; 
      RECT 30.652 173.268 36.812 173.364 ; 
      RECT 36.476 174.42 36.812 174.516 ; 
      RECT 35.54 194.74 36.592 194.836 ; 
      RECT 35.536 160.244 36.588 160.34 ; 
      RECT 35.384 159.86 36.436 159.956 ; 
      RECT 35.384 193.972 36.436 194.068 ; 
      RECT 36.044 176.148 36.38 176.244 ; 
      RECT 32.956 177.684 36.38 177.78 ; 
      RECT 34.492 186.708 36.38 186.804 ; 
      RECT 36.044 187.092 36.38 187.188 ; 
      RECT 35.192 159.476 36.244 159.572 ; 
      RECT 35.192 193.588 36.244 193.684 ; 
      RECT 34.3 183.06 36.08 183.156 ; 
      RECT 35.016 159.092 36.068 159.188 ; 
      RECT 35.016 194.932 36.068 195.028 ; 
      RECT 34.82 160.436 35.872 160.532 ; 
      RECT 34.82 194.548 35.872 194.644 ; 
      RECT 35.344 172.308 35.828 172.404 ; 
      RECT 35.26 180.756 35.792 180.852 ; 
      RECT 34.632 160.052 35.684 160.148 ; 
      RECT 34.632 194.164 35.684 194.26 ; 
      RECT 34.492 158.9 35.544 158.996 ; 
      RECT 34.492 193.78 35.544 193.876 ; 
      RECT 31.228 187.092 35.504 187.188 ; 
      RECT 35.168 191.7 35.504 191.796 ; 
      RECT 34.268 158.324 35.32 158.42 ; 
      RECT 34.268 193.396 35.32 193.492 ; 
      RECT 34.876 176.148 35.216 176.244 ; 
      RECT 30.46 178.452 34.928 178.548 ; 
      RECT 33.04 169.812 34.868 169.908 ; 
      RECT 32.348 161.204 33.416 161.3 ; 
      RECT 32.348 192.82 33.416 192.916 ; 
      RECT 32.896 175.956 33.332 176.052 ; 
      RECT 32.256 160.82 33.224 160.916 ; 
      RECT 32.256 195.316 33.224 195.412 ; 
      RECT 32.032 158.9 33 158.996 ; 
      RECT 32.148 195.7 33 195.796 ; 
      RECT 32.612 174.42 32.948 174.516 ; 
      RECT 31.816 159.284 32.808 159.38 ; 
      RECT 31.816 195.124 32.808 195.22 ; 
      RECT 30.88 184.788 32.564 184.884 ; 
      RECT 30.752 160.628 31.82 160.724 ; 
      RECT 30.752 195.7 31.82 195.796 ; 
      RECT 31.312 179.028 31.796 179.124 ; 
      RECT 31.28 191.7 31.616 191.796 ; 
      RECT 30.616 160.244 31.604 160.34 ; 
      RECT 30.348 193.972 31.604 194.068 ; 
      RECT 30.512 159.86 31.432 159.956 ; 
      RECT 30.464 195.316 31.432 195.412 ; 
      RECT 30.3 159.476 31.22 159.572 ; 
      RECT 30.884 185.364 31.22 185.46 ; 
      RECT 30.1 193.588 31.22 193.684 ; 
      RECT 30.12 159.092 31.04 159.188 ; 
      RECT 30.12 194.932 31.04 195.028 ; 
      RECT 26.272 174.42 31.028 174.516 ; 
      RECT 29.968 160.052 30.888 160.148 ; 
      RECT 29.968 194.548 30.888 194.644 ; 
      RECT 29.896 159.668 30.668 159.764 ; 
      RECT 29.896 194.164 30.668 194.26 ; 
      RECT 29.7 159.284 30.472 159.38 ; 
      RECT 29.7 193.78 30.472 193.876 ; 
      RECT 29.716 178.068 30.452 178.164 ; 
      RECT 29.492 158.9 30.264 158.996 ; 
      RECT 29.492 193.396 30.264 193.492 ; 
      RECT 27.556 167.316 30.26 167.412 ; 
      RECT 29.716 178.452 30.052 178.548 ; 
      RECT 28.64 161.012 29.692 161.108 ; 
      RECT 28.77 176.148 29.304 176.244 ; 
      RECT 27.404 168.084 27.74 168.18 ; 
  LAYER V4 ; 
      RECT 44.016 163.476 44.112 163.572 ; 
      RECT 44.016 167.64 44.112 167.736 ; 
      RECT 43.344 165.204 43.44 165.3 ; 
      RECT 43.344 167.834 43.44 167.93 ; 
      RECT 43.344 168.984 43.44 169.08 ; 
      RECT 40.848 165.204 40.944 165.3 ; 
      RECT 40.848 168.312 40.944 168.408 ; 
      RECT 38.4 168.084 38.496 168.18 ; 
      RECT 38.4 168.792 38.496 168.888 ; 
      RECT 38.4 172.884 38.496 172.98 ; 
      RECT 38.4 173.268 38.496 173.364 ; 
      RECT 37.536 166.164 37.632 166.26 ; 
      RECT 37.536 170.328 37.632 170.424 ; 
      RECT 37.536 171.54 37.632 171.636 ; 
      RECT 37.536 172.056 37.632 172.152 ; 
      RECT 37.536 173.592 37.632 173.688 ; 
      RECT 37.536 174.42 37.632 174.516 ; 
      RECT 36.672 165.78 36.768 165.876 ; 
      RECT 36.672 170.712 36.768 170.808 ; 
      RECT 36.672 171.732 36.768 171.828 ; 
      RECT 36.672 172.308 36.768 172.404 ; 
      RECT 36.672 173.268 36.768 173.364 ; 
      RECT 36.672 174.42 36.768 174.516 ; 
      RECT 36.24 176.148 36.336 176.244 ; 
      RECT 36.24 177.684 36.336 177.78 ; 
      RECT 36.24 186.708 36.336 186.804 ; 
      RECT 36.24 187.092 36.336 187.188 ; 
      RECT 35.88 160.628 35.976 160.724 ; 
      RECT 35.88 171.732 35.976 171.828 ; 
      RECT 35.88 195.124 35.976 195.22 ; 
      RECT 35.688 160.244 35.784 160.34 ; 
      RECT 35.688 172.308 35.784 172.404 ; 
      RECT 35.688 194.74 35.784 194.836 ; 
      RECT 35.496 159.86 35.592 159.956 ; 
      RECT 35.496 169.812 35.592 169.908 ; 
      RECT 35.496 193.972 35.592 194.068 ; 
      RECT 35.304 159.476 35.4 159.572 ; 
      RECT 35.304 180.756 35.4 180.852 ; 
      RECT 35.304 191.7 35.4 191.796 ; 
      RECT 35.304 193.588 35.4 193.684 ; 
      RECT 35.112 159.092 35.208 159.188 ; 
      RECT 35.112 172.884 35.208 172.98 ; 
      RECT 35.112 194.932 35.208 195.028 ; 
      RECT 34.92 160.436 35.016 160.532 ; 
      RECT 34.92 176.148 35.016 176.244 ; 
      RECT 34.92 194.548 35.016 194.644 ; 
      RECT 34.728 160.052 34.824 160.148 ; 
      RECT 34.728 169.812 34.824 169.908 ; 
      RECT 34.728 194.164 34.824 194.26 ; 
      RECT 34.536 158.9 34.632 158.996 ; 
      RECT 34.536 186.708 34.632 186.804 ; 
      RECT 34.536 193.78 34.632 193.876 ; 
      RECT 34.344 158.324 34.44 158.42 ; 
      RECT 34.344 183.06 34.44 183.156 ; 
      RECT 34.344 193.396 34.44 193.492 ; 
      RECT 33.192 161.204 33.288 161.3 ; 
      RECT 33.192 175.956 33.288 176.052 ; 
      RECT 33.192 192.82 33.288 192.916 ; 
      RECT 33 160.82 33.096 160.916 ; 
      RECT 33 177.684 33.096 177.78 ; 
      RECT 33 195.316 33.096 195.412 ; 
      RECT 32.808 158.9 32.904 158.996 ; 
      RECT 32.808 174.42 32.904 174.516 ; 
      RECT 32.808 195.7 32.904 195.796 ; 
      RECT 32.424 159.284 32.52 159.38 ; 
      RECT 32.424 184.788 32.52 184.884 ; 
      RECT 32.424 195.124 32.52 195.22 ; 
      RECT 31.656 160.628 31.752 160.724 ; 
      RECT 31.656 179.028 31.752 179.124 ; 
      RECT 31.656 195.7 31.752 195.796 ; 
      RECT 31.464 160.244 31.56 160.34 ; 
      RECT 31.464 191.7 31.56 191.796 ; 
      RECT 31.464 193.972 31.56 194.068 ; 
      RECT 31.272 159.86 31.368 159.956 ; 
      RECT 31.272 187.092 31.368 187.188 ; 
      RECT 31.272 195.316 31.368 195.412 ; 
      RECT 31.08 159.476 31.176 159.572 ; 
      RECT 31.08 185.364 31.176 185.46 ; 
      RECT 31.08 193.588 31.176 193.684 ; 
      RECT 30.888 159.092 30.984 159.188 ; 
      RECT 30.888 174.42 30.984 174.516 ; 
      RECT 30.888 194.932 30.984 195.028 ; 
      RECT 30.696 160.052 30.792 160.148 ; 
      RECT 30.696 173.268 30.792 173.364 ; 
      RECT 30.696 194.548 30.792 194.644 ; 
      RECT 30.504 159.668 30.6 159.764 ; 
      RECT 30.504 178.452 30.6 178.548 ; 
      RECT 30.504 194.164 30.6 194.26 ; 
      RECT 30.312 159.284 30.408 159.38 ; 
      RECT 30.312 178.068 30.408 178.164 ; 
      RECT 30.312 193.78 30.408 193.876 ; 
      RECT 30.12 158.9 30.216 158.996 ; 
      RECT 30.12 167.316 30.216 167.412 ; 
      RECT 30.12 193.396 30.216 193.492 ; 
      RECT 29.76 178.068 29.856 178.164 ; 
      RECT 29.76 178.452 29.856 178.548 ; 
      RECT 29.088 161.012 29.184 161.108 ; 
      RECT 29.088 176.148 29.184 176.244 ; 
      RECT 27.6 167.316 27.696 167.412 ; 
      RECT 27.6 168.084 27.696 168.18 ; 
  LAYER M5 ; 
      RECT 44.016 163.432 44.112 167.78 ; 
      RECT 43.344 165.092 43.44 169.334 ; 
      RECT 40.848 165.126 40.944 168.456 ; 
      RECT 38.4 168.04 38.496 168.932 ; 
      RECT 38.4 172.84 38.496 173.408 ; 
      RECT 37.536 166.12 37.632 170.468 ; 
      RECT 37.536 171.496 37.632 172.196 ; 
      RECT 37.536 173.548 37.632 174.56 ; 
      RECT 36.672 165.736 36.768 170.852 ; 
      RECT 36.672 171.688 36.768 172.448 ; 
      RECT 36.672 173.224 36.768 174.56 ; 
      RECT 36.24 176.104 36.336 177.824 ; 
      RECT 36.24 186.664 36.336 187.232 ; 
      RECT 35.88 161.976 35.976 192.308 ; 
      RECT 35.688 161.976 35.784 192.308 ; 
      RECT 35.496 161.976 35.592 192.308 ; 
      RECT 35.304 161.976 35.4 192.308 ; 
      RECT 35.112 161.976 35.208 192.308 ; 
      RECT 34.92 161.976 35.016 192.308 ; 
      RECT 34.728 161.976 34.824 192.308 ; 
      RECT 34.536 161.976 34.632 192.308 ; 
      RECT 34.344 161.976 34.44 192.308 ; 
      RECT 33.192 161.976 33.288 192.308 ; 
      RECT 33 161.976 33.096 192.308 ; 
      RECT 32.808 161.976 32.904 192.308 ; 
      RECT 32.424 161.976 32.52 192.308 ; 
      RECT 31.656 161.976 31.752 192.308 ; 
      RECT 31.464 161.976 31.56 192.308 ; 
      RECT 31.272 161.976 31.368 192.308 ; 
      RECT 31.08 161.976 31.176 192.308 ; 
      RECT 30.888 161.976 30.984 192.308 ; 
      RECT 30.696 161.976 30.792 192.308 ; 
      RECT 30.504 158.608 30.6 194.828 ; 
      RECT 30.312 158.46 30.408 194.644 ; 
      RECT 30.12 158.244 30.216 194.428 ; 
      RECT 29.76 178.024 29.856 178.592 ; 
      RECT 29.088 160.94 29.184 176.316 ; 
      RECT 27.6 167.272 27.696 168.224 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 63.568 354.096 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 63.568 354.096 ; 
  END 
END srambank_128x4x74_6t122 
