VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_64x4x18_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_64x4x18_6t122 0 0 ; 
  SIZE 38.448 BY 112.32 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.688 38.036 4.88 ; 
        RECT 0.404 9.008 38.036 9.2 ; 
        RECT 0.404 13.328 38.036 13.52 ; 
        RECT 0.404 17.648 38.036 17.84 ; 
        RECT 0.404 21.968 38.036 22.16 ; 
        RECT 0.404 26.288 38.036 26.48 ; 
        RECT 0.404 30.608 38.036 30.8 ; 
        RECT 0.404 34.928 38.036 35.12 ; 
        RECT 0.404 39.248 38.036 39.44 ; 
        RECT 0.432 41.196 38.016 42.06 ; 
        RECT 22.44 40.076 23.492 40.172 ; 
        RECT 22.964 55.212 23.412 55.308 ; 
        RECT 15.768 53.868 22.68 54.732 ; 
        RECT 15.768 66.54 22.68 67.404 ; 
        RECT 0.404 76.076 38.036 76.268 ; 
        RECT 0.404 80.396 38.036 80.588 ; 
        RECT 0.404 84.716 38.036 84.908 ; 
        RECT 0.404 89.036 38.036 89.228 ; 
        RECT 0.404 93.356 38.036 93.548 ; 
        RECT 0.404 97.676 38.036 97.868 ; 
        RECT 0.404 101.996 38.036 102.188 ; 
        RECT 0.404 106.316 38.036 106.508 ; 
        RECT 0.404 110.636 38.036 110.828 ; 
      LAYER M3 ; 
        RECT 37.908 0.866 37.98 5.506 ; 
        RECT 23.292 0.868 23.364 5.504 ; 
        RECT 17.676 1.012 18.036 5.468 ; 
        RECT 15.084 0.868 15.156 5.504 ; 
        RECT 0.468 0.866 0.54 5.506 ; 
        RECT 37.908 5.186 37.98 9.826 ; 
        RECT 23.292 5.188 23.364 9.824 ; 
        RECT 17.676 5.332 18.036 9.788 ; 
        RECT 15.084 5.188 15.156 9.824 ; 
        RECT 0.468 5.186 0.54 9.826 ; 
        RECT 37.908 9.506 37.98 14.146 ; 
        RECT 23.292 9.508 23.364 14.144 ; 
        RECT 17.676 9.652 18.036 14.108 ; 
        RECT 15.084 9.508 15.156 14.144 ; 
        RECT 0.468 9.506 0.54 14.146 ; 
        RECT 37.908 13.826 37.98 18.466 ; 
        RECT 23.292 13.828 23.364 18.464 ; 
        RECT 17.676 13.972 18.036 18.428 ; 
        RECT 15.084 13.828 15.156 18.464 ; 
        RECT 0.468 13.826 0.54 18.466 ; 
        RECT 37.908 18.146 37.98 22.786 ; 
        RECT 23.292 18.148 23.364 22.784 ; 
        RECT 17.676 18.292 18.036 22.748 ; 
        RECT 15.084 18.148 15.156 22.784 ; 
        RECT 0.468 18.146 0.54 22.786 ; 
        RECT 37.908 22.466 37.98 27.106 ; 
        RECT 23.292 22.468 23.364 27.104 ; 
        RECT 17.676 22.612 18.036 27.068 ; 
        RECT 15.084 22.468 15.156 27.104 ; 
        RECT 0.468 22.466 0.54 27.106 ; 
        RECT 37.908 26.786 37.98 31.426 ; 
        RECT 23.292 26.788 23.364 31.424 ; 
        RECT 17.676 26.932 18.036 31.388 ; 
        RECT 15.084 26.788 15.156 31.424 ; 
        RECT 0.468 26.786 0.54 31.426 ; 
        RECT 37.908 31.106 37.98 35.746 ; 
        RECT 23.292 31.108 23.364 35.744 ; 
        RECT 17.676 31.252 18.036 35.708 ; 
        RECT 15.084 31.108 15.156 35.744 ; 
        RECT 0.468 31.106 0.54 35.746 ; 
        RECT 37.908 35.426 37.98 40.066 ; 
        RECT 23.292 35.428 23.364 40.064 ; 
        RECT 17.676 35.572 18.036 40.028 ; 
        RECT 15.084 35.428 15.156 40.064 ; 
        RECT 0.468 35.426 0.54 40.066 ; 
        RECT 37.908 39.746 37.98 72.574 ; 
        RECT 23.292 40.064 23.364 40.43 ; 
        RECT 23.292 55.024 23.364 72.464 ; 
        RECT 17.82 41.04 18.756 71.372 ; 
        RECT 17.676 71.028 18.036 73.168 ; 
        RECT 17.676 39.92 18.036 42.06 ; 
        RECT 0.468 39.746 0.54 72.574 ; 
        RECT 37.908 72.254 37.98 76.894 ; 
        RECT 23.292 72.256 23.364 76.892 ; 
        RECT 17.676 72.4 18.036 76.856 ; 
        RECT 15.084 72.256 15.156 76.892 ; 
        RECT 0.468 72.254 0.54 76.894 ; 
        RECT 37.908 76.574 37.98 81.214 ; 
        RECT 23.292 76.576 23.364 81.212 ; 
        RECT 17.676 76.72 18.036 81.176 ; 
        RECT 15.084 76.576 15.156 81.212 ; 
        RECT 0.468 76.574 0.54 81.214 ; 
        RECT 37.908 80.894 37.98 85.534 ; 
        RECT 23.292 80.896 23.364 85.532 ; 
        RECT 17.676 81.04 18.036 85.496 ; 
        RECT 15.084 80.896 15.156 85.532 ; 
        RECT 0.468 80.894 0.54 85.534 ; 
        RECT 37.908 85.214 37.98 89.854 ; 
        RECT 23.292 85.216 23.364 89.852 ; 
        RECT 17.676 85.36 18.036 89.816 ; 
        RECT 15.084 85.216 15.156 89.852 ; 
        RECT 0.468 85.214 0.54 89.854 ; 
        RECT 37.908 89.534 37.98 94.174 ; 
        RECT 23.292 89.536 23.364 94.172 ; 
        RECT 17.676 89.68 18.036 94.136 ; 
        RECT 15.084 89.536 15.156 94.172 ; 
        RECT 0.468 89.534 0.54 94.174 ; 
        RECT 37.908 93.854 37.98 98.494 ; 
        RECT 23.292 93.856 23.364 98.492 ; 
        RECT 17.676 94 18.036 98.456 ; 
        RECT 15.084 93.856 15.156 98.492 ; 
        RECT 0.468 93.854 0.54 98.494 ; 
        RECT 37.908 98.174 37.98 102.814 ; 
        RECT 23.292 98.176 23.364 102.812 ; 
        RECT 17.676 98.32 18.036 102.776 ; 
        RECT 15.084 98.176 15.156 102.812 ; 
        RECT 0.468 98.174 0.54 102.814 ; 
        RECT 37.908 102.494 37.98 107.134 ; 
        RECT 23.292 102.496 23.364 107.132 ; 
        RECT 17.676 102.64 18.036 107.096 ; 
        RECT 15.084 102.496 15.156 107.132 ; 
        RECT 0.468 102.494 0.54 107.134 ; 
        RECT 37.908 106.814 37.98 111.454 ; 
        RECT 23.292 106.816 23.364 111.452 ; 
        RECT 17.676 106.96 18.036 111.416 ; 
        RECT 15.084 106.816 15.156 111.452 ; 
        RECT 0.468 106.814 0.54 111.454 ; 
      LAYER V3 ; 
        RECT 0.468 4.688 0.54 4.88 ; 
        RECT 15.084 4.688 15.156 4.88 ; 
        RECT 17.676 4.688 18.036 4.88 ; 
        RECT 23.292 4.688 23.364 4.88 ; 
        RECT 37.908 4.688 37.98 4.88 ; 
        RECT 0.468 9.008 0.54 9.2 ; 
        RECT 15.084 9.008 15.156 9.2 ; 
        RECT 17.676 9.008 18.036 9.2 ; 
        RECT 23.292 9.008 23.364 9.2 ; 
        RECT 37.908 9.008 37.98 9.2 ; 
        RECT 0.468 13.328 0.54 13.52 ; 
        RECT 15.084 13.328 15.156 13.52 ; 
        RECT 17.676 13.328 18.036 13.52 ; 
        RECT 23.292 13.328 23.364 13.52 ; 
        RECT 37.908 13.328 37.98 13.52 ; 
        RECT 0.468 17.648 0.54 17.84 ; 
        RECT 15.084 17.648 15.156 17.84 ; 
        RECT 17.676 17.648 18.036 17.84 ; 
        RECT 23.292 17.648 23.364 17.84 ; 
        RECT 37.908 17.648 37.98 17.84 ; 
        RECT 0.468 21.968 0.54 22.16 ; 
        RECT 15.084 21.968 15.156 22.16 ; 
        RECT 17.676 21.968 18.036 22.16 ; 
        RECT 23.292 21.968 23.364 22.16 ; 
        RECT 37.908 21.968 37.98 22.16 ; 
        RECT 0.468 26.288 0.54 26.48 ; 
        RECT 15.084 26.288 15.156 26.48 ; 
        RECT 17.676 26.288 18.036 26.48 ; 
        RECT 23.292 26.288 23.364 26.48 ; 
        RECT 37.908 26.288 37.98 26.48 ; 
        RECT 0.468 30.608 0.54 30.8 ; 
        RECT 15.084 30.608 15.156 30.8 ; 
        RECT 17.676 30.608 18.036 30.8 ; 
        RECT 23.292 30.608 23.364 30.8 ; 
        RECT 37.908 30.608 37.98 30.8 ; 
        RECT 0.468 34.928 0.54 35.12 ; 
        RECT 15.084 34.928 15.156 35.12 ; 
        RECT 17.676 34.928 18.036 35.12 ; 
        RECT 23.292 34.928 23.364 35.12 ; 
        RECT 37.908 34.928 37.98 35.12 ; 
        RECT 0.468 39.248 0.54 39.44 ; 
        RECT 15.084 39.248 15.156 39.44 ; 
        RECT 17.676 39.248 18.036 39.44 ; 
        RECT 23.292 39.248 23.364 39.44 ; 
        RECT 37.908 39.248 37.98 39.44 ; 
        RECT 0.468 41.196 0.54 42.06 ; 
        RECT 17.836 66.54 17.908 67.404 ; 
        RECT 17.836 53.868 17.908 54.732 ; 
        RECT 17.836 41.196 17.908 42.06 ; 
        RECT 18.044 66.54 18.116 67.404 ; 
        RECT 18.044 53.868 18.116 54.732 ; 
        RECT 18.044 41.196 18.116 42.06 ; 
        RECT 18.252 66.54 18.324 67.404 ; 
        RECT 18.252 53.868 18.324 54.732 ; 
        RECT 18.252 41.196 18.324 42.06 ; 
        RECT 18.46 66.54 18.532 67.404 ; 
        RECT 18.46 53.868 18.532 54.732 ; 
        RECT 18.46 41.196 18.532 42.06 ; 
        RECT 18.668 66.54 18.74 67.404 ; 
        RECT 18.668 53.868 18.74 54.732 ; 
        RECT 18.668 41.196 18.74 42.06 ; 
        RECT 23.292 55.212 23.364 55.308 ; 
        RECT 23.292 40.076 23.364 40.172 ; 
        RECT 0.468 76.076 0.54 76.268 ; 
        RECT 15.084 76.076 15.156 76.268 ; 
        RECT 17.676 76.076 18.036 76.268 ; 
        RECT 23.292 76.076 23.364 76.268 ; 
        RECT 37.908 76.076 37.98 76.268 ; 
        RECT 0.468 80.396 0.54 80.588 ; 
        RECT 15.084 80.396 15.156 80.588 ; 
        RECT 17.676 80.396 18.036 80.588 ; 
        RECT 23.292 80.396 23.364 80.588 ; 
        RECT 37.908 80.396 37.98 80.588 ; 
        RECT 0.468 84.716 0.54 84.908 ; 
        RECT 15.084 84.716 15.156 84.908 ; 
        RECT 17.676 84.716 18.036 84.908 ; 
        RECT 23.292 84.716 23.364 84.908 ; 
        RECT 37.908 84.716 37.98 84.908 ; 
        RECT 0.468 89.036 0.54 89.228 ; 
        RECT 15.084 89.036 15.156 89.228 ; 
        RECT 17.676 89.036 18.036 89.228 ; 
        RECT 23.292 89.036 23.364 89.228 ; 
        RECT 37.908 89.036 37.98 89.228 ; 
        RECT 0.468 93.356 0.54 93.548 ; 
        RECT 15.084 93.356 15.156 93.548 ; 
        RECT 17.676 93.356 18.036 93.548 ; 
        RECT 23.292 93.356 23.364 93.548 ; 
        RECT 37.908 93.356 37.98 93.548 ; 
        RECT 0.468 97.676 0.54 97.868 ; 
        RECT 15.084 97.676 15.156 97.868 ; 
        RECT 17.676 97.676 18.036 97.868 ; 
        RECT 23.292 97.676 23.364 97.868 ; 
        RECT 37.908 97.676 37.98 97.868 ; 
        RECT 0.468 101.996 0.54 102.188 ; 
        RECT 15.084 101.996 15.156 102.188 ; 
        RECT 17.676 101.996 18.036 102.188 ; 
        RECT 23.292 101.996 23.364 102.188 ; 
        RECT 37.908 101.996 37.98 102.188 ; 
        RECT 0.468 106.316 0.54 106.508 ; 
        RECT 15.084 106.316 15.156 106.508 ; 
        RECT 17.676 106.316 18.036 106.508 ; 
        RECT 23.292 106.316 23.364 106.508 ; 
        RECT 37.908 106.316 37.98 106.508 ; 
        RECT 0.468 110.636 0.54 110.828 ; 
        RECT 15.084 110.636 15.156 110.828 ; 
        RECT 17.676 110.636 18.036 110.828 ; 
        RECT 23.292 110.636 23.364 110.828 ; 
        RECT 37.908 110.636 37.98 110.828 ; 
      LAYER M5 ; 
        RECT 23.036 40.004 23.132 55.38 ; 
      LAYER V4 ; 
        RECT 23.036 55.212 23.132 55.308 ; 
        RECT 23.036 40.076 23.132 40.172 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.304 38.016 4.496 ; 
        RECT 0.404 8.624 38.016 8.816 ; 
        RECT 0.404 12.944 38.016 13.136 ; 
        RECT 0.404 17.264 38.016 17.456 ; 
        RECT 0.404 21.584 38.016 21.776 ; 
        RECT 0.404 25.904 38.016 26.096 ; 
        RECT 0.404 30.224 38.016 30.416 ; 
        RECT 0.404 34.544 38.016 34.736 ; 
        RECT 0.404 38.864 38.016 39.056 ; 
        RECT 0.432 42.924 38.016 43.788 ; 
        RECT 15.768 55.596 22.68 56.46 ; 
        RECT 15.768 68.268 22.68 69.132 ; 
        RECT 0.404 75.692 38.016 75.884 ; 
        RECT 0.404 80.012 38.016 80.204 ; 
        RECT 0.404 84.332 38.016 84.524 ; 
        RECT 0.404 88.652 38.016 88.844 ; 
        RECT 0.404 92.972 38.016 93.164 ; 
        RECT 0.404 97.292 38.016 97.484 ; 
        RECT 0.404 101.612 38.016 101.804 ; 
        RECT 0.404 105.932 38.016 106.124 ; 
        RECT 0.404 110.252 38.016 110.444 ; 
      LAYER M3 ; 
        RECT 37.764 0.866 37.836 5.506 ; 
        RECT 23.508 0.866 23.58 5.506 ; 
        RECT 20.448 1.012 20.592 5.468 ; 
        RECT 19.836 1.012 19.944 5.468 ; 
        RECT 14.868 0.866 14.94 5.506 ; 
        RECT 0.612 0.866 0.684 5.506 ; 
        RECT 37.764 5.186 37.836 9.826 ; 
        RECT 23.508 5.186 23.58 9.826 ; 
        RECT 20.448 5.332 20.592 9.788 ; 
        RECT 19.836 5.332 19.944 9.788 ; 
        RECT 14.868 5.186 14.94 9.826 ; 
        RECT 0.612 5.186 0.684 9.826 ; 
        RECT 37.764 9.506 37.836 14.146 ; 
        RECT 23.508 9.506 23.58 14.146 ; 
        RECT 20.448 9.652 20.592 14.108 ; 
        RECT 19.836 9.652 19.944 14.108 ; 
        RECT 14.868 9.506 14.94 14.146 ; 
        RECT 0.612 9.506 0.684 14.146 ; 
        RECT 37.764 13.826 37.836 18.466 ; 
        RECT 23.508 13.826 23.58 18.466 ; 
        RECT 20.448 13.972 20.592 18.428 ; 
        RECT 19.836 13.972 19.944 18.428 ; 
        RECT 14.868 13.826 14.94 18.466 ; 
        RECT 0.612 13.826 0.684 18.466 ; 
        RECT 37.764 18.146 37.836 22.786 ; 
        RECT 23.508 18.146 23.58 22.786 ; 
        RECT 20.448 18.292 20.592 22.748 ; 
        RECT 19.836 18.292 19.944 22.748 ; 
        RECT 14.868 18.146 14.94 22.786 ; 
        RECT 0.612 18.146 0.684 22.786 ; 
        RECT 37.764 22.466 37.836 27.106 ; 
        RECT 23.508 22.466 23.58 27.106 ; 
        RECT 20.448 22.612 20.592 27.068 ; 
        RECT 19.836 22.612 19.944 27.068 ; 
        RECT 14.868 22.466 14.94 27.106 ; 
        RECT 0.612 22.466 0.684 27.106 ; 
        RECT 37.764 26.786 37.836 31.426 ; 
        RECT 23.508 26.786 23.58 31.426 ; 
        RECT 20.448 26.932 20.592 31.388 ; 
        RECT 19.836 26.932 19.944 31.388 ; 
        RECT 14.868 26.786 14.94 31.426 ; 
        RECT 0.612 26.786 0.684 31.426 ; 
        RECT 37.764 31.106 37.836 35.746 ; 
        RECT 23.508 31.106 23.58 35.746 ; 
        RECT 20.448 31.252 20.592 35.708 ; 
        RECT 19.836 31.252 19.944 35.708 ; 
        RECT 14.868 31.106 14.94 35.746 ; 
        RECT 0.612 31.106 0.684 35.746 ; 
        RECT 37.764 35.426 37.836 40.066 ; 
        RECT 23.508 35.426 23.58 40.066 ; 
        RECT 20.448 35.572 20.592 40.028 ; 
        RECT 19.836 35.572 19.944 40.028 ; 
        RECT 14.868 35.426 14.94 40.066 ; 
        RECT 0.612 35.426 0.684 40.066 ; 
        RECT 37.764 39.746 37.836 72.574 ; 
        RECT 23.508 39.746 23.58 72.574 ; 
        RECT 19.692 40.64 20.628 71.372 ; 
        RECT 20.448 39.92 20.592 72.468 ; 
        RECT 19.836 39.92 19.944 72.456 ; 
        RECT 14.868 39.746 14.94 72.574 ; 
        RECT 0.612 39.746 0.684 72.574 ; 
        RECT 37.764 72.254 37.836 76.894 ; 
        RECT 23.508 72.254 23.58 76.894 ; 
        RECT 20.448 72.4 20.592 76.856 ; 
        RECT 19.836 72.4 19.944 76.856 ; 
        RECT 14.868 72.254 14.94 76.894 ; 
        RECT 0.612 72.254 0.684 76.894 ; 
        RECT 37.764 76.574 37.836 81.214 ; 
        RECT 23.508 76.574 23.58 81.214 ; 
        RECT 20.448 76.72 20.592 81.176 ; 
        RECT 19.836 76.72 19.944 81.176 ; 
        RECT 14.868 76.574 14.94 81.214 ; 
        RECT 0.612 76.574 0.684 81.214 ; 
        RECT 37.764 80.894 37.836 85.534 ; 
        RECT 23.508 80.894 23.58 85.534 ; 
        RECT 20.448 81.04 20.592 85.496 ; 
        RECT 19.836 81.04 19.944 85.496 ; 
        RECT 14.868 80.894 14.94 85.534 ; 
        RECT 0.612 80.894 0.684 85.534 ; 
        RECT 37.764 85.214 37.836 89.854 ; 
        RECT 23.508 85.214 23.58 89.854 ; 
        RECT 20.448 85.36 20.592 89.816 ; 
        RECT 19.836 85.36 19.944 89.816 ; 
        RECT 14.868 85.214 14.94 89.854 ; 
        RECT 0.612 85.214 0.684 89.854 ; 
        RECT 37.764 89.534 37.836 94.174 ; 
        RECT 23.508 89.534 23.58 94.174 ; 
        RECT 20.448 89.68 20.592 94.136 ; 
        RECT 19.836 89.68 19.944 94.136 ; 
        RECT 14.868 89.534 14.94 94.174 ; 
        RECT 0.612 89.534 0.684 94.174 ; 
        RECT 37.764 93.854 37.836 98.494 ; 
        RECT 23.508 93.854 23.58 98.494 ; 
        RECT 20.448 94 20.592 98.456 ; 
        RECT 19.836 94 19.944 98.456 ; 
        RECT 14.868 93.854 14.94 98.494 ; 
        RECT 0.612 93.854 0.684 98.494 ; 
        RECT 37.764 98.174 37.836 102.814 ; 
        RECT 23.508 98.174 23.58 102.814 ; 
        RECT 20.448 98.32 20.592 102.776 ; 
        RECT 19.836 98.32 19.944 102.776 ; 
        RECT 14.868 98.174 14.94 102.814 ; 
        RECT 0.612 98.174 0.684 102.814 ; 
        RECT 37.764 102.494 37.836 107.134 ; 
        RECT 23.508 102.494 23.58 107.134 ; 
        RECT 20.448 102.64 20.592 107.096 ; 
        RECT 19.836 102.64 19.944 107.096 ; 
        RECT 14.868 102.494 14.94 107.134 ; 
        RECT 0.612 102.494 0.684 107.134 ; 
        RECT 37.764 106.814 37.836 111.454 ; 
        RECT 23.508 106.814 23.58 111.454 ; 
        RECT 20.448 106.96 20.592 111.416 ; 
        RECT 19.836 106.96 19.944 111.416 ; 
        RECT 14.868 106.814 14.94 111.454 ; 
        RECT 0.612 106.814 0.684 111.454 ; 
      LAYER V3 ; 
        RECT 0.612 4.304 0.684 4.496 ; 
        RECT 14.868 4.304 14.94 4.496 ; 
        RECT 19.836 4.304 19.944 4.496 ; 
        RECT 20.448 4.304 20.592 4.496 ; 
        RECT 23.508 4.304 23.58 4.496 ; 
        RECT 37.764 4.304 37.836 4.496 ; 
        RECT 0.612 8.624 0.684 8.816 ; 
        RECT 14.868 8.624 14.94 8.816 ; 
        RECT 19.836 8.624 19.944 8.816 ; 
        RECT 20.448 8.624 20.592 8.816 ; 
        RECT 23.508 8.624 23.58 8.816 ; 
        RECT 37.764 8.624 37.836 8.816 ; 
        RECT 0.612 12.944 0.684 13.136 ; 
        RECT 14.868 12.944 14.94 13.136 ; 
        RECT 19.836 12.944 19.944 13.136 ; 
        RECT 20.448 12.944 20.592 13.136 ; 
        RECT 23.508 12.944 23.58 13.136 ; 
        RECT 37.764 12.944 37.836 13.136 ; 
        RECT 0.612 17.264 0.684 17.456 ; 
        RECT 14.868 17.264 14.94 17.456 ; 
        RECT 19.836 17.264 19.944 17.456 ; 
        RECT 20.448 17.264 20.592 17.456 ; 
        RECT 23.508 17.264 23.58 17.456 ; 
        RECT 37.764 17.264 37.836 17.456 ; 
        RECT 0.612 21.584 0.684 21.776 ; 
        RECT 14.868 21.584 14.94 21.776 ; 
        RECT 19.836 21.584 19.944 21.776 ; 
        RECT 20.448 21.584 20.592 21.776 ; 
        RECT 23.508 21.584 23.58 21.776 ; 
        RECT 37.764 21.584 37.836 21.776 ; 
        RECT 0.612 25.904 0.684 26.096 ; 
        RECT 14.868 25.904 14.94 26.096 ; 
        RECT 19.836 25.904 19.944 26.096 ; 
        RECT 20.448 25.904 20.592 26.096 ; 
        RECT 23.508 25.904 23.58 26.096 ; 
        RECT 37.764 25.904 37.836 26.096 ; 
        RECT 0.612 30.224 0.684 30.416 ; 
        RECT 14.868 30.224 14.94 30.416 ; 
        RECT 19.836 30.224 19.944 30.416 ; 
        RECT 20.448 30.224 20.592 30.416 ; 
        RECT 23.508 30.224 23.58 30.416 ; 
        RECT 37.764 30.224 37.836 30.416 ; 
        RECT 0.612 34.544 0.684 34.736 ; 
        RECT 14.868 34.544 14.94 34.736 ; 
        RECT 19.836 34.544 19.944 34.736 ; 
        RECT 20.448 34.544 20.592 34.736 ; 
        RECT 23.508 34.544 23.58 34.736 ; 
        RECT 37.764 34.544 37.836 34.736 ; 
        RECT 0.612 38.864 0.684 39.056 ; 
        RECT 14.868 38.864 14.94 39.056 ; 
        RECT 19.836 38.864 19.944 39.056 ; 
        RECT 20.448 38.864 20.592 39.056 ; 
        RECT 23.508 38.864 23.58 39.056 ; 
        RECT 37.764 38.864 37.836 39.056 ; 
        RECT 0.612 42.924 0.684 43.788 ; 
        RECT 19.708 68.268 19.78 69.132 ; 
        RECT 19.708 55.596 19.78 56.46 ; 
        RECT 19.708 42.924 19.78 43.788 ; 
        RECT 19.916 68.268 19.988 69.132 ; 
        RECT 19.916 55.596 19.988 56.46 ; 
        RECT 19.916 42.924 19.988 43.788 ; 
        RECT 20.124 68.268 20.196 69.132 ; 
        RECT 20.124 55.596 20.196 56.46 ; 
        RECT 20.124 42.924 20.196 43.788 ; 
        RECT 20.332 68.268 20.404 69.132 ; 
        RECT 20.332 55.596 20.404 56.46 ; 
        RECT 20.332 42.924 20.404 43.788 ; 
        RECT 20.54 68.268 20.612 69.132 ; 
        RECT 20.54 55.596 20.612 56.46 ; 
        RECT 20.54 42.924 20.612 43.788 ; 
        RECT 0.612 75.692 0.684 75.884 ; 
        RECT 14.868 75.692 14.94 75.884 ; 
        RECT 19.836 75.692 19.944 75.884 ; 
        RECT 20.448 75.692 20.592 75.884 ; 
        RECT 23.508 75.692 23.58 75.884 ; 
        RECT 37.764 75.692 37.836 75.884 ; 
        RECT 0.612 80.012 0.684 80.204 ; 
        RECT 14.868 80.012 14.94 80.204 ; 
        RECT 19.836 80.012 19.944 80.204 ; 
        RECT 20.448 80.012 20.592 80.204 ; 
        RECT 23.508 80.012 23.58 80.204 ; 
        RECT 37.764 80.012 37.836 80.204 ; 
        RECT 0.612 84.332 0.684 84.524 ; 
        RECT 14.868 84.332 14.94 84.524 ; 
        RECT 19.836 84.332 19.944 84.524 ; 
        RECT 20.448 84.332 20.592 84.524 ; 
        RECT 23.508 84.332 23.58 84.524 ; 
        RECT 37.764 84.332 37.836 84.524 ; 
        RECT 0.612 88.652 0.684 88.844 ; 
        RECT 14.868 88.652 14.94 88.844 ; 
        RECT 19.836 88.652 19.944 88.844 ; 
        RECT 20.448 88.652 20.592 88.844 ; 
        RECT 23.508 88.652 23.58 88.844 ; 
        RECT 37.764 88.652 37.836 88.844 ; 
        RECT 0.612 92.972 0.684 93.164 ; 
        RECT 14.868 92.972 14.94 93.164 ; 
        RECT 19.836 92.972 19.944 93.164 ; 
        RECT 20.448 92.972 20.592 93.164 ; 
        RECT 23.508 92.972 23.58 93.164 ; 
        RECT 37.764 92.972 37.836 93.164 ; 
        RECT 0.612 97.292 0.684 97.484 ; 
        RECT 14.868 97.292 14.94 97.484 ; 
        RECT 19.836 97.292 19.944 97.484 ; 
        RECT 20.448 97.292 20.592 97.484 ; 
        RECT 23.508 97.292 23.58 97.484 ; 
        RECT 37.764 97.292 37.836 97.484 ; 
        RECT 0.612 101.612 0.684 101.804 ; 
        RECT 14.868 101.612 14.94 101.804 ; 
        RECT 19.836 101.612 19.944 101.804 ; 
        RECT 20.448 101.612 20.592 101.804 ; 
        RECT 23.508 101.612 23.58 101.804 ; 
        RECT 37.764 101.612 37.836 101.804 ; 
        RECT 0.612 105.932 0.684 106.124 ; 
        RECT 14.868 105.932 14.94 106.124 ; 
        RECT 19.836 105.932 19.944 106.124 ; 
        RECT 20.448 105.932 20.592 106.124 ; 
        RECT 23.508 105.932 23.58 106.124 ; 
        RECT 37.764 105.932 37.836 106.124 ; 
        RECT 0.612 110.252 0.684 110.444 ; 
        RECT 14.868 110.252 14.94 110.444 ; 
        RECT 19.836 110.252 19.944 110.444 ; 
        RECT 20.448 110.252 20.592 110.444 ; 
        RECT 23.508 110.252 23.58 110.444 ; 
        RECT 37.764 110.252 37.836 110.444 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.34 44.812 29.412 44.96 ; 
      LAYER M4 ; 
        RECT 29.132 44.844 29.468 44.94 ; 
      LAYER M5 ; 
        RECT 29.328 41.04 29.424 54 ; 
      LAYER V3 ; 
        RECT 29.34 44.844 29.412 44.94 ; 
      LAYER V4 ; 
        RECT 29.328 44.844 29.424 44.94 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.476 44.824 28.548 44.972 ; 
      LAYER M4 ; 
        RECT 28.268 44.844 28.604 44.94 ; 
      LAYER M5 ; 
        RECT 28.464 41.04 28.56 54 ; 
      LAYER V3 ; 
        RECT 28.476 44.844 28.548 44.94 ; 
      LAYER V4 ; 
        RECT 28.464 44.844 28.56 44.94 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.612 42.508 27.684 42.656 ; 
      LAYER M4 ; 
        RECT 27.404 42.54 27.74 42.636 ; 
      LAYER M5 ; 
        RECT 27.6 41.04 27.696 54 ; 
      LAYER V3 ; 
        RECT 27.612 42.54 27.684 42.636 ; 
      LAYER V4 ; 
        RECT 27.6 42.54 27.696 42.636 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.748 43.468 26.82 44.192 ; 
      LAYER M4 ; 
        RECT 26.54 44.076 26.876 44.172 ; 
      LAYER M5 ; 
        RECT 26.736 41.04 26.832 54 ; 
      LAYER V3 ; 
        RECT 26.748 44.076 26.82 44.172 ; 
      LAYER V4 ; 
        RECT 26.736 44.076 26.832 44.172 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.884 42.52 25.956 42.788 ; 
      LAYER M4 ; 
        RECT 25.676 42.54 26.012 42.636 ; 
      LAYER M5 ; 
        RECT 25.872 41.04 25.968 54 ; 
      LAYER V3 ; 
        RECT 25.884 42.54 25.956 42.636 ; 
      LAYER V4 ; 
        RECT 25.872 42.54 25.968 42.636 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.02 41.452 25.092 42.464 ; 
      LAYER M4 ; 
        RECT 24.812 42.348 25.148 42.444 ; 
      LAYER M5 ; 
        RECT 25.008 41.04 25.104 54 ; 
      LAYER V3 ; 
        RECT 25.02 42.348 25.092 42.444 ; 
      LAYER V4 ; 
        RECT 25.008 42.348 25.104 42.444 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.156 45.592 24.228 45.74 ; 
      LAYER M4 ; 
        RECT 23.948 45.612 24.284 45.708 ; 
      LAYER M5 ; 
        RECT 24.144 41.04 24.24 54 ; 
      LAYER V3 ; 
        RECT 24.156 45.612 24.228 45.708 ; 
      LAYER V4 ; 
        RECT 24.144 45.612 24.24 45.708 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 20.7 42.52 20.772 42.788 ; 
      LAYER M4 ; 
        RECT 19.564 42.54 20.816 42.636 ; 
      LAYER M5 ; 
        RECT 19.608 41.04 19.704 54 ; 
      LAYER V3 ; 
        RECT 20.7 42.54 20.772 42.636 ; 
      LAYER V4 ; 
        RECT 19.608 42.54 19.704 42.636 ; 
    END 
  END ADDRESS[7] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 19.116 41.452 19.188 42.464 ; 
      LAYER M4 ; 
        RECT 18.268 42.348 19.232 42.444 ; 
      LAYER M5 ; 
        RECT 18.312 41.04 18.408 54 ; 
      LAYER V3 ; 
        RECT 19.116 42.348 19.188 42.444 ; 
      LAYER V4 ; 
        RECT 18.312 42.348 18.408 42.444 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.948 42.52 16.02 42.788 ; 
      LAYER M4 ; 
        RECT 15.74 42.54 16.076 42.636 ; 
      LAYER M5 ; 
        RECT 15.936 41.04 16.032 54 ; 
      LAYER V3 ; 
        RECT 15.948 42.54 16.02 42.636 ; 
      LAYER V4 ; 
        RECT 15.936 42.54 16.032 42.636 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.084 45.976 15.156 46.172 ; 
      LAYER M4 ; 
        RECT 14.876 45.996 15.212 46.092 ; 
      LAYER M5 ; 
        RECT 15.072 41.04 15.168 54 ; 
      LAYER V3 ; 
        RECT 15.084 45.996 15.156 46.092 ; 
      LAYER V4 ; 
        RECT 15.072 45.996 15.168 46.092 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.228 41.452 15.3 42.464 ; 
      LAYER M4 ; 
        RECT 14.164 42.348 15.344 42.444 ; 
      LAYER M5 ; 
        RECT 14.208 41.04 14.304 54 ; 
      LAYER V3 ; 
        RECT 15.228 42.348 15.3 42.444 ; 
      LAYER V4 ; 
        RECT 14.208 42.348 14.304 42.444 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 13.356 44.812 13.428 44.96 ; 
      LAYER M4 ; 
        RECT 13.148 44.844 13.484 44.94 ; 
      LAYER M5 ; 
        RECT 13.344 41.04 13.44 54 ; 
      LAYER V3 ; 
        RECT 13.356 44.844 13.428 44.94 ; 
      LAYER V4 ; 
        RECT 13.344 44.844 13.44 44.94 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 12.492 42.52 12.564 43.436 ; 
      LAYER M4 ; 
        RECT 12.284 42.54 12.62 42.636 ; 
      LAYER M5 ; 
        RECT 12.48 41.04 12.576 54 ; 
      LAYER V3 ; 
        RECT 12.492 42.54 12.564 42.636 ; 
      LAYER V4 ; 
        RECT 12.48 42.54 12.576 42.636 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 11.628 41.452 11.7 42.464 ; 
      LAYER M4 ; 
        RECT 11.42 42.348 11.756 42.444 ; 
      LAYER M5 ; 
        RECT 11.616 41.04 11.712 54 ; 
      LAYER V3 ; 
        RECT 11.628 42.348 11.7 42.444 ; 
      LAYER V4 ; 
        RECT 11.616 42.348 11.712 42.444 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 10.764 42.508 10.836 42.656 ; 
      LAYER M4 ; 
        RECT 10.556 42.54 10.892 42.636 ; 
      LAYER M5 ; 
        RECT 10.752 41.04 10.848 54 ; 
      LAYER V3 ; 
        RECT 10.764 42.54 10.836 42.636 ; 
      LAYER V4 ; 
        RECT 10.752 42.54 10.848 42.636 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 9.9 44.812 9.972 44.96 ; 
      LAYER M4 ; 
        RECT 9.692 44.844 10.028 44.94 ; 
      LAYER M5 ; 
        RECT 9.888 41.04 9.984 54 ; 
      LAYER V3 ; 
        RECT 9.9 44.844 9.972 44.94 ; 
      LAYER V4 ; 
        RECT 9.888 44.844 9.984 44.94 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.712 20.544 1.808 ; 
      LAYER M3 ; 
        RECT 20.304 1.51 20.376 2.468 ; 
      LAYER V3 ; 
        RECT 20.304 1.712 20.376 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.328 20.816 1.424 ; 
      LAYER M3 ; 
        RECT 19.404 1.08 19.476 2.7 ; 
      LAYER V3 ; 
        RECT 19.404 1.328 19.476 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 6.032 20.544 6.128 ; 
      LAYER M3 ; 
        RECT 20.304 5.83 20.376 6.788 ; 
      LAYER V3 ; 
        RECT 20.304 6.032 20.376 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 5.648 20.816 5.744 ; 
      LAYER M3 ; 
        RECT 19.404 5.4 19.476 7.02 ; 
      LAYER V3 ; 
        RECT 19.404 5.648 19.476 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 10.352 20.544 10.448 ; 
      LAYER M3 ; 
        RECT 20.304 10.15 20.376 11.108 ; 
      LAYER V3 ; 
        RECT 20.304 10.352 20.376 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 9.968 20.816 10.064 ; 
      LAYER M3 ; 
        RECT 19.404 9.72 19.476 11.34 ; 
      LAYER V3 ; 
        RECT 19.404 9.968 19.476 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.672 20.544 14.768 ; 
      LAYER M3 ; 
        RECT 20.304 14.47 20.376 15.428 ; 
      LAYER V3 ; 
        RECT 20.304 14.672 20.376 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.288 20.816 14.384 ; 
      LAYER M3 ; 
        RECT 19.404 14.04 19.476 15.66 ; 
      LAYER V3 ; 
        RECT 19.404 14.288 19.476 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.992 20.544 19.088 ; 
      LAYER M3 ; 
        RECT 20.304 18.79 20.376 19.748 ; 
      LAYER V3 ; 
        RECT 20.304 18.992 20.376 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.608 20.816 18.704 ; 
      LAYER M3 ; 
        RECT 19.404 18.36 19.476 19.98 ; 
      LAYER V3 ; 
        RECT 19.404 18.608 19.476 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 23.312 20.544 23.408 ; 
      LAYER M3 ; 
        RECT 20.304 23.11 20.376 24.068 ; 
      LAYER V3 ; 
        RECT 20.304 23.312 20.376 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 22.928 20.816 23.024 ; 
      LAYER M3 ; 
        RECT 19.404 22.68 19.476 24.3 ; 
      LAYER V3 ; 
        RECT 19.404 22.928 19.476 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.632 20.544 27.728 ; 
      LAYER M3 ; 
        RECT 20.304 27.43 20.376 28.388 ; 
      LAYER V3 ; 
        RECT 20.304 27.632 20.376 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.248 20.816 27.344 ; 
      LAYER M3 ; 
        RECT 19.404 27 19.476 28.62 ; 
      LAYER V3 ; 
        RECT 19.404 27.248 19.476 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.952 20.544 32.048 ; 
      LAYER M3 ; 
        RECT 20.304 31.75 20.376 32.708 ; 
      LAYER V3 ; 
        RECT 20.304 31.952 20.376 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.568 20.816 31.664 ; 
      LAYER M3 ; 
        RECT 19.404 31.32 19.476 32.94 ; 
      LAYER V3 ; 
        RECT 19.404 31.568 19.476 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 36.272 20.544 36.368 ; 
      LAYER M3 ; 
        RECT 20.304 36.07 20.376 37.028 ; 
      LAYER V3 ; 
        RECT 20.304 36.272 20.376 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 35.888 20.816 35.984 ; 
      LAYER M3 ; 
        RECT 19.404 35.64 19.476 37.26 ; 
      LAYER V3 ; 
        RECT 19.404 35.888 19.476 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 73.1 20.544 73.196 ; 
      LAYER M3 ; 
        RECT 20.304 72.898 20.376 73.856 ; 
      LAYER V3 ; 
        RECT 20.304 73.1 20.376 73.196 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 72.716 20.816 72.812 ; 
      LAYER M3 ; 
        RECT 19.404 72.468 19.476 74.088 ; 
      LAYER V3 ; 
        RECT 19.404 72.716 19.476 72.812 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 77.42 20.544 77.516 ; 
      LAYER M3 ; 
        RECT 20.304 77.218 20.376 78.176 ; 
      LAYER V3 ; 
        RECT 20.304 77.42 20.376 77.516 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 77.036 20.816 77.132 ; 
      LAYER M3 ; 
        RECT 19.404 76.788 19.476 78.408 ; 
      LAYER V3 ; 
        RECT 19.404 77.036 19.476 77.132 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 81.74 20.544 81.836 ; 
      LAYER M3 ; 
        RECT 20.304 81.538 20.376 82.496 ; 
      LAYER V3 ; 
        RECT 20.304 81.74 20.376 81.836 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 81.356 20.816 81.452 ; 
      LAYER M3 ; 
        RECT 19.404 81.108 19.476 82.728 ; 
      LAYER V3 ; 
        RECT 19.404 81.356 19.476 81.452 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 86.06 20.544 86.156 ; 
      LAYER M3 ; 
        RECT 20.304 85.858 20.376 86.816 ; 
      LAYER V3 ; 
        RECT 20.304 86.06 20.376 86.156 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 85.676 20.816 85.772 ; 
      LAYER M3 ; 
        RECT 19.404 85.428 19.476 87.048 ; 
      LAYER V3 ; 
        RECT 19.404 85.676 19.476 85.772 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 90.38 20.544 90.476 ; 
      LAYER M3 ; 
        RECT 20.304 90.178 20.376 91.136 ; 
      LAYER V3 ; 
        RECT 20.304 90.38 20.376 90.476 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 89.996 20.816 90.092 ; 
      LAYER M3 ; 
        RECT 19.404 89.748 19.476 91.368 ; 
      LAYER V3 ; 
        RECT 19.404 89.996 19.476 90.092 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 94.7 20.544 94.796 ; 
      LAYER M3 ; 
        RECT 20.304 94.498 20.376 95.456 ; 
      LAYER V3 ; 
        RECT 20.304 94.7 20.376 94.796 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 94.316 20.816 94.412 ; 
      LAYER M3 ; 
        RECT 19.404 94.068 19.476 95.688 ; 
      LAYER V3 ; 
        RECT 19.404 94.316 19.476 94.412 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 99.02 20.544 99.116 ; 
      LAYER M3 ; 
        RECT 20.304 98.818 20.376 99.776 ; 
      LAYER V3 ; 
        RECT 20.304 99.02 20.376 99.116 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 98.636 20.816 98.732 ; 
      LAYER M3 ; 
        RECT 19.404 98.388 19.476 100.008 ; 
      LAYER V3 ; 
        RECT 19.404 98.636 19.476 98.732 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 103.34 20.544 103.436 ; 
      LAYER M3 ; 
        RECT 20.304 103.138 20.376 104.096 ; 
      LAYER V3 ; 
        RECT 20.304 103.34 20.376 103.436 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 102.956 20.816 103.052 ; 
      LAYER M3 ; 
        RECT 19.404 102.708 19.476 104.328 ; 
      LAYER V3 ; 
        RECT 19.404 102.956 19.476 103.052 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 107.66 20.544 107.756 ; 
      LAYER M3 ; 
        RECT 20.304 107.458 20.376 108.416 ; 
      LAYER V3 ; 
        RECT 20.304 107.66 20.376 107.756 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 107.276 20.816 107.372 ; 
      LAYER M3 ; 
        RECT 19.404 107.028 19.476 108.648 ; 
      LAYER V3 ; 
        RECT 19.404 107.276 19.476 107.372 ; 
    END 
  END wd[17] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.852 38.448 74.466 ; 
        RECT 0 72.414 38.448 76.788 ; 
        RECT 0 76.734 38.448 81.108 ; 
        RECT 0 81.054 38.448 85.428 ; 
        RECT 0 85.374 38.448 89.748 ; 
        RECT 0 89.694 38.448 94.068 ; 
        RECT 0 94.014 38.448 98.388 ; 
        RECT 0 98.334 38.448 102.708 ; 
        RECT 0 102.654 38.448 107.028 ; 
        RECT 0 106.974 38.448 111.348 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.852 38.448 74.466 ; 
        RECT 0 72.414 38.448 76.788 ; 
        RECT 0 76.734 38.448 81.108 ; 
        RECT 0 81.054 38.448 85.428 ; 
        RECT 0 85.374 38.448 89.748 ; 
        RECT 0 89.694 38.448 94.068 ; 
        RECT 0 94.014 38.448 98.388 ; 
        RECT 0 98.334 38.448 102.708 ; 
        RECT 0 102.654 38.448 107.028 ; 
        RECT 0 106.974 38.448 111.348 ; 
  LAYER V1 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.852 38.448 74.466 ; 
        RECT 0 72.414 38.448 76.788 ; 
        RECT 0 76.734 38.448 81.108 ; 
        RECT 0 81.054 38.448 85.428 ; 
        RECT 0 85.374 38.448 89.748 ; 
        RECT 0 89.694 38.448 94.068 ; 
        RECT 0 94.014 38.448 98.388 ; 
        RECT 0 98.334 38.448 102.708 ; 
        RECT 0 102.654 38.448 107.028 ; 
        RECT 0 106.974 38.448 111.348 ; 
  LAYER V2 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.852 38.448 74.466 ; 
        RECT 0 72.414 38.448 76.788 ; 
        RECT 0 76.734 38.448 81.108 ; 
        RECT 0 81.054 38.448 85.428 ; 
        RECT 0 85.374 38.448 89.748 ; 
        RECT 0 89.694 38.448 94.068 ; 
        RECT 0 94.014 38.448 98.388 ; 
        RECT 0 98.334 38.448 102.708 ; 
        RECT 0 102.654 38.448 107.028 ; 
        RECT 0 106.974 38.448 111.348 ; 
  LAYER M3 ; 
      RECT 20.952 1.38 21.024 5.122 ; 
      RECT 20.808 1.38 20.88 5.122 ; 
      RECT 20.664 3.688 20.736 4.978 ; 
      RECT 20.196 4.476 20.268 4.914 ; 
      RECT 20.16 1.51 20.232 2.468 ; 
      RECT 20.016 3.834 20.088 4.448 ; 
      RECT 19.692 3.936 19.764 4.968 ; 
      RECT 17.532 1.38 17.604 5.122 ; 
      RECT 17.388 1.38 17.46 5.122 ; 
      RECT 17.244 2.104 17.316 4.376 ; 
      RECT 20.952 5.7 21.024 9.442 ; 
      RECT 20.808 5.7 20.88 9.442 ; 
      RECT 20.664 8.008 20.736 9.298 ; 
      RECT 20.196 8.796 20.268 9.234 ; 
      RECT 20.16 5.83 20.232 6.788 ; 
      RECT 20.016 8.154 20.088 8.768 ; 
      RECT 19.692 8.256 19.764 9.288 ; 
      RECT 17.532 5.7 17.604 9.442 ; 
      RECT 17.388 5.7 17.46 9.442 ; 
      RECT 17.244 6.424 17.316 8.696 ; 
      RECT 20.952 10.02 21.024 13.762 ; 
      RECT 20.808 10.02 20.88 13.762 ; 
      RECT 20.664 12.328 20.736 13.618 ; 
      RECT 20.196 13.116 20.268 13.554 ; 
      RECT 20.16 10.15 20.232 11.108 ; 
      RECT 20.016 12.474 20.088 13.088 ; 
      RECT 19.692 12.576 19.764 13.608 ; 
      RECT 17.532 10.02 17.604 13.762 ; 
      RECT 17.388 10.02 17.46 13.762 ; 
      RECT 17.244 10.744 17.316 13.016 ; 
      RECT 20.952 14.34 21.024 18.082 ; 
      RECT 20.808 14.34 20.88 18.082 ; 
      RECT 20.664 16.648 20.736 17.938 ; 
      RECT 20.196 17.436 20.268 17.874 ; 
      RECT 20.16 14.47 20.232 15.428 ; 
      RECT 20.016 16.794 20.088 17.408 ; 
      RECT 19.692 16.896 19.764 17.928 ; 
      RECT 17.532 14.34 17.604 18.082 ; 
      RECT 17.388 14.34 17.46 18.082 ; 
      RECT 17.244 15.064 17.316 17.336 ; 
      RECT 20.952 18.66 21.024 22.402 ; 
      RECT 20.808 18.66 20.88 22.402 ; 
      RECT 20.664 20.968 20.736 22.258 ; 
      RECT 20.196 21.756 20.268 22.194 ; 
      RECT 20.16 18.79 20.232 19.748 ; 
      RECT 20.016 21.114 20.088 21.728 ; 
      RECT 19.692 21.216 19.764 22.248 ; 
      RECT 17.532 18.66 17.604 22.402 ; 
      RECT 17.388 18.66 17.46 22.402 ; 
      RECT 17.244 19.384 17.316 21.656 ; 
      RECT 20.952 22.98 21.024 26.722 ; 
      RECT 20.808 22.98 20.88 26.722 ; 
      RECT 20.664 25.288 20.736 26.578 ; 
      RECT 20.196 26.076 20.268 26.514 ; 
      RECT 20.16 23.11 20.232 24.068 ; 
      RECT 20.016 25.434 20.088 26.048 ; 
      RECT 19.692 25.536 19.764 26.568 ; 
      RECT 17.532 22.98 17.604 26.722 ; 
      RECT 17.388 22.98 17.46 26.722 ; 
      RECT 17.244 23.704 17.316 25.976 ; 
      RECT 20.952 27.3 21.024 31.042 ; 
      RECT 20.808 27.3 20.88 31.042 ; 
      RECT 20.664 29.608 20.736 30.898 ; 
      RECT 20.196 30.396 20.268 30.834 ; 
      RECT 20.16 27.43 20.232 28.388 ; 
      RECT 20.016 29.754 20.088 30.368 ; 
      RECT 19.692 29.856 19.764 30.888 ; 
      RECT 17.532 27.3 17.604 31.042 ; 
      RECT 17.388 27.3 17.46 31.042 ; 
      RECT 17.244 28.024 17.316 30.296 ; 
      RECT 20.952 31.62 21.024 35.362 ; 
      RECT 20.808 31.62 20.88 35.362 ; 
      RECT 20.664 33.928 20.736 35.218 ; 
      RECT 20.196 34.716 20.268 35.154 ; 
      RECT 20.16 31.75 20.232 32.708 ; 
      RECT 20.016 34.074 20.088 34.688 ; 
      RECT 19.692 34.176 19.764 35.208 ; 
      RECT 17.532 31.62 17.604 35.362 ; 
      RECT 17.388 31.62 17.46 35.362 ; 
      RECT 17.244 32.344 17.316 34.616 ; 
      RECT 20.952 35.94 21.024 39.682 ; 
      RECT 20.808 35.94 20.88 39.682 ; 
      RECT 20.664 38.248 20.736 39.538 ; 
      RECT 20.196 39.036 20.268 39.474 ; 
      RECT 20.16 36.07 20.232 37.028 ; 
      RECT 20.016 38.394 20.088 39.008 ; 
      RECT 19.692 38.496 19.764 39.528 ; 
      RECT 17.532 35.94 17.604 39.682 ; 
      RECT 17.388 35.94 17.46 39.682 ; 
      RECT 17.244 36.664 17.316 38.936 ; 
      RECT 37.62 55.024 37.692 72.446 ; 
      RECT 37.476 49.764 37.548 50.04 ; 
      RECT 37.476 56.996 37.548 58.854 ; 
      RECT 37.332 39.746 37.404 72.574 ; 
      RECT 37.188 54.824 37.26 57.914 ; 
      RECT 37.188 58.1188 37.26 60.084 ; 
      RECT 37.188 60.284 37.26 61.77 ; 
      RECT 37.188 62.022 37.26 65.268 ; 
      RECT 37.044 55.166 37.116 57.734 ; 
      RECT 37.044 60.444 37.116 62.572 ; 
      RECT 36.9 39.746 36.972 41.146 ; 
      RECT 36.468 39.746 36.54 41.146 ; 
      RECT 36.036 39.746 36.108 41.146 ; 
      RECT 35.604 39.746 35.676 41.146 ; 
      RECT 35.172 39.746 35.244 41.146 ; 
      RECT 34.74 39.746 34.812 41.146 ; 
      RECT 34.308 39.746 34.38 41.146 ; 
      RECT 33.876 39.746 33.948 41.146 ; 
      RECT 33.444 39.746 33.516 41.146 ; 
      RECT 33.012 39.746 33.084 41.146 ; 
      RECT 32.58 39.746 32.652 41.146 ; 
      RECT 32.148 39.746 32.22 41.146 ; 
      RECT 31.716 39.746 31.788 41.146 ; 
      RECT 31.284 39.746 31.356 41.146 ; 
      RECT 30.852 39.746 30.924 41.146 ; 
      RECT 30.42 39.746 30.492 41.146 ; 
      RECT 29.988 39.746 30.06 41.146 ; 
      RECT 29.556 39.746 29.628 41.146 ; 
      RECT 29.124 39.746 29.196 41.146 ; 
      RECT 28.692 39.746 28.764 41.146 ; 
      RECT 28.26 39.746 28.332 41.146 ; 
      RECT 27.828 39.746 27.9 41.146 ; 
      RECT 27.396 39.746 27.468 41.146 ; 
      RECT 26.964 39.746 27.036 41.146 ; 
      RECT 26.532 39.746 26.604 41.146 ; 
      RECT 26.1 39.746 26.172 41.146 ; 
      RECT 25.668 39.746 25.74 41.146 ; 
      RECT 25.236 39.746 25.308 41.146 ; 
      RECT 24.804 39.746 24.876 41.146 ; 
      RECT 24.372 39.746 24.444 41.146 ; 
      RECT 24.228 54.9 24.3 57.7188 ; 
      RECT 24.228 60.688 24.3 65.412 ; 
      RECT 24.156 42.388 24.228 45.092 ; 
      RECT 24.156 48.076 24.228 49.268 ; 
      RECT 24.084 55.154 24.156 57.914 ; 
      RECT 24.084 58.118 24.156 62.084 ; 
      RECT 24.084 62.204 24.156 65.34 ; 
      RECT 23.94 39.746 24.012 72.574 ; 
      RECT 23.796 56.244 23.868 56.576 ; 
      RECT 23.724 42.82 23.796 45.344 ; 
      RECT 23.724 46.996 23.796 47.756 ; 
      RECT 23.724 50.524 23.796 50.72 ; 
      RECT 23.652 55.024 23.724 72.464 ; 
      RECT 23.292 41.308 23.364 44.516 ; 
      RECT 23.292 46.708 23.364 48.98 ; 
      RECT 23.148 46.996 23.22 48.476 ; 
      RECT 23.004 44.404 23.076 44.948 ; 
      RECT 23.004 48.364 23.076 49.268 ; 
      RECT 23.004 53.332 23.076 53.588 ; 
      RECT 22.86 44.812 22.932 44.96 ; 
      RECT 22.86 51.316 22.932 51.488 ; 
      RECT 22.86 53.452 22.932 53.6 ; 
      RECT 22.716 46.06 22.788 48.044 ; 
      RECT 22.716 48.22 22.788 48.98 ; 
      RECT 22.716 52.06 22.788 53.3 ; 
      RECT 22.572 61.18 22.644 64.1 ; 
      RECT 22.572 65.5 22.644 68.42 ; 
      RECT 21.276 44.548 21.348 45.74 ; 
      RECT 21.276 49.3 21.348 49.556 ; 
      RECT 21.276 50.38 21.348 52.22 ; 
      RECT 21.276 55.18 21.348 55.328 ; 
      RECT 21.276 63.34 21.348 64.532 ; 
      RECT 21.132 44.836 21.204 46.856 ; 
      RECT 21.132 47.932 21.204 51.14 ; 
      RECT 21.132 55.312 21.204 56.396 ; 
      RECT 21.132 56.716 21.204 57.62 ; 
      RECT 20.988 44.548 21.06 47.252 ; 
      RECT 20.988 47.644 21.06 48.98 ; 
      RECT 20.988 49.804 21.06 50.348 ; 
      RECT 20.988 52.54 21.06 55.748 ; 
      RECT 20.988 57.484 21.06 57.632 ; 
      RECT 20.988 66.148 21.06 67.484 ; 
      RECT 20.844 45.484 20.916 46.028 ; 
      RECT 20.844 53.044 20.916 56.972 ; 
      RECT 20.844 58.732 20.916 59.924 ; 
      RECT 20.844 65.5 20.916 66.548 ; 
      RECT 20.7 41.74 20.772 42.356 ; 
      RECT 20.7 44.98 20.772 52.124 ; 
      RECT 20.7 56.284 20.772 65.612 ; 
      RECT 20.7 66.436 20.772 70.868 ; 
      RECT 19.548 42.82 19.62 43.868 ; 
      RECT 19.548 44.404 19.62 44.66 ; 
      RECT 19.548 44.98 19.62 45.884 ; 
      RECT 19.548 46.06 19.62 46.82 ; 
      RECT 19.548 47.14 19.62 57.62 ; 
      RECT 19.548 57.796 19.62 63.02 ; 
      RECT 19.548 67.372 19.62 68.42 ; 
      RECT 19.404 46.816 19.476 47.9 ; 
      RECT 19.404 48.22 19.476 51.572 ; 
      RECT 19.404 52.252 19.476 55.604 ; 
      RECT 19.404 55.78 19.476 60.86 ; 
      RECT 19.404 61.684 19.476 62.372 ; 
      RECT 19.404 65.212 19.476 69.5 ; 
      RECT 19.26 47.14 19.332 48.224 ; 
      RECT 19.26 48.844 19.332 48.992 ; 
      RECT 19.26 51.964 19.332 55.892 ; 
      RECT 19.26 56.86 19.332 58.7 ; 
      RECT 19.26 60.1 19.332 63.056 ; 
      RECT 19.116 43.612 19.188 47.9 ; 
      RECT 19.116 54.268 19.188 55.136 ; 
      RECT 19.116 59.812 19.188 61.004 ; 
      RECT 18.972 46.204 19.044 48.044 ; 
      RECT 18.972 52.54 19.044 53.3 ; 
      RECT 18.972 53.464 19.044 53.612 ; 
      RECT 18.972 54.556 19.044 55.892 ; 
      RECT 18.972 56.428 19.044 61.796 ; 
      RECT 18.972 62.224 19.044 66.692 ; 
      RECT 18.828 43.9 18.9 44.66 ; 
      RECT 18.828 45.484 18.9 46.028 ; 
      RECT 18.828 47.14 18.9 59.78 ; 
      RECT 18.828 60.1 18.9 61.94 ; 
      RECT 18.828 64.42 18.9 66.26 ; 
      RECT 18.828 69.676 18.9 70.58 ; 
      RECT 18.684 39.852 18.756 40.468 ; 
      RECT 18.684 71.896 18.756 72.512 ; 
      RECT 18.54 39.852 18.612 40.052 ; 
      RECT 18.252 39.852 18.324 40.138 ; 
      RECT 18.252 72.174 18.324 72.574 ; 
      RECT 17.676 45.916 17.748 46.676 ; 
      RECT 17.676 48.868 17.748 50.348 ; 
      RECT 17.676 56.716 17.748 57.62 ; 
      RECT 17.676 58.876 17.748 63.452 ; 
      RECT 17.676 66.58 17.748 68.42 ; 
      RECT 17.676 70.732 17.748 70.88 ; 
      RECT 17.532 41.74 17.604 43.724 ; 
      RECT 17.532 58.06 17.604 58.208 ; 
      RECT 17.532 62.368 17.604 65.612 ; 
      RECT 17.388 43.612 17.46 44.66 ; 
      RECT 17.388 45.772 17.46 47.108 ; 
      RECT 17.388 47.932 17.46 48.332 ; 
      RECT 17.388 51.46 17.46 62.516 ; 
      RECT 17.388 63.052 17.46 63.956 ; 
      RECT 17.244 42.244 17.316 46.82 ; 
      RECT 17.244 61.18 17.316 61.94 ; 
      RECT 17.244 64.396 17.316 64.544 ; 
      RECT 17.244 65.5 17.316 68.708 ; 
      RECT 17.1 46.06 17.172 50.06 ; 
      RECT 17.1 63.82 17.172 63.968 ; 
      RECT 16.956 42.82 17.028 42.932 ; 
      RECT 15.66 44.404 15.732 46.028 ; 
      RECT 15.372 44.548 15.444 46.964 ; 
      RECT 15.228 43.9 15.3 44.156 ; 
      RECT 15.084 40.064 15.156 40.268 ; 
      RECT 15.084 52.54 15.156 53.3 ; 
      RECT 15.084 55.024 15.156 72.464 ; 
      RECT 14.724 55.024 14.796 72.464 ; 
      RECT 14.652 41.74 14.724 42.5 ; 
      RECT 14.652 44.836 14.724 53.876 ; 
      RECT 14.58 56.244 14.652 56.576 ; 
      RECT 14.436 39.746 14.508 72.574 ; 
      RECT 14.292 55.154 14.364 57.914 ; 
      RECT 14.292 58.118 14.364 62.084 ; 
      RECT 14.292 62.204 14.364 65.34 ; 
      RECT 14.22 41.74 14.292 43.724 ; 
      RECT 14.22 46.852 14.292 49.124 ; 
      RECT 14.22 50.38 14.292 53.3 ; 
      RECT 14.148 54.9 14.22 57.7188 ; 
      RECT 14.148 60.688 14.22 65.412 ; 
      RECT 14.004 39.746 14.076 41.146 ; 
      RECT 13.572 39.746 13.644 41.146 ; 
      RECT 13.14 39.746 13.212 41.146 ; 
      RECT 12.708 39.746 12.78 41.146 ; 
      RECT 12.276 39.746 12.348 41.146 ; 
      RECT 11.844 39.746 11.916 41.146 ; 
      RECT 11.412 39.746 11.484 41.146 ; 
      RECT 10.98 39.746 11.052 41.146 ; 
      RECT 10.548 39.746 10.62 41.146 ; 
      RECT 10.116 39.746 10.188 41.146 ; 
      RECT 9.684 39.746 9.756 41.146 ; 
      RECT 9.252 39.746 9.324 41.146 ; 
      RECT 8.82 39.746 8.892 41.146 ; 
      RECT 8.388 39.746 8.46 41.146 ; 
      RECT 7.956 39.746 8.028 41.146 ; 
      RECT 7.524 39.746 7.596 41.146 ; 
      RECT 7.092 39.746 7.164 41.146 ; 
      RECT 6.66 39.746 6.732 41.146 ; 
      RECT 6.228 39.746 6.3 41.146 ; 
      RECT 5.796 39.746 5.868 41.146 ; 
      RECT 5.364 39.746 5.436 41.146 ; 
      RECT 4.932 39.746 5.004 41.146 ; 
      RECT 4.5 39.746 4.572 41.146 ; 
      RECT 4.068 39.746 4.14 41.146 ; 
      RECT 3.636 39.746 3.708 41.146 ; 
      RECT 3.204 39.746 3.276 41.146 ; 
      RECT 2.772 39.746 2.844 41.146 ; 
      RECT 2.34 39.746 2.412 41.146 ; 
      RECT 1.908 39.746 1.98 41.146 ; 
      RECT 1.476 39.746 1.548 41.146 ; 
      RECT 1.332 55.166 1.404 57.734 ; 
      RECT 1.332 60.444 1.404 62.572 ; 
      RECT 1.26 43.9 1.332 44.804 ; 
      RECT 1.188 54.824 1.26 57.914 ; 
      RECT 1.188 58.1188 1.26 60.084 ; 
      RECT 1.188 60.284 1.26 61.77 ; 
      RECT 1.188 62.022 1.26 65.268 ; 
      RECT 1.044 39.746 1.116 72.574 ; 
      RECT 0.9 49.764 0.972 50.04 ; 
      RECT 0.9 56.996 0.972 58.854 ; 
      RECT 0.756 55.024 0.828 72.446 ; 
        RECT 20.952 72.768 21.024 76.51 ; 
        RECT 20.808 72.768 20.88 76.51 ; 
        RECT 20.664 75.076 20.736 76.366 ; 
        RECT 20.196 75.864 20.268 76.302 ; 
        RECT 20.16 72.898 20.232 73.856 ; 
        RECT 20.016 75.222 20.088 75.836 ; 
        RECT 19.692 75.324 19.764 76.356 ; 
        RECT 17.532 72.768 17.604 76.51 ; 
        RECT 17.388 72.768 17.46 76.51 ; 
        RECT 17.244 73.492 17.316 75.764 ; 
        RECT 20.952 77.088 21.024 80.83 ; 
        RECT 20.808 77.088 20.88 80.83 ; 
        RECT 20.664 79.396 20.736 80.686 ; 
        RECT 20.196 80.184 20.268 80.622 ; 
        RECT 20.16 77.218 20.232 78.176 ; 
        RECT 20.016 79.542 20.088 80.156 ; 
        RECT 19.692 79.644 19.764 80.676 ; 
        RECT 17.532 77.088 17.604 80.83 ; 
        RECT 17.388 77.088 17.46 80.83 ; 
        RECT 17.244 77.812 17.316 80.084 ; 
        RECT 20.952 81.408 21.024 85.15 ; 
        RECT 20.808 81.408 20.88 85.15 ; 
        RECT 20.664 83.716 20.736 85.006 ; 
        RECT 20.196 84.504 20.268 84.942 ; 
        RECT 20.16 81.538 20.232 82.496 ; 
        RECT 20.016 83.862 20.088 84.476 ; 
        RECT 19.692 83.964 19.764 84.996 ; 
        RECT 17.532 81.408 17.604 85.15 ; 
        RECT 17.388 81.408 17.46 85.15 ; 
        RECT 17.244 82.132 17.316 84.404 ; 
        RECT 20.952 85.728 21.024 89.47 ; 
        RECT 20.808 85.728 20.88 89.47 ; 
        RECT 20.664 88.036 20.736 89.326 ; 
        RECT 20.196 88.824 20.268 89.262 ; 
        RECT 20.16 85.858 20.232 86.816 ; 
        RECT 20.016 88.182 20.088 88.796 ; 
        RECT 19.692 88.284 19.764 89.316 ; 
        RECT 17.532 85.728 17.604 89.47 ; 
        RECT 17.388 85.728 17.46 89.47 ; 
        RECT 17.244 86.452 17.316 88.724 ; 
        RECT 20.952 90.048 21.024 93.79 ; 
        RECT 20.808 90.048 20.88 93.79 ; 
        RECT 20.664 92.356 20.736 93.646 ; 
        RECT 20.196 93.144 20.268 93.582 ; 
        RECT 20.16 90.178 20.232 91.136 ; 
        RECT 20.016 92.502 20.088 93.116 ; 
        RECT 19.692 92.604 19.764 93.636 ; 
        RECT 17.532 90.048 17.604 93.79 ; 
        RECT 17.388 90.048 17.46 93.79 ; 
        RECT 17.244 90.772 17.316 93.044 ; 
        RECT 20.952 94.368 21.024 98.11 ; 
        RECT 20.808 94.368 20.88 98.11 ; 
        RECT 20.664 96.676 20.736 97.966 ; 
        RECT 20.196 97.464 20.268 97.902 ; 
        RECT 20.16 94.498 20.232 95.456 ; 
        RECT 20.016 96.822 20.088 97.436 ; 
        RECT 19.692 96.924 19.764 97.956 ; 
        RECT 17.532 94.368 17.604 98.11 ; 
        RECT 17.388 94.368 17.46 98.11 ; 
        RECT 17.244 95.092 17.316 97.364 ; 
        RECT 20.952 98.688 21.024 102.43 ; 
        RECT 20.808 98.688 20.88 102.43 ; 
        RECT 20.664 100.996 20.736 102.286 ; 
        RECT 20.196 101.784 20.268 102.222 ; 
        RECT 20.16 98.818 20.232 99.776 ; 
        RECT 20.016 101.142 20.088 101.756 ; 
        RECT 19.692 101.244 19.764 102.276 ; 
        RECT 17.532 98.688 17.604 102.43 ; 
        RECT 17.388 98.688 17.46 102.43 ; 
        RECT 17.244 99.412 17.316 101.684 ; 
        RECT 20.952 103.008 21.024 106.75 ; 
        RECT 20.808 103.008 20.88 106.75 ; 
        RECT 20.664 105.316 20.736 106.606 ; 
        RECT 20.196 106.104 20.268 106.542 ; 
        RECT 20.16 103.138 20.232 104.096 ; 
        RECT 20.016 105.462 20.088 106.076 ; 
        RECT 19.692 105.564 19.764 106.596 ; 
        RECT 17.532 103.008 17.604 106.75 ; 
        RECT 17.388 103.008 17.46 106.75 ; 
        RECT 17.244 103.732 17.316 106.004 ; 
        RECT 20.952 107.328 21.024 111.07 ; 
        RECT 20.808 107.328 20.88 111.07 ; 
        RECT 20.664 109.636 20.736 110.926 ; 
        RECT 20.196 110.424 20.268 110.862 ; 
        RECT 20.16 107.458 20.232 108.416 ; 
        RECT 20.016 109.782 20.088 110.396 ; 
        RECT 19.692 109.884 19.764 110.916 ; 
        RECT 17.532 107.328 17.604 111.07 ; 
        RECT 17.388 107.328 17.46 111.07 ; 
        RECT 17.244 108.052 17.316 110.324 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 20.72 1.026 21.232 5.4 ; 
      RECT 20.664 3.688 21.232 4.978 ; 
      RECT 20.072 2.596 20.32 5.4 ; 
      RECT 20.016 3.834 20.32 4.448 ; 
      RECT 20.072 1.026 20.176 5.4 ; 
      RECT 20.072 1.51 20.232 2.468 ; 
      RECT 20.072 1.026 20.32 1.382 ; 
      RECT 18.884 2.828 19.708 5.4 ; 
      RECT 19.604 1.026 19.708 5.4 ; 
      RECT 18.884 3.936 19.764 4.968 ; 
      RECT 18.884 1.026 19.276 5.4 ; 
      RECT 17.216 1.026 17.548 5.4 ; 
      RECT 17.216 1.38 17.604 5.122 ; 
      RECT 38.108 1.026 38.448 5.4 ; 
      RECT 37.532 1.026 37.636 5.4 ; 
      RECT 37.1 1.026 37.204 5.4 ; 
      RECT 36.668 1.026 36.772 5.4 ; 
      RECT 36.236 1.026 36.34 5.4 ; 
      RECT 35.804 1.026 35.908 5.4 ; 
      RECT 35.372 1.026 35.476 5.4 ; 
      RECT 34.94 1.026 35.044 5.4 ; 
      RECT 34.508 1.026 34.612 5.4 ; 
      RECT 34.076 1.026 34.18 5.4 ; 
      RECT 33.644 1.026 33.748 5.4 ; 
      RECT 33.212 1.026 33.316 5.4 ; 
      RECT 32.78 1.026 32.884 5.4 ; 
      RECT 32.348 1.026 32.452 5.4 ; 
      RECT 31.916 1.026 32.02 5.4 ; 
      RECT 31.484 1.026 31.588 5.4 ; 
      RECT 31.052 1.026 31.156 5.4 ; 
      RECT 30.62 1.026 30.724 5.4 ; 
      RECT 30.188 1.026 30.292 5.4 ; 
      RECT 29.756 1.026 29.86 5.4 ; 
      RECT 29.324 1.026 29.428 5.4 ; 
      RECT 28.892 1.026 28.996 5.4 ; 
      RECT 28.46 1.026 28.564 5.4 ; 
      RECT 28.028 1.026 28.132 5.4 ; 
      RECT 27.596 1.026 27.7 5.4 ; 
      RECT 27.164 1.026 27.268 5.4 ; 
      RECT 26.732 1.026 26.836 5.4 ; 
      RECT 26.3 1.026 26.404 5.4 ; 
      RECT 25.868 1.026 25.972 5.4 ; 
      RECT 25.436 1.026 25.54 5.4 ; 
      RECT 25.004 1.026 25.108 5.4 ; 
      RECT 24.572 1.026 24.676 5.4 ; 
      RECT 24.14 1.026 24.244 5.4 ; 
      RECT 23.708 1.026 23.812 5.4 ; 
      RECT 22.856 1.026 23.164 5.4 ; 
      RECT 15.284 1.026 15.592 5.4 ; 
      RECT 14.636 1.026 14.74 5.4 ; 
      RECT 14.204 1.026 14.308 5.4 ; 
      RECT 13.772 1.026 13.876 5.4 ; 
      RECT 13.34 1.026 13.444 5.4 ; 
      RECT 12.908 1.026 13.012 5.4 ; 
      RECT 12.476 1.026 12.58 5.4 ; 
      RECT 12.044 1.026 12.148 5.4 ; 
      RECT 11.612 1.026 11.716 5.4 ; 
      RECT 11.18 1.026 11.284 5.4 ; 
      RECT 10.748 1.026 10.852 5.4 ; 
      RECT 10.316 1.026 10.42 5.4 ; 
      RECT 9.884 1.026 9.988 5.4 ; 
      RECT 9.452 1.026 9.556 5.4 ; 
      RECT 9.02 1.026 9.124 5.4 ; 
      RECT 8.588 1.026 8.692 5.4 ; 
      RECT 8.156 1.026 8.26 5.4 ; 
      RECT 7.724 1.026 7.828 5.4 ; 
      RECT 7.292 1.026 7.396 5.4 ; 
      RECT 6.86 1.026 6.964 5.4 ; 
      RECT 6.428 1.026 6.532 5.4 ; 
      RECT 5.996 1.026 6.1 5.4 ; 
      RECT 5.564 1.026 5.668 5.4 ; 
      RECT 5.132 1.026 5.236 5.4 ; 
      RECT 4.7 1.026 4.804 5.4 ; 
      RECT 4.268 1.026 4.372 5.4 ; 
      RECT 3.836 1.026 3.94 5.4 ; 
      RECT 3.404 1.026 3.508 5.4 ; 
      RECT 2.972 1.026 3.076 5.4 ; 
      RECT 2.54 1.026 2.644 5.4 ; 
      RECT 2.108 1.026 2.212 5.4 ; 
      RECT 1.676 1.026 1.78 5.4 ; 
      RECT 1.244 1.026 1.348 5.4 ; 
      RECT 0.812 1.026 0.916 5.4 ; 
      RECT 0 1.026 0.34 5.4 ; 
      RECT 20.72 5.346 21.232 9.72 ; 
      RECT 20.664 8.008 21.232 9.298 ; 
      RECT 20.072 6.916 20.32 9.72 ; 
      RECT 20.016 8.154 20.32 8.768 ; 
      RECT 20.072 5.346 20.176 9.72 ; 
      RECT 20.072 5.83 20.232 6.788 ; 
      RECT 20.072 5.346 20.32 5.702 ; 
      RECT 18.884 7.148 19.708 9.72 ; 
      RECT 19.604 5.346 19.708 9.72 ; 
      RECT 18.884 8.256 19.764 9.288 ; 
      RECT 18.884 5.346 19.276 9.72 ; 
      RECT 17.216 5.346 17.548 9.72 ; 
      RECT 17.216 5.7 17.604 9.442 ; 
      RECT 38.108 5.346 38.448 9.72 ; 
      RECT 37.532 5.346 37.636 9.72 ; 
      RECT 37.1 5.346 37.204 9.72 ; 
      RECT 36.668 5.346 36.772 9.72 ; 
      RECT 36.236 5.346 36.34 9.72 ; 
      RECT 35.804 5.346 35.908 9.72 ; 
      RECT 35.372 5.346 35.476 9.72 ; 
      RECT 34.94 5.346 35.044 9.72 ; 
      RECT 34.508 5.346 34.612 9.72 ; 
      RECT 34.076 5.346 34.18 9.72 ; 
      RECT 33.644 5.346 33.748 9.72 ; 
      RECT 33.212 5.346 33.316 9.72 ; 
      RECT 32.78 5.346 32.884 9.72 ; 
      RECT 32.348 5.346 32.452 9.72 ; 
      RECT 31.916 5.346 32.02 9.72 ; 
      RECT 31.484 5.346 31.588 9.72 ; 
      RECT 31.052 5.346 31.156 9.72 ; 
      RECT 30.62 5.346 30.724 9.72 ; 
      RECT 30.188 5.346 30.292 9.72 ; 
      RECT 29.756 5.346 29.86 9.72 ; 
      RECT 29.324 5.346 29.428 9.72 ; 
      RECT 28.892 5.346 28.996 9.72 ; 
      RECT 28.46 5.346 28.564 9.72 ; 
      RECT 28.028 5.346 28.132 9.72 ; 
      RECT 27.596 5.346 27.7 9.72 ; 
      RECT 27.164 5.346 27.268 9.72 ; 
      RECT 26.732 5.346 26.836 9.72 ; 
      RECT 26.3 5.346 26.404 9.72 ; 
      RECT 25.868 5.346 25.972 9.72 ; 
      RECT 25.436 5.346 25.54 9.72 ; 
      RECT 25.004 5.346 25.108 9.72 ; 
      RECT 24.572 5.346 24.676 9.72 ; 
      RECT 24.14 5.346 24.244 9.72 ; 
      RECT 23.708 5.346 23.812 9.72 ; 
      RECT 22.856 5.346 23.164 9.72 ; 
      RECT 15.284 5.346 15.592 9.72 ; 
      RECT 14.636 5.346 14.74 9.72 ; 
      RECT 14.204 5.346 14.308 9.72 ; 
      RECT 13.772 5.346 13.876 9.72 ; 
      RECT 13.34 5.346 13.444 9.72 ; 
      RECT 12.908 5.346 13.012 9.72 ; 
      RECT 12.476 5.346 12.58 9.72 ; 
      RECT 12.044 5.346 12.148 9.72 ; 
      RECT 11.612 5.346 11.716 9.72 ; 
      RECT 11.18 5.346 11.284 9.72 ; 
      RECT 10.748 5.346 10.852 9.72 ; 
      RECT 10.316 5.346 10.42 9.72 ; 
      RECT 9.884 5.346 9.988 9.72 ; 
      RECT 9.452 5.346 9.556 9.72 ; 
      RECT 9.02 5.346 9.124 9.72 ; 
      RECT 8.588 5.346 8.692 9.72 ; 
      RECT 8.156 5.346 8.26 9.72 ; 
      RECT 7.724 5.346 7.828 9.72 ; 
      RECT 7.292 5.346 7.396 9.72 ; 
      RECT 6.86 5.346 6.964 9.72 ; 
      RECT 6.428 5.346 6.532 9.72 ; 
      RECT 5.996 5.346 6.1 9.72 ; 
      RECT 5.564 5.346 5.668 9.72 ; 
      RECT 5.132 5.346 5.236 9.72 ; 
      RECT 4.7 5.346 4.804 9.72 ; 
      RECT 4.268 5.346 4.372 9.72 ; 
      RECT 3.836 5.346 3.94 9.72 ; 
      RECT 3.404 5.346 3.508 9.72 ; 
      RECT 2.972 5.346 3.076 9.72 ; 
      RECT 2.54 5.346 2.644 9.72 ; 
      RECT 2.108 5.346 2.212 9.72 ; 
      RECT 1.676 5.346 1.78 9.72 ; 
      RECT 1.244 5.346 1.348 9.72 ; 
      RECT 0.812 5.346 0.916 9.72 ; 
      RECT 0 5.346 0.34 9.72 ; 
      RECT 20.72 9.666 21.232 14.04 ; 
      RECT 20.664 12.328 21.232 13.618 ; 
      RECT 20.072 11.236 20.32 14.04 ; 
      RECT 20.016 12.474 20.32 13.088 ; 
      RECT 20.072 9.666 20.176 14.04 ; 
      RECT 20.072 10.15 20.232 11.108 ; 
      RECT 20.072 9.666 20.32 10.022 ; 
      RECT 18.884 11.468 19.708 14.04 ; 
      RECT 19.604 9.666 19.708 14.04 ; 
      RECT 18.884 12.576 19.764 13.608 ; 
      RECT 18.884 9.666 19.276 14.04 ; 
      RECT 17.216 9.666 17.548 14.04 ; 
      RECT 17.216 10.02 17.604 13.762 ; 
      RECT 38.108 9.666 38.448 14.04 ; 
      RECT 37.532 9.666 37.636 14.04 ; 
      RECT 37.1 9.666 37.204 14.04 ; 
      RECT 36.668 9.666 36.772 14.04 ; 
      RECT 36.236 9.666 36.34 14.04 ; 
      RECT 35.804 9.666 35.908 14.04 ; 
      RECT 35.372 9.666 35.476 14.04 ; 
      RECT 34.94 9.666 35.044 14.04 ; 
      RECT 34.508 9.666 34.612 14.04 ; 
      RECT 34.076 9.666 34.18 14.04 ; 
      RECT 33.644 9.666 33.748 14.04 ; 
      RECT 33.212 9.666 33.316 14.04 ; 
      RECT 32.78 9.666 32.884 14.04 ; 
      RECT 32.348 9.666 32.452 14.04 ; 
      RECT 31.916 9.666 32.02 14.04 ; 
      RECT 31.484 9.666 31.588 14.04 ; 
      RECT 31.052 9.666 31.156 14.04 ; 
      RECT 30.62 9.666 30.724 14.04 ; 
      RECT 30.188 9.666 30.292 14.04 ; 
      RECT 29.756 9.666 29.86 14.04 ; 
      RECT 29.324 9.666 29.428 14.04 ; 
      RECT 28.892 9.666 28.996 14.04 ; 
      RECT 28.46 9.666 28.564 14.04 ; 
      RECT 28.028 9.666 28.132 14.04 ; 
      RECT 27.596 9.666 27.7 14.04 ; 
      RECT 27.164 9.666 27.268 14.04 ; 
      RECT 26.732 9.666 26.836 14.04 ; 
      RECT 26.3 9.666 26.404 14.04 ; 
      RECT 25.868 9.666 25.972 14.04 ; 
      RECT 25.436 9.666 25.54 14.04 ; 
      RECT 25.004 9.666 25.108 14.04 ; 
      RECT 24.572 9.666 24.676 14.04 ; 
      RECT 24.14 9.666 24.244 14.04 ; 
      RECT 23.708 9.666 23.812 14.04 ; 
      RECT 22.856 9.666 23.164 14.04 ; 
      RECT 15.284 9.666 15.592 14.04 ; 
      RECT 14.636 9.666 14.74 14.04 ; 
      RECT 14.204 9.666 14.308 14.04 ; 
      RECT 13.772 9.666 13.876 14.04 ; 
      RECT 13.34 9.666 13.444 14.04 ; 
      RECT 12.908 9.666 13.012 14.04 ; 
      RECT 12.476 9.666 12.58 14.04 ; 
      RECT 12.044 9.666 12.148 14.04 ; 
      RECT 11.612 9.666 11.716 14.04 ; 
      RECT 11.18 9.666 11.284 14.04 ; 
      RECT 10.748 9.666 10.852 14.04 ; 
      RECT 10.316 9.666 10.42 14.04 ; 
      RECT 9.884 9.666 9.988 14.04 ; 
      RECT 9.452 9.666 9.556 14.04 ; 
      RECT 9.02 9.666 9.124 14.04 ; 
      RECT 8.588 9.666 8.692 14.04 ; 
      RECT 8.156 9.666 8.26 14.04 ; 
      RECT 7.724 9.666 7.828 14.04 ; 
      RECT 7.292 9.666 7.396 14.04 ; 
      RECT 6.86 9.666 6.964 14.04 ; 
      RECT 6.428 9.666 6.532 14.04 ; 
      RECT 5.996 9.666 6.1 14.04 ; 
      RECT 5.564 9.666 5.668 14.04 ; 
      RECT 5.132 9.666 5.236 14.04 ; 
      RECT 4.7 9.666 4.804 14.04 ; 
      RECT 4.268 9.666 4.372 14.04 ; 
      RECT 3.836 9.666 3.94 14.04 ; 
      RECT 3.404 9.666 3.508 14.04 ; 
      RECT 2.972 9.666 3.076 14.04 ; 
      RECT 2.54 9.666 2.644 14.04 ; 
      RECT 2.108 9.666 2.212 14.04 ; 
      RECT 1.676 9.666 1.78 14.04 ; 
      RECT 1.244 9.666 1.348 14.04 ; 
      RECT 0.812 9.666 0.916 14.04 ; 
      RECT 0 9.666 0.34 14.04 ; 
      RECT 20.72 13.986 21.232 18.36 ; 
      RECT 20.664 16.648 21.232 17.938 ; 
      RECT 20.072 15.556 20.32 18.36 ; 
      RECT 20.016 16.794 20.32 17.408 ; 
      RECT 20.072 13.986 20.176 18.36 ; 
      RECT 20.072 14.47 20.232 15.428 ; 
      RECT 20.072 13.986 20.32 14.342 ; 
      RECT 18.884 15.788 19.708 18.36 ; 
      RECT 19.604 13.986 19.708 18.36 ; 
      RECT 18.884 16.896 19.764 17.928 ; 
      RECT 18.884 13.986 19.276 18.36 ; 
      RECT 17.216 13.986 17.548 18.36 ; 
      RECT 17.216 14.34 17.604 18.082 ; 
      RECT 38.108 13.986 38.448 18.36 ; 
      RECT 37.532 13.986 37.636 18.36 ; 
      RECT 37.1 13.986 37.204 18.36 ; 
      RECT 36.668 13.986 36.772 18.36 ; 
      RECT 36.236 13.986 36.34 18.36 ; 
      RECT 35.804 13.986 35.908 18.36 ; 
      RECT 35.372 13.986 35.476 18.36 ; 
      RECT 34.94 13.986 35.044 18.36 ; 
      RECT 34.508 13.986 34.612 18.36 ; 
      RECT 34.076 13.986 34.18 18.36 ; 
      RECT 33.644 13.986 33.748 18.36 ; 
      RECT 33.212 13.986 33.316 18.36 ; 
      RECT 32.78 13.986 32.884 18.36 ; 
      RECT 32.348 13.986 32.452 18.36 ; 
      RECT 31.916 13.986 32.02 18.36 ; 
      RECT 31.484 13.986 31.588 18.36 ; 
      RECT 31.052 13.986 31.156 18.36 ; 
      RECT 30.62 13.986 30.724 18.36 ; 
      RECT 30.188 13.986 30.292 18.36 ; 
      RECT 29.756 13.986 29.86 18.36 ; 
      RECT 29.324 13.986 29.428 18.36 ; 
      RECT 28.892 13.986 28.996 18.36 ; 
      RECT 28.46 13.986 28.564 18.36 ; 
      RECT 28.028 13.986 28.132 18.36 ; 
      RECT 27.596 13.986 27.7 18.36 ; 
      RECT 27.164 13.986 27.268 18.36 ; 
      RECT 26.732 13.986 26.836 18.36 ; 
      RECT 26.3 13.986 26.404 18.36 ; 
      RECT 25.868 13.986 25.972 18.36 ; 
      RECT 25.436 13.986 25.54 18.36 ; 
      RECT 25.004 13.986 25.108 18.36 ; 
      RECT 24.572 13.986 24.676 18.36 ; 
      RECT 24.14 13.986 24.244 18.36 ; 
      RECT 23.708 13.986 23.812 18.36 ; 
      RECT 22.856 13.986 23.164 18.36 ; 
      RECT 15.284 13.986 15.592 18.36 ; 
      RECT 14.636 13.986 14.74 18.36 ; 
      RECT 14.204 13.986 14.308 18.36 ; 
      RECT 13.772 13.986 13.876 18.36 ; 
      RECT 13.34 13.986 13.444 18.36 ; 
      RECT 12.908 13.986 13.012 18.36 ; 
      RECT 12.476 13.986 12.58 18.36 ; 
      RECT 12.044 13.986 12.148 18.36 ; 
      RECT 11.612 13.986 11.716 18.36 ; 
      RECT 11.18 13.986 11.284 18.36 ; 
      RECT 10.748 13.986 10.852 18.36 ; 
      RECT 10.316 13.986 10.42 18.36 ; 
      RECT 9.884 13.986 9.988 18.36 ; 
      RECT 9.452 13.986 9.556 18.36 ; 
      RECT 9.02 13.986 9.124 18.36 ; 
      RECT 8.588 13.986 8.692 18.36 ; 
      RECT 8.156 13.986 8.26 18.36 ; 
      RECT 7.724 13.986 7.828 18.36 ; 
      RECT 7.292 13.986 7.396 18.36 ; 
      RECT 6.86 13.986 6.964 18.36 ; 
      RECT 6.428 13.986 6.532 18.36 ; 
      RECT 5.996 13.986 6.1 18.36 ; 
      RECT 5.564 13.986 5.668 18.36 ; 
      RECT 5.132 13.986 5.236 18.36 ; 
      RECT 4.7 13.986 4.804 18.36 ; 
      RECT 4.268 13.986 4.372 18.36 ; 
      RECT 3.836 13.986 3.94 18.36 ; 
      RECT 3.404 13.986 3.508 18.36 ; 
      RECT 2.972 13.986 3.076 18.36 ; 
      RECT 2.54 13.986 2.644 18.36 ; 
      RECT 2.108 13.986 2.212 18.36 ; 
      RECT 1.676 13.986 1.78 18.36 ; 
      RECT 1.244 13.986 1.348 18.36 ; 
      RECT 0.812 13.986 0.916 18.36 ; 
      RECT 0 13.986 0.34 18.36 ; 
      RECT 20.72 18.306 21.232 22.68 ; 
      RECT 20.664 20.968 21.232 22.258 ; 
      RECT 20.072 19.876 20.32 22.68 ; 
      RECT 20.016 21.114 20.32 21.728 ; 
      RECT 20.072 18.306 20.176 22.68 ; 
      RECT 20.072 18.79 20.232 19.748 ; 
      RECT 20.072 18.306 20.32 18.662 ; 
      RECT 18.884 20.108 19.708 22.68 ; 
      RECT 19.604 18.306 19.708 22.68 ; 
      RECT 18.884 21.216 19.764 22.248 ; 
      RECT 18.884 18.306 19.276 22.68 ; 
      RECT 17.216 18.306 17.548 22.68 ; 
      RECT 17.216 18.66 17.604 22.402 ; 
      RECT 38.108 18.306 38.448 22.68 ; 
      RECT 37.532 18.306 37.636 22.68 ; 
      RECT 37.1 18.306 37.204 22.68 ; 
      RECT 36.668 18.306 36.772 22.68 ; 
      RECT 36.236 18.306 36.34 22.68 ; 
      RECT 35.804 18.306 35.908 22.68 ; 
      RECT 35.372 18.306 35.476 22.68 ; 
      RECT 34.94 18.306 35.044 22.68 ; 
      RECT 34.508 18.306 34.612 22.68 ; 
      RECT 34.076 18.306 34.18 22.68 ; 
      RECT 33.644 18.306 33.748 22.68 ; 
      RECT 33.212 18.306 33.316 22.68 ; 
      RECT 32.78 18.306 32.884 22.68 ; 
      RECT 32.348 18.306 32.452 22.68 ; 
      RECT 31.916 18.306 32.02 22.68 ; 
      RECT 31.484 18.306 31.588 22.68 ; 
      RECT 31.052 18.306 31.156 22.68 ; 
      RECT 30.62 18.306 30.724 22.68 ; 
      RECT 30.188 18.306 30.292 22.68 ; 
      RECT 29.756 18.306 29.86 22.68 ; 
      RECT 29.324 18.306 29.428 22.68 ; 
      RECT 28.892 18.306 28.996 22.68 ; 
      RECT 28.46 18.306 28.564 22.68 ; 
      RECT 28.028 18.306 28.132 22.68 ; 
      RECT 27.596 18.306 27.7 22.68 ; 
      RECT 27.164 18.306 27.268 22.68 ; 
      RECT 26.732 18.306 26.836 22.68 ; 
      RECT 26.3 18.306 26.404 22.68 ; 
      RECT 25.868 18.306 25.972 22.68 ; 
      RECT 25.436 18.306 25.54 22.68 ; 
      RECT 25.004 18.306 25.108 22.68 ; 
      RECT 24.572 18.306 24.676 22.68 ; 
      RECT 24.14 18.306 24.244 22.68 ; 
      RECT 23.708 18.306 23.812 22.68 ; 
      RECT 22.856 18.306 23.164 22.68 ; 
      RECT 15.284 18.306 15.592 22.68 ; 
      RECT 14.636 18.306 14.74 22.68 ; 
      RECT 14.204 18.306 14.308 22.68 ; 
      RECT 13.772 18.306 13.876 22.68 ; 
      RECT 13.34 18.306 13.444 22.68 ; 
      RECT 12.908 18.306 13.012 22.68 ; 
      RECT 12.476 18.306 12.58 22.68 ; 
      RECT 12.044 18.306 12.148 22.68 ; 
      RECT 11.612 18.306 11.716 22.68 ; 
      RECT 11.18 18.306 11.284 22.68 ; 
      RECT 10.748 18.306 10.852 22.68 ; 
      RECT 10.316 18.306 10.42 22.68 ; 
      RECT 9.884 18.306 9.988 22.68 ; 
      RECT 9.452 18.306 9.556 22.68 ; 
      RECT 9.02 18.306 9.124 22.68 ; 
      RECT 8.588 18.306 8.692 22.68 ; 
      RECT 8.156 18.306 8.26 22.68 ; 
      RECT 7.724 18.306 7.828 22.68 ; 
      RECT 7.292 18.306 7.396 22.68 ; 
      RECT 6.86 18.306 6.964 22.68 ; 
      RECT 6.428 18.306 6.532 22.68 ; 
      RECT 5.996 18.306 6.1 22.68 ; 
      RECT 5.564 18.306 5.668 22.68 ; 
      RECT 5.132 18.306 5.236 22.68 ; 
      RECT 4.7 18.306 4.804 22.68 ; 
      RECT 4.268 18.306 4.372 22.68 ; 
      RECT 3.836 18.306 3.94 22.68 ; 
      RECT 3.404 18.306 3.508 22.68 ; 
      RECT 2.972 18.306 3.076 22.68 ; 
      RECT 2.54 18.306 2.644 22.68 ; 
      RECT 2.108 18.306 2.212 22.68 ; 
      RECT 1.676 18.306 1.78 22.68 ; 
      RECT 1.244 18.306 1.348 22.68 ; 
      RECT 0.812 18.306 0.916 22.68 ; 
      RECT 0 18.306 0.34 22.68 ; 
      RECT 20.72 22.626 21.232 27 ; 
      RECT 20.664 25.288 21.232 26.578 ; 
      RECT 20.072 24.196 20.32 27 ; 
      RECT 20.016 25.434 20.32 26.048 ; 
      RECT 20.072 22.626 20.176 27 ; 
      RECT 20.072 23.11 20.232 24.068 ; 
      RECT 20.072 22.626 20.32 22.982 ; 
      RECT 18.884 24.428 19.708 27 ; 
      RECT 19.604 22.626 19.708 27 ; 
      RECT 18.884 25.536 19.764 26.568 ; 
      RECT 18.884 22.626 19.276 27 ; 
      RECT 17.216 22.626 17.548 27 ; 
      RECT 17.216 22.98 17.604 26.722 ; 
      RECT 38.108 22.626 38.448 27 ; 
      RECT 37.532 22.626 37.636 27 ; 
      RECT 37.1 22.626 37.204 27 ; 
      RECT 36.668 22.626 36.772 27 ; 
      RECT 36.236 22.626 36.34 27 ; 
      RECT 35.804 22.626 35.908 27 ; 
      RECT 35.372 22.626 35.476 27 ; 
      RECT 34.94 22.626 35.044 27 ; 
      RECT 34.508 22.626 34.612 27 ; 
      RECT 34.076 22.626 34.18 27 ; 
      RECT 33.644 22.626 33.748 27 ; 
      RECT 33.212 22.626 33.316 27 ; 
      RECT 32.78 22.626 32.884 27 ; 
      RECT 32.348 22.626 32.452 27 ; 
      RECT 31.916 22.626 32.02 27 ; 
      RECT 31.484 22.626 31.588 27 ; 
      RECT 31.052 22.626 31.156 27 ; 
      RECT 30.62 22.626 30.724 27 ; 
      RECT 30.188 22.626 30.292 27 ; 
      RECT 29.756 22.626 29.86 27 ; 
      RECT 29.324 22.626 29.428 27 ; 
      RECT 28.892 22.626 28.996 27 ; 
      RECT 28.46 22.626 28.564 27 ; 
      RECT 28.028 22.626 28.132 27 ; 
      RECT 27.596 22.626 27.7 27 ; 
      RECT 27.164 22.626 27.268 27 ; 
      RECT 26.732 22.626 26.836 27 ; 
      RECT 26.3 22.626 26.404 27 ; 
      RECT 25.868 22.626 25.972 27 ; 
      RECT 25.436 22.626 25.54 27 ; 
      RECT 25.004 22.626 25.108 27 ; 
      RECT 24.572 22.626 24.676 27 ; 
      RECT 24.14 22.626 24.244 27 ; 
      RECT 23.708 22.626 23.812 27 ; 
      RECT 22.856 22.626 23.164 27 ; 
      RECT 15.284 22.626 15.592 27 ; 
      RECT 14.636 22.626 14.74 27 ; 
      RECT 14.204 22.626 14.308 27 ; 
      RECT 13.772 22.626 13.876 27 ; 
      RECT 13.34 22.626 13.444 27 ; 
      RECT 12.908 22.626 13.012 27 ; 
      RECT 12.476 22.626 12.58 27 ; 
      RECT 12.044 22.626 12.148 27 ; 
      RECT 11.612 22.626 11.716 27 ; 
      RECT 11.18 22.626 11.284 27 ; 
      RECT 10.748 22.626 10.852 27 ; 
      RECT 10.316 22.626 10.42 27 ; 
      RECT 9.884 22.626 9.988 27 ; 
      RECT 9.452 22.626 9.556 27 ; 
      RECT 9.02 22.626 9.124 27 ; 
      RECT 8.588 22.626 8.692 27 ; 
      RECT 8.156 22.626 8.26 27 ; 
      RECT 7.724 22.626 7.828 27 ; 
      RECT 7.292 22.626 7.396 27 ; 
      RECT 6.86 22.626 6.964 27 ; 
      RECT 6.428 22.626 6.532 27 ; 
      RECT 5.996 22.626 6.1 27 ; 
      RECT 5.564 22.626 5.668 27 ; 
      RECT 5.132 22.626 5.236 27 ; 
      RECT 4.7 22.626 4.804 27 ; 
      RECT 4.268 22.626 4.372 27 ; 
      RECT 3.836 22.626 3.94 27 ; 
      RECT 3.404 22.626 3.508 27 ; 
      RECT 2.972 22.626 3.076 27 ; 
      RECT 2.54 22.626 2.644 27 ; 
      RECT 2.108 22.626 2.212 27 ; 
      RECT 1.676 22.626 1.78 27 ; 
      RECT 1.244 22.626 1.348 27 ; 
      RECT 0.812 22.626 0.916 27 ; 
      RECT 0 22.626 0.34 27 ; 
      RECT 20.72 26.946 21.232 31.32 ; 
      RECT 20.664 29.608 21.232 30.898 ; 
      RECT 20.072 28.516 20.32 31.32 ; 
      RECT 20.016 29.754 20.32 30.368 ; 
      RECT 20.072 26.946 20.176 31.32 ; 
      RECT 20.072 27.43 20.232 28.388 ; 
      RECT 20.072 26.946 20.32 27.302 ; 
      RECT 18.884 28.748 19.708 31.32 ; 
      RECT 19.604 26.946 19.708 31.32 ; 
      RECT 18.884 29.856 19.764 30.888 ; 
      RECT 18.884 26.946 19.276 31.32 ; 
      RECT 17.216 26.946 17.548 31.32 ; 
      RECT 17.216 27.3 17.604 31.042 ; 
      RECT 38.108 26.946 38.448 31.32 ; 
      RECT 37.532 26.946 37.636 31.32 ; 
      RECT 37.1 26.946 37.204 31.32 ; 
      RECT 36.668 26.946 36.772 31.32 ; 
      RECT 36.236 26.946 36.34 31.32 ; 
      RECT 35.804 26.946 35.908 31.32 ; 
      RECT 35.372 26.946 35.476 31.32 ; 
      RECT 34.94 26.946 35.044 31.32 ; 
      RECT 34.508 26.946 34.612 31.32 ; 
      RECT 34.076 26.946 34.18 31.32 ; 
      RECT 33.644 26.946 33.748 31.32 ; 
      RECT 33.212 26.946 33.316 31.32 ; 
      RECT 32.78 26.946 32.884 31.32 ; 
      RECT 32.348 26.946 32.452 31.32 ; 
      RECT 31.916 26.946 32.02 31.32 ; 
      RECT 31.484 26.946 31.588 31.32 ; 
      RECT 31.052 26.946 31.156 31.32 ; 
      RECT 30.62 26.946 30.724 31.32 ; 
      RECT 30.188 26.946 30.292 31.32 ; 
      RECT 29.756 26.946 29.86 31.32 ; 
      RECT 29.324 26.946 29.428 31.32 ; 
      RECT 28.892 26.946 28.996 31.32 ; 
      RECT 28.46 26.946 28.564 31.32 ; 
      RECT 28.028 26.946 28.132 31.32 ; 
      RECT 27.596 26.946 27.7 31.32 ; 
      RECT 27.164 26.946 27.268 31.32 ; 
      RECT 26.732 26.946 26.836 31.32 ; 
      RECT 26.3 26.946 26.404 31.32 ; 
      RECT 25.868 26.946 25.972 31.32 ; 
      RECT 25.436 26.946 25.54 31.32 ; 
      RECT 25.004 26.946 25.108 31.32 ; 
      RECT 24.572 26.946 24.676 31.32 ; 
      RECT 24.14 26.946 24.244 31.32 ; 
      RECT 23.708 26.946 23.812 31.32 ; 
      RECT 22.856 26.946 23.164 31.32 ; 
      RECT 15.284 26.946 15.592 31.32 ; 
      RECT 14.636 26.946 14.74 31.32 ; 
      RECT 14.204 26.946 14.308 31.32 ; 
      RECT 13.772 26.946 13.876 31.32 ; 
      RECT 13.34 26.946 13.444 31.32 ; 
      RECT 12.908 26.946 13.012 31.32 ; 
      RECT 12.476 26.946 12.58 31.32 ; 
      RECT 12.044 26.946 12.148 31.32 ; 
      RECT 11.612 26.946 11.716 31.32 ; 
      RECT 11.18 26.946 11.284 31.32 ; 
      RECT 10.748 26.946 10.852 31.32 ; 
      RECT 10.316 26.946 10.42 31.32 ; 
      RECT 9.884 26.946 9.988 31.32 ; 
      RECT 9.452 26.946 9.556 31.32 ; 
      RECT 9.02 26.946 9.124 31.32 ; 
      RECT 8.588 26.946 8.692 31.32 ; 
      RECT 8.156 26.946 8.26 31.32 ; 
      RECT 7.724 26.946 7.828 31.32 ; 
      RECT 7.292 26.946 7.396 31.32 ; 
      RECT 6.86 26.946 6.964 31.32 ; 
      RECT 6.428 26.946 6.532 31.32 ; 
      RECT 5.996 26.946 6.1 31.32 ; 
      RECT 5.564 26.946 5.668 31.32 ; 
      RECT 5.132 26.946 5.236 31.32 ; 
      RECT 4.7 26.946 4.804 31.32 ; 
      RECT 4.268 26.946 4.372 31.32 ; 
      RECT 3.836 26.946 3.94 31.32 ; 
      RECT 3.404 26.946 3.508 31.32 ; 
      RECT 2.972 26.946 3.076 31.32 ; 
      RECT 2.54 26.946 2.644 31.32 ; 
      RECT 2.108 26.946 2.212 31.32 ; 
      RECT 1.676 26.946 1.78 31.32 ; 
      RECT 1.244 26.946 1.348 31.32 ; 
      RECT 0.812 26.946 0.916 31.32 ; 
      RECT 0 26.946 0.34 31.32 ; 
      RECT 20.72 31.266 21.232 35.64 ; 
      RECT 20.664 33.928 21.232 35.218 ; 
      RECT 20.072 32.836 20.32 35.64 ; 
      RECT 20.016 34.074 20.32 34.688 ; 
      RECT 20.072 31.266 20.176 35.64 ; 
      RECT 20.072 31.75 20.232 32.708 ; 
      RECT 20.072 31.266 20.32 31.622 ; 
      RECT 18.884 33.068 19.708 35.64 ; 
      RECT 19.604 31.266 19.708 35.64 ; 
      RECT 18.884 34.176 19.764 35.208 ; 
      RECT 18.884 31.266 19.276 35.64 ; 
      RECT 17.216 31.266 17.548 35.64 ; 
      RECT 17.216 31.62 17.604 35.362 ; 
      RECT 38.108 31.266 38.448 35.64 ; 
      RECT 37.532 31.266 37.636 35.64 ; 
      RECT 37.1 31.266 37.204 35.64 ; 
      RECT 36.668 31.266 36.772 35.64 ; 
      RECT 36.236 31.266 36.34 35.64 ; 
      RECT 35.804 31.266 35.908 35.64 ; 
      RECT 35.372 31.266 35.476 35.64 ; 
      RECT 34.94 31.266 35.044 35.64 ; 
      RECT 34.508 31.266 34.612 35.64 ; 
      RECT 34.076 31.266 34.18 35.64 ; 
      RECT 33.644 31.266 33.748 35.64 ; 
      RECT 33.212 31.266 33.316 35.64 ; 
      RECT 32.78 31.266 32.884 35.64 ; 
      RECT 32.348 31.266 32.452 35.64 ; 
      RECT 31.916 31.266 32.02 35.64 ; 
      RECT 31.484 31.266 31.588 35.64 ; 
      RECT 31.052 31.266 31.156 35.64 ; 
      RECT 30.62 31.266 30.724 35.64 ; 
      RECT 30.188 31.266 30.292 35.64 ; 
      RECT 29.756 31.266 29.86 35.64 ; 
      RECT 29.324 31.266 29.428 35.64 ; 
      RECT 28.892 31.266 28.996 35.64 ; 
      RECT 28.46 31.266 28.564 35.64 ; 
      RECT 28.028 31.266 28.132 35.64 ; 
      RECT 27.596 31.266 27.7 35.64 ; 
      RECT 27.164 31.266 27.268 35.64 ; 
      RECT 26.732 31.266 26.836 35.64 ; 
      RECT 26.3 31.266 26.404 35.64 ; 
      RECT 25.868 31.266 25.972 35.64 ; 
      RECT 25.436 31.266 25.54 35.64 ; 
      RECT 25.004 31.266 25.108 35.64 ; 
      RECT 24.572 31.266 24.676 35.64 ; 
      RECT 24.14 31.266 24.244 35.64 ; 
      RECT 23.708 31.266 23.812 35.64 ; 
      RECT 22.856 31.266 23.164 35.64 ; 
      RECT 15.284 31.266 15.592 35.64 ; 
      RECT 14.636 31.266 14.74 35.64 ; 
      RECT 14.204 31.266 14.308 35.64 ; 
      RECT 13.772 31.266 13.876 35.64 ; 
      RECT 13.34 31.266 13.444 35.64 ; 
      RECT 12.908 31.266 13.012 35.64 ; 
      RECT 12.476 31.266 12.58 35.64 ; 
      RECT 12.044 31.266 12.148 35.64 ; 
      RECT 11.612 31.266 11.716 35.64 ; 
      RECT 11.18 31.266 11.284 35.64 ; 
      RECT 10.748 31.266 10.852 35.64 ; 
      RECT 10.316 31.266 10.42 35.64 ; 
      RECT 9.884 31.266 9.988 35.64 ; 
      RECT 9.452 31.266 9.556 35.64 ; 
      RECT 9.02 31.266 9.124 35.64 ; 
      RECT 8.588 31.266 8.692 35.64 ; 
      RECT 8.156 31.266 8.26 35.64 ; 
      RECT 7.724 31.266 7.828 35.64 ; 
      RECT 7.292 31.266 7.396 35.64 ; 
      RECT 6.86 31.266 6.964 35.64 ; 
      RECT 6.428 31.266 6.532 35.64 ; 
      RECT 5.996 31.266 6.1 35.64 ; 
      RECT 5.564 31.266 5.668 35.64 ; 
      RECT 5.132 31.266 5.236 35.64 ; 
      RECT 4.7 31.266 4.804 35.64 ; 
      RECT 4.268 31.266 4.372 35.64 ; 
      RECT 3.836 31.266 3.94 35.64 ; 
      RECT 3.404 31.266 3.508 35.64 ; 
      RECT 2.972 31.266 3.076 35.64 ; 
      RECT 2.54 31.266 2.644 35.64 ; 
      RECT 2.108 31.266 2.212 35.64 ; 
      RECT 1.676 31.266 1.78 35.64 ; 
      RECT 1.244 31.266 1.348 35.64 ; 
      RECT 0.812 31.266 0.916 35.64 ; 
      RECT 0 31.266 0.34 35.64 ; 
      RECT 20.72 35.586 21.232 39.96 ; 
      RECT 20.664 38.248 21.232 39.538 ; 
      RECT 20.072 37.156 20.32 39.96 ; 
      RECT 20.016 38.394 20.32 39.008 ; 
      RECT 20.072 35.586 20.176 39.96 ; 
      RECT 20.072 36.07 20.232 37.028 ; 
      RECT 20.072 35.586 20.32 35.942 ; 
      RECT 18.884 37.388 19.708 39.96 ; 
      RECT 19.604 35.586 19.708 39.96 ; 
      RECT 18.884 38.496 19.764 39.528 ; 
      RECT 18.884 35.586 19.276 39.96 ; 
      RECT 17.216 35.586 17.548 39.96 ; 
      RECT 17.216 35.94 17.604 39.682 ; 
      RECT 38.108 35.586 38.448 39.96 ; 
      RECT 37.532 35.586 37.636 39.96 ; 
      RECT 37.1 35.586 37.204 39.96 ; 
      RECT 36.668 35.586 36.772 39.96 ; 
      RECT 36.236 35.586 36.34 39.96 ; 
      RECT 35.804 35.586 35.908 39.96 ; 
      RECT 35.372 35.586 35.476 39.96 ; 
      RECT 34.94 35.586 35.044 39.96 ; 
      RECT 34.508 35.586 34.612 39.96 ; 
      RECT 34.076 35.586 34.18 39.96 ; 
      RECT 33.644 35.586 33.748 39.96 ; 
      RECT 33.212 35.586 33.316 39.96 ; 
      RECT 32.78 35.586 32.884 39.96 ; 
      RECT 32.348 35.586 32.452 39.96 ; 
      RECT 31.916 35.586 32.02 39.96 ; 
      RECT 31.484 35.586 31.588 39.96 ; 
      RECT 31.052 35.586 31.156 39.96 ; 
      RECT 30.62 35.586 30.724 39.96 ; 
      RECT 30.188 35.586 30.292 39.96 ; 
      RECT 29.756 35.586 29.86 39.96 ; 
      RECT 29.324 35.586 29.428 39.96 ; 
      RECT 28.892 35.586 28.996 39.96 ; 
      RECT 28.46 35.586 28.564 39.96 ; 
      RECT 28.028 35.586 28.132 39.96 ; 
      RECT 27.596 35.586 27.7 39.96 ; 
      RECT 27.164 35.586 27.268 39.96 ; 
      RECT 26.732 35.586 26.836 39.96 ; 
      RECT 26.3 35.586 26.404 39.96 ; 
      RECT 25.868 35.586 25.972 39.96 ; 
      RECT 25.436 35.586 25.54 39.96 ; 
      RECT 25.004 35.586 25.108 39.96 ; 
      RECT 24.572 35.586 24.676 39.96 ; 
      RECT 24.14 35.586 24.244 39.96 ; 
      RECT 23.708 35.586 23.812 39.96 ; 
      RECT 22.856 35.586 23.164 39.96 ; 
      RECT 15.284 35.586 15.592 39.96 ; 
      RECT 14.636 35.586 14.74 39.96 ; 
      RECT 14.204 35.586 14.308 39.96 ; 
      RECT 13.772 35.586 13.876 39.96 ; 
      RECT 13.34 35.586 13.444 39.96 ; 
      RECT 12.908 35.586 13.012 39.96 ; 
      RECT 12.476 35.586 12.58 39.96 ; 
      RECT 12.044 35.586 12.148 39.96 ; 
      RECT 11.612 35.586 11.716 39.96 ; 
      RECT 11.18 35.586 11.284 39.96 ; 
      RECT 10.748 35.586 10.852 39.96 ; 
      RECT 10.316 35.586 10.42 39.96 ; 
      RECT 9.884 35.586 9.988 39.96 ; 
      RECT 9.452 35.586 9.556 39.96 ; 
      RECT 9.02 35.586 9.124 39.96 ; 
      RECT 8.588 35.586 8.692 39.96 ; 
      RECT 8.156 35.586 8.26 39.96 ; 
      RECT 7.724 35.586 7.828 39.96 ; 
      RECT 7.292 35.586 7.396 39.96 ; 
      RECT 6.86 35.586 6.964 39.96 ; 
      RECT 6.428 35.586 6.532 39.96 ; 
      RECT 5.996 35.586 6.1 39.96 ; 
      RECT 5.564 35.586 5.668 39.96 ; 
      RECT 5.132 35.586 5.236 39.96 ; 
      RECT 4.7 35.586 4.804 39.96 ; 
      RECT 4.268 35.586 4.372 39.96 ; 
      RECT 3.836 35.586 3.94 39.96 ; 
      RECT 3.404 35.586 3.508 39.96 ; 
      RECT 2.972 35.586 3.076 39.96 ; 
      RECT 2.54 35.586 2.644 39.96 ; 
      RECT 2.108 35.586 2.212 39.96 ; 
      RECT 1.676 35.586 1.78 39.96 ; 
      RECT 1.244 35.586 1.348 39.96 ; 
      RECT 0.812 35.586 0.916 39.96 ; 
      RECT 0 35.586 0.34 39.96 ; 
      RECT 0 73.296 38.448 74.466 ; 
      RECT 38.108 39.852 38.448 74.466 ; 
      RECT 18.164 72.702 38.448 74.466 ; 
      RECT 0 72.702 17.548 74.466 ; 
      RECT 23.708 45.868 37.636 74.466 ; 
      RECT 29.54 39.852 37.636 74.466 ; 
      RECT 18.164 72.596 23.38 74.466 ; 
      RECT 20.72 72.592 23.38 74.466 ; 
      RECT 15.068 46.3 17.548 74.466 ; 
      RECT 15.284 42.916 17.548 74.466 ; 
      RECT 0.812 45.088 14.74 74.466 ; 
      RECT 13.556 39.852 14.74 74.466 ; 
      RECT 0 39.852 0.34 74.466 ; 
      RECT 18.164 72.584 20.32 74.466 ; 
      RECT 20.072 71.5 20.32 74.466 ; 
      RECT 20.72 71.5 23.164 74.466 ; 
      RECT 18.164 71.5 19.708 74.466 ; 
      RECT 23.652 55.024 37.636 72.464 ; 
      RECT 0.812 55.024 14.796 72.464 ; 
      RECT 23.652 55.024 37.692 72.446 ; 
      RECT 0.756 55.024 14.796 72.446 ; 
      RECT 20.756 42.916 23.164 74.466 ; 
      RECT 18.884 42.592 19.564 74.466 ; 
      RECT 19.316 39.852 19.564 74.466 ; 
      RECT 16.148 42.188 17.692 70.9 ; 
      RECT 15.068 70.732 17.748 70.88 ; 
      RECT 20.7 66.436 23.164 70.868 ; 
      RECT 18.828 69.676 19.564 70.58 ; 
      RECT 18.884 67.372 19.62 68.42 ; 
      RECT 15.068 66.58 17.748 68.42 ; 
      RECT 18.828 64.42 19.564 66.26 ; 
      RECT 20.7 56.284 23.164 65.612 ; 
      RECT 15.068 58.876 17.748 63.452 ; 
      RECT 18.884 57.796 19.62 63.02 ; 
      RECT 18.828 60.1 19.62 61.94 ; 
      RECT 18.828 47.14 19.564 59.78 ; 
      RECT 18.828 47.14 19.62 57.62 ; 
      RECT 15.068 56.716 17.748 57.62 ; 
      RECT 20.9 40.558 23.38 54.896 ; 
      RECT 20.7 44.98 23.38 52.124 ; 
      RECT 15.068 48.868 17.748 50.348 ; 
      RECT 18.884 46.06 19.62 46.82 ; 
      RECT 15.284 45.916 17.748 46.676 ; 
      RECT 18.828 45.484 19.564 46.028 ; 
      RECT 18.884 44.98 19.62 45.884 ; 
      RECT 24.356 45.1 37.636 74.466 ; 
      RECT 28.676 45.088 37.636 74.466 ; 
      RECT 23.708 39.852 24.028 74.466 ; 
      RECT 15.068 42.592 15.82 45.848 ; 
      RECT 23.708 39.852 24.892 45.464 ; 
      RECT 23.708 44.32 28.348 45.464 ; 
      RECT 28.676 39.852 29.212 74.466 ; 
      RECT 10.1 43.564 13.228 74.466 ; 
      RECT 0.812 39.852 9.772 74.466 ; 
      RECT 23.708 44.32 29.212 44.696 ; 
      RECT 27.812 39.852 37.636 44.684 ; 
      RECT 12.692 39.852 14.74 44.684 ; 
      RECT 18.828 44.404 19.62 44.66 ; 
      RECT 18.828 43.9 19.564 44.66 ; 
      RECT 26.948 42.784 37.636 44.684 ; 
      RECT 23.708 42.916 26.62 45.464 ; 
      RECT 18.884 42.82 19.62 43.868 ; 
      RECT 0.812 42.784 12.364 44.684 ; 
      RECT 11.828 39.852 12.364 74.466 ; 
      RECT 26.084 39.852 27.484 43.34 ; 
      RECT 23.708 42.592 25.756 45.464 ; 
      RECT 25.22 39.852 25.756 74.466 ; 
      RECT 10.964 42.592 12.364 74.466 ; 
      RECT 0.812 39.852 10.636 44.684 ; 
      RECT 18.884 39.852 18.988 74.466 ; 
      RECT 15.428 39.852 15.82 74.466 ; 
      RECT 10.964 39.852 11.5 74.466 ; 
      RECT 25.22 39.852 27.484 42.392 ; 
      RECT 20.756 39.852 23.164 42.392 ; 
      RECT 15.428 39.852 17.548 42.392 ; 
      RECT 11.828 39.852 14.74 42.392 ; 
      RECT 25.22 39.852 37.636 42.38 ; 
      RECT 0.812 39.852 11.5 42.38 ; 
      RECT 20.7 41.74 23.38 42.356 ; 
      RECT 15.428 41.74 17.604 42.392 ; 
      RECT 23.708 39.852 37.636 41.324 ; 
      RECT 18.884 39.852 19.564 41.324 ; 
      RECT 15.068 39.852 17.548 41.324 ; 
      RECT 0.812 39.852 14.74 41.324 ; 
      RECT 18.164 39.852 19.564 40.912 ; 
      RECT 20.72 39.852 23.164 40.512 ; 
      RECT 18.164 39.852 19.708 40.512 ; 
      RECT 20.72 39.852 23.38 39.936 ; 
      RECT 25.236 39.746 25.308 74.466 ; 
      RECT 24.804 39.746 24.876 74.466 ; 
      RECT 11.844 39.746 11.916 74.466 ; 
      RECT 11.412 39.746 11.484 74.466 ; 
      RECT 20.072 39.852 20.32 40.512 ; 
        RECT 20.72 72.414 21.232 76.788 ; 
        RECT 20.664 75.076 21.232 76.366 ; 
        RECT 20.072 73.984 20.32 76.788 ; 
        RECT 20.016 75.222 20.32 75.836 ; 
        RECT 20.072 72.414 20.176 76.788 ; 
        RECT 20.072 72.898 20.232 73.856 ; 
        RECT 20.072 72.414 20.32 72.77 ; 
        RECT 18.884 74.216 19.708 76.788 ; 
        RECT 19.604 72.414 19.708 76.788 ; 
        RECT 18.884 75.324 19.764 76.356 ; 
        RECT 18.884 72.414 19.276 76.788 ; 
        RECT 17.216 72.414 17.548 76.788 ; 
        RECT 17.216 72.768 17.604 76.51 ; 
        RECT 38.108 72.414 38.448 76.788 ; 
        RECT 37.532 72.414 37.636 76.788 ; 
        RECT 37.1 72.414 37.204 76.788 ; 
        RECT 36.668 72.414 36.772 76.788 ; 
        RECT 36.236 72.414 36.34 76.788 ; 
        RECT 35.804 72.414 35.908 76.788 ; 
        RECT 35.372 72.414 35.476 76.788 ; 
        RECT 34.94 72.414 35.044 76.788 ; 
        RECT 34.508 72.414 34.612 76.788 ; 
        RECT 34.076 72.414 34.18 76.788 ; 
        RECT 33.644 72.414 33.748 76.788 ; 
        RECT 33.212 72.414 33.316 76.788 ; 
        RECT 32.78 72.414 32.884 76.788 ; 
        RECT 32.348 72.414 32.452 76.788 ; 
        RECT 31.916 72.414 32.02 76.788 ; 
        RECT 31.484 72.414 31.588 76.788 ; 
        RECT 31.052 72.414 31.156 76.788 ; 
        RECT 30.62 72.414 30.724 76.788 ; 
        RECT 30.188 72.414 30.292 76.788 ; 
        RECT 29.756 72.414 29.86 76.788 ; 
        RECT 29.324 72.414 29.428 76.788 ; 
        RECT 28.892 72.414 28.996 76.788 ; 
        RECT 28.46 72.414 28.564 76.788 ; 
        RECT 28.028 72.414 28.132 76.788 ; 
        RECT 27.596 72.414 27.7 76.788 ; 
        RECT 27.164 72.414 27.268 76.788 ; 
        RECT 26.732 72.414 26.836 76.788 ; 
        RECT 26.3 72.414 26.404 76.788 ; 
        RECT 25.868 72.414 25.972 76.788 ; 
        RECT 25.436 72.414 25.54 76.788 ; 
        RECT 25.004 72.414 25.108 76.788 ; 
        RECT 24.572 72.414 24.676 76.788 ; 
        RECT 24.14 72.414 24.244 76.788 ; 
        RECT 23.708 72.414 23.812 76.788 ; 
        RECT 22.856 72.414 23.164 76.788 ; 
        RECT 15.284 72.414 15.592 76.788 ; 
        RECT 14.636 72.414 14.74 76.788 ; 
        RECT 14.204 72.414 14.308 76.788 ; 
        RECT 13.772 72.414 13.876 76.788 ; 
        RECT 13.34 72.414 13.444 76.788 ; 
        RECT 12.908 72.414 13.012 76.788 ; 
        RECT 12.476 72.414 12.58 76.788 ; 
        RECT 12.044 72.414 12.148 76.788 ; 
        RECT 11.612 72.414 11.716 76.788 ; 
        RECT 11.18 72.414 11.284 76.788 ; 
        RECT 10.748 72.414 10.852 76.788 ; 
        RECT 10.316 72.414 10.42 76.788 ; 
        RECT 9.884 72.414 9.988 76.788 ; 
        RECT 9.452 72.414 9.556 76.788 ; 
        RECT 9.02 72.414 9.124 76.788 ; 
        RECT 8.588 72.414 8.692 76.788 ; 
        RECT 8.156 72.414 8.26 76.788 ; 
        RECT 7.724 72.414 7.828 76.788 ; 
        RECT 7.292 72.414 7.396 76.788 ; 
        RECT 6.86 72.414 6.964 76.788 ; 
        RECT 6.428 72.414 6.532 76.788 ; 
        RECT 5.996 72.414 6.1 76.788 ; 
        RECT 5.564 72.414 5.668 76.788 ; 
        RECT 5.132 72.414 5.236 76.788 ; 
        RECT 4.7 72.414 4.804 76.788 ; 
        RECT 4.268 72.414 4.372 76.788 ; 
        RECT 3.836 72.414 3.94 76.788 ; 
        RECT 3.404 72.414 3.508 76.788 ; 
        RECT 2.972 72.414 3.076 76.788 ; 
        RECT 2.54 72.414 2.644 76.788 ; 
        RECT 2.108 72.414 2.212 76.788 ; 
        RECT 1.676 72.414 1.78 76.788 ; 
        RECT 1.244 72.414 1.348 76.788 ; 
        RECT 0.812 72.414 0.916 76.788 ; 
        RECT 0 72.414 0.34 76.788 ; 
        RECT 20.72 76.734 21.232 81.108 ; 
        RECT 20.664 79.396 21.232 80.686 ; 
        RECT 20.072 78.304 20.32 81.108 ; 
        RECT 20.016 79.542 20.32 80.156 ; 
        RECT 20.072 76.734 20.176 81.108 ; 
        RECT 20.072 77.218 20.232 78.176 ; 
        RECT 20.072 76.734 20.32 77.09 ; 
        RECT 18.884 78.536 19.708 81.108 ; 
        RECT 19.604 76.734 19.708 81.108 ; 
        RECT 18.884 79.644 19.764 80.676 ; 
        RECT 18.884 76.734 19.276 81.108 ; 
        RECT 17.216 76.734 17.548 81.108 ; 
        RECT 17.216 77.088 17.604 80.83 ; 
        RECT 38.108 76.734 38.448 81.108 ; 
        RECT 37.532 76.734 37.636 81.108 ; 
        RECT 37.1 76.734 37.204 81.108 ; 
        RECT 36.668 76.734 36.772 81.108 ; 
        RECT 36.236 76.734 36.34 81.108 ; 
        RECT 35.804 76.734 35.908 81.108 ; 
        RECT 35.372 76.734 35.476 81.108 ; 
        RECT 34.94 76.734 35.044 81.108 ; 
        RECT 34.508 76.734 34.612 81.108 ; 
        RECT 34.076 76.734 34.18 81.108 ; 
        RECT 33.644 76.734 33.748 81.108 ; 
        RECT 33.212 76.734 33.316 81.108 ; 
        RECT 32.78 76.734 32.884 81.108 ; 
        RECT 32.348 76.734 32.452 81.108 ; 
        RECT 31.916 76.734 32.02 81.108 ; 
        RECT 31.484 76.734 31.588 81.108 ; 
        RECT 31.052 76.734 31.156 81.108 ; 
        RECT 30.62 76.734 30.724 81.108 ; 
        RECT 30.188 76.734 30.292 81.108 ; 
        RECT 29.756 76.734 29.86 81.108 ; 
        RECT 29.324 76.734 29.428 81.108 ; 
        RECT 28.892 76.734 28.996 81.108 ; 
        RECT 28.46 76.734 28.564 81.108 ; 
        RECT 28.028 76.734 28.132 81.108 ; 
        RECT 27.596 76.734 27.7 81.108 ; 
        RECT 27.164 76.734 27.268 81.108 ; 
        RECT 26.732 76.734 26.836 81.108 ; 
        RECT 26.3 76.734 26.404 81.108 ; 
        RECT 25.868 76.734 25.972 81.108 ; 
        RECT 25.436 76.734 25.54 81.108 ; 
        RECT 25.004 76.734 25.108 81.108 ; 
        RECT 24.572 76.734 24.676 81.108 ; 
        RECT 24.14 76.734 24.244 81.108 ; 
        RECT 23.708 76.734 23.812 81.108 ; 
        RECT 22.856 76.734 23.164 81.108 ; 
        RECT 15.284 76.734 15.592 81.108 ; 
        RECT 14.636 76.734 14.74 81.108 ; 
        RECT 14.204 76.734 14.308 81.108 ; 
        RECT 13.772 76.734 13.876 81.108 ; 
        RECT 13.34 76.734 13.444 81.108 ; 
        RECT 12.908 76.734 13.012 81.108 ; 
        RECT 12.476 76.734 12.58 81.108 ; 
        RECT 12.044 76.734 12.148 81.108 ; 
        RECT 11.612 76.734 11.716 81.108 ; 
        RECT 11.18 76.734 11.284 81.108 ; 
        RECT 10.748 76.734 10.852 81.108 ; 
        RECT 10.316 76.734 10.42 81.108 ; 
        RECT 9.884 76.734 9.988 81.108 ; 
        RECT 9.452 76.734 9.556 81.108 ; 
        RECT 9.02 76.734 9.124 81.108 ; 
        RECT 8.588 76.734 8.692 81.108 ; 
        RECT 8.156 76.734 8.26 81.108 ; 
        RECT 7.724 76.734 7.828 81.108 ; 
        RECT 7.292 76.734 7.396 81.108 ; 
        RECT 6.86 76.734 6.964 81.108 ; 
        RECT 6.428 76.734 6.532 81.108 ; 
        RECT 5.996 76.734 6.1 81.108 ; 
        RECT 5.564 76.734 5.668 81.108 ; 
        RECT 5.132 76.734 5.236 81.108 ; 
        RECT 4.7 76.734 4.804 81.108 ; 
        RECT 4.268 76.734 4.372 81.108 ; 
        RECT 3.836 76.734 3.94 81.108 ; 
        RECT 3.404 76.734 3.508 81.108 ; 
        RECT 2.972 76.734 3.076 81.108 ; 
        RECT 2.54 76.734 2.644 81.108 ; 
        RECT 2.108 76.734 2.212 81.108 ; 
        RECT 1.676 76.734 1.78 81.108 ; 
        RECT 1.244 76.734 1.348 81.108 ; 
        RECT 0.812 76.734 0.916 81.108 ; 
        RECT 0 76.734 0.34 81.108 ; 
        RECT 20.72 81.054 21.232 85.428 ; 
        RECT 20.664 83.716 21.232 85.006 ; 
        RECT 20.072 82.624 20.32 85.428 ; 
        RECT 20.016 83.862 20.32 84.476 ; 
        RECT 20.072 81.054 20.176 85.428 ; 
        RECT 20.072 81.538 20.232 82.496 ; 
        RECT 20.072 81.054 20.32 81.41 ; 
        RECT 18.884 82.856 19.708 85.428 ; 
        RECT 19.604 81.054 19.708 85.428 ; 
        RECT 18.884 83.964 19.764 84.996 ; 
        RECT 18.884 81.054 19.276 85.428 ; 
        RECT 17.216 81.054 17.548 85.428 ; 
        RECT 17.216 81.408 17.604 85.15 ; 
        RECT 38.108 81.054 38.448 85.428 ; 
        RECT 37.532 81.054 37.636 85.428 ; 
        RECT 37.1 81.054 37.204 85.428 ; 
        RECT 36.668 81.054 36.772 85.428 ; 
        RECT 36.236 81.054 36.34 85.428 ; 
        RECT 35.804 81.054 35.908 85.428 ; 
        RECT 35.372 81.054 35.476 85.428 ; 
        RECT 34.94 81.054 35.044 85.428 ; 
        RECT 34.508 81.054 34.612 85.428 ; 
        RECT 34.076 81.054 34.18 85.428 ; 
        RECT 33.644 81.054 33.748 85.428 ; 
        RECT 33.212 81.054 33.316 85.428 ; 
        RECT 32.78 81.054 32.884 85.428 ; 
        RECT 32.348 81.054 32.452 85.428 ; 
        RECT 31.916 81.054 32.02 85.428 ; 
        RECT 31.484 81.054 31.588 85.428 ; 
        RECT 31.052 81.054 31.156 85.428 ; 
        RECT 30.62 81.054 30.724 85.428 ; 
        RECT 30.188 81.054 30.292 85.428 ; 
        RECT 29.756 81.054 29.86 85.428 ; 
        RECT 29.324 81.054 29.428 85.428 ; 
        RECT 28.892 81.054 28.996 85.428 ; 
        RECT 28.46 81.054 28.564 85.428 ; 
        RECT 28.028 81.054 28.132 85.428 ; 
        RECT 27.596 81.054 27.7 85.428 ; 
        RECT 27.164 81.054 27.268 85.428 ; 
        RECT 26.732 81.054 26.836 85.428 ; 
        RECT 26.3 81.054 26.404 85.428 ; 
        RECT 25.868 81.054 25.972 85.428 ; 
        RECT 25.436 81.054 25.54 85.428 ; 
        RECT 25.004 81.054 25.108 85.428 ; 
        RECT 24.572 81.054 24.676 85.428 ; 
        RECT 24.14 81.054 24.244 85.428 ; 
        RECT 23.708 81.054 23.812 85.428 ; 
        RECT 22.856 81.054 23.164 85.428 ; 
        RECT 15.284 81.054 15.592 85.428 ; 
        RECT 14.636 81.054 14.74 85.428 ; 
        RECT 14.204 81.054 14.308 85.428 ; 
        RECT 13.772 81.054 13.876 85.428 ; 
        RECT 13.34 81.054 13.444 85.428 ; 
        RECT 12.908 81.054 13.012 85.428 ; 
        RECT 12.476 81.054 12.58 85.428 ; 
        RECT 12.044 81.054 12.148 85.428 ; 
        RECT 11.612 81.054 11.716 85.428 ; 
        RECT 11.18 81.054 11.284 85.428 ; 
        RECT 10.748 81.054 10.852 85.428 ; 
        RECT 10.316 81.054 10.42 85.428 ; 
        RECT 9.884 81.054 9.988 85.428 ; 
        RECT 9.452 81.054 9.556 85.428 ; 
        RECT 9.02 81.054 9.124 85.428 ; 
        RECT 8.588 81.054 8.692 85.428 ; 
        RECT 8.156 81.054 8.26 85.428 ; 
        RECT 7.724 81.054 7.828 85.428 ; 
        RECT 7.292 81.054 7.396 85.428 ; 
        RECT 6.86 81.054 6.964 85.428 ; 
        RECT 6.428 81.054 6.532 85.428 ; 
        RECT 5.996 81.054 6.1 85.428 ; 
        RECT 5.564 81.054 5.668 85.428 ; 
        RECT 5.132 81.054 5.236 85.428 ; 
        RECT 4.7 81.054 4.804 85.428 ; 
        RECT 4.268 81.054 4.372 85.428 ; 
        RECT 3.836 81.054 3.94 85.428 ; 
        RECT 3.404 81.054 3.508 85.428 ; 
        RECT 2.972 81.054 3.076 85.428 ; 
        RECT 2.54 81.054 2.644 85.428 ; 
        RECT 2.108 81.054 2.212 85.428 ; 
        RECT 1.676 81.054 1.78 85.428 ; 
        RECT 1.244 81.054 1.348 85.428 ; 
        RECT 0.812 81.054 0.916 85.428 ; 
        RECT 0 81.054 0.34 85.428 ; 
        RECT 20.72 85.374 21.232 89.748 ; 
        RECT 20.664 88.036 21.232 89.326 ; 
        RECT 20.072 86.944 20.32 89.748 ; 
        RECT 20.016 88.182 20.32 88.796 ; 
        RECT 20.072 85.374 20.176 89.748 ; 
        RECT 20.072 85.858 20.232 86.816 ; 
        RECT 20.072 85.374 20.32 85.73 ; 
        RECT 18.884 87.176 19.708 89.748 ; 
        RECT 19.604 85.374 19.708 89.748 ; 
        RECT 18.884 88.284 19.764 89.316 ; 
        RECT 18.884 85.374 19.276 89.748 ; 
        RECT 17.216 85.374 17.548 89.748 ; 
        RECT 17.216 85.728 17.604 89.47 ; 
        RECT 38.108 85.374 38.448 89.748 ; 
        RECT 37.532 85.374 37.636 89.748 ; 
        RECT 37.1 85.374 37.204 89.748 ; 
        RECT 36.668 85.374 36.772 89.748 ; 
        RECT 36.236 85.374 36.34 89.748 ; 
        RECT 35.804 85.374 35.908 89.748 ; 
        RECT 35.372 85.374 35.476 89.748 ; 
        RECT 34.94 85.374 35.044 89.748 ; 
        RECT 34.508 85.374 34.612 89.748 ; 
        RECT 34.076 85.374 34.18 89.748 ; 
        RECT 33.644 85.374 33.748 89.748 ; 
        RECT 33.212 85.374 33.316 89.748 ; 
        RECT 32.78 85.374 32.884 89.748 ; 
        RECT 32.348 85.374 32.452 89.748 ; 
        RECT 31.916 85.374 32.02 89.748 ; 
        RECT 31.484 85.374 31.588 89.748 ; 
        RECT 31.052 85.374 31.156 89.748 ; 
        RECT 30.62 85.374 30.724 89.748 ; 
        RECT 30.188 85.374 30.292 89.748 ; 
        RECT 29.756 85.374 29.86 89.748 ; 
        RECT 29.324 85.374 29.428 89.748 ; 
        RECT 28.892 85.374 28.996 89.748 ; 
        RECT 28.46 85.374 28.564 89.748 ; 
        RECT 28.028 85.374 28.132 89.748 ; 
        RECT 27.596 85.374 27.7 89.748 ; 
        RECT 27.164 85.374 27.268 89.748 ; 
        RECT 26.732 85.374 26.836 89.748 ; 
        RECT 26.3 85.374 26.404 89.748 ; 
        RECT 25.868 85.374 25.972 89.748 ; 
        RECT 25.436 85.374 25.54 89.748 ; 
        RECT 25.004 85.374 25.108 89.748 ; 
        RECT 24.572 85.374 24.676 89.748 ; 
        RECT 24.14 85.374 24.244 89.748 ; 
        RECT 23.708 85.374 23.812 89.748 ; 
        RECT 22.856 85.374 23.164 89.748 ; 
        RECT 15.284 85.374 15.592 89.748 ; 
        RECT 14.636 85.374 14.74 89.748 ; 
        RECT 14.204 85.374 14.308 89.748 ; 
        RECT 13.772 85.374 13.876 89.748 ; 
        RECT 13.34 85.374 13.444 89.748 ; 
        RECT 12.908 85.374 13.012 89.748 ; 
        RECT 12.476 85.374 12.58 89.748 ; 
        RECT 12.044 85.374 12.148 89.748 ; 
        RECT 11.612 85.374 11.716 89.748 ; 
        RECT 11.18 85.374 11.284 89.748 ; 
        RECT 10.748 85.374 10.852 89.748 ; 
        RECT 10.316 85.374 10.42 89.748 ; 
        RECT 9.884 85.374 9.988 89.748 ; 
        RECT 9.452 85.374 9.556 89.748 ; 
        RECT 9.02 85.374 9.124 89.748 ; 
        RECT 8.588 85.374 8.692 89.748 ; 
        RECT 8.156 85.374 8.26 89.748 ; 
        RECT 7.724 85.374 7.828 89.748 ; 
        RECT 7.292 85.374 7.396 89.748 ; 
        RECT 6.86 85.374 6.964 89.748 ; 
        RECT 6.428 85.374 6.532 89.748 ; 
        RECT 5.996 85.374 6.1 89.748 ; 
        RECT 5.564 85.374 5.668 89.748 ; 
        RECT 5.132 85.374 5.236 89.748 ; 
        RECT 4.7 85.374 4.804 89.748 ; 
        RECT 4.268 85.374 4.372 89.748 ; 
        RECT 3.836 85.374 3.94 89.748 ; 
        RECT 3.404 85.374 3.508 89.748 ; 
        RECT 2.972 85.374 3.076 89.748 ; 
        RECT 2.54 85.374 2.644 89.748 ; 
        RECT 2.108 85.374 2.212 89.748 ; 
        RECT 1.676 85.374 1.78 89.748 ; 
        RECT 1.244 85.374 1.348 89.748 ; 
        RECT 0.812 85.374 0.916 89.748 ; 
        RECT 0 85.374 0.34 89.748 ; 
        RECT 20.72 89.694 21.232 94.068 ; 
        RECT 20.664 92.356 21.232 93.646 ; 
        RECT 20.072 91.264 20.32 94.068 ; 
        RECT 20.016 92.502 20.32 93.116 ; 
        RECT 20.072 89.694 20.176 94.068 ; 
        RECT 20.072 90.178 20.232 91.136 ; 
        RECT 20.072 89.694 20.32 90.05 ; 
        RECT 18.884 91.496 19.708 94.068 ; 
        RECT 19.604 89.694 19.708 94.068 ; 
        RECT 18.884 92.604 19.764 93.636 ; 
        RECT 18.884 89.694 19.276 94.068 ; 
        RECT 17.216 89.694 17.548 94.068 ; 
        RECT 17.216 90.048 17.604 93.79 ; 
        RECT 38.108 89.694 38.448 94.068 ; 
        RECT 37.532 89.694 37.636 94.068 ; 
        RECT 37.1 89.694 37.204 94.068 ; 
        RECT 36.668 89.694 36.772 94.068 ; 
        RECT 36.236 89.694 36.34 94.068 ; 
        RECT 35.804 89.694 35.908 94.068 ; 
        RECT 35.372 89.694 35.476 94.068 ; 
        RECT 34.94 89.694 35.044 94.068 ; 
        RECT 34.508 89.694 34.612 94.068 ; 
        RECT 34.076 89.694 34.18 94.068 ; 
        RECT 33.644 89.694 33.748 94.068 ; 
        RECT 33.212 89.694 33.316 94.068 ; 
        RECT 32.78 89.694 32.884 94.068 ; 
        RECT 32.348 89.694 32.452 94.068 ; 
        RECT 31.916 89.694 32.02 94.068 ; 
        RECT 31.484 89.694 31.588 94.068 ; 
        RECT 31.052 89.694 31.156 94.068 ; 
        RECT 30.62 89.694 30.724 94.068 ; 
        RECT 30.188 89.694 30.292 94.068 ; 
        RECT 29.756 89.694 29.86 94.068 ; 
        RECT 29.324 89.694 29.428 94.068 ; 
        RECT 28.892 89.694 28.996 94.068 ; 
        RECT 28.46 89.694 28.564 94.068 ; 
        RECT 28.028 89.694 28.132 94.068 ; 
        RECT 27.596 89.694 27.7 94.068 ; 
        RECT 27.164 89.694 27.268 94.068 ; 
        RECT 26.732 89.694 26.836 94.068 ; 
        RECT 26.3 89.694 26.404 94.068 ; 
        RECT 25.868 89.694 25.972 94.068 ; 
        RECT 25.436 89.694 25.54 94.068 ; 
        RECT 25.004 89.694 25.108 94.068 ; 
        RECT 24.572 89.694 24.676 94.068 ; 
        RECT 24.14 89.694 24.244 94.068 ; 
        RECT 23.708 89.694 23.812 94.068 ; 
        RECT 22.856 89.694 23.164 94.068 ; 
        RECT 15.284 89.694 15.592 94.068 ; 
        RECT 14.636 89.694 14.74 94.068 ; 
        RECT 14.204 89.694 14.308 94.068 ; 
        RECT 13.772 89.694 13.876 94.068 ; 
        RECT 13.34 89.694 13.444 94.068 ; 
        RECT 12.908 89.694 13.012 94.068 ; 
        RECT 12.476 89.694 12.58 94.068 ; 
        RECT 12.044 89.694 12.148 94.068 ; 
        RECT 11.612 89.694 11.716 94.068 ; 
        RECT 11.18 89.694 11.284 94.068 ; 
        RECT 10.748 89.694 10.852 94.068 ; 
        RECT 10.316 89.694 10.42 94.068 ; 
        RECT 9.884 89.694 9.988 94.068 ; 
        RECT 9.452 89.694 9.556 94.068 ; 
        RECT 9.02 89.694 9.124 94.068 ; 
        RECT 8.588 89.694 8.692 94.068 ; 
        RECT 8.156 89.694 8.26 94.068 ; 
        RECT 7.724 89.694 7.828 94.068 ; 
        RECT 7.292 89.694 7.396 94.068 ; 
        RECT 6.86 89.694 6.964 94.068 ; 
        RECT 6.428 89.694 6.532 94.068 ; 
        RECT 5.996 89.694 6.1 94.068 ; 
        RECT 5.564 89.694 5.668 94.068 ; 
        RECT 5.132 89.694 5.236 94.068 ; 
        RECT 4.7 89.694 4.804 94.068 ; 
        RECT 4.268 89.694 4.372 94.068 ; 
        RECT 3.836 89.694 3.94 94.068 ; 
        RECT 3.404 89.694 3.508 94.068 ; 
        RECT 2.972 89.694 3.076 94.068 ; 
        RECT 2.54 89.694 2.644 94.068 ; 
        RECT 2.108 89.694 2.212 94.068 ; 
        RECT 1.676 89.694 1.78 94.068 ; 
        RECT 1.244 89.694 1.348 94.068 ; 
        RECT 0.812 89.694 0.916 94.068 ; 
        RECT 0 89.694 0.34 94.068 ; 
        RECT 20.72 94.014 21.232 98.388 ; 
        RECT 20.664 96.676 21.232 97.966 ; 
        RECT 20.072 95.584 20.32 98.388 ; 
        RECT 20.016 96.822 20.32 97.436 ; 
        RECT 20.072 94.014 20.176 98.388 ; 
        RECT 20.072 94.498 20.232 95.456 ; 
        RECT 20.072 94.014 20.32 94.37 ; 
        RECT 18.884 95.816 19.708 98.388 ; 
        RECT 19.604 94.014 19.708 98.388 ; 
        RECT 18.884 96.924 19.764 97.956 ; 
        RECT 18.884 94.014 19.276 98.388 ; 
        RECT 17.216 94.014 17.548 98.388 ; 
        RECT 17.216 94.368 17.604 98.11 ; 
        RECT 38.108 94.014 38.448 98.388 ; 
        RECT 37.532 94.014 37.636 98.388 ; 
        RECT 37.1 94.014 37.204 98.388 ; 
        RECT 36.668 94.014 36.772 98.388 ; 
        RECT 36.236 94.014 36.34 98.388 ; 
        RECT 35.804 94.014 35.908 98.388 ; 
        RECT 35.372 94.014 35.476 98.388 ; 
        RECT 34.94 94.014 35.044 98.388 ; 
        RECT 34.508 94.014 34.612 98.388 ; 
        RECT 34.076 94.014 34.18 98.388 ; 
        RECT 33.644 94.014 33.748 98.388 ; 
        RECT 33.212 94.014 33.316 98.388 ; 
        RECT 32.78 94.014 32.884 98.388 ; 
        RECT 32.348 94.014 32.452 98.388 ; 
        RECT 31.916 94.014 32.02 98.388 ; 
        RECT 31.484 94.014 31.588 98.388 ; 
        RECT 31.052 94.014 31.156 98.388 ; 
        RECT 30.62 94.014 30.724 98.388 ; 
        RECT 30.188 94.014 30.292 98.388 ; 
        RECT 29.756 94.014 29.86 98.388 ; 
        RECT 29.324 94.014 29.428 98.388 ; 
        RECT 28.892 94.014 28.996 98.388 ; 
        RECT 28.46 94.014 28.564 98.388 ; 
        RECT 28.028 94.014 28.132 98.388 ; 
        RECT 27.596 94.014 27.7 98.388 ; 
        RECT 27.164 94.014 27.268 98.388 ; 
        RECT 26.732 94.014 26.836 98.388 ; 
        RECT 26.3 94.014 26.404 98.388 ; 
        RECT 25.868 94.014 25.972 98.388 ; 
        RECT 25.436 94.014 25.54 98.388 ; 
        RECT 25.004 94.014 25.108 98.388 ; 
        RECT 24.572 94.014 24.676 98.388 ; 
        RECT 24.14 94.014 24.244 98.388 ; 
        RECT 23.708 94.014 23.812 98.388 ; 
        RECT 22.856 94.014 23.164 98.388 ; 
        RECT 15.284 94.014 15.592 98.388 ; 
        RECT 14.636 94.014 14.74 98.388 ; 
        RECT 14.204 94.014 14.308 98.388 ; 
        RECT 13.772 94.014 13.876 98.388 ; 
        RECT 13.34 94.014 13.444 98.388 ; 
        RECT 12.908 94.014 13.012 98.388 ; 
        RECT 12.476 94.014 12.58 98.388 ; 
        RECT 12.044 94.014 12.148 98.388 ; 
        RECT 11.612 94.014 11.716 98.388 ; 
        RECT 11.18 94.014 11.284 98.388 ; 
        RECT 10.748 94.014 10.852 98.388 ; 
        RECT 10.316 94.014 10.42 98.388 ; 
        RECT 9.884 94.014 9.988 98.388 ; 
        RECT 9.452 94.014 9.556 98.388 ; 
        RECT 9.02 94.014 9.124 98.388 ; 
        RECT 8.588 94.014 8.692 98.388 ; 
        RECT 8.156 94.014 8.26 98.388 ; 
        RECT 7.724 94.014 7.828 98.388 ; 
        RECT 7.292 94.014 7.396 98.388 ; 
        RECT 6.86 94.014 6.964 98.388 ; 
        RECT 6.428 94.014 6.532 98.388 ; 
        RECT 5.996 94.014 6.1 98.388 ; 
        RECT 5.564 94.014 5.668 98.388 ; 
        RECT 5.132 94.014 5.236 98.388 ; 
        RECT 4.7 94.014 4.804 98.388 ; 
        RECT 4.268 94.014 4.372 98.388 ; 
        RECT 3.836 94.014 3.94 98.388 ; 
        RECT 3.404 94.014 3.508 98.388 ; 
        RECT 2.972 94.014 3.076 98.388 ; 
        RECT 2.54 94.014 2.644 98.388 ; 
        RECT 2.108 94.014 2.212 98.388 ; 
        RECT 1.676 94.014 1.78 98.388 ; 
        RECT 1.244 94.014 1.348 98.388 ; 
        RECT 0.812 94.014 0.916 98.388 ; 
        RECT 0 94.014 0.34 98.388 ; 
        RECT 20.72 98.334 21.232 102.708 ; 
        RECT 20.664 100.996 21.232 102.286 ; 
        RECT 20.072 99.904 20.32 102.708 ; 
        RECT 20.016 101.142 20.32 101.756 ; 
        RECT 20.072 98.334 20.176 102.708 ; 
        RECT 20.072 98.818 20.232 99.776 ; 
        RECT 20.072 98.334 20.32 98.69 ; 
        RECT 18.884 100.136 19.708 102.708 ; 
        RECT 19.604 98.334 19.708 102.708 ; 
        RECT 18.884 101.244 19.764 102.276 ; 
        RECT 18.884 98.334 19.276 102.708 ; 
        RECT 17.216 98.334 17.548 102.708 ; 
        RECT 17.216 98.688 17.604 102.43 ; 
        RECT 38.108 98.334 38.448 102.708 ; 
        RECT 37.532 98.334 37.636 102.708 ; 
        RECT 37.1 98.334 37.204 102.708 ; 
        RECT 36.668 98.334 36.772 102.708 ; 
        RECT 36.236 98.334 36.34 102.708 ; 
        RECT 35.804 98.334 35.908 102.708 ; 
        RECT 35.372 98.334 35.476 102.708 ; 
        RECT 34.94 98.334 35.044 102.708 ; 
        RECT 34.508 98.334 34.612 102.708 ; 
        RECT 34.076 98.334 34.18 102.708 ; 
        RECT 33.644 98.334 33.748 102.708 ; 
        RECT 33.212 98.334 33.316 102.708 ; 
        RECT 32.78 98.334 32.884 102.708 ; 
        RECT 32.348 98.334 32.452 102.708 ; 
        RECT 31.916 98.334 32.02 102.708 ; 
        RECT 31.484 98.334 31.588 102.708 ; 
        RECT 31.052 98.334 31.156 102.708 ; 
        RECT 30.62 98.334 30.724 102.708 ; 
        RECT 30.188 98.334 30.292 102.708 ; 
        RECT 29.756 98.334 29.86 102.708 ; 
        RECT 29.324 98.334 29.428 102.708 ; 
        RECT 28.892 98.334 28.996 102.708 ; 
        RECT 28.46 98.334 28.564 102.708 ; 
        RECT 28.028 98.334 28.132 102.708 ; 
        RECT 27.596 98.334 27.7 102.708 ; 
        RECT 27.164 98.334 27.268 102.708 ; 
        RECT 26.732 98.334 26.836 102.708 ; 
        RECT 26.3 98.334 26.404 102.708 ; 
        RECT 25.868 98.334 25.972 102.708 ; 
        RECT 25.436 98.334 25.54 102.708 ; 
        RECT 25.004 98.334 25.108 102.708 ; 
        RECT 24.572 98.334 24.676 102.708 ; 
        RECT 24.14 98.334 24.244 102.708 ; 
        RECT 23.708 98.334 23.812 102.708 ; 
        RECT 22.856 98.334 23.164 102.708 ; 
        RECT 15.284 98.334 15.592 102.708 ; 
        RECT 14.636 98.334 14.74 102.708 ; 
        RECT 14.204 98.334 14.308 102.708 ; 
        RECT 13.772 98.334 13.876 102.708 ; 
        RECT 13.34 98.334 13.444 102.708 ; 
        RECT 12.908 98.334 13.012 102.708 ; 
        RECT 12.476 98.334 12.58 102.708 ; 
        RECT 12.044 98.334 12.148 102.708 ; 
        RECT 11.612 98.334 11.716 102.708 ; 
        RECT 11.18 98.334 11.284 102.708 ; 
        RECT 10.748 98.334 10.852 102.708 ; 
        RECT 10.316 98.334 10.42 102.708 ; 
        RECT 9.884 98.334 9.988 102.708 ; 
        RECT 9.452 98.334 9.556 102.708 ; 
        RECT 9.02 98.334 9.124 102.708 ; 
        RECT 8.588 98.334 8.692 102.708 ; 
        RECT 8.156 98.334 8.26 102.708 ; 
        RECT 7.724 98.334 7.828 102.708 ; 
        RECT 7.292 98.334 7.396 102.708 ; 
        RECT 6.86 98.334 6.964 102.708 ; 
        RECT 6.428 98.334 6.532 102.708 ; 
        RECT 5.996 98.334 6.1 102.708 ; 
        RECT 5.564 98.334 5.668 102.708 ; 
        RECT 5.132 98.334 5.236 102.708 ; 
        RECT 4.7 98.334 4.804 102.708 ; 
        RECT 4.268 98.334 4.372 102.708 ; 
        RECT 3.836 98.334 3.94 102.708 ; 
        RECT 3.404 98.334 3.508 102.708 ; 
        RECT 2.972 98.334 3.076 102.708 ; 
        RECT 2.54 98.334 2.644 102.708 ; 
        RECT 2.108 98.334 2.212 102.708 ; 
        RECT 1.676 98.334 1.78 102.708 ; 
        RECT 1.244 98.334 1.348 102.708 ; 
        RECT 0.812 98.334 0.916 102.708 ; 
        RECT 0 98.334 0.34 102.708 ; 
        RECT 20.72 102.654 21.232 107.028 ; 
        RECT 20.664 105.316 21.232 106.606 ; 
        RECT 20.072 104.224 20.32 107.028 ; 
        RECT 20.016 105.462 20.32 106.076 ; 
        RECT 20.072 102.654 20.176 107.028 ; 
        RECT 20.072 103.138 20.232 104.096 ; 
        RECT 20.072 102.654 20.32 103.01 ; 
        RECT 18.884 104.456 19.708 107.028 ; 
        RECT 19.604 102.654 19.708 107.028 ; 
        RECT 18.884 105.564 19.764 106.596 ; 
        RECT 18.884 102.654 19.276 107.028 ; 
        RECT 17.216 102.654 17.548 107.028 ; 
        RECT 17.216 103.008 17.604 106.75 ; 
        RECT 38.108 102.654 38.448 107.028 ; 
        RECT 37.532 102.654 37.636 107.028 ; 
        RECT 37.1 102.654 37.204 107.028 ; 
        RECT 36.668 102.654 36.772 107.028 ; 
        RECT 36.236 102.654 36.34 107.028 ; 
        RECT 35.804 102.654 35.908 107.028 ; 
        RECT 35.372 102.654 35.476 107.028 ; 
        RECT 34.94 102.654 35.044 107.028 ; 
        RECT 34.508 102.654 34.612 107.028 ; 
        RECT 34.076 102.654 34.18 107.028 ; 
        RECT 33.644 102.654 33.748 107.028 ; 
        RECT 33.212 102.654 33.316 107.028 ; 
        RECT 32.78 102.654 32.884 107.028 ; 
        RECT 32.348 102.654 32.452 107.028 ; 
        RECT 31.916 102.654 32.02 107.028 ; 
        RECT 31.484 102.654 31.588 107.028 ; 
        RECT 31.052 102.654 31.156 107.028 ; 
        RECT 30.62 102.654 30.724 107.028 ; 
        RECT 30.188 102.654 30.292 107.028 ; 
        RECT 29.756 102.654 29.86 107.028 ; 
        RECT 29.324 102.654 29.428 107.028 ; 
        RECT 28.892 102.654 28.996 107.028 ; 
        RECT 28.46 102.654 28.564 107.028 ; 
        RECT 28.028 102.654 28.132 107.028 ; 
        RECT 27.596 102.654 27.7 107.028 ; 
        RECT 27.164 102.654 27.268 107.028 ; 
        RECT 26.732 102.654 26.836 107.028 ; 
        RECT 26.3 102.654 26.404 107.028 ; 
        RECT 25.868 102.654 25.972 107.028 ; 
        RECT 25.436 102.654 25.54 107.028 ; 
        RECT 25.004 102.654 25.108 107.028 ; 
        RECT 24.572 102.654 24.676 107.028 ; 
        RECT 24.14 102.654 24.244 107.028 ; 
        RECT 23.708 102.654 23.812 107.028 ; 
        RECT 22.856 102.654 23.164 107.028 ; 
        RECT 15.284 102.654 15.592 107.028 ; 
        RECT 14.636 102.654 14.74 107.028 ; 
        RECT 14.204 102.654 14.308 107.028 ; 
        RECT 13.772 102.654 13.876 107.028 ; 
        RECT 13.34 102.654 13.444 107.028 ; 
        RECT 12.908 102.654 13.012 107.028 ; 
        RECT 12.476 102.654 12.58 107.028 ; 
        RECT 12.044 102.654 12.148 107.028 ; 
        RECT 11.612 102.654 11.716 107.028 ; 
        RECT 11.18 102.654 11.284 107.028 ; 
        RECT 10.748 102.654 10.852 107.028 ; 
        RECT 10.316 102.654 10.42 107.028 ; 
        RECT 9.884 102.654 9.988 107.028 ; 
        RECT 9.452 102.654 9.556 107.028 ; 
        RECT 9.02 102.654 9.124 107.028 ; 
        RECT 8.588 102.654 8.692 107.028 ; 
        RECT 8.156 102.654 8.26 107.028 ; 
        RECT 7.724 102.654 7.828 107.028 ; 
        RECT 7.292 102.654 7.396 107.028 ; 
        RECT 6.86 102.654 6.964 107.028 ; 
        RECT 6.428 102.654 6.532 107.028 ; 
        RECT 5.996 102.654 6.1 107.028 ; 
        RECT 5.564 102.654 5.668 107.028 ; 
        RECT 5.132 102.654 5.236 107.028 ; 
        RECT 4.7 102.654 4.804 107.028 ; 
        RECT 4.268 102.654 4.372 107.028 ; 
        RECT 3.836 102.654 3.94 107.028 ; 
        RECT 3.404 102.654 3.508 107.028 ; 
        RECT 2.972 102.654 3.076 107.028 ; 
        RECT 2.54 102.654 2.644 107.028 ; 
        RECT 2.108 102.654 2.212 107.028 ; 
        RECT 1.676 102.654 1.78 107.028 ; 
        RECT 1.244 102.654 1.348 107.028 ; 
        RECT 0.812 102.654 0.916 107.028 ; 
        RECT 0 102.654 0.34 107.028 ; 
        RECT 20.72 106.974 21.232 111.348 ; 
        RECT 20.664 109.636 21.232 110.926 ; 
        RECT 20.072 108.544 20.32 111.348 ; 
        RECT 20.016 109.782 20.32 110.396 ; 
        RECT 20.072 106.974 20.176 111.348 ; 
        RECT 20.072 107.458 20.232 108.416 ; 
        RECT 20.072 106.974 20.32 107.33 ; 
        RECT 18.884 108.776 19.708 111.348 ; 
        RECT 19.604 106.974 19.708 111.348 ; 
        RECT 18.884 109.884 19.764 110.916 ; 
        RECT 18.884 106.974 19.276 111.348 ; 
        RECT 17.216 106.974 17.548 111.348 ; 
        RECT 17.216 107.328 17.604 111.07 ; 
        RECT 38.108 106.974 38.448 111.348 ; 
        RECT 37.532 106.974 37.636 111.348 ; 
        RECT 37.1 106.974 37.204 111.348 ; 
        RECT 36.668 106.974 36.772 111.348 ; 
        RECT 36.236 106.974 36.34 111.348 ; 
        RECT 35.804 106.974 35.908 111.348 ; 
        RECT 35.372 106.974 35.476 111.348 ; 
        RECT 34.94 106.974 35.044 111.348 ; 
        RECT 34.508 106.974 34.612 111.348 ; 
        RECT 34.076 106.974 34.18 111.348 ; 
        RECT 33.644 106.974 33.748 111.348 ; 
        RECT 33.212 106.974 33.316 111.348 ; 
        RECT 32.78 106.974 32.884 111.348 ; 
        RECT 32.348 106.974 32.452 111.348 ; 
        RECT 31.916 106.974 32.02 111.348 ; 
        RECT 31.484 106.974 31.588 111.348 ; 
        RECT 31.052 106.974 31.156 111.348 ; 
        RECT 30.62 106.974 30.724 111.348 ; 
        RECT 30.188 106.974 30.292 111.348 ; 
        RECT 29.756 106.974 29.86 111.348 ; 
        RECT 29.324 106.974 29.428 111.348 ; 
        RECT 28.892 106.974 28.996 111.348 ; 
        RECT 28.46 106.974 28.564 111.348 ; 
        RECT 28.028 106.974 28.132 111.348 ; 
        RECT 27.596 106.974 27.7 111.348 ; 
        RECT 27.164 106.974 27.268 111.348 ; 
        RECT 26.732 106.974 26.836 111.348 ; 
        RECT 26.3 106.974 26.404 111.348 ; 
        RECT 25.868 106.974 25.972 111.348 ; 
        RECT 25.436 106.974 25.54 111.348 ; 
        RECT 25.004 106.974 25.108 111.348 ; 
        RECT 24.572 106.974 24.676 111.348 ; 
        RECT 24.14 106.974 24.244 111.348 ; 
        RECT 23.708 106.974 23.812 111.348 ; 
        RECT 22.856 106.974 23.164 111.348 ; 
        RECT 15.284 106.974 15.592 111.348 ; 
        RECT 14.636 106.974 14.74 111.348 ; 
        RECT 14.204 106.974 14.308 111.348 ; 
        RECT 13.772 106.974 13.876 111.348 ; 
        RECT 13.34 106.974 13.444 111.348 ; 
        RECT 12.908 106.974 13.012 111.348 ; 
        RECT 12.476 106.974 12.58 111.348 ; 
        RECT 12.044 106.974 12.148 111.348 ; 
        RECT 11.612 106.974 11.716 111.348 ; 
        RECT 11.18 106.974 11.284 111.348 ; 
        RECT 10.748 106.974 10.852 111.348 ; 
        RECT 10.316 106.974 10.42 111.348 ; 
        RECT 9.884 106.974 9.988 111.348 ; 
        RECT 9.452 106.974 9.556 111.348 ; 
        RECT 9.02 106.974 9.124 111.348 ; 
        RECT 8.588 106.974 8.692 111.348 ; 
        RECT 8.156 106.974 8.26 111.348 ; 
        RECT 7.724 106.974 7.828 111.348 ; 
        RECT 7.292 106.974 7.396 111.348 ; 
        RECT 6.86 106.974 6.964 111.348 ; 
        RECT 6.428 106.974 6.532 111.348 ; 
        RECT 5.996 106.974 6.1 111.348 ; 
        RECT 5.564 106.974 5.668 111.348 ; 
        RECT 5.132 106.974 5.236 111.348 ; 
        RECT 4.7 106.974 4.804 111.348 ; 
        RECT 4.268 106.974 4.372 111.348 ; 
        RECT 3.836 106.974 3.94 111.348 ; 
        RECT 3.404 106.974 3.508 111.348 ; 
        RECT 2.972 106.974 3.076 111.348 ; 
        RECT 2.54 106.974 2.644 111.348 ; 
        RECT 2.108 106.974 2.212 111.348 ; 
        RECT 1.676 106.974 1.78 111.348 ; 
        RECT 1.244 106.974 1.348 111.348 ; 
        RECT 0.812 106.974 0.916 111.348 ; 
        RECT 0 106.974 0.34 111.348 ; 
  LAYER V3 ; 
      RECT 0 4.88 38.448 5.4 ; 
      RECT 37.98 1.026 38.448 5.4 ; 
      RECT 23.364 4.496 37.908 5.4 ; 
      RECT 18.036 4.496 23.292 5.4 ; 
      RECT 15.156 1.026 17.676 5.4 ; 
      RECT 0.54 4.496 15.084 5.4 ; 
      RECT 0 1.026 0.468 5.4 ; 
      RECT 37.836 1.026 38.448 4.688 ; 
      RECT 23.58 1.026 37.764 5.4 ; 
      RECT 20.592 1.026 23.508 4.688 ; 
      RECT 19.944 1.808 20.448 5.4 ; 
      RECT 14.94 1.424 19.836 4.688 ; 
      RECT 0.684 1.026 14.868 5.4 ; 
      RECT 0 1.026 0.612 4.688 ; 
      RECT 20.376 1.026 38.448 4.304 ; 
      RECT 0 1.424 20.304 4.304 ; 
      RECT 19.476 1.026 38.448 1.712 ; 
      RECT 0 1.026 19.404 4.304 ; 
      RECT 0 1.026 38.448 1.328 ; 
      RECT 0 9.2 38.448 9.72 ; 
      RECT 37.98 5.346 38.448 9.72 ; 
      RECT 23.364 8.816 37.908 9.72 ; 
      RECT 18.036 8.816 23.292 9.72 ; 
      RECT 15.156 5.346 17.676 9.72 ; 
      RECT 0.54 8.816 15.084 9.72 ; 
      RECT 0 5.346 0.468 9.72 ; 
      RECT 37.836 5.346 38.448 9.008 ; 
      RECT 23.58 5.346 37.764 9.72 ; 
      RECT 20.592 5.346 23.508 9.008 ; 
      RECT 19.944 6.128 20.448 9.72 ; 
      RECT 14.94 5.744 19.836 9.008 ; 
      RECT 0.684 5.346 14.868 9.72 ; 
      RECT 0 5.346 0.612 9.008 ; 
      RECT 20.376 5.346 38.448 8.624 ; 
      RECT 0 5.744 20.304 8.624 ; 
      RECT 19.476 5.346 38.448 6.032 ; 
      RECT 0 5.346 19.404 8.624 ; 
      RECT 0 5.346 38.448 5.648 ; 
      RECT 0 13.52 38.448 14.04 ; 
      RECT 37.98 9.666 38.448 14.04 ; 
      RECT 23.364 13.136 37.908 14.04 ; 
      RECT 18.036 13.136 23.292 14.04 ; 
      RECT 15.156 9.666 17.676 14.04 ; 
      RECT 0.54 13.136 15.084 14.04 ; 
      RECT 0 9.666 0.468 14.04 ; 
      RECT 37.836 9.666 38.448 13.328 ; 
      RECT 23.58 9.666 37.764 14.04 ; 
      RECT 20.592 9.666 23.508 13.328 ; 
      RECT 19.944 10.448 20.448 14.04 ; 
      RECT 14.94 10.064 19.836 13.328 ; 
      RECT 0.684 9.666 14.868 14.04 ; 
      RECT 0 9.666 0.612 13.328 ; 
      RECT 20.376 9.666 38.448 12.944 ; 
      RECT 0 10.064 20.304 12.944 ; 
      RECT 19.476 9.666 38.448 10.352 ; 
      RECT 0 9.666 19.404 12.944 ; 
      RECT 0 9.666 38.448 9.968 ; 
      RECT 0 17.84 38.448 18.36 ; 
      RECT 37.98 13.986 38.448 18.36 ; 
      RECT 23.364 17.456 37.908 18.36 ; 
      RECT 18.036 17.456 23.292 18.36 ; 
      RECT 15.156 13.986 17.676 18.36 ; 
      RECT 0.54 17.456 15.084 18.36 ; 
      RECT 0 13.986 0.468 18.36 ; 
      RECT 37.836 13.986 38.448 17.648 ; 
      RECT 23.58 13.986 37.764 18.36 ; 
      RECT 20.592 13.986 23.508 17.648 ; 
      RECT 19.944 14.768 20.448 18.36 ; 
      RECT 14.94 14.384 19.836 17.648 ; 
      RECT 0.684 13.986 14.868 18.36 ; 
      RECT 0 13.986 0.612 17.648 ; 
      RECT 20.376 13.986 38.448 17.264 ; 
      RECT 0 14.384 20.304 17.264 ; 
      RECT 19.476 13.986 38.448 14.672 ; 
      RECT 0 13.986 19.404 17.264 ; 
      RECT 0 13.986 38.448 14.288 ; 
      RECT 0 22.16 38.448 22.68 ; 
      RECT 37.98 18.306 38.448 22.68 ; 
      RECT 23.364 21.776 37.908 22.68 ; 
      RECT 18.036 21.776 23.292 22.68 ; 
      RECT 15.156 18.306 17.676 22.68 ; 
      RECT 0.54 21.776 15.084 22.68 ; 
      RECT 0 18.306 0.468 22.68 ; 
      RECT 37.836 18.306 38.448 21.968 ; 
      RECT 23.58 18.306 37.764 22.68 ; 
      RECT 20.592 18.306 23.508 21.968 ; 
      RECT 19.944 19.088 20.448 22.68 ; 
      RECT 14.94 18.704 19.836 21.968 ; 
      RECT 0.684 18.306 14.868 22.68 ; 
      RECT 0 18.306 0.612 21.968 ; 
      RECT 20.376 18.306 38.448 21.584 ; 
      RECT 0 18.704 20.304 21.584 ; 
      RECT 19.476 18.306 38.448 18.992 ; 
      RECT 0 18.306 19.404 21.584 ; 
      RECT 0 18.306 38.448 18.608 ; 
      RECT 0 26.48 38.448 27 ; 
      RECT 37.98 22.626 38.448 27 ; 
      RECT 23.364 26.096 37.908 27 ; 
      RECT 18.036 26.096 23.292 27 ; 
      RECT 15.156 22.626 17.676 27 ; 
      RECT 0.54 26.096 15.084 27 ; 
      RECT 0 22.626 0.468 27 ; 
      RECT 37.836 22.626 38.448 26.288 ; 
      RECT 23.58 22.626 37.764 27 ; 
      RECT 20.592 22.626 23.508 26.288 ; 
      RECT 19.944 23.408 20.448 27 ; 
      RECT 14.94 23.024 19.836 26.288 ; 
      RECT 0.684 22.626 14.868 27 ; 
      RECT 0 22.626 0.612 26.288 ; 
      RECT 20.376 22.626 38.448 25.904 ; 
      RECT 0 23.024 20.304 25.904 ; 
      RECT 19.476 22.626 38.448 23.312 ; 
      RECT 0 22.626 19.404 25.904 ; 
      RECT 0 22.626 38.448 22.928 ; 
      RECT 0 30.8 38.448 31.32 ; 
      RECT 37.98 26.946 38.448 31.32 ; 
      RECT 23.364 30.416 37.908 31.32 ; 
      RECT 18.036 30.416 23.292 31.32 ; 
      RECT 15.156 26.946 17.676 31.32 ; 
      RECT 0.54 30.416 15.084 31.32 ; 
      RECT 0 26.946 0.468 31.32 ; 
      RECT 37.836 26.946 38.448 30.608 ; 
      RECT 23.58 26.946 37.764 31.32 ; 
      RECT 20.592 26.946 23.508 30.608 ; 
      RECT 19.944 27.728 20.448 31.32 ; 
      RECT 14.94 27.344 19.836 30.608 ; 
      RECT 0.684 26.946 14.868 31.32 ; 
      RECT 0 26.946 0.612 30.608 ; 
      RECT 20.376 26.946 38.448 30.224 ; 
      RECT 0 27.344 20.304 30.224 ; 
      RECT 19.476 26.946 38.448 27.632 ; 
      RECT 0 26.946 19.404 30.224 ; 
      RECT 0 26.946 38.448 27.248 ; 
      RECT 0 35.12 38.448 35.64 ; 
      RECT 37.98 31.266 38.448 35.64 ; 
      RECT 23.364 34.736 37.908 35.64 ; 
      RECT 18.036 34.736 23.292 35.64 ; 
      RECT 15.156 31.266 17.676 35.64 ; 
      RECT 0.54 34.736 15.084 35.64 ; 
      RECT 0 31.266 0.468 35.64 ; 
      RECT 37.836 31.266 38.448 34.928 ; 
      RECT 23.58 31.266 37.764 35.64 ; 
      RECT 20.592 31.266 23.508 34.928 ; 
      RECT 19.944 32.048 20.448 35.64 ; 
      RECT 14.94 31.664 19.836 34.928 ; 
      RECT 0.684 31.266 14.868 35.64 ; 
      RECT 0 31.266 0.612 34.928 ; 
      RECT 20.376 31.266 38.448 34.544 ; 
      RECT 0 31.664 20.304 34.544 ; 
      RECT 19.476 31.266 38.448 31.952 ; 
      RECT 0 31.266 19.404 34.544 ; 
      RECT 0 31.266 38.448 31.568 ; 
      RECT 0 39.44 38.448 39.96 ; 
      RECT 37.98 35.586 38.448 39.96 ; 
      RECT 23.364 39.056 37.908 39.96 ; 
      RECT 18.036 39.056 23.292 39.96 ; 
      RECT 15.156 35.586 17.676 39.96 ; 
      RECT 0.54 39.056 15.084 39.96 ; 
      RECT 0 35.586 0.468 39.96 ; 
      RECT 37.836 35.586 38.448 39.248 ; 
      RECT 23.58 35.586 37.764 39.96 ; 
      RECT 20.592 35.586 23.508 39.248 ; 
      RECT 19.944 36.368 20.448 39.96 ; 
      RECT 14.94 35.984 19.836 39.248 ; 
      RECT 0.684 35.586 14.868 39.96 ; 
      RECT 0 35.586 0.612 39.248 ; 
      RECT 20.376 35.586 38.448 38.864 ; 
      RECT 0 35.984 20.304 38.864 ; 
      RECT 19.476 35.586 38.448 36.272 ; 
      RECT 0 35.586 19.404 38.864 ; 
      RECT 0 35.586 38.448 35.888 ; 
      RECT 0 69.132 38.448 74.466 ; 
      RECT 29.412 39.852 38.448 74.466 ; 
      RECT 20.612 55.308 38.448 74.466 ; 
      RECT 24.228 44.94 38.448 74.466 ; 
      RECT 20.404 39.852 20.54 74.466 ; 
      RECT 20.196 39.852 20.332 74.466 ; 
      RECT 19.988 39.852 20.124 74.466 ; 
      RECT 19.78 39.852 19.916 74.466 ; 
      RECT 0 67.404 19.708 74.466 ; 
      RECT 18.74 56.46 38.448 68.268 ; 
      RECT 18.532 39.852 18.668 74.466 ; 
      RECT 18.324 39.852 18.46 74.466 ; 
      RECT 18.116 39.852 18.252 74.466 ; 
      RECT 17.908 39.852 18.044 74.466 ; 
      RECT 0 46.092 17.836 74.466 ; 
      RECT 0 54.732 19.708 66.54 ; 
      RECT 18.74 43.788 23.292 55.596 ; 
      RECT 23.364 45.708 38.448 74.466 ; 
      RECT 20.772 40.172 24.156 55.212 ; 
      RECT 16.02 42.06 19.116 53.868 ; 
      RECT 15.156 42.636 17.836 74.466 ; 
      RECT 0 44.94 15.084 74.466 ; 
      RECT 13.428 39.852 15.228 45.996 ; 
      RECT 28.548 39.852 29.34 74.466 ; 
      RECT 13.428 44.172 28.476 45.612 ; 
      RECT 9.972 42.636 13.356 74.466 ; 
      RECT 0 43.788 9.9 74.466 ; 
      RECT 27.684 39.852 38.448 44.844 ; 
      RECT 26.82 42.636 38.448 44.844 ; 
      RECT 0 43.788 26.748 44.844 ; 
      RECT 25.956 39.852 27.612 44.076 ; 
      RECT 20.612 42.636 38.448 44.076 ; 
      RECT 0.684 42.636 19.708 44.844 ; 
      RECT 18.74 42.444 19.708 74.466 ; 
      RECT 0 42.06 0.612 74.466 ; 
      RECT 19.188 39.852 20.7 42.924 ; 
      RECT 20.772 42.444 25.884 45.612 ; 
      RECT 12.564 42.444 15.948 44.844 ; 
      RECT 10.836 42.444 12.492 74.466 ; 
      RECT 0 42.06 10.764 42.924 ; 
      RECT 25.092 39.852 38.448 42.54 ; 
      RECT 19.188 40.172 25.02 42.54 ; 
      RECT 15.3 42.06 19.116 42.54 ; 
      RECT 11.7 39.852 15.228 42.54 ; 
      RECT 0 42.06 11.628 42.54 ; 
      RECT 23.364 39.852 38.448 42.348 ; 
      RECT 18.74 40.172 38.448 42.348 ; 
      RECT 0.54 39.852 17.836 42.348 ; 
      RECT 0 39.852 0.468 74.466 ; 
      RECT 0 39.852 23.292 41.196 ; 
      RECT 0 39.852 38.448 40.076 ; 
        RECT 0 76.268 38.448 76.788 ; 
        RECT 37.98 72.414 38.448 76.788 ; 
        RECT 23.364 75.884 37.908 76.788 ; 
        RECT 18.036 75.884 23.292 76.788 ; 
        RECT 15.156 72.414 17.676 76.788 ; 
        RECT 0.54 75.884 15.084 76.788 ; 
        RECT 0 72.414 0.468 76.788 ; 
        RECT 37.836 72.414 38.448 76.076 ; 
        RECT 23.58 72.414 37.764 76.788 ; 
        RECT 20.592 72.414 23.508 76.076 ; 
        RECT 19.944 73.196 20.448 76.788 ; 
        RECT 14.94 72.812 19.836 76.076 ; 
        RECT 0.684 72.414 14.868 76.788 ; 
        RECT 0 72.414 0.612 76.076 ; 
        RECT 20.376 72.414 38.448 75.692 ; 
        RECT 0 72.812 20.304 75.692 ; 
        RECT 19.476 72.414 38.448 73.1 ; 
        RECT 0 72.414 19.404 75.692 ; 
        RECT 0 72.414 38.448 72.716 ; 
        RECT 0 80.588 38.448 81.108 ; 
        RECT 37.98 76.734 38.448 81.108 ; 
        RECT 23.364 80.204 37.908 81.108 ; 
        RECT 18.036 80.204 23.292 81.108 ; 
        RECT 15.156 76.734 17.676 81.108 ; 
        RECT 0.54 80.204 15.084 81.108 ; 
        RECT 0 76.734 0.468 81.108 ; 
        RECT 37.836 76.734 38.448 80.396 ; 
        RECT 23.58 76.734 37.764 81.108 ; 
        RECT 20.592 76.734 23.508 80.396 ; 
        RECT 19.944 77.516 20.448 81.108 ; 
        RECT 14.94 77.132 19.836 80.396 ; 
        RECT 0.684 76.734 14.868 81.108 ; 
        RECT 0 76.734 0.612 80.396 ; 
        RECT 20.376 76.734 38.448 80.012 ; 
        RECT 0 77.132 20.304 80.012 ; 
        RECT 19.476 76.734 38.448 77.42 ; 
        RECT 0 76.734 19.404 80.012 ; 
        RECT 0 76.734 38.448 77.036 ; 
        RECT 0 84.908 38.448 85.428 ; 
        RECT 37.98 81.054 38.448 85.428 ; 
        RECT 23.364 84.524 37.908 85.428 ; 
        RECT 18.036 84.524 23.292 85.428 ; 
        RECT 15.156 81.054 17.676 85.428 ; 
        RECT 0.54 84.524 15.084 85.428 ; 
        RECT 0 81.054 0.468 85.428 ; 
        RECT 37.836 81.054 38.448 84.716 ; 
        RECT 23.58 81.054 37.764 85.428 ; 
        RECT 20.592 81.054 23.508 84.716 ; 
        RECT 19.944 81.836 20.448 85.428 ; 
        RECT 14.94 81.452 19.836 84.716 ; 
        RECT 0.684 81.054 14.868 85.428 ; 
        RECT 0 81.054 0.612 84.716 ; 
        RECT 20.376 81.054 38.448 84.332 ; 
        RECT 0 81.452 20.304 84.332 ; 
        RECT 19.476 81.054 38.448 81.74 ; 
        RECT 0 81.054 19.404 84.332 ; 
        RECT 0 81.054 38.448 81.356 ; 
        RECT 0 89.228 38.448 89.748 ; 
        RECT 37.98 85.374 38.448 89.748 ; 
        RECT 23.364 88.844 37.908 89.748 ; 
        RECT 18.036 88.844 23.292 89.748 ; 
        RECT 15.156 85.374 17.676 89.748 ; 
        RECT 0.54 88.844 15.084 89.748 ; 
        RECT 0 85.374 0.468 89.748 ; 
        RECT 37.836 85.374 38.448 89.036 ; 
        RECT 23.58 85.374 37.764 89.748 ; 
        RECT 20.592 85.374 23.508 89.036 ; 
        RECT 19.944 86.156 20.448 89.748 ; 
        RECT 14.94 85.772 19.836 89.036 ; 
        RECT 0.684 85.374 14.868 89.748 ; 
        RECT 0 85.374 0.612 89.036 ; 
        RECT 20.376 85.374 38.448 88.652 ; 
        RECT 0 85.772 20.304 88.652 ; 
        RECT 19.476 85.374 38.448 86.06 ; 
        RECT 0 85.374 19.404 88.652 ; 
        RECT 0 85.374 38.448 85.676 ; 
        RECT 0 93.548 38.448 94.068 ; 
        RECT 37.98 89.694 38.448 94.068 ; 
        RECT 23.364 93.164 37.908 94.068 ; 
        RECT 18.036 93.164 23.292 94.068 ; 
        RECT 15.156 89.694 17.676 94.068 ; 
        RECT 0.54 93.164 15.084 94.068 ; 
        RECT 0 89.694 0.468 94.068 ; 
        RECT 37.836 89.694 38.448 93.356 ; 
        RECT 23.58 89.694 37.764 94.068 ; 
        RECT 20.592 89.694 23.508 93.356 ; 
        RECT 19.944 90.476 20.448 94.068 ; 
        RECT 14.94 90.092 19.836 93.356 ; 
        RECT 0.684 89.694 14.868 94.068 ; 
        RECT 0 89.694 0.612 93.356 ; 
        RECT 20.376 89.694 38.448 92.972 ; 
        RECT 0 90.092 20.304 92.972 ; 
        RECT 19.476 89.694 38.448 90.38 ; 
        RECT 0 89.694 19.404 92.972 ; 
        RECT 0 89.694 38.448 89.996 ; 
        RECT 0 97.868 38.448 98.388 ; 
        RECT 37.98 94.014 38.448 98.388 ; 
        RECT 23.364 97.484 37.908 98.388 ; 
        RECT 18.036 97.484 23.292 98.388 ; 
        RECT 15.156 94.014 17.676 98.388 ; 
        RECT 0.54 97.484 15.084 98.388 ; 
        RECT 0 94.014 0.468 98.388 ; 
        RECT 37.836 94.014 38.448 97.676 ; 
        RECT 23.58 94.014 37.764 98.388 ; 
        RECT 20.592 94.014 23.508 97.676 ; 
        RECT 19.944 94.796 20.448 98.388 ; 
        RECT 14.94 94.412 19.836 97.676 ; 
        RECT 0.684 94.014 14.868 98.388 ; 
        RECT 0 94.014 0.612 97.676 ; 
        RECT 20.376 94.014 38.448 97.292 ; 
        RECT 0 94.412 20.304 97.292 ; 
        RECT 19.476 94.014 38.448 94.7 ; 
        RECT 0 94.014 19.404 97.292 ; 
        RECT 0 94.014 38.448 94.316 ; 
        RECT 0 102.188 38.448 102.708 ; 
        RECT 37.98 98.334 38.448 102.708 ; 
        RECT 23.364 101.804 37.908 102.708 ; 
        RECT 18.036 101.804 23.292 102.708 ; 
        RECT 15.156 98.334 17.676 102.708 ; 
        RECT 0.54 101.804 15.084 102.708 ; 
        RECT 0 98.334 0.468 102.708 ; 
        RECT 37.836 98.334 38.448 101.996 ; 
        RECT 23.58 98.334 37.764 102.708 ; 
        RECT 20.592 98.334 23.508 101.996 ; 
        RECT 19.944 99.116 20.448 102.708 ; 
        RECT 14.94 98.732 19.836 101.996 ; 
        RECT 0.684 98.334 14.868 102.708 ; 
        RECT 0 98.334 0.612 101.996 ; 
        RECT 20.376 98.334 38.448 101.612 ; 
        RECT 0 98.732 20.304 101.612 ; 
        RECT 19.476 98.334 38.448 99.02 ; 
        RECT 0 98.334 19.404 101.612 ; 
        RECT 0 98.334 38.448 98.636 ; 
        RECT 0 106.508 38.448 107.028 ; 
        RECT 37.98 102.654 38.448 107.028 ; 
        RECT 23.364 106.124 37.908 107.028 ; 
        RECT 18.036 106.124 23.292 107.028 ; 
        RECT 15.156 102.654 17.676 107.028 ; 
        RECT 0.54 106.124 15.084 107.028 ; 
        RECT 0 102.654 0.468 107.028 ; 
        RECT 37.836 102.654 38.448 106.316 ; 
        RECT 23.58 102.654 37.764 107.028 ; 
        RECT 20.592 102.654 23.508 106.316 ; 
        RECT 19.944 103.436 20.448 107.028 ; 
        RECT 14.94 103.052 19.836 106.316 ; 
        RECT 0.684 102.654 14.868 107.028 ; 
        RECT 0 102.654 0.612 106.316 ; 
        RECT 20.376 102.654 38.448 105.932 ; 
        RECT 0 103.052 20.304 105.932 ; 
        RECT 19.476 102.654 38.448 103.34 ; 
        RECT 0 102.654 19.404 105.932 ; 
        RECT 0 102.654 38.448 102.956 ; 
        RECT 0 110.828 38.448 111.348 ; 
        RECT 37.98 106.974 38.448 111.348 ; 
        RECT 23.364 110.444 37.908 111.348 ; 
        RECT 18.036 110.444 23.292 111.348 ; 
        RECT 15.156 106.974 17.676 111.348 ; 
        RECT 0.54 110.444 15.084 111.348 ; 
        RECT 0 106.974 0.468 111.348 ; 
        RECT 37.836 106.974 38.448 110.636 ; 
        RECT 23.58 106.974 37.764 111.348 ; 
        RECT 20.592 106.974 23.508 110.636 ; 
        RECT 19.944 107.756 20.448 111.348 ; 
        RECT 14.94 107.372 19.836 110.636 ; 
        RECT 0.684 106.974 14.868 111.348 ; 
        RECT 0 106.974 0.612 110.636 ; 
        RECT 20.376 106.974 38.448 110.252 ; 
        RECT 0 107.372 20.304 110.252 ; 
        RECT 19.476 106.974 38.448 107.66 ; 
        RECT 0 106.974 19.404 110.252 ; 
        RECT 0 106.974 38.448 107.276 ; 
  LAYER M4 ; 
      RECT 6.428 46.704 32.01 46.8 ; 
      RECT 6.428 47.856 32.01 47.952 ; 
      RECT 6.428 49.392 32.01 49.488 ; 
      RECT 6.428 49.776 32.01 49.872 ; 
      RECT 6.428 51.12 32.01 51.216 ; 
      RECT 29.996 42.54 30.332 42.636 ; 
      RECT 29.276 44.268 29.744 44.364 ; 
      RECT 29.276 46.896 29.744 46.992 ; 
      RECT 29.276 48.048 29.744 48.144 ; 
      RECT 26.714 44.268 28.992 44.364 ; 
      RECT 26.972 47.376 27.404 47.472 ; 
      RECT 21.628 48.876 26 48.972 ; 
      RECT 24.38 47.148 24.716 47.244 ; 
      RECT 21.244 51.948 24.716 52.044 ; 
      RECT 24.38 52.332 24.716 52.428 ; 
      RECT 23.668 45.228 24.004 45.324 ; 
      RECT 23.516 50.604 23.852 50.7 ; 
      RECT 22.804 44.844 23.14 44.94 ; 
      RECT 21.948 39.692 23 39.788 ; 
      RECT 21.948 74.252 23 74.348 ; 
      RECT 22.012 50.796 22.988 50.892 ; 
      RECT 22.652 51.372 22.988 51.468 ; 
      RECT 16.828 52.332 22.988 52.428 ; 
      RECT 22.652 53.484 22.988 53.58 ; 
      RECT 21.716 73.868 22.768 73.964 ; 
      RECT 21.712 39.308 22.764 39.404 ; 
      RECT 21.56 38.924 22.612 39.02 ; 
      RECT 21.56 73.1 22.612 73.196 ; 
      RECT 22.22 55.212 22.556 55.308 ; 
      RECT 19.132 56.748 22.556 56.844 ; 
      RECT 20.668 65.772 22.556 65.868 ; 
      RECT 22.22 66.156 22.556 66.252 ; 
      RECT 21.368 38.54 22.42 38.636 ; 
      RECT 21.368 72.716 22.42 72.812 ; 
      RECT 20.476 62.124 22.256 62.22 ; 
      RECT 21.192 38.156 22.244 38.252 ; 
      RECT 21.192 74.06 22.244 74.156 ; 
      RECT 20.996 39.5 22.048 39.596 ; 
      RECT 20.996 73.676 22.048 73.772 ; 
      RECT 21.52 51.372 22.004 51.468 ; 
      RECT 21.436 59.82 21.968 59.916 ; 
      RECT 20.808 39.116 21.86 39.212 ; 
      RECT 20.808 73.292 21.86 73.388 ; 
      RECT 20.668 37.964 21.72 38.06 ; 
      RECT 20.668 72.908 21.72 73.004 ; 
      RECT 17.404 66.156 21.68 66.252 ; 
      RECT 21.344 70.764 21.68 70.86 ; 
      RECT 20.444 37.388 21.496 37.484 ; 
      RECT 20.444 72.524 21.496 72.62 ; 
      RECT 21.052 55.212 21.392 55.308 ; 
      RECT 16.636 57.516 21.104 57.612 ; 
      RECT 19.216 48.876 21.044 48.972 ; 
      RECT 18.524 40.268 19.592 40.364 ; 
      RECT 18.524 71.948 19.592 72.044 ; 
      RECT 19.072 55.02 19.508 55.116 ; 
      RECT 18.432 39.884 19.4 39.98 ; 
      RECT 18.432 74.444 19.4 74.54 ; 
      RECT 18.208 37.964 19.176 38.06 ; 
      RECT 18.324 74.828 19.176 74.924 ; 
      RECT 18.788 53.484 19.124 53.58 ; 
      RECT 17.992 38.348 18.984 38.444 ; 
      RECT 17.992 74.252 18.984 74.348 ; 
      RECT 17.056 63.852 18.74 63.948 ; 
      RECT 16.928 39.692 17.996 39.788 ; 
      RECT 16.928 74.828 17.996 74.924 ; 
      RECT 17.488 58.092 17.972 58.188 ; 
      RECT 17.456 70.764 17.792 70.86 ; 
      RECT 16.792 39.308 17.78 39.404 ; 
      RECT 16.524 73.1 17.78 73.196 ; 
      RECT 16.688 38.924 17.608 39.02 ; 
      RECT 16.64 74.444 17.608 74.54 ; 
      RECT 16.476 38.54 17.396 38.636 ; 
      RECT 17.06 64.428 17.396 64.524 ; 
      RECT 16.276 72.716 17.396 72.812 ; 
      RECT 16.296 38.156 17.216 38.252 ; 
      RECT 16.296 74.06 17.216 74.156 ; 
      RECT 12.448 53.484 17.204 53.58 ; 
      RECT 16.144 39.116 17.064 39.212 ; 
      RECT 16.144 73.676 17.064 73.772 ; 
      RECT 16.072 38.732 16.844 38.828 ; 
      RECT 16.072 73.292 16.844 73.388 ; 
      RECT 15.876 38.348 16.648 38.444 ; 
      RECT 15.876 72.908 16.648 73.004 ; 
      RECT 15.892 57.132 16.628 57.228 ; 
      RECT 15.668 37.964 16.44 38.06 ; 
      RECT 15.668 72.524 16.44 72.62 ; 
      RECT 13.732 46.38 16.436 46.476 ; 
      RECT 15.892 57.516 16.228 57.612 ; 
      RECT 14.816 40.076 15.868 40.172 ; 
      RECT 15.032 55.212 15.48 55.308 ; 
      RECT 13.58 47.148 13.916 47.244 ; 
  LAYER V4 ; 
      RECT 30.192 42.54 30.288 42.636 ; 
      RECT 30.192 46.704 30.288 46.8 ; 
      RECT 29.52 44.268 29.616 44.364 ; 
      RECT 29.52 46.896 29.616 46.992 ; 
      RECT 29.52 48.048 29.616 48.144 ; 
      RECT 27.024 44.268 27.12 44.364 ; 
      RECT 27.024 47.376 27.12 47.472 ; 
      RECT 24.576 47.148 24.672 47.244 ; 
      RECT 24.576 47.856 24.672 47.952 ; 
      RECT 24.576 51.948 24.672 52.044 ; 
      RECT 24.576 52.332 24.672 52.428 ; 
      RECT 23.712 45.228 23.808 45.324 ; 
      RECT 23.712 49.392 23.808 49.488 ; 
      RECT 23.712 50.604 23.808 50.7 ; 
      RECT 23.712 51.12 23.808 51.216 ; 
      RECT 22.848 44.844 22.944 44.94 ; 
      RECT 22.848 49.776 22.944 49.872 ; 
      RECT 22.848 50.796 22.944 50.892 ; 
      RECT 22.848 51.372 22.944 51.468 ; 
      RECT 22.848 52.332 22.944 52.428 ; 
      RECT 22.848 53.484 22.944 53.58 ; 
      RECT 22.416 55.212 22.512 55.308 ; 
      RECT 22.416 56.748 22.512 56.844 ; 
      RECT 22.416 65.772 22.512 65.868 ; 
      RECT 22.416 66.156 22.512 66.252 ; 
      RECT 22.056 39.692 22.152 39.788 ; 
      RECT 22.056 50.796 22.152 50.892 ; 
      RECT 22.056 74.252 22.152 74.348 ; 
      RECT 21.864 39.308 21.96 39.404 ; 
      RECT 21.864 51.372 21.96 51.468 ; 
      RECT 21.864 73.868 21.96 73.964 ; 
      RECT 21.672 38.924 21.768 39.02 ; 
      RECT 21.672 48.876 21.768 48.972 ; 
      RECT 21.672 73.1 21.768 73.196 ; 
      RECT 21.48 38.54 21.576 38.636 ; 
      RECT 21.48 59.82 21.576 59.916 ; 
      RECT 21.48 70.764 21.576 70.86 ; 
      RECT 21.48 72.716 21.576 72.812 ; 
      RECT 21.288 38.156 21.384 38.252 ; 
      RECT 21.288 51.948 21.384 52.044 ; 
      RECT 21.288 74.06 21.384 74.156 ; 
      RECT 21.096 39.5 21.192 39.596 ; 
      RECT 21.096 55.212 21.192 55.308 ; 
      RECT 21.096 73.676 21.192 73.772 ; 
      RECT 20.904 39.116 21 39.212 ; 
      RECT 20.904 48.876 21 48.972 ; 
      RECT 20.904 73.292 21 73.388 ; 
      RECT 20.712 37.964 20.808 38.06 ; 
      RECT 20.712 65.772 20.808 65.868 ; 
      RECT 20.712 72.908 20.808 73.004 ; 
      RECT 20.52 37.388 20.616 37.484 ; 
      RECT 20.52 62.124 20.616 62.22 ; 
      RECT 20.52 72.524 20.616 72.62 ; 
      RECT 19.368 40.268 19.464 40.364 ; 
      RECT 19.368 55.02 19.464 55.116 ; 
      RECT 19.368 71.948 19.464 72.044 ; 
      RECT 19.176 39.884 19.272 39.98 ; 
      RECT 19.176 56.748 19.272 56.844 ; 
      RECT 19.176 74.444 19.272 74.54 ; 
      RECT 18.984 37.964 19.08 38.06 ; 
      RECT 18.984 53.484 19.08 53.58 ; 
      RECT 18.984 74.828 19.08 74.924 ; 
      RECT 18.6 38.348 18.696 38.444 ; 
      RECT 18.6 63.852 18.696 63.948 ; 
      RECT 18.6 74.252 18.696 74.348 ; 
      RECT 17.832 39.692 17.928 39.788 ; 
      RECT 17.832 58.092 17.928 58.188 ; 
      RECT 17.832 74.828 17.928 74.924 ; 
      RECT 17.64 39.308 17.736 39.404 ; 
      RECT 17.64 70.764 17.736 70.86 ; 
      RECT 17.64 73.1 17.736 73.196 ; 
      RECT 17.448 38.924 17.544 39.02 ; 
      RECT 17.448 66.156 17.544 66.252 ; 
      RECT 17.448 74.444 17.544 74.54 ; 
      RECT 17.256 38.54 17.352 38.636 ; 
      RECT 17.256 64.428 17.352 64.524 ; 
      RECT 17.256 72.716 17.352 72.812 ; 
      RECT 17.064 38.156 17.16 38.252 ; 
      RECT 17.064 53.484 17.16 53.58 ; 
      RECT 17.064 74.06 17.16 74.156 ; 
      RECT 16.872 39.116 16.968 39.212 ; 
      RECT 16.872 52.332 16.968 52.428 ; 
      RECT 16.872 73.676 16.968 73.772 ; 
      RECT 16.68 38.732 16.776 38.828 ; 
      RECT 16.68 57.516 16.776 57.612 ; 
      RECT 16.68 73.292 16.776 73.388 ; 
      RECT 16.488 38.348 16.584 38.444 ; 
      RECT 16.488 57.132 16.584 57.228 ; 
      RECT 16.488 72.908 16.584 73.004 ; 
      RECT 16.296 37.964 16.392 38.06 ; 
      RECT 16.296 46.38 16.392 46.476 ; 
      RECT 16.296 72.524 16.392 72.62 ; 
      RECT 15.936 57.132 16.032 57.228 ; 
      RECT 15.936 57.516 16.032 57.612 ; 
      RECT 15.268 40.076 15.364 40.172 ; 
      RECT 15.268 55.212 15.364 55.308 ; 
      RECT 13.776 46.38 13.872 46.476 ; 
      RECT 13.776 47.148 13.872 47.244 ; 
  LAYER M5 ; 
      RECT 30.192 42.496 30.288 46.844 ; 
      RECT 29.52 44.214 29.616 48.344 ; 
      RECT 27.024 44.19 27.12 47.52 ; 
      RECT 24.576 47.104 24.672 47.996 ; 
      RECT 24.576 51.904 24.672 52.472 ; 
      RECT 23.712 45.184 23.808 49.532 ; 
      RECT 23.712 50.56 23.808 51.26 ; 
      RECT 22.848 44.8 22.944 49.916 ; 
      RECT 22.848 50.752 22.944 51.512 ; 
      RECT 22.848 52.288 22.944 53.624 ; 
      RECT 22.416 55.168 22.512 56.888 ; 
      RECT 22.416 65.728 22.512 66.296 ; 
      RECT 22.056 41.04 22.152 71.372 ; 
      RECT 21.864 41.04 21.96 71.372 ; 
      RECT 21.672 41.04 21.768 71.372 ; 
      RECT 21.48 41.04 21.576 71.372 ; 
      RECT 21.288 41.04 21.384 71.372 ; 
      RECT 21.096 41.04 21.192 71.372 ; 
      RECT 20.904 41.04 21 71.372 ; 
      RECT 20.712 41.04 20.808 71.372 ; 
      RECT 20.52 41.04 20.616 71.372 ; 
      RECT 19.368 39.992 19.464 72.124 ; 
      RECT 19.176 37.908 19.272 75.224 ; 
      RECT 18.984 37.784 19.08 75.22 ; 
      RECT 18.6 37.968 18.696 75.224 ; 
      RECT 17.832 37.964 17.928 75.036 ; 
      RECT 17.64 37.964 17.736 75.036 ; 
      RECT 17.448 37.964 17.544 75.036 ; 
      RECT 17.256 37.964 17.352 75.036 ; 
      RECT 17.064 37.964 17.16 75.036 ; 
      RECT 16.872 37.848 16.968 75.036 ; 
      RECT 16.68 37.672 16.776 75.04 ; 
      RECT 16.488 37.524 16.584 75.044 ; 
      RECT 16.296 37.284 16.392 75.044 ; 
      RECT 15.936 57.088 16.032 57.656 ; 
      RECT 15.268 40.004 15.364 55.38 ; 
      RECT 13.776 46.336 13.872 47.288 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 38.016 112.176 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 38.016 112.176 ; 
  END 
END srambank_64x4x18_6t122 
