VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_128x4x20_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_128x4x20_6t122 0 0 ; 
  SIZE 64 BY 120.96 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.688 65.768 4.88 ; 
        RECT 0.376 9.008 65.768 9.2 ; 
        RECT 0.376 13.328 65.768 13.52 ; 
        RECT 0.376 17.648 65.768 17.84 ; 
        RECT 0.376 21.968 65.768 22.16 ; 
        RECT 0.376 26.288 65.768 26.48 ; 
        RECT 0.376 30.608 65.768 30.8 ; 
        RECT 0.376 34.928 65.768 35.12 ; 
        RECT 0.376 39.248 65.768 39.44 ; 
        RECT 0.376 43.568 65.768 43.76 ; 
        RECT 14.256 45.492 51.84 46.356 ; 
        RECT 36.788 59.508 37.352 59.604 ; 
        RECT 36.264 44.372 37.316 44.468 ; 
        RECT 29.592 58.164 36.504 59.028 ; 
        RECT 29.592 70.836 36.504 71.7 ; 
        RECT 0.376 80.396 65.768 80.588 ; 
        RECT 0.376 84.716 65.768 84.908 ; 
        RECT 0.376 89.036 65.768 89.228 ; 
        RECT 0.376 93.356 65.768 93.548 ; 
        RECT 0.376 97.676 65.768 97.868 ; 
        RECT 0.376 101.996 65.768 102.188 ; 
        RECT 0.376 106.316 65.768 106.508 ; 
        RECT 0.376 110.636 65.768 110.828 ; 
        RECT 0.376 114.956 65.768 115.148 ; 
        RECT 0.376 119.276 65.768 119.468 ; 
      LAYER M3 ; 
        RECT 65.576 0.866 65.648 5.506 ; 
        RECT 37.136 0.868 37.208 5.504 ; 
        RECT 31.52 1.028 31.88 5.484 ; 
        RECT 28.928 0.868 29 5.504 ; 
        RECT 0.488 0.866 0.56 5.506 ; 
        RECT 65.576 5.186 65.648 9.826 ; 
        RECT 37.136 5.188 37.208 9.824 ; 
        RECT 31.52 5.348 31.88 9.804 ; 
        RECT 28.928 5.188 29 9.824 ; 
        RECT 0.488 5.186 0.56 9.826 ; 
        RECT 65.576 9.506 65.648 14.146 ; 
        RECT 37.136 9.508 37.208 14.144 ; 
        RECT 31.52 9.668 31.88 14.124 ; 
        RECT 28.928 9.508 29 14.144 ; 
        RECT 0.488 9.506 0.56 14.146 ; 
        RECT 65.576 13.826 65.648 18.466 ; 
        RECT 37.136 13.828 37.208 18.464 ; 
        RECT 31.52 13.988 31.88 18.444 ; 
        RECT 28.928 13.828 29 18.464 ; 
        RECT 0.488 13.826 0.56 18.466 ; 
        RECT 65.576 18.146 65.648 22.786 ; 
        RECT 37.136 18.148 37.208 22.784 ; 
        RECT 31.52 18.308 31.88 22.764 ; 
        RECT 28.928 18.148 29 22.784 ; 
        RECT 0.488 18.146 0.56 22.786 ; 
        RECT 65.576 22.466 65.648 27.106 ; 
        RECT 37.136 22.468 37.208 27.104 ; 
        RECT 31.52 22.628 31.88 27.084 ; 
        RECT 28.928 22.468 29 27.104 ; 
        RECT 0.488 22.466 0.56 27.106 ; 
        RECT 65.576 26.786 65.648 31.426 ; 
        RECT 37.136 26.788 37.208 31.424 ; 
        RECT 31.52 26.948 31.88 31.404 ; 
        RECT 28.928 26.788 29 31.424 ; 
        RECT 0.488 26.786 0.56 31.426 ; 
        RECT 65.576 31.106 65.648 35.746 ; 
        RECT 37.136 31.108 37.208 35.744 ; 
        RECT 31.52 31.268 31.88 35.724 ; 
        RECT 28.928 31.108 29 35.744 ; 
        RECT 0.488 31.106 0.56 35.746 ; 
        RECT 65.576 35.426 65.648 40.066 ; 
        RECT 37.136 35.428 37.208 40.064 ; 
        RECT 31.52 35.588 31.88 40.044 ; 
        RECT 28.928 35.428 29 40.064 ; 
        RECT 0.488 35.426 0.56 40.066 ; 
        RECT 65.576 39.746 65.648 44.386 ; 
        RECT 37.136 39.748 37.208 44.384 ; 
        RECT 31.52 39.908 31.88 44.364 ; 
        RECT 28.928 39.748 29 44.384 ; 
        RECT 0.488 39.746 0.56 44.386 ; 
        RECT 65.556 44.042 65.628 76.87 ; 
        RECT 37.188 59.32 37.26 76.714 ; 
        RECT 37.116 44.174 37.188 44.726 ; 
        RECT 31.644 45.336 32.58 75.668 ; 
        RECT 31.5 75.336 31.86 76.84 ; 
        RECT 31.5 44.2 31.86 45.704 ; 
        RECT 0.468 44.042 0.54 76.87 ; 
        RECT 65.576 76.574 65.648 81.214 ; 
        RECT 37.136 76.576 37.208 81.212 ; 
        RECT 31.52 76.736 31.88 81.192 ; 
        RECT 28.928 76.576 29 81.212 ; 
        RECT 0.488 76.574 0.56 81.214 ; 
        RECT 65.576 80.894 65.648 85.534 ; 
        RECT 37.136 80.896 37.208 85.532 ; 
        RECT 31.52 81.056 31.88 85.512 ; 
        RECT 28.928 80.896 29 85.532 ; 
        RECT 0.488 80.894 0.56 85.534 ; 
        RECT 65.576 85.214 65.648 89.854 ; 
        RECT 37.136 85.216 37.208 89.852 ; 
        RECT 31.52 85.376 31.88 89.832 ; 
        RECT 28.928 85.216 29 89.852 ; 
        RECT 0.488 85.214 0.56 89.854 ; 
        RECT 65.576 89.534 65.648 94.174 ; 
        RECT 37.136 89.536 37.208 94.172 ; 
        RECT 31.52 89.696 31.88 94.152 ; 
        RECT 28.928 89.536 29 94.172 ; 
        RECT 0.488 89.534 0.56 94.174 ; 
        RECT 65.576 93.854 65.648 98.494 ; 
        RECT 37.136 93.856 37.208 98.492 ; 
        RECT 31.52 94.016 31.88 98.472 ; 
        RECT 28.928 93.856 29 98.492 ; 
        RECT 0.488 93.854 0.56 98.494 ; 
        RECT 65.576 98.174 65.648 102.814 ; 
        RECT 37.136 98.176 37.208 102.812 ; 
        RECT 31.52 98.336 31.88 102.792 ; 
        RECT 28.928 98.176 29 102.812 ; 
        RECT 0.488 98.174 0.56 102.814 ; 
        RECT 65.576 102.494 65.648 107.134 ; 
        RECT 37.136 102.496 37.208 107.132 ; 
        RECT 31.52 102.656 31.88 107.112 ; 
        RECT 28.928 102.496 29 107.132 ; 
        RECT 0.488 102.494 0.56 107.134 ; 
        RECT 65.576 106.814 65.648 111.454 ; 
        RECT 37.136 106.816 37.208 111.452 ; 
        RECT 31.52 106.976 31.88 111.432 ; 
        RECT 28.928 106.816 29 111.452 ; 
        RECT 0.488 106.814 0.56 111.454 ; 
        RECT 65.576 111.134 65.648 115.774 ; 
        RECT 37.136 111.136 37.208 115.772 ; 
        RECT 31.52 111.296 31.88 115.752 ; 
        RECT 28.928 111.136 29 115.772 ; 
        RECT 0.488 111.134 0.56 115.774 ; 
        RECT 65.576 115.454 65.648 120.094 ; 
        RECT 37.136 115.456 37.208 120.092 ; 
        RECT 31.52 115.616 31.88 120.072 ; 
        RECT 28.928 115.456 29 120.092 ; 
        RECT 0.488 115.454 0.56 120.094 ; 
      LAYER V3 ; 
        RECT 0.488 4.688 0.56 4.88 ; 
        RECT 28.928 4.688 29 4.88 ; 
        RECT 31.52 4.688 31.88 4.88 ; 
        RECT 37.136 4.688 37.208 4.88 ; 
        RECT 65.576 4.688 65.648 4.88 ; 
        RECT 0.488 9.008 0.56 9.2 ; 
        RECT 28.928 9.008 29 9.2 ; 
        RECT 31.52 9.008 31.88 9.2 ; 
        RECT 37.136 9.008 37.208 9.2 ; 
        RECT 65.576 9.008 65.648 9.2 ; 
        RECT 0.488 13.328 0.56 13.52 ; 
        RECT 28.928 13.328 29 13.52 ; 
        RECT 31.52 13.328 31.88 13.52 ; 
        RECT 37.136 13.328 37.208 13.52 ; 
        RECT 65.576 13.328 65.648 13.52 ; 
        RECT 0.488 17.648 0.56 17.84 ; 
        RECT 28.928 17.648 29 17.84 ; 
        RECT 31.52 17.648 31.88 17.84 ; 
        RECT 37.136 17.648 37.208 17.84 ; 
        RECT 65.576 17.648 65.648 17.84 ; 
        RECT 0.488 21.968 0.56 22.16 ; 
        RECT 28.928 21.968 29 22.16 ; 
        RECT 31.52 21.968 31.88 22.16 ; 
        RECT 37.136 21.968 37.208 22.16 ; 
        RECT 65.576 21.968 65.648 22.16 ; 
        RECT 0.488 26.288 0.56 26.48 ; 
        RECT 28.928 26.288 29 26.48 ; 
        RECT 31.52 26.288 31.88 26.48 ; 
        RECT 37.136 26.288 37.208 26.48 ; 
        RECT 65.576 26.288 65.648 26.48 ; 
        RECT 0.488 30.608 0.56 30.8 ; 
        RECT 28.928 30.608 29 30.8 ; 
        RECT 31.52 30.608 31.88 30.8 ; 
        RECT 37.136 30.608 37.208 30.8 ; 
        RECT 65.576 30.608 65.648 30.8 ; 
        RECT 0.488 34.928 0.56 35.12 ; 
        RECT 28.928 34.928 29 35.12 ; 
        RECT 31.52 34.928 31.88 35.12 ; 
        RECT 37.136 34.928 37.208 35.12 ; 
        RECT 65.576 34.928 65.648 35.12 ; 
        RECT 0.488 39.248 0.56 39.44 ; 
        RECT 28.928 39.248 29 39.44 ; 
        RECT 31.52 39.248 31.88 39.44 ; 
        RECT 37.136 39.248 37.208 39.44 ; 
        RECT 65.576 39.248 65.648 39.44 ; 
        RECT 0.488 43.568 0.56 43.76 ; 
        RECT 28.928 43.568 29 43.76 ; 
        RECT 31.52 43.568 31.88 43.76 ; 
        RECT 37.136 43.568 37.208 43.76 ; 
        RECT 65.576 43.568 65.648 43.76 ; 
        RECT 31.66 70.836 31.732 71.7 ; 
        RECT 31.66 58.164 31.732 59.028 ; 
        RECT 31.66 45.492 31.732 46.356 ; 
        RECT 31.868 70.836 31.94 71.7 ; 
        RECT 31.868 58.164 31.94 59.028 ; 
        RECT 31.868 45.492 31.94 46.356 ; 
        RECT 32.076 70.836 32.148 71.7 ; 
        RECT 32.076 58.164 32.148 59.028 ; 
        RECT 32.076 45.492 32.148 46.356 ; 
        RECT 32.284 70.836 32.356 71.7 ; 
        RECT 32.284 58.164 32.356 59.028 ; 
        RECT 32.284 45.492 32.356 46.356 ; 
        RECT 32.492 70.836 32.564 71.7 ; 
        RECT 32.492 58.164 32.564 59.028 ; 
        RECT 32.492 45.492 32.564 46.356 ; 
        RECT 37.116 44.372 37.188 44.468 ; 
        RECT 37.188 59.508 37.26 59.604 ; 
        RECT 0.488 80.396 0.56 80.588 ; 
        RECT 28.928 80.396 29 80.588 ; 
        RECT 31.52 80.396 31.88 80.588 ; 
        RECT 37.136 80.396 37.208 80.588 ; 
        RECT 65.576 80.396 65.648 80.588 ; 
        RECT 0.488 84.716 0.56 84.908 ; 
        RECT 28.928 84.716 29 84.908 ; 
        RECT 31.52 84.716 31.88 84.908 ; 
        RECT 37.136 84.716 37.208 84.908 ; 
        RECT 65.576 84.716 65.648 84.908 ; 
        RECT 0.488 89.036 0.56 89.228 ; 
        RECT 28.928 89.036 29 89.228 ; 
        RECT 31.52 89.036 31.88 89.228 ; 
        RECT 37.136 89.036 37.208 89.228 ; 
        RECT 65.576 89.036 65.648 89.228 ; 
        RECT 0.488 93.356 0.56 93.548 ; 
        RECT 28.928 93.356 29 93.548 ; 
        RECT 31.52 93.356 31.88 93.548 ; 
        RECT 37.136 93.356 37.208 93.548 ; 
        RECT 65.576 93.356 65.648 93.548 ; 
        RECT 0.488 97.676 0.56 97.868 ; 
        RECT 28.928 97.676 29 97.868 ; 
        RECT 31.52 97.676 31.88 97.868 ; 
        RECT 37.136 97.676 37.208 97.868 ; 
        RECT 65.576 97.676 65.648 97.868 ; 
        RECT 0.488 101.996 0.56 102.188 ; 
        RECT 28.928 101.996 29 102.188 ; 
        RECT 31.52 101.996 31.88 102.188 ; 
        RECT 37.136 101.996 37.208 102.188 ; 
        RECT 65.576 101.996 65.648 102.188 ; 
        RECT 0.488 106.316 0.56 106.508 ; 
        RECT 28.928 106.316 29 106.508 ; 
        RECT 31.52 106.316 31.88 106.508 ; 
        RECT 37.136 106.316 37.208 106.508 ; 
        RECT 65.576 106.316 65.648 106.508 ; 
        RECT 0.488 110.636 0.56 110.828 ; 
        RECT 28.928 110.636 29 110.828 ; 
        RECT 31.52 110.636 31.88 110.828 ; 
        RECT 37.136 110.636 37.208 110.828 ; 
        RECT 65.576 110.636 65.648 110.828 ; 
        RECT 0.488 114.956 0.56 115.148 ; 
        RECT 28.928 114.956 29 115.148 ; 
        RECT 31.52 114.956 31.88 115.148 ; 
        RECT 37.136 114.956 37.208 115.148 ; 
        RECT 65.576 114.956 65.648 115.148 ; 
        RECT 0.488 119.276 0.56 119.468 ; 
        RECT 28.928 119.276 29 119.468 ; 
        RECT 31.52 119.276 31.88 119.468 ; 
        RECT 37.136 119.276 37.208 119.468 ; 
        RECT 65.576 119.276 65.648 119.468 ; 
      LAYER M5 ; 
        RECT 36.864 44.3 36.96 59.676 ; 
      LAYER V4 ; 
        RECT 36.864 59.508 36.96 59.604 ; 
        RECT 36.864 45.492 36.96 46.356 ; 
        RECT 36.864 44.372 36.96 44.468 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.304 65.748 4.496 ; 
        RECT 0.376 8.624 65.748 8.816 ; 
        RECT 0.376 12.944 65.748 13.136 ; 
        RECT 0.376 17.264 65.748 17.456 ; 
        RECT 0.376 21.584 65.748 21.776 ; 
        RECT 0.376 25.904 65.748 26.096 ; 
        RECT 0.376 30.224 65.748 30.416 ; 
        RECT 0.376 34.544 65.748 34.736 ; 
        RECT 0.376 38.864 65.748 39.056 ; 
        RECT 0.376 43.184 65.748 43.376 ; 
        RECT 14.256 47.22 51.84 48.084 ; 
        RECT 29.592 59.892 36.504 60.756 ; 
        RECT 29.592 72.564 36.504 73.428 ; 
        RECT 0.376 80.012 65.748 80.204 ; 
        RECT 0.376 84.332 65.748 84.524 ; 
        RECT 0.376 88.652 65.748 88.844 ; 
        RECT 0.376 92.972 65.748 93.164 ; 
        RECT 0.376 97.292 65.748 97.484 ; 
        RECT 0.376 101.612 65.748 101.804 ; 
        RECT 0.376 105.932 65.748 106.124 ; 
        RECT 0.376 110.252 65.748 110.444 ; 
        RECT 0.376 114.572 65.748 114.764 ; 
        RECT 0.376 118.892 65.748 119.084 ; 
      LAYER M3 ; 
        RECT 65.432 0.866 65.504 5.506 ; 
        RECT 37.352 0.866 37.424 5.506 ; 
        RECT 34.292 1.012 34.436 5.468 ; 
        RECT 33.68 1.012 33.788 5.468 ; 
        RECT 28.712 0.866 28.784 5.506 ; 
        RECT 0.632 0.866 0.704 5.506 ; 
        RECT 65.432 5.186 65.504 9.826 ; 
        RECT 37.352 5.186 37.424 9.826 ; 
        RECT 34.292 5.332 34.436 9.788 ; 
        RECT 33.68 5.332 33.788 9.788 ; 
        RECT 28.712 5.186 28.784 9.826 ; 
        RECT 0.632 5.186 0.704 9.826 ; 
        RECT 65.432 9.506 65.504 14.146 ; 
        RECT 37.352 9.506 37.424 14.146 ; 
        RECT 34.292 9.652 34.436 14.108 ; 
        RECT 33.68 9.652 33.788 14.108 ; 
        RECT 28.712 9.506 28.784 14.146 ; 
        RECT 0.632 9.506 0.704 14.146 ; 
        RECT 65.432 13.826 65.504 18.466 ; 
        RECT 37.352 13.826 37.424 18.466 ; 
        RECT 34.292 13.972 34.436 18.428 ; 
        RECT 33.68 13.972 33.788 18.428 ; 
        RECT 28.712 13.826 28.784 18.466 ; 
        RECT 0.632 13.826 0.704 18.466 ; 
        RECT 65.432 18.146 65.504 22.786 ; 
        RECT 37.352 18.146 37.424 22.786 ; 
        RECT 34.292 18.292 34.436 22.748 ; 
        RECT 33.68 18.292 33.788 22.748 ; 
        RECT 28.712 18.146 28.784 22.786 ; 
        RECT 0.632 18.146 0.704 22.786 ; 
        RECT 65.432 22.466 65.504 27.106 ; 
        RECT 37.352 22.466 37.424 27.106 ; 
        RECT 34.292 22.612 34.436 27.068 ; 
        RECT 33.68 22.612 33.788 27.068 ; 
        RECT 28.712 22.466 28.784 27.106 ; 
        RECT 0.632 22.466 0.704 27.106 ; 
        RECT 65.432 26.786 65.504 31.426 ; 
        RECT 37.352 26.786 37.424 31.426 ; 
        RECT 34.292 26.932 34.436 31.388 ; 
        RECT 33.68 26.932 33.788 31.388 ; 
        RECT 28.712 26.786 28.784 31.426 ; 
        RECT 0.632 26.786 0.704 31.426 ; 
        RECT 65.432 31.106 65.504 35.746 ; 
        RECT 37.352 31.106 37.424 35.746 ; 
        RECT 34.292 31.252 34.436 35.708 ; 
        RECT 33.68 31.252 33.788 35.708 ; 
        RECT 28.712 31.106 28.784 35.746 ; 
        RECT 0.632 31.106 0.704 35.746 ; 
        RECT 65.432 35.426 65.504 40.066 ; 
        RECT 37.352 35.426 37.424 40.066 ; 
        RECT 34.292 35.572 34.436 40.028 ; 
        RECT 33.68 35.572 33.788 40.028 ; 
        RECT 28.712 35.426 28.784 40.066 ; 
        RECT 0.632 35.426 0.704 40.066 ; 
        RECT 65.432 39.746 65.504 44.386 ; 
        RECT 37.352 39.746 37.424 44.386 ; 
        RECT 34.292 39.892 34.436 44.348 ; 
        RECT 33.68 39.892 33.788 44.348 ; 
        RECT 28.712 39.746 28.784 44.386 ; 
        RECT 0.632 39.746 0.704 44.386 ; 
        RECT 65.412 44.042 65.484 76.87 ; 
        RECT 37.332 44.042 37.404 76.87 ; 
        RECT 33.516 44.936 34.452 75.668 ; 
        RECT 34.272 44.218 34.416 76.696 ; 
        RECT 33.66 44.216 33.768 76.696 ; 
        RECT 28.692 44.042 28.764 76.87 ; 
        RECT 0.612 44.042 0.684 76.87 ; 
        RECT 65.432 76.574 65.504 81.214 ; 
        RECT 37.352 76.574 37.424 81.214 ; 
        RECT 34.292 76.72 34.436 81.176 ; 
        RECT 33.68 76.72 33.788 81.176 ; 
        RECT 28.712 76.574 28.784 81.214 ; 
        RECT 0.632 76.574 0.704 81.214 ; 
        RECT 65.432 80.894 65.504 85.534 ; 
        RECT 37.352 80.894 37.424 85.534 ; 
        RECT 34.292 81.04 34.436 85.496 ; 
        RECT 33.68 81.04 33.788 85.496 ; 
        RECT 28.712 80.894 28.784 85.534 ; 
        RECT 0.632 80.894 0.704 85.534 ; 
        RECT 65.432 85.214 65.504 89.854 ; 
        RECT 37.352 85.214 37.424 89.854 ; 
        RECT 34.292 85.36 34.436 89.816 ; 
        RECT 33.68 85.36 33.788 89.816 ; 
        RECT 28.712 85.214 28.784 89.854 ; 
        RECT 0.632 85.214 0.704 89.854 ; 
        RECT 65.432 89.534 65.504 94.174 ; 
        RECT 37.352 89.534 37.424 94.174 ; 
        RECT 34.292 89.68 34.436 94.136 ; 
        RECT 33.68 89.68 33.788 94.136 ; 
        RECT 28.712 89.534 28.784 94.174 ; 
        RECT 0.632 89.534 0.704 94.174 ; 
        RECT 65.432 93.854 65.504 98.494 ; 
        RECT 37.352 93.854 37.424 98.494 ; 
        RECT 34.292 94 34.436 98.456 ; 
        RECT 33.68 94 33.788 98.456 ; 
        RECT 28.712 93.854 28.784 98.494 ; 
        RECT 0.632 93.854 0.704 98.494 ; 
        RECT 65.432 98.174 65.504 102.814 ; 
        RECT 37.352 98.174 37.424 102.814 ; 
        RECT 34.292 98.32 34.436 102.776 ; 
        RECT 33.68 98.32 33.788 102.776 ; 
        RECT 28.712 98.174 28.784 102.814 ; 
        RECT 0.632 98.174 0.704 102.814 ; 
        RECT 65.432 102.494 65.504 107.134 ; 
        RECT 37.352 102.494 37.424 107.134 ; 
        RECT 34.292 102.64 34.436 107.096 ; 
        RECT 33.68 102.64 33.788 107.096 ; 
        RECT 28.712 102.494 28.784 107.134 ; 
        RECT 0.632 102.494 0.704 107.134 ; 
        RECT 65.432 106.814 65.504 111.454 ; 
        RECT 37.352 106.814 37.424 111.454 ; 
        RECT 34.292 106.96 34.436 111.416 ; 
        RECT 33.68 106.96 33.788 111.416 ; 
        RECT 28.712 106.814 28.784 111.454 ; 
        RECT 0.632 106.814 0.704 111.454 ; 
        RECT 65.432 111.134 65.504 115.774 ; 
        RECT 37.352 111.134 37.424 115.774 ; 
        RECT 34.292 111.28 34.436 115.736 ; 
        RECT 33.68 111.28 33.788 115.736 ; 
        RECT 28.712 111.134 28.784 115.774 ; 
        RECT 0.632 111.134 0.704 115.774 ; 
        RECT 65.432 115.454 65.504 120.094 ; 
        RECT 37.352 115.454 37.424 120.094 ; 
        RECT 34.292 115.6 34.436 120.056 ; 
        RECT 33.68 115.6 33.788 120.056 ; 
        RECT 28.712 115.454 28.784 120.094 ; 
        RECT 0.632 115.454 0.704 120.094 ; 
      LAYER V3 ; 
        RECT 0.632 4.304 0.704 4.496 ; 
        RECT 28.712 4.304 28.784 4.496 ; 
        RECT 33.68 4.304 33.788 4.496 ; 
        RECT 34.292 4.304 34.436 4.496 ; 
        RECT 37.352 4.304 37.424 4.496 ; 
        RECT 65.432 4.304 65.504 4.496 ; 
        RECT 0.632 8.624 0.704 8.816 ; 
        RECT 28.712 8.624 28.784 8.816 ; 
        RECT 33.68 8.624 33.788 8.816 ; 
        RECT 34.292 8.624 34.436 8.816 ; 
        RECT 37.352 8.624 37.424 8.816 ; 
        RECT 65.432 8.624 65.504 8.816 ; 
        RECT 0.632 12.944 0.704 13.136 ; 
        RECT 28.712 12.944 28.784 13.136 ; 
        RECT 33.68 12.944 33.788 13.136 ; 
        RECT 34.292 12.944 34.436 13.136 ; 
        RECT 37.352 12.944 37.424 13.136 ; 
        RECT 65.432 12.944 65.504 13.136 ; 
        RECT 0.632 17.264 0.704 17.456 ; 
        RECT 28.712 17.264 28.784 17.456 ; 
        RECT 33.68 17.264 33.788 17.456 ; 
        RECT 34.292 17.264 34.436 17.456 ; 
        RECT 37.352 17.264 37.424 17.456 ; 
        RECT 65.432 17.264 65.504 17.456 ; 
        RECT 0.632 21.584 0.704 21.776 ; 
        RECT 28.712 21.584 28.784 21.776 ; 
        RECT 33.68 21.584 33.788 21.776 ; 
        RECT 34.292 21.584 34.436 21.776 ; 
        RECT 37.352 21.584 37.424 21.776 ; 
        RECT 65.432 21.584 65.504 21.776 ; 
        RECT 0.632 25.904 0.704 26.096 ; 
        RECT 28.712 25.904 28.784 26.096 ; 
        RECT 33.68 25.904 33.788 26.096 ; 
        RECT 34.292 25.904 34.436 26.096 ; 
        RECT 37.352 25.904 37.424 26.096 ; 
        RECT 65.432 25.904 65.504 26.096 ; 
        RECT 0.632 30.224 0.704 30.416 ; 
        RECT 28.712 30.224 28.784 30.416 ; 
        RECT 33.68 30.224 33.788 30.416 ; 
        RECT 34.292 30.224 34.436 30.416 ; 
        RECT 37.352 30.224 37.424 30.416 ; 
        RECT 65.432 30.224 65.504 30.416 ; 
        RECT 0.632 34.544 0.704 34.736 ; 
        RECT 28.712 34.544 28.784 34.736 ; 
        RECT 33.68 34.544 33.788 34.736 ; 
        RECT 34.292 34.544 34.436 34.736 ; 
        RECT 37.352 34.544 37.424 34.736 ; 
        RECT 65.432 34.544 65.504 34.736 ; 
        RECT 0.632 38.864 0.704 39.056 ; 
        RECT 28.712 38.864 28.784 39.056 ; 
        RECT 33.68 38.864 33.788 39.056 ; 
        RECT 34.292 38.864 34.436 39.056 ; 
        RECT 37.352 38.864 37.424 39.056 ; 
        RECT 65.432 38.864 65.504 39.056 ; 
        RECT 0.632 43.184 0.704 43.376 ; 
        RECT 28.712 43.184 28.784 43.376 ; 
        RECT 33.68 43.184 33.788 43.376 ; 
        RECT 34.292 43.184 34.436 43.376 ; 
        RECT 37.352 43.184 37.424 43.376 ; 
        RECT 65.432 43.184 65.504 43.376 ; 
        RECT 33.532 72.564 33.604 73.428 ; 
        RECT 33.532 59.892 33.604 60.756 ; 
        RECT 33.532 47.22 33.604 48.084 ; 
        RECT 33.74 72.564 33.812 73.428 ; 
        RECT 33.74 59.892 33.812 60.756 ; 
        RECT 33.74 47.22 33.812 48.084 ; 
        RECT 33.948 72.564 34.02 73.428 ; 
        RECT 33.948 59.892 34.02 60.756 ; 
        RECT 33.948 47.22 34.02 48.084 ; 
        RECT 34.156 72.564 34.228 73.428 ; 
        RECT 34.156 59.892 34.228 60.756 ; 
        RECT 34.156 47.22 34.228 48.084 ; 
        RECT 34.364 72.564 34.436 73.428 ; 
        RECT 34.364 59.892 34.436 60.756 ; 
        RECT 34.364 47.22 34.436 48.084 ; 
        RECT 37.332 47.222 37.404 48.086 ; 
        RECT 0.632 80.012 0.704 80.204 ; 
        RECT 28.712 80.012 28.784 80.204 ; 
        RECT 33.68 80.012 33.788 80.204 ; 
        RECT 34.292 80.012 34.436 80.204 ; 
        RECT 37.352 80.012 37.424 80.204 ; 
        RECT 65.432 80.012 65.504 80.204 ; 
        RECT 0.632 84.332 0.704 84.524 ; 
        RECT 28.712 84.332 28.784 84.524 ; 
        RECT 33.68 84.332 33.788 84.524 ; 
        RECT 34.292 84.332 34.436 84.524 ; 
        RECT 37.352 84.332 37.424 84.524 ; 
        RECT 65.432 84.332 65.504 84.524 ; 
        RECT 0.632 88.652 0.704 88.844 ; 
        RECT 28.712 88.652 28.784 88.844 ; 
        RECT 33.68 88.652 33.788 88.844 ; 
        RECT 34.292 88.652 34.436 88.844 ; 
        RECT 37.352 88.652 37.424 88.844 ; 
        RECT 65.432 88.652 65.504 88.844 ; 
        RECT 0.632 92.972 0.704 93.164 ; 
        RECT 28.712 92.972 28.784 93.164 ; 
        RECT 33.68 92.972 33.788 93.164 ; 
        RECT 34.292 92.972 34.436 93.164 ; 
        RECT 37.352 92.972 37.424 93.164 ; 
        RECT 65.432 92.972 65.504 93.164 ; 
        RECT 0.632 97.292 0.704 97.484 ; 
        RECT 28.712 97.292 28.784 97.484 ; 
        RECT 33.68 97.292 33.788 97.484 ; 
        RECT 34.292 97.292 34.436 97.484 ; 
        RECT 37.352 97.292 37.424 97.484 ; 
        RECT 65.432 97.292 65.504 97.484 ; 
        RECT 0.632 101.612 0.704 101.804 ; 
        RECT 28.712 101.612 28.784 101.804 ; 
        RECT 33.68 101.612 33.788 101.804 ; 
        RECT 34.292 101.612 34.436 101.804 ; 
        RECT 37.352 101.612 37.424 101.804 ; 
        RECT 65.432 101.612 65.504 101.804 ; 
        RECT 0.632 105.932 0.704 106.124 ; 
        RECT 28.712 105.932 28.784 106.124 ; 
        RECT 33.68 105.932 33.788 106.124 ; 
        RECT 34.292 105.932 34.436 106.124 ; 
        RECT 37.352 105.932 37.424 106.124 ; 
        RECT 65.432 105.932 65.504 106.124 ; 
        RECT 0.632 110.252 0.704 110.444 ; 
        RECT 28.712 110.252 28.784 110.444 ; 
        RECT 33.68 110.252 33.788 110.444 ; 
        RECT 34.292 110.252 34.436 110.444 ; 
        RECT 37.352 110.252 37.424 110.444 ; 
        RECT 65.432 110.252 65.504 110.444 ; 
        RECT 0.632 114.572 0.704 114.764 ; 
        RECT 28.712 114.572 28.784 114.764 ; 
        RECT 33.68 114.572 33.788 114.764 ; 
        RECT 34.292 114.572 34.436 114.764 ; 
        RECT 37.352 114.572 37.424 114.764 ; 
        RECT 65.432 114.572 65.504 114.764 ; 
        RECT 0.632 118.892 0.704 119.084 ; 
        RECT 28.712 118.892 28.784 119.084 ; 
        RECT 33.68 118.892 33.788 119.084 ; 
        RECT 34.292 118.892 34.436 119.084 ; 
        RECT 37.352 118.892 37.424 119.084 ; 
        RECT 65.432 118.892 65.504 119.084 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 43.164 49.108 43.236 49.256 ; 
      LAYER M4 ; 
        RECT 42.956 49.14 43.292 49.236 ; 
      LAYER M5 ; 
        RECT 43.152 45.336 43.248 58.296 ; 
      LAYER V3 ; 
        RECT 43.164 49.14 43.236 49.236 ; 
      LAYER V4 ; 
        RECT 43.152 49.14 43.248 49.236 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 42.3 49.12 42.372 49.268 ; 
      LAYER M4 ; 
        RECT 42.092 49.14 42.428 49.236 ; 
      LAYER M5 ; 
        RECT 42.288 45.336 42.384 58.296 ; 
      LAYER V3 ; 
        RECT 42.3 49.14 42.372 49.236 ; 
      LAYER V4 ; 
        RECT 42.288 49.14 42.384 49.236 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 41.436 46.804 41.508 46.952 ; 
      LAYER M4 ; 
        RECT 41.228 46.836 41.564 46.932 ; 
      LAYER M5 ; 
        RECT 41.424 45.336 41.52 58.296 ; 
      LAYER V3 ; 
        RECT 41.436 46.836 41.508 46.932 ; 
      LAYER V4 ; 
        RECT 41.424 46.836 41.52 46.932 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 40.572 47.764 40.644 48.488 ; 
      LAYER M4 ; 
        RECT 40.364 48.372 40.7 48.468 ; 
      LAYER M5 ; 
        RECT 40.56 45.336 40.656 58.296 ; 
      LAYER V3 ; 
        RECT 40.572 48.372 40.644 48.468 ; 
      LAYER V4 ; 
        RECT 40.56 48.372 40.656 48.468 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 39.708 46.816 39.78 47.084 ; 
      LAYER M4 ; 
        RECT 39.5 46.836 39.836 46.932 ; 
      LAYER M5 ; 
        RECT 39.696 45.336 39.792 58.296 ; 
      LAYER V3 ; 
        RECT 39.708 46.836 39.78 46.932 ; 
      LAYER V4 ; 
        RECT 39.696 46.836 39.792 46.932 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 38.844 45.748 38.916 46.76 ; 
      LAYER M4 ; 
        RECT 38.636 46.644 38.972 46.74 ; 
      LAYER M5 ; 
        RECT 38.832 45.336 38.928 58.296 ; 
      LAYER V3 ; 
        RECT 38.844 46.644 38.916 46.74 ; 
      LAYER V4 ; 
        RECT 38.832 46.644 38.928 46.74 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.98 49.888 38.052 50.036 ; 
      LAYER M4 ; 
        RECT 37.772 49.908 38.108 50.004 ; 
      LAYER M5 ; 
        RECT 37.968 45.336 38.064 58.296 ; 
      LAYER V3 ; 
        RECT 37.98 49.908 38.052 50.004 ; 
      LAYER V4 ; 
        RECT 37.968 49.908 38.064 50.004 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.116 49.276 37.188 49.64 ; 
      LAYER M4 ; 
        RECT 36.908 49.524 37.244 49.62 ; 
      LAYER M5 ; 
        RECT 37.104 45.336 37.2 58.296 ; 
      LAYER V3 ; 
        RECT 37.116 49.524 37.188 49.62 ; 
      LAYER V4 ; 
        RECT 37.104 49.524 37.2 49.62 ; 
    END 
  END ADDRESS[7] 
  PIN ADDRESS[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 34.524 46.816 34.596 47.084 ; 
      LAYER M4 ; 
        RECT 33.388 46.836 34.64 46.932 ; 
      LAYER M5 ; 
        RECT 33.432 45.336 33.528 58.296 ; 
      LAYER V3 ; 
        RECT 34.524 46.836 34.596 46.932 ; 
      LAYER V4 ; 
        RECT 33.432 46.836 33.528 46.932 ; 
    END 
  END ADDRESS[8] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 32.94 45.748 33.012 46.76 ; 
      LAYER M4 ; 
        RECT 32.092 46.644 33.056 46.74 ; 
      LAYER M5 ; 
        RECT 32.136 45.336 32.232 58.296 ; 
      LAYER V3 ; 
        RECT 32.94 46.644 33.012 46.74 ; 
      LAYER V4 ; 
        RECT 32.136 46.644 32.232 46.74 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.772 46.816 29.844 47.084 ; 
      LAYER M4 ; 
        RECT 29.564 46.836 29.9 46.932 ; 
      LAYER M5 ; 
        RECT 29.76 45.336 29.856 58.296 ; 
      LAYER V3 ; 
        RECT 29.772 46.836 29.844 46.932 ; 
      LAYER V4 ; 
        RECT 29.76 46.836 29.856 46.932 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.908 50.272 28.98 50.468 ; 
      LAYER M4 ; 
        RECT 28.7 50.292 29.036 50.388 ; 
      LAYER M5 ; 
        RECT 28.896 45.336 28.992 58.296 ; 
      LAYER V3 ; 
        RECT 28.908 50.292 28.98 50.388 ; 
      LAYER V4 ; 
        RECT 28.896 50.292 28.992 50.388 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.052 45.748 29.124 46.76 ; 
      LAYER M4 ; 
        RECT 27.988 46.644 29.168 46.74 ; 
      LAYER M5 ; 
        RECT 28.032 45.336 28.128 58.296 ; 
      LAYER V3 ; 
        RECT 29.052 46.644 29.124 46.74 ; 
      LAYER V4 ; 
        RECT 28.032 46.644 28.128 46.74 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.18 49.108 27.252 49.256 ; 
      LAYER M4 ; 
        RECT 26.972 49.14 27.308 49.236 ; 
      LAYER M5 ; 
        RECT 27.168 45.336 27.264 58.296 ; 
      LAYER V3 ; 
        RECT 27.18 49.14 27.252 49.236 ; 
      LAYER V4 ; 
        RECT 27.168 49.14 27.264 49.236 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.316 46.816 26.388 47.732 ; 
      LAYER M4 ; 
        RECT 26.108 46.836 26.444 46.932 ; 
      LAYER M5 ; 
        RECT 26.304 45.336 26.4 58.296 ; 
      LAYER V3 ; 
        RECT 26.316 46.836 26.388 46.932 ; 
      LAYER V4 ; 
        RECT 26.304 46.836 26.4 46.932 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.452 45.748 25.524 46.76 ; 
      LAYER M4 ; 
        RECT 25.244 46.644 25.58 46.74 ; 
      LAYER M5 ; 
        RECT 25.44 45.336 25.536 58.296 ; 
      LAYER V3 ; 
        RECT 25.452 46.644 25.524 46.74 ; 
      LAYER V4 ; 
        RECT 25.44 46.644 25.536 46.74 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.588 46.804 24.66 46.952 ; 
      LAYER M4 ; 
        RECT 24.38 46.836 24.716 46.932 ; 
      LAYER M5 ; 
        RECT 24.576 45.336 24.672 58.296 ; 
      LAYER V3 ; 
        RECT 24.588 46.836 24.66 46.932 ; 
      LAYER V4 ; 
        RECT 24.576 46.836 24.672 46.932 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 23.724 49.108 23.796 49.256 ; 
      LAYER M4 ; 
        RECT 23.516 49.14 23.852 49.236 ; 
      LAYER M5 ; 
        RECT 23.712 45.336 23.808 58.296 ; 
      LAYER V3 ; 
        RECT 23.724 49.14 23.796 49.236 ; 
      LAYER V4 ; 
        RECT 23.712 49.14 23.808 49.236 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.712 34.388 1.808 ; 
      LAYER M3 ; 
        RECT 34.148 1.51 34.22 2.468 ; 
      LAYER V3 ; 
        RECT 34.148 1.712 34.22 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.328 34.66 1.424 ; 
      LAYER M3 ; 
        RECT 33.248 1.08 33.32 2.7 ; 
      LAYER V3 ; 
        RECT 33.248 1.328 33.32 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 6.032 34.388 6.128 ; 
      LAYER M3 ; 
        RECT 34.148 5.83 34.22 6.788 ; 
      LAYER V3 ; 
        RECT 34.148 6.032 34.22 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 5.648 34.66 5.744 ; 
      LAYER M3 ; 
        RECT 33.248 5.4 33.32 7.02 ; 
      LAYER V3 ; 
        RECT 33.248 5.648 33.32 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 10.352 34.388 10.448 ; 
      LAYER M3 ; 
        RECT 34.148 10.15 34.22 11.108 ; 
      LAYER V3 ; 
        RECT 34.148 10.352 34.22 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 9.968 34.66 10.064 ; 
      LAYER M3 ; 
        RECT 33.248 9.72 33.32 11.34 ; 
      LAYER V3 ; 
        RECT 33.248 9.968 33.32 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.672 34.388 14.768 ; 
      LAYER M3 ; 
        RECT 34.148 14.47 34.22 15.428 ; 
      LAYER V3 ; 
        RECT 34.148 14.672 34.22 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.288 34.66 14.384 ; 
      LAYER M3 ; 
        RECT 33.248 14.04 33.32 15.66 ; 
      LAYER V3 ; 
        RECT 33.248 14.288 33.32 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.992 34.388 19.088 ; 
      LAYER M3 ; 
        RECT 34.148 18.79 34.22 19.748 ; 
      LAYER V3 ; 
        RECT 34.148 18.992 34.22 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.608 34.66 18.704 ; 
      LAYER M3 ; 
        RECT 33.248 18.36 33.32 19.98 ; 
      LAYER V3 ; 
        RECT 33.248 18.608 33.32 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 23.312 34.388 23.408 ; 
      LAYER M3 ; 
        RECT 34.148 23.11 34.22 24.068 ; 
      LAYER V3 ; 
        RECT 34.148 23.312 34.22 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 22.928 34.66 23.024 ; 
      LAYER M3 ; 
        RECT 33.248 22.68 33.32 24.3 ; 
      LAYER V3 ; 
        RECT 33.248 22.928 33.32 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.632 34.388 27.728 ; 
      LAYER M3 ; 
        RECT 34.148 27.43 34.22 28.388 ; 
      LAYER V3 ; 
        RECT 34.148 27.632 34.22 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.248 34.66 27.344 ; 
      LAYER M3 ; 
        RECT 33.248 27 33.32 28.62 ; 
      LAYER V3 ; 
        RECT 33.248 27.248 33.32 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.952 34.388 32.048 ; 
      LAYER M3 ; 
        RECT 34.148 31.75 34.22 32.708 ; 
      LAYER V3 ; 
        RECT 34.148 31.952 34.22 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.568 34.66 31.664 ; 
      LAYER M3 ; 
        RECT 33.248 31.32 33.32 32.94 ; 
      LAYER V3 ; 
        RECT 33.248 31.568 33.32 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 36.272 34.388 36.368 ; 
      LAYER M3 ; 
        RECT 34.148 36.07 34.22 37.028 ; 
      LAYER V3 ; 
        RECT 34.148 36.272 34.22 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 35.888 34.66 35.984 ; 
      LAYER M3 ; 
        RECT 33.248 35.64 33.32 37.26 ; 
      LAYER V3 ; 
        RECT 33.248 35.888 33.32 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.592 34.388 40.688 ; 
      LAYER M3 ; 
        RECT 34.148 40.39 34.22 41.348 ; 
      LAYER V3 ; 
        RECT 34.148 40.592 34.22 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.208 34.66 40.304 ; 
      LAYER M3 ; 
        RECT 33.248 39.96 33.32 41.58 ; 
      LAYER V3 ; 
        RECT 33.248 40.208 33.32 40.304 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 77.42 34.388 77.516 ; 
      LAYER M3 ; 
        RECT 34.148 77.218 34.22 78.176 ; 
      LAYER V3 ; 
        RECT 34.148 77.42 34.22 77.516 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 77.036 34.66 77.132 ; 
      LAYER M3 ; 
        RECT 33.248 76.788 33.32 78.408 ; 
      LAYER V3 ; 
        RECT 33.248 77.036 33.32 77.132 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 81.74 34.388 81.836 ; 
      LAYER M3 ; 
        RECT 34.148 81.538 34.22 82.496 ; 
      LAYER V3 ; 
        RECT 34.148 81.74 34.22 81.836 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 81.356 34.66 81.452 ; 
      LAYER M3 ; 
        RECT 33.248 81.108 33.32 82.728 ; 
      LAYER V3 ; 
        RECT 33.248 81.356 33.32 81.452 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 86.06 34.388 86.156 ; 
      LAYER M3 ; 
        RECT 34.148 85.858 34.22 86.816 ; 
      LAYER V3 ; 
        RECT 34.148 86.06 34.22 86.156 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 85.676 34.66 85.772 ; 
      LAYER M3 ; 
        RECT 33.248 85.428 33.32 87.048 ; 
      LAYER V3 ; 
        RECT 33.248 85.676 33.32 85.772 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 90.38 34.388 90.476 ; 
      LAYER M3 ; 
        RECT 34.148 90.178 34.22 91.136 ; 
      LAYER V3 ; 
        RECT 34.148 90.38 34.22 90.476 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 89.996 34.66 90.092 ; 
      LAYER M3 ; 
        RECT 33.248 89.748 33.32 91.368 ; 
      LAYER V3 ; 
        RECT 33.248 89.996 33.32 90.092 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 94.7 34.388 94.796 ; 
      LAYER M3 ; 
        RECT 34.148 94.498 34.22 95.456 ; 
      LAYER V3 ; 
        RECT 34.148 94.7 34.22 94.796 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 94.316 34.66 94.412 ; 
      LAYER M3 ; 
        RECT 33.248 94.068 33.32 95.688 ; 
      LAYER V3 ; 
        RECT 33.248 94.316 33.32 94.412 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 99.02 34.388 99.116 ; 
      LAYER M3 ; 
        RECT 34.148 98.818 34.22 99.776 ; 
      LAYER V3 ; 
        RECT 34.148 99.02 34.22 99.116 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 98.636 34.66 98.732 ; 
      LAYER M3 ; 
        RECT 33.248 98.388 33.32 100.008 ; 
      LAYER V3 ; 
        RECT 33.248 98.636 33.32 98.732 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 103.34 34.388 103.436 ; 
      LAYER M3 ; 
        RECT 34.148 103.138 34.22 104.096 ; 
      LAYER V3 ; 
        RECT 34.148 103.34 34.22 103.436 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 102.956 34.66 103.052 ; 
      LAYER M3 ; 
        RECT 33.248 102.708 33.32 104.328 ; 
      LAYER V3 ; 
        RECT 33.248 102.956 33.32 103.052 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 107.66 34.388 107.756 ; 
      LAYER M3 ; 
        RECT 34.148 107.458 34.22 108.416 ; 
      LAYER V3 ; 
        RECT 34.148 107.66 34.22 107.756 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 107.276 34.66 107.372 ; 
      LAYER M3 ; 
        RECT 33.248 107.028 33.32 108.648 ; 
      LAYER V3 ; 
        RECT 33.248 107.276 33.32 107.372 ; 
    END 
  END wd[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 111.98 34.388 112.076 ; 
      LAYER M3 ; 
        RECT 34.148 111.778 34.22 112.736 ; 
      LAYER V3 ; 
        RECT 34.148 111.98 34.22 112.076 ; 
    END 
  END dataout[18] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 111.596 34.66 111.692 ; 
      LAYER M3 ; 
        RECT 33.248 111.348 33.32 112.968 ; 
      LAYER V3 ; 
        RECT 33.248 111.596 33.32 111.692 ; 
    END 
  END wd[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 116.3 34.388 116.396 ; 
      LAYER M3 ; 
        RECT 34.148 116.098 34.22 117.056 ; 
      LAYER V3 ; 
        RECT 34.148 116.3 34.22 116.396 ; 
    END 
  END dataout[19] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 115.916 34.66 116.012 ; 
      LAYER M3 ; 
        RECT 33.248 115.668 33.32 117.288 ; 
      LAYER V3 ; 
        RECT 33.248 115.916 33.32 116.012 ; 
    END 
  END wd[19] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0 44.148 66.096 78.762 ; 
        RECT 0.02 76.734 66.116 81.108 ; 
        RECT 0.02 81.054 66.116 85.428 ; 
        RECT 0.02 85.374 66.116 89.748 ; 
        RECT 0.02 89.694 66.116 94.068 ; 
        RECT 0.02 94.014 66.116 98.388 ; 
        RECT 0.02 98.334 66.116 102.708 ; 
        RECT 0.02 102.654 66.116 107.028 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0 44.148 66.096 78.762 ; 
        RECT 0.02 76.734 66.116 81.108 ; 
        RECT 0.02 81.054 66.116 85.428 ; 
        RECT 0.02 85.374 66.116 89.748 ; 
        RECT 0.02 89.694 66.116 94.068 ; 
        RECT 0.02 94.014 66.116 98.388 ; 
        RECT 0.02 98.334 66.116 102.708 ; 
        RECT 0.02 102.654 66.116 107.028 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
  LAYER V1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0 44.148 66.096 78.762 ; 
        RECT 0.02 76.734 66.116 81.108 ; 
        RECT 0.02 81.054 66.116 85.428 ; 
        RECT 0.02 85.374 66.116 89.748 ; 
        RECT 0.02 89.694 66.116 94.068 ; 
        RECT 0.02 94.014 66.116 98.388 ; 
        RECT 0.02 98.334 66.116 102.708 ; 
        RECT 0.02 102.654 66.116 107.028 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
  LAYER V2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0 44.148 66.096 78.762 ; 
        RECT 0.02 76.734 66.116 81.108 ; 
        RECT 0.02 81.054 66.116 85.428 ; 
        RECT 0.02 85.374 66.116 89.748 ; 
        RECT 0.02 89.694 66.116 94.068 ; 
        RECT 0.02 94.014 66.116 98.388 ; 
        RECT 0.02 98.334 66.116 102.708 ; 
        RECT 0.02 102.654 66.116 107.028 ; 
        RECT 0.02 106.974 66.116 111.348 ; 
        RECT 0.02 111.294 66.116 115.668 ; 
        RECT 0.02 115.614 66.116 119.988 ; 
  LAYER M3 ; 
      RECT 34.796 1.38 34.868 5.122 ; 
      RECT 34.652 1.38 34.724 5.122 ; 
      RECT 34.508 3.688 34.58 4.978 ; 
      RECT 34.04 4.476 34.112 4.914 ; 
      RECT 34.004 1.51 34.076 2.468 ; 
      RECT 33.86 3.834 33.932 4.448 ; 
      RECT 33.536 3.936 33.608 4.968 ; 
      RECT 31.376 1.38 31.448 5.122 ; 
      RECT 31.232 1.38 31.304 5.122 ; 
      RECT 31.088 2.104 31.16 4.376 ; 
      RECT 34.796 5.7 34.868 9.442 ; 
      RECT 34.652 5.7 34.724 9.442 ; 
      RECT 34.508 8.008 34.58 9.298 ; 
      RECT 34.04 8.796 34.112 9.234 ; 
      RECT 34.004 5.83 34.076 6.788 ; 
      RECT 33.86 8.154 33.932 8.768 ; 
      RECT 33.536 8.256 33.608 9.288 ; 
      RECT 31.376 5.7 31.448 9.442 ; 
      RECT 31.232 5.7 31.304 9.442 ; 
      RECT 31.088 6.424 31.16 8.696 ; 
      RECT 34.796 10.02 34.868 13.762 ; 
      RECT 34.652 10.02 34.724 13.762 ; 
      RECT 34.508 12.328 34.58 13.618 ; 
      RECT 34.04 13.116 34.112 13.554 ; 
      RECT 34.004 10.15 34.076 11.108 ; 
      RECT 33.86 12.474 33.932 13.088 ; 
      RECT 33.536 12.576 33.608 13.608 ; 
      RECT 31.376 10.02 31.448 13.762 ; 
      RECT 31.232 10.02 31.304 13.762 ; 
      RECT 31.088 10.744 31.16 13.016 ; 
      RECT 34.796 14.34 34.868 18.082 ; 
      RECT 34.652 14.34 34.724 18.082 ; 
      RECT 34.508 16.648 34.58 17.938 ; 
      RECT 34.04 17.436 34.112 17.874 ; 
      RECT 34.004 14.47 34.076 15.428 ; 
      RECT 33.86 16.794 33.932 17.408 ; 
      RECT 33.536 16.896 33.608 17.928 ; 
      RECT 31.376 14.34 31.448 18.082 ; 
      RECT 31.232 14.34 31.304 18.082 ; 
      RECT 31.088 15.064 31.16 17.336 ; 
      RECT 34.796 18.66 34.868 22.402 ; 
      RECT 34.652 18.66 34.724 22.402 ; 
      RECT 34.508 20.968 34.58 22.258 ; 
      RECT 34.04 21.756 34.112 22.194 ; 
      RECT 34.004 18.79 34.076 19.748 ; 
      RECT 33.86 21.114 33.932 21.728 ; 
      RECT 33.536 21.216 33.608 22.248 ; 
      RECT 31.376 18.66 31.448 22.402 ; 
      RECT 31.232 18.66 31.304 22.402 ; 
      RECT 31.088 19.384 31.16 21.656 ; 
      RECT 34.796 22.98 34.868 26.722 ; 
      RECT 34.652 22.98 34.724 26.722 ; 
      RECT 34.508 25.288 34.58 26.578 ; 
      RECT 34.04 26.076 34.112 26.514 ; 
      RECT 34.004 23.11 34.076 24.068 ; 
      RECT 33.86 25.434 33.932 26.048 ; 
      RECT 33.536 25.536 33.608 26.568 ; 
      RECT 31.376 22.98 31.448 26.722 ; 
      RECT 31.232 22.98 31.304 26.722 ; 
      RECT 31.088 23.704 31.16 25.976 ; 
      RECT 34.796 27.3 34.868 31.042 ; 
      RECT 34.652 27.3 34.724 31.042 ; 
      RECT 34.508 29.608 34.58 30.898 ; 
      RECT 34.04 30.396 34.112 30.834 ; 
      RECT 34.004 27.43 34.076 28.388 ; 
      RECT 33.86 29.754 33.932 30.368 ; 
      RECT 33.536 29.856 33.608 30.888 ; 
      RECT 31.376 27.3 31.448 31.042 ; 
      RECT 31.232 27.3 31.304 31.042 ; 
      RECT 31.088 28.024 31.16 30.296 ; 
      RECT 34.796 31.62 34.868 35.362 ; 
      RECT 34.652 31.62 34.724 35.362 ; 
      RECT 34.508 33.928 34.58 35.218 ; 
      RECT 34.04 34.716 34.112 35.154 ; 
      RECT 34.004 31.75 34.076 32.708 ; 
      RECT 33.86 34.074 33.932 34.688 ; 
      RECT 33.536 34.176 33.608 35.208 ; 
      RECT 31.376 31.62 31.448 35.362 ; 
      RECT 31.232 31.62 31.304 35.362 ; 
      RECT 31.088 32.344 31.16 34.616 ; 
      RECT 34.796 35.94 34.868 39.682 ; 
      RECT 34.652 35.94 34.724 39.682 ; 
      RECT 34.508 38.248 34.58 39.538 ; 
      RECT 34.04 39.036 34.112 39.474 ; 
      RECT 34.004 36.07 34.076 37.028 ; 
      RECT 33.86 38.394 33.932 39.008 ; 
      RECT 33.536 38.496 33.608 39.528 ; 
      RECT 31.376 35.94 31.448 39.682 ; 
      RECT 31.232 35.94 31.304 39.682 ; 
      RECT 31.088 36.664 31.16 38.936 ; 
      RECT 34.796 40.26 34.868 44.002 ; 
      RECT 34.652 40.26 34.724 44.002 ; 
      RECT 34.508 42.568 34.58 43.858 ; 
      RECT 34.04 43.356 34.112 43.794 ; 
      RECT 34.004 40.39 34.076 41.348 ; 
      RECT 33.86 42.714 33.932 43.328 ; 
      RECT 33.536 42.816 33.608 43.848 ; 
      RECT 31.376 40.26 31.448 44.002 ; 
      RECT 31.232 40.26 31.304 44.002 ; 
      RECT 31.088 40.984 31.16 43.256 ; 
      RECT 65.268 59.32 65.34 76.736 ; 
      RECT 65.124 54.06 65.196 54.336 ; 
      RECT 65.124 60.54 65.196 60.872 ; 
      RECT 64.98 44.042 65.052 76.87 ; 
      RECT 64.836 59.45 64.908 62.21 ; 
      RECT 64.836 62.414 64.908 66.36 ; 
      RECT 64.836 66.52 64.908 68.988 ; 
      RECT 64.692 59.196 64.764 62.0152 ; 
      RECT 64.692 65.028 64.764 69.708 ; 
      RECT 64.548 44.042 64.62 58.428 ; 
      RECT 64.116 44.042 64.188 58.428 ; 
      RECT 63.684 44.042 63.756 58.428 ; 
      RECT 63.252 44.042 63.324 58.428 ; 
      RECT 62.82 44.042 62.892 58.428 ; 
      RECT 62.388 44.042 62.46 58.428 ; 
      RECT 61.956 44.042 62.028 58.428 ; 
      RECT 61.524 44.042 61.596 58.428 ; 
      RECT 61.092 44.042 61.164 58.428 ; 
      RECT 60.66 44.042 60.732 58.428 ; 
      RECT 60.228 44.042 60.3 58.428 ; 
      RECT 59.796 44.042 59.868 58.428 ; 
      RECT 59.364 44.042 59.436 58.428 ; 
      RECT 58.932 44.042 59.004 58.428 ; 
      RECT 58.5 44.042 58.572 58.428 ; 
      RECT 58.068 44.042 58.14 58.428 ; 
      RECT 57.636 44.042 57.708 58.428 ; 
      RECT 57.204 44.042 57.276 58.428 ; 
      RECT 56.772 44.042 56.844 58.428 ; 
      RECT 56.34 44.042 56.412 58.428 ; 
      RECT 55.908 44.042 55.98 58.428 ; 
      RECT 55.476 44.042 55.548 58.428 ; 
      RECT 55.044 44.042 55.116 58.428 ; 
      RECT 54.612 44.042 54.684 58.428 ; 
      RECT 54.18 44.042 54.252 58.428 ; 
      RECT 53.748 44.042 53.82 58.428 ; 
      RECT 53.316 44.042 53.388 58.428 ; 
      RECT 52.884 44.042 52.956 58.428 ; 
      RECT 52.452 44.042 52.524 58.428 ; 
      RECT 52.02 44.042 52.092 58.428 ; 
      RECT 51.588 44.042 51.66 58.428 ; 
      RECT 51.156 44.042 51.228 58.428 ; 
      RECT 50.724 44.042 50.796 58.428 ; 
      RECT 50.292 44.042 50.364 58.428 ; 
      RECT 49.86 44.042 49.932 58.428 ; 
      RECT 49.428 44.042 49.5 58.428 ; 
      RECT 48.996 44.042 49.068 58.428 ; 
      RECT 48.564 44.042 48.636 58.428 ; 
      RECT 48.132 44.042 48.204 58.428 ; 
      RECT 47.7 44.042 47.772 58.428 ; 
      RECT 47.268 44.042 47.34 58.428 ; 
      RECT 46.836 44.042 46.908 58.428 ; 
      RECT 46.404 44.042 46.476 58.428 ; 
      RECT 45.972 44.042 46.044 58.428 ; 
      RECT 45.54 44.042 45.612 58.428 ; 
      RECT 45.108 44.042 45.18 58.428 ; 
      RECT 44.676 44.042 44.748 58.428 ; 
      RECT 44.244 44.042 44.316 58.428 ; 
      RECT 43.812 44.042 43.884 58.428 ; 
      RECT 43.38 44.042 43.452 58.428 ; 
      RECT 42.948 44.042 43.02 58.428 ; 
      RECT 42.516 44.042 42.588 58.428 ; 
      RECT 42.084 44.042 42.156 58.428 ; 
      RECT 41.652 44.042 41.724 58.428 ; 
      RECT 41.22 44.042 41.292 58.428 ; 
      RECT 40.788 44.042 40.86 58.428 ; 
      RECT 40.356 44.042 40.428 58.428 ; 
      RECT 39.924 44.042 39.996 58.428 ; 
      RECT 39.492 44.042 39.564 58.428 ; 
      RECT 39.06 44.042 39.132 58.428 ; 
      RECT 38.628 44.042 38.7 58.428 ; 
      RECT 38.196 44.042 38.268 58.428 ; 
      RECT 38.052 59.462 38.124 62.03 ; 
      RECT 38.052 64.74 38.124 66.868 ; 
      RECT 37.98 46.684 38.052 49.388 ; 
      RECT 37.98 52.372 38.052 53.564 ; 
      RECT 37.98 56.836 38.052 57.884 ; 
      RECT 37.908 59.12 37.98 62.21 ; 
      RECT 37.908 62.4148 37.98 64.38 ; 
      RECT 37.908 64.56 37.98 66.044 ; 
      RECT 37.908 66.348 37.98 68.988 ; 
      RECT 37.764 44.042 37.836 76.87 ; 
      RECT 37.62 61.292 37.692 63.15 ; 
      RECT 37.548 47.116 37.62 49.64 ; 
      RECT 37.548 51.292 37.62 52.052 ; 
      RECT 37.548 54.82 37.62 55.016 ; 
      RECT 37.548 57.748 37.62 57.896 ; 
      RECT 37.476 59.32 37.548 76.718 ; 
      RECT 37.116 45.604 37.188 48.812 ; 
      RECT 37.116 51.004 37.188 53.276 ; 
      RECT 36.972 51.292 37.044 52.772 ; 
      RECT 36.828 48.7 36.9 49.244 ; 
      RECT 36.828 52.66 36.9 53.564 ; 
      RECT 36.828 57.628 36.9 57.884 ; 
      RECT 36.684 49.108 36.756 49.256 ; 
      RECT 36.684 55.612 36.756 55.784 ; 
      RECT 36.684 57.748 36.756 57.896 ; 
      RECT 36.54 50.356 36.612 52.34 ; 
      RECT 36.54 52.516 36.612 53.276 ; 
      RECT 36.54 56.356 36.612 57.596 ; 
      RECT 36.396 49.924 36.468 54.912 ; 
      RECT 36.396 65.476 36.468 68.396 ; 
      RECT 36.396 69.796 36.468 72.716 ; 
      RECT 35.1 48.844 35.172 50.036 ; 
      RECT 35.1 53.596 35.172 53.852 ; 
      RECT 35.1 54.676 35.172 56.516 ; 
      RECT 35.1 59.476 35.172 59.624 ; 
      RECT 35.1 67.636 35.172 68.828 ; 
      RECT 34.956 49.132 35.028 51.152 ; 
      RECT 34.956 52.228 35.028 55.436 ; 
      RECT 34.956 59.608 35.028 60.692 ; 
      RECT 34.956 61.012 35.028 61.916 ; 
      RECT 34.812 48.844 34.884 51.548 ; 
      RECT 34.812 51.94 34.884 53.276 ; 
      RECT 34.812 54.1 34.884 54.644 ; 
      RECT 34.812 56.836 34.884 60.044 ; 
      RECT 34.812 61.78 34.884 61.928 ; 
      RECT 34.812 70.444 34.884 71.78 ; 
      RECT 34.668 49.78 34.74 50.324 ; 
      RECT 34.668 57.34 34.74 61.268 ; 
      RECT 34.668 63.028 34.74 64.22 ; 
      RECT 34.668 69.796 34.74 70.844 ; 
      RECT 34.524 46.036 34.596 46.652 ; 
      RECT 34.524 49.276 34.596 56.42 ; 
      RECT 34.524 60.58 34.596 69.908 ; 
      RECT 34.524 70.732 34.596 75.164 ; 
      RECT 33.372 47.116 33.444 48.164 ; 
      RECT 33.372 48.7 33.444 48.956 ; 
      RECT 33.372 49.276 33.444 50.18 ; 
      RECT 33.372 50.356 33.444 51.116 ; 
      RECT 33.372 51.436 33.444 61.916 ; 
      RECT 33.372 62.092 33.444 67.316 ; 
      RECT 33.372 71.668 33.444 72.716 ; 
      RECT 33.228 51.112 33.3 52.196 ; 
      RECT 33.228 52.516 33.3 55.868 ; 
      RECT 33.228 56.548 33.3 59.9 ; 
      RECT 33.228 60.076 33.3 65.156 ; 
      RECT 33.228 65.98 33.3 66.668 ; 
      RECT 33.228 69.508 33.3 73.796 ; 
      RECT 33.084 51.436 33.156 52.52 ; 
      RECT 33.084 53.14 33.156 53.288 ; 
      RECT 33.084 56.26 33.156 60.188 ; 
      RECT 33.084 61.156 33.156 62.996 ; 
      RECT 33.084 64.396 33.156 67.352 ; 
      RECT 32.94 47.908 33.012 52.196 ; 
      RECT 32.94 58.564 33.012 59.432 ; 
      RECT 32.94 64.108 33.012 65.3 ; 
      RECT 32.796 50.5 32.868 52.34 ; 
      RECT 32.796 56.836 32.868 57.596 ; 
      RECT 32.796 57.76 32.868 57.908 ; 
      RECT 32.796 58.852 32.868 60.188 ; 
      RECT 32.796 60.724 32.868 66.092 ; 
      RECT 32.796 66.52 32.868 70.988 ; 
      RECT 32.652 48.196 32.724 48.956 ; 
      RECT 32.652 49.78 32.724 50.324 ; 
      RECT 32.652 51.436 32.724 64.076 ; 
      RECT 32.652 64.396 32.724 66.236 ; 
      RECT 32.652 68.716 32.724 70.556 ; 
      RECT 32.652 73.972 32.724 74.876 ; 
      RECT 32.508 44.148 32.58 44.764 ; 
      RECT 32.508 76.128 32.58 76.792 ; 
      RECT 32.364 44.148 32.436 44.348 ; 
      RECT 32.076 44.148 32.148 44.434 ; 
      RECT 32.076 76.406 32.148 76.87 ; 
      RECT 31.5 50.212 31.572 50.972 ; 
      RECT 31.5 53.164 31.572 54.644 ; 
      RECT 31.5 61.012 31.572 61.916 ; 
      RECT 31.5 63.172 31.572 67.748 ; 
      RECT 31.5 70.876 31.572 72.716 ; 
      RECT 31.5 75.028 31.572 75.176 ; 
      RECT 31.356 46.036 31.428 48.02 ; 
      RECT 31.356 62.356 31.428 62.504 ; 
      RECT 31.356 66.664 31.428 69.908 ; 
      RECT 31.212 47.908 31.284 48.956 ; 
      RECT 31.212 50.068 31.284 51.404 ; 
      RECT 31.212 52.228 31.284 52.628 ; 
      RECT 31.212 55.756 31.284 66.812 ; 
      RECT 31.212 67.348 31.284 68.252 ; 
      RECT 31.068 46.54 31.14 51.116 ; 
      RECT 31.068 65.476 31.14 66.236 ; 
      RECT 31.068 68.692 31.14 68.84 ; 
      RECT 31.068 69.796 31.14 73.004 ; 
      RECT 30.924 50.356 30.996 54.356 ; 
      RECT 30.924 68.116 30.996 68.264 ; 
      RECT 29.484 48.7 29.556 50.324 ; 
      RECT 29.196 48.844 29.268 51.26 ; 
      RECT 29.052 48.196 29.124 48.452 ; 
      RECT 28.908 44.36 28.98 44.564 ; 
      RECT 28.908 56.836 28.98 57.596 ; 
      RECT 28.836 59.32 28.908 76.714 ; 
      RECT 28.548 59.32 28.62 76.718 ; 
      RECT 28.476 46.036 28.548 46.796 ; 
      RECT 28.476 49.132 28.548 58.172 ; 
      RECT 28.404 61.292 28.476 63.15 ; 
      RECT 28.26 44.042 28.332 76.87 ; 
      RECT 28.116 59.12 28.188 62.21 ; 
      RECT 28.116 62.4148 28.188 64.38 ; 
      RECT 28.116 64.56 28.188 66.044 ; 
      RECT 28.116 66.348 28.188 68.988 ; 
      RECT 28.044 46.036 28.116 48.02 ; 
      RECT 28.044 51.148 28.116 53.42 ; 
      RECT 28.044 54.676 28.116 57.596 ; 
      RECT 27.972 59.462 28.044 62.03 ; 
      RECT 27.972 64.74 28.044 66.868 ; 
      RECT 27.828 44.042 27.9 58.428 ; 
      RECT 27.396 44.042 27.468 58.428 ; 
      RECT 26.964 44.042 27.036 58.428 ; 
      RECT 26.532 44.042 26.604 58.428 ; 
      RECT 26.1 44.042 26.172 58.428 ; 
      RECT 25.668 44.042 25.74 58.428 ; 
      RECT 25.236 44.042 25.308 58.428 ; 
      RECT 24.804 44.042 24.876 58.428 ; 
      RECT 24.372 44.042 24.444 58.428 ; 
      RECT 23.94 44.042 24.012 58.428 ; 
      RECT 23.508 44.042 23.58 58.428 ; 
      RECT 23.076 44.042 23.148 58.428 ; 
      RECT 22.644 44.042 22.716 58.428 ; 
      RECT 22.212 44.042 22.284 58.428 ; 
      RECT 21.78 44.042 21.852 58.428 ; 
      RECT 21.348 44.042 21.42 58.428 ; 
      RECT 20.916 44.042 20.988 58.428 ; 
      RECT 20.484 44.042 20.556 58.428 ; 
      RECT 20.052 44.042 20.124 58.428 ; 
      RECT 19.62 44.042 19.692 58.428 ; 
      RECT 19.188 44.042 19.26 58.428 ; 
      RECT 18.756 44.042 18.828 58.428 ; 
      RECT 18.324 44.042 18.396 58.428 ; 
      RECT 17.892 44.042 17.964 58.428 ; 
      RECT 17.46 44.042 17.532 58.428 ; 
      RECT 17.028 44.042 17.1 58.428 ; 
      RECT 16.596 44.042 16.668 58.428 ; 
      RECT 16.164 44.042 16.236 58.428 ; 
      RECT 15.732 44.042 15.804 58.428 ; 
      RECT 15.3 44.042 15.372 58.428 ; 
      RECT 14.868 44.042 14.94 58.428 ; 
      RECT 14.436 44.042 14.508 58.428 ; 
      RECT 14.004 44.042 14.076 58.428 ; 
      RECT 13.572 44.042 13.644 58.428 ; 
      RECT 13.14 44.042 13.212 58.428 ; 
      RECT 12.708 44.042 12.78 58.428 ; 
      RECT 12.276 44.042 12.348 58.428 ; 
      RECT 11.844 44.042 11.916 58.428 ; 
      RECT 11.412 44.042 11.484 58.428 ; 
      RECT 10.98 44.042 11.052 58.428 ; 
      RECT 10.548 44.042 10.62 58.428 ; 
      RECT 10.116 44.042 10.188 58.428 ; 
      RECT 9.684 44.042 9.756 58.428 ; 
      RECT 9.252 44.042 9.324 58.428 ; 
      RECT 8.82 44.042 8.892 58.428 ; 
      RECT 8.388 44.042 8.46 58.428 ; 
      RECT 7.956 44.042 8.028 58.428 ; 
      RECT 7.524 44.042 7.596 58.428 ; 
      RECT 7.092 44.042 7.164 58.428 ; 
      RECT 6.66 44.042 6.732 58.428 ; 
      RECT 6.228 44.042 6.3 58.428 ; 
      RECT 5.796 44.042 5.868 58.428 ; 
      RECT 5.364 44.042 5.436 58.428 ; 
      RECT 4.932 44.042 5.004 58.428 ; 
      RECT 4.5 44.042 4.572 58.428 ; 
      RECT 4.068 44.042 4.14 58.428 ; 
      RECT 3.636 44.042 3.708 58.428 ; 
      RECT 3.204 44.042 3.276 58.428 ; 
      RECT 2.772 44.042 2.844 58.428 ; 
      RECT 2.34 44.042 2.412 58.428 ; 
      RECT 1.908 44.042 1.98 58.428 ; 
      RECT 1.476 44.042 1.548 58.428 ; 
      RECT 1.332 59.196 1.404 62.0152 ; 
      RECT 1.332 65.028 1.404 69.708 ; 
      RECT 1.188 59.45 1.26 62.21 ; 
      RECT 1.188 62.414 1.26 66.36 ; 
      RECT 1.188 66.52 1.26 68.988 ; 
      RECT 1.044 44.042 1.116 76.87 ; 
      RECT 0.9 54.06 0.972 54.336 ; 
      RECT 0.9 60.54 0.972 60.872 ; 
      RECT 0.756 59.32 0.828 76.736 ; 
        RECT 34.796 77.088 34.868 80.83 ; 
        RECT 34.652 77.088 34.724 80.83 ; 
        RECT 34.508 79.396 34.58 80.686 ; 
        RECT 34.04 80.184 34.112 80.622 ; 
        RECT 34.004 77.218 34.076 78.176 ; 
        RECT 33.86 79.542 33.932 80.156 ; 
        RECT 33.536 79.644 33.608 80.676 ; 
        RECT 31.376 77.088 31.448 80.83 ; 
        RECT 31.232 77.088 31.304 80.83 ; 
        RECT 31.088 77.812 31.16 80.084 ; 
        RECT 34.796 81.408 34.868 85.15 ; 
        RECT 34.652 81.408 34.724 85.15 ; 
        RECT 34.508 83.716 34.58 85.006 ; 
        RECT 34.04 84.504 34.112 84.942 ; 
        RECT 34.004 81.538 34.076 82.496 ; 
        RECT 33.86 83.862 33.932 84.476 ; 
        RECT 33.536 83.964 33.608 84.996 ; 
        RECT 31.376 81.408 31.448 85.15 ; 
        RECT 31.232 81.408 31.304 85.15 ; 
        RECT 31.088 82.132 31.16 84.404 ; 
        RECT 34.796 85.728 34.868 89.47 ; 
        RECT 34.652 85.728 34.724 89.47 ; 
        RECT 34.508 88.036 34.58 89.326 ; 
        RECT 34.04 88.824 34.112 89.262 ; 
        RECT 34.004 85.858 34.076 86.816 ; 
        RECT 33.86 88.182 33.932 88.796 ; 
        RECT 33.536 88.284 33.608 89.316 ; 
        RECT 31.376 85.728 31.448 89.47 ; 
        RECT 31.232 85.728 31.304 89.47 ; 
        RECT 31.088 86.452 31.16 88.724 ; 
        RECT 34.796 90.048 34.868 93.79 ; 
        RECT 34.652 90.048 34.724 93.79 ; 
        RECT 34.508 92.356 34.58 93.646 ; 
        RECT 34.04 93.144 34.112 93.582 ; 
        RECT 34.004 90.178 34.076 91.136 ; 
        RECT 33.86 92.502 33.932 93.116 ; 
        RECT 33.536 92.604 33.608 93.636 ; 
        RECT 31.376 90.048 31.448 93.79 ; 
        RECT 31.232 90.048 31.304 93.79 ; 
        RECT 31.088 90.772 31.16 93.044 ; 
        RECT 34.796 94.368 34.868 98.11 ; 
        RECT 34.652 94.368 34.724 98.11 ; 
        RECT 34.508 96.676 34.58 97.966 ; 
        RECT 34.04 97.464 34.112 97.902 ; 
        RECT 34.004 94.498 34.076 95.456 ; 
        RECT 33.86 96.822 33.932 97.436 ; 
        RECT 33.536 96.924 33.608 97.956 ; 
        RECT 31.376 94.368 31.448 98.11 ; 
        RECT 31.232 94.368 31.304 98.11 ; 
        RECT 31.088 95.092 31.16 97.364 ; 
        RECT 34.796 98.688 34.868 102.43 ; 
        RECT 34.652 98.688 34.724 102.43 ; 
        RECT 34.508 100.996 34.58 102.286 ; 
        RECT 34.04 101.784 34.112 102.222 ; 
        RECT 34.004 98.818 34.076 99.776 ; 
        RECT 33.86 101.142 33.932 101.756 ; 
        RECT 33.536 101.244 33.608 102.276 ; 
        RECT 31.376 98.688 31.448 102.43 ; 
        RECT 31.232 98.688 31.304 102.43 ; 
        RECT 31.088 99.412 31.16 101.684 ; 
        RECT 34.796 103.008 34.868 106.75 ; 
        RECT 34.652 103.008 34.724 106.75 ; 
        RECT 34.508 105.316 34.58 106.606 ; 
        RECT 34.04 106.104 34.112 106.542 ; 
        RECT 34.004 103.138 34.076 104.096 ; 
        RECT 33.86 105.462 33.932 106.076 ; 
        RECT 33.536 105.564 33.608 106.596 ; 
        RECT 31.376 103.008 31.448 106.75 ; 
        RECT 31.232 103.008 31.304 106.75 ; 
        RECT 31.088 103.732 31.16 106.004 ; 
        RECT 34.796 107.328 34.868 111.07 ; 
        RECT 34.652 107.328 34.724 111.07 ; 
        RECT 34.508 109.636 34.58 110.926 ; 
        RECT 34.04 110.424 34.112 110.862 ; 
        RECT 34.004 107.458 34.076 108.416 ; 
        RECT 33.86 109.782 33.932 110.396 ; 
        RECT 33.536 109.884 33.608 110.916 ; 
        RECT 31.376 107.328 31.448 111.07 ; 
        RECT 31.232 107.328 31.304 111.07 ; 
        RECT 31.088 108.052 31.16 110.324 ; 
        RECT 34.796 111.648 34.868 115.39 ; 
        RECT 34.652 111.648 34.724 115.39 ; 
        RECT 34.508 113.956 34.58 115.246 ; 
        RECT 34.04 114.744 34.112 115.182 ; 
        RECT 34.004 111.778 34.076 112.736 ; 
        RECT 33.86 114.102 33.932 114.716 ; 
        RECT 33.536 114.204 33.608 115.236 ; 
        RECT 31.376 111.648 31.448 115.39 ; 
        RECT 31.232 111.648 31.304 115.39 ; 
        RECT 31.088 112.372 31.16 114.644 ; 
        RECT 34.796 115.968 34.868 119.71 ; 
        RECT 34.652 115.968 34.724 119.71 ; 
        RECT 34.508 118.276 34.58 119.566 ; 
        RECT 34.04 119.064 34.112 119.502 ; 
        RECT 34.004 116.098 34.076 117.056 ; 
        RECT 33.86 118.422 33.932 119.036 ; 
        RECT 33.536 118.524 33.608 119.556 ; 
        RECT 31.376 115.968 31.448 119.71 ; 
        RECT 31.232 115.968 31.304 119.71 ; 
        RECT 31.088 116.692 31.16 118.964 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 34.564 1.026 35.076 5.4 ; 
      RECT 34.508 3.688 35.076 4.978 ; 
      RECT 33.916 2.596 34.164 5.4 ; 
      RECT 33.86 3.834 34.164 4.448 ; 
      RECT 33.916 1.026 34.02 5.4 ; 
      RECT 33.916 1.51 34.076 2.468 ; 
      RECT 33.916 1.026 34.164 1.382 ; 
      RECT 32.728 2.828 33.552 5.4 ; 
      RECT 33.448 1.026 33.552 5.4 ; 
      RECT 32.728 3.936 33.608 4.968 ; 
      RECT 32.728 1.026 33.12 5.4 ; 
      RECT 31.06 1.026 31.392 5.4 ; 
      RECT 31.06 1.38 31.448 5.122 ; 
      RECT 65.776 1.026 66.116 5.4 ; 
      RECT 65.2 1.026 65.304 5.4 ; 
      RECT 64.768 1.026 64.872 5.4 ; 
      RECT 64.336 1.026 64.44 5.4 ; 
      RECT 63.904 1.026 64.008 5.4 ; 
      RECT 63.472 1.026 63.576 5.4 ; 
      RECT 63.04 1.026 63.144 5.4 ; 
      RECT 62.608 1.026 62.712 5.4 ; 
      RECT 62.176 1.026 62.28 5.4 ; 
      RECT 61.744 1.026 61.848 5.4 ; 
      RECT 61.312 1.026 61.416 5.4 ; 
      RECT 60.88 1.026 60.984 5.4 ; 
      RECT 60.448 1.026 60.552 5.4 ; 
      RECT 60.016 1.026 60.12 5.4 ; 
      RECT 59.584 1.026 59.688 5.4 ; 
      RECT 59.152 1.026 59.256 5.4 ; 
      RECT 58.72 1.026 58.824 5.4 ; 
      RECT 58.288 1.026 58.392 5.4 ; 
      RECT 57.856 1.026 57.96 5.4 ; 
      RECT 57.424 1.026 57.528 5.4 ; 
      RECT 56.992 1.026 57.096 5.4 ; 
      RECT 56.56 1.026 56.664 5.4 ; 
      RECT 56.128 1.026 56.232 5.4 ; 
      RECT 55.696 1.026 55.8 5.4 ; 
      RECT 55.264 1.026 55.368 5.4 ; 
      RECT 54.832 1.026 54.936 5.4 ; 
      RECT 54.4 1.026 54.504 5.4 ; 
      RECT 53.968 1.026 54.072 5.4 ; 
      RECT 53.536 1.026 53.64 5.4 ; 
      RECT 53.104 1.026 53.208 5.4 ; 
      RECT 52.672 1.026 52.776 5.4 ; 
      RECT 52.24 1.026 52.344 5.4 ; 
      RECT 51.808 1.026 51.912 5.4 ; 
      RECT 51.376 1.026 51.48 5.4 ; 
      RECT 50.944 1.026 51.048 5.4 ; 
      RECT 50.512 1.026 50.616 5.4 ; 
      RECT 50.08 1.026 50.184 5.4 ; 
      RECT 49.648 1.026 49.752 5.4 ; 
      RECT 49.216 1.026 49.32 5.4 ; 
      RECT 48.784 1.026 48.888 5.4 ; 
      RECT 48.352 1.026 48.456 5.4 ; 
      RECT 47.92 1.026 48.024 5.4 ; 
      RECT 47.488 1.026 47.592 5.4 ; 
      RECT 47.056 1.026 47.16 5.4 ; 
      RECT 46.624 1.026 46.728 5.4 ; 
      RECT 46.192 1.026 46.296 5.4 ; 
      RECT 45.76 1.026 45.864 5.4 ; 
      RECT 45.328 1.026 45.432 5.4 ; 
      RECT 44.896 1.026 45 5.4 ; 
      RECT 44.464 1.026 44.568 5.4 ; 
      RECT 44.032 1.026 44.136 5.4 ; 
      RECT 43.6 1.026 43.704 5.4 ; 
      RECT 43.168 1.026 43.272 5.4 ; 
      RECT 42.736 1.026 42.84 5.4 ; 
      RECT 42.304 1.026 42.408 5.4 ; 
      RECT 41.872 1.026 41.976 5.4 ; 
      RECT 41.44 1.026 41.544 5.4 ; 
      RECT 41.008 1.026 41.112 5.4 ; 
      RECT 40.576 1.026 40.68 5.4 ; 
      RECT 40.144 1.026 40.248 5.4 ; 
      RECT 39.712 1.026 39.816 5.4 ; 
      RECT 39.28 1.026 39.384 5.4 ; 
      RECT 38.848 1.026 38.952 5.4 ; 
      RECT 38.416 1.026 38.52 5.4 ; 
      RECT 37.984 1.026 38.088 5.4 ; 
      RECT 37.552 1.026 37.656 5.4 ; 
      RECT 36.7 1.026 37.008 5.4 ; 
      RECT 29.128 1.026 29.436 5.4 ; 
      RECT 28.48 1.026 28.584 5.4 ; 
      RECT 28.048 1.026 28.152 5.4 ; 
      RECT 27.616 1.026 27.72 5.4 ; 
      RECT 27.184 1.026 27.288 5.4 ; 
      RECT 26.752 1.026 26.856 5.4 ; 
      RECT 26.32 1.026 26.424 5.4 ; 
      RECT 25.888 1.026 25.992 5.4 ; 
      RECT 25.456 1.026 25.56 5.4 ; 
      RECT 25.024 1.026 25.128 5.4 ; 
      RECT 24.592 1.026 24.696 5.4 ; 
      RECT 24.16 1.026 24.264 5.4 ; 
      RECT 23.728 1.026 23.832 5.4 ; 
      RECT 23.296 1.026 23.4 5.4 ; 
      RECT 22.864 1.026 22.968 5.4 ; 
      RECT 22.432 1.026 22.536 5.4 ; 
      RECT 22 1.026 22.104 5.4 ; 
      RECT 21.568 1.026 21.672 5.4 ; 
      RECT 21.136 1.026 21.24 5.4 ; 
      RECT 20.704 1.026 20.808 5.4 ; 
      RECT 20.272 1.026 20.376 5.4 ; 
      RECT 19.84 1.026 19.944 5.4 ; 
      RECT 19.408 1.026 19.512 5.4 ; 
      RECT 18.976 1.026 19.08 5.4 ; 
      RECT 18.544 1.026 18.648 5.4 ; 
      RECT 18.112 1.026 18.216 5.4 ; 
      RECT 17.68 1.026 17.784 5.4 ; 
      RECT 17.248 1.026 17.352 5.4 ; 
      RECT 16.816 1.026 16.92 5.4 ; 
      RECT 16.384 1.026 16.488 5.4 ; 
      RECT 15.952 1.026 16.056 5.4 ; 
      RECT 15.52 1.026 15.624 5.4 ; 
      RECT 15.088 1.026 15.192 5.4 ; 
      RECT 14.656 1.026 14.76 5.4 ; 
      RECT 14.224 1.026 14.328 5.4 ; 
      RECT 13.792 1.026 13.896 5.4 ; 
      RECT 13.36 1.026 13.464 5.4 ; 
      RECT 12.928 1.026 13.032 5.4 ; 
      RECT 12.496 1.026 12.6 5.4 ; 
      RECT 12.064 1.026 12.168 5.4 ; 
      RECT 11.632 1.026 11.736 5.4 ; 
      RECT 11.2 1.026 11.304 5.4 ; 
      RECT 10.768 1.026 10.872 5.4 ; 
      RECT 10.336 1.026 10.44 5.4 ; 
      RECT 9.904 1.026 10.008 5.4 ; 
      RECT 9.472 1.026 9.576 5.4 ; 
      RECT 9.04 1.026 9.144 5.4 ; 
      RECT 8.608 1.026 8.712 5.4 ; 
      RECT 8.176 1.026 8.28 5.4 ; 
      RECT 7.744 1.026 7.848 5.4 ; 
      RECT 7.312 1.026 7.416 5.4 ; 
      RECT 6.88 1.026 6.984 5.4 ; 
      RECT 6.448 1.026 6.552 5.4 ; 
      RECT 6.016 1.026 6.12 5.4 ; 
      RECT 5.584 1.026 5.688 5.4 ; 
      RECT 5.152 1.026 5.256 5.4 ; 
      RECT 4.72 1.026 4.824 5.4 ; 
      RECT 4.288 1.026 4.392 5.4 ; 
      RECT 3.856 1.026 3.96 5.4 ; 
      RECT 3.424 1.026 3.528 5.4 ; 
      RECT 2.992 1.026 3.096 5.4 ; 
      RECT 2.56 1.026 2.664 5.4 ; 
      RECT 2.128 1.026 2.232 5.4 ; 
      RECT 1.696 1.026 1.8 5.4 ; 
      RECT 1.264 1.026 1.368 5.4 ; 
      RECT 0.832 1.026 0.936 5.4 ; 
      RECT 0.02 1.026 0.36 5.4 ; 
      RECT 34.564 5.346 35.076 9.72 ; 
      RECT 34.508 8.008 35.076 9.298 ; 
      RECT 33.916 6.916 34.164 9.72 ; 
      RECT 33.86 8.154 34.164 8.768 ; 
      RECT 33.916 5.346 34.02 9.72 ; 
      RECT 33.916 5.83 34.076 6.788 ; 
      RECT 33.916 5.346 34.164 5.702 ; 
      RECT 32.728 7.148 33.552 9.72 ; 
      RECT 33.448 5.346 33.552 9.72 ; 
      RECT 32.728 8.256 33.608 9.288 ; 
      RECT 32.728 5.346 33.12 9.72 ; 
      RECT 31.06 5.346 31.392 9.72 ; 
      RECT 31.06 5.7 31.448 9.442 ; 
      RECT 65.776 5.346 66.116 9.72 ; 
      RECT 65.2 5.346 65.304 9.72 ; 
      RECT 64.768 5.346 64.872 9.72 ; 
      RECT 64.336 5.346 64.44 9.72 ; 
      RECT 63.904 5.346 64.008 9.72 ; 
      RECT 63.472 5.346 63.576 9.72 ; 
      RECT 63.04 5.346 63.144 9.72 ; 
      RECT 62.608 5.346 62.712 9.72 ; 
      RECT 62.176 5.346 62.28 9.72 ; 
      RECT 61.744 5.346 61.848 9.72 ; 
      RECT 61.312 5.346 61.416 9.72 ; 
      RECT 60.88 5.346 60.984 9.72 ; 
      RECT 60.448 5.346 60.552 9.72 ; 
      RECT 60.016 5.346 60.12 9.72 ; 
      RECT 59.584 5.346 59.688 9.72 ; 
      RECT 59.152 5.346 59.256 9.72 ; 
      RECT 58.72 5.346 58.824 9.72 ; 
      RECT 58.288 5.346 58.392 9.72 ; 
      RECT 57.856 5.346 57.96 9.72 ; 
      RECT 57.424 5.346 57.528 9.72 ; 
      RECT 56.992 5.346 57.096 9.72 ; 
      RECT 56.56 5.346 56.664 9.72 ; 
      RECT 56.128 5.346 56.232 9.72 ; 
      RECT 55.696 5.346 55.8 9.72 ; 
      RECT 55.264 5.346 55.368 9.72 ; 
      RECT 54.832 5.346 54.936 9.72 ; 
      RECT 54.4 5.346 54.504 9.72 ; 
      RECT 53.968 5.346 54.072 9.72 ; 
      RECT 53.536 5.346 53.64 9.72 ; 
      RECT 53.104 5.346 53.208 9.72 ; 
      RECT 52.672 5.346 52.776 9.72 ; 
      RECT 52.24 5.346 52.344 9.72 ; 
      RECT 51.808 5.346 51.912 9.72 ; 
      RECT 51.376 5.346 51.48 9.72 ; 
      RECT 50.944 5.346 51.048 9.72 ; 
      RECT 50.512 5.346 50.616 9.72 ; 
      RECT 50.08 5.346 50.184 9.72 ; 
      RECT 49.648 5.346 49.752 9.72 ; 
      RECT 49.216 5.346 49.32 9.72 ; 
      RECT 48.784 5.346 48.888 9.72 ; 
      RECT 48.352 5.346 48.456 9.72 ; 
      RECT 47.92 5.346 48.024 9.72 ; 
      RECT 47.488 5.346 47.592 9.72 ; 
      RECT 47.056 5.346 47.16 9.72 ; 
      RECT 46.624 5.346 46.728 9.72 ; 
      RECT 46.192 5.346 46.296 9.72 ; 
      RECT 45.76 5.346 45.864 9.72 ; 
      RECT 45.328 5.346 45.432 9.72 ; 
      RECT 44.896 5.346 45 9.72 ; 
      RECT 44.464 5.346 44.568 9.72 ; 
      RECT 44.032 5.346 44.136 9.72 ; 
      RECT 43.6 5.346 43.704 9.72 ; 
      RECT 43.168 5.346 43.272 9.72 ; 
      RECT 42.736 5.346 42.84 9.72 ; 
      RECT 42.304 5.346 42.408 9.72 ; 
      RECT 41.872 5.346 41.976 9.72 ; 
      RECT 41.44 5.346 41.544 9.72 ; 
      RECT 41.008 5.346 41.112 9.72 ; 
      RECT 40.576 5.346 40.68 9.72 ; 
      RECT 40.144 5.346 40.248 9.72 ; 
      RECT 39.712 5.346 39.816 9.72 ; 
      RECT 39.28 5.346 39.384 9.72 ; 
      RECT 38.848 5.346 38.952 9.72 ; 
      RECT 38.416 5.346 38.52 9.72 ; 
      RECT 37.984 5.346 38.088 9.72 ; 
      RECT 37.552 5.346 37.656 9.72 ; 
      RECT 36.7 5.346 37.008 9.72 ; 
      RECT 29.128 5.346 29.436 9.72 ; 
      RECT 28.48 5.346 28.584 9.72 ; 
      RECT 28.048 5.346 28.152 9.72 ; 
      RECT 27.616 5.346 27.72 9.72 ; 
      RECT 27.184 5.346 27.288 9.72 ; 
      RECT 26.752 5.346 26.856 9.72 ; 
      RECT 26.32 5.346 26.424 9.72 ; 
      RECT 25.888 5.346 25.992 9.72 ; 
      RECT 25.456 5.346 25.56 9.72 ; 
      RECT 25.024 5.346 25.128 9.72 ; 
      RECT 24.592 5.346 24.696 9.72 ; 
      RECT 24.16 5.346 24.264 9.72 ; 
      RECT 23.728 5.346 23.832 9.72 ; 
      RECT 23.296 5.346 23.4 9.72 ; 
      RECT 22.864 5.346 22.968 9.72 ; 
      RECT 22.432 5.346 22.536 9.72 ; 
      RECT 22 5.346 22.104 9.72 ; 
      RECT 21.568 5.346 21.672 9.72 ; 
      RECT 21.136 5.346 21.24 9.72 ; 
      RECT 20.704 5.346 20.808 9.72 ; 
      RECT 20.272 5.346 20.376 9.72 ; 
      RECT 19.84 5.346 19.944 9.72 ; 
      RECT 19.408 5.346 19.512 9.72 ; 
      RECT 18.976 5.346 19.08 9.72 ; 
      RECT 18.544 5.346 18.648 9.72 ; 
      RECT 18.112 5.346 18.216 9.72 ; 
      RECT 17.68 5.346 17.784 9.72 ; 
      RECT 17.248 5.346 17.352 9.72 ; 
      RECT 16.816 5.346 16.92 9.72 ; 
      RECT 16.384 5.346 16.488 9.72 ; 
      RECT 15.952 5.346 16.056 9.72 ; 
      RECT 15.52 5.346 15.624 9.72 ; 
      RECT 15.088 5.346 15.192 9.72 ; 
      RECT 14.656 5.346 14.76 9.72 ; 
      RECT 14.224 5.346 14.328 9.72 ; 
      RECT 13.792 5.346 13.896 9.72 ; 
      RECT 13.36 5.346 13.464 9.72 ; 
      RECT 12.928 5.346 13.032 9.72 ; 
      RECT 12.496 5.346 12.6 9.72 ; 
      RECT 12.064 5.346 12.168 9.72 ; 
      RECT 11.632 5.346 11.736 9.72 ; 
      RECT 11.2 5.346 11.304 9.72 ; 
      RECT 10.768 5.346 10.872 9.72 ; 
      RECT 10.336 5.346 10.44 9.72 ; 
      RECT 9.904 5.346 10.008 9.72 ; 
      RECT 9.472 5.346 9.576 9.72 ; 
      RECT 9.04 5.346 9.144 9.72 ; 
      RECT 8.608 5.346 8.712 9.72 ; 
      RECT 8.176 5.346 8.28 9.72 ; 
      RECT 7.744 5.346 7.848 9.72 ; 
      RECT 7.312 5.346 7.416 9.72 ; 
      RECT 6.88 5.346 6.984 9.72 ; 
      RECT 6.448 5.346 6.552 9.72 ; 
      RECT 6.016 5.346 6.12 9.72 ; 
      RECT 5.584 5.346 5.688 9.72 ; 
      RECT 5.152 5.346 5.256 9.72 ; 
      RECT 4.72 5.346 4.824 9.72 ; 
      RECT 4.288 5.346 4.392 9.72 ; 
      RECT 3.856 5.346 3.96 9.72 ; 
      RECT 3.424 5.346 3.528 9.72 ; 
      RECT 2.992 5.346 3.096 9.72 ; 
      RECT 2.56 5.346 2.664 9.72 ; 
      RECT 2.128 5.346 2.232 9.72 ; 
      RECT 1.696 5.346 1.8 9.72 ; 
      RECT 1.264 5.346 1.368 9.72 ; 
      RECT 0.832 5.346 0.936 9.72 ; 
      RECT 0.02 5.346 0.36 9.72 ; 
      RECT 34.564 9.666 35.076 14.04 ; 
      RECT 34.508 12.328 35.076 13.618 ; 
      RECT 33.916 11.236 34.164 14.04 ; 
      RECT 33.86 12.474 34.164 13.088 ; 
      RECT 33.916 9.666 34.02 14.04 ; 
      RECT 33.916 10.15 34.076 11.108 ; 
      RECT 33.916 9.666 34.164 10.022 ; 
      RECT 32.728 11.468 33.552 14.04 ; 
      RECT 33.448 9.666 33.552 14.04 ; 
      RECT 32.728 12.576 33.608 13.608 ; 
      RECT 32.728 9.666 33.12 14.04 ; 
      RECT 31.06 9.666 31.392 14.04 ; 
      RECT 31.06 10.02 31.448 13.762 ; 
      RECT 65.776 9.666 66.116 14.04 ; 
      RECT 65.2 9.666 65.304 14.04 ; 
      RECT 64.768 9.666 64.872 14.04 ; 
      RECT 64.336 9.666 64.44 14.04 ; 
      RECT 63.904 9.666 64.008 14.04 ; 
      RECT 63.472 9.666 63.576 14.04 ; 
      RECT 63.04 9.666 63.144 14.04 ; 
      RECT 62.608 9.666 62.712 14.04 ; 
      RECT 62.176 9.666 62.28 14.04 ; 
      RECT 61.744 9.666 61.848 14.04 ; 
      RECT 61.312 9.666 61.416 14.04 ; 
      RECT 60.88 9.666 60.984 14.04 ; 
      RECT 60.448 9.666 60.552 14.04 ; 
      RECT 60.016 9.666 60.12 14.04 ; 
      RECT 59.584 9.666 59.688 14.04 ; 
      RECT 59.152 9.666 59.256 14.04 ; 
      RECT 58.72 9.666 58.824 14.04 ; 
      RECT 58.288 9.666 58.392 14.04 ; 
      RECT 57.856 9.666 57.96 14.04 ; 
      RECT 57.424 9.666 57.528 14.04 ; 
      RECT 56.992 9.666 57.096 14.04 ; 
      RECT 56.56 9.666 56.664 14.04 ; 
      RECT 56.128 9.666 56.232 14.04 ; 
      RECT 55.696 9.666 55.8 14.04 ; 
      RECT 55.264 9.666 55.368 14.04 ; 
      RECT 54.832 9.666 54.936 14.04 ; 
      RECT 54.4 9.666 54.504 14.04 ; 
      RECT 53.968 9.666 54.072 14.04 ; 
      RECT 53.536 9.666 53.64 14.04 ; 
      RECT 53.104 9.666 53.208 14.04 ; 
      RECT 52.672 9.666 52.776 14.04 ; 
      RECT 52.24 9.666 52.344 14.04 ; 
      RECT 51.808 9.666 51.912 14.04 ; 
      RECT 51.376 9.666 51.48 14.04 ; 
      RECT 50.944 9.666 51.048 14.04 ; 
      RECT 50.512 9.666 50.616 14.04 ; 
      RECT 50.08 9.666 50.184 14.04 ; 
      RECT 49.648 9.666 49.752 14.04 ; 
      RECT 49.216 9.666 49.32 14.04 ; 
      RECT 48.784 9.666 48.888 14.04 ; 
      RECT 48.352 9.666 48.456 14.04 ; 
      RECT 47.92 9.666 48.024 14.04 ; 
      RECT 47.488 9.666 47.592 14.04 ; 
      RECT 47.056 9.666 47.16 14.04 ; 
      RECT 46.624 9.666 46.728 14.04 ; 
      RECT 46.192 9.666 46.296 14.04 ; 
      RECT 45.76 9.666 45.864 14.04 ; 
      RECT 45.328 9.666 45.432 14.04 ; 
      RECT 44.896 9.666 45 14.04 ; 
      RECT 44.464 9.666 44.568 14.04 ; 
      RECT 44.032 9.666 44.136 14.04 ; 
      RECT 43.6 9.666 43.704 14.04 ; 
      RECT 43.168 9.666 43.272 14.04 ; 
      RECT 42.736 9.666 42.84 14.04 ; 
      RECT 42.304 9.666 42.408 14.04 ; 
      RECT 41.872 9.666 41.976 14.04 ; 
      RECT 41.44 9.666 41.544 14.04 ; 
      RECT 41.008 9.666 41.112 14.04 ; 
      RECT 40.576 9.666 40.68 14.04 ; 
      RECT 40.144 9.666 40.248 14.04 ; 
      RECT 39.712 9.666 39.816 14.04 ; 
      RECT 39.28 9.666 39.384 14.04 ; 
      RECT 38.848 9.666 38.952 14.04 ; 
      RECT 38.416 9.666 38.52 14.04 ; 
      RECT 37.984 9.666 38.088 14.04 ; 
      RECT 37.552 9.666 37.656 14.04 ; 
      RECT 36.7 9.666 37.008 14.04 ; 
      RECT 29.128 9.666 29.436 14.04 ; 
      RECT 28.48 9.666 28.584 14.04 ; 
      RECT 28.048 9.666 28.152 14.04 ; 
      RECT 27.616 9.666 27.72 14.04 ; 
      RECT 27.184 9.666 27.288 14.04 ; 
      RECT 26.752 9.666 26.856 14.04 ; 
      RECT 26.32 9.666 26.424 14.04 ; 
      RECT 25.888 9.666 25.992 14.04 ; 
      RECT 25.456 9.666 25.56 14.04 ; 
      RECT 25.024 9.666 25.128 14.04 ; 
      RECT 24.592 9.666 24.696 14.04 ; 
      RECT 24.16 9.666 24.264 14.04 ; 
      RECT 23.728 9.666 23.832 14.04 ; 
      RECT 23.296 9.666 23.4 14.04 ; 
      RECT 22.864 9.666 22.968 14.04 ; 
      RECT 22.432 9.666 22.536 14.04 ; 
      RECT 22 9.666 22.104 14.04 ; 
      RECT 21.568 9.666 21.672 14.04 ; 
      RECT 21.136 9.666 21.24 14.04 ; 
      RECT 20.704 9.666 20.808 14.04 ; 
      RECT 20.272 9.666 20.376 14.04 ; 
      RECT 19.84 9.666 19.944 14.04 ; 
      RECT 19.408 9.666 19.512 14.04 ; 
      RECT 18.976 9.666 19.08 14.04 ; 
      RECT 18.544 9.666 18.648 14.04 ; 
      RECT 18.112 9.666 18.216 14.04 ; 
      RECT 17.68 9.666 17.784 14.04 ; 
      RECT 17.248 9.666 17.352 14.04 ; 
      RECT 16.816 9.666 16.92 14.04 ; 
      RECT 16.384 9.666 16.488 14.04 ; 
      RECT 15.952 9.666 16.056 14.04 ; 
      RECT 15.52 9.666 15.624 14.04 ; 
      RECT 15.088 9.666 15.192 14.04 ; 
      RECT 14.656 9.666 14.76 14.04 ; 
      RECT 14.224 9.666 14.328 14.04 ; 
      RECT 13.792 9.666 13.896 14.04 ; 
      RECT 13.36 9.666 13.464 14.04 ; 
      RECT 12.928 9.666 13.032 14.04 ; 
      RECT 12.496 9.666 12.6 14.04 ; 
      RECT 12.064 9.666 12.168 14.04 ; 
      RECT 11.632 9.666 11.736 14.04 ; 
      RECT 11.2 9.666 11.304 14.04 ; 
      RECT 10.768 9.666 10.872 14.04 ; 
      RECT 10.336 9.666 10.44 14.04 ; 
      RECT 9.904 9.666 10.008 14.04 ; 
      RECT 9.472 9.666 9.576 14.04 ; 
      RECT 9.04 9.666 9.144 14.04 ; 
      RECT 8.608 9.666 8.712 14.04 ; 
      RECT 8.176 9.666 8.28 14.04 ; 
      RECT 7.744 9.666 7.848 14.04 ; 
      RECT 7.312 9.666 7.416 14.04 ; 
      RECT 6.88 9.666 6.984 14.04 ; 
      RECT 6.448 9.666 6.552 14.04 ; 
      RECT 6.016 9.666 6.12 14.04 ; 
      RECT 5.584 9.666 5.688 14.04 ; 
      RECT 5.152 9.666 5.256 14.04 ; 
      RECT 4.72 9.666 4.824 14.04 ; 
      RECT 4.288 9.666 4.392 14.04 ; 
      RECT 3.856 9.666 3.96 14.04 ; 
      RECT 3.424 9.666 3.528 14.04 ; 
      RECT 2.992 9.666 3.096 14.04 ; 
      RECT 2.56 9.666 2.664 14.04 ; 
      RECT 2.128 9.666 2.232 14.04 ; 
      RECT 1.696 9.666 1.8 14.04 ; 
      RECT 1.264 9.666 1.368 14.04 ; 
      RECT 0.832 9.666 0.936 14.04 ; 
      RECT 0.02 9.666 0.36 14.04 ; 
      RECT 34.564 13.986 35.076 18.36 ; 
      RECT 34.508 16.648 35.076 17.938 ; 
      RECT 33.916 15.556 34.164 18.36 ; 
      RECT 33.86 16.794 34.164 17.408 ; 
      RECT 33.916 13.986 34.02 18.36 ; 
      RECT 33.916 14.47 34.076 15.428 ; 
      RECT 33.916 13.986 34.164 14.342 ; 
      RECT 32.728 15.788 33.552 18.36 ; 
      RECT 33.448 13.986 33.552 18.36 ; 
      RECT 32.728 16.896 33.608 17.928 ; 
      RECT 32.728 13.986 33.12 18.36 ; 
      RECT 31.06 13.986 31.392 18.36 ; 
      RECT 31.06 14.34 31.448 18.082 ; 
      RECT 65.776 13.986 66.116 18.36 ; 
      RECT 65.2 13.986 65.304 18.36 ; 
      RECT 64.768 13.986 64.872 18.36 ; 
      RECT 64.336 13.986 64.44 18.36 ; 
      RECT 63.904 13.986 64.008 18.36 ; 
      RECT 63.472 13.986 63.576 18.36 ; 
      RECT 63.04 13.986 63.144 18.36 ; 
      RECT 62.608 13.986 62.712 18.36 ; 
      RECT 62.176 13.986 62.28 18.36 ; 
      RECT 61.744 13.986 61.848 18.36 ; 
      RECT 61.312 13.986 61.416 18.36 ; 
      RECT 60.88 13.986 60.984 18.36 ; 
      RECT 60.448 13.986 60.552 18.36 ; 
      RECT 60.016 13.986 60.12 18.36 ; 
      RECT 59.584 13.986 59.688 18.36 ; 
      RECT 59.152 13.986 59.256 18.36 ; 
      RECT 58.72 13.986 58.824 18.36 ; 
      RECT 58.288 13.986 58.392 18.36 ; 
      RECT 57.856 13.986 57.96 18.36 ; 
      RECT 57.424 13.986 57.528 18.36 ; 
      RECT 56.992 13.986 57.096 18.36 ; 
      RECT 56.56 13.986 56.664 18.36 ; 
      RECT 56.128 13.986 56.232 18.36 ; 
      RECT 55.696 13.986 55.8 18.36 ; 
      RECT 55.264 13.986 55.368 18.36 ; 
      RECT 54.832 13.986 54.936 18.36 ; 
      RECT 54.4 13.986 54.504 18.36 ; 
      RECT 53.968 13.986 54.072 18.36 ; 
      RECT 53.536 13.986 53.64 18.36 ; 
      RECT 53.104 13.986 53.208 18.36 ; 
      RECT 52.672 13.986 52.776 18.36 ; 
      RECT 52.24 13.986 52.344 18.36 ; 
      RECT 51.808 13.986 51.912 18.36 ; 
      RECT 51.376 13.986 51.48 18.36 ; 
      RECT 50.944 13.986 51.048 18.36 ; 
      RECT 50.512 13.986 50.616 18.36 ; 
      RECT 50.08 13.986 50.184 18.36 ; 
      RECT 49.648 13.986 49.752 18.36 ; 
      RECT 49.216 13.986 49.32 18.36 ; 
      RECT 48.784 13.986 48.888 18.36 ; 
      RECT 48.352 13.986 48.456 18.36 ; 
      RECT 47.92 13.986 48.024 18.36 ; 
      RECT 47.488 13.986 47.592 18.36 ; 
      RECT 47.056 13.986 47.16 18.36 ; 
      RECT 46.624 13.986 46.728 18.36 ; 
      RECT 46.192 13.986 46.296 18.36 ; 
      RECT 45.76 13.986 45.864 18.36 ; 
      RECT 45.328 13.986 45.432 18.36 ; 
      RECT 44.896 13.986 45 18.36 ; 
      RECT 44.464 13.986 44.568 18.36 ; 
      RECT 44.032 13.986 44.136 18.36 ; 
      RECT 43.6 13.986 43.704 18.36 ; 
      RECT 43.168 13.986 43.272 18.36 ; 
      RECT 42.736 13.986 42.84 18.36 ; 
      RECT 42.304 13.986 42.408 18.36 ; 
      RECT 41.872 13.986 41.976 18.36 ; 
      RECT 41.44 13.986 41.544 18.36 ; 
      RECT 41.008 13.986 41.112 18.36 ; 
      RECT 40.576 13.986 40.68 18.36 ; 
      RECT 40.144 13.986 40.248 18.36 ; 
      RECT 39.712 13.986 39.816 18.36 ; 
      RECT 39.28 13.986 39.384 18.36 ; 
      RECT 38.848 13.986 38.952 18.36 ; 
      RECT 38.416 13.986 38.52 18.36 ; 
      RECT 37.984 13.986 38.088 18.36 ; 
      RECT 37.552 13.986 37.656 18.36 ; 
      RECT 36.7 13.986 37.008 18.36 ; 
      RECT 29.128 13.986 29.436 18.36 ; 
      RECT 28.48 13.986 28.584 18.36 ; 
      RECT 28.048 13.986 28.152 18.36 ; 
      RECT 27.616 13.986 27.72 18.36 ; 
      RECT 27.184 13.986 27.288 18.36 ; 
      RECT 26.752 13.986 26.856 18.36 ; 
      RECT 26.32 13.986 26.424 18.36 ; 
      RECT 25.888 13.986 25.992 18.36 ; 
      RECT 25.456 13.986 25.56 18.36 ; 
      RECT 25.024 13.986 25.128 18.36 ; 
      RECT 24.592 13.986 24.696 18.36 ; 
      RECT 24.16 13.986 24.264 18.36 ; 
      RECT 23.728 13.986 23.832 18.36 ; 
      RECT 23.296 13.986 23.4 18.36 ; 
      RECT 22.864 13.986 22.968 18.36 ; 
      RECT 22.432 13.986 22.536 18.36 ; 
      RECT 22 13.986 22.104 18.36 ; 
      RECT 21.568 13.986 21.672 18.36 ; 
      RECT 21.136 13.986 21.24 18.36 ; 
      RECT 20.704 13.986 20.808 18.36 ; 
      RECT 20.272 13.986 20.376 18.36 ; 
      RECT 19.84 13.986 19.944 18.36 ; 
      RECT 19.408 13.986 19.512 18.36 ; 
      RECT 18.976 13.986 19.08 18.36 ; 
      RECT 18.544 13.986 18.648 18.36 ; 
      RECT 18.112 13.986 18.216 18.36 ; 
      RECT 17.68 13.986 17.784 18.36 ; 
      RECT 17.248 13.986 17.352 18.36 ; 
      RECT 16.816 13.986 16.92 18.36 ; 
      RECT 16.384 13.986 16.488 18.36 ; 
      RECT 15.952 13.986 16.056 18.36 ; 
      RECT 15.52 13.986 15.624 18.36 ; 
      RECT 15.088 13.986 15.192 18.36 ; 
      RECT 14.656 13.986 14.76 18.36 ; 
      RECT 14.224 13.986 14.328 18.36 ; 
      RECT 13.792 13.986 13.896 18.36 ; 
      RECT 13.36 13.986 13.464 18.36 ; 
      RECT 12.928 13.986 13.032 18.36 ; 
      RECT 12.496 13.986 12.6 18.36 ; 
      RECT 12.064 13.986 12.168 18.36 ; 
      RECT 11.632 13.986 11.736 18.36 ; 
      RECT 11.2 13.986 11.304 18.36 ; 
      RECT 10.768 13.986 10.872 18.36 ; 
      RECT 10.336 13.986 10.44 18.36 ; 
      RECT 9.904 13.986 10.008 18.36 ; 
      RECT 9.472 13.986 9.576 18.36 ; 
      RECT 9.04 13.986 9.144 18.36 ; 
      RECT 8.608 13.986 8.712 18.36 ; 
      RECT 8.176 13.986 8.28 18.36 ; 
      RECT 7.744 13.986 7.848 18.36 ; 
      RECT 7.312 13.986 7.416 18.36 ; 
      RECT 6.88 13.986 6.984 18.36 ; 
      RECT 6.448 13.986 6.552 18.36 ; 
      RECT 6.016 13.986 6.12 18.36 ; 
      RECT 5.584 13.986 5.688 18.36 ; 
      RECT 5.152 13.986 5.256 18.36 ; 
      RECT 4.72 13.986 4.824 18.36 ; 
      RECT 4.288 13.986 4.392 18.36 ; 
      RECT 3.856 13.986 3.96 18.36 ; 
      RECT 3.424 13.986 3.528 18.36 ; 
      RECT 2.992 13.986 3.096 18.36 ; 
      RECT 2.56 13.986 2.664 18.36 ; 
      RECT 2.128 13.986 2.232 18.36 ; 
      RECT 1.696 13.986 1.8 18.36 ; 
      RECT 1.264 13.986 1.368 18.36 ; 
      RECT 0.832 13.986 0.936 18.36 ; 
      RECT 0.02 13.986 0.36 18.36 ; 
      RECT 34.564 18.306 35.076 22.68 ; 
      RECT 34.508 20.968 35.076 22.258 ; 
      RECT 33.916 19.876 34.164 22.68 ; 
      RECT 33.86 21.114 34.164 21.728 ; 
      RECT 33.916 18.306 34.02 22.68 ; 
      RECT 33.916 18.79 34.076 19.748 ; 
      RECT 33.916 18.306 34.164 18.662 ; 
      RECT 32.728 20.108 33.552 22.68 ; 
      RECT 33.448 18.306 33.552 22.68 ; 
      RECT 32.728 21.216 33.608 22.248 ; 
      RECT 32.728 18.306 33.12 22.68 ; 
      RECT 31.06 18.306 31.392 22.68 ; 
      RECT 31.06 18.66 31.448 22.402 ; 
      RECT 65.776 18.306 66.116 22.68 ; 
      RECT 65.2 18.306 65.304 22.68 ; 
      RECT 64.768 18.306 64.872 22.68 ; 
      RECT 64.336 18.306 64.44 22.68 ; 
      RECT 63.904 18.306 64.008 22.68 ; 
      RECT 63.472 18.306 63.576 22.68 ; 
      RECT 63.04 18.306 63.144 22.68 ; 
      RECT 62.608 18.306 62.712 22.68 ; 
      RECT 62.176 18.306 62.28 22.68 ; 
      RECT 61.744 18.306 61.848 22.68 ; 
      RECT 61.312 18.306 61.416 22.68 ; 
      RECT 60.88 18.306 60.984 22.68 ; 
      RECT 60.448 18.306 60.552 22.68 ; 
      RECT 60.016 18.306 60.12 22.68 ; 
      RECT 59.584 18.306 59.688 22.68 ; 
      RECT 59.152 18.306 59.256 22.68 ; 
      RECT 58.72 18.306 58.824 22.68 ; 
      RECT 58.288 18.306 58.392 22.68 ; 
      RECT 57.856 18.306 57.96 22.68 ; 
      RECT 57.424 18.306 57.528 22.68 ; 
      RECT 56.992 18.306 57.096 22.68 ; 
      RECT 56.56 18.306 56.664 22.68 ; 
      RECT 56.128 18.306 56.232 22.68 ; 
      RECT 55.696 18.306 55.8 22.68 ; 
      RECT 55.264 18.306 55.368 22.68 ; 
      RECT 54.832 18.306 54.936 22.68 ; 
      RECT 54.4 18.306 54.504 22.68 ; 
      RECT 53.968 18.306 54.072 22.68 ; 
      RECT 53.536 18.306 53.64 22.68 ; 
      RECT 53.104 18.306 53.208 22.68 ; 
      RECT 52.672 18.306 52.776 22.68 ; 
      RECT 52.24 18.306 52.344 22.68 ; 
      RECT 51.808 18.306 51.912 22.68 ; 
      RECT 51.376 18.306 51.48 22.68 ; 
      RECT 50.944 18.306 51.048 22.68 ; 
      RECT 50.512 18.306 50.616 22.68 ; 
      RECT 50.08 18.306 50.184 22.68 ; 
      RECT 49.648 18.306 49.752 22.68 ; 
      RECT 49.216 18.306 49.32 22.68 ; 
      RECT 48.784 18.306 48.888 22.68 ; 
      RECT 48.352 18.306 48.456 22.68 ; 
      RECT 47.92 18.306 48.024 22.68 ; 
      RECT 47.488 18.306 47.592 22.68 ; 
      RECT 47.056 18.306 47.16 22.68 ; 
      RECT 46.624 18.306 46.728 22.68 ; 
      RECT 46.192 18.306 46.296 22.68 ; 
      RECT 45.76 18.306 45.864 22.68 ; 
      RECT 45.328 18.306 45.432 22.68 ; 
      RECT 44.896 18.306 45 22.68 ; 
      RECT 44.464 18.306 44.568 22.68 ; 
      RECT 44.032 18.306 44.136 22.68 ; 
      RECT 43.6 18.306 43.704 22.68 ; 
      RECT 43.168 18.306 43.272 22.68 ; 
      RECT 42.736 18.306 42.84 22.68 ; 
      RECT 42.304 18.306 42.408 22.68 ; 
      RECT 41.872 18.306 41.976 22.68 ; 
      RECT 41.44 18.306 41.544 22.68 ; 
      RECT 41.008 18.306 41.112 22.68 ; 
      RECT 40.576 18.306 40.68 22.68 ; 
      RECT 40.144 18.306 40.248 22.68 ; 
      RECT 39.712 18.306 39.816 22.68 ; 
      RECT 39.28 18.306 39.384 22.68 ; 
      RECT 38.848 18.306 38.952 22.68 ; 
      RECT 38.416 18.306 38.52 22.68 ; 
      RECT 37.984 18.306 38.088 22.68 ; 
      RECT 37.552 18.306 37.656 22.68 ; 
      RECT 36.7 18.306 37.008 22.68 ; 
      RECT 29.128 18.306 29.436 22.68 ; 
      RECT 28.48 18.306 28.584 22.68 ; 
      RECT 28.048 18.306 28.152 22.68 ; 
      RECT 27.616 18.306 27.72 22.68 ; 
      RECT 27.184 18.306 27.288 22.68 ; 
      RECT 26.752 18.306 26.856 22.68 ; 
      RECT 26.32 18.306 26.424 22.68 ; 
      RECT 25.888 18.306 25.992 22.68 ; 
      RECT 25.456 18.306 25.56 22.68 ; 
      RECT 25.024 18.306 25.128 22.68 ; 
      RECT 24.592 18.306 24.696 22.68 ; 
      RECT 24.16 18.306 24.264 22.68 ; 
      RECT 23.728 18.306 23.832 22.68 ; 
      RECT 23.296 18.306 23.4 22.68 ; 
      RECT 22.864 18.306 22.968 22.68 ; 
      RECT 22.432 18.306 22.536 22.68 ; 
      RECT 22 18.306 22.104 22.68 ; 
      RECT 21.568 18.306 21.672 22.68 ; 
      RECT 21.136 18.306 21.24 22.68 ; 
      RECT 20.704 18.306 20.808 22.68 ; 
      RECT 20.272 18.306 20.376 22.68 ; 
      RECT 19.84 18.306 19.944 22.68 ; 
      RECT 19.408 18.306 19.512 22.68 ; 
      RECT 18.976 18.306 19.08 22.68 ; 
      RECT 18.544 18.306 18.648 22.68 ; 
      RECT 18.112 18.306 18.216 22.68 ; 
      RECT 17.68 18.306 17.784 22.68 ; 
      RECT 17.248 18.306 17.352 22.68 ; 
      RECT 16.816 18.306 16.92 22.68 ; 
      RECT 16.384 18.306 16.488 22.68 ; 
      RECT 15.952 18.306 16.056 22.68 ; 
      RECT 15.52 18.306 15.624 22.68 ; 
      RECT 15.088 18.306 15.192 22.68 ; 
      RECT 14.656 18.306 14.76 22.68 ; 
      RECT 14.224 18.306 14.328 22.68 ; 
      RECT 13.792 18.306 13.896 22.68 ; 
      RECT 13.36 18.306 13.464 22.68 ; 
      RECT 12.928 18.306 13.032 22.68 ; 
      RECT 12.496 18.306 12.6 22.68 ; 
      RECT 12.064 18.306 12.168 22.68 ; 
      RECT 11.632 18.306 11.736 22.68 ; 
      RECT 11.2 18.306 11.304 22.68 ; 
      RECT 10.768 18.306 10.872 22.68 ; 
      RECT 10.336 18.306 10.44 22.68 ; 
      RECT 9.904 18.306 10.008 22.68 ; 
      RECT 9.472 18.306 9.576 22.68 ; 
      RECT 9.04 18.306 9.144 22.68 ; 
      RECT 8.608 18.306 8.712 22.68 ; 
      RECT 8.176 18.306 8.28 22.68 ; 
      RECT 7.744 18.306 7.848 22.68 ; 
      RECT 7.312 18.306 7.416 22.68 ; 
      RECT 6.88 18.306 6.984 22.68 ; 
      RECT 6.448 18.306 6.552 22.68 ; 
      RECT 6.016 18.306 6.12 22.68 ; 
      RECT 5.584 18.306 5.688 22.68 ; 
      RECT 5.152 18.306 5.256 22.68 ; 
      RECT 4.72 18.306 4.824 22.68 ; 
      RECT 4.288 18.306 4.392 22.68 ; 
      RECT 3.856 18.306 3.96 22.68 ; 
      RECT 3.424 18.306 3.528 22.68 ; 
      RECT 2.992 18.306 3.096 22.68 ; 
      RECT 2.56 18.306 2.664 22.68 ; 
      RECT 2.128 18.306 2.232 22.68 ; 
      RECT 1.696 18.306 1.8 22.68 ; 
      RECT 1.264 18.306 1.368 22.68 ; 
      RECT 0.832 18.306 0.936 22.68 ; 
      RECT 0.02 18.306 0.36 22.68 ; 
      RECT 34.564 22.626 35.076 27 ; 
      RECT 34.508 25.288 35.076 26.578 ; 
      RECT 33.916 24.196 34.164 27 ; 
      RECT 33.86 25.434 34.164 26.048 ; 
      RECT 33.916 22.626 34.02 27 ; 
      RECT 33.916 23.11 34.076 24.068 ; 
      RECT 33.916 22.626 34.164 22.982 ; 
      RECT 32.728 24.428 33.552 27 ; 
      RECT 33.448 22.626 33.552 27 ; 
      RECT 32.728 25.536 33.608 26.568 ; 
      RECT 32.728 22.626 33.12 27 ; 
      RECT 31.06 22.626 31.392 27 ; 
      RECT 31.06 22.98 31.448 26.722 ; 
      RECT 65.776 22.626 66.116 27 ; 
      RECT 65.2 22.626 65.304 27 ; 
      RECT 64.768 22.626 64.872 27 ; 
      RECT 64.336 22.626 64.44 27 ; 
      RECT 63.904 22.626 64.008 27 ; 
      RECT 63.472 22.626 63.576 27 ; 
      RECT 63.04 22.626 63.144 27 ; 
      RECT 62.608 22.626 62.712 27 ; 
      RECT 62.176 22.626 62.28 27 ; 
      RECT 61.744 22.626 61.848 27 ; 
      RECT 61.312 22.626 61.416 27 ; 
      RECT 60.88 22.626 60.984 27 ; 
      RECT 60.448 22.626 60.552 27 ; 
      RECT 60.016 22.626 60.12 27 ; 
      RECT 59.584 22.626 59.688 27 ; 
      RECT 59.152 22.626 59.256 27 ; 
      RECT 58.72 22.626 58.824 27 ; 
      RECT 58.288 22.626 58.392 27 ; 
      RECT 57.856 22.626 57.96 27 ; 
      RECT 57.424 22.626 57.528 27 ; 
      RECT 56.992 22.626 57.096 27 ; 
      RECT 56.56 22.626 56.664 27 ; 
      RECT 56.128 22.626 56.232 27 ; 
      RECT 55.696 22.626 55.8 27 ; 
      RECT 55.264 22.626 55.368 27 ; 
      RECT 54.832 22.626 54.936 27 ; 
      RECT 54.4 22.626 54.504 27 ; 
      RECT 53.968 22.626 54.072 27 ; 
      RECT 53.536 22.626 53.64 27 ; 
      RECT 53.104 22.626 53.208 27 ; 
      RECT 52.672 22.626 52.776 27 ; 
      RECT 52.24 22.626 52.344 27 ; 
      RECT 51.808 22.626 51.912 27 ; 
      RECT 51.376 22.626 51.48 27 ; 
      RECT 50.944 22.626 51.048 27 ; 
      RECT 50.512 22.626 50.616 27 ; 
      RECT 50.08 22.626 50.184 27 ; 
      RECT 49.648 22.626 49.752 27 ; 
      RECT 49.216 22.626 49.32 27 ; 
      RECT 48.784 22.626 48.888 27 ; 
      RECT 48.352 22.626 48.456 27 ; 
      RECT 47.92 22.626 48.024 27 ; 
      RECT 47.488 22.626 47.592 27 ; 
      RECT 47.056 22.626 47.16 27 ; 
      RECT 46.624 22.626 46.728 27 ; 
      RECT 46.192 22.626 46.296 27 ; 
      RECT 45.76 22.626 45.864 27 ; 
      RECT 45.328 22.626 45.432 27 ; 
      RECT 44.896 22.626 45 27 ; 
      RECT 44.464 22.626 44.568 27 ; 
      RECT 44.032 22.626 44.136 27 ; 
      RECT 43.6 22.626 43.704 27 ; 
      RECT 43.168 22.626 43.272 27 ; 
      RECT 42.736 22.626 42.84 27 ; 
      RECT 42.304 22.626 42.408 27 ; 
      RECT 41.872 22.626 41.976 27 ; 
      RECT 41.44 22.626 41.544 27 ; 
      RECT 41.008 22.626 41.112 27 ; 
      RECT 40.576 22.626 40.68 27 ; 
      RECT 40.144 22.626 40.248 27 ; 
      RECT 39.712 22.626 39.816 27 ; 
      RECT 39.28 22.626 39.384 27 ; 
      RECT 38.848 22.626 38.952 27 ; 
      RECT 38.416 22.626 38.52 27 ; 
      RECT 37.984 22.626 38.088 27 ; 
      RECT 37.552 22.626 37.656 27 ; 
      RECT 36.7 22.626 37.008 27 ; 
      RECT 29.128 22.626 29.436 27 ; 
      RECT 28.48 22.626 28.584 27 ; 
      RECT 28.048 22.626 28.152 27 ; 
      RECT 27.616 22.626 27.72 27 ; 
      RECT 27.184 22.626 27.288 27 ; 
      RECT 26.752 22.626 26.856 27 ; 
      RECT 26.32 22.626 26.424 27 ; 
      RECT 25.888 22.626 25.992 27 ; 
      RECT 25.456 22.626 25.56 27 ; 
      RECT 25.024 22.626 25.128 27 ; 
      RECT 24.592 22.626 24.696 27 ; 
      RECT 24.16 22.626 24.264 27 ; 
      RECT 23.728 22.626 23.832 27 ; 
      RECT 23.296 22.626 23.4 27 ; 
      RECT 22.864 22.626 22.968 27 ; 
      RECT 22.432 22.626 22.536 27 ; 
      RECT 22 22.626 22.104 27 ; 
      RECT 21.568 22.626 21.672 27 ; 
      RECT 21.136 22.626 21.24 27 ; 
      RECT 20.704 22.626 20.808 27 ; 
      RECT 20.272 22.626 20.376 27 ; 
      RECT 19.84 22.626 19.944 27 ; 
      RECT 19.408 22.626 19.512 27 ; 
      RECT 18.976 22.626 19.08 27 ; 
      RECT 18.544 22.626 18.648 27 ; 
      RECT 18.112 22.626 18.216 27 ; 
      RECT 17.68 22.626 17.784 27 ; 
      RECT 17.248 22.626 17.352 27 ; 
      RECT 16.816 22.626 16.92 27 ; 
      RECT 16.384 22.626 16.488 27 ; 
      RECT 15.952 22.626 16.056 27 ; 
      RECT 15.52 22.626 15.624 27 ; 
      RECT 15.088 22.626 15.192 27 ; 
      RECT 14.656 22.626 14.76 27 ; 
      RECT 14.224 22.626 14.328 27 ; 
      RECT 13.792 22.626 13.896 27 ; 
      RECT 13.36 22.626 13.464 27 ; 
      RECT 12.928 22.626 13.032 27 ; 
      RECT 12.496 22.626 12.6 27 ; 
      RECT 12.064 22.626 12.168 27 ; 
      RECT 11.632 22.626 11.736 27 ; 
      RECT 11.2 22.626 11.304 27 ; 
      RECT 10.768 22.626 10.872 27 ; 
      RECT 10.336 22.626 10.44 27 ; 
      RECT 9.904 22.626 10.008 27 ; 
      RECT 9.472 22.626 9.576 27 ; 
      RECT 9.04 22.626 9.144 27 ; 
      RECT 8.608 22.626 8.712 27 ; 
      RECT 8.176 22.626 8.28 27 ; 
      RECT 7.744 22.626 7.848 27 ; 
      RECT 7.312 22.626 7.416 27 ; 
      RECT 6.88 22.626 6.984 27 ; 
      RECT 6.448 22.626 6.552 27 ; 
      RECT 6.016 22.626 6.12 27 ; 
      RECT 5.584 22.626 5.688 27 ; 
      RECT 5.152 22.626 5.256 27 ; 
      RECT 4.72 22.626 4.824 27 ; 
      RECT 4.288 22.626 4.392 27 ; 
      RECT 3.856 22.626 3.96 27 ; 
      RECT 3.424 22.626 3.528 27 ; 
      RECT 2.992 22.626 3.096 27 ; 
      RECT 2.56 22.626 2.664 27 ; 
      RECT 2.128 22.626 2.232 27 ; 
      RECT 1.696 22.626 1.8 27 ; 
      RECT 1.264 22.626 1.368 27 ; 
      RECT 0.832 22.626 0.936 27 ; 
      RECT 0.02 22.626 0.36 27 ; 
      RECT 34.564 26.946 35.076 31.32 ; 
      RECT 34.508 29.608 35.076 30.898 ; 
      RECT 33.916 28.516 34.164 31.32 ; 
      RECT 33.86 29.754 34.164 30.368 ; 
      RECT 33.916 26.946 34.02 31.32 ; 
      RECT 33.916 27.43 34.076 28.388 ; 
      RECT 33.916 26.946 34.164 27.302 ; 
      RECT 32.728 28.748 33.552 31.32 ; 
      RECT 33.448 26.946 33.552 31.32 ; 
      RECT 32.728 29.856 33.608 30.888 ; 
      RECT 32.728 26.946 33.12 31.32 ; 
      RECT 31.06 26.946 31.392 31.32 ; 
      RECT 31.06 27.3 31.448 31.042 ; 
      RECT 65.776 26.946 66.116 31.32 ; 
      RECT 65.2 26.946 65.304 31.32 ; 
      RECT 64.768 26.946 64.872 31.32 ; 
      RECT 64.336 26.946 64.44 31.32 ; 
      RECT 63.904 26.946 64.008 31.32 ; 
      RECT 63.472 26.946 63.576 31.32 ; 
      RECT 63.04 26.946 63.144 31.32 ; 
      RECT 62.608 26.946 62.712 31.32 ; 
      RECT 62.176 26.946 62.28 31.32 ; 
      RECT 61.744 26.946 61.848 31.32 ; 
      RECT 61.312 26.946 61.416 31.32 ; 
      RECT 60.88 26.946 60.984 31.32 ; 
      RECT 60.448 26.946 60.552 31.32 ; 
      RECT 60.016 26.946 60.12 31.32 ; 
      RECT 59.584 26.946 59.688 31.32 ; 
      RECT 59.152 26.946 59.256 31.32 ; 
      RECT 58.72 26.946 58.824 31.32 ; 
      RECT 58.288 26.946 58.392 31.32 ; 
      RECT 57.856 26.946 57.96 31.32 ; 
      RECT 57.424 26.946 57.528 31.32 ; 
      RECT 56.992 26.946 57.096 31.32 ; 
      RECT 56.56 26.946 56.664 31.32 ; 
      RECT 56.128 26.946 56.232 31.32 ; 
      RECT 55.696 26.946 55.8 31.32 ; 
      RECT 55.264 26.946 55.368 31.32 ; 
      RECT 54.832 26.946 54.936 31.32 ; 
      RECT 54.4 26.946 54.504 31.32 ; 
      RECT 53.968 26.946 54.072 31.32 ; 
      RECT 53.536 26.946 53.64 31.32 ; 
      RECT 53.104 26.946 53.208 31.32 ; 
      RECT 52.672 26.946 52.776 31.32 ; 
      RECT 52.24 26.946 52.344 31.32 ; 
      RECT 51.808 26.946 51.912 31.32 ; 
      RECT 51.376 26.946 51.48 31.32 ; 
      RECT 50.944 26.946 51.048 31.32 ; 
      RECT 50.512 26.946 50.616 31.32 ; 
      RECT 50.08 26.946 50.184 31.32 ; 
      RECT 49.648 26.946 49.752 31.32 ; 
      RECT 49.216 26.946 49.32 31.32 ; 
      RECT 48.784 26.946 48.888 31.32 ; 
      RECT 48.352 26.946 48.456 31.32 ; 
      RECT 47.92 26.946 48.024 31.32 ; 
      RECT 47.488 26.946 47.592 31.32 ; 
      RECT 47.056 26.946 47.16 31.32 ; 
      RECT 46.624 26.946 46.728 31.32 ; 
      RECT 46.192 26.946 46.296 31.32 ; 
      RECT 45.76 26.946 45.864 31.32 ; 
      RECT 45.328 26.946 45.432 31.32 ; 
      RECT 44.896 26.946 45 31.32 ; 
      RECT 44.464 26.946 44.568 31.32 ; 
      RECT 44.032 26.946 44.136 31.32 ; 
      RECT 43.6 26.946 43.704 31.32 ; 
      RECT 43.168 26.946 43.272 31.32 ; 
      RECT 42.736 26.946 42.84 31.32 ; 
      RECT 42.304 26.946 42.408 31.32 ; 
      RECT 41.872 26.946 41.976 31.32 ; 
      RECT 41.44 26.946 41.544 31.32 ; 
      RECT 41.008 26.946 41.112 31.32 ; 
      RECT 40.576 26.946 40.68 31.32 ; 
      RECT 40.144 26.946 40.248 31.32 ; 
      RECT 39.712 26.946 39.816 31.32 ; 
      RECT 39.28 26.946 39.384 31.32 ; 
      RECT 38.848 26.946 38.952 31.32 ; 
      RECT 38.416 26.946 38.52 31.32 ; 
      RECT 37.984 26.946 38.088 31.32 ; 
      RECT 37.552 26.946 37.656 31.32 ; 
      RECT 36.7 26.946 37.008 31.32 ; 
      RECT 29.128 26.946 29.436 31.32 ; 
      RECT 28.48 26.946 28.584 31.32 ; 
      RECT 28.048 26.946 28.152 31.32 ; 
      RECT 27.616 26.946 27.72 31.32 ; 
      RECT 27.184 26.946 27.288 31.32 ; 
      RECT 26.752 26.946 26.856 31.32 ; 
      RECT 26.32 26.946 26.424 31.32 ; 
      RECT 25.888 26.946 25.992 31.32 ; 
      RECT 25.456 26.946 25.56 31.32 ; 
      RECT 25.024 26.946 25.128 31.32 ; 
      RECT 24.592 26.946 24.696 31.32 ; 
      RECT 24.16 26.946 24.264 31.32 ; 
      RECT 23.728 26.946 23.832 31.32 ; 
      RECT 23.296 26.946 23.4 31.32 ; 
      RECT 22.864 26.946 22.968 31.32 ; 
      RECT 22.432 26.946 22.536 31.32 ; 
      RECT 22 26.946 22.104 31.32 ; 
      RECT 21.568 26.946 21.672 31.32 ; 
      RECT 21.136 26.946 21.24 31.32 ; 
      RECT 20.704 26.946 20.808 31.32 ; 
      RECT 20.272 26.946 20.376 31.32 ; 
      RECT 19.84 26.946 19.944 31.32 ; 
      RECT 19.408 26.946 19.512 31.32 ; 
      RECT 18.976 26.946 19.08 31.32 ; 
      RECT 18.544 26.946 18.648 31.32 ; 
      RECT 18.112 26.946 18.216 31.32 ; 
      RECT 17.68 26.946 17.784 31.32 ; 
      RECT 17.248 26.946 17.352 31.32 ; 
      RECT 16.816 26.946 16.92 31.32 ; 
      RECT 16.384 26.946 16.488 31.32 ; 
      RECT 15.952 26.946 16.056 31.32 ; 
      RECT 15.52 26.946 15.624 31.32 ; 
      RECT 15.088 26.946 15.192 31.32 ; 
      RECT 14.656 26.946 14.76 31.32 ; 
      RECT 14.224 26.946 14.328 31.32 ; 
      RECT 13.792 26.946 13.896 31.32 ; 
      RECT 13.36 26.946 13.464 31.32 ; 
      RECT 12.928 26.946 13.032 31.32 ; 
      RECT 12.496 26.946 12.6 31.32 ; 
      RECT 12.064 26.946 12.168 31.32 ; 
      RECT 11.632 26.946 11.736 31.32 ; 
      RECT 11.2 26.946 11.304 31.32 ; 
      RECT 10.768 26.946 10.872 31.32 ; 
      RECT 10.336 26.946 10.44 31.32 ; 
      RECT 9.904 26.946 10.008 31.32 ; 
      RECT 9.472 26.946 9.576 31.32 ; 
      RECT 9.04 26.946 9.144 31.32 ; 
      RECT 8.608 26.946 8.712 31.32 ; 
      RECT 8.176 26.946 8.28 31.32 ; 
      RECT 7.744 26.946 7.848 31.32 ; 
      RECT 7.312 26.946 7.416 31.32 ; 
      RECT 6.88 26.946 6.984 31.32 ; 
      RECT 6.448 26.946 6.552 31.32 ; 
      RECT 6.016 26.946 6.12 31.32 ; 
      RECT 5.584 26.946 5.688 31.32 ; 
      RECT 5.152 26.946 5.256 31.32 ; 
      RECT 4.72 26.946 4.824 31.32 ; 
      RECT 4.288 26.946 4.392 31.32 ; 
      RECT 3.856 26.946 3.96 31.32 ; 
      RECT 3.424 26.946 3.528 31.32 ; 
      RECT 2.992 26.946 3.096 31.32 ; 
      RECT 2.56 26.946 2.664 31.32 ; 
      RECT 2.128 26.946 2.232 31.32 ; 
      RECT 1.696 26.946 1.8 31.32 ; 
      RECT 1.264 26.946 1.368 31.32 ; 
      RECT 0.832 26.946 0.936 31.32 ; 
      RECT 0.02 26.946 0.36 31.32 ; 
      RECT 34.564 31.266 35.076 35.64 ; 
      RECT 34.508 33.928 35.076 35.218 ; 
      RECT 33.916 32.836 34.164 35.64 ; 
      RECT 33.86 34.074 34.164 34.688 ; 
      RECT 33.916 31.266 34.02 35.64 ; 
      RECT 33.916 31.75 34.076 32.708 ; 
      RECT 33.916 31.266 34.164 31.622 ; 
      RECT 32.728 33.068 33.552 35.64 ; 
      RECT 33.448 31.266 33.552 35.64 ; 
      RECT 32.728 34.176 33.608 35.208 ; 
      RECT 32.728 31.266 33.12 35.64 ; 
      RECT 31.06 31.266 31.392 35.64 ; 
      RECT 31.06 31.62 31.448 35.362 ; 
      RECT 65.776 31.266 66.116 35.64 ; 
      RECT 65.2 31.266 65.304 35.64 ; 
      RECT 64.768 31.266 64.872 35.64 ; 
      RECT 64.336 31.266 64.44 35.64 ; 
      RECT 63.904 31.266 64.008 35.64 ; 
      RECT 63.472 31.266 63.576 35.64 ; 
      RECT 63.04 31.266 63.144 35.64 ; 
      RECT 62.608 31.266 62.712 35.64 ; 
      RECT 62.176 31.266 62.28 35.64 ; 
      RECT 61.744 31.266 61.848 35.64 ; 
      RECT 61.312 31.266 61.416 35.64 ; 
      RECT 60.88 31.266 60.984 35.64 ; 
      RECT 60.448 31.266 60.552 35.64 ; 
      RECT 60.016 31.266 60.12 35.64 ; 
      RECT 59.584 31.266 59.688 35.64 ; 
      RECT 59.152 31.266 59.256 35.64 ; 
      RECT 58.72 31.266 58.824 35.64 ; 
      RECT 58.288 31.266 58.392 35.64 ; 
      RECT 57.856 31.266 57.96 35.64 ; 
      RECT 57.424 31.266 57.528 35.64 ; 
      RECT 56.992 31.266 57.096 35.64 ; 
      RECT 56.56 31.266 56.664 35.64 ; 
      RECT 56.128 31.266 56.232 35.64 ; 
      RECT 55.696 31.266 55.8 35.64 ; 
      RECT 55.264 31.266 55.368 35.64 ; 
      RECT 54.832 31.266 54.936 35.64 ; 
      RECT 54.4 31.266 54.504 35.64 ; 
      RECT 53.968 31.266 54.072 35.64 ; 
      RECT 53.536 31.266 53.64 35.64 ; 
      RECT 53.104 31.266 53.208 35.64 ; 
      RECT 52.672 31.266 52.776 35.64 ; 
      RECT 52.24 31.266 52.344 35.64 ; 
      RECT 51.808 31.266 51.912 35.64 ; 
      RECT 51.376 31.266 51.48 35.64 ; 
      RECT 50.944 31.266 51.048 35.64 ; 
      RECT 50.512 31.266 50.616 35.64 ; 
      RECT 50.08 31.266 50.184 35.64 ; 
      RECT 49.648 31.266 49.752 35.64 ; 
      RECT 49.216 31.266 49.32 35.64 ; 
      RECT 48.784 31.266 48.888 35.64 ; 
      RECT 48.352 31.266 48.456 35.64 ; 
      RECT 47.92 31.266 48.024 35.64 ; 
      RECT 47.488 31.266 47.592 35.64 ; 
      RECT 47.056 31.266 47.16 35.64 ; 
      RECT 46.624 31.266 46.728 35.64 ; 
      RECT 46.192 31.266 46.296 35.64 ; 
      RECT 45.76 31.266 45.864 35.64 ; 
      RECT 45.328 31.266 45.432 35.64 ; 
      RECT 44.896 31.266 45 35.64 ; 
      RECT 44.464 31.266 44.568 35.64 ; 
      RECT 44.032 31.266 44.136 35.64 ; 
      RECT 43.6 31.266 43.704 35.64 ; 
      RECT 43.168 31.266 43.272 35.64 ; 
      RECT 42.736 31.266 42.84 35.64 ; 
      RECT 42.304 31.266 42.408 35.64 ; 
      RECT 41.872 31.266 41.976 35.64 ; 
      RECT 41.44 31.266 41.544 35.64 ; 
      RECT 41.008 31.266 41.112 35.64 ; 
      RECT 40.576 31.266 40.68 35.64 ; 
      RECT 40.144 31.266 40.248 35.64 ; 
      RECT 39.712 31.266 39.816 35.64 ; 
      RECT 39.28 31.266 39.384 35.64 ; 
      RECT 38.848 31.266 38.952 35.64 ; 
      RECT 38.416 31.266 38.52 35.64 ; 
      RECT 37.984 31.266 38.088 35.64 ; 
      RECT 37.552 31.266 37.656 35.64 ; 
      RECT 36.7 31.266 37.008 35.64 ; 
      RECT 29.128 31.266 29.436 35.64 ; 
      RECT 28.48 31.266 28.584 35.64 ; 
      RECT 28.048 31.266 28.152 35.64 ; 
      RECT 27.616 31.266 27.72 35.64 ; 
      RECT 27.184 31.266 27.288 35.64 ; 
      RECT 26.752 31.266 26.856 35.64 ; 
      RECT 26.32 31.266 26.424 35.64 ; 
      RECT 25.888 31.266 25.992 35.64 ; 
      RECT 25.456 31.266 25.56 35.64 ; 
      RECT 25.024 31.266 25.128 35.64 ; 
      RECT 24.592 31.266 24.696 35.64 ; 
      RECT 24.16 31.266 24.264 35.64 ; 
      RECT 23.728 31.266 23.832 35.64 ; 
      RECT 23.296 31.266 23.4 35.64 ; 
      RECT 22.864 31.266 22.968 35.64 ; 
      RECT 22.432 31.266 22.536 35.64 ; 
      RECT 22 31.266 22.104 35.64 ; 
      RECT 21.568 31.266 21.672 35.64 ; 
      RECT 21.136 31.266 21.24 35.64 ; 
      RECT 20.704 31.266 20.808 35.64 ; 
      RECT 20.272 31.266 20.376 35.64 ; 
      RECT 19.84 31.266 19.944 35.64 ; 
      RECT 19.408 31.266 19.512 35.64 ; 
      RECT 18.976 31.266 19.08 35.64 ; 
      RECT 18.544 31.266 18.648 35.64 ; 
      RECT 18.112 31.266 18.216 35.64 ; 
      RECT 17.68 31.266 17.784 35.64 ; 
      RECT 17.248 31.266 17.352 35.64 ; 
      RECT 16.816 31.266 16.92 35.64 ; 
      RECT 16.384 31.266 16.488 35.64 ; 
      RECT 15.952 31.266 16.056 35.64 ; 
      RECT 15.52 31.266 15.624 35.64 ; 
      RECT 15.088 31.266 15.192 35.64 ; 
      RECT 14.656 31.266 14.76 35.64 ; 
      RECT 14.224 31.266 14.328 35.64 ; 
      RECT 13.792 31.266 13.896 35.64 ; 
      RECT 13.36 31.266 13.464 35.64 ; 
      RECT 12.928 31.266 13.032 35.64 ; 
      RECT 12.496 31.266 12.6 35.64 ; 
      RECT 12.064 31.266 12.168 35.64 ; 
      RECT 11.632 31.266 11.736 35.64 ; 
      RECT 11.2 31.266 11.304 35.64 ; 
      RECT 10.768 31.266 10.872 35.64 ; 
      RECT 10.336 31.266 10.44 35.64 ; 
      RECT 9.904 31.266 10.008 35.64 ; 
      RECT 9.472 31.266 9.576 35.64 ; 
      RECT 9.04 31.266 9.144 35.64 ; 
      RECT 8.608 31.266 8.712 35.64 ; 
      RECT 8.176 31.266 8.28 35.64 ; 
      RECT 7.744 31.266 7.848 35.64 ; 
      RECT 7.312 31.266 7.416 35.64 ; 
      RECT 6.88 31.266 6.984 35.64 ; 
      RECT 6.448 31.266 6.552 35.64 ; 
      RECT 6.016 31.266 6.12 35.64 ; 
      RECT 5.584 31.266 5.688 35.64 ; 
      RECT 5.152 31.266 5.256 35.64 ; 
      RECT 4.72 31.266 4.824 35.64 ; 
      RECT 4.288 31.266 4.392 35.64 ; 
      RECT 3.856 31.266 3.96 35.64 ; 
      RECT 3.424 31.266 3.528 35.64 ; 
      RECT 2.992 31.266 3.096 35.64 ; 
      RECT 2.56 31.266 2.664 35.64 ; 
      RECT 2.128 31.266 2.232 35.64 ; 
      RECT 1.696 31.266 1.8 35.64 ; 
      RECT 1.264 31.266 1.368 35.64 ; 
      RECT 0.832 31.266 0.936 35.64 ; 
      RECT 0.02 31.266 0.36 35.64 ; 
      RECT 34.564 35.586 35.076 39.96 ; 
      RECT 34.508 38.248 35.076 39.538 ; 
      RECT 33.916 37.156 34.164 39.96 ; 
      RECT 33.86 38.394 34.164 39.008 ; 
      RECT 33.916 35.586 34.02 39.96 ; 
      RECT 33.916 36.07 34.076 37.028 ; 
      RECT 33.916 35.586 34.164 35.942 ; 
      RECT 32.728 37.388 33.552 39.96 ; 
      RECT 33.448 35.586 33.552 39.96 ; 
      RECT 32.728 38.496 33.608 39.528 ; 
      RECT 32.728 35.586 33.12 39.96 ; 
      RECT 31.06 35.586 31.392 39.96 ; 
      RECT 31.06 35.94 31.448 39.682 ; 
      RECT 65.776 35.586 66.116 39.96 ; 
      RECT 65.2 35.586 65.304 39.96 ; 
      RECT 64.768 35.586 64.872 39.96 ; 
      RECT 64.336 35.586 64.44 39.96 ; 
      RECT 63.904 35.586 64.008 39.96 ; 
      RECT 63.472 35.586 63.576 39.96 ; 
      RECT 63.04 35.586 63.144 39.96 ; 
      RECT 62.608 35.586 62.712 39.96 ; 
      RECT 62.176 35.586 62.28 39.96 ; 
      RECT 61.744 35.586 61.848 39.96 ; 
      RECT 61.312 35.586 61.416 39.96 ; 
      RECT 60.88 35.586 60.984 39.96 ; 
      RECT 60.448 35.586 60.552 39.96 ; 
      RECT 60.016 35.586 60.12 39.96 ; 
      RECT 59.584 35.586 59.688 39.96 ; 
      RECT 59.152 35.586 59.256 39.96 ; 
      RECT 58.72 35.586 58.824 39.96 ; 
      RECT 58.288 35.586 58.392 39.96 ; 
      RECT 57.856 35.586 57.96 39.96 ; 
      RECT 57.424 35.586 57.528 39.96 ; 
      RECT 56.992 35.586 57.096 39.96 ; 
      RECT 56.56 35.586 56.664 39.96 ; 
      RECT 56.128 35.586 56.232 39.96 ; 
      RECT 55.696 35.586 55.8 39.96 ; 
      RECT 55.264 35.586 55.368 39.96 ; 
      RECT 54.832 35.586 54.936 39.96 ; 
      RECT 54.4 35.586 54.504 39.96 ; 
      RECT 53.968 35.586 54.072 39.96 ; 
      RECT 53.536 35.586 53.64 39.96 ; 
      RECT 53.104 35.586 53.208 39.96 ; 
      RECT 52.672 35.586 52.776 39.96 ; 
      RECT 52.24 35.586 52.344 39.96 ; 
      RECT 51.808 35.586 51.912 39.96 ; 
      RECT 51.376 35.586 51.48 39.96 ; 
      RECT 50.944 35.586 51.048 39.96 ; 
      RECT 50.512 35.586 50.616 39.96 ; 
      RECT 50.08 35.586 50.184 39.96 ; 
      RECT 49.648 35.586 49.752 39.96 ; 
      RECT 49.216 35.586 49.32 39.96 ; 
      RECT 48.784 35.586 48.888 39.96 ; 
      RECT 48.352 35.586 48.456 39.96 ; 
      RECT 47.92 35.586 48.024 39.96 ; 
      RECT 47.488 35.586 47.592 39.96 ; 
      RECT 47.056 35.586 47.16 39.96 ; 
      RECT 46.624 35.586 46.728 39.96 ; 
      RECT 46.192 35.586 46.296 39.96 ; 
      RECT 45.76 35.586 45.864 39.96 ; 
      RECT 45.328 35.586 45.432 39.96 ; 
      RECT 44.896 35.586 45 39.96 ; 
      RECT 44.464 35.586 44.568 39.96 ; 
      RECT 44.032 35.586 44.136 39.96 ; 
      RECT 43.6 35.586 43.704 39.96 ; 
      RECT 43.168 35.586 43.272 39.96 ; 
      RECT 42.736 35.586 42.84 39.96 ; 
      RECT 42.304 35.586 42.408 39.96 ; 
      RECT 41.872 35.586 41.976 39.96 ; 
      RECT 41.44 35.586 41.544 39.96 ; 
      RECT 41.008 35.586 41.112 39.96 ; 
      RECT 40.576 35.586 40.68 39.96 ; 
      RECT 40.144 35.586 40.248 39.96 ; 
      RECT 39.712 35.586 39.816 39.96 ; 
      RECT 39.28 35.586 39.384 39.96 ; 
      RECT 38.848 35.586 38.952 39.96 ; 
      RECT 38.416 35.586 38.52 39.96 ; 
      RECT 37.984 35.586 38.088 39.96 ; 
      RECT 37.552 35.586 37.656 39.96 ; 
      RECT 36.7 35.586 37.008 39.96 ; 
      RECT 29.128 35.586 29.436 39.96 ; 
      RECT 28.48 35.586 28.584 39.96 ; 
      RECT 28.048 35.586 28.152 39.96 ; 
      RECT 27.616 35.586 27.72 39.96 ; 
      RECT 27.184 35.586 27.288 39.96 ; 
      RECT 26.752 35.586 26.856 39.96 ; 
      RECT 26.32 35.586 26.424 39.96 ; 
      RECT 25.888 35.586 25.992 39.96 ; 
      RECT 25.456 35.586 25.56 39.96 ; 
      RECT 25.024 35.586 25.128 39.96 ; 
      RECT 24.592 35.586 24.696 39.96 ; 
      RECT 24.16 35.586 24.264 39.96 ; 
      RECT 23.728 35.586 23.832 39.96 ; 
      RECT 23.296 35.586 23.4 39.96 ; 
      RECT 22.864 35.586 22.968 39.96 ; 
      RECT 22.432 35.586 22.536 39.96 ; 
      RECT 22 35.586 22.104 39.96 ; 
      RECT 21.568 35.586 21.672 39.96 ; 
      RECT 21.136 35.586 21.24 39.96 ; 
      RECT 20.704 35.586 20.808 39.96 ; 
      RECT 20.272 35.586 20.376 39.96 ; 
      RECT 19.84 35.586 19.944 39.96 ; 
      RECT 19.408 35.586 19.512 39.96 ; 
      RECT 18.976 35.586 19.08 39.96 ; 
      RECT 18.544 35.586 18.648 39.96 ; 
      RECT 18.112 35.586 18.216 39.96 ; 
      RECT 17.68 35.586 17.784 39.96 ; 
      RECT 17.248 35.586 17.352 39.96 ; 
      RECT 16.816 35.586 16.92 39.96 ; 
      RECT 16.384 35.586 16.488 39.96 ; 
      RECT 15.952 35.586 16.056 39.96 ; 
      RECT 15.52 35.586 15.624 39.96 ; 
      RECT 15.088 35.586 15.192 39.96 ; 
      RECT 14.656 35.586 14.76 39.96 ; 
      RECT 14.224 35.586 14.328 39.96 ; 
      RECT 13.792 35.586 13.896 39.96 ; 
      RECT 13.36 35.586 13.464 39.96 ; 
      RECT 12.928 35.586 13.032 39.96 ; 
      RECT 12.496 35.586 12.6 39.96 ; 
      RECT 12.064 35.586 12.168 39.96 ; 
      RECT 11.632 35.586 11.736 39.96 ; 
      RECT 11.2 35.586 11.304 39.96 ; 
      RECT 10.768 35.586 10.872 39.96 ; 
      RECT 10.336 35.586 10.44 39.96 ; 
      RECT 9.904 35.586 10.008 39.96 ; 
      RECT 9.472 35.586 9.576 39.96 ; 
      RECT 9.04 35.586 9.144 39.96 ; 
      RECT 8.608 35.586 8.712 39.96 ; 
      RECT 8.176 35.586 8.28 39.96 ; 
      RECT 7.744 35.586 7.848 39.96 ; 
      RECT 7.312 35.586 7.416 39.96 ; 
      RECT 6.88 35.586 6.984 39.96 ; 
      RECT 6.448 35.586 6.552 39.96 ; 
      RECT 6.016 35.586 6.12 39.96 ; 
      RECT 5.584 35.586 5.688 39.96 ; 
      RECT 5.152 35.586 5.256 39.96 ; 
      RECT 4.72 35.586 4.824 39.96 ; 
      RECT 4.288 35.586 4.392 39.96 ; 
      RECT 3.856 35.586 3.96 39.96 ; 
      RECT 3.424 35.586 3.528 39.96 ; 
      RECT 2.992 35.586 3.096 39.96 ; 
      RECT 2.56 35.586 2.664 39.96 ; 
      RECT 2.128 35.586 2.232 39.96 ; 
      RECT 1.696 35.586 1.8 39.96 ; 
      RECT 1.264 35.586 1.368 39.96 ; 
      RECT 0.832 35.586 0.936 39.96 ; 
      RECT 0.02 35.586 0.36 39.96 ; 
      RECT 34.564 39.906 35.076 44.28 ; 
      RECT 34.508 42.568 35.076 43.858 ; 
      RECT 33.916 41.476 34.164 44.28 ; 
      RECT 33.86 42.714 34.164 43.328 ; 
      RECT 33.916 39.906 34.02 44.28 ; 
      RECT 33.916 40.39 34.076 41.348 ; 
      RECT 33.916 39.906 34.164 40.262 ; 
      RECT 32.728 41.708 33.552 44.28 ; 
      RECT 33.448 39.906 33.552 44.28 ; 
      RECT 32.728 42.816 33.608 43.848 ; 
      RECT 32.728 39.906 33.12 44.28 ; 
      RECT 31.06 39.906 31.392 44.28 ; 
      RECT 31.06 40.26 31.448 44.002 ; 
      RECT 65.776 39.906 66.116 44.28 ; 
      RECT 65.2 39.906 65.304 44.28 ; 
      RECT 64.768 39.906 64.872 44.28 ; 
      RECT 64.336 39.906 64.44 44.28 ; 
      RECT 63.904 39.906 64.008 44.28 ; 
      RECT 63.472 39.906 63.576 44.28 ; 
      RECT 63.04 39.906 63.144 44.28 ; 
      RECT 62.608 39.906 62.712 44.28 ; 
      RECT 62.176 39.906 62.28 44.28 ; 
      RECT 61.744 39.906 61.848 44.28 ; 
      RECT 61.312 39.906 61.416 44.28 ; 
      RECT 60.88 39.906 60.984 44.28 ; 
      RECT 60.448 39.906 60.552 44.28 ; 
      RECT 60.016 39.906 60.12 44.28 ; 
      RECT 59.584 39.906 59.688 44.28 ; 
      RECT 59.152 39.906 59.256 44.28 ; 
      RECT 58.72 39.906 58.824 44.28 ; 
      RECT 58.288 39.906 58.392 44.28 ; 
      RECT 57.856 39.906 57.96 44.28 ; 
      RECT 57.424 39.906 57.528 44.28 ; 
      RECT 56.992 39.906 57.096 44.28 ; 
      RECT 56.56 39.906 56.664 44.28 ; 
      RECT 56.128 39.906 56.232 44.28 ; 
      RECT 55.696 39.906 55.8 44.28 ; 
      RECT 55.264 39.906 55.368 44.28 ; 
      RECT 54.832 39.906 54.936 44.28 ; 
      RECT 54.4 39.906 54.504 44.28 ; 
      RECT 53.968 39.906 54.072 44.28 ; 
      RECT 53.536 39.906 53.64 44.28 ; 
      RECT 53.104 39.906 53.208 44.28 ; 
      RECT 52.672 39.906 52.776 44.28 ; 
      RECT 52.24 39.906 52.344 44.28 ; 
      RECT 51.808 39.906 51.912 44.28 ; 
      RECT 51.376 39.906 51.48 44.28 ; 
      RECT 50.944 39.906 51.048 44.28 ; 
      RECT 50.512 39.906 50.616 44.28 ; 
      RECT 50.08 39.906 50.184 44.28 ; 
      RECT 49.648 39.906 49.752 44.28 ; 
      RECT 49.216 39.906 49.32 44.28 ; 
      RECT 48.784 39.906 48.888 44.28 ; 
      RECT 48.352 39.906 48.456 44.28 ; 
      RECT 47.92 39.906 48.024 44.28 ; 
      RECT 47.488 39.906 47.592 44.28 ; 
      RECT 47.056 39.906 47.16 44.28 ; 
      RECT 46.624 39.906 46.728 44.28 ; 
      RECT 46.192 39.906 46.296 44.28 ; 
      RECT 45.76 39.906 45.864 44.28 ; 
      RECT 45.328 39.906 45.432 44.28 ; 
      RECT 44.896 39.906 45 44.28 ; 
      RECT 44.464 39.906 44.568 44.28 ; 
      RECT 44.032 39.906 44.136 44.28 ; 
      RECT 43.6 39.906 43.704 44.28 ; 
      RECT 43.168 39.906 43.272 44.28 ; 
      RECT 42.736 39.906 42.84 44.28 ; 
      RECT 42.304 39.906 42.408 44.28 ; 
      RECT 41.872 39.906 41.976 44.28 ; 
      RECT 41.44 39.906 41.544 44.28 ; 
      RECT 41.008 39.906 41.112 44.28 ; 
      RECT 40.576 39.906 40.68 44.28 ; 
      RECT 40.144 39.906 40.248 44.28 ; 
      RECT 39.712 39.906 39.816 44.28 ; 
      RECT 39.28 39.906 39.384 44.28 ; 
      RECT 38.848 39.906 38.952 44.28 ; 
      RECT 38.416 39.906 38.52 44.28 ; 
      RECT 37.984 39.906 38.088 44.28 ; 
      RECT 37.552 39.906 37.656 44.28 ; 
      RECT 36.7 39.906 37.008 44.28 ; 
      RECT 29.128 39.906 29.436 44.28 ; 
      RECT 28.48 39.906 28.584 44.28 ; 
      RECT 28.048 39.906 28.152 44.28 ; 
      RECT 27.616 39.906 27.72 44.28 ; 
      RECT 27.184 39.906 27.288 44.28 ; 
      RECT 26.752 39.906 26.856 44.28 ; 
      RECT 26.32 39.906 26.424 44.28 ; 
      RECT 25.888 39.906 25.992 44.28 ; 
      RECT 25.456 39.906 25.56 44.28 ; 
      RECT 25.024 39.906 25.128 44.28 ; 
      RECT 24.592 39.906 24.696 44.28 ; 
      RECT 24.16 39.906 24.264 44.28 ; 
      RECT 23.728 39.906 23.832 44.28 ; 
      RECT 23.296 39.906 23.4 44.28 ; 
      RECT 22.864 39.906 22.968 44.28 ; 
      RECT 22.432 39.906 22.536 44.28 ; 
      RECT 22 39.906 22.104 44.28 ; 
      RECT 21.568 39.906 21.672 44.28 ; 
      RECT 21.136 39.906 21.24 44.28 ; 
      RECT 20.704 39.906 20.808 44.28 ; 
      RECT 20.272 39.906 20.376 44.28 ; 
      RECT 19.84 39.906 19.944 44.28 ; 
      RECT 19.408 39.906 19.512 44.28 ; 
      RECT 18.976 39.906 19.08 44.28 ; 
      RECT 18.544 39.906 18.648 44.28 ; 
      RECT 18.112 39.906 18.216 44.28 ; 
      RECT 17.68 39.906 17.784 44.28 ; 
      RECT 17.248 39.906 17.352 44.28 ; 
      RECT 16.816 39.906 16.92 44.28 ; 
      RECT 16.384 39.906 16.488 44.28 ; 
      RECT 15.952 39.906 16.056 44.28 ; 
      RECT 15.52 39.906 15.624 44.28 ; 
      RECT 15.088 39.906 15.192 44.28 ; 
      RECT 14.656 39.906 14.76 44.28 ; 
      RECT 14.224 39.906 14.328 44.28 ; 
      RECT 13.792 39.906 13.896 44.28 ; 
      RECT 13.36 39.906 13.464 44.28 ; 
      RECT 12.928 39.906 13.032 44.28 ; 
      RECT 12.496 39.906 12.6 44.28 ; 
      RECT 12.064 39.906 12.168 44.28 ; 
      RECT 11.632 39.906 11.736 44.28 ; 
      RECT 11.2 39.906 11.304 44.28 ; 
      RECT 10.768 39.906 10.872 44.28 ; 
      RECT 10.336 39.906 10.44 44.28 ; 
      RECT 9.904 39.906 10.008 44.28 ; 
      RECT 9.472 39.906 9.576 44.28 ; 
      RECT 9.04 39.906 9.144 44.28 ; 
      RECT 8.608 39.906 8.712 44.28 ; 
      RECT 8.176 39.906 8.28 44.28 ; 
      RECT 7.744 39.906 7.848 44.28 ; 
      RECT 7.312 39.906 7.416 44.28 ; 
      RECT 6.88 39.906 6.984 44.28 ; 
      RECT 6.448 39.906 6.552 44.28 ; 
      RECT 6.016 39.906 6.12 44.28 ; 
      RECT 5.584 39.906 5.688 44.28 ; 
      RECT 5.152 39.906 5.256 44.28 ; 
      RECT 4.72 39.906 4.824 44.28 ; 
      RECT 4.288 39.906 4.392 44.28 ; 
      RECT 3.856 39.906 3.96 44.28 ; 
      RECT 3.424 39.906 3.528 44.28 ; 
      RECT 2.992 39.906 3.096 44.28 ; 
      RECT 2.56 39.906 2.664 44.28 ; 
      RECT 2.128 39.906 2.232 44.28 ; 
      RECT 1.696 39.906 1.8 44.28 ; 
      RECT 1.264 39.906 1.368 44.28 ; 
      RECT 0.832 39.906 0.936 44.28 ; 
      RECT 0.02 39.906 0.36 44.28 ; 
      RECT 0 76.998 66.096 78.762 ; 
      RECT 65.756 44.148 66.096 78.762 ; 
      RECT 37.532 50.164 65.284 78.762 ; 
      RECT 43.364 44.148 65.284 78.762 ; 
      RECT 28.892 76.968 37.204 78.762 ; 
      RECT 31.988 76.842 37.204 78.762 ; 
      RECT 0.812 49.384 28.564 78.762 ; 
      RECT 27.38 44.148 28.564 78.762 ; 
      RECT 0 44.148 0.34 78.762 ; 
      RECT 28.892 50.596 31.372 78.762 ; 
      RECT 31.988 76.824 37.06 78.762 ; 
      RECT 34.58 49.768 37.06 78.762 ; 
      RECT 34.544 75.796 37.06 78.762 ; 
      RECT 33.896 75.796 34.144 78.762 ; 
      RECT 31.988 75.796 33.532 78.762 ; 
      RECT 37.532 59.32 65.34 76.736 ; 
      RECT 0.756 59.32 28.564 76.736 ; 
      RECT 37.476 59.32 65.34 76.718 ; 
      RECT 0.756 59.32 28.62 76.718 ; 
      RECT 28.836 59.32 31.372 76.714 ; 
      RECT 32.708 46.888 33.388 78.762 ; 
      RECT 33.14 44.148 33.388 78.762 ; 
      RECT 29.972 45.832 31.516 75.208 ; 
      RECT 28.836 75.028 31.572 75.176 ; 
      RECT 34.524 70.732 37.06 75.164 ; 
      RECT 32.652 73.972 33.388 74.876 ; 
      RECT 32.708 71.668 33.444 72.716 ; 
      RECT 28.836 70.876 31.572 72.716 ; 
      RECT 32.652 68.716 33.388 70.556 ; 
      RECT 34.524 60.58 37.06 69.908 ; 
      RECT 28.836 63.172 31.572 67.748 ; 
      RECT 32.708 62.092 33.444 67.316 ; 
      RECT 32.652 64.396 33.444 66.236 ; 
      RECT 32.652 51.436 33.388 64.076 ; 
      RECT 32.652 51.436 33.444 61.916 ; 
      RECT 28.836 61.012 31.572 61.916 ; 
      RECT 34.58 49.768 37.204 59.192 ; 
      RECT 34.524 49.276 36.988 56.42 ; 
      RECT 28.892 53.164 31.572 54.644 ; 
      RECT 32.708 50.356 33.444 51.116 ; 
      RECT 29.108 50.212 31.572 50.972 ; 
      RECT 32.652 49.78 33.388 50.324 ; 
      RECT 29.108 47.212 31.516 75.208 ; 
      RECT 32.708 49.276 33.444 50.18 ; 
      RECT 38.18 49.396 65.284 78.762 ; 
      RECT 42.5 49.384 65.284 78.762 ; 
      RECT 37.532 44.148 37.852 78.762 ; 
      RECT 28.892 46.888 29.644 50.144 ; 
      RECT 37.532 44.148 38.716 49.76 ; 
      RECT 37.532 48.616 42.172 49.76 ; 
      RECT 42.5 44.148 43.036 78.762 ; 
      RECT 23.924 47.86 27.052 78.762 ; 
      RECT 0.812 44.148 23.596 78.762 ; 
      RECT 34.58 47.212 36.988 78.762 ; 
      RECT 34.724 44.854 37.204 49.148 ; 
      RECT 37.532 48.616 43.036 48.992 ; 
      RECT 41.636 44.148 65.284 48.98 ; 
      RECT 26.516 44.148 28.564 48.98 ; 
      RECT 32.652 48.7 33.444 48.956 ; 
      RECT 32.652 48.196 33.388 48.956 ; 
      RECT 40.772 47.08 65.284 48.98 ; 
      RECT 37.532 47.212 40.444 49.76 ; 
      RECT 32.708 47.116 33.444 48.164 ; 
      RECT 0.812 47.08 26.188 48.98 ; 
      RECT 25.652 44.148 26.188 78.762 ; 
      RECT 39.908 44.148 41.308 47.636 ; 
      RECT 37.532 46.888 39.58 49.76 ; 
      RECT 39.044 44.148 39.58 78.762 ; 
      RECT 24.788 46.888 26.188 78.762 ; 
      RECT 0.812 44.148 24.46 48.98 ; 
      RECT 32.708 44.148 32.812 78.762 ; 
      RECT 29.252 44.148 29.644 78.762 ; 
      RECT 24.788 44.148 25.324 78.762 ; 
      RECT 39.044 44.148 41.308 46.688 ; 
      RECT 34.58 44.148 36.988 46.688 ; 
      RECT 29.252 44.148 31.372 46.688 ; 
      RECT 25.652 44.148 28.564 46.688 ; 
      RECT 39.044 44.148 65.284 46.676 ; 
      RECT 0.812 44.148 25.324 46.676 ; 
      RECT 34.524 46.036 37.204 46.652 ; 
      RECT 37.532 44.148 65.284 45.62 ; 
      RECT 32.708 44.148 33.388 45.62 ; 
      RECT 28.892 44.148 31.372 45.62 ; 
      RECT 0.812 44.148 28.564 45.62 ; 
      RECT 31.988 44.148 33.388 45.208 ; 
      RECT 34.544 44.148 36.988 44.808 ; 
      RECT 31.988 44.148 33.532 44.808 ; 
      RECT 39.06 44.042 39.132 78.762 ; 
      RECT 38.628 44.042 38.7 78.762 ; 
      RECT 27.396 44.092 27.468 78.762 ; 
      RECT 26.964 44.092 27.036 78.762 ; 
      RECT 26.532 44.092 26.604 78.762 ; 
      RECT 26.1 44.092 26.172 78.762 ; 
      RECT 25.668 44.042 25.74 78.762 ; 
      RECT 25.236 44.042 25.308 78.762 ; 
      RECT 24.804 44.092 24.876 78.762 ; 
      RECT 24.372 44.092 24.444 78.762 ; 
      RECT 23.94 44.092 24.012 78.762 ; 
      RECT 23.508 44.092 23.58 78.762 ; 
      RECT 33.896 44.148 34.144 44.808 ; 
        RECT 34.564 76.734 35.076 81.108 ; 
        RECT 34.508 79.396 35.076 80.686 ; 
        RECT 33.916 78.304 34.164 81.108 ; 
        RECT 33.86 79.542 34.164 80.156 ; 
        RECT 33.916 76.734 34.02 81.108 ; 
        RECT 33.916 77.218 34.076 78.176 ; 
        RECT 33.916 76.734 34.164 77.09 ; 
        RECT 32.728 78.536 33.552 81.108 ; 
        RECT 33.448 76.734 33.552 81.108 ; 
        RECT 32.728 79.644 33.608 80.676 ; 
        RECT 32.728 76.734 33.12 81.108 ; 
        RECT 31.06 76.734 31.392 81.108 ; 
        RECT 31.06 77.088 31.448 80.83 ; 
        RECT 65.776 76.734 66.116 81.108 ; 
        RECT 65.2 76.734 65.304 81.108 ; 
        RECT 64.768 76.734 64.872 81.108 ; 
        RECT 64.336 76.734 64.44 81.108 ; 
        RECT 63.904 76.734 64.008 81.108 ; 
        RECT 63.472 76.734 63.576 81.108 ; 
        RECT 63.04 76.734 63.144 81.108 ; 
        RECT 62.608 76.734 62.712 81.108 ; 
        RECT 62.176 76.734 62.28 81.108 ; 
        RECT 61.744 76.734 61.848 81.108 ; 
        RECT 61.312 76.734 61.416 81.108 ; 
        RECT 60.88 76.734 60.984 81.108 ; 
        RECT 60.448 76.734 60.552 81.108 ; 
        RECT 60.016 76.734 60.12 81.108 ; 
        RECT 59.584 76.734 59.688 81.108 ; 
        RECT 59.152 76.734 59.256 81.108 ; 
        RECT 58.72 76.734 58.824 81.108 ; 
        RECT 58.288 76.734 58.392 81.108 ; 
        RECT 57.856 76.734 57.96 81.108 ; 
        RECT 57.424 76.734 57.528 81.108 ; 
        RECT 56.992 76.734 57.096 81.108 ; 
        RECT 56.56 76.734 56.664 81.108 ; 
        RECT 56.128 76.734 56.232 81.108 ; 
        RECT 55.696 76.734 55.8 81.108 ; 
        RECT 55.264 76.734 55.368 81.108 ; 
        RECT 54.832 76.734 54.936 81.108 ; 
        RECT 54.4 76.734 54.504 81.108 ; 
        RECT 53.968 76.734 54.072 81.108 ; 
        RECT 53.536 76.734 53.64 81.108 ; 
        RECT 53.104 76.734 53.208 81.108 ; 
        RECT 52.672 76.734 52.776 81.108 ; 
        RECT 52.24 76.734 52.344 81.108 ; 
        RECT 51.808 76.734 51.912 81.108 ; 
        RECT 51.376 76.734 51.48 81.108 ; 
        RECT 50.944 76.734 51.048 81.108 ; 
        RECT 50.512 76.734 50.616 81.108 ; 
        RECT 50.08 76.734 50.184 81.108 ; 
        RECT 49.648 76.734 49.752 81.108 ; 
        RECT 49.216 76.734 49.32 81.108 ; 
        RECT 48.784 76.734 48.888 81.108 ; 
        RECT 48.352 76.734 48.456 81.108 ; 
        RECT 47.92 76.734 48.024 81.108 ; 
        RECT 47.488 76.734 47.592 81.108 ; 
        RECT 47.056 76.734 47.16 81.108 ; 
        RECT 46.624 76.734 46.728 81.108 ; 
        RECT 46.192 76.734 46.296 81.108 ; 
        RECT 45.76 76.734 45.864 81.108 ; 
        RECT 45.328 76.734 45.432 81.108 ; 
        RECT 44.896 76.734 45 81.108 ; 
        RECT 44.464 76.734 44.568 81.108 ; 
        RECT 44.032 76.734 44.136 81.108 ; 
        RECT 43.6 76.734 43.704 81.108 ; 
        RECT 43.168 76.734 43.272 81.108 ; 
        RECT 42.736 76.734 42.84 81.108 ; 
        RECT 42.304 76.734 42.408 81.108 ; 
        RECT 41.872 76.734 41.976 81.108 ; 
        RECT 41.44 76.734 41.544 81.108 ; 
        RECT 41.008 76.734 41.112 81.108 ; 
        RECT 40.576 76.734 40.68 81.108 ; 
        RECT 40.144 76.734 40.248 81.108 ; 
        RECT 39.712 76.734 39.816 81.108 ; 
        RECT 39.28 76.734 39.384 81.108 ; 
        RECT 38.848 76.734 38.952 81.108 ; 
        RECT 38.416 76.734 38.52 81.108 ; 
        RECT 37.984 76.734 38.088 81.108 ; 
        RECT 37.552 76.734 37.656 81.108 ; 
        RECT 36.7 76.734 37.008 81.108 ; 
        RECT 29.128 76.734 29.436 81.108 ; 
        RECT 28.48 76.734 28.584 81.108 ; 
        RECT 28.048 76.734 28.152 81.108 ; 
        RECT 27.616 76.734 27.72 81.108 ; 
        RECT 27.184 76.734 27.288 81.108 ; 
        RECT 26.752 76.734 26.856 81.108 ; 
        RECT 26.32 76.734 26.424 81.108 ; 
        RECT 25.888 76.734 25.992 81.108 ; 
        RECT 25.456 76.734 25.56 81.108 ; 
        RECT 25.024 76.734 25.128 81.108 ; 
        RECT 24.592 76.734 24.696 81.108 ; 
        RECT 24.16 76.734 24.264 81.108 ; 
        RECT 23.728 76.734 23.832 81.108 ; 
        RECT 23.296 76.734 23.4 81.108 ; 
        RECT 22.864 76.734 22.968 81.108 ; 
        RECT 22.432 76.734 22.536 81.108 ; 
        RECT 22 76.734 22.104 81.108 ; 
        RECT 21.568 76.734 21.672 81.108 ; 
        RECT 21.136 76.734 21.24 81.108 ; 
        RECT 20.704 76.734 20.808 81.108 ; 
        RECT 20.272 76.734 20.376 81.108 ; 
        RECT 19.84 76.734 19.944 81.108 ; 
        RECT 19.408 76.734 19.512 81.108 ; 
        RECT 18.976 76.734 19.08 81.108 ; 
        RECT 18.544 76.734 18.648 81.108 ; 
        RECT 18.112 76.734 18.216 81.108 ; 
        RECT 17.68 76.734 17.784 81.108 ; 
        RECT 17.248 76.734 17.352 81.108 ; 
        RECT 16.816 76.734 16.92 81.108 ; 
        RECT 16.384 76.734 16.488 81.108 ; 
        RECT 15.952 76.734 16.056 81.108 ; 
        RECT 15.52 76.734 15.624 81.108 ; 
        RECT 15.088 76.734 15.192 81.108 ; 
        RECT 14.656 76.734 14.76 81.108 ; 
        RECT 14.224 76.734 14.328 81.108 ; 
        RECT 13.792 76.734 13.896 81.108 ; 
        RECT 13.36 76.734 13.464 81.108 ; 
        RECT 12.928 76.734 13.032 81.108 ; 
        RECT 12.496 76.734 12.6 81.108 ; 
        RECT 12.064 76.734 12.168 81.108 ; 
        RECT 11.632 76.734 11.736 81.108 ; 
        RECT 11.2 76.734 11.304 81.108 ; 
        RECT 10.768 76.734 10.872 81.108 ; 
        RECT 10.336 76.734 10.44 81.108 ; 
        RECT 9.904 76.734 10.008 81.108 ; 
        RECT 9.472 76.734 9.576 81.108 ; 
        RECT 9.04 76.734 9.144 81.108 ; 
        RECT 8.608 76.734 8.712 81.108 ; 
        RECT 8.176 76.734 8.28 81.108 ; 
        RECT 7.744 76.734 7.848 81.108 ; 
        RECT 7.312 76.734 7.416 81.108 ; 
        RECT 6.88 76.734 6.984 81.108 ; 
        RECT 6.448 76.734 6.552 81.108 ; 
        RECT 6.016 76.734 6.12 81.108 ; 
        RECT 5.584 76.734 5.688 81.108 ; 
        RECT 5.152 76.734 5.256 81.108 ; 
        RECT 4.72 76.734 4.824 81.108 ; 
        RECT 4.288 76.734 4.392 81.108 ; 
        RECT 3.856 76.734 3.96 81.108 ; 
        RECT 3.424 76.734 3.528 81.108 ; 
        RECT 2.992 76.734 3.096 81.108 ; 
        RECT 2.56 76.734 2.664 81.108 ; 
        RECT 2.128 76.734 2.232 81.108 ; 
        RECT 1.696 76.734 1.8 81.108 ; 
        RECT 1.264 76.734 1.368 81.108 ; 
        RECT 0.832 76.734 0.936 81.108 ; 
        RECT 0.02 76.734 0.36 81.108 ; 
        RECT 34.564 81.054 35.076 85.428 ; 
        RECT 34.508 83.716 35.076 85.006 ; 
        RECT 33.916 82.624 34.164 85.428 ; 
        RECT 33.86 83.862 34.164 84.476 ; 
        RECT 33.916 81.054 34.02 85.428 ; 
        RECT 33.916 81.538 34.076 82.496 ; 
        RECT 33.916 81.054 34.164 81.41 ; 
        RECT 32.728 82.856 33.552 85.428 ; 
        RECT 33.448 81.054 33.552 85.428 ; 
        RECT 32.728 83.964 33.608 84.996 ; 
        RECT 32.728 81.054 33.12 85.428 ; 
        RECT 31.06 81.054 31.392 85.428 ; 
        RECT 31.06 81.408 31.448 85.15 ; 
        RECT 65.776 81.054 66.116 85.428 ; 
        RECT 65.2 81.054 65.304 85.428 ; 
        RECT 64.768 81.054 64.872 85.428 ; 
        RECT 64.336 81.054 64.44 85.428 ; 
        RECT 63.904 81.054 64.008 85.428 ; 
        RECT 63.472 81.054 63.576 85.428 ; 
        RECT 63.04 81.054 63.144 85.428 ; 
        RECT 62.608 81.054 62.712 85.428 ; 
        RECT 62.176 81.054 62.28 85.428 ; 
        RECT 61.744 81.054 61.848 85.428 ; 
        RECT 61.312 81.054 61.416 85.428 ; 
        RECT 60.88 81.054 60.984 85.428 ; 
        RECT 60.448 81.054 60.552 85.428 ; 
        RECT 60.016 81.054 60.12 85.428 ; 
        RECT 59.584 81.054 59.688 85.428 ; 
        RECT 59.152 81.054 59.256 85.428 ; 
        RECT 58.72 81.054 58.824 85.428 ; 
        RECT 58.288 81.054 58.392 85.428 ; 
        RECT 57.856 81.054 57.96 85.428 ; 
        RECT 57.424 81.054 57.528 85.428 ; 
        RECT 56.992 81.054 57.096 85.428 ; 
        RECT 56.56 81.054 56.664 85.428 ; 
        RECT 56.128 81.054 56.232 85.428 ; 
        RECT 55.696 81.054 55.8 85.428 ; 
        RECT 55.264 81.054 55.368 85.428 ; 
        RECT 54.832 81.054 54.936 85.428 ; 
        RECT 54.4 81.054 54.504 85.428 ; 
        RECT 53.968 81.054 54.072 85.428 ; 
        RECT 53.536 81.054 53.64 85.428 ; 
        RECT 53.104 81.054 53.208 85.428 ; 
        RECT 52.672 81.054 52.776 85.428 ; 
        RECT 52.24 81.054 52.344 85.428 ; 
        RECT 51.808 81.054 51.912 85.428 ; 
        RECT 51.376 81.054 51.48 85.428 ; 
        RECT 50.944 81.054 51.048 85.428 ; 
        RECT 50.512 81.054 50.616 85.428 ; 
        RECT 50.08 81.054 50.184 85.428 ; 
        RECT 49.648 81.054 49.752 85.428 ; 
        RECT 49.216 81.054 49.32 85.428 ; 
        RECT 48.784 81.054 48.888 85.428 ; 
        RECT 48.352 81.054 48.456 85.428 ; 
        RECT 47.92 81.054 48.024 85.428 ; 
        RECT 47.488 81.054 47.592 85.428 ; 
        RECT 47.056 81.054 47.16 85.428 ; 
        RECT 46.624 81.054 46.728 85.428 ; 
        RECT 46.192 81.054 46.296 85.428 ; 
        RECT 45.76 81.054 45.864 85.428 ; 
        RECT 45.328 81.054 45.432 85.428 ; 
        RECT 44.896 81.054 45 85.428 ; 
        RECT 44.464 81.054 44.568 85.428 ; 
        RECT 44.032 81.054 44.136 85.428 ; 
        RECT 43.6 81.054 43.704 85.428 ; 
        RECT 43.168 81.054 43.272 85.428 ; 
        RECT 42.736 81.054 42.84 85.428 ; 
        RECT 42.304 81.054 42.408 85.428 ; 
        RECT 41.872 81.054 41.976 85.428 ; 
        RECT 41.44 81.054 41.544 85.428 ; 
        RECT 41.008 81.054 41.112 85.428 ; 
        RECT 40.576 81.054 40.68 85.428 ; 
        RECT 40.144 81.054 40.248 85.428 ; 
        RECT 39.712 81.054 39.816 85.428 ; 
        RECT 39.28 81.054 39.384 85.428 ; 
        RECT 38.848 81.054 38.952 85.428 ; 
        RECT 38.416 81.054 38.52 85.428 ; 
        RECT 37.984 81.054 38.088 85.428 ; 
        RECT 37.552 81.054 37.656 85.428 ; 
        RECT 36.7 81.054 37.008 85.428 ; 
        RECT 29.128 81.054 29.436 85.428 ; 
        RECT 28.48 81.054 28.584 85.428 ; 
        RECT 28.048 81.054 28.152 85.428 ; 
        RECT 27.616 81.054 27.72 85.428 ; 
        RECT 27.184 81.054 27.288 85.428 ; 
        RECT 26.752 81.054 26.856 85.428 ; 
        RECT 26.32 81.054 26.424 85.428 ; 
        RECT 25.888 81.054 25.992 85.428 ; 
        RECT 25.456 81.054 25.56 85.428 ; 
        RECT 25.024 81.054 25.128 85.428 ; 
        RECT 24.592 81.054 24.696 85.428 ; 
        RECT 24.16 81.054 24.264 85.428 ; 
        RECT 23.728 81.054 23.832 85.428 ; 
        RECT 23.296 81.054 23.4 85.428 ; 
        RECT 22.864 81.054 22.968 85.428 ; 
        RECT 22.432 81.054 22.536 85.428 ; 
        RECT 22 81.054 22.104 85.428 ; 
        RECT 21.568 81.054 21.672 85.428 ; 
        RECT 21.136 81.054 21.24 85.428 ; 
        RECT 20.704 81.054 20.808 85.428 ; 
        RECT 20.272 81.054 20.376 85.428 ; 
        RECT 19.84 81.054 19.944 85.428 ; 
        RECT 19.408 81.054 19.512 85.428 ; 
        RECT 18.976 81.054 19.08 85.428 ; 
        RECT 18.544 81.054 18.648 85.428 ; 
        RECT 18.112 81.054 18.216 85.428 ; 
        RECT 17.68 81.054 17.784 85.428 ; 
        RECT 17.248 81.054 17.352 85.428 ; 
        RECT 16.816 81.054 16.92 85.428 ; 
        RECT 16.384 81.054 16.488 85.428 ; 
        RECT 15.952 81.054 16.056 85.428 ; 
        RECT 15.52 81.054 15.624 85.428 ; 
        RECT 15.088 81.054 15.192 85.428 ; 
        RECT 14.656 81.054 14.76 85.428 ; 
        RECT 14.224 81.054 14.328 85.428 ; 
        RECT 13.792 81.054 13.896 85.428 ; 
        RECT 13.36 81.054 13.464 85.428 ; 
        RECT 12.928 81.054 13.032 85.428 ; 
        RECT 12.496 81.054 12.6 85.428 ; 
        RECT 12.064 81.054 12.168 85.428 ; 
        RECT 11.632 81.054 11.736 85.428 ; 
        RECT 11.2 81.054 11.304 85.428 ; 
        RECT 10.768 81.054 10.872 85.428 ; 
        RECT 10.336 81.054 10.44 85.428 ; 
        RECT 9.904 81.054 10.008 85.428 ; 
        RECT 9.472 81.054 9.576 85.428 ; 
        RECT 9.04 81.054 9.144 85.428 ; 
        RECT 8.608 81.054 8.712 85.428 ; 
        RECT 8.176 81.054 8.28 85.428 ; 
        RECT 7.744 81.054 7.848 85.428 ; 
        RECT 7.312 81.054 7.416 85.428 ; 
        RECT 6.88 81.054 6.984 85.428 ; 
        RECT 6.448 81.054 6.552 85.428 ; 
        RECT 6.016 81.054 6.12 85.428 ; 
        RECT 5.584 81.054 5.688 85.428 ; 
        RECT 5.152 81.054 5.256 85.428 ; 
        RECT 4.72 81.054 4.824 85.428 ; 
        RECT 4.288 81.054 4.392 85.428 ; 
        RECT 3.856 81.054 3.96 85.428 ; 
        RECT 3.424 81.054 3.528 85.428 ; 
        RECT 2.992 81.054 3.096 85.428 ; 
        RECT 2.56 81.054 2.664 85.428 ; 
        RECT 2.128 81.054 2.232 85.428 ; 
        RECT 1.696 81.054 1.8 85.428 ; 
        RECT 1.264 81.054 1.368 85.428 ; 
        RECT 0.832 81.054 0.936 85.428 ; 
        RECT 0.02 81.054 0.36 85.428 ; 
        RECT 34.564 85.374 35.076 89.748 ; 
        RECT 34.508 88.036 35.076 89.326 ; 
        RECT 33.916 86.944 34.164 89.748 ; 
        RECT 33.86 88.182 34.164 88.796 ; 
        RECT 33.916 85.374 34.02 89.748 ; 
        RECT 33.916 85.858 34.076 86.816 ; 
        RECT 33.916 85.374 34.164 85.73 ; 
        RECT 32.728 87.176 33.552 89.748 ; 
        RECT 33.448 85.374 33.552 89.748 ; 
        RECT 32.728 88.284 33.608 89.316 ; 
        RECT 32.728 85.374 33.12 89.748 ; 
        RECT 31.06 85.374 31.392 89.748 ; 
        RECT 31.06 85.728 31.448 89.47 ; 
        RECT 65.776 85.374 66.116 89.748 ; 
        RECT 65.2 85.374 65.304 89.748 ; 
        RECT 64.768 85.374 64.872 89.748 ; 
        RECT 64.336 85.374 64.44 89.748 ; 
        RECT 63.904 85.374 64.008 89.748 ; 
        RECT 63.472 85.374 63.576 89.748 ; 
        RECT 63.04 85.374 63.144 89.748 ; 
        RECT 62.608 85.374 62.712 89.748 ; 
        RECT 62.176 85.374 62.28 89.748 ; 
        RECT 61.744 85.374 61.848 89.748 ; 
        RECT 61.312 85.374 61.416 89.748 ; 
        RECT 60.88 85.374 60.984 89.748 ; 
        RECT 60.448 85.374 60.552 89.748 ; 
        RECT 60.016 85.374 60.12 89.748 ; 
        RECT 59.584 85.374 59.688 89.748 ; 
        RECT 59.152 85.374 59.256 89.748 ; 
        RECT 58.72 85.374 58.824 89.748 ; 
        RECT 58.288 85.374 58.392 89.748 ; 
        RECT 57.856 85.374 57.96 89.748 ; 
        RECT 57.424 85.374 57.528 89.748 ; 
        RECT 56.992 85.374 57.096 89.748 ; 
        RECT 56.56 85.374 56.664 89.748 ; 
        RECT 56.128 85.374 56.232 89.748 ; 
        RECT 55.696 85.374 55.8 89.748 ; 
        RECT 55.264 85.374 55.368 89.748 ; 
        RECT 54.832 85.374 54.936 89.748 ; 
        RECT 54.4 85.374 54.504 89.748 ; 
        RECT 53.968 85.374 54.072 89.748 ; 
        RECT 53.536 85.374 53.64 89.748 ; 
        RECT 53.104 85.374 53.208 89.748 ; 
        RECT 52.672 85.374 52.776 89.748 ; 
        RECT 52.24 85.374 52.344 89.748 ; 
        RECT 51.808 85.374 51.912 89.748 ; 
        RECT 51.376 85.374 51.48 89.748 ; 
        RECT 50.944 85.374 51.048 89.748 ; 
        RECT 50.512 85.374 50.616 89.748 ; 
        RECT 50.08 85.374 50.184 89.748 ; 
        RECT 49.648 85.374 49.752 89.748 ; 
        RECT 49.216 85.374 49.32 89.748 ; 
        RECT 48.784 85.374 48.888 89.748 ; 
        RECT 48.352 85.374 48.456 89.748 ; 
        RECT 47.92 85.374 48.024 89.748 ; 
        RECT 47.488 85.374 47.592 89.748 ; 
        RECT 47.056 85.374 47.16 89.748 ; 
        RECT 46.624 85.374 46.728 89.748 ; 
        RECT 46.192 85.374 46.296 89.748 ; 
        RECT 45.76 85.374 45.864 89.748 ; 
        RECT 45.328 85.374 45.432 89.748 ; 
        RECT 44.896 85.374 45 89.748 ; 
        RECT 44.464 85.374 44.568 89.748 ; 
        RECT 44.032 85.374 44.136 89.748 ; 
        RECT 43.6 85.374 43.704 89.748 ; 
        RECT 43.168 85.374 43.272 89.748 ; 
        RECT 42.736 85.374 42.84 89.748 ; 
        RECT 42.304 85.374 42.408 89.748 ; 
        RECT 41.872 85.374 41.976 89.748 ; 
        RECT 41.44 85.374 41.544 89.748 ; 
        RECT 41.008 85.374 41.112 89.748 ; 
        RECT 40.576 85.374 40.68 89.748 ; 
        RECT 40.144 85.374 40.248 89.748 ; 
        RECT 39.712 85.374 39.816 89.748 ; 
        RECT 39.28 85.374 39.384 89.748 ; 
        RECT 38.848 85.374 38.952 89.748 ; 
        RECT 38.416 85.374 38.52 89.748 ; 
        RECT 37.984 85.374 38.088 89.748 ; 
        RECT 37.552 85.374 37.656 89.748 ; 
        RECT 36.7 85.374 37.008 89.748 ; 
        RECT 29.128 85.374 29.436 89.748 ; 
        RECT 28.48 85.374 28.584 89.748 ; 
        RECT 28.048 85.374 28.152 89.748 ; 
        RECT 27.616 85.374 27.72 89.748 ; 
        RECT 27.184 85.374 27.288 89.748 ; 
        RECT 26.752 85.374 26.856 89.748 ; 
        RECT 26.32 85.374 26.424 89.748 ; 
        RECT 25.888 85.374 25.992 89.748 ; 
        RECT 25.456 85.374 25.56 89.748 ; 
        RECT 25.024 85.374 25.128 89.748 ; 
        RECT 24.592 85.374 24.696 89.748 ; 
        RECT 24.16 85.374 24.264 89.748 ; 
        RECT 23.728 85.374 23.832 89.748 ; 
        RECT 23.296 85.374 23.4 89.748 ; 
        RECT 22.864 85.374 22.968 89.748 ; 
        RECT 22.432 85.374 22.536 89.748 ; 
        RECT 22 85.374 22.104 89.748 ; 
        RECT 21.568 85.374 21.672 89.748 ; 
        RECT 21.136 85.374 21.24 89.748 ; 
        RECT 20.704 85.374 20.808 89.748 ; 
        RECT 20.272 85.374 20.376 89.748 ; 
        RECT 19.84 85.374 19.944 89.748 ; 
        RECT 19.408 85.374 19.512 89.748 ; 
        RECT 18.976 85.374 19.08 89.748 ; 
        RECT 18.544 85.374 18.648 89.748 ; 
        RECT 18.112 85.374 18.216 89.748 ; 
        RECT 17.68 85.374 17.784 89.748 ; 
        RECT 17.248 85.374 17.352 89.748 ; 
        RECT 16.816 85.374 16.92 89.748 ; 
        RECT 16.384 85.374 16.488 89.748 ; 
        RECT 15.952 85.374 16.056 89.748 ; 
        RECT 15.52 85.374 15.624 89.748 ; 
        RECT 15.088 85.374 15.192 89.748 ; 
        RECT 14.656 85.374 14.76 89.748 ; 
        RECT 14.224 85.374 14.328 89.748 ; 
        RECT 13.792 85.374 13.896 89.748 ; 
        RECT 13.36 85.374 13.464 89.748 ; 
        RECT 12.928 85.374 13.032 89.748 ; 
        RECT 12.496 85.374 12.6 89.748 ; 
        RECT 12.064 85.374 12.168 89.748 ; 
        RECT 11.632 85.374 11.736 89.748 ; 
        RECT 11.2 85.374 11.304 89.748 ; 
        RECT 10.768 85.374 10.872 89.748 ; 
        RECT 10.336 85.374 10.44 89.748 ; 
        RECT 9.904 85.374 10.008 89.748 ; 
        RECT 9.472 85.374 9.576 89.748 ; 
        RECT 9.04 85.374 9.144 89.748 ; 
        RECT 8.608 85.374 8.712 89.748 ; 
        RECT 8.176 85.374 8.28 89.748 ; 
        RECT 7.744 85.374 7.848 89.748 ; 
        RECT 7.312 85.374 7.416 89.748 ; 
        RECT 6.88 85.374 6.984 89.748 ; 
        RECT 6.448 85.374 6.552 89.748 ; 
        RECT 6.016 85.374 6.12 89.748 ; 
        RECT 5.584 85.374 5.688 89.748 ; 
        RECT 5.152 85.374 5.256 89.748 ; 
        RECT 4.72 85.374 4.824 89.748 ; 
        RECT 4.288 85.374 4.392 89.748 ; 
        RECT 3.856 85.374 3.96 89.748 ; 
        RECT 3.424 85.374 3.528 89.748 ; 
        RECT 2.992 85.374 3.096 89.748 ; 
        RECT 2.56 85.374 2.664 89.748 ; 
        RECT 2.128 85.374 2.232 89.748 ; 
        RECT 1.696 85.374 1.8 89.748 ; 
        RECT 1.264 85.374 1.368 89.748 ; 
        RECT 0.832 85.374 0.936 89.748 ; 
        RECT 0.02 85.374 0.36 89.748 ; 
        RECT 34.564 89.694 35.076 94.068 ; 
        RECT 34.508 92.356 35.076 93.646 ; 
        RECT 33.916 91.264 34.164 94.068 ; 
        RECT 33.86 92.502 34.164 93.116 ; 
        RECT 33.916 89.694 34.02 94.068 ; 
        RECT 33.916 90.178 34.076 91.136 ; 
        RECT 33.916 89.694 34.164 90.05 ; 
        RECT 32.728 91.496 33.552 94.068 ; 
        RECT 33.448 89.694 33.552 94.068 ; 
        RECT 32.728 92.604 33.608 93.636 ; 
        RECT 32.728 89.694 33.12 94.068 ; 
        RECT 31.06 89.694 31.392 94.068 ; 
        RECT 31.06 90.048 31.448 93.79 ; 
        RECT 65.776 89.694 66.116 94.068 ; 
        RECT 65.2 89.694 65.304 94.068 ; 
        RECT 64.768 89.694 64.872 94.068 ; 
        RECT 64.336 89.694 64.44 94.068 ; 
        RECT 63.904 89.694 64.008 94.068 ; 
        RECT 63.472 89.694 63.576 94.068 ; 
        RECT 63.04 89.694 63.144 94.068 ; 
        RECT 62.608 89.694 62.712 94.068 ; 
        RECT 62.176 89.694 62.28 94.068 ; 
        RECT 61.744 89.694 61.848 94.068 ; 
        RECT 61.312 89.694 61.416 94.068 ; 
        RECT 60.88 89.694 60.984 94.068 ; 
        RECT 60.448 89.694 60.552 94.068 ; 
        RECT 60.016 89.694 60.12 94.068 ; 
        RECT 59.584 89.694 59.688 94.068 ; 
        RECT 59.152 89.694 59.256 94.068 ; 
        RECT 58.72 89.694 58.824 94.068 ; 
        RECT 58.288 89.694 58.392 94.068 ; 
        RECT 57.856 89.694 57.96 94.068 ; 
        RECT 57.424 89.694 57.528 94.068 ; 
        RECT 56.992 89.694 57.096 94.068 ; 
        RECT 56.56 89.694 56.664 94.068 ; 
        RECT 56.128 89.694 56.232 94.068 ; 
        RECT 55.696 89.694 55.8 94.068 ; 
        RECT 55.264 89.694 55.368 94.068 ; 
        RECT 54.832 89.694 54.936 94.068 ; 
        RECT 54.4 89.694 54.504 94.068 ; 
        RECT 53.968 89.694 54.072 94.068 ; 
        RECT 53.536 89.694 53.64 94.068 ; 
        RECT 53.104 89.694 53.208 94.068 ; 
        RECT 52.672 89.694 52.776 94.068 ; 
        RECT 52.24 89.694 52.344 94.068 ; 
        RECT 51.808 89.694 51.912 94.068 ; 
        RECT 51.376 89.694 51.48 94.068 ; 
        RECT 50.944 89.694 51.048 94.068 ; 
        RECT 50.512 89.694 50.616 94.068 ; 
        RECT 50.08 89.694 50.184 94.068 ; 
        RECT 49.648 89.694 49.752 94.068 ; 
        RECT 49.216 89.694 49.32 94.068 ; 
        RECT 48.784 89.694 48.888 94.068 ; 
        RECT 48.352 89.694 48.456 94.068 ; 
        RECT 47.92 89.694 48.024 94.068 ; 
        RECT 47.488 89.694 47.592 94.068 ; 
        RECT 47.056 89.694 47.16 94.068 ; 
        RECT 46.624 89.694 46.728 94.068 ; 
        RECT 46.192 89.694 46.296 94.068 ; 
        RECT 45.76 89.694 45.864 94.068 ; 
        RECT 45.328 89.694 45.432 94.068 ; 
        RECT 44.896 89.694 45 94.068 ; 
        RECT 44.464 89.694 44.568 94.068 ; 
        RECT 44.032 89.694 44.136 94.068 ; 
        RECT 43.6 89.694 43.704 94.068 ; 
        RECT 43.168 89.694 43.272 94.068 ; 
        RECT 42.736 89.694 42.84 94.068 ; 
        RECT 42.304 89.694 42.408 94.068 ; 
        RECT 41.872 89.694 41.976 94.068 ; 
        RECT 41.44 89.694 41.544 94.068 ; 
        RECT 41.008 89.694 41.112 94.068 ; 
        RECT 40.576 89.694 40.68 94.068 ; 
        RECT 40.144 89.694 40.248 94.068 ; 
        RECT 39.712 89.694 39.816 94.068 ; 
        RECT 39.28 89.694 39.384 94.068 ; 
        RECT 38.848 89.694 38.952 94.068 ; 
        RECT 38.416 89.694 38.52 94.068 ; 
        RECT 37.984 89.694 38.088 94.068 ; 
        RECT 37.552 89.694 37.656 94.068 ; 
        RECT 36.7 89.694 37.008 94.068 ; 
        RECT 29.128 89.694 29.436 94.068 ; 
        RECT 28.48 89.694 28.584 94.068 ; 
        RECT 28.048 89.694 28.152 94.068 ; 
        RECT 27.616 89.694 27.72 94.068 ; 
        RECT 27.184 89.694 27.288 94.068 ; 
        RECT 26.752 89.694 26.856 94.068 ; 
        RECT 26.32 89.694 26.424 94.068 ; 
        RECT 25.888 89.694 25.992 94.068 ; 
        RECT 25.456 89.694 25.56 94.068 ; 
        RECT 25.024 89.694 25.128 94.068 ; 
        RECT 24.592 89.694 24.696 94.068 ; 
        RECT 24.16 89.694 24.264 94.068 ; 
        RECT 23.728 89.694 23.832 94.068 ; 
        RECT 23.296 89.694 23.4 94.068 ; 
        RECT 22.864 89.694 22.968 94.068 ; 
        RECT 22.432 89.694 22.536 94.068 ; 
        RECT 22 89.694 22.104 94.068 ; 
        RECT 21.568 89.694 21.672 94.068 ; 
        RECT 21.136 89.694 21.24 94.068 ; 
        RECT 20.704 89.694 20.808 94.068 ; 
        RECT 20.272 89.694 20.376 94.068 ; 
        RECT 19.84 89.694 19.944 94.068 ; 
        RECT 19.408 89.694 19.512 94.068 ; 
        RECT 18.976 89.694 19.08 94.068 ; 
        RECT 18.544 89.694 18.648 94.068 ; 
        RECT 18.112 89.694 18.216 94.068 ; 
        RECT 17.68 89.694 17.784 94.068 ; 
        RECT 17.248 89.694 17.352 94.068 ; 
        RECT 16.816 89.694 16.92 94.068 ; 
        RECT 16.384 89.694 16.488 94.068 ; 
        RECT 15.952 89.694 16.056 94.068 ; 
        RECT 15.52 89.694 15.624 94.068 ; 
        RECT 15.088 89.694 15.192 94.068 ; 
        RECT 14.656 89.694 14.76 94.068 ; 
        RECT 14.224 89.694 14.328 94.068 ; 
        RECT 13.792 89.694 13.896 94.068 ; 
        RECT 13.36 89.694 13.464 94.068 ; 
        RECT 12.928 89.694 13.032 94.068 ; 
        RECT 12.496 89.694 12.6 94.068 ; 
        RECT 12.064 89.694 12.168 94.068 ; 
        RECT 11.632 89.694 11.736 94.068 ; 
        RECT 11.2 89.694 11.304 94.068 ; 
        RECT 10.768 89.694 10.872 94.068 ; 
        RECT 10.336 89.694 10.44 94.068 ; 
        RECT 9.904 89.694 10.008 94.068 ; 
        RECT 9.472 89.694 9.576 94.068 ; 
        RECT 9.04 89.694 9.144 94.068 ; 
        RECT 8.608 89.694 8.712 94.068 ; 
        RECT 8.176 89.694 8.28 94.068 ; 
        RECT 7.744 89.694 7.848 94.068 ; 
        RECT 7.312 89.694 7.416 94.068 ; 
        RECT 6.88 89.694 6.984 94.068 ; 
        RECT 6.448 89.694 6.552 94.068 ; 
        RECT 6.016 89.694 6.12 94.068 ; 
        RECT 5.584 89.694 5.688 94.068 ; 
        RECT 5.152 89.694 5.256 94.068 ; 
        RECT 4.72 89.694 4.824 94.068 ; 
        RECT 4.288 89.694 4.392 94.068 ; 
        RECT 3.856 89.694 3.96 94.068 ; 
        RECT 3.424 89.694 3.528 94.068 ; 
        RECT 2.992 89.694 3.096 94.068 ; 
        RECT 2.56 89.694 2.664 94.068 ; 
        RECT 2.128 89.694 2.232 94.068 ; 
        RECT 1.696 89.694 1.8 94.068 ; 
        RECT 1.264 89.694 1.368 94.068 ; 
        RECT 0.832 89.694 0.936 94.068 ; 
        RECT 0.02 89.694 0.36 94.068 ; 
        RECT 34.564 94.014 35.076 98.388 ; 
        RECT 34.508 96.676 35.076 97.966 ; 
        RECT 33.916 95.584 34.164 98.388 ; 
        RECT 33.86 96.822 34.164 97.436 ; 
        RECT 33.916 94.014 34.02 98.388 ; 
        RECT 33.916 94.498 34.076 95.456 ; 
        RECT 33.916 94.014 34.164 94.37 ; 
        RECT 32.728 95.816 33.552 98.388 ; 
        RECT 33.448 94.014 33.552 98.388 ; 
        RECT 32.728 96.924 33.608 97.956 ; 
        RECT 32.728 94.014 33.12 98.388 ; 
        RECT 31.06 94.014 31.392 98.388 ; 
        RECT 31.06 94.368 31.448 98.11 ; 
        RECT 65.776 94.014 66.116 98.388 ; 
        RECT 65.2 94.014 65.304 98.388 ; 
        RECT 64.768 94.014 64.872 98.388 ; 
        RECT 64.336 94.014 64.44 98.388 ; 
        RECT 63.904 94.014 64.008 98.388 ; 
        RECT 63.472 94.014 63.576 98.388 ; 
        RECT 63.04 94.014 63.144 98.388 ; 
        RECT 62.608 94.014 62.712 98.388 ; 
        RECT 62.176 94.014 62.28 98.388 ; 
        RECT 61.744 94.014 61.848 98.388 ; 
        RECT 61.312 94.014 61.416 98.388 ; 
        RECT 60.88 94.014 60.984 98.388 ; 
        RECT 60.448 94.014 60.552 98.388 ; 
        RECT 60.016 94.014 60.12 98.388 ; 
        RECT 59.584 94.014 59.688 98.388 ; 
        RECT 59.152 94.014 59.256 98.388 ; 
        RECT 58.72 94.014 58.824 98.388 ; 
        RECT 58.288 94.014 58.392 98.388 ; 
        RECT 57.856 94.014 57.96 98.388 ; 
        RECT 57.424 94.014 57.528 98.388 ; 
        RECT 56.992 94.014 57.096 98.388 ; 
        RECT 56.56 94.014 56.664 98.388 ; 
        RECT 56.128 94.014 56.232 98.388 ; 
        RECT 55.696 94.014 55.8 98.388 ; 
        RECT 55.264 94.014 55.368 98.388 ; 
        RECT 54.832 94.014 54.936 98.388 ; 
        RECT 54.4 94.014 54.504 98.388 ; 
        RECT 53.968 94.014 54.072 98.388 ; 
        RECT 53.536 94.014 53.64 98.388 ; 
        RECT 53.104 94.014 53.208 98.388 ; 
        RECT 52.672 94.014 52.776 98.388 ; 
        RECT 52.24 94.014 52.344 98.388 ; 
        RECT 51.808 94.014 51.912 98.388 ; 
        RECT 51.376 94.014 51.48 98.388 ; 
        RECT 50.944 94.014 51.048 98.388 ; 
        RECT 50.512 94.014 50.616 98.388 ; 
        RECT 50.08 94.014 50.184 98.388 ; 
        RECT 49.648 94.014 49.752 98.388 ; 
        RECT 49.216 94.014 49.32 98.388 ; 
        RECT 48.784 94.014 48.888 98.388 ; 
        RECT 48.352 94.014 48.456 98.388 ; 
        RECT 47.92 94.014 48.024 98.388 ; 
        RECT 47.488 94.014 47.592 98.388 ; 
        RECT 47.056 94.014 47.16 98.388 ; 
        RECT 46.624 94.014 46.728 98.388 ; 
        RECT 46.192 94.014 46.296 98.388 ; 
        RECT 45.76 94.014 45.864 98.388 ; 
        RECT 45.328 94.014 45.432 98.388 ; 
        RECT 44.896 94.014 45 98.388 ; 
        RECT 44.464 94.014 44.568 98.388 ; 
        RECT 44.032 94.014 44.136 98.388 ; 
        RECT 43.6 94.014 43.704 98.388 ; 
        RECT 43.168 94.014 43.272 98.388 ; 
        RECT 42.736 94.014 42.84 98.388 ; 
        RECT 42.304 94.014 42.408 98.388 ; 
        RECT 41.872 94.014 41.976 98.388 ; 
        RECT 41.44 94.014 41.544 98.388 ; 
        RECT 41.008 94.014 41.112 98.388 ; 
        RECT 40.576 94.014 40.68 98.388 ; 
        RECT 40.144 94.014 40.248 98.388 ; 
        RECT 39.712 94.014 39.816 98.388 ; 
        RECT 39.28 94.014 39.384 98.388 ; 
        RECT 38.848 94.014 38.952 98.388 ; 
        RECT 38.416 94.014 38.52 98.388 ; 
        RECT 37.984 94.014 38.088 98.388 ; 
        RECT 37.552 94.014 37.656 98.388 ; 
        RECT 36.7 94.014 37.008 98.388 ; 
        RECT 29.128 94.014 29.436 98.388 ; 
        RECT 28.48 94.014 28.584 98.388 ; 
        RECT 28.048 94.014 28.152 98.388 ; 
        RECT 27.616 94.014 27.72 98.388 ; 
        RECT 27.184 94.014 27.288 98.388 ; 
        RECT 26.752 94.014 26.856 98.388 ; 
        RECT 26.32 94.014 26.424 98.388 ; 
        RECT 25.888 94.014 25.992 98.388 ; 
        RECT 25.456 94.014 25.56 98.388 ; 
        RECT 25.024 94.014 25.128 98.388 ; 
        RECT 24.592 94.014 24.696 98.388 ; 
        RECT 24.16 94.014 24.264 98.388 ; 
        RECT 23.728 94.014 23.832 98.388 ; 
        RECT 23.296 94.014 23.4 98.388 ; 
        RECT 22.864 94.014 22.968 98.388 ; 
        RECT 22.432 94.014 22.536 98.388 ; 
        RECT 22 94.014 22.104 98.388 ; 
        RECT 21.568 94.014 21.672 98.388 ; 
        RECT 21.136 94.014 21.24 98.388 ; 
        RECT 20.704 94.014 20.808 98.388 ; 
        RECT 20.272 94.014 20.376 98.388 ; 
        RECT 19.84 94.014 19.944 98.388 ; 
        RECT 19.408 94.014 19.512 98.388 ; 
        RECT 18.976 94.014 19.08 98.388 ; 
        RECT 18.544 94.014 18.648 98.388 ; 
        RECT 18.112 94.014 18.216 98.388 ; 
        RECT 17.68 94.014 17.784 98.388 ; 
        RECT 17.248 94.014 17.352 98.388 ; 
        RECT 16.816 94.014 16.92 98.388 ; 
        RECT 16.384 94.014 16.488 98.388 ; 
        RECT 15.952 94.014 16.056 98.388 ; 
        RECT 15.52 94.014 15.624 98.388 ; 
        RECT 15.088 94.014 15.192 98.388 ; 
        RECT 14.656 94.014 14.76 98.388 ; 
        RECT 14.224 94.014 14.328 98.388 ; 
        RECT 13.792 94.014 13.896 98.388 ; 
        RECT 13.36 94.014 13.464 98.388 ; 
        RECT 12.928 94.014 13.032 98.388 ; 
        RECT 12.496 94.014 12.6 98.388 ; 
        RECT 12.064 94.014 12.168 98.388 ; 
        RECT 11.632 94.014 11.736 98.388 ; 
        RECT 11.2 94.014 11.304 98.388 ; 
        RECT 10.768 94.014 10.872 98.388 ; 
        RECT 10.336 94.014 10.44 98.388 ; 
        RECT 9.904 94.014 10.008 98.388 ; 
        RECT 9.472 94.014 9.576 98.388 ; 
        RECT 9.04 94.014 9.144 98.388 ; 
        RECT 8.608 94.014 8.712 98.388 ; 
        RECT 8.176 94.014 8.28 98.388 ; 
        RECT 7.744 94.014 7.848 98.388 ; 
        RECT 7.312 94.014 7.416 98.388 ; 
        RECT 6.88 94.014 6.984 98.388 ; 
        RECT 6.448 94.014 6.552 98.388 ; 
        RECT 6.016 94.014 6.12 98.388 ; 
        RECT 5.584 94.014 5.688 98.388 ; 
        RECT 5.152 94.014 5.256 98.388 ; 
        RECT 4.72 94.014 4.824 98.388 ; 
        RECT 4.288 94.014 4.392 98.388 ; 
        RECT 3.856 94.014 3.96 98.388 ; 
        RECT 3.424 94.014 3.528 98.388 ; 
        RECT 2.992 94.014 3.096 98.388 ; 
        RECT 2.56 94.014 2.664 98.388 ; 
        RECT 2.128 94.014 2.232 98.388 ; 
        RECT 1.696 94.014 1.8 98.388 ; 
        RECT 1.264 94.014 1.368 98.388 ; 
        RECT 0.832 94.014 0.936 98.388 ; 
        RECT 0.02 94.014 0.36 98.388 ; 
        RECT 34.564 98.334 35.076 102.708 ; 
        RECT 34.508 100.996 35.076 102.286 ; 
        RECT 33.916 99.904 34.164 102.708 ; 
        RECT 33.86 101.142 34.164 101.756 ; 
        RECT 33.916 98.334 34.02 102.708 ; 
        RECT 33.916 98.818 34.076 99.776 ; 
        RECT 33.916 98.334 34.164 98.69 ; 
        RECT 32.728 100.136 33.552 102.708 ; 
        RECT 33.448 98.334 33.552 102.708 ; 
        RECT 32.728 101.244 33.608 102.276 ; 
        RECT 32.728 98.334 33.12 102.708 ; 
        RECT 31.06 98.334 31.392 102.708 ; 
        RECT 31.06 98.688 31.448 102.43 ; 
        RECT 65.776 98.334 66.116 102.708 ; 
        RECT 65.2 98.334 65.304 102.708 ; 
        RECT 64.768 98.334 64.872 102.708 ; 
        RECT 64.336 98.334 64.44 102.708 ; 
        RECT 63.904 98.334 64.008 102.708 ; 
        RECT 63.472 98.334 63.576 102.708 ; 
        RECT 63.04 98.334 63.144 102.708 ; 
        RECT 62.608 98.334 62.712 102.708 ; 
        RECT 62.176 98.334 62.28 102.708 ; 
        RECT 61.744 98.334 61.848 102.708 ; 
        RECT 61.312 98.334 61.416 102.708 ; 
        RECT 60.88 98.334 60.984 102.708 ; 
        RECT 60.448 98.334 60.552 102.708 ; 
        RECT 60.016 98.334 60.12 102.708 ; 
        RECT 59.584 98.334 59.688 102.708 ; 
        RECT 59.152 98.334 59.256 102.708 ; 
        RECT 58.72 98.334 58.824 102.708 ; 
        RECT 58.288 98.334 58.392 102.708 ; 
        RECT 57.856 98.334 57.96 102.708 ; 
        RECT 57.424 98.334 57.528 102.708 ; 
        RECT 56.992 98.334 57.096 102.708 ; 
        RECT 56.56 98.334 56.664 102.708 ; 
        RECT 56.128 98.334 56.232 102.708 ; 
        RECT 55.696 98.334 55.8 102.708 ; 
        RECT 55.264 98.334 55.368 102.708 ; 
        RECT 54.832 98.334 54.936 102.708 ; 
        RECT 54.4 98.334 54.504 102.708 ; 
        RECT 53.968 98.334 54.072 102.708 ; 
        RECT 53.536 98.334 53.64 102.708 ; 
        RECT 53.104 98.334 53.208 102.708 ; 
        RECT 52.672 98.334 52.776 102.708 ; 
        RECT 52.24 98.334 52.344 102.708 ; 
        RECT 51.808 98.334 51.912 102.708 ; 
        RECT 51.376 98.334 51.48 102.708 ; 
        RECT 50.944 98.334 51.048 102.708 ; 
        RECT 50.512 98.334 50.616 102.708 ; 
        RECT 50.08 98.334 50.184 102.708 ; 
        RECT 49.648 98.334 49.752 102.708 ; 
        RECT 49.216 98.334 49.32 102.708 ; 
        RECT 48.784 98.334 48.888 102.708 ; 
        RECT 48.352 98.334 48.456 102.708 ; 
        RECT 47.92 98.334 48.024 102.708 ; 
        RECT 47.488 98.334 47.592 102.708 ; 
        RECT 47.056 98.334 47.16 102.708 ; 
        RECT 46.624 98.334 46.728 102.708 ; 
        RECT 46.192 98.334 46.296 102.708 ; 
        RECT 45.76 98.334 45.864 102.708 ; 
        RECT 45.328 98.334 45.432 102.708 ; 
        RECT 44.896 98.334 45 102.708 ; 
        RECT 44.464 98.334 44.568 102.708 ; 
        RECT 44.032 98.334 44.136 102.708 ; 
        RECT 43.6 98.334 43.704 102.708 ; 
        RECT 43.168 98.334 43.272 102.708 ; 
        RECT 42.736 98.334 42.84 102.708 ; 
        RECT 42.304 98.334 42.408 102.708 ; 
        RECT 41.872 98.334 41.976 102.708 ; 
        RECT 41.44 98.334 41.544 102.708 ; 
        RECT 41.008 98.334 41.112 102.708 ; 
        RECT 40.576 98.334 40.68 102.708 ; 
        RECT 40.144 98.334 40.248 102.708 ; 
        RECT 39.712 98.334 39.816 102.708 ; 
        RECT 39.28 98.334 39.384 102.708 ; 
        RECT 38.848 98.334 38.952 102.708 ; 
        RECT 38.416 98.334 38.52 102.708 ; 
        RECT 37.984 98.334 38.088 102.708 ; 
        RECT 37.552 98.334 37.656 102.708 ; 
        RECT 36.7 98.334 37.008 102.708 ; 
        RECT 29.128 98.334 29.436 102.708 ; 
        RECT 28.48 98.334 28.584 102.708 ; 
        RECT 28.048 98.334 28.152 102.708 ; 
        RECT 27.616 98.334 27.72 102.708 ; 
        RECT 27.184 98.334 27.288 102.708 ; 
        RECT 26.752 98.334 26.856 102.708 ; 
        RECT 26.32 98.334 26.424 102.708 ; 
        RECT 25.888 98.334 25.992 102.708 ; 
        RECT 25.456 98.334 25.56 102.708 ; 
        RECT 25.024 98.334 25.128 102.708 ; 
        RECT 24.592 98.334 24.696 102.708 ; 
        RECT 24.16 98.334 24.264 102.708 ; 
        RECT 23.728 98.334 23.832 102.708 ; 
        RECT 23.296 98.334 23.4 102.708 ; 
        RECT 22.864 98.334 22.968 102.708 ; 
        RECT 22.432 98.334 22.536 102.708 ; 
        RECT 22 98.334 22.104 102.708 ; 
        RECT 21.568 98.334 21.672 102.708 ; 
        RECT 21.136 98.334 21.24 102.708 ; 
        RECT 20.704 98.334 20.808 102.708 ; 
        RECT 20.272 98.334 20.376 102.708 ; 
        RECT 19.84 98.334 19.944 102.708 ; 
        RECT 19.408 98.334 19.512 102.708 ; 
        RECT 18.976 98.334 19.08 102.708 ; 
        RECT 18.544 98.334 18.648 102.708 ; 
        RECT 18.112 98.334 18.216 102.708 ; 
        RECT 17.68 98.334 17.784 102.708 ; 
        RECT 17.248 98.334 17.352 102.708 ; 
        RECT 16.816 98.334 16.92 102.708 ; 
        RECT 16.384 98.334 16.488 102.708 ; 
        RECT 15.952 98.334 16.056 102.708 ; 
        RECT 15.52 98.334 15.624 102.708 ; 
        RECT 15.088 98.334 15.192 102.708 ; 
        RECT 14.656 98.334 14.76 102.708 ; 
        RECT 14.224 98.334 14.328 102.708 ; 
        RECT 13.792 98.334 13.896 102.708 ; 
        RECT 13.36 98.334 13.464 102.708 ; 
        RECT 12.928 98.334 13.032 102.708 ; 
        RECT 12.496 98.334 12.6 102.708 ; 
        RECT 12.064 98.334 12.168 102.708 ; 
        RECT 11.632 98.334 11.736 102.708 ; 
        RECT 11.2 98.334 11.304 102.708 ; 
        RECT 10.768 98.334 10.872 102.708 ; 
        RECT 10.336 98.334 10.44 102.708 ; 
        RECT 9.904 98.334 10.008 102.708 ; 
        RECT 9.472 98.334 9.576 102.708 ; 
        RECT 9.04 98.334 9.144 102.708 ; 
        RECT 8.608 98.334 8.712 102.708 ; 
        RECT 8.176 98.334 8.28 102.708 ; 
        RECT 7.744 98.334 7.848 102.708 ; 
        RECT 7.312 98.334 7.416 102.708 ; 
        RECT 6.88 98.334 6.984 102.708 ; 
        RECT 6.448 98.334 6.552 102.708 ; 
        RECT 6.016 98.334 6.12 102.708 ; 
        RECT 5.584 98.334 5.688 102.708 ; 
        RECT 5.152 98.334 5.256 102.708 ; 
        RECT 4.72 98.334 4.824 102.708 ; 
        RECT 4.288 98.334 4.392 102.708 ; 
        RECT 3.856 98.334 3.96 102.708 ; 
        RECT 3.424 98.334 3.528 102.708 ; 
        RECT 2.992 98.334 3.096 102.708 ; 
        RECT 2.56 98.334 2.664 102.708 ; 
        RECT 2.128 98.334 2.232 102.708 ; 
        RECT 1.696 98.334 1.8 102.708 ; 
        RECT 1.264 98.334 1.368 102.708 ; 
        RECT 0.832 98.334 0.936 102.708 ; 
        RECT 0.02 98.334 0.36 102.708 ; 
        RECT 34.564 102.654 35.076 107.028 ; 
        RECT 34.508 105.316 35.076 106.606 ; 
        RECT 33.916 104.224 34.164 107.028 ; 
        RECT 33.86 105.462 34.164 106.076 ; 
        RECT 33.916 102.654 34.02 107.028 ; 
        RECT 33.916 103.138 34.076 104.096 ; 
        RECT 33.916 102.654 34.164 103.01 ; 
        RECT 32.728 104.456 33.552 107.028 ; 
        RECT 33.448 102.654 33.552 107.028 ; 
        RECT 32.728 105.564 33.608 106.596 ; 
        RECT 32.728 102.654 33.12 107.028 ; 
        RECT 31.06 102.654 31.392 107.028 ; 
        RECT 31.06 103.008 31.448 106.75 ; 
        RECT 65.776 102.654 66.116 107.028 ; 
        RECT 65.2 102.654 65.304 107.028 ; 
        RECT 64.768 102.654 64.872 107.028 ; 
        RECT 64.336 102.654 64.44 107.028 ; 
        RECT 63.904 102.654 64.008 107.028 ; 
        RECT 63.472 102.654 63.576 107.028 ; 
        RECT 63.04 102.654 63.144 107.028 ; 
        RECT 62.608 102.654 62.712 107.028 ; 
        RECT 62.176 102.654 62.28 107.028 ; 
        RECT 61.744 102.654 61.848 107.028 ; 
        RECT 61.312 102.654 61.416 107.028 ; 
        RECT 60.88 102.654 60.984 107.028 ; 
        RECT 60.448 102.654 60.552 107.028 ; 
        RECT 60.016 102.654 60.12 107.028 ; 
        RECT 59.584 102.654 59.688 107.028 ; 
        RECT 59.152 102.654 59.256 107.028 ; 
        RECT 58.72 102.654 58.824 107.028 ; 
        RECT 58.288 102.654 58.392 107.028 ; 
        RECT 57.856 102.654 57.96 107.028 ; 
        RECT 57.424 102.654 57.528 107.028 ; 
        RECT 56.992 102.654 57.096 107.028 ; 
        RECT 56.56 102.654 56.664 107.028 ; 
        RECT 56.128 102.654 56.232 107.028 ; 
        RECT 55.696 102.654 55.8 107.028 ; 
        RECT 55.264 102.654 55.368 107.028 ; 
        RECT 54.832 102.654 54.936 107.028 ; 
        RECT 54.4 102.654 54.504 107.028 ; 
        RECT 53.968 102.654 54.072 107.028 ; 
        RECT 53.536 102.654 53.64 107.028 ; 
        RECT 53.104 102.654 53.208 107.028 ; 
        RECT 52.672 102.654 52.776 107.028 ; 
        RECT 52.24 102.654 52.344 107.028 ; 
        RECT 51.808 102.654 51.912 107.028 ; 
        RECT 51.376 102.654 51.48 107.028 ; 
        RECT 50.944 102.654 51.048 107.028 ; 
        RECT 50.512 102.654 50.616 107.028 ; 
        RECT 50.08 102.654 50.184 107.028 ; 
        RECT 49.648 102.654 49.752 107.028 ; 
        RECT 49.216 102.654 49.32 107.028 ; 
        RECT 48.784 102.654 48.888 107.028 ; 
        RECT 48.352 102.654 48.456 107.028 ; 
        RECT 47.92 102.654 48.024 107.028 ; 
        RECT 47.488 102.654 47.592 107.028 ; 
        RECT 47.056 102.654 47.16 107.028 ; 
        RECT 46.624 102.654 46.728 107.028 ; 
        RECT 46.192 102.654 46.296 107.028 ; 
        RECT 45.76 102.654 45.864 107.028 ; 
        RECT 45.328 102.654 45.432 107.028 ; 
        RECT 44.896 102.654 45 107.028 ; 
        RECT 44.464 102.654 44.568 107.028 ; 
        RECT 44.032 102.654 44.136 107.028 ; 
        RECT 43.6 102.654 43.704 107.028 ; 
        RECT 43.168 102.654 43.272 107.028 ; 
        RECT 42.736 102.654 42.84 107.028 ; 
        RECT 42.304 102.654 42.408 107.028 ; 
        RECT 41.872 102.654 41.976 107.028 ; 
        RECT 41.44 102.654 41.544 107.028 ; 
        RECT 41.008 102.654 41.112 107.028 ; 
        RECT 40.576 102.654 40.68 107.028 ; 
        RECT 40.144 102.654 40.248 107.028 ; 
        RECT 39.712 102.654 39.816 107.028 ; 
        RECT 39.28 102.654 39.384 107.028 ; 
        RECT 38.848 102.654 38.952 107.028 ; 
        RECT 38.416 102.654 38.52 107.028 ; 
        RECT 37.984 102.654 38.088 107.028 ; 
        RECT 37.552 102.654 37.656 107.028 ; 
        RECT 36.7 102.654 37.008 107.028 ; 
        RECT 29.128 102.654 29.436 107.028 ; 
        RECT 28.48 102.654 28.584 107.028 ; 
        RECT 28.048 102.654 28.152 107.028 ; 
        RECT 27.616 102.654 27.72 107.028 ; 
        RECT 27.184 102.654 27.288 107.028 ; 
        RECT 26.752 102.654 26.856 107.028 ; 
        RECT 26.32 102.654 26.424 107.028 ; 
        RECT 25.888 102.654 25.992 107.028 ; 
        RECT 25.456 102.654 25.56 107.028 ; 
        RECT 25.024 102.654 25.128 107.028 ; 
        RECT 24.592 102.654 24.696 107.028 ; 
        RECT 24.16 102.654 24.264 107.028 ; 
        RECT 23.728 102.654 23.832 107.028 ; 
        RECT 23.296 102.654 23.4 107.028 ; 
        RECT 22.864 102.654 22.968 107.028 ; 
        RECT 22.432 102.654 22.536 107.028 ; 
        RECT 22 102.654 22.104 107.028 ; 
        RECT 21.568 102.654 21.672 107.028 ; 
        RECT 21.136 102.654 21.24 107.028 ; 
        RECT 20.704 102.654 20.808 107.028 ; 
        RECT 20.272 102.654 20.376 107.028 ; 
        RECT 19.84 102.654 19.944 107.028 ; 
        RECT 19.408 102.654 19.512 107.028 ; 
        RECT 18.976 102.654 19.08 107.028 ; 
        RECT 18.544 102.654 18.648 107.028 ; 
        RECT 18.112 102.654 18.216 107.028 ; 
        RECT 17.68 102.654 17.784 107.028 ; 
        RECT 17.248 102.654 17.352 107.028 ; 
        RECT 16.816 102.654 16.92 107.028 ; 
        RECT 16.384 102.654 16.488 107.028 ; 
        RECT 15.952 102.654 16.056 107.028 ; 
        RECT 15.52 102.654 15.624 107.028 ; 
        RECT 15.088 102.654 15.192 107.028 ; 
        RECT 14.656 102.654 14.76 107.028 ; 
        RECT 14.224 102.654 14.328 107.028 ; 
        RECT 13.792 102.654 13.896 107.028 ; 
        RECT 13.36 102.654 13.464 107.028 ; 
        RECT 12.928 102.654 13.032 107.028 ; 
        RECT 12.496 102.654 12.6 107.028 ; 
        RECT 12.064 102.654 12.168 107.028 ; 
        RECT 11.632 102.654 11.736 107.028 ; 
        RECT 11.2 102.654 11.304 107.028 ; 
        RECT 10.768 102.654 10.872 107.028 ; 
        RECT 10.336 102.654 10.44 107.028 ; 
        RECT 9.904 102.654 10.008 107.028 ; 
        RECT 9.472 102.654 9.576 107.028 ; 
        RECT 9.04 102.654 9.144 107.028 ; 
        RECT 8.608 102.654 8.712 107.028 ; 
        RECT 8.176 102.654 8.28 107.028 ; 
        RECT 7.744 102.654 7.848 107.028 ; 
        RECT 7.312 102.654 7.416 107.028 ; 
        RECT 6.88 102.654 6.984 107.028 ; 
        RECT 6.448 102.654 6.552 107.028 ; 
        RECT 6.016 102.654 6.12 107.028 ; 
        RECT 5.584 102.654 5.688 107.028 ; 
        RECT 5.152 102.654 5.256 107.028 ; 
        RECT 4.72 102.654 4.824 107.028 ; 
        RECT 4.288 102.654 4.392 107.028 ; 
        RECT 3.856 102.654 3.96 107.028 ; 
        RECT 3.424 102.654 3.528 107.028 ; 
        RECT 2.992 102.654 3.096 107.028 ; 
        RECT 2.56 102.654 2.664 107.028 ; 
        RECT 2.128 102.654 2.232 107.028 ; 
        RECT 1.696 102.654 1.8 107.028 ; 
        RECT 1.264 102.654 1.368 107.028 ; 
        RECT 0.832 102.654 0.936 107.028 ; 
        RECT 0.02 102.654 0.36 107.028 ; 
        RECT 34.564 106.974 35.076 111.348 ; 
        RECT 34.508 109.636 35.076 110.926 ; 
        RECT 33.916 108.544 34.164 111.348 ; 
        RECT 33.86 109.782 34.164 110.396 ; 
        RECT 33.916 106.974 34.02 111.348 ; 
        RECT 33.916 107.458 34.076 108.416 ; 
        RECT 33.916 106.974 34.164 107.33 ; 
        RECT 32.728 108.776 33.552 111.348 ; 
        RECT 33.448 106.974 33.552 111.348 ; 
        RECT 32.728 109.884 33.608 110.916 ; 
        RECT 32.728 106.974 33.12 111.348 ; 
        RECT 31.06 106.974 31.392 111.348 ; 
        RECT 31.06 107.328 31.448 111.07 ; 
        RECT 65.776 106.974 66.116 111.348 ; 
        RECT 65.2 106.974 65.304 111.348 ; 
        RECT 64.768 106.974 64.872 111.348 ; 
        RECT 64.336 106.974 64.44 111.348 ; 
        RECT 63.904 106.974 64.008 111.348 ; 
        RECT 63.472 106.974 63.576 111.348 ; 
        RECT 63.04 106.974 63.144 111.348 ; 
        RECT 62.608 106.974 62.712 111.348 ; 
        RECT 62.176 106.974 62.28 111.348 ; 
        RECT 61.744 106.974 61.848 111.348 ; 
        RECT 61.312 106.974 61.416 111.348 ; 
        RECT 60.88 106.974 60.984 111.348 ; 
        RECT 60.448 106.974 60.552 111.348 ; 
        RECT 60.016 106.974 60.12 111.348 ; 
        RECT 59.584 106.974 59.688 111.348 ; 
        RECT 59.152 106.974 59.256 111.348 ; 
        RECT 58.72 106.974 58.824 111.348 ; 
        RECT 58.288 106.974 58.392 111.348 ; 
        RECT 57.856 106.974 57.96 111.348 ; 
        RECT 57.424 106.974 57.528 111.348 ; 
        RECT 56.992 106.974 57.096 111.348 ; 
        RECT 56.56 106.974 56.664 111.348 ; 
        RECT 56.128 106.974 56.232 111.348 ; 
        RECT 55.696 106.974 55.8 111.348 ; 
        RECT 55.264 106.974 55.368 111.348 ; 
        RECT 54.832 106.974 54.936 111.348 ; 
        RECT 54.4 106.974 54.504 111.348 ; 
        RECT 53.968 106.974 54.072 111.348 ; 
        RECT 53.536 106.974 53.64 111.348 ; 
        RECT 53.104 106.974 53.208 111.348 ; 
        RECT 52.672 106.974 52.776 111.348 ; 
        RECT 52.24 106.974 52.344 111.348 ; 
        RECT 51.808 106.974 51.912 111.348 ; 
        RECT 51.376 106.974 51.48 111.348 ; 
        RECT 50.944 106.974 51.048 111.348 ; 
        RECT 50.512 106.974 50.616 111.348 ; 
        RECT 50.08 106.974 50.184 111.348 ; 
        RECT 49.648 106.974 49.752 111.348 ; 
        RECT 49.216 106.974 49.32 111.348 ; 
        RECT 48.784 106.974 48.888 111.348 ; 
        RECT 48.352 106.974 48.456 111.348 ; 
        RECT 47.92 106.974 48.024 111.348 ; 
        RECT 47.488 106.974 47.592 111.348 ; 
        RECT 47.056 106.974 47.16 111.348 ; 
        RECT 46.624 106.974 46.728 111.348 ; 
        RECT 46.192 106.974 46.296 111.348 ; 
        RECT 45.76 106.974 45.864 111.348 ; 
        RECT 45.328 106.974 45.432 111.348 ; 
        RECT 44.896 106.974 45 111.348 ; 
        RECT 44.464 106.974 44.568 111.348 ; 
        RECT 44.032 106.974 44.136 111.348 ; 
        RECT 43.6 106.974 43.704 111.348 ; 
        RECT 43.168 106.974 43.272 111.348 ; 
        RECT 42.736 106.974 42.84 111.348 ; 
        RECT 42.304 106.974 42.408 111.348 ; 
        RECT 41.872 106.974 41.976 111.348 ; 
        RECT 41.44 106.974 41.544 111.348 ; 
        RECT 41.008 106.974 41.112 111.348 ; 
        RECT 40.576 106.974 40.68 111.348 ; 
        RECT 40.144 106.974 40.248 111.348 ; 
        RECT 39.712 106.974 39.816 111.348 ; 
        RECT 39.28 106.974 39.384 111.348 ; 
        RECT 38.848 106.974 38.952 111.348 ; 
        RECT 38.416 106.974 38.52 111.348 ; 
        RECT 37.984 106.974 38.088 111.348 ; 
        RECT 37.552 106.974 37.656 111.348 ; 
        RECT 36.7 106.974 37.008 111.348 ; 
        RECT 29.128 106.974 29.436 111.348 ; 
        RECT 28.48 106.974 28.584 111.348 ; 
        RECT 28.048 106.974 28.152 111.348 ; 
        RECT 27.616 106.974 27.72 111.348 ; 
        RECT 27.184 106.974 27.288 111.348 ; 
        RECT 26.752 106.974 26.856 111.348 ; 
        RECT 26.32 106.974 26.424 111.348 ; 
        RECT 25.888 106.974 25.992 111.348 ; 
        RECT 25.456 106.974 25.56 111.348 ; 
        RECT 25.024 106.974 25.128 111.348 ; 
        RECT 24.592 106.974 24.696 111.348 ; 
        RECT 24.16 106.974 24.264 111.348 ; 
        RECT 23.728 106.974 23.832 111.348 ; 
        RECT 23.296 106.974 23.4 111.348 ; 
        RECT 22.864 106.974 22.968 111.348 ; 
        RECT 22.432 106.974 22.536 111.348 ; 
        RECT 22 106.974 22.104 111.348 ; 
        RECT 21.568 106.974 21.672 111.348 ; 
        RECT 21.136 106.974 21.24 111.348 ; 
        RECT 20.704 106.974 20.808 111.348 ; 
        RECT 20.272 106.974 20.376 111.348 ; 
        RECT 19.84 106.974 19.944 111.348 ; 
        RECT 19.408 106.974 19.512 111.348 ; 
        RECT 18.976 106.974 19.08 111.348 ; 
        RECT 18.544 106.974 18.648 111.348 ; 
        RECT 18.112 106.974 18.216 111.348 ; 
        RECT 17.68 106.974 17.784 111.348 ; 
        RECT 17.248 106.974 17.352 111.348 ; 
        RECT 16.816 106.974 16.92 111.348 ; 
        RECT 16.384 106.974 16.488 111.348 ; 
        RECT 15.952 106.974 16.056 111.348 ; 
        RECT 15.52 106.974 15.624 111.348 ; 
        RECT 15.088 106.974 15.192 111.348 ; 
        RECT 14.656 106.974 14.76 111.348 ; 
        RECT 14.224 106.974 14.328 111.348 ; 
        RECT 13.792 106.974 13.896 111.348 ; 
        RECT 13.36 106.974 13.464 111.348 ; 
        RECT 12.928 106.974 13.032 111.348 ; 
        RECT 12.496 106.974 12.6 111.348 ; 
        RECT 12.064 106.974 12.168 111.348 ; 
        RECT 11.632 106.974 11.736 111.348 ; 
        RECT 11.2 106.974 11.304 111.348 ; 
        RECT 10.768 106.974 10.872 111.348 ; 
        RECT 10.336 106.974 10.44 111.348 ; 
        RECT 9.904 106.974 10.008 111.348 ; 
        RECT 9.472 106.974 9.576 111.348 ; 
        RECT 9.04 106.974 9.144 111.348 ; 
        RECT 8.608 106.974 8.712 111.348 ; 
        RECT 8.176 106.974 8.28 111.348 ; 
        RECT 7.744 106.974 7.848 111.348 ; 
        RECT 7.312 106.974 7.416 111.348 ; 
        RECT 6.88 106.974 6.984 111.348 ; 
        RECT 6.448 106.974 6.552 111.348 ; 
        RECT 6.016 106.974 6.12 111.348 ; 
        RECT 5.584 106.974 5.688 111.348 ; 
        RECT 5.152 106.974 5.256 111.348 ; 
        RECT 4.72 106.974 4.824 111.348 ; 
        RECT 4.288 106.974 4.392 111.348 ; 
        RECT 3.856 106.974 3.96 111.348 ; 
        RECT 3.424 106.974 3.528 111.348 ; 
        RECT 2.992 106.974 3.096 111.348 ; 
        RECT 2.56 106.974 2.664 111.348 ; 
        RECT 2.128 106.974 2.232 111.348 ; 
        RECT 1.696 106.974 1.8 111.348 ; 
        RECT 1.264 106.974 1.368 111.348 ; 
        RECT 0.832 106.974 0.936 111.348 ; 
        RECT 0.02 106.974 0.36 111.348 ; 
        RECT 34.564 111.294 35.076 115.668 ; 
        RECT 34.508 113.956 35.076 115.246 ; 
        RECT 33.916 112.864 34.164 115.668 ; 
        RECT 33.86 114.102 34.164 114.716 ; 
        RECT 33.916 111.294 34.02 115.668 ; 
        RECT 33.916 111.778 34.076 112.736 ; 
        RECT 33.916 111.294 34.164 111.65 ; 
        RECT 32.728 113.096 33.552 115.668 ; 
        RECT 33.448 111.294 33.552 115.668 ; 
        RECT 32.728 114.204 33.608 115.236 ; 
        RECT 32.728 111.294 33.12 115.668 ; 
        RECT 31.06 111.294 31.392 115.668 ; 
        RECT 31.06 111.648 31.448 115.39 ; 
        RECT 65.776 111.294 66.116 115.668 ; 
        RECT 65.2 111.294 65.304 115.668 ; 
        RECT 64.768 111.294 64.872 115.668 ; 
        RECT 64.336 111.294 64.44 115.668 ; 
        RECT 63.904 111.294 64.008 115.668 ; 
        RECT 63.472 111.294 63.576 115.668 ; 
        RECT 63.04 111.294 63.144 115.668 ; 
        RECT 62.608 111.294 62.712 115.668 ; 
        RECT 62.176 111.294 62.28 115.668 ; 
        RECT 61.744 111.294 61.848 115.668 ; 
        RECT 61.312 111.294 61.416 115.668 ; 
        RECT 60.88 111.294 60.984 115.668 ; 
        RECT 60.448 111.294 60.552 115.668 ; 
        RECT 60.016 111.294 60.12 115.668 ; 
        RECT 59.584 111.294 59.688 115.668 ; 
        RECT 59.152 111.294 59.256 115.668 ; 
        RECT 58.72 111.294 58.824 115.668 ; 
        RECT 58.288 111.294 58.392 115.668 ; 
        RECT 57.856 111.294 57.96 115.668 ; 
        RECT 57.424 111.294 57.528 115.668 ; 
        RECT 56.992 111.294 57.096 115.668 ; 
        RECT 56.56 111.294 56.664 115.668 ; 
        RECT 56.128 111.294 56.232 115.668 ; 
        RECT 55.696 111.294 55.8 115.668 ; 
        RECT 55.264 111.294 55.368 115.668 ; 
        RECT 54.832 111.294 54.936 115.668 ; 
        RECT 54.4 111.294 54.504 115.668 ; 
        RECT 53.968 111.294 54.072 115.668 ; 
        RECT 53.536 111.294 53.64 115.668 ; 
        RECT 53.104 111.294 53.208 115.668 ; 
        RECT 52.672 111.294 52.776 115.668 ; 
        RECT 52.24 111.294 52.344 115.668 ; 
        RECT 51.808 111.294 51.912 115.668 ; 
        RECT 51.376 111.294 51.48 115.668 ; 
        RECT 50.944 111.294 51.048 115.668 ; 
        RECT 50.512 111.294 50.616 115.668 ; 
        RECT 50.08 111.294 50.184 115.668 ; 
        RECT 49.648 111.294 49.752 115.668 ; 
        RECT 49.216 111.294 49.32 115.668 ; 
        RECT 48.784 111.294 48.888 115.668 ; 
        RECT 48.352 111.294 48.456 115.668 ; 
        RECT 47.92 111.294 48.024 115.668 ; 
        RECT 47.488 111.294 47.592 115.668 ; 
        RECT 47.056 111.294 47.16 115.668 ; 
        RECT 46.624 111.294 46.728 115.668 ; 
        RECT 46.192 111.294 46.296 115.668 ; 
        RECT 45.76 111.294 45.864 115.668 ; 
        RECT 45.328 111.294 45.432 115.668 ; 
        RECT 44.896 111.294 45 115.668 ; 
        RECT 44.464 111.294 44.568 115.668 ; 
        RECT 44.032 111.294 44.136 115.668 ; 
        RECT 43.6 111.294 43.704 115.668 ; 
        RECT 43.168 111.294 43.272 115.668 ; 
        RECT 42.736 111.294 42.84 115.668 ; 
        RECT 42.304 111.294 42.408 115.668 ; 
        RECT 41.872 111.294 41.976 115.668 ; 
        RECT 41.44 111.294 41.544 115.668 ; 
        RECT 41.008 111.294 41.112 115.668 ; 
        RECT 40.576 111.294 40.68 115.668 ; 
        RECT 40.144 111.294 40.248 115.668 ; 
        RECT 39.712 111.294 39.816 115.668 ; 
        RECT 39.28 111.294 39.384 115.668 ; 
        RECT 38.848 111.294 38.952 115.668 ; 
        RECT 38.416 111.294 38.52 115.668 ; 
        RECT 37.984 111.294 38.088 115.668 ; 
        RECT 37.552 111.294 37.656 115.668 ; 
        RECT 36.7 111.294 37.008 115.668 ; 
        RECT 29.128 111.294 29.436 115.668 ; 
        RECT 28.48 111.294 28.584 115.668 ; 
        RECT 28.048 111.294 28.152 115.668 ; 
        RECT 27.616 111.294 27.72 115.668 ; 
        RECT 27.184 111.294 27.288 115.668 ; 
        RECT 26.752 111.294 26.856 115.668 ; 
        RECT 26.32 111.294 26.424 115.668 ; 
        RECT 25.888 111.294 25.992 115.668 ; 
        RECT 25.456 111.294 25.56 115.668 ; 
        RECT 25.024 111.294 25.128 115.668 ; 
        RECT 24.592 111.294 24.696 115.668 ; 
        RECT 24.16 111.294 24.264 115.668 ; 
        RECT 23.728 111.294 23.832 115.668 ; 
        RECT 23.296 111.294 23.4 115.668 ; 
        RECT 22.864 111.294 22.968 115.668 ; 
        RECT 22.432 111.294 22.536 115.668 ; 
        RECT 22 111.294 22.104 115.668 ; 
        RECT 21.568 111.294 21.672 115.668 ; 
        RECT 21.136 111.294 21.24 115.668 ; 
        RECT 20.704 111.294 20.808 115.668 ; 
        RECT 20.272 111.294 20.376 115.668 ; 
        RECT 19.84 111.294 19.944 115.668 ; 
        RECT 19.408 111.294 19.512 115.668 ; 
        RECT 18.976 111.294 19.08 115.668 ; 
        RECT 18.544 111.294 18.648 115.668 ; 
        RECT 18.112 111.294 18.216 115.668 ; 
        RECT 17.68 111.294 17.784 115.668 ; 
        RECT 17.248 111.294 17.352 115.668 ; 
        RECT 16.816 111.294 16.92 115.668 ; 
        RECT 16.384 111.294 16.488 115.668 ; 
        RECT 15.952 111.294 16.056 115.668 ; 
        RECT 15.52 111.294 15.624 115.668 ; 
        RECT 15.088 111.294 15.192 115.668 ; 
        RECT 14.656 111.294 14.76 115.668 ; 
        RECT 14.224 111.294 14.328 115.668 ; 
        RECT 13.792 111.294 13.896 115.668 ; 
        RECT 13.36 111.294 13.464 115.668 ; 
        RECT 12.928 111.294 13.032 115.668 ; 
        RECT 12.496 111.294 12.6 115.668 ; 
        RECT 12.064 111.294 12.168 115.668 ; 
        RECT 11.632 111.294 11.736 115.668 ; 
        RECT 11.2 111.294 11.304 115.668 ; 
        RECT 10.768 111.294 10.872 115.668 ; 
        RECT 10.336 111.294 10.44 115.668 ; 
        RECT 9.904 111.294 10.008 115.668 ; 
        RECT 9.472 111.294 9.576 115.668 ; 
        RECT 9.04 111.294 9.144 115.668 ; 
        RECT 8.608 111.294 8.712 115.668 ; 
        RECT 8.176 111.294 8.28 115.668 ; 
        RECT 7.744 111.294 7.848 115.668 ; 
        RECT 7.312 111.294 7.416 115.668 ; 
        RECT 6.88 111.294 6.984 115.668 ; 
        RECT 6.448 111.294 6.552 115.668 ; 
        RECT 6.016 111.294 6.12 115.668 ; 
        RECT 5.584 111.294 5.688 115.668 ; 
        RECT 5.152 111.294 5.256 115.668 ; 
        RECT 4.72 111.294 4.824 115.668 ; 
        RECT 4.288 111.294 4.392 115.668 ; 
        RECT 3.856 111.294 3.96 115.668 ; 
        RECT 3.424 111.294 3.528 115.668 ; 
        RECT 2.992 111.294 3.096 115.668 ; 
        RECT 2.56 111.294 2.664 115.668 ; 
        RECT 2.128 111.294 2.232 115.668 ; 
        RECT 1.696 111.294 1.8 115.668 ; 
        RECT 1.264 111.294 1.368 115.668 ; 
        RECT 0.832 111.294 0.936 115.668 ; 
        RECT 0.02 111.294 0.36 115.668 ; 
        RECT 34.564 115.614 35.076 119.988 ; 
        RECT 34.508 118.276 35.076 119.566 ; 
        RECT 33.916 117.184 34.164 119.988 ; 
        RECT 33.86 118.422 34.164 119.036 ; 
        RECT 33.916 115.614 34.02 119.988 ; 
        RECT 33.916 116.098 34.076 117.056 ; 
        RECT 33.916 115.614 34.164 115.97 ; 
        RECT 32.728 117.416 33.552 119.988 ; 
        RECT 33.448 115.614 33.552 119.988 ; 
        RECT 32.728 118.524 33.608 119.556 ; 
        RECT 32.728 115.614 33.12 119.988 ; 
        RECT 31.06 115.614 31.392 119.988 ; 
        RECT 31.06 115.968 31.448 119.71 ; 
        RECT 65.776 115.614 66.116 119.988 ; 
        RECT 65.2 115.614 65.304 119.988 ; 
        RECT 64.768 115.614 64.872 119.988 ; 
        RECT 64.336 115.614 64.44 119.988 ; 
        RECT 63.904 115.614 64.008 119.988 ; 
        RECT 63.472 115.614 63.576 119.988 ; 
        RECT 63.04 115.614 63.144 119.988 ; 
        RECT 62.608 115.614 62.712 119.988 ; 
        RECT 62.176 115.614 62.28 119.988 ; 
        RECT 61.744 115.614 61.848 119.988 ; 
        RECT 61.312 115.614 61.416 119.988 ; 
        RECT 60.88 115.614 60.984 119.988 ; 
        RECT 60.448 115.614 60.552 119.988 ; 
        RECT 60.016 115.614 60.12 119.988 ; 
        RECT 59.584 115.614 59.688 119.988 ; 
        RECT 59.152 115.614 59.256 119.988 ; 
        RECT 58.72 115.614 58.824 119.988 ; 
        RECT 58.288 115.614 58.392 119.988 ; 
        RECT 57.856 115.614 57.96 119.988 ; 
        RECT 57.424 115.614 57.528 119.988 ; 
        RECT 56.992 115.614 57.096 119.988 ; 
        RECT 56.56 115.614 56.664 119.988 ; 
        RECT 56.128 115.614 56.232 119.988 ; 
        RECT 55.696 115.614 55.8 119.988 ; 
        RECT 55.264 115.614 55.368 119.988 ; 
        RECT 54.832 115.614 54.936 119.988 ; 
        RECT 54.4 115.614 54.504 119.988 ; 
        RECT 53.968 115.614 54.072 119.988 ; 
        RECT 53.536 115.614 53.64 119.988 ; 
        RECT 53.104 115.614 53.208 119.988 ; 
        RECT 52.672 115.614 52.776 119.988 ; 
        RECT 52.24 115.614 52.344 119.988 ; 
        RECT 51.808 115.614 51.912 119.988 ; 
        RECT 51.376 115.614 51.48 119.988 ; 
        RECT 50.944 115.614 51.048 119.988 ; 
        RECT 50.512 115.614 50.616 119.988 ; 
        RECT 50.08 115.614 50.184 119.988 ; 
        RECT 49.648 115.614 49.752 119.988 ; 
        RECT 49.216 115.614 49.32 119.988 ; 
        RECT 48.784 115.614 48.888 119.988 ; 
        RECT 48.352 115.614 48.456 119.988 ; 
        RECT 47.92 115.614 48.024 119.988 ; 
        RECT 47.488 115.614 47.592 119.988 ; 
        RECT 47.056 115.614 47.16 119.988 ; 
        RECT 46.624 115.614 46.728 119.988 ; 
        RECT 46.192 115.614 46.296 119.988 ; 
        RECT 45.76 115.614 45.864 119.988 ; 
        RECT 45.328 115.614 45.432 119.988 ; 
        RECT 44.896 115.614 45 119.988 ; 
        RECT 44.464 115.614 44.568 119.988 ; 
        RECT 44.032 115.614 44.136 119.988 ; 
        RECT 43.6 115.614 43.704 119.988 ; 
        RECT 43.168 115.614 43.272 119.988 ; 
        RECT 42.736 115.614 42.84 119.988 ; 
        RECT 42.304 115.614 42.408 119.988 ; 
        RECT 41.872 115.614 41.976 119.988 ; 
        RECT 41.44 115.614 41.544 119.988 ; 
        RECT 41.008 115.614 41.112 119.988 ; 
        RECT 40.576 115.614 40.68 119.988 ; 
        RECT 40.144 115.614 40.248 119.988 ; 
        RECT 39.712 115.614 39.816 119.988 ; 
        RECT 39.28 115.614 39.384 119.988 ; 
        RECT 38.848 115.614 38.952 119.988 ; 
        RECT 38.416 115.614 38.52 119.988 ; 
        RECT 37.984 115.614 38.088 119.988 ; 
        RECT 37.552 115.614 37.656 119.988 ; 
        RECT 36.7 115.614 37.008 119.988 ; 
        RECT 29.128 115.614 29.436 119.988 ; 
        RECT 28.48 115.614 28.584 119.988 ; 
        RECT 28.048 115.614 28.152 119.988 ; 
        RECT 27.616 115.614 27.72 119.988 ; 
        RECT 27.184 115.614 27.288 119.988 ; 
        RECT 26.752 115.614 26.856 119.988 ; 
        RECT 26.32 115.614 26.424 119.988 ; 
        RECT 25.888 115.614 25.992 119.988 ; 
        RECT 25.456 115.614 25.56 119.988 ; 
        RECT 25.024 115.614 25.128 119.988 ; 
        RECT 24.592 115.614 24.696 119.988 ; 
        RECT 24.16 115.614 24.264 119.988 ; 
        RECT 23.728 115.614 23.832 119.988 ; 
        RECT 23.296 115.614 23.4 119.988 ; 
        RECT 22.864 115.614 22.968 119.988 ; 
        RECT 22.432 115.614 22.536 119.988 ; 
        RECT 22 115.614 22.104 119.988 ; 
        RECT 21.568 115.614 21.672 119.988 ; 
        RECT 21.136 115.614 21.24 119.988 ; 
        RECT 20.704 115.614 20.808 119.988 ; 
        RECT 20.272 115.614 20.376 119.988 ; 
        RECT 19.84 115.614 19.944 119.988 ; 
        RECT 19.408 115.614 19.512 119.988 ; 
        RECT 18.976 115.614 19.08 119.988 ; 
        RECT 18.544 115.614 18.648 119.988 ; 
        RECT 18.112 115.614 18.216 119.988 ; 
        RECT 17.68 115.614 17.784 119.988 ; 
        RECT 17.248 115.614 17.352 119.988 ; 
        RECT 16.816 115.614 16.92 119.988 ; 
        RECT 16.384 115.614 16.488 119.988 ; 
        RECT 15.952 115.614 16.056 119.988 ; 
        RECT 15.52 115.614 15.624 119.988 ; 
        RECT 15.088 115.614 15.192 119.988 ; 
        RECT 14.656 115.614 14.76 119.988 ; 
        RECT 14.224 115.614 14.328 119.988 ; 
        RECT 13.792 115.614 13.896 119.988 ; 
        RECT 13.36 115.614 13.464 119.988 ; 
        RECT 12.928 115.614 13.032 119.988 ; 
        RECT 12.496 115.614 12.6 119.988 ; 
        RECT 12.064 115.614 12.168 119.988 ; 
        RECT 11.632 115.614 11.736 119.988 ; 
        RECT 11.2 115.614 11.304 119.988 ; 
        RECT 10.768 115.614 10.872 119.988 ; 
        RECT 10.336 115.614 10.44 119.988 ; 
        RECT 9.904 115.614 10.008 119.988 ; 
        RECT 9.472 115.614 9.576 119.988 ; 
        RECT 9.04 115.614 9.144 119.988 ; 
        RECT 8.608 115.614 8.712 119.988 ; 
        RECT 8.176 115.614 8.28 119.988 ; 
        RECT 7.744 115.614 7.848 119.988 ; 
        RECT 7.312 115.614 7.416 119.988 ; 
        RECT 6.88 115.614 6.984 119.988 ; 
        RECT 6.448 115.614 6.552 119.988 ; 
        RECT 6.016 115.614 6.12 119.988 ; 
        RECT 5.584 115.614 5.688 119.988 ; 
        RECT 5.152 115.614 5.256 119.988 ; 
        RECT 4.72 115.614 4.824 119.988 ; 
        RECT 4.288 115.614 4.392 119.988 ; 
        RECT 3.856 115.614 3.96 119.988 ; 
        RECT 3.424 115.614 3.528 119.988 ; 
        RECT 2.992 115.614 3.096 119.988 ; 
        RECT 2.56 115.614 2.664 119.988 ; 
        RECT 2.128 115.614 2.232 119.988 ; 
        RECT 1.696 115.614 1.8 119.988 ; 
        RECT 1.264 115.614 1.368 119.988 ; 
        RECT 0.832 115.614 0.936 119.988 ; 
        RECT 0.02 115.614 0.36 119.988 ; 
  LAYER V3 SPACING 0.072 ; 
      RECT 0.02 4.88 66.116 5.4 ; 
      RECT 65.648 1.026 66.116 5.4 ; 
      RECT 37.208 4.496 65.576 5.4 ; 
      RECT 31.88 4.496 37.136 5.4 ; 
      RECT 29 1.026 31.52 5.4 ; 
      RECT 0.56 4.496 28.928 5.4 ; 
      RECT 0.02 1.026 0.488 5.4 ; 
      RECT 65.504 1.026 66.116 4.688 ; 
      RECT 37.424 1.026 65.432 5.4 ; 
      RECT 34.436 1.026 37.352 4.688 ; 
      RECT 33.788 1.808 34.292 5.4 ; 
      RECT 28.784 1.424 33.68 4.688 ; 
      RECT 0.704 1.026 28.712 5.4 ; 
      RECT 0.02 1.026 0.632 4.688 ; 
      RECT 34.22 1.026 66.116 4.304 ; 
      RECT 0.02 1.424 34.148 4.304 ; 
      RECT 33.32 1.026 66.116 1.712 ; 
      RECT 0.02 1.026 33.248 4.304 ; 
      RECT 0.02 1.026 66.116 1.328 ; 
      RECT 0.02 9.2 66.116 9.72 ; 
      RECT 65.648 5.346 66.116 9.72 ; 
      RECT 37.208 8.816 65.576 9.72 ; 
      RECT 31.88 8.816 37.136 9.72 ; 
      RECT 29 5.346 31.52 9.72 ; 
      RECT 0.56 8.816 28.928 9.72 ; 
      RECT 0.02 5.346 0.488 9.72 ; 
      RECT 65.504 5.346 66.116 9.008 ; 
      RECT 37.424 5.346 65.432 9.72 ; 
      RECT 34.436 5.346 37.352 9.008 ; 
      RECT 33.788 6.128 34.292 9.72 ; 
      RECT 28.784 5.744 33.68 9.008 ; 
      RECT 0.704 5.346 28.712 9.72 ; 
      RECT 0.02 5.346 0.632 9.008 ; 
      RECT 34.22 5.346 66.116 8.624 ; 
      RECT 0.02 5.744 34.148 8.624 ; 
      RECT 33.32 5.346 66.116 6.032 ; 
      RECT 0.02 5.346 33.248 8.624 ; 
      RECT 0.02 5.346 66.116 5.648 ; 
      RECT 0.02 13.52 66.116 14.04 ; 
      RECT 65.648 9.666 66.116 14.04 ; 
      RECT 37.208 13.136 65.576 14.04 ; 
      RECT 31.88 13.136 37.136 14.04 ; 
      RECT 29 9.666 31.52 14.04 ; 
      RECT 0.56 13.136 28.928 14.04 ; 
      RECT 0.02 9.666 0.488 14.04 ; 
      RECT 65.504 9.666 66.116 13.328 ; 
      RECT 37.424 9.666 65.432 14.04 ; 
      RECT 34.436 9.666 37.352 13.328 ; 
      RECT 33.788 10.448 34.292 14.04 ; 
      RECT 28.784 10.064 33.68 13.328 ; 
      RECT 0.704 9.666 28.712 14.04 ; 
      RECT 0.02 9.666 0.632 13.328 ; 
      RECT 34.22 9.666 66.116 12.944 ; 
      RECT 0.02 10.064 34.148 12.944 ; 
      RECT 33.32 9.666 66.116 10.352 ; 
      RECT 0.02 9.666 33.248 12.944 ; 
      RECT 0.02 9.666 66.116 9.968 ; 
      RECT 0.02 17.84 66.116 18.36 ; 
      RECT 65.648 13.986 66.116 18.36 ; 
      RECT 37.208 17.456 65.576 18.36 ; 
      RECT 31.88 17.456 37.136 18.36 ; 
      RECT 29 13.986 31.52 18.36 ; 
      RECT 0.56 17.456 28.928 18.36 ; 
      RECT 0.02 13.986 0.488 18.36 ; 
      RECT 65.504 13.986 66.116 17.648 ; 
      RECT 37.424 13.986 65.432 18.36 ; 
      RECT 34.436 13.986 37.352 17.648 ; 
      RECT 33.788 14.768 34.292 18.36 ; 
      RECT 28.784 14.384 33.68 17.648 ; 
      RECT 0.704 13.986 28.712 18.36 ; 
      RECT 0.02 13.986 0.632 17.648 ; 
      RECT 34.22 13.986 66.116 17.264 ; 
      RECT 0.02 14.384 34.148 17.264 ; 
      RECT 33.32 13.986 66.116 14.672 ; 
      RECT 0.02 13.986 33.248 17.264 ; 
      RECT 0.02 13.986 66.116 14.288 ; 
      RECT 0.02 22.16 66.116 22.68 ; 
      RECT 65.648 18.306 66.116 22.68 ; 
      RECT 37.208 21.776 65.576 22.68 ; 
      RECT 31.88 21.776 37.136 22.68 ; 
      RECT 29 18.306 31.52 22.68 ; 
      RECT 0.56 21.776 28.928 22.68 ; 
      RECT 0.02 18.306 0.488 22.68 ; 
      RECT 65.504 18.306 66.116 21.968 ; 
      RECT 37.424 18.306 65.432 22.68 ; 
      RECT 34.436 18.306 37.352 21.968 ; 
      RECT 33.788 19.088 34.292 22.68 ; 
      RECT 28.784 18.704 33.68 21.968 ; 
      RECT 0.704 18.306 28.712 22.68 ; 
      RECT 0.02 18.306 0.632 21.968 ; 
      RECT 34.22 18.306 66.116 21.584 ; 
      RECT 0.02 18.704 34.148 21.584 ; 
      RECT 33.32 18.306 66.116 18.992 ; 
      RECT 0.02 18.306 33.248 21.584 ; 
      RECT 0.02 18.306 66.116 18.608 ; 
      RECT 0.02 26.48 66.116 27 ; 
      RECT 65.648 22.626 66.116 27 ; 
      RECT 37.208 26.096 65.576 27 ; 
      RECT 31.88 26.096 37.136 27 ; 
      RECT 29 22.626 31.52 27 ; 
      RECT 0.56 26.096 28.928 27 ; 
      RECT 0.02 22.626 0.488 27 ; 
      RECT 65.504 22.626 66.116 26.288 ; 
      RECT 37.424 22.626 65.432 27 ; 
      RECT 34.436 22.626 37.352 26.288 ; 
      RECT 33.788 23.408 34.292 27 ; 
      RECT 28.784 23.024 33.68 26.288 ; 
      RECT 0.704 22.626 28.712 27 ; 
      RECT 0.02 22.626 0.632 26.288 ; 
      RECT 34.22 22.626 66.116 25.904 ; 
      RECT 0.02 23.024 34.148 25.904 ; 
      RECT 33.32 22.626 66.116 23.312 ; 
      RECT 0.02 22.626 33.248 25.904 ; 
      RECT 0.02 22.626 66.116 22.928 ; 
      RECT 0.02 30.8 66.116 31.32 ; 
      RECT 65.648 26.946 66.116 31.32 ; 
      RECT 37.208 30.416 65.576 31.32 ; 
      RECT 31.88 30.416 37.136 31.32 ; 
      RECT 29 26.946 31.52 31.32 ; 
      RECT 0.56 30.416 28.928 31.32 ; 
      RECT 0.02 26.946 0.488 31.32 ; 
      RECT 65.504 26.946 66.116 30.608 ; 
      RECT 37.424 26.946 65.432 31.32 ; 
      RECT 34.436 26.946 37.352 30.608 ; 
      RECT 33.788 27.728 34.292 31.32 ; 
      RECT 28.784 27.344 33.68 30.608 ; 
      RECT 0.704 26.946 28.712 31.32 ; 
      RECT 0.02 26.946 0.632 30.608 ; 
      RECT 34.22 26.946 66.116 30.224 ; 
      RECT 0.02 27.344 34.148 30.224 ; 
      RECT 33.32 26.946 66.116 27.632 ; 
      RECT 0.02 26.946 33.248 30.224 ; 
      RECT 0.02 26.946 66.116 27.248 ; 
      RECT 0.02 35.12 66.116 35.64 ; 
      RECT 65.648 31.266 66.116 35.64 ; 
      RECT 37.208 34.736 65.576 35.64 ; 
      RECT 31.88 34.736 37.136 35.64 ; 
      RECT 29 31.266 31.52 35.64 ; 
      RECT 0.56 34.736 28.928 35.64 ; 
      RECT 0.02 31.266 0.488 35.64 ; 
      RECT 65.504 31.266 66.116 34.928 ; 
      RECT 37.424 31.266 65.432 35.64 ; 
      RECT 34.436 31.266 37.352 34.928 ; 
      RECT 33.788 32.048 34.292 35.64 ; 
      RECT 28.784 31.664 33.68 34.928 ; 
      RECT 0.704 31.266 28.712 35.64 ; 
      RECT 0.02 31.266 0.632 34.928 ; 
      RECT 34.22 31.266 66.116 34.544 ; 
      RECT 0.02 31.664 34.148 34.544 ; 
      RECT 33.32 31.266 66.116 31.952 ; 
      RECT 0.02 31.266 33.248 34.544 ; 
      RECT 0.02 31.266 66.116 31.568 ; 
      RECT 0.02 39.44 66.116 39.96 ; 
      RECT 65.648 35.586 66.116 39.96 ; 
      RECT 37.208 39.056 65.576 39.96 ; 
      RECT 31.88 39.056 37.136 39.96 ; 
      RECT 29 35.586 31.52 39.96 ; 
      RECT 0.56 39.056 28.928 39.96 ; 
      RECT 0.02 35.586 0.488 39.96 ; 
      RECT 65.504 35.586 66.116 39.248 ; 
      RECT 37.424 35.586 65.432 39.96 ; 
      RECT 34.436 35.586 37.352 39.248 ; 
      RECT 33.788 36.368 34.292 39.96 ; 
      RECT 28.784 35.984 33.68 39.248 ; 
      RECT 0.704 35.586 28.712 39.96 ; 
      RECT 0.02 35.586 0.632 39.248 ; 
      RECT 34.22 35.586 66.116 38.864 ; 
      RECT 0.02 35.984 34.148 38.864 ; 
      RECT 33.32 35.586 66.116 36.272 ; 
      RECT 0.02 35.586 33.248 38.864 ; 
      RECT 0.02 35.586 66.116 35.888 ; 
      RECT 0.02 43.76 66.116 44.28 ; 
      RECT 65.648 39.906 66.116 44.28 ; 
      RECT 37.208 43.376 65.576 44.28 ; 
      RECT 31.88 43.376 37.136 44.28 ; 
      RECT 29 39.906 31.52 44.28 ; 
      RECT 0.56 43.376 28.928 44.28 ; 
      RECT 0.02 39.906 0.488 44.28 ; 
      RECT 65.504 39.906 66.116 43.568 ; 
      RECT 37.424 39.906 65.432 44.28 ; 
      RECT 34.436 39.906 37.352 43.568 ; 
      RECT 33.788 40.688 34.292 44.28 ; 
      RECT 28.784 40.304 33.68 43.568 ; 
      RECT 0.704 39.906 28.712 44.28 ; 
      RECT 0.02 39.906 0.632 43.568 ; 
      RECT 34.22 39.906 66.116 43.184 ; 
      RECT 0.02 40.304 34.148 43.184 ; 
      RECT 33.32 39.906 66.116 40.592 ; 
      RECT 0.02 39.906 33.248 43.184 ; 
      RECT 0.02 39.906 66.116 40.208 ; 
      RECT 0 73.428 66.096 78.762 ; 
      RECT 43.236 44.148 66.096 78.762 ; 
      RECT 34.436 59.604 66.096 78.762 ; 
      RECT 38.052 49.236 66.096 78.762 ; 
      RECT 34.228 44.148 34.364 78.762 ; 
      RECT 34.02 44.148 34.156 78.762 ; 
      RECT 33.812 44.148 33.948 78.762 ; 
      RECT 33.604 44.148 33.74 78.762 ; 
      RECT 0 71.7 33.532 78.762 ; 
      RECT 32.564 60.756 66.096 72.564 ; 
      RECT 32.356 44.148 32.492 78.762 ; 
      RECT 32.148 44.148 32.284 78.762 ; 
      RECT 31.94 44.148 32.076 78.762 ; 
      RECT 31.732 44.148 31.868 78.762 ; 
      RECT 0 50.388 31.66 78.762 ; 
      RECT 0 59.028 33.532 70.836 ; 
      RECT 32.564 48.084 37.116 59.892 ; 
      RECT 37.26 50.004 66.096 78.762 ; 
      RECT 0 59.028 37.188 59.892 ; 
      RECT 32.564 50.004 66.096 59.508 ; 
      RECT 29.844 46.356 32.94 58.164 ; 
      RECT 28.98 46.932 31.66 78.762 ; 
      RECT 0 49.236 28.908 78.762 ; 
      RECT 27.252 44.148 29.052 50.292 ; 
      RECT 0 49.62 37.98 50.292 ; 
      RECT 37.188 49.236 66.096 49.908 ; 
      RECT 42.372 44.148 43.164 78.762 ; 
      RECT 27.252 48.468 42.3 49.524 ; 
      RECT 23.796 46.932 27.18 78.762 ; 
      RECT 0 44.148 23.724 78.762 ; 
      RECT 41.508 44.148 66.096 49.14 ; 
      RECT 40.644 46.932 66.096 49.14 ; 
      RECT 0 48.086 40.572 49.14 ; 
      RECT 39.78 44.148 41.436 48.372 ; 
      RECT 37.404 46.932 66.096 48.372 ; 
      RECT 34.436 46.932 37.332 49.524 ; 
      RECT 32.564 46.74 33.532 78.762 ; 
      RECT 33.012 44.148 34.524 47.22 ; 
      RECT 34.596 46.74 39.708 47.222 ; 
      RECT 26.388 46.74 29.772 49.14 ; 
      RECT 24.66 46.74 26.316 78.762 ; 
      RECT 0 44.148 24.588 49.14 ; 
      RECT 38.916 44.148 66.096 46.836 ; 
      RECT 33.012 44.468 38.844 46.836 ; 
      RECT 29.124 46.356 32.94 46.836 ; 
      RECT 25.524 44.148 29.052 46.836 ; 
      RECT 0 44.148 25.452 46.836 ; 
      RECT 37.188 44.148 66.096 46.644 ; 
      RECT 32.564 44.468 66.096 46.644 ; 
      RECT 0 44.148 31.66 46.644 ; 
      RECT 0 44.148 37.116 45.492 ; 
      RECT 0 44.148 66.096 44.372 ; 
        RECT 0.02 80.588 66.116 81.108 ; 
        RECT 65.648 76.734 66.116 81.108 ; 
        RECT 37.208 80.204 65.576 81.108 ; 
        RECT 31.88 80.204 37.136 81.108 ; 
        RECT 29 76.734 31.52 81.108 ; 
        RECT 0.56 80.204 28.928 81.108 ; 
        RECT 0.02 76.734 0.488 81.108 ; 
        RECT 65.504 76.734 66.116 80.396 ; 
        RECT 37.424 76.734 65.432 81.108 ; 
        RECT 34.436 76.734 37.352 80.396 ; 
        RECT 33.788 77.516 34.292 81.108 ; 
        RECT 28.784 77.132 33.68 80.396 ; 
        RECT 0.704 76.734 28.712 81.108 ; 
        RECT 0.02 76.734 0.632 80.396 ; 
        RECT 34.22 76.734 66.116 80.012 ; 
        RECT 0.02 77.132 34.148 80.012 ; 
        RECT 33.32 76.734 66.116 77.42 ; 
        RECT 0.02 76.734 33.248 80.012 ; 
        RECT 0.02 76.734 66.116 77.036 ; 
        RECT 0.02 84.908 66.116 85.428 ; 
        RECT 65.648 81.054 66.116 85.428 ; 
        RECT 37.208 84.524 65.576 85.428 ; 
        RECT 31.88 84.524 37.136 85.428 ; 
        RECT 29 81.054 31.52 85.428 ; 
        RECT 0.56 84.524 28.928 85.428 ; 
        RECT 0.02 81.054 0.488 85.428 ; 
        RECT 65.504 81.054 66.116 84.716 ; 
        RECT 37.424 81.054 65.432 85.428 ; 
        RECT 34.436 81.054 37.352 84.716 ; 
        RECT 33.788 81.836 34.292 85.428 ; 
        RECT 28.784 81.452 33.68 84.716 ; 
        RECT 0.704 81.054 28.712 85.428 ; 
        RECT 0.02 81.054 0.632 84.716 ; 
        RECT 34.22 81.054 66.116 84.332 ; 
        RECT 0.02 81.452 34.148 84.332 ; 
        RECT 33.32 81.054 66.116 81.74 ; 
        RECT 0.02 81.054 33.248 84.332 ; 
        RECT 0.02 81.054 66.116 81.356 ; 
        RECT 0.02 89.228 66.116 89.748 ; 
        RECT 65.648 85.374 66.116 89.748 ; 
        RECT 37.208 88.844 65.576 89.748 ; 
        RECT 31.88 88.844 37.136 89.748 ; 
        RECT 29 85.374 31.52 89.748 ; 
        RECT 0.56 88.844 28.928 89.748 ; 
        RECT 0.02 85.374 0.488 89.748 ; 
        RECT 65.504 85.374 66.116 89.036 ; 
        RECT 37.424 85.374 65.432 89.748 ; 
        RECT 34.436 85.374 37.352 89.036 ; 
        RECT 33.788 86.156 34.292 89.748 ; 
        RECT 28.784 85.772 33.68 89.036 ; 
        RECT 0.704 85.374 28.712 89.748 ; 
        RECT 0.02 85.374 0.632 89.036 ; 
        RECT 34.22 85.374 66.116 88.652 ; 
        RECT 0.02 85.772 34.148 88.652 ; 
        RECT 33.32 85.374 66.116 86.06 ; 
        RECT 0.02 85.374 33.248 88.652 ; 
        RECT 0.02 85.374 66.116 85.676 ; 
        RECT 0.02 93.548 66.116 94.068 ; 
        RECT 65.648 89.694 66.116 94.068 ; 
        RECT 37.208 93.164 65.576 94.068 ; 
        RECT 31.88 93.164 37.136 94.068 ; 
        RECT 29 89.694 31.52 94.068 ; 
        RECT 0.56 93.164 28.928 94.068 ; 
        RECT 0.02 89.694 0.488 94.068 ; 
        RECT 65.504 89.694 66.116 93.356 ; 
        RECT 37.424 89.694 65.432 94.068 ; 
        RECT 34.436 89.694 37.352 93.356 ; 
        RECT 33.788 90.476 34.292 94.068 ; 
        RECT 28.784 90.092 33.68 93.356 ; 
        RECT 0.704 89.694 28.712 94.068 ; 
        RECT 0.02 89.694 0.632 93.356 ; 
        RECT 34.22 89.694 66.116 92.972 ; 
        RECT 0.02 90.092 34.148 92.972 ; 
        RECT 33.32 89.694 66.116 90.38 ; 
        RECT 0.02 89.694 33.248 92.972 ; 
        RECT 0.02 89.694 66.116 89.996 ; 
        RECT 0.02 97.868 66.116 98.388 ; 
        RECT 65.648 94.014 66.116 98.388 ; 
        RECT 37.208 97.484 65.576 98.388 ; 
        RECT 31.88 97.484 37.136 98.388 ; 
        RECT 29 94.014 31.52 98.388 ; 
        RECT 0.56 97.484 28.928 98.388 ; 
        RECT 0.02 94.014 0.488 98.388 ; 
        RECT 65.504 94.014 66.116 97.676 ; 
        RECT 37.424 94.014 65.432 98.388 ; 
        RECT 34.436 94.014 37.352 97.676 ; 
        RECT 33.788 94.796 34.292 98.388 ; 
        RECT 28.784 94.412 33.68 97.676 ; 
        RECT 0.704 94.014 28.712 98.388 ; 
        RECT 0.02 94.014 0.632 97.676 ; 
        RECT 34.22 94.014 66.116 97.292 ; 
        RECT 0.02 94.412 34.148 97.292 ; 
        RECT 33.32 94.014 66.116 94.7 ; 
        RECT 0.02 94.014 33.248 97.292 ; 
        RECT 0.02 94.014 66.116 94.316 ; 
        RECT 0.02 102.188 66.116 102.708 ; 
        RECT 65.648 98.334 66.116 102.708 ; 
        RECT 37.208 101.804 65.576 102.708 ; 
        RECT 31.88 101.804 37.136 102.708 ; 
        RECT 29 98.334 31.52 102.708 ; 
        RECT 0.56 101.804 28.928 102.708 ; 
        RECT 0.02 98.334 0.488 102.708 ; 
        RECT 65.504 98.334 66.116 101.996 ; 
        RECT 37.424 98.334 65.432 102.708 ; 
        RECT 34.436 98.334 37.352 101.996 ; 
        RECT 33.788 99.116 34.292 102.708 ; 
        RECT 28.784 98.732 33.68 101.996 ; 
        RECT 0.704 98.334 28.712 102.708 ; 
        RECT 0.02 98.334 0.632 101.996 ; 
        RECT 34.22 98.334 66.116 101.612 ; 
        RECT 0.02 98.732 34.148 101.612 ; 
        RECT 33.32 98.334 66.116 99.02 ; 
        RECT 0.02 98.334 33.248 101.612 ; 
        RECT 0.02 98.334 66.116 98.636 ; 
        RECT 0.02 106.508 66.116 107.028 ; 
        RECT 65.648 102.654 66.116 107.028 ; 
        RECT 37.208 106.124 65.576 107.028 ; 
        RECT 31.88 106.124 37.136 107.028 ; 
        RECT 29 102.654 31.52 107.028 ; 
        RECT 0.56 106.124 28.928 107.028 ; 
        RECT 0.02 102.654 0.488 107.028 ; 
        RECT 65.504 102.654 66.116 106.316 ; 
        RECT 37.424 102.654 65.432 107.028 ; 
        RECT 34.436 102.654 37.352 106.316 ; 
        RECT 33.788 103.436 34.292 107.028 ; 
        RECT 28.784 103.052 33.68 106.316 ; 
        RECT 0.704 102.654 28.712 107.028 ; 
        RECT 0.02 102.654 0.632 106.316 ; 
        RECT 34.22 102.654 66.116 105.932 ; 
        RECT 0.02 103.052 34.148 105.932 ; 
        RECT 33.32 102.654 66.116 103.34 ; 
        RECT 0.02 102.654 33.248 105.932 ; 
        RECT 0.02 102.654 66.116 102.956 ; 
        RECT 0.02 110.828 66.116 111.348 ; 
        RECT 65.648 106.974 66.116 111.348 ; 
        RECT 37.208 110.444 65.576 111.348 ; 
        RECT 31.88 110.444 37.136 111.348 ; 
        RECT 29 106.974 31.52 111.348 ; 
        RECT 0.56 110.444 28.928 111.348 ; 
        RECT 0.02 106.974 0.488 111.348 ; 
        RECT 65.504 106.974 66.116 110.636 ; 
        RECT 37.424 106.974 65.432 111.348 ; 
        RECT 34.436 106.974 37.352 110.636 ; 
        RECT 33.788 107.756 34.292 111.348 ; 
        RECT 28.784 107.372 33.68 110.636 ; 
        RECT 0.704 106.974 28.712 111.348 ; 
        RECT 0.02 106.974 0.632 110.636 ; 
        RECT 34.22 106.974 66.116 110.252 ; 
        RECT 0.02 107.372 34.148 110.252 ; 
        RECT 33.32 106.974 66.116 107.66 ; 
        RECT 0.02 106.974 33.248 110.252 ; 
        RECT 0.02 106.974 66.116 107.276 ; 
        RECT 0.02 115.148 66.116 115.668 ; 
        RECT 65.648 111.294 66.116 115.668 ; 
        RECT 37.208 114.764 65.576 115.668 ; 
        RECT 31.88 114.764 37.136 115.668 ; 
        RECT 29 111.294 31.52 115.668 ; 
        RECT 0.56 114.764 28.928 115.668 ; 
        RECT 0.02 111.294 0.488 115.668 ; 
        RECT 65.504 111.294 66.116 114.956 ; 
        RECT 37.424 111.294 65.432 115.668 ; 
        RECT 34.436 111.294 37.352 114.956 ; 
        RECT 33.788 112.076 34.292 115.668 ; 
        RECT 28.784 111.692 33.68 114.956 ; 
        RECT 0.704 111.294 28.712 115.668 ; 
        RECT 0.02 111.294 0.632 114.956 ; 
        RECT 34.22 111.294 66.116 114.572 ; 
        RECT 0.02 111.692 34.148 114.572 ; 
        RECT 33.32 111.294 66.116 111.98 ; 
        RECT 0.02 111.294 33.248 114.572 ; 
        RECT 0.02 111.294 66.116 111.596 ; 
        RECT 0.02 119.468 66.116 119.988 ; 
        RECT 65.648 115.614 66.116 119.988 ; 
        RECT 37.208 119.084 65.576 119.988 ; 
        RECT 31.88 119.084 37.136 119.988 ; 
        RECT 29 115.614 31.52 119.988 ; 
        RECT 0.56 119.084 28.928 119.988 ; 
        RECT 0.02 115.614 0.488 119.988 ; 
        RECT 65.504 115.614 66.116 119.276 ; 
        RECT 37.424 115.614 65.432 119.988 ; 
        RECT 34.436 115.614 37.352 119.276 ; 
        RECT 33.788 116.396 34.292 119.988 ; 
        RECT 28.784 116.012 33.68 119.276 ; 
        RECT 0.704 115.614 28.712 119.988 ; 
        RECT 0.02 115.614 0.632 119.276 ; 
        RECT 34.22 115.614 66.116 118.892 ; 
        RECT 0.02 116.012 34.148 118.892 ; 
        RECT 33.32 115.614 66.116 116.3 ; 
        RECT 0.02 115.614 33.248 118.892 ; 
        RECT 0.02 115.614 66.116 115.916 ; 
  LAYER M4 ; 
      RECT 6.276 51 60.038 51.096 ; 
      RECT 6.276 52.152 60.038 52.248 ; 
      RECT 6.276 53.688 60.038 53.784 ; 
      RECT 6.276 54.072 60.038 54.168 ; 
      RECT 6.276 55.416 60.038 55.512 ; 
      RECT 6.276 56.952 60.038 57.048 ; 
      RECT 43.82 46.836 44.156 46.932 ; 
      RECT 43.068 48.564 43.588 48.66 ; 
      RECT 43.1 51.194 43.568 51.29 ; 
      RECT 43.1 52.344 43.568 52.44 ; 
      RECT 40.544 48.564 42.828 48.66 ; 
      RECT 40.784 51.672 41.216 51.768 ; 
      RECT 35.452 53.172 39.824 53.268 ; 
      RECT 38.204 51.444 38.54 51.54 ; 
      RECT 35.068 56.244 38.54 56.34 ; 
      RECT 38.204 56.628 38.54 56.724 ; 
      RECT 37.492 49.524 37.828 49.62 ; 
      RECT 37.34 54.9 37.676 54.996 ; 
      RECT 37.34 57.78 37.676 57.876 ; 
      RECT 36.628 49.14 36.964 49.236 ; 
      RECT 35.772 43.988 36.824 44.084 ; 
      RECT 35.772 78.484 36.824 78.58 ; 
      RECT 35.836 55.092 36.812 55.188 ; 
      RECT 36.476 55.668 36.812 55.764 ; 
      RECT 30.652 56.628 36.812 56.724 ; 
      RECT 36.476 57.78 36.812 57.876 ; 
      RECT 35.54 78.1 36.592 78.196 ; 
      RECT 35.536 43.604 36.588 43.7 ; 
      RECT 35.384 43.22 36.436 43.316 ; 
      RECT 35.384 77.332 36.436 77.428 ; 
      RECT 36.044 59.508 36.38 59.604 ; 
      RECT 32.956 61.044 36.38 61.14 ; 
      RECT 34.492 70.068 36.38 70.164 ; 
      RECT 36.044 70.452 36.38 70.548 ; 
      RECT 35.192 42.836 36.244 42.932 ; 
      RECT 35.192 76.948 36.244 77.044 ; 
      RECT 34.3 66.42 36.08 66.516 ; 
      RECT 35.016 42.452 36.068 42.548 ; 
      RECT 35.016 78.292 36.068 78.388 ; 
      RECT 34.82 43.796 35.872 43.892 ; 
      RECT 34.82 77.908 35.872 78.004 ; 
      RECT 35.344 55.668 35.828 55.764 ; 
      RECT 35.26 64.116 35.792 64.212 ; 
      RECT 34.632 43.412 35.684 43.508 ; 
      RECT 34.632 77.524 35.684 77.62 ; 
      RECT 34.492 42.26 35.544 42.356 ; 
      RECT 34.492 77.14 35.544 77.236 ; 
      RECT 31.228 70.452 35.504 70.548 ; 
      RECT 35.168 75.06 35.504 75.156 ; 
      RECT 34.268 41.684 35.32 41.78 ; 
      RECT 34.268 76.756 35.32 76.852 ; 
      RECT 34.876 59.508 35.216 59.604 ; 
      RECT 30.46 61.812 34.928 61.908 ; 
      RECT 33.04 53.172 34.868 53.268 ; 
      RECT 32.348 44.564 33.416 44.66 ; 
      RECT 32.348 76.18 33.416 76.276 ; 
      RECT 32.896 59.316 33.332 59.412 ; 
      RECT 32.256 44.18 33.224 44.276 ; 
      RECT 32.256 78.676 33.224 78.772 ; 
      RECT 32.032 42.26 33 42.356 ; 
      RECT 32.148 79.06 33 79.156 ; 
      RECT 32.612 57.78 32.948 57.876 ; 
      RECT 31.816 42.644 32.808 42.74 ; 
      RECT 31.816 78.484 32.808 78.58 ; 
      RECT 30.88 68.148 32.564 68.244 ; 
      RECT 30.752 43.988 31.82 44.084 ; 
      RECT 30.752 79.06 31.82 79.156 ; 
      RECT 31.312 62.388 31.796 62.484 ; 
      RECT 31.28 75.06 31.616 75.156 ; 
      RECT 30.616 43.604 31.604 43.7 ; 
      RECT 30.348 77.332 31.604 77.428 ; 
      RECT 30.512 43.22 31.432 43.316 ; 
      RECT 30.464 78.676 31.432 78.772 ; 
      RECT 30.3 42.836 31.22 42.932 ; 
      RECT 30.884 68.724 31.22 68.82 ; 
      RECT 30.1 76.948 31.22 77.044 ; 
      RECT 30.12 42.452 31.04 42.548 ; 
      RECT 30.12 78.292 31.04 78.388 ; 
      RECT 26.272 57.78 31.028 57.876 ; 
      RECT 29.968 43.412 30.888 43.508 ; 
      RECT 29.968 77.908 30.888 78.004 ; 
      RECT 29.896 43.028 30.668 43.124 ; 
      RECT 29.896 77.524 30.668 77.62 ; 
      RECT 29.7 42.644 30.472 42.74 ; 
      RECT 29.7 77.14 30.472 77.236 ; 
      RECT 29.716 61.428 30.452 61.524 ; 
      RECT 29.492 42.26 30.264 42.356 ; 
      RECT 29.492 76.756 30.264 76.852 ; 
      RECT 27.556 50.676 30.26 50.772 ; 
      RECT 29.716 61.812 30.052 61.908 ; 
      RECT 28.64 44.372 29.692 44.468 ; 
      RECT 28.77 59.508 29.304 59.604 ; 
      RECT 27.404 51.444 27.74 51.54 ; 
  LAYER V4 ; 
      RECT 44.016 46.836 44.112 46.932 ; 
      RECT 44.016 51 44.112 51.096 ; 
      RECT 43.344 48.564 43.44 48.66 ; 
      RECT 43.344 51.194 43.44 51.29 ; 
      RECT 43.344 52.344 43.44 52.44 ; 
      RECT 40.848 48.564 40.944 48.66 ; 
      RECT 40.848 51.672 40.944 51.768 ; 
      RECT 38.4 51.444 38.496 51.54 ; 
      RECT 38.4 52.152 38.496 52.248 ; 
      RECT 38.4 56.244 38.496 56.34 ; 
      RECT 38.4 56.628 38.496 56.724 ; 
      RECT 37.536 49.524 37.632 49.62 ; 
      RECT 37.536 53.688 37.632 53.784 ; 
      RECT 37.536 54.9 37.632 54.996 ; 
      RECT 37.536 55.416 37.632 55.512 ; 
      RECT 37.536 56.952 37.632 57.048 ; 
      RECT 37.536 57.78 37.632 57.876 ; 
      RECT 36.672 49.14 36.768 49.236 ; 
      RECT 36.672 54.072 36.768 54.168 ; 
      RECT 36.672 55.092 36.768 55.188 ; 
      RECT 36.672 55.668 36.768 55.764 ; 
      RECT 36.672 56.628 36.768 56.724 ; 
      RECT 36.672 57.78 36.768 57.876 ; 
      RECT 36.24 59.508 36.336 59.604 ; 
      RECT 36.24 61.044 36.336 61.14 ; 
      RECT 36.24 70.068 36.336 70.164 ; 
      RECT 36.24 70.452 36.336 70.548 ; 
      RECT 35.88 43.988 35.976 44.084 ; 
      RECT 35.88 55.092 35.976 55.188 ; 
      RECT 35.88 78.484 35.976 78.58 ; 
      RECT 35.688 43.604 35.784 43.7 ; 
      RECT 35.688 55.668 35.784 55.764 ; 
      RECT 35.688 78.1 35.784 78.196 ; 
      RECT 35.496 43.22 35.592 43.316 ; 
      RECT 35.496 53.172 35.592 53.268 ; 
      RECT 35.496 77.332 35.592 77.428 ; 
      RECT 35.304 42.836 35.4 42.932 ; 
      RECT 35.304 64.116 35.4 64.212 ; 
      RECT 35.304 75.06 35.4 75.156 ; 
      RECT 35.304 76.948 35.4 77.044 ; 
      RECT 35.112 42.452 35.208 42.548 ; 
      RECT 35.112 56.244 35.208 56.34 ; 
      RECT 35.112 78.292 35.208 78.388 ; 
      RECT 34.92 43.796 35.016 43.892 ; 
      RECT 34.92 59.508 35.016 59.604 ; 
      RECT 34.92 77.908 35.016 78.004 ; 
      RECT 34.728 43.412 34.824 43.508 ; 
      RECT 34.728 53.172 34.824 53.268 ; 
      RECT 34.728 77.524 34.824 77.62 ; 
      RECT 34.536 42.26 34.632 42.356 ; 
      RECT 34.536 70.068 34.632 70.164 ; 
      RECT 34.536 77.14 34.632 77.236 ; 
      RECT 34.344 41.684 34.44 41.78 ; 
      RECT 34.344 66.42 34.44 66.516 ; 
      RECT 34.344 76.756 34.44 76.852 ; 
      RECT 33.192 44.564 33.288 44.66 ; 
      RECT 33.192 59.316 33.288 59.412 ; 
      RECT 33.192 76.18 33.288 76.276 ; 
      RECT 33 44.18 33.096 44.276 ; 
      RECT 33 61.044 33.096 61.14 ; 
      RECT 33 78.676 33.096 78.772 ; 
      RECT 32.808 42.26 32.904 42.356 ; 
      RECT 32.808 57.78 32.904 57.876 ; 
      RECT 32.808 79.06 32.904 79.156 ; 
      RECT 32.424 42.644 32.52 42.74 ; 
      RECT 32.424 68.148 32.52 68.244 ; 
      RECT 32.424 78.484 32.52 78.58 ; 
      RECT 31.656 43.988 31.752 44.084 ; 
      RECT 31.656 62.388 31.752 62.484 ; 
      RECT 31.656 79.06 31.752 79.156 ; 
      RECT 31.464 43.604 31.56 43.7 ; 
      RECT 31.464 75.06 31.56 75.156 ; 
      RECT 31.464 77.332 31.56 77.428 ; 
      RECT 31.272 43.22 31.368 43.316 ; 
      RECT 31.272 70.452 31.368 70.548 ; 
      RECT 31.272 78.676 31.368 78.772 ; 
      RECT 31.08 42.836 31.176 42.932 ; 
      RECT 31.08 68.724 31.176 68.82 ; 
      RECT 31.08 76.948 31.176 77.044 ; 
      RECT 30.888 42.452 30.984 42.548 ; 
      RECT 30.888 57.78 30.984 57.876 ; 
      RECT 30.888 78.292 30.984 78.388 ; 
      RECT 30.696 43.412 30.792 43.508 ; 
      RECT 30.696 56.628 30.792 56.724 ; 
      RECT 30.696 77.908 30.792 78.004 ; 
      RECT 30.504 43.028 30.6 43.124 ; 
      RECT 30.504 61.812 30.6 61.908 ; 
      RECT 30.504 77.524 30.6 77.62 ; 
      RECT 30.312 42.644 30.408 42.74 ; 
      RECT 30.312 61.428 30.408 61.524 ; 
      RECT 30.312 77.14 30.408 77.236 ; 
      RECT 30.12 42.26 30.216 42.356 ; 
      RECT 30.12 50.676 30.216 50.772 ; 
      RECT 30.12 76.756 30.216 76.852 ; 
      RECT 29.76 61.428 29.856 61.524 ; 
      RECT 29.76 61.812 29.856 61.908 ; 
      RECT 29.088 44.372 29.184 44.468 ; 
      RECT 29.088 59.508 29.184 59.604 ; 
      RECT 27.6 50.676 27.696 50.772 ; 
      RECT 27.6 51.444 27.696 51.54 ; 
  LAYER M5 ; 
      RECT 44.016 46.792 44.112 51.14 ; 
      RECT 43.344 48.452 43.44 52.694 ; 
      RECT 40.848 48.486 40.944 51.816 ; 
      RECT 38.4 51.4 38.496 52.292 ; 
      RECT 38.4 56.2 38.496 56.768 ; 
      RECT 37.536 49.48 37.632 53.828 ; 
      RECT 37.536 54.856 37.632 55.556 ; 
      RECT 37.536 56.908 37.632 57.92 ; 
      RECT 36.672 49.096 36.768 54.212 ; 
      RECT 36.672 55.048 36.768 55.808 ; 
      RECT 36.672 56.584 36.768 57.92 ; 
      RECT 36.24 59.464 36.336 61.184 ; 
      RECT 36.24 70.024 36.336 70.592 ; 
      RECT 35.88 45.336 35.976 75.668 ; 
      RECT 35.688 45.336 35.784 75.668 ; 
      RECT 35.496 45.336 35.592 75.668 ; 
      RECT 35.304 45.336 35.4 75.668 ; 
      RECT 35.112 45.336 35.208 75.668 ; 
      RECT 34.92 45.336 35.016 75.668 ; 
      RECT 34.728 45.336 34.824 75.668 ; 
      RECT 34.536 45.336 34.632 75.668 ; 
      RECT 34.344 45.336 34.44 75.668 ; 
      RECT 33.192 45.336 33.288 75.668 ; 
      RECT 33 45.336 33.096 75.668 ; 
      RECT 32.808 45.336 32.904 75.668 ; 
      RECT 32.424 45.336 32.52 75.668 ; 
      RECT 31.656 45.336 31.752 75.668 ; 
      RECT 31.464 45.336 31.56 75.668 ; 
      RECT 31.272 45.336 31.368 75.668 ; 
      RECT 31.08 45.336 31.176 75.668 ; 
      RECT 30.888 45.336 30.984 75.668 ; 
      RECT 30.696 45.336 30.792 75.668 ; 
      RECT 30.504 41.968 30.6 78.188 ; 
      RECT 30.312 41.82 30.408 78.004 ; 
      RECT 30.12 41.604 30.216 77.788 ; 
      RECT 29.76 61.384 29.856 61.952 ; 
      RECT 29.088 44.3 29.184 59.676 ; 
      RECT 27.6 50.632 27.696 51.584 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 63.568 120.816 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 63.568 120.816 ; 
  END 
END srambank_128x4x20_6t122 
