VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_256x4x64_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_256x4x64_6t122 0 0 ;
  SIZE 30.348 BY 77.76 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1040 1.1720 30.2580 1.2200 ;
        RECT 0.1040 2.2520 30.2580 2.3000 ;
        RECT 0.1040 3.3320 30.2580 3.3800 ;
        RECT 0.1040 4.4120 30.2580 4.4600 ;
        RECT 0.1040 5.4920 30.2580 5.5400 ;
        RECT 0.1040 6.5720 30.2580 6.6200 ;
        RECT 0.1040 7.6520 30.2580 7.7000 ;
        RECT 0.1040 8.7320 30.2580 8.7800 ;
        RECT 0.1040 9.8120 30.2580 9.8600 ;
        RECT 0.1040 10.8920 30.2580 10.9400 ;
        RECT 0.1040 11.9720 30.2580 12.0200 ;
        RECT 0.1040 13.0520 30.2580 13.1000 ;
        RECT 0.1040 14.1320 30.2580 14.1800 ;
        RECT 0.1040 15.2120 30.2580 15.2600 ;
        RECT 0.1040 16.2920 30.2580 16.3400 ;
        RECT 0.1040 17.3720 30.2580 17.4200 ;
        RECT 0.1040 18.4520 30.2580 18.5000 ;
        RECT 0.1040 19.5320 30.2580 19.5800 ;
        RECT 0.1040 20.6120 30.2580 20.6600 ;
        RECT 0.1040 21.6920 30.2580 21.7400 ;
        RECT 0.1040 22.7720 30.2580 22.8200 ;
        RECT 0.1040 23.8520 30.2580 23.9000 ;
        RECT 0.1040 24.9320 30.2580 24.9800 ;
        RECT 0.1040 26.0120 30.2580 26.0600 ;
        RECT 0.1040 27.0920 30.2580 27.1400 ;
        RECT 0.1040 28.1720 30.2580 28.2200 ;
        RECT 0.1040 29.2520 30.2580 29.3000 ;
        RECT 0.1040 30.3320 30.2580 30.3800 ;
        RECT 0.1040 31.4120 30.2580 31.4600 ;
        RECT 0.1040 32.4920 30.2580 32.5400 ;
        RECT 0.1040 33.5720 30.2580 33.6200 ;
        RECT 0.1040 34.6520 30.2580 34.7000 ;
        RECT 0.1040 43.8590 30.2580 43.9070 ;
        RECT 0.1040 44.9390 30.2580 44.9870 ;
        RECT 0.1040 46.0190 30.2580 46.0670 ;
        RECT 0.1040 47.0990 30.2580 47.1470 ;
        RECT 0.1040 48.1790 30.2580 48.2270 ;
        RECT 0.1040 49.2590 30.2580 49.3070 ;
        RECT 0.1040 50.3390 30.2580 50.3870 ;
        RECT 0.1040 51.4190 30.2580 51.4670 ;
        RECT 0.1040 52.4990 30.2580 52.5470 ;
        RECT 0.1040 53.5790 30.2580 53.6270 ;
        RECT 0.1040 54.6590 30.2580 54.7070 ;
        RECT 0.1040 55.7390 30.2580 55.7870 ;
        RECT 0.1040 56.8190 30.2580 56.8670 ;
        RECT 0.1040 57.8990 30.2580 57.9470 ;
        RECT 0.1040 58.9790 30.2580 59.0270 ;
        RECT 0.1040 60.0590 30.2580 60.1070 ;
        RECT 0.1040 61.1390 30.2580 61.1870 ;
        RECT 0.1040 62.2190 30.2580 62.2670 ;
        RECT 0.1040 63.2990 30.2580 63.3470 ;
        RECT 0.1040 64.3790 30.2580 64.4270 ;
        RECT 0.1040 65.4590 30.2580 65.5070 ;
        RECT 0.1040 66.5390 30.2580 66.5870 ;
        RECT 0.1040 67.6190 30.2580 67.6670 ;
        RECT 0.1040 68.6990 30.2580 68.7470 ;
        RECT 0.1040 69.7790 30.2580 69.8270 ;
        RECT 0.1040 70.8590 30.2580 70.9070 ;
        RECT 0.1040 71.9390 30.2580 71.9870 ;
        RECT 0.1040 73.0190 30.2580 73.0670 ;
        RECT 0.1040 74.0990 30.2580 74.1470 ;
        RECT 0.1040 75.1790 30.2580 75.2270 ;
        RECT 0.1040 76.2590 30.2580 76.3070 ;
        RECT 0.1040 77.3390 30.2580 77.3870 ;
      LAYER M3  ;
        RECT 30.2180 0.2165 30.2360 1.3765 ;
        RECT 16.1960 0.2170 16.2140 1.3760 ;
        RECT 14.7920 0.2530 14.8820 1.3685 ;
        RECT 14.1440 0.2170 14.1620 1.3760 ;
        RECT 0.1220 0.2165 0.1400 1.3765 ;
        RECT 30.2180 1.2965 30.2360 2.4565 ;
        RECT 16.1960 1.2970 16.2140 2.4560 ;
        RECT 14.7920 1.3330 14.8820 2.4485 ;
        RECT 14.1440 1.2970 14.1620 2.4560 ;
        RECT 0.1220 1.2965 0.1400 2.4565 ;
        RECT 30.2180 2.3765 30.2360 3.5365 ;
        RECT 16.1960 2.3770 16.2140 3.5360 ;
        RECT 14.7920 2.4130 14.8820 3.5285 ;
        RECT 14.1440 2.3770 14.1620 3.5360 ;
        RECT 0.1220 2.3765 0.1400 3.5365 ;
        RECT 30.2180 3.4565 30.2360 4.6165 ;
        RECT 16.1960 3.4570 16.2140 4.6160 ;
        RECT 14.7920 3.4930 14.8820 4.6085 ;
        RECT 14.1440 3.4570 14.1620 4.6160 ;
        RECT 0.1220 3.4565 0.1400 4.6165 ;
        RECT 30.2180 4.5365 30.2360 5.6965 ;
        RECT 16.1960 4.5370 16.2140 5.6960 ;
        RECT 14.7920 4.5730 14.8820 5.6885 ;
        RECT 14.1440 4.5370 14.1620 5.6960 ;
        RECT 0.1220 4.5365 0.1400 5.6965 ;
        RECT 30.2180 5.6165 30.2360 6.7765 ;
        RECT 16.1960 5.6170 16.2140 6.7760 ;
        RECT 14.7920 5.6530 14.8820 6.7685 ;
        RECT 14.1440 5.6170 14.1620 6.7760 ;
        RECT 0.1220 5.6165 0.1400 6.7765 ;
        RECT 30.2180 6.6965 30.2360 7.8565 ;
        RECT 16.1960 6.6970 16.2140 7.8560 ;
        RECT 14.7920 6.7330 14.8820 7.8485 ;
        RECT 14.1440 6.6970 14.1620 7.8560 ;
        RECT 0.1220 6.6965 0.1400 7.8565 ;
        RECT 30.2180 7.7765 30.2360 8.9365 ;
        RECT 16.1960 7.7770 16.2140 8.9360 ;
        RECT 14.7920 7.8130 14.8820 8.9285 ;
        RECT 14.1440 7.7770 14.1620 8.9360 ;
        RECT 0.1220 7.7765 0.1400 8.9365 ;
        RECT 30.2180 8.8565 30.2360 10.0165 ;
        RECT 16.1960 8.8570 16.2140 10.0160 ;
        RECT 14.7920 8.8930 14.8820 10.0085 ;
        RECT 14.1440 8.8570 14.1620 10.0160 ;
        RECT 0.1220 8.8565 0.1400 10.0165 ;
        RECT 30.2180 9.9365 30.2360 11.0965 ;
        RECT 16.1960 9.9370 16.2140 11.0960 ;
        RECT 14.7920 9.9730 14.8820 11.0885 ;
        RECT 14.1440 9.9370 14.1620 11.0960 ;
        RECT 0.1220 9.9365 0.1400 11.0965 ;
        RECT 30.2180 11.0165 30.2360 12.1765 ;
        RECT 16.1960 11.0170 16.2140 12.1760 ;
        RECT 14.7920 11.0530 14.8820 12.1685 ;
        RECT 14.1440 11.0170 14.1620 12.1760 ;
        RECT 0.1220 11.0165 0.1400 12.1765 ;
        RECT 30.2180 12.0965 30.2360 13.2565 ;
        RECT 16.1960 12.0970 16.2140 13.2560 ;
        RECT 14.7920 12.1330 14.8820 13.2485 ;
        RECT 14.1440 12.0970 14.1620 13.2560 ;
        RECT 0.1220 12.0965 0.1400 13.2565 ;
        RECT 30.2180 13.1765 30.2360 14.3365 ;
        RECT 16.1960 13.1770 16.2140 14.3360 ;
        RECT 14.7920 13.2130 14.8820 14.3285 ;
        RECT 14.1440 13.1770 14.1620 14.3360 ;
        RECT 0.1220 13.1765 0.1400 14.3365 ;
        RECT 30.2180 14.2565 30.2360 15.4165 ;
        RECT 16.1960 14.2570 16.2140 15.4160 ;
        RECT 14.7920 14.2930 14.8820 15.4085 ;
        RECT 14.1440 14.2570 14.1620 15.4160 ;
        RECT 0.1220 14.2565 0.1400 15.4165 ;
        RECT 30.2180 15.3365 30.2360 16.4965 ;
        RECT 16.1960 15.3370 16.2140 16.4960 ;
        RECT 14.7920 15.3730 14.8820 16.4885 ;
        RECT 14.1440 15.3370 14.1620 16.4960 ;
        RECT 0.1220 15.3365 0.1400 16.4965 ;
        RECT 30.2180 16.4165 30.2360 17.5765 ;
        RECT 16.1960 16.4170 16.2140 17.5760 ;
        RECT 14.7920 16.4530 14.8820 17.5685 ;
        RECT 14.1440 16.4170 14.1620 17.5760 ;
        RECT 0.1220 16.4165 0.1400 17.5765 ;
        RECT 30.2180 17.4965 30.2360 18.6565 ;
        RECT 16.1960 17.4970 16.2140 18.6560 ;
        RECT 14.7920 17.5330 14.8820 18.6485 ;
        RECT 14.1440 17.4970 14.1620 18.6560 ;
        RECT 0.1220 17.4965 0.1400 18.6565 ;
        RECT 30.2180 18.5765 30.2360 19.7365 ;
        RECT 16.1960 18.5770 16.2140 19.7360 ;
        RECT 14.7920 18.6130 14.8820 19.7285 ;
        RECT 14.1440 18.5770 14.1620 19.7360 ;
        RECT 0.1220 18.5765 0.1400 19.7365 ;
        RECT 30.2180 19.6565 30.2360 20.8165 ;
        RECT 16.1960 19.6570 16.2140 20.8160 ;
        RECT 14.7920 19.6930 14.8820 20.8085 ;
        RECT 14.1440 19.6570 14.1620 20.8160 ;
        RECT 0.1220 19.6565 0.1400 20.8165 ;
        RECT 30.2180 20.7365 30.2360 21.8965 ;
        RECT 16.1960 20.7370 16.2140 21.8960 ;
        RECT 14.7920 20.7730 14.8820 21.8885 ;
        RECT 14.1440 20.7370 14.1620 21.8960 ;
        RECT 0.1220 20.7365 0.1400 21.8965 ;
        RECT 30.2180 21.8165 30.2360 22.9765 ;
        RECT 16.1960 21.8170 16.2140 22.9760 ;
        RECT 14.7920 21.8530 14.8820 22.9685 ;
        RECT 14.1440 21.8170 14.1620 22.9760 ;
        RECT 0.1220 21.8165 0.1400 22.9765 ;
        RECT 30.2180 22.8965 30.2360 24.0565 ;
        RECT 16.1960 22.8970 16.2140 24.0560 ;
        RECT 14.7920 22.9330 14.8820 24.0485 ;
        RECT 14.1440 22.8970 14.1620 24.0560 ;
        RECT 0.1220 22.8965 0.1400 24.0565 ;
        RECT 30.2180 23.9765 30.2360 25.1365 ;
        RECT 16.1960 23.9770 16.2140 25.1360 ;
        RECT 14.7920 24.0130 14.8820 25.1285 ;
        RECT 14.1440 23.9770 14.1620 25.1360 ;
        RECT 0.1220 23.9765 0.1400 25.1365 ;
        RECT 30.2180 25.0565 30.2360 26.2165 ;
        RECT 16.1960 25.0570 16.2140 26.2160 ;
        RECT 14.7920 25.0930 14.8820 26.2085 ;
        RECT 14.1440 25.0570 14.1620 26.2160 ;
        RECT 0.1220 25.0565 0.1400 26.2165 ;
        RECT 30.2180 26.1365 30.2360 27.2965 ;
        RECT 16.1960 26.1370 16.2140 27.2960 ;
        RECT 14.7920 26.1730 14.8820 27.2885 ;
        RECT 14.1440 26.1370 14.1620 27.2960 ;
        RECT 0.1220 26.1365 0.1400 27.2965 ;
        RECT 30.2180 27.2165 30.2360 28.3765 ;
        RECT 16.1960 27.2170 16.2140 28.3760 ;
        RECT 14.7920 27.2530 14.8820 28.3685 ;
        RECT 14.1440 27.2170 14.1620 28.3760 ;
        RECT 0.1220 27.2165 0.1400 28.3765 ;
        RECT 30.2180 28.2965 30.2360 29.4565 ;
        RECT 16.1960 28.2970 16.2140 29.4560 ;
        RECT 14.7920 28.3330 14.8820 29.4485 ;
        RECT 14.1440 28.2970 14.1620 29.4560 ;
        RECT 0.1220 28.2965 0.1400 29.4565 ;
        RECT 30.2180 29.3765 30.2360 30.5365 ;
        RECT 16.1960 29.3770 16.2140 30.5360 ;
        RECT 14.7920 29.4130 14.8820 30.5285 ;
        RECT 14.1440 29.3770 14.1620 30.5360 ;
        RECT 0.1220 29.3765 0.1400 30.5365 ;
        RECT 30.2180 30.4565 30.2360 31.6165 ;
        RECT 16.1960 30.4570 16.2140 31.6160 ;
        RECT 14.7920 30.4930 14.8820 31.6085 ;
        RECT 14.1440 30.4570 14.1620 31.6160 ;
        RECT 0.1220 30.4565 0.1400 31.6165 ;
        RECT 30.2180 31.5365 30.2360 32.6965 ;
        RECT 16.1960 31.5370 16.2140 32.6960 ;
        RECT 14.7920 31.5730 14.8820 32.6885 ;
        RECT 14.1440 31.5370 14.1620 32.6960 ;
        RECT 0.1220 31.5365 0.1400 32.6965 ;
        RECT 30.2180 32.6165 30.2360 33.7765 ;
        RECT 16.1960 32.6170 16.2140 33.7760 ;
        RECT 14.7920 32.6530 14.8820 33.7685 ;
        RECT 14.1440 32.6170 14.1620 33.7760 ;
        RECT 0.1220 32.6165 0.1400 33.7765 ;
        RECT 30.2180 33.6965 30.2360 34.8565 ;
        RECT 16.1960 33.6970 16.2140 34.8560 ;
        RECT 14.7920 33.7330 14.8820 34.8485 ;
        RECT 14.1440 33.6970 14.1620 34.8560 ;
        RECT 0.1220 33.6965 0.1400 34.8565 ;
        RECT 14.0490 38.6450 14.0670 44.7085 ;
        RECT 30.2180 42.9035 30.2360 44.0635 ;
        RECT 16.1960 42.9040 16.2140 44.0630 ;
        RECT 14.7920 42.9400 14.8820 44.0555 ;
        RECT 14.1440 42.9040 14.1620 44.0630 ;
        RECT 0.1220 42.9035 0.1400 44.0635 ;
        RECT 30.2180 43.9835 30.2360 45.1435 ;
        RECT 16.1960 43.9840 16.2140 45.1430 ;
        RECT 14.7920 44.0200 14.8820 45.1355 ;
        RECT 14.1440 43.9840 14.1620 45.1430 ;
        RECT 0.1220 43.9835 0.1400 45.1435 ;
        RECT 30.2180 45.0635 30.2360 46.2235 ;
        RECT 16.1960 45.0640 16.2140 46.2230 ;
        RECT 14.7920 45.1000 14.8820 46.2155 ;
        RECT 14.1440 45.0640 14.1620 46.2230 ;
        RECT 0.1220 45.0635 0.1400 46.2235 ;
        RECT 30.2180 46.1435 30.2360 47.3035 ;
        RECT 16.1960 46.1440 16.2140 47.3030 ;
        RECT 14.7920 46.1800 14.8820 47.2955 ;
        RECT 14.1440 46.1440 14.1620 47.3030 ;
        RECT 0.1220 46.1435 0.1400 47.3035 ;
        RECT 30.2180 47.2235 30.2360 48.3835 ;
        RECT 16.1960 47.2240 16.2140 48.3830 ;
        RECT 14.7920 47.2600 14.8820 48.3755 ;
        RECT 14.1440 47.2240 14.1620 48.3830 ;
        RECT 0.1220 47.2235 0.1400 48.3835 ;
        RECT 30.2180 48.3035 30.2360 49.4635 ;
        RECT 16.1960 48.3040 16.2140 49.4630 ;
        RECT 14.7920 48.3400 14.8820 49.4555 ;
        RECT 14.1440 48.3040 14.1620 49.4630 ;
        RECT 0.1220 48.3035 0.1400 49.4635 ;
        RECT 30.2180 49.3835 30.2360 50.5435 ;
        RECT 16.1960 49.3840 16.2140 50.5430 ;
        RECT 14.7920 49.4200 14.8820 50.5355 ;
        RECT 14.1440 49.3840 14.1620 50.5430 ;
        RECT 0.1220 49.3835 0.1400 50.5435 ;
        RECT 30.2180 50.4635 30.2360 51.6235 ;
        RECT 16.1960 50.4640 16.2140 51.6230 ;
        RECT 14.7920 50.5000 14.8820 51.6155 ;
        RECT 14.1440 50.4640 14.1620 51.6230 ;
        RECT 0.1220 50.4635 0.1400 51.6235 ;
        RECT 30.2180 51.5435 30.2360 52.7035 ;
        RECT 16.1960 51.5440 16.2140 52.7030 ;
        RECT 14.7920 51.5800 14.8820 52.6955 ;
        RECT 14.1440 51.5440 14.1620 52.7030 ;
        RECT 0.1220 51.5435 0.1400 52.7035 ;
        RECT 30.2180 52.6235 30.2360 53.7835 ;
        RECT 16.1960 52.6240 16.2140 53.7830 ;
        RECT 14.7920 52.6600 14.8820 53.7755 ;
        RECT 14.1440 52.6240 14.1620 53.7830 ;
        RECT 0.1220 52.6235 0.1400 53.7835 ;
        RECT 30.2180 53.7035 30.2360 54.8635 ;
        RECT 16.1960 53.7040 16.2140 54.8630 ;
        RECT 14.7920 53.7400 14.8820 54.8555 ;
        RECT 14.1440 53.7040 14.1620 54.8630 ;
        RECT 0.1220 53.7035 0.1400 54.8635 ;
        RECT 30.2180 54.7835 30.2360 55.9435 ;
        RECT 16.1960 54.7840 16.2140 55.9430 ;
        RECT 14.7920 54.8200 14.8820 55.9355 ;
        RECT 14.1440 54.7840 14.1620 55.9430 ;
        RECT 0.1220 54.7835 0.1400 55.9435 ;
        RECT 30.2180 55.8635 30.2360 57.0235 ;
        RECT 16.1960 55.8640 16.2140 57.0230 ;
        RECT 14.7920 55.9000 14.8820 57.0155 ;
        RECT 14.1440 55.8640 14.1620 57.0230 ;
        RECT 0.1220 55.8635 0.1400 57.0235 ;
        RECT 30.2180 56.9435 30.2360 58.1035 ;
        RECT 16.1960 56.9440 16.2140 58.1030 ;
        RECT 14.7920 56.9800 14.8820 58.0955 ;
        RECT 14.1440 56.9440 14.1620 58.1030 ;
        RECT 0.1220 56.9435 0.1400 58.1035 ;
        RECT 30.2180 58.0235 30.2360 59.1835 ;
        RECT 16.1960 58.0240 16.2140 59.1830 ;
        RECT 14.7920 58.0600 14.8820 59.1755 ;
        RECT 14.1440 58.0240 14.1620 59.1830 ;
        RECT 0.1220 58.0235 0.1400 59.1835 ;
        RECT 30.2180 59.1035 30.2360 60.2635 ;
        RECT 16.1960 59.1040 16.2140 60.2630 ;
        RECT 14.7920 59.1400 14.8820 60.2555 ;
        RECT 14.1440 59.1040 14.1620 60.2630 ;
        RECT 0.1220 59.1035 0.1400 60.2635 ;
        RECT 30.2180 60.1835 30.2360 61.3435 ;
        RECT 16.1960 60.1840 16.2140 61.3430 ;
        RECT 14.7920 60.2200 14.8820 61.3355 ;
        RECT 14.1440 60.1840 14.1620 61.3430 ;
        RECT 0.1220 60.1835 0.1400 61.3435 ;
        RECT 30.2180 61.2635 30.2360 62.4235 ;
        RECT 16.1960 61.2640 16.2140 62.4230 ;
        RECT 14.7920 61.3000 14.8820 62.4155 ;
        RECT 14.1440 61.2640 14.1620 62.4230 ;
        RECT 0.1220 61.2635 0.1400 62.4235 ;
        RECT 30.2180 62.3435 30.2360 63.5035 ;
        RECT 16.1960 62.3440 16.2140 63.5030 ;
        RECT 14.7920 62.3800 14.8820 63.4955 ;
        RECT 14.1440 62.3440 14.1620 63.5030 ;
        RECT 0.1220 62.3435 0.1400 63.5035 ;
        RECT 30.2180 63.4235 30.2360 64.5835 ;
        RECT 16.1960 63.4240 16.2140 64.5830 ;
        RECT 14.7920 63.4600 14.8820 64.5755 ;
        RECT 14.1440 63.4240 14.1620 64.5830 ;
        RECT 0.1220 63.4235 0.1400 64.5835 ;
        RECT 30.2180 64.5035 30.2360 65.6635 ;
        RECT 16.1960 64.5040 16.2140 65.6630 ;
        RECT 14.7920 64.5400 14.8820 65.6555 ;
        RECT 14.1440 64.5040 14.1620 65.6630 ;
        RECT 0.1220 64.5035 0.1400 65.6635 ;
        RECT 30.2180 65.5835 30.2360 66.7435 ;
        RECT 16.1960 65.5840 16.2140 66.7430 ;
        RECT 14.7920 65.6200 14.8820 66.7355 ;
        RECT 14.1440 65.5840 14.1620 66.7430 ;
        RECT 0.1220 65.5835 0.1400 66.7435 ;
        RECT 30.2180 66.6635 30.2360 67.8235 ;
        RECT 16.1960 66.6640 16.2140 67.8230 ;
        RECT 14.7920 66.7000 14.8820 67.8155 ;
        RECT 14.1440 66.6640 14.1620 67.8230 ;
        RECT 0.1220 66.6635 0.1400 67.8235 ;
        RECT 30.2180 67.7435 30.2360 68.9035 ;
        RECT 16.1960 67.7440 16.2140 68.9030 ;
        RECT 14.7920 67.7800 14.8820 68.8955 ;
        RECT 14.1440 67.7440 14.1620 68.9030 ;
        RECT 0.1220 67.7435 0.1400 68.9035 ;
        RECT 30.2180 68.8235 30.2360 69.9835 ;
        RECT 16.1960 68.8240 16.2140 69.9830 ;
        RECT 14.7920 68.8600 14.8820 69.9755 ;
        RECT 14.1440 68.8240 14.1620 69.9830 ;
        RECT 0.1220 68.8235 0.1400 69.9835 ;
        RECT 30.2180 69.9035 30.2360 71.0635 ;
        RECT 16.1960 69.9040 16.2140 71.0630 ;
        RECT 14.7920 69.9400 14.8820 71.0555 ;
        RECT 14.1440 69.9040 14.1620 71.0630 ;
        RECT 0.1220 69.9035 0.1400 71.0635 ;
        RECT 30.2180 70.9835 30.2360 72.1435 ;
        RECT 16.1960 70.9840 16.2140 72.1430 ;
        RECT 14.7920 71.0200 14.8820 72.1355 ;
        RECT 14.1440 70.9840 14.1620 72.1430 ;
        RECT 0.1220 70.9835 0.1400 72.1435 ;
        RECT 30.2180 72.0635 30.2360 73.2235 ;
        RECT 16.1960 72.0640 16.2140 73.2230 ;
        RECT 14.7920 72.1000 14.8820 73.2155 ;
        RECT 14.1440 72.0640 14.1620 73.2230 ;
        RECT 0.1220 72.0635 0.1400 73.2235 ;
        RECT 30.2180 73.1435 30.2360 74.3035 ;
        RECT 16.1960 73.1440 16.2140 74.3030 ;
        RECT 14.7920 73.1800 14.8820 74.2955 ;
        RECT 14.1440 73.1440 14.1620 74.3030 ;
        RECT 0.1220 73.1435 0.1400 74.3035 ;
        RECT 30.2180 74.2235 30.2360 75.3835 ;
        RECT 16.1960 74.2240 16.2140 75.3830 ;
        RECT 14.7920 74.2600 14.8820 75.3755 ;
        RECT 14.1440 74.2240 14.1620 75.3830 ;
        RECT 0.1220 74.2235 0.1400 75.3835 ;
        RECT 30.2180 75.3035 30.2360 76.4635 ;
        RECT 16.1960 75.3040 16.2140 76.4630 ;
        RECT 14.7920 75.3400 14.8820 76.4555 ;
        RECT 14.1440 75.3040 14.1620 76.4630 ;
        RECT 0.1220 75.3035 0.1400 76.4635 ;
        RECT 30.2180 76.3835 30.2360 77.5435 ;
        RECT 16.1960 76.3840 16.2140 77.5430 ;
        RECT 14.7920 76.4200 14.8820 77.5355 ;
        RECT 14.1440 76.3840 14.1620 77.5430 ;
        RECT 0.1220 76.3835 0.1400 77.5435 ;
      LAYER V3  ;
        RECT 0.1220 1.1720 0.1400 1.2200 ;
        RECT 14.1440 1.1720 14.1620 1.2200 ;
        RECT 14.7920 1.1720 14.8820 1.2200 ;
        RECT 16.1960 1.1720 16.2140 1.2200 ;
        RECT 30.2180 1.1720 30.2360 1.2200 ;
        RECT 0.1220 2.2520 0.1400 2.3000 ;
        RECT 14.1440 2.2520 14.1620 2.3000 ;
        RECT 14.7920 2.2520 14.8820 2.3000 ;
        RECT 16.1960 2.2520 16.2140 2.3000 ;
        RECT 30.2180 2.2520 30.2360 2.3000 ;
        RECT 0.1220 3.3320 0.1400 3.3800 ;
        RECT 14.1440 3.3320 14.1620 3.3800 ;
        RECT 14.7920 3.3320 14.8820 3.3800 ;
        RECT 16.1960 3.3320 16.2140 3.3800 ;
        RECT 30.2180 3.3320 30.2360 3.3800 ;
        RECT 0.1220 4.4120 0.1400 4.4600 ;
        RECT 14.1440 4.4120 14.1620 4.4600 ;
        RECT 14.7920 4.4120 14.8820 4.4600 ;
        RECT 16.1960 4.4120 16.2140 4.4600 ;
        RECT 30.2180 4.4120 30.2360 4.4600 ;
        RECT 0.1220 5.4920 0.1400 5.5400 ;
        RECT 14.1440 5.4920 14.1620 5.5400 ;
        RECT 14.7920 5.4920 14.8820 5.5400 ;
        RECT 16.1960 5.4920 16.2140 5.5400 ;
        RECT 30.2180 5.4920 30.2360 5.5400 ;
        RECT 0.1220 6.5720 0.1400 6.6200 ;
        RECT 14.1440 6.5720 14.1620 6.6200 ;
        RECT 14.7920 6.5720 14.8820 6.6200 ;
        RECT 16.1960 6.5720 16.2140 6.6200 ;
        RECT 30.2180 6.5720 30.2360 6.6200 ;
        RECT 0.1220 7.6520 0.1400 7.7000 ;
        RECT 14.1440 7.6520 14.1620 7.7000 ;
        RECT 14.7920 7.6520 14.8820 7.7000 ;
        RECT 16.1960 7.6520 16.2140 7.7000 ;
        RECT 30.2180 7.6520 30.2360 7.7000 ;
        RECT 0.1220 8.7320 0.1400 8.7800 ;
        RECT 14.1440 8.7320 14.1620 8.7800 ;
        RECT 14.7920 8.7320 14.8820 8.7800 ;
        RECT 16.1960 8.7320 16.2140 8.7800 ;
        RECT 30.2180 8.7320 30.2360 8.7800 ;
        RECT 0.1220 9.8120 0.1400 9.8600 ;
        RECT 14.1440 9.8120 14.1620 9.8600 ;
        RECT 14.7920 9.8120 14.8820 9.8600 ;
        RECT 16.1960 9.8120 16.2140 9.8600 ;
        RECT 30.2180 9.8120 30.2360 9.8600 ;
        RECT 0.1220 10.8920 0.1400 10.9400 ;
        RECT 14.1440 10.8920 14.1620 10.9400 ;
        RECT 14.7920 10.8920 14.8820 10.9400 ;
        RECT 16.1960 10.8920 16.2140 10.9400 ;
        RECT 30.2180 10.8920 30.2360 10.9400 ;
        RECT 0.1220 11.9720 0.1400 12.0200 ;
        RECT 14.1440 11.9720 14.1620 12.0200 ;
        RECT 14.7920 11.9720 14.8820 12.0200 ;
        RECT 16.1960 11.9720 16.2140 12.0200 ;
        RECT 30.2180 11.9720 30.2360 12.0200 ;
        RECT 0.1220 13.0520 0.1400 13.1000 ;
        RECT 14.1440 13.0520 14.1620 13.1000 ;
        RECT 14.7920 13.0520 14.8820 13.1000 ;
        RECT 16.1960 13.0520 16.2140 13.1000 ;
        RECT 30.2180 13.0520 30.2360 13.1000 ;
        RECT 0.1220 14.1320 0.1400 14.1800 ;
        RECT 14.1440 14.1320 14.1620 14.1800 ;
        RECT 14.7920 14.1320 14.8820 14.1800 ;
        RECT 16.1960 14.1320 16.2140 14.1800 ;
        RECT 30.2180 14.1320 30.2360 14.1800 ;
        RECT 0.1220 15.2120 0.1400 15.2600 ;
        RECT 14.1440 15.2120 14.1620 15.2600 ;
        RECT 14.7920 15.2120 14.8820 15.2600 ;
        RECT 16.1960 15.2120 16.2140 15.2600 ;
        RECT 30.2180 15.2120 30.2360 15.2600 ;
        RECT 0.1220 16.2920 0.1400 16.3400 ;
        RECT 14.1440 16.2920 14.1620 16.3400 ;
        RECT 14.7920 16.2920 14.8820 16.3400 ;
        RECT 16.1960 16.2920 16.2140 16.3400 ;
        RECT 30.2180 16.2920 30.2360 16.3400 ;
        RECT 0.1220 17.3720 0.1400 17.4200 ;
        RECT 14.1440 17.3720 14.1620 17.4200 ;
        RECT 14.7920 17.3720 14.8820 17.4200 ;
        RECT 16.1960 17.3720 16.2140 17.4200 ;
        RECT 30.2180 17.3720 30.2360 17.4200 ;
        RECT 0.1220 18.4520 0.1400 18.5000 ;
        RECT 14.1440 18.4520 14.1620 18.5000 ;
        RECT 14.7920 18.4520 14.8820 18.5000 ;
        RECT 16.1960 18.4520 16.2140 18.5000 ;
        RECT 30.2180 18.4520 30.2360 18.5000 ;
        RECT 0.1220 19.5320 0.1400 19.5800 ;
        RECT 14.1440 19.5320 14.1620 19.5800 ;
        RECT 14.7920 19.5320 14.8820 19.5800 ;
        RECT 16.1960 19.5320 16.2140 19.5800 ;
        RECT 30.2180 19.5320 30.2360 19.5800 ;
        RECT 0.1220 20.6120 0.1400 20.6600 ;
        RECT 14.1440 20.6120 14.1620 20.6600 ;
        RECT 14.7920 20.6120 14.8820 20.6600 ;
        RECT 16.1960 20.6120 16.2140 20.6600 ;
        RECT 30.2180 20.6120 30.2360 20.6600 ;
        RECT 0.1220 21.6920 0.1400 21.7400 ;
        RECT 14.1440 21.6920 14.1620 21.7400 ;
        RECT 14.7920 21.6920 14.8820 21.7400 ;
        RECT 16.1960 21.6920 16.2140 21.7400 ;
        RECT 30.2180 21.6920 30.2360 21.7400 ;
        RECT 0.1220 22.7720 0.1400 22.8200 ;
        RECT 14.1440 22.7720 14.1620 22.8200 ;
        RECT 14.7920 22.7720 14.8820 22.8200 ;
        RECT 16.1960 22.7720 16.2140 22.8200 ;
        RECT 30.2180 22.7720 30.2360 22.8200 ;
        RECT 0.1220 23.8520 0.1400 23.9000 ;
        RECT 14.1440 23.8520 14.1620 23.9000 ;
        RECT 14.7920 23.8520 14.8820 23.9000 ;
        RECT 16.1960 23.8520 16.2140 23.9000 ;
        RECT 30.2180 23.8520 30.2360 23.9000 ;
        RECT 0.1220 24.9320 0.1400 24.9800 ;
        RECT 14.1440 24.9320 14.1620 24.9800 ;
        RECT 14.7920 24.9320 14.8820 24.9800 ;
        RECT 16.1960 24.9320 16.2140 24.9800 ;
        RECT 30.2180 24.9320 30.2360 24.9800 ;
        RECT 0.1220 26.0120 0.1400 26.0600 ;
        RECT 14.1440 26.0120 14.1620 26.0600 ;
        RECT 14.7920 26.0120 14.8820 26.0600 ;
        RECT 16.1960 26.0120 16.2140 26.0600 ;
        RECT 30.2180 26.0120 30.2360 26.0600 ;
        RECT 0.1220 27.0920 0.1400 27.1400 ;
        RECT 14.1440 27.0920 14.1620 27.1400 ;
        RECT 14.7920 27.0920 14.8820 27.1400 ;
        RECT 16.1960 27.0920 16.2140 27.1400 ;
        RECT 30.2180 27.0920 30.2360 27.1400 ;
        RECT 0.1220 28.1720 0.1400 28.2200 ;
        RECT 14.1440 28.1720 14.1620 28.2200 ;
        RECT 14.7920 28.1720 14.8820 28.2200 ;
        RECT 16.1960 28.1720 16.2140 28.2200 ;
        RECT 30.2180 28.1720 30.2360 28.2200 ;
        RECT 0.1220 29.2520 0.1400 29.3000 ;
        RECT 14.1440 29.2520 14.1620 29.3000 ;
        RECT 14.7920 29.2520 14.8820 29.3000 ;
        RECT 16.1960 29.2520 16.2140 29.3000 ;
        RECT 30.2180 29.2520 30.2360 29.3000 ;
        RECT 0.1220 30.3320 0.1400 30.3800 ;
        RECT 14.1440 30.3320 14.1620 30.3800 ;
        RECT 14.7920 30.3320 14.8820 30.3800 ;
        RECT 16.1960 30.3320 16.2140 30.3800 ;
        RECT 30.2180 30.3320 30.2360 30.3800 ;
        RECT 0.1220 31.4120 0.1400 31.4600 ;
        RECT 14.1440 31.4120 14.1620 31.4600 ;
        RECT 14.7920 31.4120 14.8820 31.4600 ;
        RECT 16.1960 31.4120 16.2140 31.4600 ;
        RECT 30.2180 31.4120 30.2360 31.4600 ;
        RECT 0.1220 32.4920 0.1400 32.5400 ;
        RECT 14.1440 32.4920 14.1620 32.5400 ;
        RECT 14.7920 32.4920 14.8820 32.5400 ;
        RECT 16.1960 32.4920 16.2140 32.5400 ;
        RECT 30.2180 32.4920 30.2360 32.5400 ;
        RECT 0.1220 33.5720 0.1400 33.6200 ;
        RECT 14.1440 33.5720 14.1620 33.6200 ;
        RECT 14.7920 33.5720 14.8820 33.6200 ;
        RECT 16.1960 33.5720 16.2140 33.6200 ;
        RECT 30.2180 33.5720 30.2360 33.6200 ;
        RECT 0.1220 34.6520 0.1400 34.7000 ;
        RECT 14.1440 34.6520 14.1620 34.7000 ;
        RECT 14.7920 34.6520 14.8820 34.7000 ;
        RECT 16.1960 34.6520 16.2140 34.7000 ;
        RECT 30.2180 34.6520 30.2360 34.7000 ;
        RECT 0.1220 43.8590 0.1400 43.9070 ;
        RECT 14.1440 43.8590 14.1620 43.9070 ;
        RECT 14.7920 43.8590 14.8820 43.9070 ;
        RECT 16.1960 43.8590 16.2140 43.9070 ;
        RECT 30.2180 43.8590 30.2360 43.9070 ;
        RECT 0.1220 44.9390 0.1400 44.9870 ;
        RECT 14.1440 44.9390 14.1620 44.9870 ;
        RECT 14.7920 44.9390 14.8820 44.9870 ;
        RECT 16.1960 44.9390 16.2140 44.9870 ;
        RECT 30.2180 44.9390 30.2360 44.9870 ;
        RECT 0.1220 46.0190 0.1400 46.0670 ;
        RECT 14.1440 46.0190 14.1620 46.0670 ;
        RECT 14.7920 46.0190 14.8820 46.0670 ;
        RECT 16.1960 46.0190 16.2140 46.0670 ;
        RECT 30.2180 46.0190 30.2360 46.0670 ;
        RECT 0.1220 47.0990 0.1400 47.1470 ;
        RECT 14.1440 47.0990 14.1620 47.1470 ;
        RECT 14.7920 47.0990 14.8820 47.1470 ;
        RECT 16.1960 47.0990 16.2140 47.1470 ;
        RECT 30.2180 47.0990 30.2360 47.1470 ;
        RECT 0.1220 48.1790 0.1400 48.2270 ;
        RECT 14.1440 48.1790 14.1620 48.2270 ;
        RECT 14.7920 48.1790 14.8820 48.2270 ;
        RECT 16.1960 48.1790 16.2140 48.2270 ;
        RECT 30.2180 48.1790 30.2360 48.2270 ;
        RECT 0.1220 49.2590 0.1400 49.3070 ;
        RECT 14.1440 49.2590 14.1620 49.3070 ;
        RECT 14.7920 49.2590 14.8820 49.3070 ;
        RECT 16.1960 49.2590 16.2140 49.3070 ;
        RECT 30.2180 49.2590 30.2360 49.3070 ;
        RECT 0.1220 50.3390 0.1400 50.3870 ;
        RECT 14.1440 50.3390 14.1620 50.3870 ;
        RECT 14.7920 50.3390 14.8820 50.3870 ;
        RECT 16.1960 50.3390 16.2140 50.3870 ;
        RECT 30.2180 50.3390 30.2360 50.3870 ;
        RECT 0.1220 51.4190 0.1400 51.4670 ;
        RECT 14.1440 51.4190 14.1620 51.4670 ;
        RECT 14.7920 51.4190 14.8820 51.4670 ;
        RECT 16.1960 51.4190 16.2140 51.4670 ;
        RECT 30.2180 51.4190 30.2360 51.4670 ;
        RECT 0.1220 52.4990 0.1400 52.5470 ;
        RECT 14.1440 52.4990 14.1620 52.5470 ;
        RECT 14.7920 52.4990 14.8820 52.5470 ;
        RECT 16.1960 52.4990 16.2140 52.5470 ;
        RECT 30.2180 52.4990 30.2360 52.5470 ;
        RECT 0.1220 53.5790 0.1400 53.6270 ;
        RECT 14.1440 53.5790 14.1620 53.6270 ;
        RECT 14.7920 53.5790 14.8820 53.6270 ;
        RECT 16.1960 53.5790 16.2140 53.6270 ;
        RECT 30.2180 53.5790 30.2360 53.6270 ;
        RECT 0.1220 54.6590 0.1400 54.7070 ;
        RECT 14.1440 54.6590 14.1620 54.7070 ;
        RECT 14.7920 54.6590 14.8820 54.7070 ;
        RECT 16.1960 54.6590 16.2140 54.7070 ;
        RECT 30.2180 54.6590 30.2360 54.7070 ;
        RECT 0.1220 55.7390 0.1400 55.7870 ;
        RECT 14.1440 55.7390 14.1620 55.7870 ;
        RECT 14.7920 55.7390 14.8820 55.7870 ;
        RECT 16.1960 55.7390 16.2140 55.7870 ;
        RECT 30.2180 55.7390 30.2360 55.7870 ;
        RECT 0.1220 56.8190 0.1400 56.8670 ;
        RECT 14.1440 56.8190 14.1620 56.8670 ;
        RECT 14.7920 56.8190 14.8820 56.8670 ;
        RECT 16.1960 56.8190 16.2140 56.8670 ;
        RECT 30.2180 56.8190 30.2360 56.8670 ;
        RECT 0.1220 57.8990 0.1400 57.9470 ;
        RECT 14.1440 57.8990 14.1620 57.9470 ;
        RECT 14.7920 57.8990 14.8820 57.9470 ;
        RECT 16.1960 57.8990 16.2140 57.9470 ;
        RECT 30.2180 57.8990 30.2360 57.9470 ;
        RECT 0.1220 58.9790 0.1400 59.0270 ;
        RECT 14.1440 58.9790 14.1620 59.0270 ;
        RECT 14.7920 58.9790 14.8820 59.0270 ;
        RECT 16.1960 58.9790 16.2140 59.0270 ;
        RECT 30.2180 58.9790 30.2360 59.0270 ;
        RECT 0.1220 60.0590 0.1400 60.1070 ;
        RECT 14.1440 60.0590 14.1620 60.1070 ;
        RECT 14.7920 60.0590 14.8820 60.1070 ;
        RECT 16.1960 60.0590 16.2140 60.1070 ;
        RECT 30.2180 60.0590 30.2360 60.1070 ;
        RECT 0.1220 61.1390 0.1400 61.1870 ;
        RECT 14.1440 61.1390 14.1620 61.1870 ;
        RECT 14.7920 61.1390 14.8820 61.1870 ;
        RECT 16.1960 61.1390 16.2140 61.1870 ;
        RECT 30.2180 61.1390 30.2360 61.1870 ;
        RECT 0.1220 62.2190 0.1400 62.2670 ;
        RECT 14.1440 62.2190 14.1620 62.2670 ;
        RECT 14.7920 62.2190 14.8820 62.2670 ;
        RECT 16.1960 62.2190 16.2140 62.2670 ;
        RECT 30.2180 62.2190 30.2360 62.2670 ;
        RECT 0.1220 63.2990 0.1400 63.3470 ;
        RECT 14.1440 63.2990 14.1620 63.3470 ;
        RECT 14.7920 63.2990 14.8820 63.3470 ;
        RECT 16.1960 63.2990 16.2140 63.3470 ;
        RECT 30.2180 63.2990 30.2360 63.3470 ;
        RECT 0.1220 64.3790 0.1400 64.4270 ;
        RECT 14.1440 64.3790 14.1620 64.4270 ;
        RECT 14.7920 64.3790 14.8820 64.4270 ;
        RECT 16.1960 64.3790 16.2140 64.4270 ;
        RECT 30.2180 64.3790 30.2360 64.4270 ;
        RECT 0.1220 65.4590 0.1400 65.5070 ;
        RECT 14.1440 65.4590 14.1620 65.5070 ;
        RECT 14.7920 65.4590 14.8820 65.5070 ;
        RECT 16.1960 65.4590 16.2140 65.5070 ;
        RECT 30.2180 65.4590 30.2360 65.5070 ;
        RECT 0.1220 66.5390 0.1400 66.5870 ;
        RECT 14.1440 66.5390 14.1620 66.5870 ;
        RECT 14.7920 66.5390 14.8820 66.5870 ;
        RECT 16.1960 66.5390 16.2140 66.5870 ;
        RECT 30.2180 66.5390 30.2360 66.5870 ;
        RECT 0.1220 67.6190 0.1400 67.6670 ;
        RECT 14.1440 67.6190 14.1620 67.6670 ;
        RECT 14.7920 67.6190 14.8820 67.6670 ;
        RECT 16.1960 67.6190 16.2140 67.6670 ;
        RECT 30.2180 67.6190 30.2360 67.6670 ;
        RECT 0.1220 68.6990 0.1400 68.7470 ;
        RECT 14.1440 68.6990 14.1620 68.7470 ;
        RECT 14.7920 68.6990 14.8820 68.7470 ;
        RECT 16.1960 68.6990 16.2140 68.7470 ;
        RECT 30.2180 68.6990 30.2360 68.7470 ;
        RECT 0.1220 69.7790 0.1400 69.8270 ;
        RECT 14.1440 69.7790 14.1620 69.8270 ;
        RECT 14.7920 69.7790 14.8820 69.8270 ;
        RECT 16.1960 69.7790 16.2140 69.8270 ;
        RECT 30.2180 69.7790 30.2360 69.8270 ;
        RECT 0.1220 70.8590 0.1400 70.9070 ;
        RECT 14.1440 70.8590 14.1620 70.9070 ;
        RECT 14.7920 70.8590 14.8820 70.9070 ;
        RECT 16.1960 70.8590 16.2140 70.9070 ;
        RECT 30.2180 70.8590 30.2360 70.9070 ;
        RECT 0.1220 71.9390 0.1400 71.9870 ;
        RECT 14.1440 71.9390 14.1620 71.9870 ;
        RECT 14.7920 71.9390 14.8820 71.9870 ;
        RECT 16.1960 71.9390 16.2140 71.9870 ;
        RECT 30.2180 71.9390 30.2360 71.9870 ;
        RECT 0.1220 73.0190 0.1400 73.0670 ;
        RECT 14.1440 73.0190 14.1620 73.0670 ;
        RECT 14.7920 73.0190 14.8820 73.0670 ;
        RECT 16.1960 73.0190 16.2140 73.0670 ;
        RECT 30.2180 73.0190 30.2360 73.0670 ;
        RECT 0.1220 74.0990 0.1400 74.1470 ;
        RECT 14.1440 74.0990 14.1620 74.1470 ;
        RECT 14.7920 74.0990 14.8820 74.1470 ;
        RECT 16.1960 74.0990 16.2140 74.1470 ;
        RECT 30.2180 74.0990 30.2360 74.1470 ;
        RECT 0.1220 75.1790 0.1400 75.2270 ;
        RECT 14.1440 75.1790 14.1620 75.2270 ;
        RECT 14.7920 75.1790 14.8820 75.2270 ;
        RECT 16.1960 75.1790 16.2140 75.2270 ;
        RECT 30.2180 75.1790 30.2360 75.2270 ;
        RECT 0.1220 76.2590 0.1400 76.3070 ;
        RECT 14.1440 76.2590 14.1620 76.3070 ;
        RECT 14.7920 76.2590 14.8820 76.3070 ;
        RECT 16.1960 76.2590 16.2140 76.3070 ;
        RECT 30.2180 76.2590 30.2360 76.3070 ;
        RECT 0.1220 77.3390 0.1400 77.3870 ;
        RECT 14.1440 77.3390 14.1620 77.3870 ;
        RECT 14.7920 77.3390 14.8820 77.3870 ;
        RECT 16.1960 77.3390 16.2140 77.3870 ;
        RECT 30.2180 77.3390 30.2360 77.3870 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1040 1.0760 30.2580 1.1240 ;
        RECT 0.1040 2.1560 30.2580 2.2040 ;
        RECT 0.1040 3.2360 30.2580 3.2840 ;
        RECT 0.1040 4.3160 30.2580 4.3640 ;
        RECT 0.1040 5.3960 30.2580 5.4440 ;
        RECT 0.1040 6.4760 30.2580 6.5240 ;
        RECT 0.1040 7.5560 30.2580 7.6040 ;
        RECT 0.1040 8.6360 30.2580 8.6840 ;
        RECT 0.1040 9.7160 30.2580 9.7640 ;
        RECT 0.1040 10.7960 30.2580 10.8440 ;
        RECT 0.1040 11.8760 30.2580 11.9240 ;
        RECT 0.1040 12.9560 30.2580 13.0040 ;
        RECT 0.1040 14.0360 30.2580 14.0840 ;
        RECT 0.1040 15.1160 30.2580 15.1640 ;
        RECT 0.1040 16.1960 30.2580 16.2440 ;
        RECT 0.1040 17.2760 30.2580 17.3240 ;
        RECT 0.1040 18.3560 30.2580 18.4040 ;
        RECT 0.1040 19.4360 30.2580 19.4840 ;
        RECT 0.1040 20.5160 30.2580 20.5640 ;
        RECT 0.1040 21.5960 30.2580 21.6440 ;
        RECT 0.1040 22.6760 30.2580 22.7240 ;
        RECT 0.1040 23.7560 30.2580 23.8040 ;
        RECT 0.1040 24.8360 30.2580 24.8840 ;
        RECT 0.1040 25.9160 30.2580 25.9640 ;
        RECT 0.1040 26.9960 30.2580 27.0440 ;
        RECT 0.1040 28.0760 30.2580 28.1240 ;
        RECT 0.1040 29.1560 30.2580 29.2040 ;
        RECT 0.1040 30.2360 30.2580 30.2840 ;
        RECT 0.1040 31.3160 30.2580 31.3640 ;
        RECT 0.1040 32.3960 30.2580 32.4440 ;
        RECT 0.1040 33.4760 30.2580 33.5240 ;
        RECT 0.1040 34.5560 30.2580 34.6040 ;
        RECT 10.4760 35.6215 19.8720 35.8375 ;
        RECT 14.3100 38.7895 16.0380 39.0055 ;
        RECT 14.3100 41.9575 16.0380 42.1735 ;
        RECT 0.1040 43.7630 30.2580 43.8110 ;
        RECT 0.1040 44.8430 30.2580 44.8910 ;
        RECT 0.1040 45.9230 30.2580 45.9710 ;
        RECT 0.1040 47.0030 30.2580 47.0510 ;
        RECT 0.1040 48.0830 30.2580 48.1310 ;
        RECT 0.1040 49.1630 30.2580 49.2110 ;
        RECT 0.1040 50.2430 30.2580 50.2910 ;
        RECT 0.1040 51.3230 30.2580 51.3710 ;
        RECT 0.1040 52.4030 30.2580 52.4510 ;
        RECT 0.1040 53.4830 30.2580 53.5310 ;
        RECT 0.1040 54.5630 30.2580 54.6110 ;
        RECT 0.1040 55.6430 30.2580 55.6910 ;
        RECT 0.1040 56.7230 30.2580 56.7710 ;
        RECT 0.1040 57.8030 30.2580 57.8510 ;
        RECT 0.1040 58.8830 30.2580 58.9310 ;
        RECT 0.1040 59.9630 30.2580 60.0110 ;
        RECT 0.1040 61.0430 30.2580 61.0910 ;
        RECT 0.1040 62.1230 30.2580 62.1710 ;
        RECT 0.1040 63.2030 30.2580 63.2510 ;
        RECT 0.1040 64.2830 30.2580 64.3310 ;
        RECT 0.1040 65.3630 30.2580 65.4110 ;
        RECT 0.1040 66.4430 30.2580 66.4910 ;
        RECT 0.1040 67.5230 30.2580 67.5710 ;
        RECT 0.1040 68.6030 30.2580 68.6510 ;
        RECT 0.1040 69.6830 30.2580 69.7310 ;
        RECT 0.1040 70.7630 30.2580 70.8110 ;
        RECT 0.1040 71.8430 30.2580 71.8910 ;
        RECT 0.1040 72.9230 30.2580 72.9710 ;
        RECT 0.1040 74.0030 30.2580 74.0510 ;
        RECT 0.1040 75.0830 30.2580 75.1310 ;
        RECT 0.1040 76.1630 30.2580 76.2110 ;
        RECT 0.1040 77.2430 30.2580 77.2910 ;
      LAYER M3  ;
        RECT 30.1820 0.2165 30.2000 1.3765 ;
        RECT 16.2500 0.2165 16.2680 1.3765 ;
        RECT 15.4850 0.2530 15.5210 1.3675 ;
        RECT 15.2600 0.2530 15.2870 1.3675 ;
        RECT 14.0900 0.2165 14.1080 1.3765 ;
        RECT 0.1580 0.2165 0.1760 1.3765 ;
        RECT 30.1820 1.2965 30.2000 2.4565 ;
        RECT 16.2500 1.2965 16.2680 2.4565 ;
        RECT 15.4850 1.3330 15.5210 2.4475 ;
        RECT 15.2600 1.3330 15.2870 2.4475 ;
        RECT 14.0900 1.2965 14.1080 2.4565 ;
        RECT 0.1580 1.2965 0.1760 2.4565 ;
        RECT 30.1820 2.3765 30.2000 3.5365 ;
        RECT 16.2500 2.3765 16.2680 3.5365 ;
        RECT 15.4850 2.4130 15.5210 3.5275 ;
        RECT 15.2600 2.4130 15.2870 3.5275 ;
        RECT 14.0900 2.3765 14.1080 3.5365 ;
        RECT 0.1580 2.3765 0.1760 3.5365 ;
        RECT 30.1820 3.4565 30.2000 4.6165 ;
        RECT 16.2500 3.4565 16.2680 4.6165 ;
        RECT 15.4850 3.4930 15.5210 4.6075 ;
        RECT 15.2600 3.4930 15.2870 4.6075 ;
        RECT 14.0900 3.4565 14.1080 4.6165 ;
        RECT 0.1580 3.4565 0.1760 4.6165 ;
        RECT 30.1820 4.5365 30.2000 5.6965 ;
        RECT 16.2500 4.5365 16.2680 5.6965 ;
        RECT 15.4850 4.5730 15.5210 5.6875 ;
        RECT 15.2600 4.5730 15.2870 5.6875 ;
        RECT 14.0900 4.5365 14.1080 5.6965 ;
        RECT 0.1580 4.5365 0.1760 5.6965 ;
        RECT 30.1820 5.6165 30.2000 6.7765 ;
        RECT 16.2500 5.6165 16.2680 6.7765 ;
        RECT 15.4850 5.6530 15.5210 6.7675 ;
        RECT 15.2600 5.6530 15.2870 6.7675 ;
        RECT 14.0900 5.6165 14.1080 6.7765 ;
        RECT 0.1580 5.6165 0.1760 6.7765 ;
        RECT 30.1820 6.6965 30.2000 7.8565 ;
        RECT 16.2500 6.6965 16.2680 7.8565 ;
        RECT 15.4850 6.7330 15.5210 7.8475 ;
        RECT 15.2600 6.7330 15.2870 7.8475 ;
        RECT 14.0900 6.6965 14.1080 7.8565 ;
        RECT 0.1580 6.6965 0.1760 7.8565 ;
        RECT 30.1820 7.7765 30.2000 8.9365 ;
        RECT 16.2500 7.7765 16.2680 8.9365 ;
        RECT 15.4850 7.8130 15.5210 8.9275 ;
        RECT 15.2600 7.8130 15.2870 8.9275 ;
        RECT 14.0900 7.7765 14.1080 8.9365 ;
        RECT 0.1580 7.7765 0.1760 8.9365 ;
        RECT 30.1820 8.8565 30.2000 10.0165 ;
        RECT 16.2500 8.8565 16.2680 10.0165 ;
        RECT 15.4850 8.8930 15.5210 10.0075 ;
        RECT 15.2600 8.8930 15.2870 10.0075 ;
        RECT 14.0900 8.8565 14.1080 10.0165 ;
        RECT 0.1580 8.8565 0.1760 10.0165 ;
        RECT 30.1820 9.9365 30.2000 11.0965 ;
        RECT 16.2500 9.9365 16.2680 11.0965 ;
        RECT 15.4850 9.9730 15.5210 11.0875 ;
        RECT 15.2600 9.9730 15.2870 11.0875 ;
        RECT 14.0900 9.9365 14.1080 11.0965 ;
        RECT 0.1580 9.9365 0.1760 11.0965 ;
        RECT 30.1820 11.0165 30.2000 12.1765 ;
        RECT 16.2500 11.0165 16.2680 12.1765 ;
        RECT 15.4850 11.0530 15.5210 12.1675 ;
        RECT 15.2600 11.0530 15.2870 12.1675 ;
        RECT 14.0900 11.0165 14.1080 12.1765 ;
        RECT 0.1580 11.0165 0.1760 12.1765 ;
        RECT 30.1820 12.0965 30.2000 13.2565 ;
        RECT 16.2500 12.0965 16.2680 13.2565 ;
        RECT 15.4850 12.1330 15.5210 13.2475 ;
        RECT 15.2600 12.1330 15.2870 13.2475 ;
        RECT 14.0900 12.0965 14.1080 13.2565 ;
        RECT 0.1580 12.0965 0.1760 13.2565 ;
        RECT 30.1820 13.1765 30.2000 14.3365 ;
        RECT 16.2500 13.1765 16.2680 14.3365 ;
        RECT 15.4850 13.2130 15.5210 14.3275 ;
        RECT 15.2600 13.2130 15.2870 14.3275 ;
        RECT 14.0900 13.1765 14.1080 14.3365 ;
        RECT 0.1580 13.1765 0.1760 14.3365 ;
        RECT 30.1820 14.2565 30.2000 15.4165 ;
        RECT 16.2500 14.2565 16.2680 15.4165 ;
        RECT 15.4850 14.2930 15.5210 15.4075 ;
        RECT 15.2600 14.2930 15.2870 15.4075 ;
        RECT 14.0900 14.2565 14.1080 15.4165 ;
        RECT 0.1580 14.2565 0.1760 15.4165 ;
        RECT 30.1820 15.3365 30.2000 16.4965 ;
        RECT 16.2500 15.3365 16.2680 16.4965 ;
        RECT 15.4850 15.3730 15.5210 16.4875 ;
        RECT 15.2600 15.3730 15.2870 16.4875 ;
        RECT 14.0900 15.3365 14.1080 16.4965 ;
        RECT 0.1580 15.3365 0.1760 16.4965 ;
        RECT 30.1820 16.4165 30.2000 17.5765 ;
        RECT 16.2500 16.4165 16.2680 17.5765 ;
        RECT 15.4850 16.4530 15.5210 17.5675 ;
        RECT 15.2600 16.4530 15.2870 17.5675 ;
        RECT 14.0900 16.4165 14.1080 17.5765 ;
        RECT 0.1580 16.4165 0.1760 17.5765 ;
        RECT 30.1820 17.4965 30.2000 18.6565 ;
        RECT 16.2500 17.4965 16.2680 18.6565 ;
        RECT 15.4850 17.5330 15.5210 18.6475 ;
        RECT 15.2600 17.5330 15.2870 18.6475 ;
        RECT 14.0900 17.4965 14.1080 18.6565 ;
        RECT 0.1580 17.4965 0.1760 18.6565 ;
        RECT 30.1820 18.5765 30.2000 19.7365 ;
        RECT 16.2500 18.5765 16.2680 19.7365 ;
        RECT 15.4850 18.6130 15.5210 19.7275 ;
        RECT 15.2600 18.6130 15.2870 19.7275 ;
        RECT 14.0900 18.5765 14.1080 19.7365 ;
        RECT 0.1580 18.5765 0.1760 19.7365 ;
        RECT 30.1820 19.6565 30.2000 20.8165 ;
        RECT 16.2500 19.6565 16.2680 20.8165 ;
        RECT 15.4850 19.6930 15.5210 20.8075 ;
        RECT 15.2600 19.6930 15.2870 20.8075 ;
        RECT 14.0900 19.6565 14.1080 20.8165 ;
        RECT 0.1580 19.6565 0.1760 20.8165 ;
        RECT 30.1820 20.7365 30.2000 21.8965 ;
        RECT 16.2500 20.7365 16.2680 21.8965 ;
        RECT 15.4850 20.7730 15.5210 21.8875 ;
        RECT 15.2600 20.7730 15.2870 21.8875 ;
        RECT 14.0900 20.7365 14.1080 21.8965 ;
        RECT 0.1580 20.7365 0.1760 21.8965 ;
        RECT 30.1820 21.8165 30.2000 22.9765 ;
        RECT 16.2500 21.8165 16.2680 22.9765 ;
        RECT 15.4850 21.8530 15.5210 22.9675 ;
        RECT 15.2600 21.8530 15.2870 22.9675 ;
        RECT 14.0900 21.8165 14.1080 22.9765 ;
        RECT 0.1580 21.8165 0.1760 22.9765 ;
        RECT 30.1820 22.8965 30.2000 24.0565 ;
        RECT 16.2500 22.8965 16.2680 24.0565 ;
        RECT 15.4850 22.9330 15.5210 24.0475 ;
        RECT 15.2600 22.9330 15.2870 24.0475 ;
        RECT 14.0900 22.8965 14.1080 24.0565 ;
        RECT 0.1580 22.8965 0.1760 24.0565 ;
        RECT 30.1820 23.9765 30.2000 25.1365 ;
        RECT 16.2500 23.9765 16.2680 25.1365 ;
        RECT 15.4850 24.0130 15.5210 25.1275 ;
        RECT 15.2600 24.0130 15.2870 25.1275 ;
        RECT 14.0900 23.9765 14.1080 25.1365 ;
        RECT 0.1580 23.9765 0.1760 25.1365 ;
        RECT 30.1820 25.0565 30.2000 26.2165 ;
        RECT 16.2500 25.0565 16.2680 26.2165 ;
        RECT 15.4850 25.0930 15.5210 26.2075 ;
        RECT 15.2600 25.0930 15.2870 26.2075 ;
        RECT 14.0900 25.0565 14.1080 26.2165 ;
        RECT 0.1580 25.0565 0.1760 26.2165 ;
        RECT 30.1820 26.1365 30.2000 27.2965 ;
        RECT 16.2500 26.1365 16.2680 27.2965 ;
        RECT 15.4850 26.1730 15.5210 27.2875 ;
        RECT 15.2600 26.1730 15.2870 27.2875 ;
        RECT 14.0900 26.1365 14.1080 27.2965 ;
        RECT 0.1580 26.1365 0.1760 27.2965 ;
        RECT 30.1820 27.2165 30.2000 28.3765 ;
        RECT 16.2500 27.2165 16.2680 28.3765 ;
        RECT 15.4850 27.2530 15.5210 28.3675 ;
        RECT 15.2600 27.2530 15.2870 28.3675 ;
        RECT 14.0900 27.2165 14.1080 28.3765 ;
        RECT 0.1580 27.2165 0.1760 28.3765 ;
        RECT 30.1820 28.2965 30.2000 29.4565 ;
        RECT 16.2500 28.2965 16.2680 29.4565 ;
        RECT 15.4850 28.3330 15.5210 29.4475 ;
        RECT 15.2600 28.3330 15.2870 29.4475 ;
        RECT 14.0900 28.2965 14.1080 29.4565 ;
        RECT 0.1580 28.2965 0.1760 29.4565 ;
        RECT 30.1820 29.3765 30.2000 30.5365 ;
        RECT 16.2500 29.3765 16.2680 30.5365 ;
        RECT 15.4850 29.4130 15.5210 30.5275 ;
        RECT 15.2600 29.4130 15.2870 30.5275 ;
        RECT 14.0900 29.3765 14.1080 30.5365 ;
        RECT 0.1580 29.3765 0.1760 30.5365 ;
        RECT 30.1820 30.4565 30.2000 31.6165 ;
        RECT 16.2500 30.4565 16.2680 31.6165 ;
        RECT 15.4850 30.4930 15.5210 31.6075 ;
        RECT 15.2600 30.4930 15.2870 31.6075 ;
        RECT 14.0900 30.4565 14.1080 31.6165 ;
        RECT 0.1580 30.4565 0.1760 31.6165 ;
        RECT 30.1820 31.5365 30.2000 32.6965 ;
        RECT 16.2500 31.5365 16.2680 32.6965 ;
        RECT 15.4850 31.5730 15.5210 32.6875 ;
        RECT 15.2600 31.5730 15.2870 32.6875 ;
        RECT 14.0900 31.5365 14.1080 32.6965 ;
        RECT 0.1580 31.5365 0.1760 32.6965 ;
        RECT 30.1820 32.6165 30.2000 33.7765 ;
        RECT 16.2500 32.6165 16.2680 33.7765 ;
        RECT 15.4850 32.6530 15.5210 33.7675 ;
        RECT 15.2600 32.6530 15.2870 33.7675 ;
        RECT 14.0900 32.6165 14.1080 33.7765 ;
        RECT 0.1580 32.6165 0.1760 33.7765 ;
        RECT 30.1820 33.6965 30.2000 34.8565 ;
        RECT 16.2500 33.6965 16.2680 34.8565 ;
        RECT 15.4850 33.7330 15.5210 34.8475 ;
        RECT 15.2600 33.7330 15.2870 34.8475 ;
        RECT 14.0900 33.6965 14.1080 34.8565 ;
        RECT 0.1580 33.6965 0.1760 34.8565 ;
        RECT 16.2450 34.8270 16.2630 43.0340 ;
        RECT 15.2910 35.0505 15.5250 42.7335 ;
        RECT 14.0850 34.8270 14.1030 44.7085 ;
        RECT 30.1820 42.9035 30.2000 44.0635 ;
        RECT 16.2500 42.9035 16.2680 44.0635 ;
        RECT 15.4850 42.9400 15.5210 44.0545 ;
        RECT 15.2600 42.9400 15.2870 44.0545 ;
        RECT 14.0900 42.9035 14.1080 44.0635 ;
        RECT 0.1580 42.9035 0.1760 44.0635 ;
        RECT 30.1820 43.9835 30.2000 45.1435 ;
        RECT 16.2500 43.9835 16.2680 45.1435 ;
        RECT 15.4850 44.0200 15.5210 45.1345 ;
        RECT 15.2600 44.0200 15.2870 45.1345 ;
        RECT 14.0900 43.9835 14.1080 45.1435 ;
        RECT 0.1580 43.9835 0.1760 45.1435 ;
        RECT 30.1820 45.0635 30.2000 46.2235 ;
        RECT 16.2500 45.0635 16.2680 46.2235 ;
        RECT 15.4850 45.1000 15.5210 46.2145 ;
        RECT 15.2600 45.1000 15.2870 46.2145 ;
        RECT 14.0900 45.0635 14.1080 46.2235 ;
        RECT 0.1580 45.0635 0.1760 46.2235 ;
        RECT 30.1820 46.1435 30.2000 47.3035 ;
        RECT 16.2500 46.1435 16.2680 47.3035 ;
        RECT 15.4850 46.1800 15.5210 47.2945 ;
        RECT 15.2600 46.1800 15.2870 47.2945 ;
        RECT 14.0900 46.1435 14.1080 47.3035 ;
        RECT 0.1580 46.1435 0.1760 47.3035 ;
        RECT 30.1820 47.2235 30.2000 48.3835 ;
        RECT 16.2500 47.2235 16.2680 48.3835 ;
        RECT 15.4850 47.2600 15.5210 48.3745 ;
        RECT 15.2600 47.2600 15.2870 48.3745 ;
        RECT 14.0900 47.2235 14.1080 48.3835 ;
        RECT 0.1580 47.2235 0.1760 48.3835 ;
        RECT 30.1820 48.3035 30.2000 49.4635 ;
        RECT 16.2500 48.3035 16.2680 49.4635 ;
        RECT 15.4850 48.3400 15.5210 49.4545 ;
        RECT 15.2600 48.3400 15.2870 49.4545 ;
        RECT 14.0900 48.3035 14.1080 49.4635 ;
        RECT 0.1580 48.3035 0.1760 49.4635 ;
        RECT 30.1820 49.3835 30.2000 50.5435 ;
        RECT 16.2500 49.3835 16.2680 50.5435 ;
        RECT 15.4850 49.4200 15.5210 50.5345 ;
        RECT 15.2600 49.4200 15.2870 50.5345 ;
        RECT 14.0900 49.3835 14.1080 50.5435 ;
        RECT 0.1580 49.3835 0.1760 50.5435 ;
        RECT 30.1820 50.4635 30.2000 51.6235 ;
        RECT 16.2500 50.4635 16.2680 51.6235 ;
        RECT 15.4850 50.5000 15.5210 51.6145 ;
        RECT 15.2600 50.5000 15.2870 51.6145 ;
        RECT 14.0900 50.4635 14.1080 51.6235 ;
        RECT 0.1580 50.4635 0.1760 51.6235 ;
        RECT 30.1820 51.5435 30.2000 52.7035 ;
        RECT 16.2500 51.5435 16.2680 52.7035 ;
        RECT 15.4850 51.5800 15.5210 52.6945 ;
        RECT 15.2600 51.5800 15.2870 52.6945 ;
        RECT 14.0900 51.5435 14.1080 52.7035 ;
        RECT 0.1580 51.5435 0.1760 52.7035 ;
        RECT 30.1820 52.6235 30.2000 53.7835 ;
        RECT 16.2500 52.6235 16.2680 53.7835 ;
        RECT 15.4850 52.6600 15.5210 53.7745 ;
        RECT 15.2600 52.6600 15.2870 53.7745 ;
        RECT 14.0900 52.6235 14.1080 53.7835 ;
        RECT 0.1580 52.6235 0.1760 53.7835 ;
        RECT 30.1820 53.7035 30.2000 54.8635 ;
        RECT 16.2500 53.7035 16.2680 54.8635 ;
        RECT 15.4850 53.7400 15.5210 54.8545 ;
        RECT 15.2600 53.7400 15.2870 54.8545 ;
        RECT 14.0900 53.7035 14.1080 54.8635 ;
        RECT 0.1580 53.7035 0.1760 54.8635 ;
        RECT 30.1820 54.7835 30.2000 55.9435 ;
        RECT 16.2500 54.7835 16.2680 55.9435 ;
        RECT 15.4850 54.8200 15.5210 55.9345 ;
        RECT 15.2600 54.8200 15.2870 55.9345 ;
        RECT 14.0900 54.7835 14.1080 55.9435 ;
        RECT 0.1580 54.7835 0.1760 55.9435 ;
        RECT 30.1820 55.8635 30.2000 57.0235 ;
        RECT 16.2500 55.8635 16.2680 57.0235 ;
        RECT 15.4850 55.9000 15.5210 57.0145 ;
        RECT 15.2600 55.9000 15.2870 57.0145 ;
        RECT 14.0900 55.8635 14.1080 57.0235 ;
        RECT 0.1580 55.8635 0.1760 57.0235 ;
        RECT 30.1820 56.9435 30.2000 58.1035 ;
        RECT 16.2500 56.9435 16.2680 58.1035 ;
        RECT 15.4850 56.9800 15.5210 58.0945 ;
        RECT 15.2600 56.9800 15.2870 58.0945 ;
        RECT 14.0900 56.9435 14.1080 58.1035 ;
        RECT 0.1580 56.9435 0.1760 58.1035 ;
        RECT 30.1820 58.0235 30.2000 59.1835 ;
        RECT 16.2500 58.0235 16.2680 59.1835 ;
        RECT 15.4850 58.0600 15.5210 59.1745 ;
        RECT 15.2600 58.0600 15.2870 59.1745 ;
        RECT 14.0900 58.0235 14.1080 59.1835 ;
        RECT 0.1580 58.0235 0.1760 59.1835 ;
        RECT 30.1820 59.1035 30.2000 60.2635 ;
        RECT 16.2500 59.1035 16.2680 60.2635 ;
        RECT 15.4850 59.1400 15.5210 60.2545 ;
        RECT 15.2600 59.1400 15.2870 60.2545 ;
        RECT 14.0900 59.1035 14.1080 60.2635 ;
        RECT 0.1580 59.1035 0.1760 60.2635 ;
        RECT 30.1820 60.1835 30.2000 61.3435 ;
        RECT 16.2500 60.1835 16.2680 61.3435 ;
        RECT 15.4850 60.2200 15.5210 61.3345 ;
        RECT 15.2600 60.2200 15.2870 61.3345 ;
        RECT 14.0900 60.1835 14.1080 61.3435 ;
        RECT 0.1580 60.1835 0.1760 61.3435 ;
        RECT 30.1820 61.2635 30.2000 62.4235 ;
        RECT 16.2500 61.2635 16.2680 62.4235 ;
        RECT 15.4850 61.3000 15.5210 62.4145 ;
        RECT 15.2600 61.3000 15.2870 62.4145 ;
        RECT 14.0900 61.2635 14.1080 62.4235 ;
        RECT 0.1580 61.2635 0.1760 62.4235 ;
        RECT 30.1820 62.3435 30.2000 63.5035 ;
        RECT 16.2500 62.3435 16.2680 63.5035 ;
        RECT 15.4850 62.3800 15.5210 63.4945 ;
        RECT 15.2600 62.3800 15.2870 63.4945 ;
        RECT 14.0900 62.3435 14.1080 63.5035 ;
        RECT 0.1580 62.3435 0.1760 63.5035 ;
        RECT 30.1820 63.4235 30.2000 64.5835 ;
        RECT 16.2500 63.4235 16.2680 64.5835 ;
        RECT 15.4850 63.4600 15.5210 64.5745 ;
        RECT 15.2600 63.4600 15.2870 64.5745 ;
        RECT 14.0900 63.4235 14.1080 64.5835 ;
        RECT 0.1580 63.4235 0.1760 64.5835 ;
        RECT 30.1820 64.5035 30.2000 65.6635 ;
        RECT 16.2500 64.5035 16.2680 65.6635 ;
        RECT 15.4850 64.5400 15.5210 65.6545 ;
        RECT 15.2600 64.5400 15.2870 65.6545 ;
        RECT 14.0900 64.5035 14.1080 65.6635 ;
        RECT 0.1580 64.5035 0.1760 65.6635 ;
        RECT 30.1820 65.5835 30.2000 66.7435 ;
        RECT 16.2500 65.5835 16.2680 66.7435 ;
        RECT 15.4850 65.6200 15.5210 66.7345 ;
        RECT 15.2600 65.6200 15.2870 66.7345 ;
        RECT 14.0900 65.5835 14.1080 66.7435 ;
        RECT 0.1580 65.5835 0.1760 66.7435 ;
        RECT 30.1820 66.6635 30.2000 67.8235 ;
        RECT 16.2500 66.6635 16.2680 67.8235 ;
        RECT 15.4850 66.7000 15.5210 67.8145 ;
        RECT 15.2600 66.7000 15.2870 67.8145 ;
        RECT 14.0900 66.6635 14.1080 67.8235 ;
        RECT 0.1580 66.6635 0.1760 67.8235 ;
        RECT 30.1820 67.7435 30.2000 68.9035 ;
        RECT 16.2500 67.7435 16.2680 68.9035 ;
        RECT 15.4850 67.7800 15.5210 68.8945 ;
        RECT 15.2600 67.7800 15.2870 68.8945 ;
        RECT 14.0900 67.7435 14.1080 68.9035 ;
        RECT 0.1580 67.7435 0.1760 68.9035 ;
        RECT 30.1820 68.8235 30.2000 69.9835 ;
        RECT 16.2500 68.8235 16.2680 69.9835 ;
        RECT 15.4850 68.8600 15.5210 69.9745 ;
        RECT 15.2600 68.8600 15.2870 69.9745 ;
        RECT 14.0900 68.8235 14.1080 69.9835 ;
        RECT 0.1580 68.8235 0.1760 69.9835 ;
        RECT 30.1820 69.9035 30.2000 71.0635 ;
        RECT 16.2500 69.9035 16.2680 71.0635 ;
        RECT 15.4850 69.9400 15.5210 71.0545 ;
        RECT 15.2600 69.9400 15.2870 71.0545 ;
        RECT 14.0900 69.9035 14.1080 71.0635 ;
        RECT 0.1580 69.9035 0.1760 71.0635 ;
        RECT 30.1820 70.9835 30.2000 72.1435 ;
        RECT 16.2500 70.9835 16.2680 72.1435 ;
        RECT 15.4850 71.0200 15.5210 72.1345 ;
        RECT 15.2600 71.0200 15.2870 72.1345 ;
        RECT 14.0900 70.9835 14.1080 72.1435 ;
        RECT 0.1580 70.9835 0.1760 72.1435 ;
        RECT 30.1820 72.0635 30.2000 73.2235 ;
        RECT 16.2500 72.0635 16.2680 73.2235 ;
        RECT 15.4850 72.1000 15.5210 73.2145 ;
        RECT 15.2600 72.1000 15.2870 73.2145 ;
        RECT 14.0900 72.0635 14.1080 73.2235 ;
        RECT 0.1580 72.0635 0.1760 73.2235 ;
        RECT 30.1820 73.1435 30.2000 74.3035 ;
        RECT 16.2500 73.1435 16.2680 74.3035 ;
        RECT 15.4850 73.1800 15.5210 74.2945 ;
        RECT 15.2600 73.1800 15.2870 74.2945 ;
        RECT 14.0900 73.1435 14.1080 74.3035 ;
        RECT 0.1580 73.1435 0.1760 74.3035 ;
        RECT 30.1820 74.2235 30.2000 75.3835 ;
        RECT 16.2500 74.2235 16.2680 75.3835 ;
        RECT 15.4850 74.2600 15.5210 75.3745 ;
        RECT 15.2600 74.2600 15.2870 75.3745 ;
        RECT 14.0900 74.2235 14.1080 75.3835 ;
        RECT 0.1580 74.2235 0.1760 75.3835 ;
        RECT 30.1820 75.3035 30.2000 76.4635 ;
        RECT 16.2500 75.3035 16.2680 76.4635 ;
        RECT 15.4850 75.3400 15.5210 76.4545 ;
        RECT 15.2600 75.3400 15.2870 76.4545 ;
        RECT 14.0900 75.3035 14.1080 76.4635 ;
        RECT 0.1580 75.3035 0.1760 76.4635 ;
        RECT 30.1820 76.3835 30.2000 77.5435 ;
        RECT 16.2500 76.3835 16.2680 77.5435 ;
        RECT 15.4850 76.4200 15.5210 77.5345 ;
        RECT 15.2600 76.4200 15.2870 77.5345 ;
        RECT 14.0900 76.3835 14.1080 77.5435 ;
        RECT 0.1580 76.3835 0.1760 77.5435 ;
      LAYER V3  ;
        RECT 0.1580 1.0760 0.1760 1.1240 ;
        RECT 14.0900 1.0760 14.1080 1.1240 ;
        RECT 15.2600 1.0760 15.2870 1.1240 ;
        RECT 15.4850 1.0760 15.5210 1.1240 ;
        RECT 16.2500 1.0760 16.2680 1.1240 ;
        RECT 30.1820 1.0760 30.2000 1.1240 ;
        RECT 0.1580 2.1560 0.1760 2.2040 ;
        RECT 14.0900 2.1560 14.1080 2.2040 ;
        RECT 15.2600 2.1560 15.2870 2.2040 ;
        RECT 15.4850 2.1560 15.5210 2.2040 ;
        RECT 16.2500 2.1560 16.2680 2.2040 ;
        RECT 30.1820 2.1560 30.2000 2.2040 ;
        RECT 0.1580 3.2360 0.1760 3.2840 ;
        RECT 14.0900 3.2360 14.1080 3.2840 ;
        RECT 15.2600 3.2360 15.2870 3.2840 ;
        RECT 15.4850 3.2360 15.5210 3.2840 ;
        RECT 16.2500 3.2360 16.2680 3.2840 ;
        RECT 30.1820 3.2360 30.2000 3.2840 ;
        RECT 0.1580 4.3160 0.1760 4.3640 ;
        RECT 14.0900 4.3160 14.1080 4.3640 ;
        RECT 15.2600 4.3160 15.2870 4.3640 ;
        RECT 15.4850 4.3160 15.5210 4.3640 ;
        RECT 16.2500 4.3160 16.2680 4.3640 ;
        RECT 30.1820 4.3160 30.2000 4.3640 ;
        RECT 0.1580 5.3960 0.1760 5.4440 ;
        RECT 14.0900 5.3960 14.1080 5.4440 ;
        RECT 15.2600 5.3960 15.2870 5.4440 ;
        RECT 15.4850 5.3960 15.5210 5.4440 ;
        RECT 16.2500 5.3960 16.2680 5.4440 ;
        RECT 30.1820 5.3960 30.2000 5.4440 ;
        RECT 0.1580 6.4760 0.1760 6.5240 ;
        RECT 14.0900 6.4760 14.1080 6.5240 ;
        RECT 15.2600 6.4760 15.2870 6.5240 ;
        RECT 15.4850 6.4760 15.5210 6.5240 ;
        RECT 16.2500 6.4760 16.2680 6.5240 ;
        RECT 30.1820 6.4760 30.2000 6.5240 ;
        RECT 0.1580 7.5560 0.1760 7.6040 ;
        RECT 14.0900 7.5560 14.1080 7.6040 ;
        RECT 15.2600 7.5560 15.2870 7.6040 ;
        RECT 15.4850 7.5560 15.5210 7.6040 ;
        RECT 16.2500 7.5560 16.2680 7.6040 ;
        RECT 30.1820 7.5560 30.2000 7.6040 ;
        RECT 0.1580 8.6360 0.1760 8.6840 ;
        RECT 14.0900 8.6360 14.1080 8.6840 ;
        RECT 15.2600 8.6360 15.2870 8.6840 ;
        RECT 15.4850 8.6360 15.5210 8.6840 ;
        RECT 16.2500 8.6360 16.2680 8.6840 ;
        RECT 30.1820 8.6360 30.2000 8.6840 ;
        RECT 0.1580 9.7160 0.1760 9.7640 ;
        RECT 14.0900 9.7160 14.1080 9.7640 ;
        RECT 15.2600 9.7160 15.2870 9.7640 ;
        RECT 15.4850 9.7160 15.5210 9.7640 ;
        RECT 16.2500 9.7160 16.2680 9.7640 ;
        RECT 30.1820 9.7160 30.2000 9.7640 ;
        RECT 0.1580 10.7960 0.1760 10.8440 ;
        RECT 14.0900 10.7960 14.1080 10.8440 ;
        RECT 15.2600 10.7960 15.2870 10.8440 ;
        RECT 15.4850 10.7960 15.5210 10.8440 ;
        RECT 16.2500 10.7960 16.2680 10.8440 ;
        RECT 30.1820 10.7960 30.2000 10.8440 ;
        RECT 0.1580 11.8760 0.1760 11.9240 ;
        RECT 14.0900 11.8760 14.1080 11.9240 ;
        RECT 15.2600 11.8760 15.2870 11.9240 ;
        RECT 15.4850 11.8760 15.5210 11.9240 ;
        RECT 16.2500 11.8760 16.2680 11.9240 ;
        RECT 30.1820 11.8760 30.2000 11.9240 ;
        RECT 0.1580 12.9560 0.1760 13.0040 ;
        RECT 14.0900 12.9560 14.1080 13.0040 ;
        RECT 15.2600 12.9560 15.2870 13.0040 ;
        RECT 15.4850 12.9560 15.5210 13.0040 ;
        RECT 16.2500 12.9560 16.2680 13.0040 ;
        RECT 30.1820 12.9560 30.2000 13.0040 ;
        RECT 0.1580 14.0360 0.1760 14.0840 ;
        RECT 14.0900 14.0360 14.1080 14.0840 ;
        RECT 15.2600 14.0360 15.2870 14.0840 ;
        RECT 15.4850 14.0360 15.5210 14.0840 ;
        RECT 16.2500 14.0360 16.2680 14.0840 ;
        RECT 30.1820 14.0360 30.2000 14.0840 ;
        RECT 0.1580 15.1160 0.1760 15.1640 ;
        RECT 14.0900 15.1160 14.1080 15.1640 ;
        RECT 15.2600 15.1160 15.2870 15.1640 ;
        RECT 15.4850 15.1160 15.5210 15.1640 ;
        RECT 16.2500 15.1160 16.2680 15.1640 ;
        RECT 30.1820 15.1160 30.2000 15.1640 ;
        RECT 0.1580 16.1960 0.1760 16.2440 ;
        RECT 14.0900 16.1960 14.1080 16.2440 ;
        RECT 15.2600 16.1960 15.2870 16.2440 ;
        RECT 15.4850 16.1960 15.5210 16.2440 ;
        RECT 16.2500 16.1960 16.2680 16.2440 ;
        RECT 30.1820 16.1960 30.2000 16.2440 ;
        RECT 0.1580 17.2760 0.1760 17.3240 ;
        RECT 14.0900 17.2760 14.1080 17.3240 ;
        RECT 15.2600 17.2760 15.2870 17.3240 ;
        RECT 15.4850 17.2760 15.5210 17.3240 ;
        RECT 16.2500 17.2760 16.2680 17.3240 ;
        RECT 30.1820 17.2760 30.2000 17.3240 ;
        RECT 0.1580 18.3560 0.1760 18.4040 ;
        RECT 14.0900 18.3560 14.1080 18.4040 ;
        RECT 15.2600 18.3560 15.2870 18.4040 ;
        RECT 15.4850 18.3560 15.5210 18.4040 ;
        RECT 16.2500 18.3560 16.2680 18.4040 ;
        RECT 30.1820 18.3560 30.2000 18.4040 ;
        RECT 0.1580 19.4360 0.1760 19.4840 ;
        RECT 14.0900 19.4360 14.1080 19.4840 ;
        RECT 15.2600 19.4360 15.2870 19.4840 ;
        RECT 15.4850 19.4360 15.5210 19.4840 ;
        RECT 16.2500 19.4360 16.2680 19.4840 ;
        RECT 30.1820 19.4360 30.2000 19.4840 ;
        RECT 0.1580 20.5160 0.1760 20.5640 ;
        RECT 14.0900 20.5160 14.1080 20.5640 ;
        RECT 15.2600 20.5160 15.2870 20.5640 ;
        RECT 15.4850 20.5160 15.5210 20.5640 ;
        RECT 16.2500 20.5160 16.2680 20.5640 ;
        RECT 30.1820 20.5160 30.2000 20.5640 ;
        RECT 0.1580 21.5960 0.1760 21.6440 ;
        RECT 14.0900 21.5960 14.1080 21.6440 ;
        RECT 15.2600 21.5960 15.2870 21.6440 ;
        RECT 15.4850 21.5960 15.5210 21.6440 ;
        RECT 16.2500 21.5960 16.2680 21.6440 ;
        RECT 30.1820 21.5960 30.2000 21.6440 ;
        RECT 0.1580 22.6760 0.1760 22.7240 ;
        RECT 14.0900 22.6760 14.1080 22.7240 ;
        RECT 15.2600 22.6760 15.2870 22.7240 ;
        RECT 15.4850 22.6760 15.5210 22.7240 ;
        RECT 16.2500 22.6760 16.2680 22.7240 ;
        RECT 30.1820 22.6760 30.2000 22.7240 ;
        RECT 0.1580 23.7560 0.1760 23.8040 ;
        RECT 14.0900 23.7560 14.1080 23.8040 ;
        RECT 15.2600 23.7560 15.2870 23.8040 ;
        RECT 15.4850 23.7560 15.5210 23.8040 ;
        RECT 16.2500 23.7560 16.2680 23.8040 ;
        RECT 30.1820 23.7560 30.2000 23.8040 ;
        RECT 0.1580 24.8360 0.1760 24.8840 ;
        RECT 14.0900 24.8360 14.1080 24.8840 ;
        RECT 15.2600 24.8360 15.2870 24.8840 ;
        RECT 15.4850 24.8360 15.5210 24.8840 ;
        RECT 16.2500 24.8360 16.2680 24.8840 ;
        RECT 30.1820 24.8360 30.2000 24.8840 ;
        RECT 0.1580 25.9160 0.1760 25.9640 ;
        RECT 14.0900 25.9160 14.1080 25.9640 ;
        RECT 15.2600 25.9160 15.2870 25.9640 ;
        RECT 15.4850 25.9160 15.5210 25.9640 ;
        RECT 16.2500 25.9160 16.2680 25.9640 ;
        RECT 30.1820 25.9160 30.2000 25.9640 ;
        RECT 0.1580 26.9960 0.1760 27.0440 ;
        RECT 14.0900 26.9960 14.1080 27.0440 ;
        RECT 15.2600 26.9960 15.2870 27.0440 ;
        RECT 15.4850 26.9960 15.5210 27.0440 ;
        RECT 16.2500 26.9960 16.2680 27.0440 ;
        RECT 30.1820 26.9960 30.2000 27.0440 ;
        RECT 0.1580 28.0760 0.1760 28.1240 ;
        RECT 14.0900 28.0760 14.1080 28.1240 ;
        RECT 15.2600 28.0760 15.2870 28.1240 ;
        RECT 15.4850 28.0760 15.5210 28.1240 ;
        RECT 16.2500 28.0760 16.2680 28.1240 ;
        RECT 30.1820 28.0760 30.2000 28.1240 ;
        RECT 0.1580 29.1560 0.1760 29.2040 ;
        RECT 14.0900 29.1560 14.1080 29.2040 ;
        RECT 15.2600 29.1560 15.2870 29.2040 ;
        RECT 15.4850 29.1560 15.5210 29.2040 ;
        RECT 16.2500 29.1560 16.2680 29.2040 ;
        RECT 30.1820 29.1560 30.2000 29.2040 ;
        RECT 0.1580 30.2360 0.1760 30.2840 ;
        RECT 14.0900 30.2360 14.1080 30.2840 ;
        RECT 15.2600 30.2360 15.2870 30.2840 ;
        RECT 15.4850 30.2360 15.5210 30.2840 ;
        RECT 16.2500 30.2360 16.2680 30.2840 ;
        RECT 30.1820 30.2360 30.2000 30.2840 ;
        RECT 0.1580 31.3160 0.1760 31.3640 ;
        RECT 14.0900 31.3160 14.1080 31.3640 ;
        RECT 15.2600 31.3160 15.2870 31.3640 ;
        RECT 15.4850 31.3160 15.5210 31.3640 ;
        RECT 16.2500 31.3160 16.2680 31.3640 ;
        RECT 30.1820 31.3160 30.2000 31.3640 ;
        RECT 0.1580 32.3960 0.1760 32.4440 ;
        RECT 14.0900 32.3960 14.1080 32.4440 ;
        RECT 15.2600 32.3960 15.2870 32.4440 ;
        RECT 15.4850 32.3960 15.5210 32.4440 ;
        RECT 16.2500 32.3960 16.2680 32.4440 ;
        RECT 30.1820 32.3960 30.2000 32.4440 ;
        RECT 0.1580 33.4760 0.1760 33.5240 ;
        RECT 14.0900 33.4760 14.1080 33.5240 ;
        RECT 15.2600 33.4760 15.2870 33.5240 ;
        RECT 15.4850 33.4760 15.5210 33.5240 ;
        RECT 16.2500 33.4760 16.2680 33.5240 ;
        RECT 30.1820 33.4760 30.2000 33.5240 ;
        RECT 0.1580 34.5560 0.1760 34.6040 ;
        RECT 14.0900 34.5560 14.1080 34.6040 ;
        RECT 15.2600 34.5560 15.2870 34.6040 ;
        RECT 15.4850 34.5560 15.5210 34.6040 ;
        RECT 16.2500 34.5560 16.2680 34.6040 ;
        RECT 30.1820 34.5560 30.2000 34.6040 ;
        RECT 14.0850 35.6215 14.1030 35.8375 ;
        RECT 15.2950 41.9575 15.3130 42.1735 ;
        RECT 15.2950 38.7895 15.3130 39.0055 ;
        RECT 15.2950 35.6215 15.3130 35.8375 ;
        RECT 15.3470 41.9575 15.3650 42.1735 ;
        RECT 15.3470 38.7895 15.3650 39.0055 ;
        RECT 15.3470 35.6215 15.3650 35.8375 ;
        RECT 15.3990 41.9575 15.4170 42.1735 ;
        RECT 15.3990 38.7895 15.4170 39.0055 ;
        RECT 15.3990 35.6215 15.4170 35.8375 ;
        RECT 15.4510 41.9575 15.4690 42.1735 ;
        RECT 15.4510 38.7895 15.4690 39.0055 ;
        RECT 15.4510 35.6215 15.4690 35.8375 ;
        RECT 15.5030 41.9575 15.5210 42.1735 ;
        RECT 15.5030 38.7895 15.5210 39.0055 ;
        RECT 15.5030 35.6215 15.5210 35.8375 ;
        RECT 16.2450 35.6215 16.2630 35.8375 ;
        RECT 0.1580 43.7630 0.1760 43.8110 ;
        RECT 14.0900 43.7630 14.1080 43.8110 ;
        RECT 15.2600 43.7630 15.2870 43.8110 ;
        RECT 15.4850 43.7630 15.5210 43.8110 ;
        RECT 16.2500 43.7630 16.2680 43.8110 ;
        RECT 30.1820 43.7630 30.2000 43.8110 ;
        RECT 0.1580 44.8430 0.1760 44.8910 ;
        RECT 14.0900 44.8430 14.1080 44.8910 ;
        RECT 15.2600 44.8430 15.2870 44.8910 ;
        RECT 15.4850 44.8430 15.5210 44.8910 ;
        RECT 16.2500 44.8430 16.2680 44.8910 ;
        RECT 30.1820 44.8430 30.2000 44.8910 ;
        RECT 0.1580 45.9230 0.1760 45.9710 ;
        RECT 14.0900 45.9230 14.1080 45.9710 ;
        RECT 15.2600 45.9230 15.2870 45.9710 ;
        RECT 15.4850 45.9230 15.5210 45.9710 ;
        RECT 16.2500 45.9230 16.2680 45.9710 ;
        RECT 30.1820 45.9230 30.2000 45.9710 ;
        RECT 0.1580 47.0030 0.1760 47.0510 ;
        RECT 14.0900 47.0030 14.1080 47.0510 ;
        RECT 15.2600 47.0030 15.2870 47.0510 ;
        RECT 15.4850 47.0030 15.5210 47.0510 ;
        RECT 16.2500 47.0030 16.2680 47.0510 ;
        RECT 30.1820 47.0030 30.2000 47.0510 ;
        RECT 0.1580 48.0830 0.1760 48.1310 ;
        RECT 14.0900 48.0830 14.1080 48.1310 ;
        RECT 15.2600 48.0830 15.2870 48.1310 ;
        RECT 15.4850 48.0830 15.5210 48.1310 ;
        RECT 16.2500 48.0830 16.2680 48.1310 ;
        RECT 30.1820 48.0830 30.2000 48.1310 ;
        RECT 0.1580 49.1630 0.1760 49.2110 ;
        RECT 14.0900 49.1630 14.1080 49.2110 ;
        RECT 15.2600 49.1630 15.2870 49.2110 ;
        RECT 15.4850 49.1630 15.5210 49.2110 ;
        RECT 16.2500 49.1630 16.2680 49.2110 ;
        RECT 30.1820 49.1630 30.2000 49.2110 ;
        RECT 0.1580 50.2430 0.1760 50.2910 ;
        RECT 14.0900 50.2430 14.1080 50.2910 ;
        RECT 15.2600 50.2430 15.2870 50.2910 ;
        RECT 15.4850 50.2430 15.5210 50.2910 ;
        RECT 16.2500 50.2430 16.2680 50.2910 ;
        RECT 30.1820 50.2430 30.2000 50.2910 ;
        RECT 0.1580 51.3230 0.1760 51.3710 ;
        RECT 14.0900 51.3230 14.1080 51.3710 ;
        RECT 15.2600 51.3230 15.2870 51.3710 ;
        RECT 15.4850 51.3230 15.5210 51.3710 ;
        RECT 16.2500 51.3230 16.2680 51.3710 ;
        RECT 30.1820 51.3230 30.2000 51.3710 ;
        RECT 0.1580 52.4030 0.1760 52.4510 ;
        RECT 14.0900 52.4030 14.1080 52.4510 ;
        RECT 15.2600 52.4030 15.2870 52.4510 ;
        RECT 15.4850 52.4030 15.5210 52.4510 ;
        RECT 16.2500 52.4030 16.2680 52.4510 ;
        RECT 30.1820 52.4030 30.2000 52.4510 ;
        RECT 0.1580 53.4830 0.1760 53.5310 ;
        RECT 14.0900 53.4830 14.1080 53.5310 ;
        RECT 15.2600 53.4830 15.2870 53.5310 ;
        RECT 15.4850 53.4830 15.5210 53.5310 ;
        RECT 16.2500 53.4830 16.2680 53.5310 ;
        RECT 30.1820 53.4830 30.2000 53.5310 ;
        RECT 0.1580 54.5630 0.1760 54.6110 ;
        RECT 14.0900 54.5630 14.1080 54.6110 ;
        RECT 15.2600 54.5630 15.2870 54.6110 ;
        RECT 15.4850 54.5630 15.5210 54.6110 ;
        RECT 16.2500 54.5630 16.2680 54.6110 ;
        RECT 30.1820 54.5630 30.2000 54.6110 ;
        RECT 0.1580 55.6430 0.1760 55.6910 ;
        RECT 14.0900 55.6430 14.1080 55.6910 ;
        RECT 15.2600 55.6430 15.2870 55.6910 ;
        RECT 15.4850 55.6430 15.5210 55.6910 ;
        RECT 16.2500 55.6430 16.2680 55.6910 ;
        RECT 30.1820 55.6430 30.2000 55.6910 ;
        RECT 0.1580 56.7230 0.1760 56.7710 ;
        RECT 14.0900 56.7230 14.1080 56.7710 ;
        RECT 15.2600 56.7230 15.2870 56.7710 ;
        RECT 15.4850 56.7230 15.5210 56.7710 ;
        RECT 16.2500 56.7230 16.2680 56.7710 ;
        RECT 30.1820 56.7230 30.2000 56.7710 ;
        RECT 0.1580 57.8030 0.1760 57.8510 ;
        RECT 14.0900 57.8030 14.1080 57.8510 ;
        RECT 15.2600 57.8030 15.2870 57.8510 ;
        RECT 15.4850 57.8030 15.5210 57.8510 ;
        RECT 16.2500 57.8030 16.2680 57.8510 ;
        RECT 30.1820 57.8030 30.2000 57.8510 ;
        RECT 0.1580 58.8830 0.1760 58.9310 ;
        RECT 14.0900 58.8830 14.1080 58.9310 ;
        RECT 15.2600 58.8830 15.2870 58.9310 ;
        RECT 15.4850 58.8830 15.5210 58.9310 ;
        RECT 16.2500 58.8830 16.2680 58.9310 ;
        RECT 30.1820 58.8830 30.2000 58.9310 ;
        RECT 0.1580 59.9630 0.1760 60.0110 ;
        RECT 14.0900 59.9630 14.1080 60.0110 ;
        RECT 15.2600 59.9630 15.2870 60.0110 ;
        RECT 15.4850 59.9630 15.5210 60.0110 ;
        RECT 16.2500 59.9630 16.2680 60.0110 ;
        RECT 30.1820 59.9630 30.2000 60.0110 ;
        RECT 0.1580 61.0430 0.1760 61.0910 ;
        RECT 14.0900 61.0430 14.1080 61.0910 ;
        RECT 15.2600 61.0430 15.2870 61.0910 ;
        RECT 15.4850 61.0430 15.5210 61.0910 ;
        RECT 16.2500 61.0430 16.2680 61.0910 ;
        RECT 30.1820 61.0430 30.2000 61.0910 ;
        RECT 0.1580 62.1230 0.1760 62.1710 ;
        RECT 14.0900 62.1230 14.1080 62.1710 ;
        RECT 15.2600 62.1230 15.2870 62.1710 ;
        RECT 15.4850 62.1230 15.5210 62.1710 ;
        RECT 16.2500 62.1230 16.2680 62.1710 ;
        RECT 30.1820 62.1230 30.2000 62.1710 ;
        RECT 0.1580 63.2030 0.1760 63.2510 ;
        RECT 14.0900 63.2030 14.1080 63.2510 ;
        RECT 15.2600 63.2030 15.2870 63.2510 ;
        RECT 15.4850 63.2030 15.5210 63.2510 ;
        RECT 16.2500 63.2030 16.2680 63.2510 ;
        RECT 30.1820 63.2030 30.2000 63.2510 ;
        RECT 0.1580 64.2830 0.1760 64.3310 ;
        RECT 14.0900 64.2830 14.1080 64.3310 ;
        RECT 15.2600 64.2830 15.2870 64.3310 ;
        RECT 15.4850 64.2830 15.5210 64.3310 ;
        RECT 16.2500 64.2830 16.2680 64.3310 ;
        RECT 30.1820 64.2830 30.2000 64.3310 ;
        RECT 0.1580 65.3630 0.1760 65.4110 ;
        RECT 14.0900 65.3630 14.1080 65.4110 ;
        RECT 15.2600 65.3630 15.2870 65.4110 ;
        RECT 15.4850 65.3630 15.5210 65.4110 ;
        RECT 16.2500 65.3630 16.2680 65.4110 ;
        RECT 30.1820 65.3630 30.2000 65.4110 ;
        RECT 0.1580 66.4430 0.1760 66.4910 ;
        RECT 14.0900 66.4430 14.1080 66.4910 ;
        RECT 15.2600 66.4430 15.2870 66.4910 ;
        RECT 15.4850 66.4430 15.5210 66.4910 ;
        RECT 16.2500 66.4430 16.2680 66.4910 ;
        RECT 30.1820 66.4430 30.2000 66.4910 ;
        RECT 0.1580 67.5230 0.1760 67.5710 ;
        RECT 14.0900 67.5230 14.1080 67.5710 ;
        RECT 15.2600 67.5230 15.2870 67.5710 ;
        RECT 15.4850 67.5230 15.5210 67.5710 ;
        RECT 16.2500 67.5230 16.2680 67.5710 ;
        RECT 30.1820 67.5230 30.2000 67.5710 ;
        RECT 0.1580 68.6030 0.1760 68.6510 ;
        RECT 14.0900 68.6030 14.1080 68.6510 ;
        RECT 15.2600 68.6030 15.2870 68.6510 ;
        RECT 15.4850 68.6030 15.5210 68.6510 ;
        RECT 16.2500 68.6030 16.2680 68.6510 ;
        RECT 30.1820 68.6030 30.2000 68.6510 ;
        RECT 0.1580 69.6830 0.1760 69.7310 ;
        RECT 14.0900 69.6830 14.1080 69.7310 ;
        RECT 15.2600 69.6830 15.2870 69.7310 ;
        RECT 15.4850 69.6830 15.5210 69.7310 ;
        RECT 16.2500 69.6830 16.2680 69.7310 ;
        RECT 30.1820 69.6830 30.2000 69.7310 ;
        RECT 0.1580 70.7630 0.1760 70.8110 ;
        RECT 14.0900 70.7630 14.1080 70.8110 ;
        RECT 15.2600 70.7630 15.2870 70.8110 ;
        RECT 15.4850 70.7630 15.5210 70.8110 ;
        RECT 16.2500 70.7630 16.2680 70.8110 ;
        RECT 30.1820 70.7630 30.2000 70.8110 ;
        RECT 0.1580 71.8430 0.1760 71.8910 ;
        RECT 14.0900 71.8430 14.1080 71.8910 ;
        RECT 15.2600 71.8430 15.2870 71.8910 ;
        RECT 15.4850 71.8430 15.5210 71.8910 ;
        RECT 16.2500 71.8430 16.2680 71.8910 ;
        RECT 30.1820 71.8430 30.2000 71.8910 ;
        RECT 0.1580 72.9230 0.1760 72.9710 ;
        RECT 14.0900 72.9230 14.1080 72.9710 ;
        RECT 15.2600 72.9230 15.2870 72.9710 ;
        RECT 15.4850 72.9230 15.5210 72.9710 ;
        RECT 16.2500 72.9230 16.2680 72.9710 ;
        RECT 30.1820 72.9230 30.2000 72.9710 ;
        RECT 0.1580 74.0030 0.1760 74.0510 ;
        RECT 14.0900 74.0030 14.1080 74.0510 ;
        RECT 15.2600 74.0030 15.2870 74.0510 ;
        RECT 15.4850 74.0030 15.5210 74.0510 ;
        RECT 16.2500 74.0030 16.2680 74.0510 ;
        RECT 30.1820 74.0030 30.2000 74.0510 ;
        RECT 0.1580 75.0830 0.1760 75.1310 ;
        RECT 14.0900 75.0830 14.1080 75.1310 ;
        RECT 15.2600 75.0830 15.2870 75.1310 ;
        RECT 15.4850 75.0830 15.5210 75.1310 ;
        RECT 16.2500 75.0830 16.2680 75.1310 ;
        RECT 30.1820 75.0830 30.2000 75.1310 ;
        RECT 0.1580 76.1630 0.1760 76.2110 ;
        RECT 14.0900 76.1630 14.1080 76.2110 ;
        RECT 15.2600 76.1630 15.2870 76.2110 ;
        RECT 15.4850 76.1630 15.5210 76.2110 ;
        RECT 16.2500 76.1630 16.2680 76.2110 ;
        RECT 30.1820 76.1630 30.2000 76.2110 ;
        RECT 0.1580 77.2430 0.1760 77.2910 ;
        RECT 14.0900 77.2430 14.1080 77.2910 ;
        RECT 15.2600 77.2430 15.2870 77.2910 ;
        RECT 15.4850 77.2430 15.5210 77.2910 ;
        RECT 16.2500 77.2430 16.2680 77.2910 ;
        RECT 30.1820 77.2430 30.2000 77.2910 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.7030 36.0935 17.7210 36.1305 ;
      LAYER M4  ;
        RECT 17.6510 36.1015 17.7350 36.1255 ;
      LAYER M5  ;
        RECT 17.7000 35.1505 17.7240 38.3905 ;
      LAYER V3  ;
        RECT 17.7030 36.1015 17.7210 36.1255 ;
      LAYER V4  ;
        RECT 17.7000 36.1015 17.7240 36.1255 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.4870 36.0965 17.5050 36.1335 ;
      LAYER M4  ;
        RECT 17.4350 36.1015 17.5190 36.1255 ;
      LAYER M5  ;
        RECT 17.4840 35.1505 17.5080 38.3905 ;
      LAYER V3  ;
        RECT 17.4870 36.1015 17.5050 36.1255 ;
      LAYER V4  ;
        RECT 17.4840 36.1015 17.5080 36.1255 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.2710 35.5175 17.2890 35.5545 ;
      LAYER M4  ;
        RECT 17.2190 35.5255 17.3030 35.5495 ;
      LAYER M5  ;
        RECT 17.2680 35.1505 17.2920 38.3905 ;
      LAYER V3  ;
        RECT 17.2710 35.5255 17.2890 35.5495 ;
      LAYER V4  ;
        RECT 17.2680 35.5255 17.2920 35.5495 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.0550 35.7575 17.0730 35.9385 ;
      LAYER M4  ;
        RECT 17.0030 35.9095 17.0870 35.9335 ;
      LAYER M5  ;
        RECT 17.0520 35.1505 17.0760 38.3905 ;
      LAYER V3  ;
        RECT 17.0550 35.9095 17.0730 35.9335 ;
      LAYER V4  ;
        RECT 17.0520 35.9095 17.0760 35.9335 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.8390 35.5205 16.8570 35.5875 ;
      LAYER M4  ;
        RECT 16.7870 35.5255 16.8710 35.5495 ;
      LAYER M5  ;
        RECT 16.8360 35.1505 16.8600 38.3905 ;
      LAYER V3  ;
        RECT 16.8390 35.5255 16.8570 35.5495 ;
      LAYER V4  ;
        RECT 16.8360 35.5255 16.8600 35.5495 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.6230 35.2535 16.6410 35.5065 ;
      LAYER M4  ;
        RECT 16.5710 35.4775 16.6550 35.5015 ;
      LAYER M5  ;
        RECT 16.6200 35.1505 16.6440 38.3905 ;
      LAYER V3  ;
        RECT 16.6230 35.4775 16.6410 35.5015 ;
      LAYER V4  ;
        RECT 16.6200 35.4775 16.6440 35.5015 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.4070 36.2885 16.4250 36.3255 ;
      LAYER M4  ;
        RECT 16.3550 36.2935 16.4390 36.3175 ;
      LAYER M5  ;
        RECT 16.4040 35.1505 16.4280 38.3905 ;
      LAYER V3  ;
        RECT 16.4070 36.2935 16.4250 36.3175 ;
      LAYER V4  ;
        RECT 16.4040 36.2935 16.4280 36.3175 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.1910 36.1355 16.2090 36.2265 ;
      LAYER M4  ;
        RECT 16.1390 36.1975 16.2230 36.2215 ;
      LAYER M5  ;
        RECT 16.1880 35.1505 16.2120 38.3905 ;
      LAYER V3  ;
        RECT 16.1910 36.1975 16.2090 36.2215 ;
      LAYER V4  ;
        RECT 16.1880 36.1975 16.2120 36.2215 ;
    END
  END ADDRESS[7]
  PIN ADDRESS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.8310 35.7935 15.8490 35.9385 ;
      LAYER M4  ;
        RECT 15.8200 35.9095 16.0070 35.9335 ;
      LAYER M5  ;
        RECT 15.9720 34.8915 15.9960 38.3905 ;
      LAYER V3  ;
        RECT 15.8310 35.9095 15.8490 35.9335 ;
      LAYER V4  ;
        RECT 15.9720 35.9095 15.9960 35.9335 ;
    END
  END ADDRESS[8]
  PIN ADDRESS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.5430 35.5205 15.5610 35.5875 ;
      LAYER M4  ;
        RECT 15.2590 35.5255 15.5720 35.5495 ;
      LAYER M5  ;
        RECT 15.2700 35.1505 15.2940 38.3905 ;
      LAYER V3  ;
        RECT 15.5430 35.5255 15.5610 35.5495 ;
      LAYER V4  ;
        RECT 15.2700 35.5255 15.2940 35.5495 ;
    END
  END ADDRESS[9]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.1470 35.2535 15.1650 35.5065 ;
      LAYER M4  ;
        RECT 14.9350 35.4775 15.1760 35.5015 ;
      LAYER M5  ;
        RECT 14.9460 35.1505 14.9700 38.3905 ;
      LAYER V3  ;
        RECT 15.1470 35.4775 15.1650 35.5015 ;
      LAYER V4  ;
        RECT 14.9460 35.4775 14.9700 35.5015 ;
    END
  END banksel
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.1390 36.3845 14.1570 36.4335 ;
      LAYER M4  ;
        RECT 14.0870 36.3895 14.1710 36.4135 ;
      LAYER M5  ;
        RECT 14.1360 35.1505 14.1600 38.3905 ;
      LAYER V3  ;
        RECT 14.1390 36.3895 14.1570 36.4135 ;
      LAYER V4  ;
        RECT 14.1360 36.3895 14.1600 36.4135 ;
    END
  END clk
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.3550 35.5205 14.3730 35.5875 ;
      LAYER M4  ;
        RECT 14.3030 35.5255 14.3870 35.5495 ;
      LAYER M5  ;
        RECT 14.3520 35.1505 14.3760 38.3905 ;
      LAYER V3  ;
        RECT 14.3550 35.5255 14.3730 35.5495 ;
      LAYER V4  ;
        RECT 14.3520 35.5255 14.3760 35.5495 ;
    END
  END write
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.1750 35.2535 14.1930 35.5065 ;
      LAYER M4  ;
        RECT 13.9090 35.4775 14.2040 35.5015 ;
      LAYER M5  ;
        RECT 13.9200 35.1505 13.9440 38.3905 ;
      LAYER V3  ;
        RECT 14.1750 35.4775 14.1930 35.5015 ;
      LAYER V4  ;
        RECT 13.9200 35.4775 13.9440 35.5015 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.7070 36.0935 13.7250 36.1305 ;
      LAYER M4  ;
        RECT 13.6550 36.1015 13.7390 36.1255 ;
      LAYER M5  ;
        RECT 13.7040 35.1505 13.7280 38.3905 ;
      LAYER V3  ;
        RECT 13.7070 36.1015 13.7250 36.1255 ;
      LAYER V4  ;
        RECT 13.7040 36.1015 13.7280 36.1255 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.4910 35.5205 13.5090 35.7495 ;
      LAYER M4  ;
        RECT 13.4390 35.5255 13.5230 35.5495 ;
      LAYER M5  ;
        RECT 13.4880 35.1505 13.5120 38.3905 ;
      LAYER V3  ;
        RECT 13.4910 35.5255 13.5090 35.5495 ;
      LAYER V4  ;
        RECT 13.4880 35.5255 13.5120 35.5495 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.2750 35.2535 13.2930 35.5065 ;
      LAYER M4  ;
        RECT 13.2230 35.4775 13.3070 35.5015 ;
      LAYER M5  ;
        RECT 13.2720 35.1505 13.2960 38.3905 ;
      LAYER V3  ;
        RECT 13.2750 35.4775 13.2930 35.5015 ;
      LAYER V4  ;
        RECT 13.2720 35.4775 13.2960 35.5015 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.0590 35.5175 13.0770 35.5545 ;
      LAYER M4  ;
        RECT 13.0070 35.5255 13.0910 35.5495 ;
      LAYER M5  ;
        RECT 13.0560 35.1505 13.0800 38.3905 ;
      LAYER V3  ;
        RECT 13.0590 35.5255 13.0770 35.5495 ;
      LAYER V4  ;
        RECT 13.0560 35.5255 13.0800 35.5495 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 12.8430 36.0935 12.8610 36.1305 ;
      LAYER M4  ;
        RECT 12.7910 36.1015 12.8750 36.1255 ;
      LAYER M5  ;
        RECT 12.8400 35.1505 12.8640 38.3905 ;
      LAYER V3  ;
        RECT 12.8430 36.1015 12.8610 36.1255 ;
      LAYER V4  ;
        RECT 12.8400 36.1015 12.8640 36.1255 ;
    END
  END sdel[4]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 15.4975 15.4670 15.7370 ;
      LAYER M4  ;
        RECT 14.8610 15.5480 15.5090 15.5720 ;
      LAYER V3  ;
        RECT 15.4490 15.5480 15.4670 15.5720 ;
    END
  END dataout[14]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 14.4175 15.4670 14.6570 ;
      LAYER M4  ;
        RECT 14.8610 14.4680 15.5090 14.4920 ;
      LAYER V3  ;
        RECT 15.4490 14.4680 15.4670 14.4920 ;
    END
  END dataout[13]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 13.3375 15.4670 13.5770 ;
      LAYER M4  ;
        RECT 14.8610 13.3880 15.5090 13.4120 ;
      LAYER V3  ;
        RECT 15.4490 13.3880 15.4670 13.4120 ;
    END
  END dataout[12]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 12.2575 15.4670 12.4970 ;
      LAYER M4  ;
        RECT 14.8610 12.3080 15.5090 12.3320 ;
      LAYER V3  ;
        RECT 15.4490 12.3080 15.4670 12.3320 ;
    END
  END dataout[11]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 11.1775 15.4670 11.4170 ;
      LAYER M4  ;
        RECT 14.8610 11.2280 15.5090 11.2520 ;
      LAYER V3  ;
        RECT 15.4490 11.2280 15.4670 11.2520 ;
    END
  END dataout[10]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 0.3775 15.4670 0.6170 ;
      LAYER M4  ;
        RECT 14.8610 0.4280 15.5090 0.4520 ;
      LAYER V3  ;
        RECT 15.4490 0.4280 15.4670 0.4520 ;
    END
  END dataout[0]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 16.5775 15.4670 16.8170 ;
      LAYER M4  ;
        RECT 14.8610 16.6280 15.5090 16.6520 ;
      LAYER V3  ;
        RECT 15.4490 16.6280 15.4670 16.6520 ;
    END
  END dataout[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 17.6575 15.4670 17.8970 ;
      LAYER M4  ;
        RECT 14.8610 17.7080 15.5090 17.7320 ;
      LAYER V3  ;
        RECT 15.4490 17.7080 15.4670 17.7320 ;
    END
  END dataout[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 18.7375 15.4670 18.9770 ;
      LAYER M4  ;
        RECT 14.8610 18.7880 15.5090 18.8120 ;
      LAYER V3  ;
        RECT 15.4490 18.7880 15.4670 18.8120 ;
    END
  END dataout[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 19.8175 15.4670 20.0570 ;
      LAYER M4  ;
        RECT 14.8610 19.8680 15.5090 19.8920 ;
      LAYER V3  ;
        RECT 15.4490 19.8680 15.4670 19.8920 ;
    END
  END dataout[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 20.8975 15.4670 21.1370 ;
      LAYER M4  ;
        RECT 14.8610 20.9480 15.5090 20.9720 ;
      LAYER V3  ;
        RECT 15.4490 20.9480 15.4670 20.9720 ;
    END
  END dataout[19]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 1.4575 15.4670 1.6970 ;
      LAYER M4  ;
        RECT 14.8610 1.5080 15.5090 1.5320 ;
      LAYER V3  ;
        RECT 15.4490 1.5080 15.4670 1.5320 ;
    END
  END dataout[1]
  PIN dataout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 21.9775 15.4670 22.2170 ;
      LAYER M4  ;
        RECT 14.8610 22.0280 15.5090 22.0520 ;
      LAYER V3  ;
        RECT 15.4490 22.0280 15.4670 22.0520 ;
    END
  END dataout[20]
  PIN dataout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 23.0575 15.4670 23.2970 ;
      LAYER M4  ;
        RECT 14.8610 23.1080 15.5090 23.1320 ;
      LAYER V3  ;
        RECT 15.4490 23.1080 15.4670 23.1320 ;
    END
  END dataout[21]
  PIN dataout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 24.1375 15.4670 24.3770 ;
      LAYER M4  ;
        RECT 14.8610 24.1880 15.5090 24.2120 ;
      LAYER V3  ;
        RECT 15.4490 24.1880 15.4670 24.2120 ;
    END
  END dataout[22]
  PIN dataout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 25.2175 15.4670 25.4570 ;
      LAYER M4  ;
        RECT 14.8610 25.2680 15.5090 25.2920 ;
      LAYER V3  ;
        RECT 15.4490 25.2680 15.4670 25.2920 ;
    END
  END dataout[23]
  PIN dataout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 26.2975 15.4670 26.5370 ;
      LAYER M4  ;
        RECT 14.8610 26.3480 15.5090 26.3720 ;
      LAYER V3  ;
        RECT 15.4490 26.3480 15.4670 26.3720 ;
    END
  END dataout[24]
  PIN dataout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 27.3775 15.4670 27.6170 ;
      LAYER M4  ;
        RECT 14.8610 27.4280 15.5090 27.4520 ;
      LAYER V3  ;
        RECT 15.4490 27.4280 15.4670 27.4520 ;
    END
  END dataout[25]
  PIN dataout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 28.4575 15.4670 28.6970 ;
      LAYER M4  ;
        RECT 14.8610 28.5080 15.5090 28.5320 ;
      LAYER V3  ;
        RECT 15.4490 28.5080 15.4670 28.5320 ;
    END
  END dataout[26]
  PIN dataout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 29.5375 15.4670 29.7770 ;
      LAYER M4  ;
        RECT 14.8610 29.5880 15.5090 29.6120 ;
      LAYER V3  ;
        RECT 15.4490 29.5880 15.4670 29.6120 ;
    END
  END dataout[27]
  PIN dataout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 30.6175 15.4670 30.8570 ;
      LAYER M4  ;
        RECT 14.8610 30.6680 15.5090 30.6920 ;
      LAYER V3  ;
        RECT 15.4490 30.6680 15.4670 30.6920 ;
    END
  END dataout[28]
  PIN dataout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 31.6975 15.4670 31.9370 ;
      LAYER M4  ;
        RECT 14.8610 31.7480 15.5090 31.7720 ;
      LAYER V3  ;
        RECT 15.4490 31.7480 15.4670 31.7720 ;
    END
  END dataout[29]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 2.5375 15.4670 2.7770 ;
      LAYER M4  ;
        RECT 14.8610 2.5880 15.5090 2.6120 ;
      LAYER V3  ;
        RECT 15.4490 2.5880 15.4670 2.6120 ;
    END
  END dataout[2]
  PIN dataout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 32.7775 15.4670 33.0170 ;
      LAYER M4  ;
        RECT 14.8610 32.8280 15.5090 32.8520 ;
      LAYER V3  ;
        RECT 15.4490 32.8280 15.4670 32.8520 ;
    END
  END dataout[30]
  PIN dataout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 33.8575 15.4670 34.0970 ;
      LAYER M4  ;
        RECT 14.8610 33.9080 15.5090 33.9320 ;
      LAYER V3  ;
        RECT 15.4490 33.9080 15.4670 33.9320 ;
    END
  END dataout[31]
  PIN dataout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 43.0645 15.4670 43.3040 ;
      LAYER M4  ;
        RECT 14.8610 43.1150 15.5090 43.1390 ;
      LAYER V3  ;
        RECT 15.4490 43.1150 15.4670 43.1390 ;
    END
  END dataout[32]
  PIN dataout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 44.1445 15.4670 44.3840 ;
      LAYER M4  ;
        RECT 14.8610 44.1950 15.5090 44.2190 ;
      LAYER V3  ;
        RECT 15.4490 44.1950 15.4670 44.2190 ;
    END
  END dataout[33]
  PIN dataout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 45.2245 15.4670 45.4640 ;
      LAYER M4  ;
        RECT 14.8610 45.2750 15.5090 45.2990 ;
      LAYER V3  ;
        RECT 15.4490 45.2750 15.4670 45.2990 ;
    END
  END dataout[34]
  PIN dataout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 46.3045 15.4670 46.5440 ;
      LAYER M4  ;
        RECT 14.8610 46.3550 15.5090 46.3790 ;
      LAYER V3  ;
        RECT 15.4490 46.3550 15.4670 46.3790 ;
    END
  END dataout[35]
  PIN dataout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 47.3845 15.4670 47.6240 ;
      LAYER M4  ;
        RECT 14.8610 47.4350 15.5090 47.4590 ;
      LAYER V3  ;
        RECT 15.4490 47.4350 15.4670 47.4590 ;
    END
  END dataout[36]
  PIN dataout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 48.4645 15.4670 48.7040 ;
      LAYER M4  ;
        RECT 14.8610 48.5150 15.5090 48.5390 ;
      LAYER V3  ;
        RECT 15.4490 48.5150 15.4670 48.5390 ;
    END
  END dataout[37]
  PIN dataout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 49.5445 15.4670 49.7840 ;
      LAYER M4  ;
        RECT 14.8610 49.5950 15.5090 49.6190 ;
      LAYER V3  ;
        RECT 15.4490 49.5950 15.4670 49.6190 ;
    END
  END dataout[38]
  PIN dataout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 50.6245 15.4670 50.8640 ;
      LAYER M4  ;
        RECT 14.8610 50.6750 15.5090 50.6990 ;
      LAYER V3  ;
        RECT 15.4490 50.6750 15.4670 50.6990 ;
    END
  END dataout[39]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 3.6175 15.4670 3.8570 ;
      LAYER M4  ;
        RECT 14.8610 3.6680 15.5090 3.6920 ;
      LAYER V3  ;
        RECT 15.4490 3.6680 15.4670 3.6920 ;
    END
  END dataout[3]
  PIN dataout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 51.7045 15.4670 51.9440 ;
      LAYER M4  ;
        RECT 14.8610 51.7550 15.5090 51.7790 ;
      LAYER V3  ;
        RECT 15.4490 51.7550 15.4670 51.7790 ;
    END
  END dataout[40]
  PIN dataout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 52.7845 15.4670 53.0240 ;
      LAYER M4  ;
        RECT 14.8610 52.8350 15.5090 52.8590 ;
      LAYER V3  ;
        RECT 15.4490 52.8350 15.4670 52.8590 ;
    END
  END dataout[41]
  PIN dataout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 53.8645 15.4670 54.1040 ;
      LAYER M4  ;
        RECT 14.8610 53.9150 15.5090 53.9390 ;
      LAYER V3  ;
        RECT 15.4490 53.9150 15.4670 53.9390 ;
    END
  END dataout[42]
  PIN dataout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 54.9445 15.4670 55.1840 ;
      LAYER M4  ;
        RECT 14.8610 54.9950 15.5090 55.0190 ;
      LAYER V3  ;
        RECT 15.4490 54.9950 15.4670 55.0190 ;
    END
  END dataout[43]
  PIN dataout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 56.0245 15.4670 56.2640 ;
      LAYER M4  ;
        RECT 14.8610 56.0750 15.5090 56.0990 ;
      LAYER V3  ;
        RECT 15.4490 56.0750 15.4670 56.0990 ;
    END
  END dataout[44]
  PIN dataout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 57.1045 15.4670 57.3440 ;
      LAYER M4  ;
        RECT 14.8610 57.1550 15.5090 57.1790 ;
      LAYER V3  ;
        RECT 15.4490 57.1550 15.4670 57.1790 ;
    END
  END dataout[45]
  PIN dataout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 58.1845 15.4670 58.4240 ;
      LAYER M4  ;
        RECT 14.8610 58.2350 15.5090 58.2590 ;
      LAYER V3  ;
        RECT 15.4490 58.2350 15.4670 58.2590 ;
    END
  END dataout[46]
  PIN dataout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 59.2645 15.4670 59.5040 ;
      LAYER M4  ;
        RECT 14.8610 59.3150 15.5090 59.3390 ;
      LAYER V3  ;
        RECT 15.4490 59.3150 15.4670 59.3390 ;
    END
  END dataout[47]
  PIN dataout[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 60.3445 15.4670 60.5840 ;
      LAYER M4  ;
        RECT 14.8610 60.3950 15.5090 60.4190 ;
      LAYER V3  ;
        RECT 15.4490 60.3950 15.4670 60.4190 ;
    END
  END dataout[48]
  PIN dataout[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 61.4245 15.4670 61.6640 ;
      LAYER M4  ;
        RECT 14.8610 61.4750 15.5090 61.4990 ;
      LAYER V3  ;
        RECT 15.4490 61.4750 15.4670 61.4990 ;
    END
  END dataout[49]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 4.6975 15.4670 4.9370 ;
      LAYER M4  ;
        RECT 14.8610 4.7480 15.5090 4.7720 ;
      LAYER V3  ;
        RECT 15.4490 4.7480 15.4670 4.7720 ;
    END
  END dataout[4]
  PIN dataout[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 62.5045 15.4670 62.7440 ;
      LAYER M4  ;
        RECT 14.8610 62.5550 15.5090 62.5790 ;
      LAYER V3  ;
        RECT 15.4490 62.5550 15.4670 62.5790 ;
    END
  END dataout[50]
  PIN dataout[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 63.5845 15.4670 63.8240 ;
      LAYER M4  ;
        RECT 14.8610 63.6350 15.5090 63.6590 ;
      LAYER V3  ;
        RECT 15.4490 63.6350 15.4670 63.6590 ;
    END
  END dataout[51]
  PIN dataout[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 64.6645 15.4670 64.9040 ;
      LAYER M4  ;
        RECT 14.8610 64.7150 15.5090 64.7390 ;
      LAYER V3  ;
        RECT 15.4490 64.7150 15.4670 64.7390 ;
    END
  END dataout[52]
  PIN dataout[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 65.7445 15.4670 65.9840 ;
      LAYER M4  ;
        RECT 14.8610 65.7950 15.5090 65.8190 ;
      LAYER V3  ;
        RECT 15.4490 65.7950 15.4670 65.8190 ;
    END
  END dataout[53]
  PIN dataout[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 66.8245 15.4670 67.0640 ;
      LAYER M4  ;
        RECT 14.8610 66.8750 15.5090 66.8990 ;
      LAYER V3  ;
        RECT 15.4490 66.8750 15.4670 66.8990 ;
    END
  END dataout[54]
  PIN dataout[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 67.9045 15.4670 68.1440 ;
      LAYER M4  ;
        RECT 14.8610 67.9550 15.5090 67.9790 ;
      LAYER V3  ;
        RECT 15.4490 67.9550 15.4670 67.9790 ;
    END
  END dataout[55]
  PIN dataout[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 68.9845 15.4670 69.2240 ;
      LAYER M4  ;
        RECT 14.8610 69.0350 15.5090 69.0590 ;
      LAYER V3  ;
        RECT 15.4490 69.0350 15.4670 69.0590 ;
    END
  END dataout[56]
  PIN dataout[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 70.0645 15.4670 70.3040 ;
      LAYER M4  ;
        RECT 14.8610 70.1150 15.5090 70.1390 ;
      LAYER V3  ;
        RECT 15.4490 70.1150 15.4670 70.1390 ;
    END
  END dataout[57]
  PIN dataout[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 71.1445 15.4670 71.3840 ;
      LAYER M4  ;
        RECT 14.8610 71.1950 15.5090 71.2190 ;
      LAYER V3  ;
        RECT 15.4490 71.1950 15.4670 71.2190 ;
    END
  END dataout[58]
  PIN dataout[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 72.2245 15.4670 72.4640 ;
      LAYER M4  ;
        RECT 14.8610 72.2750 15.5090 72.2990 ;
      LAYER V3  ;
        RECT 15.4490 72.2750 15.4670 72.2990 ;
    END
  END dataout[59]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 5.7775 15.4670 6.0170 ;
      LAYER M4  ;
        RECT 14.8610 5.8280 15.5090 5.8520 ;
      LAYER V3  ;
        RECT 15.4490 5.8280 15.4670 5.8520 ;
    END
  END dataout[5]
  PIN dataout[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 73.3045 15.4670 73.5440 ;
      LAYER M4  ;
        RECT 14.8610 73.3550 15.5090 73.3790 ;
      LAYER V3  ;
        RECT 15.4490 73.3550 15.4670 73.3790 ;
    END
  END dataout[60]
  PIN dataout[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 74.3845 15.4670 74.6240 ;
      LAYER M4  ;
        RECT 14.8610 74.4350 15.5090 74.4590 ;
      LAYER V3  ;
        RECT 15.4490 74.4350 15.4670 74.4590 ;
    END
  END dataout[61]
  PIN dataout[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 75.4645 15.4670 75.7040 ;
      LAYER M4  ;
        RECT 14.8610 75.5150 15.5090 75.5390 ;
      LAYER V3  ;
        RECT 15.4490 75.5150 15.4670 75.5390 ;
    END
  END dataout[62]
  PIN dataout[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 76.5445 15.4670 76.7840 ;
      LAYER M4  ;
        RECT 14.8610 76.5950 15.5090 76.6190 ;
      LAYER V3  ;
        RECT 15.4490 76.5950 15.4670 76.6190 ;
    END
  END dataout[63]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 6.8575 15.4670 7.0970 ;
      LAYER M4  ;
        RECT 14.8610 6.9080 15.5090 6.9320 ;
      LAYER V3  ;
        RECT 15.4490 6.9080 15.4670 6.9320 ;
    END
  END dataout[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 7.9375 15.4670 8.1770 ;
      LAYER M4  ;
        RECT 14.8610 7.9880 15.5090 8.0120 ;
      LAYER V3  ;
        RECT 15.4490 7.9880 15.4670 8.0120 ;
    END
  END dataout[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 9.0175 15.4670 9.2570 ;
      LAYER M4  ;
        RECT 14.8610 9.0680 15.5090 9.0920 ;
      LAYER V3  ;
        RECT 15.4490 9.0680 15.4670 9.0920 ;
    END
  END dataout[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 10.0975 15.4670 10.3370 ;
      LAYER M4  ;
        RECT 14.8610 10.1480 15.5090 10.1720 ;
      LAYER V3  ;
        RECT 15.4490 10.1480 15.4670 10.1720 ;
    END
  END dataout[9]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 0.2700 15.2420 0.6750 ;
      LAYER M4  ;
        RECT 14.8610 0.3320 15.4970 0.3560 ;
      LAYER V3  ;
        RECT 15.2240 0.3320 15.2420 0.3560 ;
    END
  END wd[0]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 11.0700 15.2420 11.4750 ;
      LAYER M4  ;
        RECT 14.8610 11.1320 15.4970 11.1560 ;
      LAYER V3  ;
        RECT 15.2240 11.1320 15.2420 11.1560 ;
    END
  END wd[10]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 12.1500 15.2420 12.5550 ;
      LAYER M4  ;
        RECT 14.8610 12.2120 15.4970 12.2360 ;
      LAYER V3  ;
        RECT 15.2240 12.2120 15.2420 12.2360 ;
    END
  END wd[11]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 13.2300 15.2420 13.6350 ;
      LAYER M4  ;
        RECT 14.8610 13.2920 15.4970 13.3160 ;
      LAYER V3  ;
        RECT 15.2240 13.2920 15.2420 13.3160 ;
    END
  END wd[12]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 14.3100 15.2420 14.7150 ;
      LAYER M4  ;
        RECT 14.8610 14.3720 15.4970 14.3960 ;
      LAYER V3  ;
        RECT 15.2240 14.3720 15.2420 14.3960 ;
    END
  END wd[13]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 15.3900 15.2420 15.7950 ;
      LAYER M4  ;
        RECT 14.8610 15.4520 15.4970 15.4760 ;
      LAYER V3  ;
        RECT 15.2240 15.4520 15.2420 15.4760 ;
    END
  END wd[14]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 16.4700 15.2420 16.8750 ;
      LAYER M4  ;
        RECT 14.8610 16.5320 15.4970 16.5560 ;
      LAYER V3  ;
        RECT 15.2240 16.5320 15.2420 16.5560 ;
    END
  END wd[15]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 17.5500 15.2420 17.9550 ;
      LAYER M4  ;
        RECT 14.8610 17.6120 15.4970 17.6360 ;
      LAYER V3  ;
        RECT 15.2240 17.6120 15.2420 17.6360 ;
    END
  END wd[16]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 18.6300 15.2420 19.0350 ;
      LAYER M4  ;
        RECT 14.8610 18.6920 15.4970 18.7160 ;
      LAYER V3  ;
        RECT 15.2240 18.6920 15.2420 18.7160 ;
    END
  END wd[17]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 19.7100 15.2420 20.1150 ;
      LAYER M4  ;
        RECT 14.8610 19.7720 15.4970 19.7960 ;
      LAYER V3  ;
        RECT 15.2240 19.7720 15.2420 19.7960 ;
    END
  END wd[18]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 20.7900 15.2420 21.1950 ;
      LAYER M4  ;
        RECT 14.8610 20.8520 15.4970 20.8760 ;
      LAYER V3  ;
        RECT 15.2240 20.8520 15.2420 20.8760 ;
    END
  END wd[19]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 1.3500 15.2420 1.7550 ;
      LAYER M4  ;
        RECT 14.8610 1.4120 15.4970 1.4360 ;
      LAYER V3  ;
        RECT 15.2240 1.4120 15.2420 1.4360 ;
    END
  END wd[1]
  PIN wd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 21.8700 15.2420 22.2750 ;
      LAYER M4  ;
        RECT 14.8610 21.9320 15.4970 21.9560 ;
      LAYER V3  ;
        RECT 15.2240 21.9320 15.2420 21.9560 ;
    END
  END wd[20]
  PIN wd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 22.9500 15.2420 23.3550 ;
      LAYER M4  ;
        RECT 14.8610 23.0120 15.4970 23.0360 ;
      LAYER V3  ;
        RECT 15.2240 23.0120 15.2420 23.0360 ;
    END
  END wd[21]
  PIN wd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 24.0300 15.2420 24.4350 ;
      LAYER M4  ;
        RECT 14.8610 24.0920 15.4970 24.1160 ;
      LAYER V3  ;
        RECT 15.2240 24.0920 15.2420 24.1160 ;
    END
  END wd[22]
  PIN wd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 25.1100 15.2420 25.5150 ;
      LAYER M4  ;
        RECT 14.8610 25.1720 15.4970 25.1960 ;
      LAYER V3  ;
        RECT 15.2240 25.1720 15.2420 25.1960 ;
    END
  END wd[23]
  PIN wd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 26.1900 15.2420 26.5950 ;
      LAYER M4  ;
        RECT 14.8610 26.2520 15.4970 26.2760 ;
      LAYER V3  ;
        RECT 15.2240 26.2520 15.2420 26.2760 ;
    END
  END wd[24]
  PIN wd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 27.2700 15.2420 27.6750 ;
      LAYER M4  ;
        RECT 14.8610 27.3320 15.4970 27.3560 ;
      LAYER V3  ;
        RECT 15.2240 27.3320 15.2420 27.3560 ;
    END
  END wd[25]
  PIN wd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 28.3500 15.2420 28.7550 ;
      LAYER M4  ;
        RECT 14.8610 28.4120 15.4970 28.4360 ;
      LAYER V3  ;
        RECT 15.2240 28.4120 15.2420 28.4360 ;
    END
  END wd[26]
  PIN wd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 29.4300 15.2420 29.8350 ;
      LAYER M4  ;
        RECT 14.8610 29.4920 15.4970 29.5160 ;
      LAYER V3  ;
        RECT 15.2240 29.4920 15.2420 29.5160 ;
    END
  END wd[27]
  PIN wd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 30.5100 15.2420 30.9150 ;
      LAYER M4  ;
        RECT 14.8610 30.5720 15.4970 30.5960 ;
      LAYER V3  ;
        RECT 15.2240 30.5720 15.2420 30.5960 ;
    END
  END wd[28]
  PIN wd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 31.5900 15.2420 31.9950 ;
      LAYER M4  ;
        RECT 14.8610 31.6520 15.4970 31.6760 ;
      LAYER V3  ;
        RECT 15.2240 31.6520 15.2420 31.6760 ;
    END
  END wd[29]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 2.4300 15.2420 2.8350 ;
      LAYER M4  ;
        RECT 14.8610 2.4920 15.4970 2.5160 ;
      LAYER V3  ;
        RECT 15.2240 2.4920 15.2420 2.5160 ;
    END
  END wd[2]
  PIN wd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 32.6700 15.2420 33.0750 ;
      LAYER M4  ;
        RECT 14.8610 32.7320 15.4970 32.7560 ;
      LAYER V3  ;
        RECT 15.2240 32.7320 15.2420 32.7560 ;
    END
  END wd[30]
  PIN wd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 33.7500 15.2420 34.1550 ;
      LAYER M4  ;
        RECT 14.8610 33.8120 15.4970 33.8360 ;
      LAYER V3  ;
        RECT 15.2240 33.8120 15.2420 33.8360 ;
    END
  END wd[31]
  PIN wd[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 42.9570 15.2420 43.3620 ;
      LAYER M4  ;
        RECT 14.8610 43.0190 15.4970 43.0430 ;
      LAYER V3  ;
        RECT 15.2240 43.0190 15.2420 43.0430 ;
    END
  END wd[32]
  PIN wd[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 44.0370 15.2420 44.4420 ;
      LAYER M4  ;
        RECT 14.8610 44.0990 15.4970 44.1230 ;
      LAYER V3  ;
        RECT 15.2240 44.0990 15.2420 44.1230 ;
    END
  END wd[33]
  PIN wd[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 45.1170 15.2420 45.5220 ;
      LAYER M4  ;
        RECT 14.8610 45.1790 15.4970 45.2030 ;
      LAYER V3  ;
        RECT 15.2240 45.1790 15.2420 45.2030 ;
    END
  END wd[34]
  PIN wd[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 46.1970 15.2420 46.6020 ;
      LAYER M4  ;
        RECT 14.8610 46.2590 15.4970 46.2830 ;
      LAYER V3  ;
        RECT 15.2240 46.2590 15.2420 46.2830 ;
    END
  END wd[35]
  PIN wd[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 47.2770 15.2420 47.6820 ;
      LAYER M4  ;
        RECT 14.8610 47.3390 15.4970 47.3630 ;
      LAYER V3  ;
        RECT 15.2240 47.3390 15.2420 47.3630 ;
    END
  END wd[36]
  PIN wd[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 48.3570 15.2420 48.7620 ;
      LAYER M4  ;
        RECT 14.8610 48.4190 15.4970 48.4430 ;
      LAYER V3  ;
        RECT 15.2240 48.4190 15.2420 48.4430 ;
    END
  END wd[37]
  PIN wd[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 49.4370 15.2420 49.8420 ;
      LAYER M4  ;
        RECT 14.8610 49.4990 15.4970 49.5230 ;
      LAYER V3  ;
        RECT 15.2240 49.4990 15.2420 49.5230 ;
    END
  END wd[38]
  PIN wd[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 50.5170 15.2420 50.9220 ;
      LAYER M4  ;
        RECT 14.8610 50.5790 15.4970 50.6030 ;
      LAYER V3  ;
        RECT 15.2240 50.5790 15.2420 50.6030 ;
    END
  END wd[39]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 3.5100 15.2420 3.9150 ;
      LAYER M4  ;
        RECT 14.8610 3.5720 15.4970 3.5960 ;
      LAYER V3  ;
        RECT 15.2240 3.5720 15.2420 3.5960 ;
    END
  END wd[3]
  PIN wd[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 51.5970 15.2420 52.0020 ;
      LAYER M4  ;
        RECT 14.8610 51.6590 15.4970 51.6830 ;
      LAYER V3  ;
        RECT 15.2240 51.6590 15.2420 51.6830 ;
    END
  END wd[40]
  PIN wd[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 52.6770 15.2420 53.0820 ;
      LAYER M4  ;
        RECT 14.8610 52.7390 15.4970 52.7630 ;
      LAYER V3  ;
        RECT 15.2240 52.7390 15.2420 52.7630 ;
    END
  END wd[41]
  PIN wd[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 53.7570 15.2420 54.1620 ;
      LAYER M4  ;
        RECT 14.8610 53.8190 15.4970 53.8430 ;
      LAYER V3  ;
        RECT 15.2240 53.8190 15.2420 53.8430 ;
    END
  END wd[42]
  PIN wd[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 54.8370 15.2420 55.2420 ;
      LAYER M4  ;
        RECT 14.8610 54.8990 15.4970 54.9230 ;
      LAYER V3  ;
        RECT 15.2240 54.8990 15.2420 54.9230 ;
    END
  END wd[43]
  PIN wd[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 55.9170 15.2420 56.3220 ;
      LAYER M4  ;
        RECT 14.8610 55.9790 15.4970 56.0030 ;
      LAYER V3  ;
        RECT 15.2240 55.9790 15.2420 56.0030 ;
    END
  END wd[44]
  PIN wd[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 56.9970 15.2420 57.4020 ;
      LAYER M4  ;
        RECT 14.8610 57.0590 15.4970 57.0830 ;
      LAYER V3  ;
        RECT 15.2240 57.0590 15.2420 57.0830 ;
    END
  END wd[45]
  PIN wd[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 58.0770 15.2420 58.4820 ;
      LAYER M4  ;
        RECT 14.8610 58.1390 15.4970 58.1630 ;
      LAYER V3  ;
        RECT 15.2240 58.1390 15.2420 58.1630 ;
    END
  END wd[46]
  PIN wd[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 59.1570 15.2420 59.5620 ;
      LAYER M4  ;
        RECT 14.8610 59.2190 15.4970 59.2430 ;
      LAYER V3  ;
        RECT 15.2240 59.2190 15.2420 59.2430 ;
    END
  END wd[47]
  PIN wd[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 60.2370 15.2420 60.6420 ;
      LAYER M4  ;
        RECT 14.8610 60.2990 15.4970 60.3230 ;
      LAYER V3  ;
        RECT 15.2240 60.2990 15.2420 60.3230 ;
    END
  END wd[48]
  PIN wd[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 61.3170 15.2420 61.7220 ;
      LAYER M4  ;
        RECT 14.8610 61.3790 15.4970 61.4030 ;
      LAYER V3  ;
        RECT 15.2240 61.3790 15.2420 61.4030 ;
    END
  END wd[49]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 4.5900 15.2420 4.9950 ;
      LAYER M4  ;
        RECT 14.8610 4.6520 15.4970 4.6760 ;
      LAYER V3  ;
        RECT 15.2240 4.6520 15.2420 4.6760 ;
    END
  END wd[4]
  PIN wd[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 62.3970 15.2420 62.8020 ;
      LAYER M4  ;
        RECT 14.8610 62.4590 15.4970 62.4830 ;
      LAYER V3  ;
        RECT 15.2240 62.4590 15.2420 62.4830 ;
    END
  END wd[50]
  PIN wd[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 63.4770 15.2420 63.8820 ;
      LAYER M4  ;
        RECT 14.8610 63.5390 15.4970 63.5630 ;
      LAYER V3  ;
        RECT 15.2240 63.5390 15.2420 63.5630 ;
    END
  END wd[51]
  PIN wd[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 64.5570 15.2420 64.9620 ;
      LAYER M4  ;
        RECT 14.8610 64.6190 15.4970 64.6430 ;
      LAYER V3  ;
        RECT 15.2240 64.6190 15.2420 64.6430 ;
    END
  END wd[52]
  PIN wd[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 65.6370 15.2420 66.0420 ;
      LAYER M4  ;
        RECT 14.8610 65.6990 15.4970 65.7230 ;
      LAYER V3  ;
        RECT 15.2240 65.6990 15.2420 65.7230 ;
    END
  END wd[53]
  PIN wd[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 66.7170 15.2420 67.1220 ;
      LAYER M4  ;
        RECT 14.8610 66.7790 15.4970 66.8030 ;
      LAYER V3  ;
        RECT 15.2240 66.7790 15.2420 66.8030 ;
    END
  END wd[54]
  PIN wd[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 67.7970 15.2420 68.2020 ;
      LAYER M4  ;
        RECT 14.8610 67.8590 15.4970 67.8830 ;
      LAYER V3  ;
        RECT 15.2240 67.8590 15.2420 67.8830 ;
    END
  END wd[55]
  PIN wd[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 68.8770 15.2420 69.2820 ;
      LAYER M4  ;
        RECT 14.8610 68.9390 15.4970 68.9630 ;
      LAYER V3  ;
        RECT 15.2240 68.9390 15.2420 68.9630 ;
    END
  END wd[56]
  PIN wd[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 69.9570 15.2420 70.3620 ;
      LAYER M4  ;
        RECT 14.8610 70.0190 15.4970 70.0430 ;
      LAYER V3  ;
        RECT 15.2240 70.0190 15.2420 70.0430 ;
    END
  END wd[57]
  PIN wd[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 71.0370 15.2420 71.4420 ;
      LAYER M4  ;
        RECT 14.8610 71.0990 15.4970 71.1230 ;
      LAYER V3  ;
        RECT 15.2240 71.0990 15.2420 71.1230 ;
    END
  END wd[58]
  PIN wd[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 72.1170 15.2420 72.5220 ;
      LAYER M4  ;
        RECT 14.8610 72.1790 15.4970 72.2030 ;
      LAYER V3  ;
        RECT 15.2240 72.1790 15.2420 72.2030 ;
    END
  END wd[59]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 5.6700 15.2420 6.0750 ;
      LAYER M4  ;
        RECT 14.8610 5.7320 15.4970 5.7560 ;
      LAYER V3  ;
        RECT 15.2240 5.7320 15.2420 5.7560 ;
    END
  END wd[5]
  PIN wd[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 73.1970 15.2420 73.6020 ;
      LAYER M4  ;
        RECT 14.8610 73.2590 15.4970 73.2830 ;
      LAYER V3  ;
        RECT 15.2240 73.2590 15.2420 73.2830 ;
    END
  END wd[60]
  PIN wd[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 74.2770 15.2420 74.6820 ;
      LAYER M4  ;
        RECT 14.8610 74.3390 15.4970 74.3630 ;
      LAYER V3  ;
        RECT 15.2240 74.3390 15.2420 74.3630 ;
    END
  END wd[61]
  PIN wd[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 75.3570 15.2420 75.7620 ;
      LAYER M4  ;
        RECT 14.8610 75.4190 15.4970 75.4430 ;
      LAYER V3  ;
        RECT 15.2240 75.4190 15.2420 75.4430 ;
    END
  END wd[62]
  PIN wd[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 76.4370 15.2420 76.8420 ;
      LAYER M4  ;
        RECT 14.8610 76.4990 15.4970 76.5230 ;
      LAYER V3  ;
        RECT 15.2240 76.4990 15.2420 76.5230 ;
    END
  END wd[63]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 6.7500 15.2420 7.1550 ;
      LAYER M4  ;
        RECT 14.8610 6.8120 15.4970 6.8360 ;
      LAYER V3  ;
        RECT 15.2240 6.8120 15.2420 6.8360 ;
    END
  END wd[6]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 7.8300 15.2420 8.2350 ;
      LAYER M4  ;
        RECT 14.8610 7.8920 15.4970 7.9160 ;
      LAYER V3  ;
        RECT 15.2240 7.8920 15.2420 7.9160 ;
    END
  END wd[7]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 8.9100 15.2420 9.3150 ;
      LAYER M4  ;
        RECT 14.8610 8.9720 15.4970 8.9960 ;
      LAYER V3  ;
        RECT 15.2240 8.9720 15.2420 8.9960 ;
    END
  END wd[8]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 9.9900 15.2420 10.3950 ;
      LAYER M4  ;
        RECT 14.8610 10.0520 15.4970 10.0760 ;
      LAYER V3  ;
        RECT 15.2240 10.0520 15.2420 10.0760 ;
    END
  END wd[9]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0050 17.5365 30.3530 18.6300 ;
      RECT 0.0050 18.6165 30.3530 19.7100 ;
      RECT 0.0050 19.6965 30.3530 20.7900 ;
      RECT 0.0050 20.7765 30.3530 21.8700 ;
      RECT 0.0050 21.8565 30.3530 22.9500 ;
      RECT 0.0050 22.9365 30.3530 24.0300 ;
      RECT 0.0050 24.0165 30.3530 25.1100 ;
      RECT 0.0050 25.0965 30.3530 26.1900 ;
      RECT 0.0050 26.1765 30.3530 27.2700 ;
      RECT 0.0050 27.2565 30.3530 28.3500 ;
      RECT 0.0050 28.3365 30.3530 29.4300 ;
      RECT 0.0050 29.4165 30.3530 30.5100 ;
      RECT 0.0050 30.4965 30.3530 31.5900 ;
      RECT 0.0050 31.5765 30.3530 32.6700 ;
      RECT 0.0050 32.6565 30.3530 33.7500 ;
      RECT 0.0050 33.7365 30.3530 34.8300 ;
      RECT 0.0000 34.8535 30.3480 43.5070 ;
        RECT 0.0050 42.9435 30.3530 44.0370 ;
        RECT 0.0050 44.0235 30.3530 45.1170 ;
        RECT 0.0050 45.1035 30.3530 46.1970 ;
        RECT 0.0050 46.1835 30.3530 47.2770 ;
        RECT 0.0050 47.2635 30.3530 48.3570 ;
        RECT 0.0050 48.3435 30.3530 49.4370 ;
        RECT 0.0050 49.4235 30.3530 50.5170 ;
        RECT 0.0050 50.5035 30.3530 51.5970 ;
        RECT 0.0050 51.5835 30.3530 52.6770 ;
        RECT 0.0050 52.6635 30.3530 53.7570 ;
        RECT 0.0050 53.7435 30.3530 54.8370 ;
        RECT 0.0050 54.8235 30.3530 55.9170 ;
        RECT 0.0050 55.9035 30.3530 56.9970 ;
        RECT 0.0050 56.9835 30.3530 58.0770 ;
        RECT 0.0050 58.0635 30.3530 59.1570 ;
        RECT 0.0050 59.1435 30.3530 60.2370 ;
        RECT 0.0050 60.2235 30.3530 61.3170 ;
        RECT 0.0050 61.3035 30.3530 62.3970 ;
        RECT 0.0050 62.3835 30.3530 63.4770 ;
        RECT 0.0050 63.4635 30.3530 64.5570 ;
        RECT 0.0050 64.5435 30.3530 65.6370 ;
        RECT 0.0050 65.6235 30.3530 66.7170 ;
        RECT 0.0050 66.7035 30.3530 67.7970 ;
        RECT 0.0050 67.7835 30.3530 68.8770 ;
        RECT 0.0050 68.8635 30.3530 69.9570 ;
        RECT 0.0050 69.9435 30.3530 71.0370 ;
        RECT 0.0050 71.0235 30.3530 72.1170 ;
        RECT 0.0050 72.1035 30.3530 73.1970 ;
        RECT 0.0050 73.1835 30.3530 74.2770 ;
        RECT 0.0050 74.2635 30.3530 75.3570 ;
        RECT 0.0050 75.3435 30.3530 76.4370 ;
        RECT 0.0050 76.4235 30.3530 77.5170 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0050 17.5365 30.3530 18.6300 ;
      RECT 0.0050 18.6165 30.3530 19.7100 ;
      RECT 0.0050 19.6965 30.3530 20.7900 ;
      RECT 0.0050 20.7765 30.3530 21.8700 ;
      RECT 0.0050 21.8565 30.3530 22.9500 ;
      RECT 0.0050 22.9365 30.3530 24.0300 ;
      RECT 0.0050 24.0165 30.3530 25.1100 ;
      RECT 0.0050 25.0965 30.3530 26.1900 ;
      RECT 0.0050 26.1765 30.3530 27.2700 ;
      RECT 0.0050 27.2565 30.3530 28.3500 ;
      RECT 0.0050 28.3365 30.3530 29.4300 ;
      RECT 0.0050 29.4165 30.3530 30.5100 ;
      RECT 0.0050 30.4965 30.3530 31.5900 ;
      RECT 0.0050 31.5765 30.3530 32.6700 ;
      RECT 0.0050 32.6565 30.3530 33.7500 ;
      RECT 0.0050 33.7365 30.3530 34.8300 ;
      RECT 0.0000 34.8535 30.3480 43.5070 ;
        RECT 0.0050 42.9435 30.3530 44.0370 ;
        RECT 0.0050 44.0235 30.3530 45.1170 ;
        RECT 0.0050 45.1035 30.3530 46.1970 ;
        RECT 0.0050 46.1835 30.3530 47.2770 ;
        RECT 0.0050 47.2635 30.3530 48.3570 ;
        RECT 0.0050 48.3435 30.3530 49.4370 ;
        RECT 0.0050 49.4235 30.3530 50.5170 ;
        RECT 0.0050 50.5035 30.3530 51.5970 ;
        RECT 0.0050 51.5835 30.3530 52.6770 ;
        RECT 0.0050 52.6635 30.3530 53.7570 ;
        RECT 0.0050 53.7435 30.3530 54.8370 ;
        RECT 0.0050 54.8235 30.3530 55.9170 ;
        RECT 0.0050 55.9035 30.3530 56.9970 ;
        RECT 0.0050 56.9835 30.3530 58.0770 ;
        RECT 0.0050 58.0635 30.3530 59.1570 ;
        RECT 0.0050 59.1435 30.3530 60.2370 ;
        RECT 0.0050 60.2235 30.3530 61.3170 ;
        RECT 0.0050 61.3035 30.3530 62.3970 ;
        RECT 0.0050 62.3835 30.3530 63.4770 ;
        RECT 0.0050 63.4635 30.3530 64.5570 ;
        RECT 0.0050 64.5435 30.3530 65.6370 ;
        RECT 0.0050 65.6235 30.3530 66.7170 ;
        RECT 0.0050 66.7035 30.3530 67.7970 ;
        RECT 0.0050 67.7835 30.3530 68.8770 ;
        RECT 0.0050 68.8635 30.3530 69.9570 ;
        RECT 0.0050 69.9435 30.3530 71.0370 ;
        RECT 0.0050 71.0235 30.3530 72.1170 ;
        RECT 0.0050 72.1035 30.3530 73.1970 ;
        RECT 0.0050 73.1835 30.3530 74.2770 ;
        RECT 0.0050 74.2635 30.3530 75.3570 ;
        RECT 0.0050 75.3435 30.3530 76.4370 ;
        RECT 0.0050 76.4235 30.3530 77.5170 ;
  LAYER V1 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0050 17.5365 30.3530 18.6300 ;
      RECT 0.0050 18.6165 30.3530 19.7100 ;
      RECT 0.0050 19.6965 30.3530 20.7900 ;
      RECT 0.0050 20.7765 30.3530 21.8700 ;
      RECT 0.0050 21.8565 30.3530 22.9500 ;
      RECT 0.0050 22.9365 30.3530 24.0300 ;
      RECT 0.0050 24.0165 30.3530 25.1100 ;
      RECT 0.0050 25.0965 30.3530 26.1900 ;
      RECT 0.0050 26.1765 30.3530 27.2700 ;
      RECT 0.0050 27.2565 30.3530 28.3500 ;
      RECT 0.0050 28.3365 30.3530 29.4300 ;
      RECT 0.0050 29.4165 30.3530 30.5100 ;
      RECT 0.0050 30.4965 30.3530 31.5900 ;
      RECT 0.0050 31.5765 30.3530 32.6700 ;
      RECT 0.0050 32.6565 30.3530 33.7500 ;
      RECT 0.0050 33.7365 30.3530 34.8300 ;
      RECT 0.0000 34.8535 30.3480 43.5070 ;
        RECT 0.0050 42.9435 30.3530 44.0370 ;
        RECT 0.0050 44.0235 30.3530 45.1170 ;
        RECT 0.0050 45.1035 30.3530 46.1970 ;
        RECT 0.0050 46.1835 30.3530 47.2770 ;
        RECT 0.0050 47.2635 30.3530 48.3570 ;
        RECT 0.0050 48.3435 30.3530 49.4370 ;
        RECT 0.0050 49.4235 30.3530 50.5170 ;
        RECT 0.0050 50.5035 30.3530 51.5970 ;
        RECT 0.0050 51.5835 30.3530 52.6770 ;
        RECT 0.0050 52.6635 30.3530 53.7570 ;
        RECT 0.0050 53.7435 30.3530 54.8370 ;
        RECT 0.0050 54.8235 30.3530 55.9170 ;
        RECT 0.0050 55.9035 30.3530 56.9970 ;
        RECT 0.0050 56.9835 30.3530 58.0770 ;
        RECT 0.0050 58.0635 30.3530 59.1570 ;
        RECT 0.0050 59.1435 30.3530 60.2370 ;
        RECT 0.0050 60.2235 30.3530 61.3170 ;
        RECT 0.0050 61.3035 30.3530 62.3970 ;
        RECT 0.0050 62.3835 30.3530 63.4770 ;
        RECT 0.0050 63.4635 30.3530 64.5570 ;
        RECT 0.0050 64.5435 30.3530 65.6370 ;
        RECT 0.0050 65.6235 30.3530 66.7170 ;
        RECT 0.0050 66.7035 30.3530 67.7970 ;
        RECT 0.0050 67.7835 30.3530 68.8770 ;
        RECT 0.0050 68.8635 30.3530 69.9570 ;
        RECT 0.0050 69.9435 30.3530 71.0370 ;
        RECT 0.0050 71.0235 30.3530 72.1170 ;
        RECT 0.0050 72.1035 30.3530 73.1970 ;
        RECT 0.0050 73.1835 30.3530 74.2770 ;
        RECT 0.0050 74.2635 30.3530 75.3570 ;
        RECT 0.0050 75.3435 30.3530 76.4370 ;
        RECT 0.0050 76.4235 30.3530 77.5170 ;
  LAYER V2 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0050 11.0565 30.3530 12.1500 ;
      RECT 0.0050 12.1365 30.3530 13.2300 ;
      RECT 0.0050 13.2165 30.3530 14.3100 ;
      RECT 0.0050 14.2965 30.3530 15.3900 ;
      RECT 0.0050 15.3765 30.3530 16.4700 ;
      RECT 0.0050 16.4565 30.3530 17.5500 ;
      RECT 0.0050 17.5365 30.3530 18.6300 ;
      RECT 0.0050 18.6165 30.3530 19.7100 ;
      RECT 0.0050 19.6965 30.3530 20.7900 ;
      RECT 0.0050 20.7765 30.3530 21.8700 ;
      RECT 0.0050 21.8565 30.3530 22.9500 ;
      RECT 0.0050 22.9365 30.3530 24.0300 ;
      RECT 0.0050 24.0165 30.3530 25.1100 ;
      RECT 0.0050 25.0965 30.3530 26.1900 ;
      RECT 0.0050 26.1765 30.3530 27.2700 ;
      RECT 0.0050 27.2565 30.3530 28.3500 ;
      RECT 0.0050 28.3365 30.3530 29.4300 ;
      RECT 0.0050 29.4165 30.3530 30.5100 ;
      RECT 0.0050 30.4965 30.3530 31.5900 ;
      RECT 0.0050 31.5765 30.3530 32.6700 ;
      RECT 0.0050 32.6565 30.3530 33.7500 ;
      RECT 0.0050 33.7365 30.3530 34.8300 ;
      RECT 0.0000 34.8535 30.3480 43.5070 ;
        RECT 0.0050 42.9435 30.3530 44.0370 ;
        RECT 0.0050 44.0235 30.3530 45.1170 ;
        RECT 0.0050 45.1035 30.3530 46.1970 ;
        RECT 0.0050 46.1835 30.3530 47.2770 ;
        RECT 0.0050 47.2635 30.3530 48.3570 ;
        RECT 0.0050 48.3435 30.3530 49.4370 ;
        RECT 0.0050 49.4235 30.3530 50.5170 ;
        RECT 0.0050 50.5035 30.3530 51.5970 ;
        RECT 0.0050 51.5835 30.3530 52.6770 ;
        RECT 0.0050 52.6635 30.3530 53.7570 ;
        RECT 0.0050 53.7435 30.3530 54.8370 ;
        RECT 0.0050 54.8235 30.3530 55.9170 ;
        RECT 0.0050 55.9035 30.3530 56.9970 ;
        RECT 0.0050 56.9835 30.3530 58.0770 ;
        RECT 0.0050 58.0635 30.3530 59.1570 ;
        RECT 0.0050 59.1435 30.3530 60.2370 ;
        RECT 0.0050 60.2235 30.3530 61.3170 ;
        RECT 0.0050 61.3035 30.3530 62.3970 ;
        RECT 0.0050 62.3835 30.3530 63.4770 ;
        RECT 0.0050 63.4635 30.3530 64.5570 ;
        RECT 0.0050 64.5435 30.3530 65.6370 ;
        RECT 0.0050 65.6235 30.3530 66.7170 ;
        RECT 0.0050 66.7035 30.3530 67.7970 ;
        RECT 0.0050 67.7835 30.3530 68.8770 ;
        RECT 0.0050 68.8635 30.3530 69.9570 ;
        RECT 0.0050 69.9435 30.3530 71.0370 ;
        RECT 0.0050 71.0235 30.3530 72.1170 ;
        RECT 0.0050 72.1035 30.3530 73.1970 ;
        RECT 0.0050 73.1835 30.3530 74.2770 ;
        RECT 0.0050 74.2635 30.3530 75.3570 ;
        RECT 0.0050 75.3435 30.3530 76.4370 ;
        RECT 0.0050 76.4235 30.3530 77.5170 ;
  LAYER M3  ;
      RECT 15.6110 0.3450 15.6290 1.2805 ;
      RECT 15.5750 0.3450 15.5930 1.2805 ;
      RECT 15.5390 0.9220 15.5570 1.2445 ;
      RECT 15.4220 1.1190 15.4400 1.2285 ;
      RECT 15.4130 0.3775 15.4310 0.6170 ;
      RECT 15.3770 0.9585 15.3950 1.1120 ;
      RECT 15.2960 0.9840 15.3140 1.2420 ;
      RECT 14.7560 0.3450 14.7740 1.2805 ;
      RECT 14.7200 0.3450 14.7380 1.2805 ;
      RECT 14.6840 0.5260 14.7020 1.0940 ;
      RECT 15.6110 1.4250 15.6290 2.3605 ;
      RECT 15.5750 1.4250 15.5930 2.3605 ;
      RECT 15.5390 2.0020 15.5570 2.3245 ;
      RECT 15.4220 2.1990 15.4400 2.3085 ;
      RECT 15.4130 1.4575 15.4310 1.6970 ;
      RECT 15.3770 2.0385 15.3950 2.1920 ;
      RECT 15.2960 2.0640 15.3140 2.3220 ;
      RECT 14.7560 1.4250 14.7740 2.3605 ;
      RECT 14.7200 1.4250 14.7380 2.3605 ;
      RECT 14.6840 1.6060 14.7020 2.1740 ;
      RECT 15.6110 2.5050 15.6290 3.4405 ;
      RECT 15.5750 2.5050 15.5930 3.4405 ;
      RECT 15.5390 3.0820 15.5570 3.4045 ;
      RECT 15.4220 3.2790 15.4400 3.3885 ;
      RECT 15.4130 2.5375 15.4310 2.7770 ;
      RECT 15.3770 3.1185 15.3950 3.2720 ;
      RECT 15.2960 3.1440 15.3140 3.4020 ;
      RECT 14.7560 2.5050 14.7740 3.4405 ;
      RECT 14.7200 2.5050 14.7380 3.4405 ;
      RECT 14.6840 2.6860 14.7020 3.2540 ;
      RECT 15.6110 3.5850 15.6290 4.5205 ;
      RECT 15.5750 3.5850 15.5930 4.5205 ;
      RECT 15.5390 4.1620 15.5570 4.4845 ;
      RECT 15.4220 4.3590 15.4400 4.4685 ;
      RECT 15.4130 3.6175 15.4310 3.8570 ;
      RECT 15.3770 4.1985 15.3950 4.3520 ;
      RECT 15.2960 4.2240 15.3140 4.4820 ;
      RECT 14.7560 3.5850 14.7740 4.5205 ;
      RECT 14.7200 3.5850 14.7380 4.5205 ;
      RECT 14.6840 3.7660 14.7020 4.3340 ;
      RECT 15.6110 4.6650 15.6290 5.6005 ;
      RECT 15.5750 4.6650 15.5930 5.6005 ;
      RECT 15.5390 5.2420 15.5570 5.5645 ;
      RECT 15.4220 5.4390 15.4400 5.5485 ;
      RECT 15.4130 4.6975 15.4310 4.9370 ;
      RECT 15.3770 5.2785 15.3950 5.4320 ;
      RECT 15.2960 5.3040 15.3140 5.5620 ;
      RECT 14.7560 4.6650 14.7740 5.6005 ;
      RECT 14.7200 4.6650 14.7380 5.6005 ;
      RECT 14.6840 4.8460 14.7020 5.4140 ;
      RECT 15.6110 5.7450 15.6290 6.6805 ;
      RECT 15.5750 5.7450 15.5930 6.6805 ;
      RECT 15.5390 6.3220 15.5570 6.6445 ;
      RECT 15.4220 6.5190 15.4400 6.6285 ;
      RECT 15.4130 5.7775 15.4310 6.0170 ;
      RECT 15.3770 6.3585 15.3950 6.5120 ;
      RECT 15.2960 6.3840 15.3140 6.6420 ;
      RECT 14.7560 5.7450 14.7740 6.6805 ;
      RECT 14.7200 5.7450 14.7380 6.6805 ;
      RECT 14.6840 5.9260 14.7020 6.4940 ;
      RECT 15.6110 6.8250 15.6290 7.7605 ;
      RECT 15.5750 6.8250 15.5930 7.7605 ;
      RECT 15.5390 7.4020 15.5570 7.7245 ;
      RECT 15.4220 7.5990 15.4400 7.7085 ;
      RECT 15.4130 6.8575 15.4310 7.0970 ;
      RECT 15.3770 7.4385 15.3950 7.5920 ;
      RECT 15.2960 7.4640 15.3140 7.7220 ;
      RECT 14.7560 6.8250 14.7740 7.7605 ;
      RECT 14.7200 6.8250 14.7380 7.7605 ;
      RECT 14.6840 7.0060 14.7020 7.5740 ;
      RECT 15.6110 7.9050 15.6290 8.8405 ;
      RECT 15.5750 7.9050 15.5930 8.8405 ;
      RECT 15.5390 8.4820 15.5570 8.8045 ;
      RECT 15.4220 8.6790 15.4400 8.7885 ;
      RECT 15.4130 7.9375 15.4310 8.1770 ;
      RECT 15.3770 8.5185 15.3950 8.6720 ;
      RECT 15.2960 8.5440 15.3140 8.8020 ;
      RECT 14.7560 7.9050 14.7740 8.8405 ;
      RECT 14.7200 7.9050 14.7380 8.8405 ;
      RECT 14.6840 8.0860 14.7020 8.6540 ;
      RECT 15.6110 8.9850 15.6290 9.9205 ;
      RECT 15.5750 8.9850 15.5930 9.9205 ;
      RECT 15.5390 9.5620 15.5570 9.8845 ;
      RECT 15.4220 9.7590 15.4400 9.8685 ;
      RECT 15.4130 9.0175 15.4310 9.2570 ;
      RECT 15.3770 9.5985 15.3950 9.7520 ;
      RECT 15.2960 9.6240 15.3140 9.8820 ;
      RECT 14.7560 8.9850 14.7740 9.9205 ;
      RECT 14.7200 8.9850 14.7380 9.9205 ;
      RECT 14.6840 9.1660 14.7020 9.7340 ;
      RECT 15.6110 10.0650 15.6290 11.0005 ;
      RECT 15.5750 10.0650 15.5930 11.0005 ;
      RECT 15.5390 10.6420 15.5570 10.9645 ;
      RECT 15.4220 10.8390 15.4400 10.9485 ;
      RECT 15.4130 10.0975 15.4310 10.3370 ;
      RECT 15.3770 10.6785 15.3950 10.8320 ;
      RECT 15.2960 10.7040 15.3140 10.9620 ;
      RECT 14.7560 10.0650 14.7740 11.0005 ;
      RECT 14.7200 10.0650 14.7380 11.0005 ;
      RECT 14.6840 10.2460 14.7020 10.8140 ;
      RECT 15.6110 11.1450 15.6290 12.0805 ;
      RECT 15.5750 11.1450 15.5930 12.0805 ;
      RECT 15.5390 11.7220 15.5570 12.0445 ;
      RECT 15.4220 11.9190 15.4400 12.0285 ;
      RECT 15.4130 11.1775 15.4310 11.4170 ;
      RECT 15.3770 11.7585 15.3950 11.9120 ;
      RECT 15.2960 11.7840 15.3140 12.0420 ;
      RECT 14.7560 11.1450 14.7740 12.0805 ;
      RECT 14.7200 11.1450 14.7380 12.0805 ;
      RECT 14.6840 11.3260 14.7020 11.8940 ;
      RECT 15.6110 12.2250 15.6290 13.1605 ;
      RECT 15.5750 12.2250 15.5930 13.1605 ;
      RECT 15.5390 12.8020 15.5570 13.1245 ;
      RECT 15.4220 12.9990 15.4400 13.1085 ;
      RECT 15.4130 12.2575 15.4310 12.4970 ;
      RECT 15.3770 12.8385 15.3950 12.9920 ;
      RECT 15.2960 12.8640 15.3140 13.1220 ;
      RECT 14.7560 12.2250 14.7740 13.1605 ;
      RECT 14.7200 12.2250 14.7380 13.1605 ;
      RECT 14.6840 12.4060 14.7020 12.9740 ;
      RECT 15.6110 13.3050 15.6290 14.2405 ;
      RECT 15.5750 13.3050 15.5930 14.2405 ;
      RECT 15.5390 13.8820 15.5570 14.2045 ;
      RECT 15.4220 14.0790 15.4400 14.1885 ;
      RECT 15.4130 13.3375 15.4310 13.5770 ;
      RECT 15.3770 13.9185 15.3950 14.0720 ;
      RECT 15.2960 13.9440 15.3140 14.2020 ;
      RECT 14.7560 13.3050 14.7740 14.2405 ;
      RECT 14.7200 13.3050 14.7380 14.2405 ;
      RECT 14.6840 13.4860 14.7020 14.0540 ;
      RECT 15.6110 14.3850 15.6290 15.3205 ;
      RECT 15.5750 14.3850 15.5930 15.3205 ;
      RECT 15.5390 14.9620 15.5570 15.2845 ;
      RECT 15.4220 15.1590 15.4400 15.2685 ;
      RECT 15.4130 14.4175 15.4310 14.6570 ;
      RECT 15.3770 14.9985 15.3950 15.1520 ;
      RECT 15.2960 15.0240 15.3140 15.2820 ;
      RECT 14.7560 14.3850 14.7740 15.3205 ;
      RECT 14.7200 14.3850 14.7380 15.3205 ;
      RECT 14.6840 14.5660 14.7020 15.1340 ;
      RECT 15.6110 15.4650 15.6290 16.4005 ;
      RECT 15.5750 15.4650 15.5930 16.4005 ;
      RECT 15.5390 16.0420 15.5570 16.3645 ;
      RECT 15.4220 16.2390 15.4400 16.3485 ;
      RECT 15.4130 15.4975 15.4310 15.7370 ;
      RECT 15.3770 16.0785 15.3950 16.2320 ;
      RECT 15.2960 16.1040 15.3140 16.3620 ;
      RECT 14.7560 15.4650 14.7740 16.4005 ;
      RECT 14.7200 15.4650 14.7380 16.4005 ;
      RECT 14.6840 15.6460 14.7020 16.2140 ;
      RECT 15.6110 16.5450 15.6290 17.4805 ;
      RECT 15.5750 16.5450 15.5930 17.4805 ;
      RECT 15.5390 17.1220 15.5570 17.4445 ;
      RECT 15.4220 17.3190 15.4400 17.4285 ;
      RECT 15.4130 16.5775 15.4310 16.8170 ;
      RECT 15.3770 17.1585 15.3950 17.3120 ;
      RECT 15.2960 17.1840 15.3140 17.4420 ;
      RECT 14.7560 16.5450 14.7740 17.4805 ;
      RECT 14.7200 16.5450 14.7380 17.4805 ;
      RECT 14.6840 16.7260 14.7020 17.2940 ;
      RECT 15.6110 17.6250 15.6290 18.5605 ;
      RECT 15.5750 17.6250 15.5930 18.5605 ;
      RECT 15.5390 18.2020 15.5570 18.5245 ;
      RECT 15.4220 18.3990 15.4400 18.5085 ;
      RECT 15.4130 17.6575 15.4310 17.8970 ;
      RECT 15.3770 18.2385 15.3950 18.3920 ;
      RECT 15.2960 18.2640 15.3140 18.5220 ;
      RECT 14.7560 17.6250 14.7740 18.5605 ;
      RECT 14.7200 17.6250 14.7380 18.5605 ;
      RECT 14.6840 17.8060 14.7020 18.3740 ;
      RECT 15.6110 18.7050 15.6290 19.6405 ;
      RECT 15.5750 18.7050 15.5930 19.6405 ;
      RECT 15.5390 19.2820 15.5570 19.6045 ;
      RECT 15.4220 19.4790 15.4400 19.5885 ;
      RECT 15.4130 18.7375 15.4310 18.9770 ;
      RECT 15.3770 19.3185 15.3950 19.4720 ;
      RECT 15.2960 19.3440 15.3140 19.6020 ;
      RECT 14.7560 18.7050 14.7740 19.6405 ;
      RECT 14.7200 18.7050 14.7380 19.6405 ;
      RECT 14.6840 18.8860 14.7020 19.4540 ;
      RECT 15.6110 19.7850 15.6290 20.7205 ;
      RECT 15.5750 19.7850 15.5930 20.7205 ;
      RECT 15.5390 20.3620 15.5570 20.6845 ;
      RECT 15.4220 20.5590 15.4400 20.6685 ;
      RECT 15.4130 19.8175 15.4310 20.0570 ;
      RECT 15.3770 20.3985 15.3950 20.5520 ;
      RECT 15.2960 20.4240 15.3140 20.6820 ;
      RECT 14.7560 19.7850 14.7740 20.7205 ;
      RECT 14.7200 19.7850 14.7380 20.7205 ;
      RECT 14.6840 19.9660 14.7020 20.5340 ;
      RECT 15.6110 20.8650 15.6290 21.8005 ;
      RECT 15.5750 20.8650 15.5930 21.8005 ;
      RECT 15.5390 21.4420 15.5570 21.7645 ;
      RECT 15.4220 21.6390 15.4400 21.7485 ;
      RECT 15.4130 20.8975 15.4310 21.1370 ;
      RECT 15.3770 21.4785 15.3950 21.6320 ;
      RECT 15.2960 21.5040 15.3140 21.7620 ;
      RECT 14.7560 20.8650 14.7740 21.8005 ;
      RECT 14.7200 20.8650 14.7380 21.8005 ;
      RECT 14.6840 21.0460 14.7020 21.6140 ;
      RECT 15.6110 21.9450 15.6290 22.8805 ;
      RECT 15.5750 21.9450 15.5930 22.8805 ;
      RECT 15.5390 22.5220 15.5570 22.8445 ;
      RECT 15.4220 22.7190 15.4400 22.8285 ;
      RECT 15.4130 21.9775 15.4310 22.2170 ;
      RECT 15.3770 22.5585 15.3950 22.7120 ;
      RECT 15.2960 22.5840 15.3140 22.8420 ;
      RECT 14.7560 21.9450 14.7740 22.8805 ;
      RECT 14.7200 21.9450 14.7380 22.8805 ;
      RECT 14.6840 22.1260 14.7020 22.6940 ;
      RECT 15.6110 23.0250 15.6290 23.9605 ;
      RECT 15.5750 23.0250 15.5930 23.9605 ;
      RECT 15.5390 23.6020 15.5570 23.9245 ;
      RECT 15.4220 23.7990 15.4400 23.9085 ;
      RECT 15.4130 23.0575 15.4310 23.2970 ;
      RECT 15.3770 23.6385 15.3950 23.7920 ;
      RECT 15.2960 23.6640 15.3140 23.9220 ;
      RECT 14.7560 23.0250 14.7740 23.9605 ;
      RECT 14.7200 23.0250 14.7380 23.9605 ;
      RECT 14.6840 23.2060 14.7020 23.7740 ;
      RECT 15.6110 24.1050 15.6290 25.0405 ;
      RECT 15.5750 24.1050 15.5930 25.0405 ;
      RECT 15.5390 24.6820 15.5570 25.0045 ;
      RECT 15.4220 24.8790 15.4400 24.9885 ;
      RECT 15.4130 24.1375 15.4310 24.3770 ;
      RECT 15.3770 24.7185 15.3950 24.8720 ;
      RECT 15.2960 24.7440 15.3140 25.0020 ;
      RECT 14.7560 24.1050 14.7740 25.0405 ;
      RECT 14.7200 24.1050 14.7380 25.0405 ;
      RECT 14.6840 24.2860 14.7020 24.8540 ;
      RECT 15.6110 25.1850 15.6290 26.1205 ;
      RECT 15.5750 25.1850 15.5930 26.1205 ;
      RECT 15.5390 25.7620 15.5570 26.0845 ;
      RECT 15.4220 25.9590 15.4400 26.0685 ;
      RECT 15.4130 25.2175 15.4310 25.4570 ;
      RECT 15.3770 25.7985 15.3950 25.9520 ;
      RECT 15.2960 25.8240 15.3140 26.0820 ;
      RECT 14.7560 25.1850 14.7740 26.1205 ;
      RECT 14.7200 25.1850 14.7380 26.1205 ;
      RECT 14.6840 25.3660 14.7020 25.9340 ;
      RECT 15.6110 26.2650 15.6290 27.2005 ;
      RECT 15.5750 26.2650 15.5930 27.2005 ;
      RECT 15.5390 26.8420 15.5570 27.1645 ;
      RECT 15.4220 27.0390 15.4400 27.1485 ;
      RECT 15.4130 26.2975 15.4310 26.5370 ;
      RECT 15.3770 26.8785 15.3950 27.0320 ;
      RECT 15.2960 26.9040 15.3140 27.1620 ;
      RECT 14.7560 26.2650 14.7740 27.2005 ;
      RECT 14.7200 26.2650 14.7380 27.2005 ;
      RECT 14.6840 26.4460 14.7020 27.0140 ;
      RECT 15.6110 27.3450 15.6290 28.2805 ;
      RECT 15.5750 27.3450 15.5930 28.2805 ;
      RECT 15.5390 27.9220 15.5570 28.2445 ;
      RECT 15.4220 28.1190 15.4400 28.2285 ;
      RECT 15.4130 27.3775 15.4310 27.6170 ;
      RECT 15.3770 27.9585 15.3950 28.1120 ;
      RECT 15.2960 27.9840 15.3140 28.2420 ;
      RECT 14.7560 27.3450 14.7740 28.2805 ;
      RECT 14.7200 27.3450 14.7380 28.2805 ;
      RECT 14.6840 27.5260 14.7020 28.0940 ;
      RECT 15.6110 28.4250 15.6290 29.3605 ;
      RECT 15.5750 28.4250 15.5930 29.3605 ;
      RECT 15.5390 29.0020 15.5570 29.3245 ;
      RECT 15.4220 29.1990 15.4400 29.3085 ;
      RECT 15.4130 28.4575 15.4310 28.6970 ;
      RECT 15.3770 29.0385 15.3950 29.1920 ;
      RECT 15.2960 29.0640 15.3140 29.3220 ;
      RECT 14.7560 28.4250 14.7740 29.3605 ;
      RECT 14.7200 28.4250 14.7380 29.3605 ;
      RECT 14.6840 28.6060 14.7020 29.1740 ;
      RECT 15.6110 29.5050 15.6290 30.4405 ;
      RECT 15.5750 29.5050 15.5930 30.4405 ;
      RECT 15.5390 30.0820 15.5570 30.4045 ;
      RECT 15.4220 30.2790 15.4400 30.3885 ;
      RECT 15.4130 29.5375 15.4310 29.7770 ;
      RECT 15.3770 30.1185 15.3950 30.2720 ;
      RECT 15.2960 30.1440 15.3140 30.4020 ;
      RECT 14.7560 29.5050 14.7740 30.4405 ;
      RECT 14.7200 29.5050 14.7380 30.4405 ;
      RECT 14.6840 29.6860 14.7020 30.2540 ;
      RECT 15.6110 30.5850 15.6290 31.5205 ;
      RECT 15.5750 30.5850 15.5930 31.5205 ;
      RECT 15.5390 31.1620 15.5570 31.4845 ;
      RECT 15.4220 31.3590 15.4400 31.4685 ;
      RECT 15.4130 30.6175 15.4310 30.8570 ;
      RECT 15.3770 31.1985 15.3950 31.3520 ;
      RECT 15.2960 31.2240 15.3140 31.4820 ;
      RECT 14.7560 30.5850 14.7740 31.5205 ;
      RECT 14.7200 30.5850 14.7380 31.5205 ;
      RECT 14.6840 30.7660 14.7020 31.3340 ;
      RECT 15.6110 31.6650 15.6290 32.6005 ;
      RECT 15.5750 31.6650 15.5930 32.6005 ;
      RECT 15.5390 32.2420 15.5570 32.5645 ;
      RECT 15.4220 32.4390 15.4400 32.5485 ;
      RECT 15.4130 31.6975 15.4310 31.9370 ;
      RECT 15.3770 32.2785 15.3950 32.4320 ;
      RECT 15.2960 32.3040 15.3140 32.5620 ;
      RECT 14.7560 31.6650 14.7740 32.6005 ;
      RECT 14.7200 31.6650 14.7380 32.6005 ;
      RECT 14.6840 31.8460 14.7020 32.4140 ;
      RECT 15.6110 32.7450 15.6290 33.6805 ;
      RECT 15.5750 32.7450 15.5930 33.6805 ;
      RECT 15.5390 33.3220 15.5570 33.6445 ;
      RECT 15.4220 33.5190 15.4400 33.6285 ;
      RECT 15.4130 32.7775 15.4310 33.0170 ;
      RECT 15.3770 33.3585 15.3950 33.5120 ;
      RECT 15.2960 33.3840 15.3140 33.6420 ;
      RECT 14.7560 32.7450 14.7740 33.6805 ;
      RECT 14.7200 32.7450 14.7380 33.6805 ;
      RECT 14.6840 32.9260 14.7020 33.4940 ;
      RECT 15.6110 33.8250 15.6290 34.7605 ;
      RECT 15.5750 33.8250 15.5930 34.7605 ;
      RECT 15.5390 34.4020 15.5570 34.7245 ;
      RECT 15.4220 34.5990 15.4400 34.7085 ;
      RECT 15.4130 33.8575 15.4310 34.0970 ;
      RECT 15.3770 34.4385 15.3950 34.5920 ;
      RECT 15.2960 34.4640 15.3140 34.7220 ;
      RECT 14.7560 33.8250 14.7740 34.7605 ;
      RECT 14.7200 33.8250 14.7380 34.7605 ;
      RECT 14.6840 34.0060 14.7020 34.5740 ;
      RECT 30.2130 34.6635 30.2310 43.0340 ;
      RECT 30.1770 34.6635 30.1950 43.0340 ;
      RECT 30.0690 34.6635 30.0870 38.4045 ;
      RECT 29.9610 34.6635 29.9790 38.4045 ;
      RECT 29.8530 34.6635 29.8710 38.4045 ;
      RECT 29.7450 34.6635 29.7630 38.4045 ;
      RECT 29.6370 34.6635 29.6550 38.4045 ;
      RECT 29.5290 34.6635 29.5470 38.4045 ;
      RECT 29.4210 34.6635 29.4390 38.4045 ;
      RECT 29.3130 34.6635 29.3310 38.4045 ;
      RECT 29.2050 34.6635 29.2230 38.4045 ;
      RECT 29.0970 34.6635 29.1150 38.4045 ;
      RECT 28.9890 34.6635 29.0070 38.4045 ;
      RECT 28.8810 34.6635 28.8990 38.4045 ;
      RECT 28.7730 34.6635 28.7910 38.4045 ;
      RECT 28.6650 34.6635 28.6830 38.4045 ;
      RECT 28.5570 34.6635 28.5750 38.4045 ;
      RECT 28.4490 34.6635 28.4670 38.4045 ;
      RECT 28.3410 34.6635 28.3590 38.4045 ;
      RECT 28.2330 34.6635 28.2510 38.4045 ;
      RECT 28.1250 34.6635 28.1430 38.4045 ;
      RECT 28.0170 34.6635 28.0350 38.4045 ;
      RECT 27.9090 34.6635 27.9270 38.4045 ;
      RECT 27.8010 34.6635 27.8190 38.4045 ;
      RECT 27.6930 34.6635 27.7110 38.4045 ;
      RECT 27.5850 34.6635 27.6030 38.4045 ;
      RECT 27.4770 34.6635 27.4950 38.4045 ;
      RECT 27.3690 34.6635 27.3870 38.4045 ;
      RECT 27.2610 34.6635 27.2790 38.4045 ;
      RECT 27.1530 34.6635 27.1710 38.4045 ;
      RECT 27.0450 34.6635 27.0630 38.4045 ;
      RECT 26.9370 34.6635 26.9550 38.4045 ;
      RECT 26.8290 34.6635 26.8470 38.4045 ;
      RECT 26.7210 34.6635 26.7390 38.4045 ;
      RECT 26.6130 34.6635 26.6310 38.4045 ;
      RECT 26.5050 34.6635 26.5230 38.4045 ;
      RECT 26.3970 34.6635 26.4150 38.4045 ;
      RECT 26.2890 34.6635 26.3070 38.4045 ;
      RECT 26.1810 34.6635 26.1990 38.4045 ;
      RECT 26.0730 34.6635 26.0910 38.4045 ;
      RECT 25.9650 34.6635 25.9830 38.4045 ;
      RECT 25.8570 34.6635 25.8750 38.4045 ;
      RECT 25.7490 34.6635 25.7670 38.4045 ;
      RECT 25.6410 34.6635 25.6590 38.4045 ;
      RECT 25.5330 34.6635 25.5510 38.4045 ;
      RECT 25.4250 34.6635 25.4430 38.4045 ;
      RECT 25.3170 34.6635 25.3350 38.4045 ;
      RECT 25.2090 34.6635 25.2270 38.4045 ;
      RECT 25.1010 34.6635 25.1190 38.4045 ;
      RECT 24.9930 34.6635 25.0110 38.4045 ;
      RECT 24.8850 34.6635 24.9030 38.4045 ;
      RECT 24.7770 34.6635 24.7950 38.4045 ;
      RECT 24.6690 34.6635 24.6870 38.4045 ;
      RECT 24.5610 34.6635 24.5790 38.4045 ;
      RECT 24.4530 34.6635 24.4710 38.4045 ;
      RECT 24.3450 34.6635 24.3630 38.4045 ;
      RECT 24.2370 34.6635 24.2550 38.4045 ;
      RECT 24.1290 34.6635 24.1470 38.4045 ;
      RECT 24.0210 34.6635 24.0390 38.4045 ;
      RECT 23.9130 34.6635 23.9310 38.4045 ;
      RECT 23.8050 34.6635 23.8230 38.4045 ;
      RECT 23.6970 34.6635 23.7150 38.4045 ;
      RECT 23.5890 34.6635 23.6070 38.4045 ;
      RECT 23.4810 34.6635 23.4990 38.4045 ;
      RECT 23.3730 34.6635 23.3910 38.4045 ;
      RECT 23.2650 34.6635 23.2830 38.4045 ;
      RECT 23.1570 34.6635 23.1750 38.4045 ;
      RECT 23.0490 34.6635 23.0670 38.4045 ;
      RECT 22.9410 34.6635 22.9590 38.4045 ;
      RECT 22.8330 34.6635 22.8510 38.4045 ;
      RECT 22.7250 34.6635 22.7430 38.4045 ;
      RECT 22.6170 34.6635 22.6350 38.4045 ;
      RECT 22.5090 34.6635 22.5270 38.4045 ;
      RECT 22.4010 34.6635 22.4190 38.4045 ;
      RECT 22.2930 34.6635 22.3110 38.4045 ;
      RECT 22.1850 34.6635 22.2030 38.4045 ;
      RECT 22.0770 34.6635 22.0950 38.4045 ;
      RECT 21.9690 34.6635 21.9870 38.4045 ;
      RECT 21.8610 34.6635 21.8790 38.4045 ;
      RECT 21.7530 34.6635 21.7710 38.4045 ;
      RECT 21.6450 34.6635 21.6630 38.4045 ;
      RECT 21.5370 34.6635 21.5550 38.4045 ;
      RECT 21.4290 34.6635 21.4470 38.4045 ;
      RECT 21.3210 34.6635 21.3390 38.4045 ;
      RECT 21.2130 34.6635 21.2310 38.4045 ;
      RECT 21.1050 34.6635 21.1230 38.4045 ;
      RECT 20.9970 34.6635 21.0150 38.4045 ;
      RECT 20.8890 34.6635 20.9070 38.4045 ;
      RECT 20.7810 34.6635 20.7990 38.4045 ;
      RECT 20.6730 34.6635 20.6910 38.4045 ;
      RECT 20.5650 34.6635 20.5830 38.4045 ;
      RECT 20.4570 34.6635 20.4750 38.4045 ;
      RECT 20.3490 34.6635 20.3670 38.4045 ;
      RECT 20.2410 34.6635 20.2590 38.4045 ;
      RECT 20.1330 34.6635 20.1510 38.4045 ;
      RECT 20.0250 34.6635 20.0430 38.4045 ;
      RECT 19.9170 34.6635 19.9350 38.4045 ;
      RECT 19.8090 34.8270 19.8270 35.1770 ;
      RECT 19.7010 34.6635 19.7190 38.4045 ;
      RECT 19.5930 34.6635 19.6110 38.4045 ;
      RECT 19.4850 34.6635 19.5030 38.4045 ;
      RECT 19.3770 34.6635 19.3950 38.4045 ;
      RECT 19.2690 34.6635 19.2870 38.4045 ;
      RECT 19.1610 34.6635 19.1790 38.4045 ;
      RECT 19.0530 34.6635 19.0710 38.4045 ;
      RECT 18.9450 34.6635 18.9630 38.4045 ;
      RECT 18.8370 34.6635 18.8550 38.4045 ;
      RECT 18.7290 34.6635 18.7470 38.4045 ;
      RECT 18.6210 34.6635 18.6390 38.4045 ;
      RECT 18.5130 34.6635 18.5310 38.4045 ;
      RECT 18.4050 34.6635 18.4230 38.4045 ;
      RECT 18.2970 34.6635 18.3150 38.4045 ;
      RECT 18.1890 34.6635 18.2070 38.4045 ;
      RECT 18.0810 34.6635 18.0990 38.4045 ;
      RECT 17.9730 34.6635 17.9910 38.4045 ;
      RECT 17.8650 34.6635 17.8830 38.4045 ;
      RECT 17.7570 34.6635 17.7750 38.4045 ;
      RECT 17.6490 34.6635 17.6670 38.4045 ;
      RECT 17.5410 34.6635 17.5590 38.4045 ;
      RECT 17.4330 34.6635 17.4510 38.4045 ;
      RECT 17.3250 34.6635 17.3430 38.4045 ;
      RECT 17.2170 34.6635 17.2350 38.4045 ;
      RECT 17.1090 34.6635 17.1270 38.4045 ;
      RECT 17.0010 34.6635 17.0190 38.4045 ;
      RECT 16.8930 34.6635 16.9110 38.4045 ;
      RECT 16.7850 34.6635 16.8030 38.4045 ;
      RECT 16.6770 34.6635 16.6950 38.4045 ;
      RECT 16.5690 34.6635 16.5870 38.4045 ;
      RECT 16.4610 34.6635 16.4790 38.4045 ;
      RECT 16.4250 38.6155 16.4430 39.3202 ;
      RECT 16.4250 40.0585 16.4430 41.2195 ;
      RECT 16.4070 35.4875 16.4250 36.1635 ;
      RECT 16.4070 36.9095 16.4250 37.2075 ;
      RECT 16.4070 38.0255 16.4250 38.2875 ;
      RECT 16.3890 38.6790 16.4070 39.3690 ;
      RECT 16.3890 39.4200 16.4070 40.4055 ;
      RECT 16.3890 40.4465 16.4070 41.0635 ;
      RECT 16.3530 34.6635 16.3710 43.0340 ;
      RECT 16.3170 38.9515 16.3350 39.0345 ;
      RECT 16.2990 35.5955 16.3170 36.2265 ;
      RECT 16.2990 36.6395 16.3170 36.8295 ;
      RECT 16.2990 37.5215 16.3170 37.5705 ;
      RECT 16.2990 38.2535 16.3170 38.2905 ;
      RECT 16.2810 38.6465 16.2990 42.2395 ;
      RECT 16.1910 34.8600 16.2090 34.9980 ;
      RECT 16.1910 35.2175 16.2090 36.0195 ;
      RECT 16.1910 36.5675 16.2090 37.1355 ;
      RECT 16.1910 38.6465 16.2090 42.2395 ;
      RECT 16.1550 36.6395 16.1730 37.0095 ;
      RECT 16.1190 35.9915 16.1370 36.1275 ;
      RECT 16.1190 36.9815 16.1370 37.2075 ;
      RECT 16.1190 38.2235 16.1370 38.2875 ;
      RECT 16.0830 36.0935 16.1010 36.1305 ;
      RECT 16.0830 37.7195 16.1010 37.7625 ;
      RECT 16.0830 38.2535 16.1010 38.2905 ;
      RECT 16.0470 36.4055 16.0650 36.9015 ;
      RECT 16.0470 36.9455 16.0650 37.1355 ;
      RECT 16.0470 37.9055 16.0650 38.2155 ;
      RECT 16.0110 36.2975 16.0290 37.5445 ;
      RECT 15.0390 34.8535 15.0570 35.0075 ;
      RECT 15.0030 34.8535 15.0210 34.9035 ;
      RECT 14.9310 34.8535 14.9490 34.9250 ;
      RECT 14.2830 35.9915 14.3010 36.3975 ;
      RECT 14.2470 37.1015 14.2650 37.1385 ;
      RECT 14.2110 36.0275 14.2290 36.6315 ;
      RECT 14.1750 35.8655 14.1930 35.9295 ;
      RECT 14.1390 34.9065 14.1570 34.9575 ;
      RECT 14.1390 38.0255 14.1570 38.2155 ;
      RECT 14.1390 38.6465 14.1570 42.2395 ;
      RECT 14.0310 35.3255 14.0490 35.5155 ;
      RECT 14.0310 36.0995 14.0490 38.3595 ;
      RECT 14.0130 38.9515 14.0310 39.0345 ;
      RECT 13.9770 34.8270 13.9950 43.0340 ;
      RECT 13.9410 38.6790 13.9590 39.3690 ;
      RECT 13.9410 39.4200 13.9590 40.4055 ;
      RECT 13.9410 40.4465 13.9590 41.0635 ;
      RECT 13.9230 35.3255 13.9410 35.8215 ;
      RECT 13.9230 36.6035 13.9410 37.1715 ;
      RECT 13.9230 37.4855 13.9410 38.2155 ;
      RECT 13.9050 38.6155 13.9230 39.3202 ;
      RECT 13.9050 40.0585 13.9230 41.2195 ;
      RECT 13.8690 34.8270 13.8870 35.1770 ;
      RECT 13.8690 38.3710 13.8870 43.0340 ;
      RECT 13.7610 34.8270 13.7790 35.1770 ;
      RECT 13.6530 34.8270 13.6710 35.1770 ;
      RECT 13.5450 34.8270 13.5630 35.1770 ;
      RECT 13.4370 34.8270 13.4550 35.1770 ;
      RECT 13.3290 34.8270 13.3470 35.1770 ;
      RECT 13.2210 34.8270 13.2390 35.1770 ;
      RECT 13.1130 34.8270 13.1310 35.1770 ;
      RECT 13.0050 34.8270 13.0230 35.1770 ;
      RECT 12.8970 34.8270 12.9150 35.1770 ;
      RECT 12.7890 34.8270 12.8070 35.1770 ;
      RECT 12.6810 34.8270 12.6990 35.1770 ;
      RECT 12.5730 34.8270 12.5910 35.1770 ;
      RECT 12.4650 34.8270 12.4830 35.1770 ;
      RECT 12.3570 34.8270 12.3750 35.1770 ;
      RECT 12.2490 34.8270 12.2670 35.1770 ;
      RECT 12.1410 34.8270 12.1590 35.1770 ;
      RECT 12.0330 34.8270 12.0510 35.1770 ;
      RECT 11.9250 34.8270 11.9430 35.1770 ;
      RECT 11.8170 34.8270 11.8350 35.1770 ;
      RECT 11.7090 34.8270 11.7270 35.1770 ;
      RECT 11.6010 34.8270 11.6190 35.1770 ;
      RECT 11.4930 34.8270 11.5110 35.1770 ;
      RECT 11.3850 34.8270 11.4030 35.1770 ;
      RECT 11.2770 34.8270 11.2950 35.1770 ;
      RECT 11.1690 34.8270 11.1870 35.1770 ;
      RECT 11.0610 34.8270 11.0790 35.1770 ;
      RECT 10.9530 34.8270 10.9710 35.1770 ;
      RECT 10.8450 34.8270 10.8630 35.1770 ;
      RECT 10.7370 34.8270 10.7550 35.1770 ;
      RECT 10.6290 34.8270 10.6470 35.1770 ;
      RECT 10.5210 34.8270 10.5390 35.1770 ;
      RECT 10.4130 34.8270 10.4310 35.1770 ;
      RECT 10.3050 34.8270 10.3230 35.1770 ;
      RECT 10.1970 34.8270 10.2150 35.1770 ;
      RECT 10.0890 34.8270 10.1070 35.1770 ;
      RECT 9.9810 34.8270 9.9990 35.1770 ;
      RECT 9.8730 34.8270 9.8910 35.1770 ;
      RECT 9.7650 34.8270 9.7830 35.1770 ;
      RECT 9.6570 34.8270 9.6750 35.1770 ;
      RECT 9.5490 34.8270 9.5670 35.1770 ;
      RECT 9.4410 34.8270 9.4590 35.1770 ;
      RECT 9.3330 34.8270 9.3510 35.1770 ;
      RECT 9.2250 34.8270 9.2430 35.1770 ;
      RECT 9.1170 34.8270 9.1350 35.1770 ;
      RECT 9.0090 34.8270 9.0270 35.1770 ;
      RECT 8.9010 34.8270 8.9190 35.1770 ;
      RECT 8.7930 34.8270 8.8110 35.1770 ;
      RECT 8.6850 34.8270 8.7030 35.1770 ;
      RECT 8.5770 34.8270 8.5950 35.1770 ;
      RECT 8.4690 34.8270 8.4870 35.1770 ;
      RECT 8.3610 34.8270 8.3790 35.1770 ;
      RECT 8.2530 34.8270 8.2710 35.1770 ;
      RECT 8.1450 34.8270 8.1630 35.1770 ;
      RECT 8.0370 34.8270 8.0550 35.1770 ;
      RECT 7.9290 34.8270 7.9470 35.1770 ;
      RECT 7.8210 34.8270 7.8390 35.1770 ;
      RECT 7.7130 34.8270 7.7310 35.1770 ;
      RECT 7.6050 34.8270 7.6230 35.1770 ;
      RECT 7.4970 34.8270 7.5150 35.1770 ;
      RECT 7.3890 34.8270 7.4070 35.1770 ;
      RECT 7.2810 34.8270 7.2990 35.1770 ;
      RECT 7.1730 34.8270 7.1910 35.1770 ;
      RECT 7.0650 34.8270 7.0830 35.1770 ;
      RECT 6.9570 34.8270 6.9750 35.1770 ;
      RECT 6.8490 34.8270 6.8670 35.1770 ;
      RECT 6.7410 34.8270 6.7590 35.1770 ;
      RECT 6.6330 34.8270 6.6510 35.1770 ;
      RECT 6.5250 34.8270 6.5430 35.1770 ;
      RECT 6.4170 34.8270 6.4350 35.1770 ;
      RECT 6.3090 34.8270 6.3270 35.1770 ;
      RECT 6.2010 34.8270 6.2190 35.1770 ;
      RECT 6.0930 34.8270 6.1110 35.1770 ;
      RECT 5.9850 34.8270 6.0030 35.1770 ;
      RECT 5.8770 34.8270 5.8950 35.1770 ;
      RECT 5.7690 34.8270 5.7870 35.1770 ;
      RECT 5.6610 34.8270 5.6790 35.1770 ;
      RECT 5.5530 34.8270 5.5710 35.1770 ;
      RECT 5.4450 34.8270 5.4630 35.1770 ;
      RECT 5.3370 34.8270 5.3550 35.1770 ;
      RECT 5.2290 34.8270 5.2470 35.1770 ;
      RECT 5.1210 34.8270 5.1390 35.1770 ;
      RECT 5.0130 34.8270 5.0310 35.1770 ;
      RECT 4.9050 34.8270 4.9230 35.1770 ;
      RECT 4.7970 34.8270 4.8150 35.1770 ;
      RECT 4.6890 34.8270 4.7070 35.1770 ;
      RECT 4.5810 34.8270 4.5990 35.1770 ;
      RECT 4.4730 34.8270 4.4910 35.1770 ;
      RECT 4.3650 34.8270 4.3830 35.1770 ;
      RECT 4.2570 34.8270 4.2750 35.1770 ;
      RECT 4.1490 34.8270 4.1670 35.1770 ;
      RECT 4.0410 34.8270 4.0590 35.1770 ;
      RECT 3.9330 34.8270 3.9510 35.1770 ;
      RECT 3.8250 34.8270 3.8430 35.1770 ;
      RECT 3.7170 34.8270 3.7350 35.1770 ;
      RECT 3.6090 34.8270 3.6270 35.1770 ;
      RECT 3.5010 34.8270 3.5190 35.1770 ;
      RECT 3.3930 34.8270 3.4110 35.1770 ;
      RECT 3.2850 34.8270 3.3030 35.1770 ;
      RECT 3.1770 34.8270 3.1950 35.1770 ;
      RECT 3.0690 34.8270 3.0870 35.1770 ;
      RECT 2.9610 34.8270 2.9790 35.1770 ;
      RECT 2.8530 34.8270 2.8710 35.1770 ;
      RECT 2.7450 34.8270 2.7630 35.1770 ;
      RECT 2.6370 34.8270 2.6550 35.1770 ;
      RECT 2.5290 34.8270 2.5470 35.1770 ;
      RECT 2.4210 34.8270 2.4390 35.1770 ;
      RECT 2.3130 34.8270 2.3310 35.1770 ;
      RECT 2.2050 34.8270 2.2230 35.1770 ;
      RECT 2.0970 34.8270 2.1150 35.1770 ;
      RECT 1.9890 34.8270 2.0070 35.1770 ;
      RECT 1.8810 34.8270 1.8990 35.1770 ;
      RECT 1.7730 34.8270 1.7910 35.1770 ;
      RECT 1.6650 34.8270 1.6830 35.1770 ;
      RECT 1.5570 34.8270 1.5750 35.1770 ;
      RECT 1.4490 34.8270 1.4670 35.1770 ;
      RECT 1.3410 34.8270 1.3590 35.1770 ;
      RECT 1.2330 34.8270 1.2510 35.1770 ;
      RECT 1.1250 34.8270 1.1430 35.1770 ;
      RECT 1.0170 34.8270 1.0350 35.1770 ;
      RECT 0.9090 34.8270 0.9270 35.1770 ;
      RECT 0.8010 34.8270 0.8190 35.1770 ;
      RECT 0.6930 34.8270 0.7110 35.1770 ;
      RECT 0.5850 34.8270 0.6030 35.1770 ;
      RECT 0.4770 34.8270 0.4950 35.1770 ;
      RECT 0.3690 34.8270 0.3870 35.1770 ;
      RECT 0.2610 34.8270 0.2790 35.1770 ;
      RECT 0.1530 34.8270 0.1710 43.0340 ;
      RECT 0.1170 34.8270 0.1350 43.0340 ;
        RECT 15.6110 43.0320 15.6290 43.9675 ;
        RECT 15.5750 43.0320 15.5930 43.9675 ;
        RECT 15.5390 43.6090 15.5570 43.9315 ;
        RECT 15.4220 43.8060 15.4400 43.9155 ;
        RECT 15.4130 43.0645 15.4310 43.3040 ;
        RECT 15.3770 43.6455 15.3950 43.7990 ;
        RECT 15.2960 43.6710 15.3140 43.9290 ;
        RECT 14.7560 43.0320 14.7740 43.9675 ;
        RECT 14.7200 43.0320 14.7380 43.9675 ;
        RECT 14.6840 43.2130 14.7020 43.7810 ;
        RECT 15.6110 44.1120 15.6290 45.0475 ;
        RECT 15.5750 44.1120 15.5930 45.0475 ;
        RECT 15.5390 44.6890 15.5570 45.0115 ;
        RECT 15.4220 44.8860 15.4400 44.9955 ;
        RECT 15.4130 44.1445 15.4310 44.3840 ;
        RECT 15.3770 44.7255 15.3950 44.8790 ;
        RECT 15.2960 44.7510 15.3140 45.0090 ;
        RECT 14.7560 44.1120 14.7740 45.0475 ;
        RECT 14.7200 44.1120 14.7380 45.0475 ;
        RECT 14.6840 44.2930 14.7020 44.8610 ;
        RECT 15.6110 45.1920 15.6290 46.1275 ;
        RECT 15.5750 45.1920 15.5930 46.1275 ;
        RECT 15.5390 45.7690 15.5570 46.0915 ;
        RECT 15.4220 45.9660 15.4400 46.0755 ;
        RECT 15.4130 45.2245 15.4310 45.4640 ;
        RECT 15.3770 45.8055 15.3950 45.9590 ;
        RECT 15.2960 45.8310 15.3140 46.0890 ;
        RECT 14.7560 45.1920 14.7740 46.1275 ;
        RECT 14.7200 45.1920 14.7380 46.1275 ;
        RECT 14.6840 45.3730 14.7020 45.9410 ;
        RECT 15.6110 46.2720 15.6290 47.2075 ;
        RECT 15.5750 46.2720 15.5930 47.2075 ;
        RECT 15.5390 46.8490 15.5570 47.1715 ;
        RECT 15.4220 47.0460 15.4400 47.1555 ;
        RECT 15.4130 46.3045 15.4310 46.5440 ;
        RECT 15.3770 46.8855 15.3950 47.0390 ;
        RECT 15.2960 46.9110 15.3140 47.1690 ;
        RECT 14.7560 46.2720 14.7740 47.2075 ;
        RECT 14.7200 46.2720 14.7380 47.2075 ;
        RECT 14.6840 46.4530 14.7020 47.0210 ;
        RECT 15.6110 47.3520 15.6290 48.2875 ;
        RECT 15.5750 47.3520 15.5930 48.2875 ;
        RECT 15.5390 47.9290 15.5570 48.2515 ;
        RECT 15.4220 48.1260 15.4400 48.2355 ;
        RECT 15.4130 47.3845 15.4310 47.6240 ;
        RECT 15.3770 47.9655 15.3950 48.1190 ;
        RECT 15.2960 47.9910 15.3140 48.2490 ;
        RECT 14.7560 47.3520 14.7740 48.2875 ;
        RECT 14.7200 47.3520 14.7380 48.2875 ;
        RECT 14.6840 47.5330 14.7020 48.1010 ;
        RECT 15.6110 48.4320 15.6290 49.3675 ;
        RECT 15.5750 48.4320 15.5930 49.3675 ;
        RECT 15.5390 49.0090 15.5570 49.3315 ;
        RECT 15.4220 49.2060 15.4400 49.3155 ;
        RECT 15.4130 48.4645 15.4310 48.7040 ;
        RECT 15.3770 49.0455 15.3950 49.1990 ;
        RECT 15.2960 49.0710 15.3140 49.3290 ;
        RECT 14.7560 48.4320 14.7740 49.3675 ;
        RECT 14.7200 48.4320 14.7380 49.3675 ;
        RECT 14.6840 48.6130 14.7020 49.1810 ;
        RECT 15.6110 49.5120 15.6290 50.4475 ;
        RECT 15.5750 49.5120 15.5930 50.4475 ;
        RECT 15.5390 50.0890 15.5570 50.4115 ;
        RECT 15.4220 50.2860 15.4400 50.3955 ;
        RECT 15.4130 49.5445 15.4310 49.7840 ;
        RECT 15.3770 50.1255 15.3950 50.2790 ;
        RECT 15.2960 50.1510 15.3140 50.4090 ;
        RECT 14.7560 49.5120 14.7740 50.4475 ;
        RECT 14.7200 49.5120 14.7380 50.4475 ;
        RECT 14.6840 49.6930 14.7020 50.2610 ;
        RECT 15.6110 50.5920 15.6290 51.5275 ;
        RECT 15.5750 50.5920 15.5930 51.5275 ;
        RECT 15.5390 51.1690 15.5570 51.4915 ;
        RECT 15.4220 51.3660 15.4400 51.4755 ;
        RECT 15.4130 50.6245 15.4310 50.8640 ;
        RECT 15.3770 51.2055 15.3950 51.3590 ;
        RECT 15.2960 51.2310 15.3140 51.4890 ;
        RECT 14.7560 50.5920 14.7740 51.5275 ;
        RECT 14.7200 50.5920 14.7380 51.5275 ;
        RECT 14.6840 50.7730 14.7020 51.3410 ;
        RECT 15.6110 51.6720 15.6290 52.6075 ;
        RECT 15.5750 51.6720 15.5930 52.6075 ;
        RECT 15.5390 52.2490 15.5570 52.5715 ;
        RECT 15.4220 52.4460 15.4400 52.5555 ;
        RECT 15.4130 51.7045 15.4310 51.9440 ;
        RECT 15.3770 52.2855 15.3950 52.4390 ;
        RECT 15.2960 52.3110 15.3140 52.5690 ;
        RECT 14.7560 51.6720 14.7740 52.6075 ;
        RECT 14.7200 51.6720 14.7380 52.6075 ;
        RECT 14.6840 51.8530 14.7020 52.4210 ;
        RECT 15.6110 52.7520 15.6290 53.6875 ;
        RECT 15.5750 52.7520 15.5930 53.6875 ;
        RECT 15.5390 53.3290 15.5570 53.6515 ;
        RECT 15.4220 53.5260 15.4400 53.6355 ;
        RECT 15.4130 52.7845 15.4310 53.0240 ;
        RECT 15.3770 53.3655 15.3950 53.5190 ;
        RECT 15.2960 53.3910 15.3140 53.6490 ;
        RECT 14.7560 52.7520 14.7740 53.6875 ;
        RECT 14.7200 52.7520 14.7380 53.6875 ;
        RECT 14.6840 52.9330 14.7020 53.5010 ;
        RECT 15.6110 53.8320 15.6290 54.7675 ;
        RECT 15.5750 53.8320 15.5930 54.7675 ;
        RECT 15.5390 54.4090 15.5570 54.7315 ;
        RECT 15.4220 54.6060 15.4400 54.7155 ;
        RECT 15.4130 53.8645 15.4310 54.1040 ;
        RECT 15.3770 54.4455 15.3950 54.5990 ;
        RECT 15.2960 54.4710 15.3140 54.7290 ;
        RECT 14.7560 53.8320 14.7740 54.7675 ;
        RECT 14.7200 53.8320 14.7380 54.7675 ;
        RECT 14.6840 54.0130 14.7020 54.5810 ;
        RECT 15.6110 54.9120 15.6290 55.8475 ;
        RECT 15.5750 54.9120 15.5930 55.8475 ;
        RECT 15.5390 55.4890 15.5570 55.8115 ;
        RECT 15.4220 55.6860 15.4400 55.7955 ;
        RECT 15.4130 54.9445 15.4310 55.1840 ;
        RECT 15.3770 55.5255 15.3950 55.6790 ;
        RECT 15.2960 55.5510 15.3140 55.8090 ;
        RECT 14.7560 54.9120 14.7740 55.8475 ;
        RECT 14.7200 54.9120 14.7380 55.8475 ;
        RECT 14.6840 55.0930 14.7020 55.6610 ;
        RECT 15.6110 55.9920 15.6290 56.9275 ;
        RECT 15.5750 55.9920 15.5930 56.9275 ;
        RECT 15.5390 56.5690 15.5570 56.8915 ;
        RECT 15.4220 56.7660 15.4400 56.8755 ;
        RECT 15.4130 56.0245 15.4310 56.2640 ;
        RECT 15.3770 56.6055 15.3950 56.7590 ;
        RECT 15.2960 56.6310 15.3140 56.8890 ;
        RECT 14.7560 55.9920 14.7740 56.9275 ;
        RECT 14.7200 55.9920 14.7380 56.9275 ;
        RECT 14.6840 56.1730 14.7020 56.7410 ;
        RECT 15.6110 57.0720 15.6290 58.0075 ;
        RECT 15.5750 57.0720 15.5930 58.0075 ;
        RECT 15.5390 57.6490 15.5570 57.9715 ;
        RECT 15.4220 57.8460 15.4400 57.9555 ;
        RECT 15.4130 57.1045 15.4310 57.3440 ;
        RECT 15.3770 57.6855 15.3950 57.8390 ;
        RECT 15.2960 57.7110 15.3140 57.9690 ;
        RECT 14.7560 57.0720 14.7740 58.0075 ;
        RECT 14.7200 57.0720 14.7380 58.0075 ;
        RECT 14.6840 57.2530 14.7020 57.8210 ;
        RECT 15.6110 58.1520 15.6290 59.0875 ;
        RECT 15.5750 58.1520 15.5930 59.0875 ;
        RECT 15.5390 58.7290 15.5570 59.0515 ;
        RECT 15.4220 58.9260 15.4400 59.0355 ;
        RECT 15.4130 58.1845 15.4310 58.4240 ;
        RECT 15.3770 58.7655 15.3950 58.9190 ;
        RECT 15.2960 58.7910 15.3140 59.0490 ;
        RECT 14.7560 58.1520 14.7740 59.0875 ;
        RECT 14.7200 58.1520 14.7380 59.0875 ;
        RECT 14.6840 58.3330 14.7020 58.9010 ;
        RECT 15.6110 59.2320 15.6290 60.1675 ;
        RECT 15.5750 59.2320 15.5930 60.1675 ;
        RECT 15.5390 59.8090 15.5570 60.1315 ;
        RECT 15.4220 60.0060 15.4400 60.1155 ;
        RECT 15.4130 59.2645 15.4310 59.5040 ;
        RECT 15.3770 59.8455 15.3950 59.9990 ;
        RECT 15.2960 59.8710 15.3140 60.1290 ;
        RECT 14.7560 59.2320 14.7740 60.1675 ;
        RECT 14.7200 59.2320 14.7380 60.1675 ;
        RECT 14.6840 59.4130 14.7020 59.9810 ;
        RECT 15.6110 60.3120 15.6290 61.2475 ;
        RECT 15.5750 60.3120 15.5930 61.2475 ;
        RECT 15.5390 60.8890 15.5570 61.2115 ;
        RECT 15.4220 61.0860 15.4400 61.1955 ;
        RECT 15.4130 60.3445 15.4310 60.5840 ;
        RECT 15.3770 60.9255 15.3950 61.0790 ;
        RECT 15.2960 60.9510 15.3140 61.2090 ;
        RECT 14.7560 60.3120 14.7740 61.2475 ;
        RECT 14.7200 60.3120 14.7380 61.2475 ;
        RECT 14.6840 60.4930 14.7020 61.0610 ;
        RECT 15.6110 61.3920 15.6290 62.3275 ;
        RECT 15.5750 61.3920 15.5930 62.3275 ;
        RECT 15.5390 61.9690 15.5570 62.2915 ;
        RECT 15.4220 62.1660 15.4400 62.2755 ;
        RECT 15.4130 61.4245 15.4310 61.6640 ;
        RECT 15.3770 62.0055 15.3950 62.1590 ;
        RECT 15.2960 62.0310 15.3140 62.2890 ;
        RECT 14.7560 61.3920 14.7740 62.3275 ;
        RECT 14.7200 61.3920 14.7380 62.3275 ;
        RECT 14.6840 61.5730 14.7020 62.1410 ;
        RECT 15.6110 62.4720 15.6290 63.4075 ;
        RECT 15.5750 62.4720 15.5930 63.4075 ;
        RECT 15.5390 63.0490 15.5570 63.3715 ;
        RECT 15.4220 63.2460 15.4400 63.3555 ;
        RECT 15.4130 62.5045 15.4310 62.7440 ;
        RECT 15.3770 63.0855 15.3950 63.2390 ;
        RECT 15.2960 63.1110 15.3140 63.3690 ;
        RECT 14.7560 62.4720 14.7740 63.4075 ;
        RECT 14.7200 62.4720 14.7380 63.4075 ;
        RECT 14.6840 62.6530 14.7020 63.2210 ;
        RECT 15.6110 63.5520 15.6290 64.4875 ;
        RECT 15.5750 63.5520 15.5930 64.4875 ;
        RECT 15.5390 64.1290 15.5570 64.4515 ;
        RECT 15.4220 64.3260 15.4400 64.4355 ;
        RECT 15.4130 63.5845 15.4310 63.8240 ;
        RECT 15.3770 64.1655 15.3950 64.3190 ;
        RECT 15.2960 64.1910 15.3140 64.4490 ;
        RECT 14.7560 63.5520 14.7740 64.4875 ;
        RECT 14.7200 63.5520 14.7380 64.4875 ;
        RECT 14.6840 63.7330 14.7020 64.3010 ;
        RECT 15.6110 64.6320 15.6290 65.5675 ;
        RECT 15.5750 64.6320 15.5930 65.5675 ;
        RECT 15.5390 65.2090 15.5570 65.5315 ;
        RECT 15.4220 65.4060 15.4400 65.5155 ;
        RECT 15.4130 64.6645 15.4310 64.9040 ;
        RECT 15.3770 65.2455 15.3950 65.3990 ;
        RECT 15.2960 65.2710 15.3140 65.5290 ;
        RECT 14.7560 64.6320 14.7740 65.5675 ;
        RECT 14.7200 64.6320 14.7380 65.5675 ;
        RECT 14.6840 64.8130 14.7020 65.3810 ;
        RECT 15.6110 65.7120 15.6290 66.6475 ;
        RECT 15.5750 65.7120 15.5930 66.6475 ;
        RECT 15.5390 66.2890 15.5570 66.6115 ;
        RECT 15.4220 66.4860 15.4400 66.5955 ;
        RECT 15.4130 65.7445 15.4310 65.9840 ;
        RECT 15.3770 66.3255 15.3950 66.4790 ;
        RECT 15.2960 66.3510 15.3140 66.6090 ;
        RECT 14.7560 65.7120 14.7740 66.6475 ;
        RECT 14.7200 65.7120 14.7380 66.6475 ;
        RECT 14.6840 65.8930 14.7020 66.4610 ;
        RECT 15.6110 66.7920 15.6290 67.7275 ;
        RECT 15.5750 66.7920 15.5930 67.7275 ;
        RECT 15.5390 67.3690 15.5570 67.6915 ;
        RECT 15.4220 67.5660 15.4400 67.6755 ;
        RECT 15.4130 66.8245 15.4310 67.0640 ;
        RECT 15.3770 67.4055 15.3950 67.5590 ;
        RECT 15.2960 67.4310 15.3140 67.6890 ;
        RECT 14.7560 66.7920 14.7740 67.7275 ;
        RECT 14.7200 66.7920 14.7380 67.7275 ;
        RECT 14.6840 66.9730 14.7020 67.5410 ;
        RECT 15.6110 67.8720 15.6290 68.8075 ;
        RECT 15.5750 67.8720 15.5930 68.8075 ;
        RECT 15.5390 68.4490 15.5570 68.7715 ;
        RECT 15.4220 68.6460 15.4400 68.7555 ;
        RECT 15.4130 67.9045 15.4310 68.1440 ;
        RECT 15.3770 68.4855 15.3950 68.6390 ;
        RECT 15.2960 68.5110 15.3140 68.7690 ;
        RECT 14.7560 67.8720 14.7740 68.8075 ;
        RECT 14.7200 67.8720 14.7380 68.8075 ;
        RECT 14.6840 68.0530 14.7020 68.6210 ;
        RECT 15.6110 68.9520 15.6290 69.8875 ;
        RECT 15.5750 68.9520 15.5930 69.8875 ;
        RECT 15.5390 69.5290 15.5570 69.8515 ;
        RECT 15.4220 69.7260 15.4400 69.8355 ;
        RECT 15.4130 68.9845 15.4310 69.2240 ;
        RECT 15.3770 69.5655 15.3950 69.7190 ;
        RECT 15.2960 69.5910 15.3140 69.8490 ;
        RECT 14.7560 68.9520 14.7740 69.8875 ;
        RECT 14.7200 68.9520 14.7380 69.8875 ;
        RECT 14.6840 69.1330 14.7020 69.7010 ;
        RECT 15.6110 70.0320 15.6290 70.9675 ;
        RECT 15.5750 70.0320 15.5930 70.9675 ;
        RECT 15.5390 70.6090 15.5570 70.9315 ;
        RECT 15.4220 70.8060 15.4400 70.9155 ;
        RECT 15.4130 70.0645 15.4310 70.3040 ;
        RECT 15.3770 70.6455 15.3950 70.7990 ;
        RECT 15.2960 70.6710 15.3140 70.9290 ;
        RECT 14.7560 70.0320 14.7740 70.9675 ;
        RECT 14.7200 70.0320 14.7380 70.9675 ;
        RECT 14.6840 70.2130 14.7020 70.7810 ;
        RECT 15.6110 71.1120 15.6290 72.0475 ;
        RECT 15.5750 71.1120 15.5930 72.0475 ;
        RECT 15.5390 71.6890 15.5570 72.0115 ;
        RECT 15.4220 71.8860 15.4400 71.9955 ;
        RECT 15.4130 71.1445 15.4310 71.3840 ;
        RECT 15.3770 71.7255 15.3950 71.8790 ;
        RECT 15.2960 71.7510 15.3140 72.0090 ;
        RECT 14.7560 71.1120 14.7740 72.0475 ;
        RECT 14.7200 71.1120 14.7380 72.0475 ;
        RECT 14.6840 71.2930 14.7020 71.8610 ;
        RECT 15.6110 72.1920 15.6290 73.1275 ;
        RECT 15.5750 72.1920 15.5930 73.1275 ;
        RECT 15.5390 72.7690 15.5570 73.0915 ;
        RECT 15.4220 72.9660 15.4400 73.0755 ;
        RECT 15.4130 72.2245 15.4310 72.4640 ;
        RECT 15.3770 72.8055 15.3950 72.9590 ;
        RECT 15.2960 72.8310 15.3140 73.0890 ;
        RECT 14.7560 72.1920 14.7740 73.1275 ;
        RECT 14.7200 72.1920 14.7380 73.1275 ;
        RECT 14.6840 72.3730 14.7020 72.9410 ;
        RECT 15.6110 73.2720 15.6290 74.2075 ;
        RECT 15.5750 73.2720 15.5930 74.2075 ;
        RECT 15.5390 73.8490 15.5570 74.1715 ;
        RECT 15.4220 74.0460 15.4400 74.1555 ;
        RECT 15.4130 73.3045 15.4310 73.5440 ;
        RECT 15.3770 73.8855 15.3950 74.0390 ;
        RECT 15.2960 73.9110 15.3140 74.1690 ;
        RECT 14.7560 73.2720 14.7740 74.2075 ;
        RECT 14.7200 73.2720 14.7380 74.2075 ;
        RECT 14.6840 73.4530 14.7020 74.0210 ;
        RECT 15.6110 74.3520 15.6290 75.2875 ;
        RECT 15.5750 74.3520 15.5930 75.2875 ;
        RECT 15.5390 74.9290 15.5570 75.2515 ;
        RECT 15.4220 75.1260 15.4400 75.2355 ;
        RECT 15.4130 74.3845 15.4310 74.6240 ;
        RECT 15.3770 74.9655 15.3950 75.1190 ;
        RECT 15.2960 74.9910 15.3140 75.2490 ;
        RECT 14.7560 74.3520 14.7740 75.2875 ;
        RECT 14.7200 74.3520 14.7380 75.2875 ;
        RECT 14.6840 74.5330 14.7020 75.1010 ;
        RECT 15.6110 75.4320 15.6290 76.3675 ;
        RECT 15.5750 75.4320 15.5930 76.3675 ;
        RECT 15.5390 76.0090 15.5570 76.3315 ;
        RECT 15.4220 76.2060 15.4400 76.3155 ;
        RECT 15.4130 75.4645 15.4310 75.7040 ;
        RECT 15.3770 76.0455 15.3950 76.1990 ;
        RECT 15.2960 76.0710 15.3140 76.3290 ;
        RECT 14.7560 75.4320 14.7740 76.3675 ;
        RECT 14.7200 75.4320 14.7380 76.3675 ;
        RECT 14.6840 75.6130 14.7020 76.1810 ;
        RECT 15.6110 76.5120 15.6290 77.4475 ;
        RECT 15.5750 76.5120 15.5930 77.4475 ;
        RECT 15.5390 77.0890 15.5570 77.4115 ;
        RECT 15.4220 77.2860 15.4400 77.3955 ;
        RECT 15.4130 76.5445 15.4310 76.7840 ;
        RECT 15.3770 77.1255 15.3950 77.2790 ;
        RECT 15.2960 77.1510 15.3140 77.4090 ;
        RECT 14.7560 76.5120 14.7740 77.4475 ;
        RECT 14.7200 76.5120 14.7380 77.4475 ;
        RECT 14.6840 76.6930 14.7020 77.2610 ;
  LAYER M3 SPACING 0.018  ;
      RECT 15.5530 0.2565 15.6810 1.3500 ;
      RECT 15.5390 0.9220 15.6810 1.2445 ;
      RECT 15.3190 0.6490 15.4530 1.3500 ;
      RECT 15.2960 0.9840 15.4530 1.2420 ;
      RECT 15.3190 0.2565 15.4170 1.3500 ;
      RECT 15.3190 0.3775 15.4310 0.6170 ;
      RECT 15.3190 0.2565 15.4530 0.3455 ;
      RECT 15.0940 0.7070 15.2280 1.3500 ;
      RECT 15.0940 0.2565 15.1920 1.3500 ;
      RECT 14.6770 0.2565 14.7600 1.3500 ;
      RECT 14.6770 0.3450 14.7740 1.2805 ;
      RECT 30.2680 0.2565 30.3530 1.3500 ;
      RECT 30.1240 0.2565 30.1500 1.3500 ;
      RECT 30.0160 0.2565 30.0420 1.3500 ;
      RECT 29.9080 0.2565 29.9340 1.3500 ;
      RECT 29.8000 0.2565 29.8260 1.3500 ;
      RECT 29.6920 0.2565 29.7180 1.3500 ;
      RECT 29.5840 0.2565 29.6100 1.3500 ;
      RECT 29.4760 0.2565 29.5020 1.3500 ;
      RECT 29.3680 0.2565 29.3940 1.3500 ;
      RECT 29.2600 0.2565 29.2860 1.3500 ;
      RECT 29.1520 0.2565 29.1780 1.3500 ;
      RECT 29.0440 0.2565 29.0700 1.3500 ;
      RECT 28.9360 0.2565 28.9620 1.3500 ;
      RECT 28.8280 0.2565 28.8540 1.3500 ;
      RECT 28.7200 0.2565 28.7460 1.3500 ;
      RECT 28.6120 0.2565 28.6380 1.3500 ;
      RECT 28.5040 0.2565 28.5300 1.3500 ;
      RECT 28.3960 0.2565 28.4220 1.3500 ;
      RECT 28.2880 0.2565 28.3140 1.3500 ;
      RECT 28.1800 0.2565 28.2060 1.3500 ;
      RECT 28.0720 0.2565 28.0980 1.3500 ;
      RECT 27.9640 0.2565 27.9900 1.3500 ;
      RECT 27.8560 0.2565 27.8820 1.3500 ;
      RECT 27.7480 0.2565 27.7740 1.3500 ;
      RECT 27.6400 0.2565 27.6660 1.3500 ;
      RECT 27.5320 0.2565 27.5580 1.3500 ;
      RECT 27.4240 0.2565 27.4500 1.3500 ;
      RECT 27.3160 0.2565 27.3420 1.3500 ;
      RECT 27.2080 0.2565 27.2340 1.3500 ;
      RECT 27.1000 0.2565 27.1260 1.3500 ;
      RECT 26.9920 0.2565 27.0180 1.3500 ;
      RECT 26.8840 0.2565 26.9100 1.3500 ;
      RECT 26.7760 0.2565 26.8020 1.3500 ;
      RECT 26.6680 0.2565 26.6940 1.3500 ;
      RECT 26.5600 0.2565 26.5860 1.3500 ;
      RECT 26.4520 0.2565 26.4780 1.3500 ;
      RECT 26.3440 0.2565 26.3700 1.3500 ;
      RECT 26.2360 0.2565 26.2620 1.3500 ;
      RECT 26.1280 0.2565 26.1540 1.3500 ;
      RECT 26.0200 0.2565 26.0460 1.3500 ;
      RECT 25.9120 0.2565 25.9380 1.3500 ;
      RECT 25.8040 0.2565 25.8300 1.3500 ;
      RECT 25.6960 0.2565 25.7220 1.3500 ;
      RECT 25.5880 0.2565 25.6140 1.3500 ;
      RECT 25.4800 0.2565 25.5060 1.3500 ;
      RECT 25.3720 0.2565 25.3980 1.3500 ;
      RECT 25.2640 0.2565 25.2900 1.3500 ;
      RECT 25.1560 0.2565 25.1820 1.3500 ;
      RECT 25.0480 0.2565 25.0740 1.3500 ;
      RECT 24.9400 0.2565 24.9660 1.3500 ;
      RECT 24.8320 0.2565 24.8580 1.3500 ;
      RECT 24.7240 0.2565 24.7500 1.3500 ;
      RECT 24.6160 0.2565 24.6420 1.3500 ;
      RECT 24.5080 0.2565 24.5340 1.3500 ;
      RECT 24.4000 0.2565 24.4260 1.3500 ;
      RECT 24.2920 0.2565 24.3180 1.3500 ;
      RECT 24.1840 0.2565 24.2100 1.3500 ;
      RECT 24.0760 0.2565 24.1020 1.3500 ;
      RECT 23.9680 0.2565 23.9940 1.3500 ;
      RECT 23.8600 0.2565 23.8860 1.3500 ;
      RECT 23.7520 0.2565 23.7780 1.3500 ;
      RECT 23.6440 0.2565 23.6700 1.3500 ;
      RECT 23.5360 0.2565 23.5620 1.3500 ;
      RECT 23.4280 0.2565 23.4540 1.3500 ;
      RECT 23.3200 0.2565 23.3460 1.3500 ;
      RECT 23.2120 0.2565 23.2380 1.3500 ;
      RECT 23.1040 0.2565 23.1300 1.3500 ;
      RECT 22.9960 0.2565 23.0220 1.3500 ;
      RECT 22.8880 0.2565 22.9140 1.3500 ;
      RECT 22.7800 0.2565 22.8060 1.3500 ;
      RECT 22.6720 0.2565 22.6980 1.3500 ;
      RECT 22.5640 0.2565 22.5900 1.3500 ;
      RECT 22.4560 0.2565 22.4820 1.3500 ;
      RECT 22.3480 0.2565 22.3740 1.3500 ;
      RECT 22.2400 0.2565 22.2660 1.3500 ;
      RECT 22.1320 0.2565 22.1580 1.3500 ;
      RECT 22.0240 0.2565 22.0500 1.3500 ;
      RECT 21.9160 0.2565 21.9420 1.3500 ;
      RECT 21.8080 0.2565 21.8340 1.3500 ;
      RECT 21.7000 0.2565 21.7260 1.3500 ;
      RECT 21.5920 0.2565 21.6180 1.3500 ;
      RECT 21.4840 0.2565 21.5100 1.3500 ;
      RECT 21.3760 0.2565 21.4020 1.3500 ;
      RECT 21.2680 0.2565 21.2940 1.3500 ;
      RECT 21.1600 0.2565 21.1860 1.3500 ;
      RECT 21.0520 0.2565 21.0780 1.3500 ;
      RECT 20.9440 0.2565 20.9700 1.3500 ;
      RECT 20.8360 0.2565 20.8620 1.3500 ;
      RECT 20.7280 0.2565 20.7540 1.3500 ;
      RECT 20.6200 0.2565 20.6460 1.3500 ;
      RECT 20.5120 0.2565 20.5380 1.3500 ;
      RECT 20.4040 0.2565 20.4300 1.3500 ;
      RECT 20.2960 0.2565 20.3220 1.3500 ;
      RECT 20.1880 0.2565 20.2140 1.3500 ;
      RECT 20.0800 0.2565 20.1060 1.3500 ;
      RECT 19.9720 0.2565 19.9980 1.3500 ;
      RECT 19.8640 0.2565 19.8900 1.3500 ;
      RECT 19.7560 0.2565 19.7820 1.3500 ;
      RECT 19.6480 0.2565 19.6740 1.3500 ;
      RECT 19.5400 0.2565 19.5660 1.3500 ;
      RECT 19.4320 0.2565 19.4580 1.3500 ;
      RECT 19.3240 0.2565 19.3500 1.3500 ;
      RECT 19.2160 0.2565 19.2420 1.3500 ;
      RECT 19.1080 0.2565 19.1340 1.3500 ;
      RECT 19.0000 0.2565 19.0260 1.3500 ;
      RECT 18.8920 0.2565 18.9180 1.3500 ;
      RECT 18.7840 0.2565 18.8100 1.3500 ;
      RECT 18.6760 0.2565 18.7020 1.3500 ;
      RECT 18.5680 0.2565 18.5940 1.3500 ;
      RECT 18.4600 0.2565 18.4860 1.3500 ;
      RECT 18.3520 0.2565 18.3780 1.3500 ;
      RECT 18.2440 0.2565 18.2700 1.3500 ;
      RECT 18.1360 0.2565 18.1620 1.3500 ;
      RECT 18.0280 0.2565 18.0540 1.3500 ;
      RECT 17.9200 0.2565 17.9460 1.3500 ;
      RECT 17.8120 0.2565 17.8380 1.3500 ;
      RECT 17.7040 0.2565 17.7300 1.3500 ;
      RECT 17.5960 0.2565 17.6220 1.3500 ;
      RECT 17.4880 0.2565 17.5140 1.3500 ;
      RECT 17.3800 0.2565 17.4060 1.3500 ;
      RECT 17.2720 0.2565 17.2980 1.3500 ;
      RECT 17.1640 0.2565 17.1900 1.3500 ;
      RECT 17.0560 0.2565 17.0820 1.3500 ;
      RECT 16.9480 0.2565 16.9740 1.3500 ;
      RECT 16.8400 0.2565 16.8660 1.3500 ;
      RECT 16.7320 0.2565 16.7580 1.3500 ;
      RECT 16.6240 0.2565 16.6500 1.3500 ;
      RECT 16.5160 0.2565 16.5420 1.3500 ;
      RECT 16.4080 0.2565 16.4340 1.3500 ;
      RECT 16.3000 0.2565 16.3260 1.3500 ;
      RECT 16.0870 0.2565 16.1640 1.3500 ;
      RECT 14.1940 0.2565 14.2710 1.3500 ;
      RECT 14.0320 0.2565 14.0580 1.3500 ;
      RECT 13.9240 0.2565 13.9500 1.3500 ;
      RECT 13.8160 0.2565 13.8420 1.3500 ;
      RECT 13.7080 0.2565 13.7340 1.3500 ;
      RECT 13.6000 0.2565 13.6260 1.3500 ;
      RECT 13.4920 0.2565 13.5180 1.3500 ;
      RECT 13.3840 0.2565 13.4100 1.3500 ;
      RECT 13.2760 0.2565 13.3020 1.3500 ;
      RECT 13.1680 0.2565 13.1940 1.3500 ;
      RECT 13.0600 0.2565 13.0860 1.3500 ;
      RECT 12.9520 0.2565 12.9780 1.3500 ;
      RECT 12.8440 0.2565 12.8700 1.3500 ;
      RECT 12.7360 0.2565 12.7620 1.3500 ;
      RECT 12.6280 0.2565 12.6540 1.3500 ;
      RECT 12.5200 0.2565 12.5460 1.3500 ;
      RECT 12.4120 0.2565 12.4380 1.3500 ;
      RECT 12.3040 0.2565 12.3300 1.3500 ;
      RECT 12.1960 0.2565 12.2220 1.3500 ;
      RECT 12.0880 0.2565 12.1140 1.3500 ;
      RECT 11.9800 0.2565 12.0060 1.3500 ;
      RECT 11.8720 0.2565 11.8980 1.3500 ;
      RECT 11.7640 0.2565 11.7900 1.3500 ;
      RECT 11.6560 0.2565 11.6820 1.3500 ;
      RECT 11.5480 0.2565 11.5740 1.3500 ;
      RECT 11.4400 0.2565 11.4660 1.3500 ;
      RECT 11.3320 0.2565 11.3580 1.3500 ;
      RECT 11.2240 0.2565 11.2500 1.3500 ;
      RECT 11.1160 0.2565 11.1420 1.3500 ;
      RECT 11.0080 0.2565 11.0340 1.3500 ;
      RECT 10.9000 0.2565 10.9260 1.3500 ;
      RECT 10.7920 0.2565 10.8180 1.3500 ;
      RECT 10.6840 0.2565 10.7100 1.3500 ;
      RECT 10.5760 0.2565 10.6020 1.3500 ;
      RECT 10.4680 0.2565 10.4940 1.3500 ;
      RECT 10.3600 0.2565 10.3860 1.3500 ;
      RECT 10.2520 0.2565 10.2780 1.3500 ;
      RECT 10.1440 0.2565 10.1700 1.3500 ;
      RECT 10.0360 0.2565 10.0620 1.3500 ;
      RECT 9.9280 0.2565 9.9540 1.3500 ;
      RECT 9.8200 0.2565 9.8460 1.3500 ;
      RECT 9.7120 0.2565 9.7380 1.3500 ;
      RECT 9.6040 0.2565 9.6300 1.3500 ;
      RECT 9.4960 0.2565 9.5220 1.3500 ;
      RECT 9.3880 0.2565 9.4140 1.3500 ;
      RECT 9.2800 0.2565 9.3060 1.3500 ;
      RECT 9.1720 0.2565 9.1980 1.3500 ;
      RECT 9.0640 0.2565 9.0900 1.3500 ;
      RECT 8.9560 0.2565 8.9820 1.3500 ;
      RECT 8.8480 0.2565 8.8740 1.3500 ;
      RECT 8.7400 0.2565 8.7660 1.3500 ;
      RECT 8.6320 0.2565 8.6580 1.3500 ;
      RECT 8.5240 0.2565 8.5500 1.3500 ;
      RECT 8.4160 0.2565 8.4420 1.3500 ;
      RECT 8.3080 0.2565 8.3340 1.3500 ;
      RECT 8.2000 0.2565 8.2260 1.3500 ;
      RECT 8.0920 0.2565 8.1180 1.3500 ;
      RECT 7.9840 0.2565 8.0100 1.3500 ;
      RECT 7.8760 0.2565 7.9020 1.3500 ;
      RECT 7.7680 0.2565 7.7940 1.3500 ;
      RECT 7.6600 0.2565 7.6860 1.3500 ;
      RECT 7.5520 0.2565 7.5780 1.3500 ;
      RECT 7.4440 0.2565 7.4700 1.3500 ;
      RECT 7.3360 0.2565 7.3620 1.3500 ;
      RECT 7.2280 0.2565 7.2540 1.3500 ;
      RECT 7.1200 0.2565 7.1460 1.3500 ;
      RECT 7.0120 0.2565 7.0380 1.3500 ;
      RECT 6.9040 0.2565 6.9300 1.3500 ;
      RECT 6.7960 0.2565 6.8220 1.3500 ;
      RECT 6.6880 0.2565 6.7140 1.3500 ;
      RECT 6.5800 0.2565 6.6060 1.3500 ;
      RECT 6.4720 0.2565 6.4980 1.3500 ;
      RECT 6.3640 0.2565 6.3900 1.3500 ;
      RECT 6.2560 0.2565 6.2820 1.3500 ;
      RECT 6.1480 0.2565 6.1740 1.3500 ;
      RECT 6.0400 0.2565 6.0660 1.3500 ;
      RECT 5.9320 0.2565 5.9580 1.3500 ;
      RECT 5.8240 0.2565 5.8500 1.3500 ;
      RECT 5.7160 0.2565 5.7420 1.3500 ;
      RECT 5.6080 0.2565 5.6340 1.3500 ;
      RECT 5.5000 0.2565 5.5260 1.3500 ;
      RECT 5.3920 0.2565 5.4180 1.3500 ;
      RECT 5.2840 0.2565 5.3100 1.3500 ;
      RECT 5.1760 0.2565 5.2020 1.3500 ;
      RECT 5.0680 0.2565 5.0940 1.3500 ;
      RECT 4.9600 0.2565 4.9860 1.3500 ;
      RECT 4.8520 0.2565 4.8780 1.3500 ;
      RECT 4.7440 0.2565 4.7700 1.3500 ;
      RECT 4.6360 0.2565 4.6620 1.3500 ;
      RECT 4.5280 0.2565 4.5540 1.3500 ;
      RECT 4.4200 0.2565 4.4460 1.3500 ;
      RECT 4.3120 0.2565 4.3380 1.3500 ;
      RECT 4.2040 0.2565 4.2300 1.3500 ;
      RECT 4.0960 0.2565 4.1220 1.3500 ;
      RECT 3.9880 0.2565 4.0140 1.3500 ;
      RECT 3.8800 0.2565 3.9060 1.3500 ;
      RECT 3.7720 0.2565 3.7980 1.3500 ;
      RECT 3.6640 0.2565 3.6900 1.3500 ;
      RECT 3.5560 0.2565 3.5820 1.3500 ;
      RECT 3.4480 0.2565 3.4740 1.3500 ;
      RECT 3.3400 0.2565 3.3660 1.3500 ;
      RECT 3.2320 0.2565 3.2580 1.3500 ;
      RECT 3.1240 0.2565 3.1500 1.3500 ;
      RECT 3.0160 0.2565 3.0420 1.3500 ;
      RECT 2.9080 0.2565 2.9340 1.3500 ;
      RECT 2.8000 0.2565 2.8260 1.3500 ;
      RECT 2.6920 0.2565 2.7180 1.3500 ;
      RECT 2.5840 0.2565 2.6100 1.3500 ;
      RECT 2.4760 0.2565 2.5020 1.3500 ;
      RECT 2.3680 0.2565 2.3940 1.3500 ;
      RECT 2.2600 0.2565 2.2860 1.3500 ;
      RECT 2.1520 0.2565 2.1780 1.3500 ;
      RECT 2.0440 0.2565 2.0700 1.3500 ;
      RECT 1.9360 0.2565 1.9620 1.3500 ;
      RECT 1.8280 0.2565 1.8540 1.3500 ;
      RECT 1.7200 0.2565 1.7460 1.3500 ;
      RECT 1.6120 0.2565 1.6380 1.3500 ;
      RECT 1.5040 0.2565 1.5300 1.3500 ;
      RECT 1.3960 0.2565 1.4220 1.3500 ;
      RECT 1.2880 0.2565 1.3140 1.3500 ;
      RECT 1.1800 0.2565 1.2060 1.3500 ;
      RECT 1.0720 0.2565 1.0980 1.3500 ;
      RECT 0.9640 0.2565 0.9900 1.3500 ;
      RECT 0.8560 0.2565 0.8820 1.3500 ;
      RECT 0.7480 0.2565 0.7740 1.3500 ;
      RECT 0.6400 0.2565 0.6660 1.3500 ;
      RECT 0.5320 0.2565 0.5580 1.3500 ;
      RECT 0.4240 0.2565 0.4500 1.3500 ;
      RECT 0.3160 0.2565 0.3420 1.3500 ;
      RECT 0.2080 0.2565 0.2340 1.3500 ;
      RECT 0.0050 0.2565 0.0900 1.3500 ;
      RECT 15.5530 1.3365 15.6810 2.4300 ;
      RECT 15.5390 2.0020 15.6810 2.3245 ;
      RECT 15.3190 1.7290 15.4530 2.4300 ;
      RECT 15.2960 2.0640 15.4530 2.3220 ;
      RECT 15.3190 1.3365 15.4170 2.4300 ;
      RECT 15.3190 1.4575 15.4310 1.6970 ;
      RECT 15.3190 1.3365 15.4530 1.4255 ;
      RECT 15.0940 1.7870 15.2280 2.4300 ;
      RECT 15.0940 1.3365 15.1920 2.4300 ;
      RECT 14.6770 1.3365 14.7600 2.4300 ;
      RECT 14.6770 1.4250 14.7740 2.3605 ;
      RECT 30.2680 1.3365 30.3530 2.4300 ;
      RECT 30.1240 1.3365 30.1500 2.4300 ;
      RECT 30.0160 1.3365 30.0420 2.4300 ;
      RECT 29.9080 1.3365 29.9340 2.4300 ;
      RECT 29.8000 1.3365 29.8260 2.4300 ;
      RECT 29.6920 1.3365 29.7180 2.4300 ;
      RECT 29.5840 1.3365 29.6100 2.4300 ;
      RECT 29.4760 1.3365 29.5020 2.4300 ;
      RECT 29.3680 1.3365 29.3940 2.4300 ;
      RECT 29.2600 1.3365 29.2860 2.4300 ;
      RECT 29.1520 1.3365 29.1780 2.4300 ;
      RECT 29.0440 1.3365 29.0700 2.4300 ;
      RECT 28.9360 1.3365 28.9620 2.4300 ;
      RECT 28.8280 1.3365 28.8540 2.4300 ;
      RECT 28.7200 1.3365 28.7460 2.4300 ;
      RECT 28.6120 1.3365 28.6380 2.4300 ;
      RECT 28.5040 1.3365 28.5300 2.4300 ;
      RECT 28.3960 1.3365 28.4220 2.4300 ;
      RECT 28.2880 1.3365 28.3140 2.4300 ;
      RECT 28.1800 1.3365 28.2060 2.4300 ;
      RECT 28.0720 1.3365 28.0980 2.4300 ;
      RECT 27.9640 1.3365 27.9900 2.4300 ;
      RECT 27.8560 1.3365 27.8820 2.4300 ;
      RECT 27.7480 1.3365 27.7740 2.4300 ;
      RECT 27.6400 1.3365 27.6660 2.4300 ;
      RECT 27.5320 1.3365 27.5580 2.4300 ;
      RECT 27.4240 1.3365 27.4500 2.4300 ;
      RECT 27.3160 1.3365 27.3420 2.4300 ;
      RECT 27.2080 1.3365 27.2340 2.4300 ;
      RECT 27.1000 1.3365 27.1260 2.4300 ;
      RECT 26.9920 1.3365 27.0180 2.4300 ;
      RECT 26.8840 1.3365 26.9100 2.4300 ;
      RECT 26.7760 1.3365 26.8020 2.4300 ;
      RECT 26.6680 1.3365 26.6940 2.4300 ;
      RECT 26.5600 1.3365 26.5860 2.4300 ;
      RECT 26.4520 1.3365 26.4780 2.4300 ;
      RECT 26.3440 1.3365 26.3700 2.4300 ;
      RECT 26.2360 1.3365 26.2620 2.4300 ;
      RECT 26.1280 1.3365 26.1540 2.4300 ;
      RECT 26.0200 1.3365 26.0460 2.4300 ;
      RECT 25.9120 1.3365 25.9380 2.4300 ;
      RECT 25.8040 1.3365 25.8300 2.4300 ;
      RECT 25.6960 1.3365 25.7220 2.4300 ;
      RECT 25.5880 1.3365 25.6140 2.4300 ;
      RECT 25.4800 1.3365 25.5060 2.4300 ;
      RECT 25.3720 1.3365 25.3980 2.4300 ;
      RECT 25.2640 1.3365 25.2900 2.4300 ;
      RECT 25.1560 1.3365 25.1820 2.4300 ;
      RECT 25.0480 1.3365 25.0740 2.4300 ;
      RECT 24.9400 1.3365 24.9660 2.4300 ;
      RECT 24.8320 1.3365 24.8580 2.4300 ;
      RECT 24.7240 1.3365 24.7500 2.4300 ;
      RECT 24.6160 1.3365 24.6420 2.4300 ;
      RECT 24.5080 1.3365 24.5340 2.4300 ;
      RECT 24.4000 1.3365 24.4260 2.4300 ;
      RECT 24.2920 1.3365 24.3180 2.4300 ;
      RECT 24.1840 1.3365 24.2100 2.4300 ;
      RECT 24.0760 1.3365 24.1020 2.4300 ;
      RECT 23.9680 1.3365 23.9940 2.4300 ;
      RECT 23.8600 1.3365 23.8860 2.4300 ;
      RECT 23.7520 1.3365 23.7780 2.4300 ;
      RECT 23.6440 1.3365 23.6700 2.4300 ;
      RECT 23.5360 1.3365 23.5620 2.4300 ;
      RECT 23.4280 1.3365 23.4540 2.4300 ;
      RECT 23.3200 1.3365 23.3460 2.4300 ;
      RECT 23.2120 1.3365 23.2380 2.4300 ;
      RECT 23.1040 1.3365 23.1300 2.4300 ;
      RECT 22.9960 1.3365 23.0220 2.4300 ;
      RECT 22.8880 1.3365 22.9140 2.4300 ;
      RECT 22.7800 1.3365 22.8060 2.4300 ;
      RECT 22.6720 1.3365 22.6980 2.4300 ;
      RECT 22.5640 1.3365 22.5900 2.4300 ;
      RECT 22.4560 1.3365 22.4820 2.4300 ;
      RECT 22.3480 1.3365 22.3740 2.4300 ;
      RECT 22.2400 1.3365 22.2660 2.4300 ;
      RECT 22.1320 1.3365 22.1580 2.4300 ;
      RECT 22.0240 1.3365 22.0500 2.4300 ;
      RECT 21.9160 1.3365 21.9420 2.4300 ;
      RECT 21.8080 1.3365 21.8340 2.4300 ;
      RECT 21.7000 1.3365 21.7260 2.4300 ;
      RECT 21.5920 1.3365 21.6180 2.4300 ;
      RECT 21.4840 1.3365 21.5100 2.4300 ;
      RECT 21.3760 1.3365 21.4020 2.4300 ;
      RECT 21.2680 1.3365 21.2940 2.4300 ;
      RECT 21.1600 1.3365 21.1860 2.4300 ;
      RECT 21.0520 1.3365 21.0780 2.4300 ;
      RECT 20.9440 1.3365 20.9700 2.4300 ;
      RECT 20.8360 1.3365 20.8620 2.4300 ;
      RECT 20.7280 1.3365 20.7540 2.4300 ;
      RECT 20.6200 1.3365 20.6460 2.4300 ;
      RECT 20.5120 1.3365 20.5380 2.4300 ;
      RECT 20.4040 1.3365 20.4300 2.4300 ;
      RECT 20.2960 1.3365 20.3220 2.4300 ;
      RECT 20.1880 1.3365 20.2140 2.4300 ;
      RECT 20.0800 1.3365 20.1060 2.4300 ;
      RECT 19.9720 1.3365 19.9980 2.4300 ;
      RECT 19.8640 1.3365 19.8900 2.4300 ;
      RECT 19.7560 1.3365 19.7820 2.4300 ;
      RECT 19.6480 1.3365 19.6740 2.4300 ;
      RECT 19.5400 1.3365 19.5660 2.4300 ;
      RECT 19.4320 1.3365 19.4580 2.4300 ;
      RECT 19.3240 1.3365 19.3500 2.4300 ;
      RECT 19.2160 1.3365 19.2420 2.4300 ;
      RECT 19.1080 1.3365 19.1340 2.4300 ;
      RECT 19.0000 1.3365 19.0260 2.4300 ;
      RECT 18.8920 1.3365 18.9180 2.4300 ;
      RECT 18.7840 1.3365 18.8100 2.4300 ;
      RECT 18.6760 1.3365 18.7020 2.4300 ;
      RECT 18.5680 1.3365 18.5940 2.4300 ;
      RECT 18.4600 1.3365 18.4860 2.4300 ;
      RECT 18.3520 1.3365 18.3780 2.4300 ;
      RECT 18.2440 1.3365 18.2700 2.4300 ;
      RECT 18.1360 1.3365 18.1620 2.4300 ;
      RECT 18.0280 1.3365 18.0540 2.4300 ;
      RECT 17.9200 1.3365 17.9460 2.4300 ;
      RECT 17.8120 1.3365 17.8380 2.4300 ;
      RECT 17.7040 1.3365 17.7300 2.4300 ;
      RECT 17.5960 1.3365 17.6220 2.4300 ;
      RECT 17.4880 1.3365 17.5140 2.4300 ;
      RECT 17.3800 1.3365 17.4060 2.4300 ;
      RECT 17.2720 1.3365 17.2980 2.4300 ;
      RECT 17.1640 1.3365 17.1900 2.4300 ;
      RECT 17.0560 1.3365 17.0820 2.4300 ;
      RECT 16.9480 1.3365 16.9740 2.4300 ;
      RECT 16.8400 1.3365 16.8660 2.4300 ;
      RECT 16.7320 1.3365 16.7580 2.4300 ;
      RECT 16.6240 1.3365 16.6500 2.4300 ;
      RECT 16.5160 1.3365 16.5420 2.4300 ;
      RECT 16.4080 1.3365 16.4340 2.4300 ;
      RECT 16.3000 1.3365 16.3260 2.4300 ;
      RECT 16.0870 1.3365 16.1640 2.4300 ;
      RECT 14.1940 1.3365 14.2710 2.4300 ;
      RECT 14.0320 1.3365 14.0580 2.4300 ;
      RECT 13.9240 1.3365 13.9500 2.4300 ;
      RECT 13.8160 1.3365 13.8420 2.4300 ;
      RECT 13.7080 1.3365 13.7340 2.4300 ;
      RECT 13.6000 1.3365 13.6260 2.4300 ;
      RECT 13.4920 1.3365 13.5180 2.4300 ;
      RECT 13.3840 1.3365 13.4100 2.4300 ;
      RECT 13.2760 1.3365 13.3020 2.4300 ;
      RECT 13.1680 1.3365 13.1940 2.4300 ;
      RECT 13.0600 1.3365 13.0860 2.4300 ;
      RECT 12.9520 1.3365 12.9780 2.4300 ;
      RECT 12.8440 1.3365 12.8700 2.4300 ;
      RECT 12.7360 1.3365 12.7620 2.4300 ;
      RECT 12.6280 1.3365 12.6540 2.4300 ;
      RECT 12.5200 1.3365 12.5460 2.4300 ;
      RECT 12.4120 1.3365 12.4380 2.4300 ;
      RECT 12.3040 1.3365 12.3300 2.4300 ;
      RECT 12.1960 1.3365 12.2220 2.4300 ;
      RECT 12.0880 1.3365 12.1140 2.4300 ;
      RECT 11.9800 1.3365 12.0060 2.4300 ;
      RECT 11.8720 1.3365 11.8980 2.4300 ;
      RECT 11.7640 1.3365 11.7900 2.4300 ;
      RECT 11.6560 1.3365 11.6820 2.4300 ;
      RECT 11.5480 1.3365 11.5740 2.4300 ;
      RECT 11.4400 1.3365 11.4660 2.4300 ;
      RECT 11.3320 1.3365 11.3580 2.4300 ;
      RECT 11.2240 1.3365 11.2500 2.4300 ;
      RECT 11.1160 1.3365 11.1420 2.4300 ;
      RECT 11.0080 1.3365 11.0340 2.4300 ;
      RECT 10.9000 1.3365 10.9260 2.4300 ;
      RECT 10.7920 1.3365 10.8180 2.4300 ;
      RECT 10.6840 1.3365 10.7100 2.4300 ;
      RECT 10.5760 1.3365 10.6020 2.4300 ;
      RECT 10.4680 1.3365 10.4940 2.4300 ;
      RECT 10.3600 1.3365 10.3860 2.4300 ;
      RECT 10.2520 1.3365 10.2780 2.4300 ;
      RECT 10.1440 1.3365 10.1700 2.4300 ;
      RECT 10.0360 1.3365 10.0620 2.4300 ;
      RECT 9.9280 1.3365 9.9540 2.4300 ;
      RECT 9.8200 1.3365 9.8460 2.4300 ;
      RECT 9.7120 1.3365 9.7380 2.4300 ;
      RECT 9.6040 1.3365 9.6300 2.4300 ;
      RECT 9.4960 1.3365 9.5220 2.4300 ;
      RECT 9.3880 1.3365 9.4140 2.4300 ;
      RECT 9.2800 1.3365 9.3060 2.4300 ;
      RECT 9.1720 1.3365 9.1980 2.4300 ;
      RECT 9.0640 1.3365 9.0900 2.4300 ;
      RECT 8.9560 1.3365 8.9820 2.4300 ;
      RECT 8.8480 1.3365 8.8740 2.4300 ;
      RECT 8.7400 1.3365 8.7660 2.4300 ;
      RECT 8.6320 1.3365 8.6580 2.4300 ;
      RECT 8.5240 1.3365 8.5500 2.4300 ;
      RECT 8.4160 1.3365 8.4420 2.4300 ;
      RECT 8.3080 1.3365 8.3340 2.4300 ;
      RECT 8.2000 1.3365 8.2260 2.4300 ;
      RECT 8.0920 1.3365 8.1180 2.4300 ;
      RECT 7.9840 1.3365 8.0100 2.4300 ;
      RECT 7.8760 1.3365 7.9020 2.4300 ;
      RECT 7.7680 1.3365 7.7940 2.4300 ;
      RECT 7.6600 1.3365 7.6860 2.4300 ;
      RECT 7.5520 1.3365 7.5780 2.4300 ;
      RECT 7.4440 1.3365 7.4700 2.4300 ;
      RECT 7.3360 1.3365 7.3620 2.4300 ;
      RECT 7.2280 1.3365 7.2540 2.4300 ;
      RECT 7.1200 1.3365 7.1460 2.4300 ;
      RECT 7.0120 1.3365 7.0380 2.4300 ;
      RECT 6.9040 1.3365 6.9300 2.4300 ;
      RECT 6.7960 1.3365 6.8220 2.4300 ;
      RECT 6.6880 1.3365 6.7140 2.4300 ;
      RECT 6.5800 1.3365 6.6060 2.4300 ;
      RECT 6.4720 1.3365 6.4980 2.4300 ;
      RECT 6.3640 1.3365 6.3900 2.4300 ;
      RECT 6.2560 1.3365 6.2820 2.4300 ;
      RECT 6.1480 1.3365 6.1740 2.4300 ;
      RECT 6.0400 1.3365 6.0660 2.4300 ;
      RECT 5.9320 1.3365 5.9580 2.4300 ;
      RECT 5.8240 1.3365 5.8500 2.4300 ;
      RECT 5.7160 1.3365 5.7420 2.4300 ;
      RECT 5.6080 1.3365 5.6340 2.4300 ;
      RECT 5.5000 1.3365 5.5260 2.4300 ;
      RECT 5.3920 1.3365 5.4180 2.4300 ;
      RECT 5.2840 1.3365 5.3100 2.4300 ;
      RECT 5.1760 1.3365 5.2020 2.4300 ;
      RECT 5.0680 1.3365 5.0940 2.4300 ;
      RECT 4.9600 1.3365 4.9860 2.4300 ;
      RECT 4.8520 1.3365 4.8780 2.4300 ;
      RECT 4.7440 1.3365 4.7700 2.4300 ;
      RECT 4.6360 1.3365 4.6620 2.4300 ;
      RECT 4.5280 1.3365 4.5540 2.4300 ;
      RECT 4.4200 1.3365 4.4460 2.4300 ;
      RECT 4.3120 1.3365 4.3380 2.4300 ;
      RECT 4.2040 1.3365 4.2300 2.4300 ;
      RECT 4.0960 1.3365 4.1220 2.4300 ;
      RECT 3.9880 1.3365 4.0140 2.4300 ;
      RECT 3.8800 1.3365 3.9060 2.4300 ;
      RECT 3.7720 1.3365 3.7980 2.4300 ;
      RECT 3.6640 1.3365 3.6900 2.4300 ;
      RECT 3.5560 1.3365 3.5820 2.4300 ;
      RECT 3.4480 1.3365 3.4740 2.4300 ;
      RECT 3.3400 1.3365 3.3660 2.4300 ;
      RECT 3.2320 1.3365 3.2580 2.4300 ;
      RECT 3.1240 1.3365 3.1500 2.4300 ;
      RECT 3.0160 1.3365 3.0420 2.4300 ;
      RECT 2.9080 1.3365 2.9340 2.4300 ;
      RECT 2.8000 1.3365 2.8260 2.4300 ;
      RECT 2.6920 1.3365 2.7180 2.4300 ;
      RECT 2.5840 1.3365 2.6100 2.4300 ;
      RECT 2.4760 1.3365 2.5020 2.4300 ;
      RECT 2.3680 1.3365 2.3940 2.4300 ;
      RECT 2.2600 1.3365 2.2860 2.4300 ;
      RECT 2.1520 1.3365 2.1780 2.4300 ;
      RECT 2.0440 1.3365 2.0700 2.4300 ;
      RECT 1.9360 1.3365 1.9620 2.4300 ;
      RECT 1.8280 1.3365 1.8540 2.4300 ;
      RECT 1.7200 1.3365 1.7460 2.4300 ;
      RECT 1.6120 1.3365 1.6380 2.4300 ;
      RECT 1.5040 1.3365 1.5300 2.4300 ;
      RECT 1.3960 1.3365 1.4220 2.4300 ;
      RECT 1.2880 1.3365 1.3140 2.4300 ;
      RECT 1.1800 1.3365 1.2060 2.4300 ;
      RECT 1.0720 1.3365 1.0980 2.4300 ;
      RECT 0.9640 1.3365 0.9900 2.4300 ;
      RECT 0.8560 1.3365 0.8820 2.4300 ;
      RECT 0.7480 1.3365 0.7740 2.4300 ;
      RECT 0.6400 1.3365 0.6660 2.4300 ;
      RECT 0.5320 1.3365 0.5580 2.4300 ;
      RECT 0.4240 1.3365 0.4500 2.4300 ;
      RECT 0.3160 1.3365 0.3420 2.4300 ;
      RECT 0.2080 1.3365 0.2340 2.4300 ;
      RECT 0.0050 1.3365 0.0900 2.4300 ;
      RECT 15.5530 2.4165 15.6810 3.5100 ;
      RECT 15.5390 3.0820 15.6810 3.4045 ;
      RECT 15.3190 2.8090 15.4530 3.5100 ;
      RECT 15.2960 3.1440 15.4530 3.4020 ;
      RECT 15.3190 2.4165 15.4170 3.5100 ;
      RECT 15.3190 2.5375 15.4310 2.7770 ;
      RECT 15.3190 2.4165 15.4530 2.5055 ;
      RECT 15.0940 2.8670 15.2280 3.5100 ;
      RECT 15.0940 2.4165 15.1920 3.5100 ;
      RECT 14.6770 2.4165 14.7600 3.5100 ;
      RECT 14.6770 2.5050 14.7740 3.4405 ;
      RECT 30.2680 2.4165 30.3530 3.5100 ;
      RECT 30.1240 2.4165 30.1500 3.5100 ;
      RECT 30.0160 2.4165 30.0420 3.5100 ;
      RECT 29.9080 2.4165 29.9340 3.5100 ;
      RECT 29.8000 2.4165 29.8260 3.5100 ;
      RECT 29.6920 2.4165 29.7180 3.5100 ;
      RECT 29.5840 2.4165 29.6100 3.5100 ;
      RECT 29.4760 2.4165 29.5020 3.5100 ;
      RECT 29.3680 2.4165 29.3940 3.5100 ;
      RECT 29.2600 2.4165 29.2860 3.5100 ;
      RECT 29.1520 2.4165 29.1780 3.5100 ;
      RECT 29.0440 2.4165 29.0700 3.5100 ;
      RECT 28.9360 2.4165 28.9620 3.5100 ;
      RECT 28.8280 2.4165 28.8540 3.5100 ;
      RECT 28.7200 2.4165 28.7460 3.5100 ;
      RECT 28.6120 2.4165 28.6380 3.5100 ;
      RECT 28.5040 2.4165 28.5300 3.5100 ;
      RECT 28.3960 2.4165 28.4220 3.5100 ;
      RECT 28.2880 2.4165 28.3140 3.5100 ;
      RECT 28.1800 2.4165 28.2060 3.5100 ;
      RECT 28.0720 2.4165 28.0980 3.5100 ;
      RECT 27.9640 2.4165 27.9900 3.5100 ;
      RECT 27.8560 2.4165 27.8820 3.5100 ;
      RECT 27.7480 2.4165 27.7740 3.5100 ;
      RECT 27.6400 2.4165 27.6660 3.5100 ;
      RECT 27.5320 2.4165 27.5580 3.5100 ;
      RECT 27.4240 2.4165 27.4500 3.5100 ;
      RECT 27.3160 2.4165 27.3420 3.5100 ;
      RECT 27.2080 2.4165 27.2340 3.5100 ;
      RECT 27.1000 2.4165 27.1260 3.5100 ;
      RECT 26.9920 2.4165 27.0180 3.5100 ;
      RECT 26.8840 2.4165 26.9100 3.5100 ;
      RECT 26.7760 2.4165 26.8020 3.5100 ;
      RECT 26.6680 2.4165 26.6940 3.5100 ;
      RECT 26.5600 2.4165 26.5860 3.5100 ;
      RECT 26.4520 2.4165 26.4780 3.5100 ;
      RECT 26.3440 2.4165 26.3700 3.5100 ;
      RECT 26.2360 2.4165 26.2620 3.5100 ;
      RECT 26.1280 2.4165 26.1540 3.5100 ;
      RECT 26.0200 2.4165 26.0460 3.5100 ;
      RECT 25.9120 2.4165 25.9380 3.5100 ;
      RECT 25.8040 2.4165 25.8300 3.5100 ;
      RECT 25.6960 2.4165 25.7220 3.5100 ;
      RECT 25.5880 2.4165 25.6140 3.5100 ;
      RECT 25.4800 2.4165 25.5060 3.5100 ;
      RECT 25.3720 2.4165 25.3980 3.5100 ;
      RECT 25.2640 2.4165 25.2900 3.5100 ;
      RECT 25.1560 2.4165 25.1820 3.5100 ;
      RECT 25.0480 2.4165 25.0740 3.5100 ;
      RECT 24.9400 2.4165 24.9660 3.5100 ;
      RECT 24.8320 2.4165 24.8580 3.5100 ;
      RECT 24.7240 2.4165 24.7500 3.5100 ;
      RECT 24.6160 2.4165 24.6420 3.5100 ;
      RECT 24.5080 2.4165 24.5340 3.5100 ;
      RECT 24.4000 2.4165 24.4260 3.5100 ;
      RECT 24.2920 2.4165 24.3180 3.5100 ;
      RECT 24.1840 2.4165 24.2100 3.5100 ;
      RECT 24.0760 2.4165 24.1020 3.5100 ;
      RECT 23.9680 2.4165 23.9940 3.5100 ;
      RECT 23.8600 2.4165 23.8860 3.5100 ;
      RECT 23.7520 2.4165 23.7780 3.5100 ;
      RECT 23.6440 2.4165 23.6700 3.5100 ;
      RECT 23.5360 2.4165 23.5620 3.5100 ;
      RECT 23.4280 2.4165 23.4540 3.5100 ;
      RECT 23.3200 2.4165 23.3460 3.5100 ;
      RECT 23.2120 2.4165 23.2380 3.5100 ;
      RECT 23.1040 2.4165 23.1300 3.5100 ;
      RECT 22.9960 2.4165 23.0220 3.5100 ;
      RECT 22.8880 2.4165 22.9140 3.5100 ;
      RECT 22.7800 2.4165 22.8060 3.5100 ;
      RECT 22.6720 2.4165 22.6980 3.5100 ;
      RECT 22.5640 2.4165 22.5900 3.5100 ;
      RECT 22.4560 2.4165 22.4820 3.5100 ;
      RECT 22.3480 2.4165 22.3740 3.5100 ;
      RECT 22.2400 2.4165 22.2660 3.5100 ;
      RECT 22.1320 2.4165 22.1580 3.5100 ;
      RECT 22.0240 2.4165 22.0500 3.5100 ;
      RECT 21.9160 2.4165 21.9420 3.5100 ;
      RECT 21.8080 2.4165 21.8340 3.5100 ;
      RECT 21.7000 2.4165 21.7260 3.5100 ;
      RECT 21.5920 2.4165 21.6180 3.5100 ;
      RECT 21.4840 2.4165 21.5100 3.5100 ;
      RECT 21.3760 2.4165 21.4020 3.5100 ;
      RECT 21.2680 2.4165 21.2940 3.5100 ;
      RECT 21.1600 2.4165 21.1860 3.5100 ;
      RECT 21.0520 2.4165 21.0780 3.5100 ;
      RECT 20.9440 2.4165 20.9700 3.5100 ;
      RECT 20.8360 2.4165 20.8620 3.5100 ;
      RECT 20.7280 2.4165 20.7540 3.5100 ;
      RECT 20.6200 2.4165 20.6460 3.5100 ;
      RECT 20.5120 2.4165 20.5380 3.5100 ;
      RECT 20.4040 2.4165 20.4300 3.5100 ;
      RECT 20.2960 2.4165 20.3220 3.5100 ;
      RECT 20.1880 2.4165 20.2140 3.5100 ;
      RECT 20.0800 2.4165 20.1060 3.5100 ;
      RECT 19.9720 2.4165 19.9980 3.5100 ;
      RECT 19.8640 2.4165 19.8900 3.5100 ;
      RECT 19.7560 2.4165 19.7820 3.5100 ;
      RECT 19.6480 2.4165 19.6740 3.5100 ;
      RECT 19.5400 2.4165 19.5660 3.5100 ;
      RECT 19.4320 2.4165 19.4580 3.5100 ;
      RECT 19.3240 2.4165 19.3500 3.5100 ;
      RECT 19.2160 2.4165 19.2420 3.5100 ;
      RECT 19.1080 2.4165 19.1340 3.5100 ;
      RECT 19.0000 2.4165 19.0260 3.5100 ;
      RECT 18.8920 2.4165 18.9180 3.5100 ;
      RECT 18.7840 2.4165 18.8100 3.5100 ;
      RECT 18.6760 2.4165 18.7020 3.5100 ;
      RECT 18.5680 2.4165 18.5940 3.5100 ;
      RECT 18.4600 2.4165 18.4860 3.5100 ;
      RECT 18.3520 2.4165 18.3780 3.5100 ;
      RECT 18.2440 2.4165 18.2700 3.5100 ;
      RECT 18.1360 2.4165 18.1620 3.5100 ;
      RECT 18.0280 2.4165 18.0540 3.5100 ;
      RECT 17.9200 2.4165 17.9460 3.5100 ;
      RECT 17.8120 2.4165 17.8380 3.5100 ;
      RECT 17.7040 2.4165 17.7300 3.5100 ;
      RECT 17.5960 2.4165 17.6220 3.5100 ;
      RECT 17.4880 2.4165 17.5140 3.5100 ;
      RECT 17.3800 2.4165 17.4060 3.5100 ;
      RECT 17.2720 2.4165 17.2980 3.5100 ;
      RECT 17.1640 2.4165 17.1900 3.5100 ;
      RECT 17.0560 2.4165 17.0820 3.5100 ;
      RECT 16.9480 2.4165 16.9740 3.5100 ;
      RECT 16.8400 2.4165 16.8660 3.5100 ;
      RECT 16.7320 2.4165 16.7580 3.5100 ;
      RECT 16.6240 2.4165 16.6500 3.5100 ;
      RECT 16.5160 2.4165 16.5420 3.5100 ;
      RECT 16.4080 2.4165 16.4340 3.5100 ;
      RECT 16.3000 2.4165 16.3260 3.5100 ;
      RECT 16.0870 2.4165 16.1640 3.5100 ;
      RECT 14.1940 2.4165 14.2710 3.5100 ;
      RECT 14.0320 2.4165 14.0580 3.5100 ;
      RECT 13.9240 2.4165 13.9500 3.5100 ;
      RECT 13.8160 2.4165 13.8420 3.5100 ;
      RECT 13.7080 2.4165 13.7340 3.5100 ;
      RECT 13.6000 2.4165 13.6260 3.5100 ;
      RECT 13.4920 2.4165 13.5180 3.5100 ;
      RECT 13.3840 2.4165 13.4100 3.5100 ;
      RECT 13.2760 2.4165 13.3020 3.5100 ;
      RECT 13.1680 2.4165 13.1940 3.5100 ;
      RECT 13.0600 2.4165 13.0860 3.5100 ;
      RECT 12.9520 2.4165 12.9780 3.5100 ;
      RECT 12.8440 2.4165 12.8700 3.5100 ;
      RECT 12.7360 2.4165 12.7620 3.5100 ;
      RECT 12.6280 2.4165 12.6540 3.5100 ;
      RECT 12.5200 2.4165 12.5460 3.5100 ;
      RECT 12.4120 2.4165 12.4380 3.5100 ;
      RECT 12.3040 2.4165 12.3300 3.5100 ;
      RECT 12.1960 2.4165 12.2220 3.5100 ;
      RECT 12.0880 2.4165 12.1140 3.5100 ;
      RECT 11.9800 2.4165 12.0060 3.5100 ;
      RECT 11.8720 2.4165 11.8980 3.5100 ;
      RECT 11.7640 2.4165 11.7900 3.5100 ;
      RECT 11.6560 2.4165 11.6820 3.5100 ;
      RECT 11.5480 2.4165 11.5740 3.5100 ;
      RECT 11.4400 2.4165 11.4660 3.5100 ;
      RECT 11.3320 2.4165 11.3580 3.5100 ;
      RECT 11.2240 2.4165 11.2500 3.5100 ;
      RECT 11.1160 2.4165 11.1420 3.5100 ;
      RECT 11.0080 2.4165 11.0340 3.5100 ;
      RECT 10.9000 2.4165 10.9260 3.5100 ;
      RECT 10.7920 2.4165 10.8180 3.5100 ;
      RECT 10.6840 2.4165 10.7100 3.5100 ;
      RECT 10.5760 2.4165 10.6020 3.5100 ;
      RECT 10.4680 2.4165 10.4940 3.5100 ;
      RECT 10.3600 2.4165 10.3860 3.5100 ;
      RECT 10.2520 2.4165 10.2780 3.5100 ;
      RECT 10.1440 2.4165 10.1700 3.5100 ;
      RECT 10.0360 2.4165 10.0620 3.5100 ;
      RECT 9.9280 2.4165 9.9540 3.5100 ;
      RECT 9.8200 2.4165 9.8460 3.5100 ;
      RECT 9.7120 2.4165 9.7380 3.5100 ;
      RECT 9.6040 2.4165 9.6300 3.5100 ;
      RECT 9.4960 2.4165 9.5220 3.5100 ;
      RECT 9.3880 2.4165 9.4140 3.5100 ;
      RECT 9.2800 2.4165 9.3060 3.5100 ;
      RECT 9.1720 2.4165 9.1980 3.5100 ;
      RECT 9.0640 2.4165 9.0900 3.5100 ;
      RECT 8.9560 2.4165 8.9820 3.5100 ;
      RECT 8.8480 2.4165 8.8740 3.5100 ;
      RECT 8.7400 2.4165 8.7660 3.5100 ;
      RECT 8.6320 2.4165 8.6580 3.5100 ;
      RECT 8.5240 2.4165 8.5500 3.5100 ;
      RECT 8.4160 2.4165 8.4420 3.5100 ;
      RECT 8.3080 2.4165 8.3340 3.5100 ;
      RECT 8.2000 2.4165 8.2260 3.5100 ;
      RECT 8.0920 2.4165 8.1180 3.5100 ;
      RECT 7.9840 2.4165 8.0100 3.5100 ;
      RECT 7.8760 2.4165 7.9020 3.5100 ;
      RECT 7.7680 2.4165 7.7940 3.5100 ;
      RECT 7.6600 2.4165 7.6860 3.5100 ;
      RECT 7.5520 2.4165 7.5780 3.5100 ;
      RECT 7.4440 2.4165 7.4700 3.5100 ;
      RECT 7.3360 2.4165 7.3620 3.5100 ;
      RECT 7.2280 2.4165 7.2540 3.5100 ;
      RECT 7.1200 2.4165 7.1460 3.5100 ;
      RECT 7.0120 2.4165 7.0380 3.5100 ;
      RECT 6.9040 2.4165 6.9300 3.5100 ;
      RECT 6.7960 2.4165 6.8220 3.5100 ;
      RECT 6.6880 2.4165 6.7140 3.5100 ;
      RECT 6.5800 2.4165 6.6060 3.5100 ;
      RECT 6.4720 2.4165 6.4980 3.5100 ;
      RECT 6.3640 2.4165 6.3900 3.5100 ;
      RECT 6.2560 2.4165 6.2820 3.5100 ;
      RECT 6.1480 2.4165 6.1740 3.5100 ;
      RECT 6.0400 2.4165 6.0660 3.5100 ;
      RECT 5.9320 2.4165 5.9580 3.5100 ;
      RECT 5.8240 2.4165 5.8500 3.5100 ;
      RECT 5.7160 2.4165 5.7420 3.5100 ;
      RECT 5.6080 2.4165 5.6340 3.5100 ;
      RECT 5.5000 2.4165 5.5260 3.5100 ;
      RECT 5.3920 2.4165 5.4180 3.5100 ;
      RECT 5.2840 2.4165 5.3100 3.5100 ;
      RECT 5.1760 2.4165 5.2020 3.5100 ;
      RECT 5.0680 2.4165 5.0940 3.5100 ;
      RECT 4.9600 2.4165 4.9860 3.5100 ;
      RECT 4.8520 2.4165 4.8780 3.5100 ;
      RECT 4.7440 2.4165 4.7700 3.5100 ;
      RECT 4.6360 2.4165 4.6620 3.5100 ;
      RECT 4.5280 2.4165 4.5540 3.5100 ;
      RECT 4.4200 2.4165 4.4460 3.5100 ;
      RECT 4.3120 2.4165 4.3380 3.5100 ;
      RECT 4.2040 2.4165 4.2300 3.5100 ;
      RECT 4.0960 2.4165 4.1220 3.5100 ;
      RECT 3.9880 2.4165 4.0140 3.5100 ;
      RECT 3.8800 2.4165 3.9060 3.5100 ;
      RECT 3.7720 2.4165 3.7980 3.5100 ;
      RECT 3.6640 2.4165 3.6900 3.5100 ;
      RECT 3.5560 2.4165 3.5820 3.5100 ;
      RECT 3.4480 2.4165 3.4740 3.5100 ;
      RECT 3.3400 2.4165 3.3660 3.5100 ;
      RECT 3.2320 2.4165 3.2580 3.5100 ;
      RECT 3.1240 2.4165 3.1500 3.5100 ;
      RECT 3.0160 2.4165 3.0420 3.5100 ;
      RECT 2.9080 2.4165 2.9340 3.5100 ;
      RECT 2.8000 2.4165 2.8260 3.5100 ;
      RECT 2.6920 2.4165 2.7180 3.5100 ;
      RECT 2.5840 2.4165 2.6100 3.5100 ;
      RECT 2.4760 2.4165 2.5020 3.5100 ;
      RECT 2.3680 2.4165 2.3940 3.5100 ;
      RECT 2.2600 2.4165 2.2860 3.5100 ;
      RECT 2.1520 2.4165 2.1780 3.5100 ;
      RECT 2.0440 2.4165 2.0700 3.5100 ;
      RECT 1.9360 2.4165 1.9620 3.5100 ;
      RECT 1.8280 2.4165 1.8540 3.5100 ;
      RECT 1.7200 2.4165 1.7460 3.5100 ;
      RECT 1.6120 2.4165 1.6380 3.5100 ;
      RECT 1.5040 2.4165 1.5300 3.5100 ;
      RECT 1.3960 2.4165 1.4220 3.5100 ;
      RECT 1.2880 2.4165 1.3140 3.5100 ;
      RECT 1.1800 2.4165 1.2060 3.5100 ;
      RECT 1.0720 2.4165 1.0980 3.5100 ;
      RECT 0.9640 2.4165 0.9900 3.5100 ;
      RECT 0.8560 2.4165 0.8820 3.5100 ;
      RECT 0.7480 2.4165 0.7740 3.5100 ;
      RECT 0.6400 2.4165 0.6660 3.5100 ;
      RECT 0.5320 2.4165 0.5580 3.5100 ;
      RECT 0.4240 2.4165 0.4500 3.5100 ;
      RECT 0.3160 2.4165 0.3420 3.5100 ;
      RECT 0.2080 2.4165 0.2340 3.5100 ;
      RECT 0.0050 2.4165 0.0900 3.5100 ;
      RECT 15.5530 3.4965 15.6810 4.5900 ;
      RECT 15.5390 4.1620 15.6810 4.4845 ;
      RECT 15.3190 3.8890 15.4530 4.5900 ;
      RECT 15.2960 4.2240 15.4530 4.4820 ;
      RECT 15.3190 3.4965 15.4170 4.5900 ;
      RECT 15.3190 3.6175 15.4310 3.8570 ;
      RECT 15.3190 3.4965 15.4530 3.5855 ;
      RECT 15.0940 3.9470 15.2280 4.5900 ;
      RECT 15.0940 3.4965 15.1920 4.5900 ;
      RECT 14.6770 3.4965 14.7600 4.5900 ;
      RECT 14.6770 3.5850 14.7740 4.5205 ;
      RECT 30.2680 3.4965 30.3530 4.5900 ;
      RECT 30.1240 3.4965 30.1500 4.5900 ;
      RECT 30.0160 3.4965 30.0420 4.5900 ;
      RECT 29.9080 3.4965 29.9340 4.5900 ;
      RECT 29.8000 3.4965 29.8260 4.5900 ;
      RECT 29.6920 3.4965 29.7180 4.5900 ;
      RECT 29.5840 3.4965 29.6100 4.5900 ;
      RECT 29.4760 3.4965 29.5020 4.5900 ;
      RECT 29.3680 3.4965 29.3940 4.5900 ;
      RECT 29.2600 3.4965 29.2860 4.5900 ;
      RECT 29.1520 3.4965 29.1780 4.5900 ;
      RECT 29.0440 3.4965 29.0700 4.5900 ;
      RECT 28.9360 3.4965 28.9620 4.5900 ;
      RECT 28.8280 3.4965 28.8540 4.5900 ;
      RECT 28.7200 3.4965 28.7460 4.5900 ;
      RECT 28.6120 3.4965 28.6380 4.5900 ;
      RECT 28.5040 3.4965 28.5300 4.5900 ;
      RECT 28.3960 3.4965 28.4220 4.5900 ;
      RECT 28.2880 3.4965 28.3140 4.5900 ;
      RECT 28.1800 3.4965 28.2060 4.5900 ;
      RECT 28.0720 3.4965 28.0980 4.5900 ;
      RECT 27.9640 3.4965 27.9900 4.5900 ;
      RECT 27.8560 3.4965 27.8820 4.5900 ;
      RECT 27.7480 3.4965 27.7740 4.5900 ;
      RECT 27.6400 3.4965 27.6660 4.5900 ;
      RECT 27.5320 3.4965 27.5580 4.5900 ;
      RECT 27.4240 3.4965 27.4500 4.5900 ;
      RECT 27.3160 3.4965 27.3420 4.5900 ;
      RECT 27.2080 3.4965 27.2340 4.5900 ;
      RECT 27.1000 3.4965 27.1260 4.5900 ;
      RECT 26.9920 3.4965 27.0180 4.5900 ;
      RECT 26.8840 3.4965 26.9100 4.5900 ;
      RECT 26.7760 3.4965 26.8020 4.5900 ;
      RECT 26.6680 3.4965 26.6940 4.5900 ;
      RECT 26.5600 3.4965 26.5860 4.5900 ;
      RECT 26.4520 3.4965 26.4780 4.5900 ;
      RECT 26.3440 3.4965 26.3700 4.5900 ;
      RECT 26.2360 3.4965 26.2620 4.5900 ;
      RECT 26.1280 3.4965 26.1540 4.5900 ;
      RECT 26.0200 3.4965 26.0460 4.5900 ;
      RECT 25.9120 3.4965 25.9380 4.5900 ;
      RECT 25.8040 3.4965 25.8300 4.5900 ;
      RECT 25.6960 3.4965 25.7220 4.5900 ;
      RECT 25.5880 3.4965 25.6140 4.5900 ;
      RECT 25.4800 3.4965 25.5060 4.5900 ;
      RECT 25.3720 3.4965 25.3980 4.5900 ;
      RECT 25.2640 3.4965 25.2900 4.5900 ;
      RECT 25.1560 3.4965 25.1820 4.5900 ;
      RECT 25.0480 3.4965 25.0740 4.5900 ;
      RECT 24.9400 3.4965 24.9660 4.5900 ;
      RECT 24.8320 3.4965 24.8580 4.5900 ;
      RECT 24.7240 3.4965 24.7500 4.5900 ;
      RECT 24.6160 3.4965 24.6420 4.5900 ;
      RECT 24.5080 3.4965 24.5340 4.5900 ;
      RECT 24.4000 3.4965 24.4260 4.5900 ;
      RECT 24.2920 3.4965 24.3180 4.5900 ;
      RECT 24.1840 3.4965 24.2100 4.5900 ;
      RECT 24.0760 3.4965 24.1020 4.5900 ;
      RECT 23.9680 3.4965 23.9940 4.5900 ;
      RECT 23.8600 3.4965 23.8860 4.5900 ;
      RECT 23.7520 3.4965 23.7780 4.5900 ;
      RECT 23.6440 3.4965 23.6700 4.5900 ;
      RECT 23.5360 3.4965 23.5620 4.5900 ;
      RECT 23.4280 3.4965 23.4540 4.5900 ;
      RECT 23.3200 3.4965 23.3460 4.5900 ;
      RECT 23.2120 3.4965 23.2380 4.5900 ;
      RECT 23.1040 3.4965 23.1300 4.5900 ;
      RECT 22.9960 3.4965 23.0220 4.5900 ;
      RECT 22.8880 3.4965 22.9140 4.5900 ;
      RECT 22.7800 3.4965 22.8060 4.5900 ;
      RECT 22.6720 3.4965 22.6980 4.5900 ;
      RECT 22.5640 3.4965 22.5900 4.5900 ;
      RECT 22.4560 3.4965 22.4820 4.5900 ;
      RECT 22.3480 3.4965 22.3740 4.5900 ;
      RECT 22.2400 3.4965 22.2660 4.5900 ;
      RECT 22.1320 3.4965 22.1580 4.5900 ;
      RECT 22.0240 3.4965 22.0500 4.5900 ;
      RECT 21.9160 3.4965 21.9420 4.5900 ;
      RECT 21.8080 3.4965 21.8340 4.5900 ;
      RECT 21.7000 3.4965 21.7260 4.5900 ;
      RECT 21.5920 3.4965 21.6180 4.5900 ;
      RECT 21.4840 3.4965 21.5100 4.5900 ;
      RECT 21.3760 3.4965 21.4020 4.5900 ;
      RECT 21.2680 3.4965 21.2940 4.5900 ;
      RECT 21.1600 3.4965 21.1860 4.5900 ;
      RECT 21.0520 3.4965 21.0780 4.5900 ;
      RECT 20.9440 3.4965 20.9700 4.5900 ;
      RECT 20.8360 3.4965 20.8620 4.5900 ;
      RECT 20.7280 3.4965 20.7540 4.5900 ;
      RECT 20.6200 3.4965 20.6460 4.5900 ;
      RECT 20.5120 3.4965 20.5380 4.5900 ;
      RECT 20.4040 3.4965 20.4300 4.5900 ;
      RECT 20.2960 3.4965 20.3220 4.5900 ;
      RECT 20.1880 3.4965 20.2140 4.5900 ;
      RECT 20.0800 3.4965 20.1060 4.5900 ;
      RECT 19.9720 3.4965 19.9980 4.5900 ;
      RECT 19.8640 3.4965 19.8900 4.5900 ;
      RECT 19.7560 3.4965 19.7820 4.5900 ;
      RECT 19.6480 3.4965 19.6740 4.5900 ;
      RECT 19.5400 3.4965 19.5660 4.5900 ;
      RECT 19.4320 3.4965 19.4580 4.5900 ;
      RECT 19.3240 3.4965 19.3500 4.5900 ;
      RECT 19.2160 3.4965 19.2420 4.5900 ;
      RECT 19.1080 3.4965 19.1340 4.5900 ;
      RECT 19.0000 3.4965 19.0260 4.5900 ;
      RECT 18.8920 3.4965 18.9180 4.5900 ;
      RECT 18.7840 3.4965 18.8100 4.5900 ;
      RECT 18.6760 3.4965 18.7020 4.5900 ;
      RECT 18.5680 3.4965 18.5940 4.5900 ;
      RECT 18.4600 3.4965 18.4860 4.5900 ;
      RECT 18.3520 3.4965 18.3780 4.5900 ;
      RECT 18.2440 3.4965 18.2700 4.5900 ;
      RECT 18.1360 3.4965 18.1620 4.5900 ;
      RECT 18.0280 3.4965 18.0540 4.5900 ;
      RECT 17.9200 3.4965 17.9460 4.5900 ;
      RECT 17.8120 3.4965 17.8380 4.5900 ;
      RECT 17.7040 3.4965 17.7300 4.5900 ;
      RECT 17.5960 3.4965 17.6220 4.5900 ;
      RECT 17.4880 3.4965 17.5140 4.5900 ;
      RECT 17.3800 3.4965 17.4060 4.5900 ;
      RECT 17.2720 3.4965 17.2980 4.5900 ;
      RECT 17.1640 3.4965 17.1900 4.5900 ;
      RECT 17.0560 3.4965 17.0820 4.5900 ;
      RECT 16.9480 3.4965 16.9740 4.5900 ;
      RECT 16.8400 3.4965 16.8660 4.5900 ;
      RECT 16.7320 3.4965 16.7580 4.5900 ;
      RECT 16.6240 3.4965 16.6500 4.5900 ;
      RECT 16.5160 3.4965 16.5420 4.5900 ;
      RECT 16.4080 3.4965 16.4340 4.5900 ;
      RECT 16.3000 3.4965 16.3260 4.5900 ;
      RECT 16.0870 3.4965 16.1640 4.5900 ;
      RECT 14.1940 3.4965 14.2710 4.5900 ;
      RECT 14.0320 3.4965 14.0580 4.5900 ;
      RECT 13.9240 3.4965 13.9500 4.5900 ;
      RECT 13.8160 3.4965 13.8420 4.5900 ;
      RECT 13.7080 3.4965 13.7340 4.5900 ;
      RECT 13.6000 3.4965 13.6260 4.5900 ;
      RECT 13.4920 3.4965 13.5180 4.5900 ;
      RECT 13.3840 3.4965 13.4100 4.5900 ;
      RECT 13.2760 3.4965 13.3020 4.5900 ;
      RECT 13.1680 3.4965 13.1940 4.5900 ;
      RECT 13.0600 3.4965 13.0860 4.5900 ;
      RECT 12.9520 3.4965 12.9780 4.5900 ;
      RECT 12.8440 3.4965 12.8700 4.5900 ;
      RECT 12.7360 3.4965 12.7620 4.5900 ;
      RECT 12.6280 3.4965 12.6540 4.5900 ;
      RECT 12.5200 3.4965 12.5460 4.5900 ;
      RECT 12.4120 3.4965 12.4380 4.5900 ;
      RECT 12.3040 3.4965 12.3300 4.5900 ;
      RECT 12.1960 3.4965 12.2220 4.5900 ;
      RECT 12.0880 3.4965 12.1140 4.5900 ;
      RECT 11.9800 3.4965 12.0060 4.5900 ;
      RECT 11.8720 3.4965 11.8980 4.5900 ;
      RECT 11.7640 3.4965 11.7900 4.5900 ;
      RECT 11.6560 3.4965 11.6820 4.5900 ;
      RECT 11.5480 3.4965 11.5740 4.5900 ;
      RECT 11.4400 3.4965 11.4660 4.5900 ;
      RECT 11.3320 3.4965 11.3580 4.5900 ;
      RECT 11.2240 3.4965 11.2500 4.5900 ;
      RECT 11.1160 3.4965 11.1420 4.5900 ;
      RECT 11.0080 3.4965 11.0340 4.5900 ;
      RECT 10.9000 3.4965 10.9260 4.5900 ;
      RECT 10.7920 3.4965 10.8180 4.5900 ;
      RECT 10.6840 3.4965 10.7100 4.5900 ;
      RECT 10.5760 3.4965 10.6020 4.5900 ;
      RECT 10.4680 3.4965 10.4940 4.5900 ;
      RECT 10.3600 3.4965 10.3860 4.5900 ;
      RECT 10.2520 3.4965 10.2780 4.5900 ;
      RECT 10.1440 3.4965 10.1700 4.5900 ;
      RECT 10.0360 3.4965 10.0620 4.5900 ;
      RECT 9.9280 3.4965 9.9540 4.5900 ;
      RECT 9.8200 3.4965 9.8460 4.5900 ;
      RECT 9.7120 3.4965 9.7380 4.5900 ;
      RECT 9.6040 3.4965 9.6300 4.5900 ;
      RECT 9.4960 3.4965 9.5220 4.5900 ;
      RECT 9.3880 3.4965 9.4140 4.5900 ;
      RECT 9.2800 3.4965 9.3060 4.5900 ;
      RECT 9.1720 3.4965 9.1980 4.5900 ;
      RECT 9.0640 3.4965 9.0900 4.5900 ;
      RECT 8.9560 3.4965 8.9820 4.5900 ;
      RECT 8.8480 3.4965 8.8740 4.5900 ;
      RECT 8.7400 3.4965 8.7660 4.5900 ;
      RECT 8.6320 3.4965 8.6580 4.5900 ;
      RECT 8.5240 3.4965 8.5500 4.5900 ;
      RECT 8.4160 3.4965 8.4420 4.5900 ;
      RECT 8.3080 3.4965 8.3340 4.5900 ;
      RECT 8.2000 3.4965 8.2260 4.5900 ;
      RECT 8.0920 3.4965 8.1180 4.5900 ;
      RECT 7.9840 3.4965 8.0100 4.5900 ;
      RECT 7.8760 3.4965 7.9020 4.5900 ;
      RECT 7.7680 3.4965 7.7940 4.5900 ;
      RECT 7.6600 3.4965 7.6860 4.5900 ;
      RECT 7.5520 3.4965 7.5780 4.5900 ;
      RECT 7.4440 3.4965 7.4700 4.5900 ;
      RECT 7.3360 3.4965 7.3620 4.5900 ;
      RECT 7.2280 3.4965 7.2540 4.5900 ;
      RECT 7.1200 3.4965 7.1460 4.5900 ;
      RECT 7.0120 3.4965 7.0380 4.5900 ;
      RECT 6.9040 3.4965 6.9300 4.5900 ;
      RECT 6.7960 3.4965 6.8220 4.5900 ;
      RECT 6.6880 3.4965 6.7140 4.5900 ;
      RECT 6.5800 3.4965 6.6060 4.5900 ;
      RECT 6.4720 3.4965 6.4980 4.5900 ;
      RECT 6.3640 3.4965 6.3900 4.5900 ;
      RECT 6.2560 3.4965 6.2820 4.5900 ;
      RECT 6.1480 3.4965 6.1740 4.5900 ;
      RECT 6.0400 3.4965 6.0660 4.5900 ;
      RECT 5.9320 3.4965 5.9580 4.5900 ;
      RECT 5.8240 3.4965 5.8500 4.5900 ;
      RECT 5.7160 3.4965 5.7420 4.5900 ;
      RECT 5.6080 3.4965 5.6340 4.5900 ;
      RECT 5.5000 3.4965 5.5260 4.5900 ;
      RECT 5.3920 3.4965 5.4180 4.5900 ;
      RECT 5.2840 3.4965 5.3100 4.5900 ;
      RECT 5.1760 3.4965 5.2020 4.5900 ;
      RECT 5.0680 3.4965 5.0940 4.5900 ;
      RECT 4.9600 3.4965 4.9860 4.5900 ;
      RECT 4.8520 3.4965 4.8780 4.5900 ;
      RECT 4.7440 3.4965 4.7700 4.5900 ;
      RECT 4.6360 3.4965 4.6620 4.5900 ;
      RECT 4.5280 3.4965 4.5540 4.5900 ;
      RECT 4.4200 3.4965 4.4460 4.5900 ;
      RECT 4.3120 3.4965 4.3380 4.5900 ;
      RECT 4.2040 3.4965 4.2300 4.5900 ;
      RECT 4.0960 3.4965 4.1220 4.5900 ;
      RECT 3.9880 3.4965 4.0140 4.5900 ;
      RECT 3.8800 3.4965 3.9060 4.5900 ;
      RECT 3.7720 3.4965 3.7980 4.5900 ;
      RECT 3.6640 3.4965 3.6900 4.5900 ;
      RECT 3.5560 3.4965 3.5820 4.5900 ;
      RECT 3.4480 3.4965 3.4740 4.5900 ;
      RECT 3.3400 3.4965 3.3660 4.5900 ;
      RECT 3.2320 3.4965 3.2580 4.5900 ;
      RECT 3.1240 3.4965 3.1500 4.5900 ;
      RECT 3.0160 3.4965 3.0420 4.5900 ;
      RECT 2.9080 3.4965 2.9340 4.5900 ;
      RECT 2.8000 3.4965 2.8260 4.5900 ;
      RECT 2.6920 3.4965 2.7180 4.5900 ;
      RECT 2.5840 3.4965 2.6100 4.5900 ;
      RECT 2.4760 3.4965 2.5020 4.5900 ;
      RECT 2.3680 3.4965 2.3940 4.5900 ;
      RECT 2.2600 3.4965 2.2860 4.5900 ;
      RECT 2.1520 3.4965 2.1780 4.5900 ;
      RECT 2.0440 3.4965 2.0700 4.5900 ;
      RECT 1.9360 3.4965 1.9620 4.5900 ;
      RECT 1.8280 3.4965 1.8540 4.5900 ;
      RECT 1.7200 3.4965 1.7460 4.5900 ;
      RECT 1.6120 3.4965 1.6380 4.5900 ;
      RECT 1.5040 3.4965 1.5300 4.5900 ;
      RECT 1.3960 3.4965 1.4220 4.5900 ;
      RECT 1.2880 3.4965 1.3140 4.5900 ;
      RECT 1.1800 3.4965 1.2060 4.5900 ;
      RECT 1.0720 3.4965 1.0980 4.5900 ;
      RECT 0.9640 3.4965 0.9900 4.5900 ;
      RECT 0.8560 3.4965 0.8820 4.5900 ;
      RECT 0.7480 3.4965 0.7740 4.5900 ;
      RECT 0.6400 3.4965 0.6660 4.5900 ;
      RECT 0.5320 3.4965 0.5580 4.5900 ;
      RECT 0.4240 3.4965 0.4500 4.5900 ;
      RECT 0.3160 3.4965 0.3420 4.5900 ;
      RECT 0.2080 3.4965 0.2340 4.5900 ;
      RECT 0.0050 3.4965 0.0900 4.5900 ;
      RECT 15.5530 4.5765 15.6810 5.6700 ;
      RECT 15.5390 5.2420 15.6810 5.5645 ;
      RECT 15.3190 4.9690 15.4530 5.6700 ;
      RECT 15.2960 5.3040 15.4530 5.5620 ;
      RECT 15.3190 4.5765 15.4170 5.6700 ;
      RECT 15.3190 4.6975 15.4310 4.9370 ;
      RECT 15.3190 4.5765 15.4530 4.6655 ;
      RECT 15.0940 5.0270 15.2280 5.6700 ;
      RECT 15.0940 4.5765 15.1920 5.6700 ;
      RECT 14.6770 4.5765 14.7600 5.6700 ;
      RECT 14.6770 4.6650 14.7740 5.6005 ;
      RECT 30.2680 4.5765 30.3530 5.6700 ;
      RECT 30.1240 4.5765 30.1500 5.6700 ;
      RECT 30.0160 4.5765 30.0420 5.6700 ;
      RECT 29.9080 4.5765 29.9340 5.6700 ;
      RECT 29.8000 4.5765 29.8260 5.6700 ;
      RECT 29.6920 4.5765 29.7180 5.6700 ;
      RECT 29.5840 4.5765 29.6100 5.6700 ;
      RECT 29.4760 4.5765 29.5020 5.6700 ;
      RECT 29.3680 4.5765 29.3940 5.6700 ;
      RECT 29.2600 4.5765 29.2860 5.6700 ;
      RECT 29.1520 4.5765 29.1780 5.6700 ;
      RECT 29.0440 4.5765 29.0700 5.6700 ;
      RECT 28.9360 4.5765 28.9620 5.6700 ;
      RECT 28.8280 4.5765 28.8540 5.6700 ;
      RECT 28.7200 4.5765 28.7460 5.6700 ;
      RECT 28.6120 4.5765 28.6380 5.6700 ;
      RECT 28.5040 4.5765 28.5300 5.6700 ;
      RECT 28.3960 4.5765 28.4220 5.6700 ;
      RECT 28.2880 4.5765 28.3140 5.6700 ;
      RECT 28.1800 4.5765 28.2060 5.6700 ;
      RECT 28.0720 4.5765 28.0980 5.6700 ;
      RECT 27.9640 4.5765 27.9900 5.6700 ;
      RECT 27.8560 4.5765 27.8820 5.6700 ;
      RECT 27.7480 4.5765 27.7740 5.6700 ;
      RECT 27.6400 4.5765 27.6660 5.6700 ;
      RECT 27.5320 4.5765 27.5580 5.6700 ;
      RECT 27.4240 4.5765 27.4500 5.6700 ;
      RECT 27.3160 4.5765 27.3420 5.6700 ;
      RECT 27.2080 4.5765 27.2340 5.6700 ;
      RECT 27.1000 4.5765 27.1260 5.6700 ;
      RECT 26.9920 4.5765 27.0180 5.6700 ;
      RECT 26.8840 4.5765 26.9100 5.6700 ;
      RECT 26.7760 4.5765 26.8020 5.6700 ;
      RECT 26.6680 4.5765 26.6940 5.6700 ;
      RECT 26.5600 4.5765 26.5860 5.6700 ;
      RECT 26.4520 4.5765 26.4780 5.6700 ;
      RECT 26.3440 4.5765 26.3700 5.6700 ;
      RECT 26.2360 4.5765 26.2620 5.6700 ;
      RECT 26.1280 4.5765 26.1540 5.6700 ;
      RECT 26.0200 4.5765 26.0460 5.6700 ;
      RECT 25.9120 4.5765 25.9380 5.6700 ;
      RECT 25.8040 4.5765 25.8300 5.6700 ;
      RECT 25.6960 4.5765 25.7220 5.6700 ;
      RECT 25.5880 4.5765 25.6140 5.6700 ;
      RECT 25.4800 4.5765 25.5060 5.6700 ;
      RECT 25.3720 4.5765 25.3980 5.6700 ;
      RECT 25.2640 4.5765 25.2900 5.6700 ;
      RECT 25.1560 4.5765 25.1820 5.6700 ;
      RECT 25.0480 4.5765 25.0740 5.6700 ;
      RECT 24.9400 4.5765 24.9660 5.6700 ;
      RECT 24.8320 4.5765 24.8580 5.6700 ;
      RECT 24.7240 4.5765 24.7500 5.6700 ;
      RECT 24.6160 4.5765 24.6420 5.6700 ;
      RECT 24.5080 4.5765 24.5340 5.6700 ;
      RECT 24.4000 4.5765 24.4260 5.6700 ;
      RECT 24.2920 4.5765 24.3180 5.6700 ;
      RECT 24.1840 4.5765 24.2100 5.6700 ;
      RECT 24.0760 4.5765 24.1020 5.6700 ;
      RECT 23.9680 4.5765 23.9940 5.6700 ;
      RECT 23.8600 4.5765 23.8860 5.6700 ;
      RECT 23.7520 4.5765 23.7780 5.6700 ;
      RECT 23.6440 4.5765 23.6700 5.6700 ;
      RECT 23.5360 4.5765 23.5620 5.6700 ;
      RECT 23.4280 4.5765 23.4540 5.6700 ;
      RECT 23.3200 4.5765 23.3460 5.6700 ;
      RECT 23.2120 4.5765 23.2380 5.6700 ;
      RECT 23.1040 4.5765 23.1300 5.6700 ;
      RECT 22.9960 4.5765 23.0220 5.6700 ;
      RECT 22.8880 4.5765 22.9140 5.6700 ;
      RECT 22.7800 4.5765 22.8060 5.6700 ;
      RECT 22.6720 4.5765 22.6980 5.6700 ;
      RECT 22.5640 4.5765 22.5900 5.6700 ;
      RECT 22.4560 4.5765 22.4820 5.6700 ;
      RECT 22.3480 4.5765 22.3740 5.6700 ;
      RECT 22.2400 4.5765 22.2660 5.6700 ;
      RECT 22.1320 4.5765 22.1580 5.6700 ;
      RECT 22.0240 4.5765 22.0500 5.6700 ;
      RECT 21.9160 4.5765 21.9420 5.6700 ;
      RECT 21.8080 4.5765 21.8340 5.6700 ;
      RECT 21.7000 4.5765 21.7260 5.6700 ;
      RECT 21.5920 4.5765 21.6180 5.6700 ;
      RECT 21.4840 4.5765 21.5100 5.6700 ;
      RECT 21.3760 4.5765 21.4020 5.6700 ;
      RECT 21.2680 4.5765 21.2940 5.6700 ;
      RECT 21.1600 4.5765 21.1860 5.6700 ;
      RECT 21.0520 4.5765 21.0780 5.6700 ;
      RECT 20.9440 4.5765 20.9700 5.6700 ;
      RECT 20.8360 4.5765 20.8620 5.6700 ;
      RECT 20.7280 4.5765 20.7540 5.6700 ;
      RECT 20.6200 4.5765 20.6460 5.6700 ;
      RECT 20.5120 4.5765 20.5380 5.6700 ;
      RECT 20.4040 4.5765 20.4300 5.6700 ;
      RECT 20.2960 4.5765 20.3220 5.6700 ;
      RECT 20.1880 4.5765 20.2140 5.6700 ;
      RECT 20.0800 4.5765 20.1060 5.6700 ;
      RECT 19.9720 4.5765 19.9980 5.6700 ;
      RECT 19.8640 4.5765 19.8900 5.6700 ;
      RECT 19.7560 4.5765 19.7820 5.6700 ;
      RECT 19.6480 4.5765 19.6740 5.6700 ;
      RECT 19.5400 4.5765 19.5660 5.6700 ;
      RECT 19.4320 4.5765 19.4580 5.6700 ;
      RECT 19.3240 4.5765 19.3500 5.6700 ;
      RECT 19.2160 4.5765 19.2420 5.6700 ;
      RECT 19.1080 4.5765 19.1340 5.6700 ;
      RECT 19.0000 4.5765 19.0260 5.6700 ;
      RECT 18.8920 4.5765 18.9180 5.6700 ;
      RECT 18.7840 4.5765 18.8100 5.6700 ;
      RECT 18.6760 4.5765 18.7020 5.6700 ;
      RECT 18.5680 4.5765 18.5940 5.6700 ;
      RECT 18.4600 4.5765 18.4860 5.6700 ;
      RECT 18.3520 4.5765 18.3780 5.6700 ;
      RECT 18.2440 4.5765 18.2700 5.6700 ;
      RECT 18.1360 4.5765 18.1620 5.6700 ;
      RECT 18.0280 4.5765 18.0540 5.6700 ;
      RECT 17.9200 4.5765 17.9460 5.6700 ;
      RECT 17.8120 4.5765 17.8380 5.6700 ;
      RECT 17.7040 4.5765 17.7300 5.6700 ;
      RECT 17.5960 4.5765 17.6220 5.6700 ;
      RECT 17.4880 4.5765 17.5140 5.6700 ;
      RECT 17.3800 4.5765 17.4060 5.6700 ;
      RECT 17.2720 4.5765 17.2980 5.6700 ;
      RECT 17.1640 4.5765 17.1900 5.6700 ;
      RECT 17.0560 4.5765 17.0820 5.6700 ;
      RECT 16.9480 4.5765 16.9740 5.6700 ;
      RECT 16.8400 4.5765 16.8660 5.6700 ;
      RECT 16.7320 4.5765 16.7580 5.6700 ;
      RECT 16.6240 4.5765 16.6500 5.6700 ;
      RECT 16.5160 4.5765 16.5420 5.6700 ;
      RECT 16.4080 4.5765 16.4340 5.6700 ;
      RECT 16.3000 4.5765 16.3260 5.6700 ;
      RECT 16.0870 4.5765 16.1640 5.6700 ;
      RECT 14.1940 4.5765 14.2710 5.6700 ;
      RECT 14.0320 4.5765 14.0580 5.6700 ;
      RECT 13.9240 4.5765 13.9500 5.6700 ;
      RECT 13.8160 4.5765 13.8420 5.6700 ;
      RECT 13.7080 4.5765 13.7340 5.6700 ;
      RECT 13.6000 4.5765 13.6260 5.6700 ;
      RECT 13.4920 4.5765 13.5180 5.6700 ;
      RECT 13.3840 4.5765 13.4100 5.6700 ;
      RECT 13.2760 4.5765 13.3020 5.6700 ;
      RECT 13.1680 4.5765 13.1940 5.6700 ;
      RECT 13.0600 4.5765 13.0860 5.6700 ;
      RECT 12.9520 4.5765 12.9780 5.6700 ;
      RECT 12.8440 4.5765 12.8700 5.6700 ;
      RECT 12.7360 4.5765 12.7620 5.6700 ;
      RECT 12.6280 4.5765 12.6540 5.6700 ;
      RECT 12.5200 4.5765 12.5460 5.6700 ;
      RECT 12.4120 4.5765 12.4380 5.6700 ;
      RECT 12.3040 4.5765 12.3300 5.6700 ;
      RECT 12.1960 4.5765 12.2220 5.6700 ;
      RECT 12.0880 4.5765 12.1140 5.6700 ;
      RECT 11.9800 4.5765 12.0060 5.6700 ;
      RECT 11.8720 4.5765 11.8980 5.6700 ;
      RECT 11.7640 4.5765 11.7900 5.6700 ;
      RECT 11.6560 4.5765 11.6820 5.6700 ;
      RECT 11.5480 4.5765 11.5740 5.6700 ;
      RECT 11.4400 4.5765 11.4660 5.6700 ;
      RECT 11.3320 4.5765 11.3580 5.6700 ;
      RECT 11.2240 4.5765 11.2500 5.6700 ;
      RECT 11.1160 4.5765 11.1420 5.6700 ;
      RECT 11.0080 4.5765 11.0340 5.6700 ;
      RECT 10.9000 4.5765 10.9260 5.6700 ;
      RECT 10.7920 4.5765 10.8180 5.6700 ;
      RECT 10.6840 4.5765 10.7100 5.6700 ;
      RECT 10.5760 4.5765 10.6020 5.6700 ;
      RECT 10.4680 4.5765 10.4940 5.6700 ;
      RECT 10.3600 4.5765 10.3860 5.6700 ;
      RECT 10.2520 4.5765 10.2780 5.6700 ;
      RECT 10.1440 4.5765 10.1700 5.6700 ;
      RECT 10.0360 4.5765 10.0620 5.6700 ;
      RECT 9.9280 4.5765 9.9540 5.6700 ;
      RECT 9.8200 4.5765 9.8460 5.6700 ;
      RECT 9.7120 4.5765 9.7380 5.6700 ;
      RECT 9.6040 4.5765 9.6300 5.6700 ;
      RECT 9.4960 4.5765 9.5220 5.6700 ;
      RECT 9.3880 4.5765 9.4140 5.6700 ;
      RECT 9.2800 4.5765 9.3060 5.6700 ;
      RECT 9.1720 4.5765 9.1980 5.6700 ;
      RECT 9.0640 4.5765 9.0900 5.6700 ;
      RECT 8.9560 4.5765 8.9820 5.6700 ;
      RECT 8.8480 4.5765 8.8740 5.6700 ;
      RECT 8.7400 4.5765 8.7660 5.6700 ;
      RECT 8.6320 4.5765 8.6580 5.6700 ;
      RECT 8.5240 4.5765 8.5500 5.6700 ;
      RECT 8.4160 4.5765 8.4420 5.6700 ;
      RECT 8.3080 4.5765 8.3340 5.6700 ;
      RECT 8.2000 4.5765 8.2260 5.6700 ;
      RECT 8.0920 4.5765 8.1180 5.6700 ;
      RECT 7.9840 4.5765 8.0100 5.6700 ;
      RECT 7.8760 4.5765 7.9020 5.6700 ;
      RECT 7.7680 4.5765 7.7940 5.6700 ;
      RECT 7.6600 4.5765 7.6860 5.6700 ;
      RECT 7.5520 4.5765 7.5780 5.6700 ;
      RECT 7.4440 4.5765 7.4700 5.6700 ;
      RECT 7.3360 4.5765 7.3620 5.6700 ;
      RECT 7.2280 4.5765 7.2540 5.6700 ;
      RECT 7.1200 4.5765 7.1460 5.6700 ;
      RECT 7.0120 4.5765 7.0380 5.6700 ;
      RECT 6.9040 4.5765 6.9300 5.6700 ;
      RECT 6.7960 4.5765 6.8220 5.6700 ;
      RECT 6.6880 4.5765 6.7140 5.6700 ;
      RECT 6.5800 4.5765 6.6060 5.6700 ;
      RECT 6.4720 4.5765 6.4980 5.6700 ;
      RECT 6.3640 4.5765 6.3900 5.6700 ;
      RECT 6.2560 4.5765 6.2820 5.6700 ;
      RECT 6.1480 4.5765 6.1740 5.6700 ;
      RECT 6.0400 4.5765 6.0660 5.6700 ;
      RECT 5.9320 4.5765 5.9580 5.6700 ;
      RECT 5.8240 4.5765 5.8500 5.6700 ;
      RECT 5.7160 4.5765 5.7420 5.6700 ;
      RECT 5.6080 4.5765 5.6340 5.6700 ;
      RECT 5.5000 4.5765 5.5260 5.6700 ;
      RECT 5.3920 4.5765 5.4180 5.6700 ;
      RECT 5.2840 4.5765 5.3100 5.6700 ;
      RECT 5.1760 4.5765 5.2020 5.6700 ;
      RECT 5.0680 4.5765 5.0940 5.6700 ;
      RECT 4.9600 4.5765 4.9860 5.6700 ;
      RECT 4.8520 4.5765 4.8780 5.6700 ;
      RECT 4.7440 4.5765 4.7700 5.6700 ;
      RECT 4.6360 4.5765 4.6620 5.6700 ;
      RECT 4.5280 4.5765 4.5540 5.6700 ;
      RECT 4.4200 4.5765 4.4460 5.6700 ;
      RECT 4.3120 4.5765 4.3380 5.6700 ;
      RECT 4.2040 4.5765 4.2300 5.6700 ;
      RECT 4.0960 4.5765 4.1220 5.6700 ;
      RECT 3.9880 4.5765 4.0140 5.6700 ;
      RECT 3.8800 4.5765 3.9060 5.6700 ;
      RECT 3.7720 4.5765 3.7980 5.6700 ;
      RECT 3.6640 4.5765 3.6900 5.6700 ;
      RECT 3.5560 4.5765 3.5820 5.6700 ;
      RECT 3.4480 4.5765 3.4740 5.6700 ;
      RECT 3.3400 4.5765 3.3660 5.6700 ;
      RECT 3.2320 4.5765 3.2580 5.6700 ;
      RECT 3.1240 4.5765 3.1500 5.6700 ;
      RECT 3.0160 4.5765 3.0420 5.6700 ;
      RECT 2.9080 4.5765 2.9340 5.6700 ;
      RECT 2.8000 4.5765 2.8260 5.6700 ;
      RECT 2.6920 4.5765 2.7180 5.6700 ;
      RECT 2.5840 4.5765 2.6100 5.6700 ;
      RECT 2.4760 4.5765 2.5020 5.6700 ;
      RECT 2.3680 4.5765 2.3940 5.6700 ;
      RECT 2.2600 4.5765 2.2860 5.6700 ;
      RECT 2.1520 4.5765 2.1780 5.6700 ;
      RECT 2.0440 4.5765 2.0700 5.6700 ;
      RECT 1.9360 4.5765 1.9620 5.6700 ;
      RECT 1.8280 4.5765 1.8540 5.6700 ;
      RECT 1.7200 4.5765 1.7460 5.6700 ;
      RECT 1.6120 4.5765 1.6380 5.6700 ;
      RECT 1.5040 4.5765 1.5300 5.6700 ;
      RECT 1.3960 4.5765 1.4220 5.6700 ;
      RECT 1.2880 4.5765 1.3140 5.6700 ;
      RECT 1.1800 4.5765 1.2060 5.6700 ;
      RECT 1.0720 4.5765 1.0980 5.6700 ;
      RECT 0.9640 4.5765 0.9900 5.6700 ;
      RECT 0.8560 4.5765 0.8820 5.6700 ;
      RECT 0.7480 4.5765 0.7740 5.6700 ;
      RECT 0.6400 4.5765 0.6660 5.6700 ;
      RECT 0.5320 4.5765 0.5580 5.6700 ;
      RECT 0.4240 4.5765 0.4500 5.6700 ;
      RECT 0.3160 4.5765 0.3420 5.6700 ;
      RECT 0.2080 4.5765 0.2340 5.6700 ;
      RECT 0.0050 4.5765 0.0900 5.6700 ;
      RECT 15.5530 5.6565 15.6810 6.7500 ;
      RECT 15.5390 6.3220 15.6810 6.6445 ;
      RECT 15.3190 6.0490 15.4530 6.7500 ;
      RECT 15.2960 6.3840 15.4530 6.6420 ;
      RECT 15.3190 5.6565 15.4170 6.7500 ;
      RECT 15.3190 5.7775 15.4310 6.0170 ;
      RECT 15.3190 5.6565 15.4530 5.7455 ;
      RECT 15.0940 6.1070 15.2280 6.7500 ;
      RECT 15.0940 5.6565 15.1920 6.7500 ;
      RECT 14.6770 5.6565 14.7600 6.7500 ;
      RECT 14.6770 5.7450 14.7740 6.6805 ;
      RECT 30.2680 5.6565 30.3530 6.7500 ;
      RECT 30.1240 5.6565 30.1500 6.7500 ;
      RECT 30.0160 5.6565 30.0420 6.7500 ;
      RECT 29.9080 5.6565 29.9340 6.7500 ;
      RECT 29.8000 5.6565 29.8260 6.7500 ;
      RECT 29.6920 5.6565 29.7180 6.7500 ;
      RECT 29.5840 5.6565 29.6100 6.7500 ;
      RECT 29.4760 5.6565 29.5020 6.7500 ;
      RECT 29.3680 5.6565 29.3940 6.7500 ;
      RECT 29.2600 5.6565 29.2860 6.7500 ;
      RECT 29.1520 5.6565 29.1780 6.7500 ;
      RECT 29.0440 5.6565 29.0700 6.7500 ;
      RECT 28.9360 5.6565 28.9620 6.7500 ;
      RECT 28.8280 5.6565 28.8540 6.7500 ;
      RECT 28.7200 5.6565 28.7460 6.7500 ;
      RECT 28.6120 5.6565 28.6380 6.7500 ;
      RECT 28.5040 5.6565 28.5300 6.7500 ;
      RECT 28.3960 5.6565 28.4220 6.7500 ;
      RECT 28.2880 5.6565 28.3140 6.7500 ;
      RECT 28.1800 5.6565 28.2060 6.7500 ;
      RECT 28.0720 5.6565 28.0980 6.7500 ;
      RECT 27.9640 5.6565 27.9900 6.7500 ;
      RECT 27.8560 5.6565 27.8820 6.7500 ;
      RECT 27.7480 5.6565 27.7740 6.7500 ;
      RECT 27.6400 5.6565 27.6660 6.7500 ;
      RECT 27.5320 5.6565 27.5580 6.7500 ;
      RECT 27.4240 5.6565 27.4500 6.7500 ;
      RECT 27.3160 5.6565 27.3420 6.7500 ;
      RECT 27.2080 5.6565 27.2340 6.7500 ;
      RECT 27.1000 5.6565 27.1260 6.7500 ;
      RECT 26.9920 5.6565 27.0180 6.7500 ;
      RECT 26.8840 5.6565 26.9100 6.7500 ;
      RECT 26.7760 5.6565 26.8020 6.7500 ;
      RECT 26.6680 5.6565 26.6940 6.7500 ;
      RECT 26.5600 5.6565 26.5860 6.7500 ;
      RECT 26.4520 5.6565 26.4780 6.7500 ;
      RECT 26.3440 5.6565 26.3700 6.7500 ;
      RECT 26.2360 5.6565 26.2620 6.7500 ;
      RECT 26.1280 5.6565 26.1540 6.7500 ;
      RECT 26.0200 5.6565 26.0460 6.7500 ;
      RECT 25.9120 5.6565 25.9380 6.7500 ;
      RECT 25.8040 5.6565 25.8300 6.7500 ;
      RECT 25.6960 5.6565 25.7220 6.7500 ;
      RECT 25.5880 5.6565 25.6140 6.7500 ;
      RECT 25.4800 5.6565 25.5060 6.7500 ;
      RECT 25.3720 5.6565 25.3980 6.7500 ;
      RECT 25.2640 5.6565 25.2900 6.7500 ;
      RECT 25.1560 5.6565 25.1820 6.7500 ;
      RECT 25.0480 5.6565 25.0740 6.7500 ;
      RECT 24.9400 5.6565 24.9660 6.7500 ;
      RECT 24.8320 5.6565 24.8580 6.7500 ;
      RECT 24.7240 5.6565 24.7500 6.7500 ;
      RECT 24.6160 5.6565 24.6420 6.7500 ;
      RECT 24.5080 5.6565 24.5340 6.7500 ;
      RECT 24.4000 5.6565 24.4260 6.7500 ;
      RECT 24.2920 5.6565 24.3180 6.7500 ;
      RECT 24.1840 5.6565 24.2100 6.7500 ;
      RECT 24.0760 5.6565 24.1020 6.7500 ;
      RECT 23.9680 5.6565 23.9940 6.7500 ;
      RECT 23.8600 5.6565 23.8860 6.7500 ;
      RECT 23.7520 5.6565 23.7780 6.7500 ;
      RECT 23.6440 5.6565 23.6700 6.7500 ;
      RECT 23.5360 5.6565 23.5620 6.7500 ;
      RECT 23.4280 5.6565 23.4540 6.7500 ;
      RECT 23.3200 5.6565 23.3460 6.7500 ;
      RECT 23.2120 5.6565 23.2380 6.7500 ;
      RECT 23.1040 5.6565 23.1300 6.7500 ;
      RECT 22.9960 5.6565 23.0220 6.7500 ;
      RECT 22.8880 5.6565 22.9140 6.7500 ;
      RECT 22.7800 5.6565 22.8060 6.7500 ;
      RECT 22.6720 5.6565 22.6980 6.7500 ;
      RECT 22.5640 5.6565 22.5900 6.7500 ;
      RECT 22.4560 5.6565 22.4820 6.7500 ;
      RECT 22.3480 5.6565 22.3740 6.7500 ;
      RECT 22.2400 5.6565 22.2660 6.7500 ;
      RECT 22.1320 5.6565 22.1580 6.7500 ;
      RECT 22.0240 5.6565 22.0500 6.7500 ;
      RECT 21.9160 5.6565 21.9420 6.7500 ;
      RECT 21.8080 5.6565 21.8340 6.7500 ;
      RECT 21.7000 5.6565 21.7260 6.7500 ;
      RECT 21.5920 5.6565 21.6180 6.7500 ;
      RECT 21.4840 5.6565 21.5100 6.7500 ;
      RECT 21.3760 5.6565 21.4020 6.7500 ;
      RECT 21.2680 5.6565 21.2940 6.7500 ;
      RECT 21.1600 5.6565 21.1860 6.7500 ;
      RECT 21.0520 5.6565 21.0780 6.7500 ;
      RECT 20.9440 5.6565 20.9700 6.7500 ;
      RECT 20.8360 5.6565 20.8620 6.7500 ;
      RECT 20.7280 5.6565 20.7540 6.7500 ;
      RECT 20.6200 5.6565 20.6460 6.7500 ;
      RECT 20.5120 5.6565 20.5380 6.7500 ;
      RECT 20.4040 5.6565 20.4300 6.7500 ;
      RECT 20.2960 5.6565 20.3220 6.7500 ;
      RECT 20.1880 5.6565 20.2140 6.7500 ;
      RECT 20.0800 5.6565 20.1060 6.7500 ;
      RECT 19.9720 5.6565 19.9980 6.7500 ;
      RECT 19.8640 5.6565 19.8900 6.7500 ;
      RECT 19.7560 5.6565 19.7820 6.7500 ;
      RECT 19.6480 5.6565 19.6740 6.7500 ;
      RECT 19.5400 5.6565 19.5660 6.7500 ;
      RECT 19.4320 5.6565 19.4580 6.7500 ;
      RECT 19.3240 5.6565 19.3500 6.7500 ;
      RECT 19.2160 5.6565 19.2420 6.7500 ;
      RECT 19.1080 5.6565 19.1340 6.7500 ;
      RECT 19.0000 5.6565 19.0260 6.7500 ;
      RECT 18.8920 5.6565 18.9180 6.7500 ;
      RECT 18.7840 5.6565 18.8100 6.7500 ;
      RECT 18.6760 5.6565 18.7020 6.7500 ;
      RECT 18.5680 5.6565 18.5940 6.7500 ;
      RECT 18.4600 5.6565 18.4860 6.7500 ;
      RECT 18.3520 5.6565 18.3780 6.7500 ;
      RECT 18.2440 5.6565 18.2700 6.7500 ;
      RECT 18.1360 5.6565 18.1620 6.7500 ;
      RECT 18.0280 5.6565 18.0540 6.7500 ;
      RECT 17.9200 5.6565 17.9460 6.7500 ;
      RECT 17.8120 5.6565 17.8380 6.7500 ;
      RECT 17.7040 5.6565 17.7300 6.7500 ;
      RECT 17.5960 5.6565 17.6220 6.7500 ;
      RECT 17.4880 5.6565 17.5140 6.7500 ;
      RECT 17.3800 5.6565 17.4060 6.7500 ;
      RECT 17.2720 5.6565 17.2980 6.7500 ;
      RECT 17.1640 5.6565 17.1900 6.7500 ;
      RECT 17.0560 5.6565 17.0820 6.7500 ;
      RECT 16.9480 5.6565 16.9740 6.7500 ;
      RECT 16.8400 5.6565 16.8660 6.7500 ;
      RECT 16.7320 5.6565 16.7580 6.7500 ;
      RECT 16.6240 5.6565 16.6500 6.7500 ;
      RECT 16.5160 5.6565 16.5420 6.7500 ;
      RECT 16.4080 5.6565 16.4340 6.7500 ;
      RECT 16.3000 5.6565 16.3260 6.7500 ;
      RECT 16.0870 5.6565 16.1640 6.7500 ;
      RECT 14.1940 5.6565 14.2710 6.7500 ;
      RECT 14.0320 5.6565 14.0580 6.7500 ;
      RECT 13.9240 5.6565 13.9500 6.7500 ;
      RECT 13.8160 5.6565 13.8420 6.7500 ;
      RECT 13.7080 5.6565 13.7340 6.7500 ;
      RECT 13.6000 5.6565 13.6260 6.7500 ;
      RECT 13.4920 5.6565 13.5180 6.7500 ;
      RECT 13.3840 5.6565 13.4100 6.7500 ;
      RECT 13.2760 5.6565 13.3020 6.7500 ;
      RECT 13.1680 5.6565 13.1940 6.7500 ;
      RECT 13.0600 5.6565 13.0860 6.7500 ;
      RECT 12.9520 5.6565 12.9780 6.7500 ;
      RECT 12.8440 5.6565 12.8700 6.7500 ;
      RECT 12.7360 5.6565 12.7620 6.7500 ;
      RECT 12.6280 5.6565 12.6540 6.7500 ;
      RECT 12.5200 5.6565 12.5460 6.7500 ;
      RECT 12.4120 5.6565 12.4380 6.7500 ;
      RECT 12.3040 5.6565 12.3300 6.7500 ;
      RECT 12.1960 5.6565 12.2220 6.7500 ;
      RECT 12.0880 5.6565 12.1140 6.7500 ;
      RECT 11.9800 5.6565 12.0060 6.7500 ;
      RECT 11.8720 5.6565 11.8980 6.7500 ;
      RECT 11.7640 5.6565 11.7900 6.7500 ;
      RECT 11.6560 5.6565 11.6820 6.7500 ;
      RECT 11.5480 5.6565 11.5740 6.7500 ;
      RECT 11.4400 5.6565 11.4660 6.7500 ;
      RECT 11.3320 5.6565 11.3580 6.7500 ;
      RECT 11.2240 5.6565 11.2500 6.7500 ;
      RECT 11.1160 5.6565 11.1420 6.7500 ;
      RECT 11.0080 5.6565 11.0340 6.7500 ;
      RECT 10.9000 5.6565 10.9260 6.7500 ;
      RECT 10.7920 5.6565 10.8180 6.7500 ;
      RECT 10.6840 5.6565 10.7100 6.7500 ;
      RECT 10.5760 5.6565 10.6020 6.7500 ;
      RECT 10.4680 5.6565 10.4940 6.7500 ;
      RECT 10.3600 5.6565 10.3860 6.7500 ;
      RECT 10.2520 5.6565 10.2780 6.7500 ;
      RECT 10.1440 5.6565 10.1700 6.7500 ;
      RECT 10.0360 5.6565 10.0620 6.7500 ;
      RECT 9.9280 5.6565 9.9540 6.7500 ;
      RECT 9.8200 5.6565 9.8460 6.7500 ;
      RECT 9.7120 5.6565 9.7380 6.7500 ;
      RECT 9.6040 5.6565 9.6300 6.7500 ;
      RECT 9.4960 5.6565 9.5220 6.7500 ;
      RECT 9.3880 5.6565 9.4140 6.7500 ;
      RECT 9.2800 5.6565 9.3060 6.7500 ;
      RECT 9.1720 5.6565 9.1980 6.7500 ;
      RECT 9.0640 5.6565 9.0900 6.7500 ;
      RECT 8.9560 5.6565 8.9820 6.7500 ;
      RECT 8.8480 5.6565 8.8740 6.7500 ;
      RECT 8.7400 5.6565 8.7660 6.7500 ;
      RECT 8.6320 5.6565 8.6580 6.7500 ;
      RECT 8.5240 5.6565 8.5500 6.7500 ;
      RECT 8.4160 5.6565 8.4420 6.7500 ;
      RECT 8.3080 5.6565 8.3340 6.7500 ;
      RECT 8.2000 5.6565 8.2260 6.7500 ;
      RECT 8.0920 5.6565 8.1180 6.7500 ;
      RECT 7.9840 5.6565 8.0100 6.7500 ;
      RECT 7.8760 5.6565 7.9020 6.7500 ;
      RECT 7.7680 5.6565 7.7940 6.7500 ;
      RECT 7.6600 5.6565 7.6860 6.7500 ;
      RECT 7.5520 5.6565 7.5780 6.7500 ;
      RECT 7.4440 5.6565 7.4700 6.7500 ;
      RECT 7.3360 5.6565 7.3620 6.7500 ;
      RECT 7.2280 5.6565 7.2540 6.7500 ;
      RECT 7.1200 5.6565 7.1460 6.7500 ;
      RECT 7.0120 5.6565 7.0380 6.7500 ;
      RECT 6.9040 5.6565 6.9300 6.7500 ;
      RECT 6.7960 5.6565 6.8220 6.7500 ;
      RECT 6.6880 5.6565 6.7140 6.7500 ;
      RECT 6.5800 5.6565 6.6060 6.7500 ;
      RECT 6.4720 5.6565 6.4980 6.7500 ;
      RECT 6.3640 5.6565 6.3900 6.7500 ;
      RECT 6.2560 5.6565 6.2820 6.7500 ;
      RECT 6.1480 5.6565 6.1740 6.7500 ;
      RECT 6.0400 5.6565 6.0660 6.7500 ;
      RECT 5.9320 5.6565 5.9580 6.7500 ;
      RECT 5.8240 5.6565 5.8500 6.7500 ;
      RECT 5.7160 5.6565 5.7420 6.7500 ;
      RECT 5.6080 5.6565 5.6340 6.7500 ;
      RECT 5.5000 5.6565 5.5260 6.7500 ;
      RECT 5.3920 5.6565 5.4180 6.7500 ;
      RECT 5.2840 5.6565 5.3100 6.7500 ;
      RECT 5.1760 5.6565 5.2020 6.7500 ;
      RECT 5.0680 5.6565 5.0940 6.7500 ;
      RECT 4.9600 5.6565 4.9860 6.7500 ;
      RECT 4.8520 5.6565 4.8780 6.7500 ;
      RECT 4.7440 5.6565 4.7700 6.7500 ;
      RECT 4.6360 5.6565 4.6620 6.7500 ;
      RECT 4.5280 5.6565 4.5540 6.7500 ;
      RECT 4.4200 5.6565 4.4460 6.7500 ;
      RECT 4.3120 5.6565 4.3380 6.7500 ;
      RECT 4.2040 5.6565 4.2300 6.7500 ;
      RECT 4.0960 5.6565 4.1220 6.7500 ;
      RECT 3.9880 5.6565 4.0140 6.7500 ;
      RECT 3.8800 5.6565 3.9060 6.7500 ;
      RECT 3.7720 5.6565 3.7980 6.7500 ;
      RECT 3.6640 5.6565 3.6900 6.7500 ;
      RECT 3.5560 5.6565 3.5820 6.7500 ;
      RECT 3.4480 5.6565 3.4740 6.7500 ;
      RECT 3.3400 5.6565 3.3660 6.7500 ;
      RECT 3.2320 5.6565 3.2580 6.7500 ;
      RECT 3.1240 5.6565 3.1500 6.7500 ;
      RECT 3.0160 5.6565 3.0420 6.7500 ;
      RECT 2.9080 5.6565 2.9340 6.7500 ;
      RECT 2.8000 5.6565 2.8260 6.7500 ;
      RECT 2.6920 5.6565 2.7180 6.7500 ;
      RECT 2.5840 5.6565 2.6100 6.7500 ;
      RECT 2.4760 5.6565 2.5020 6.7500 ;
      RECT 2.3680 5.6565 2.3940 6.7500 ;
      RECT 2.2600 5.6565 2.2860 6.7500 ;
      RECT 2.1520 5.6565 2.1780 6.7500 ;
      RECT 2.0440 5.6565 2.0700 6.7500 ;
      RECT 1.9360 5.6565 1.9620 6.7500 ;
      RECT 1.8280 5.6565 1.8540 6.7500 ;
      RECT 1.7200 5.6565 1.7460 6.7500 ;
      RECT 1.6120 5.6565 1.6380 6.7500 ;
      RECT 1.5040 5.6565 1.5300 6.7500 ;
      RECT 1.3960 5.6565 1.4220 6.7500 ;
      RECT 1.2880 5.6565 1.3140 6.7500 ;
      RECT 1.1800 5.6565 1.2060 6.7500 ;
      RECT 1.0720 5.6565 1.0980 6.7500 ;
      RECT 0.9640 5.6565 0.9900 6.7500 ;
      RECT 0.8560 5.6565 0.8820 6.7500 ;
      RECT 0.7480 5.6565 0.7740 6.7500 ;
      RECT 0.6400 5.6565 0.6660 6.7500 ;
      RECT 0.5320 5.6565 0.5580 6.7500 ;
      RECT 0.4240 5.6565 0.4500 6.7500 ;
      RECT 0.3160 5.6565 0.3420 6.7500 ;
      RECT 0.2080 5.6565 0.2340 6.7500 ;
      RECT 0.0050 5.6565 0.0900 6.7500 ;
      RECT 15.5530 6.7365 15.6810 7.8300 ;
      RECT 15.5390 7.4020 15.6810 7.7245 ;
      RECT 15.3190 7.1290 15.4530 7.8300 ;
      RECT 15.2960 7.4640 15.4530 7.7220 ;
      RECT 15.3190 6.7365 15.4170 7.8300 ;
      RECT 15.3190 6.8575 15.4310 7.0970 ;
      RECT 15.3190 6.7365 15.4530 6.8255 ;
      RECT 15.0940 7.1870 15.2280 7.8300 ;
      RECT 15.0940 6.7365 15.1920 7.8300 ;
      RECT 14.6770 6.7365 14.7600 7.8300 ;
      RECT 14.6770 6.8250 14.7740 7.7605 ;
      RECT 30.2680 6.7365 30.3530 7.8300 ;
      RECT 30.1240 6.7365 30.1500 7.8300 ;
      RECT 30.0160 6.7365 30.0420 7.8300 ;
      RECT 29.9080 6.7365 29.9340 7.8300 ;
      RECT 29.8000 6.7365 29.8260 7.8300 ;
      RECT 29.6920 6.7365 29.7180 7.8300 ;
      RECT 29.5840 6.7365 29.6100 7.8300 ;
      RECT 29.4760 6.7365 29.5020 7.8300 ;
      RECT 29.3680 6.7365 29.3940 7.8300 ;
      RECT 29.2600 6.7365 29.2860 7.8300 ;
      RECT 29.1520 6.7365 29.1780 7.8300 ;
      RECT 29.0440 6.7365 29.0700 7.8300 ;
      RECT 28.9360 6.7365 28.9620 7.8300 ;
      RECT 28.8280 6.7365 28.8540 7.8300 ;
      RECT 28.7200 6.7365 28.7460 7.8300 ;
      RECT 28.6120 6.7365 28.6380 7.8300 ;
      RECT 28.5040 6.7365 28.5300 7.8300 ;
      RECT 28.3960 6.7365 28.4220 7.8300 ;
      RECT 28.2880 6.7365 28.3140 7.8300 ;
      RECT 28.1800 6.7365 28.2060 7.8300 ;
      RECT 28.0720 6.7365 28.0980 7.8300 ;
      RECT 27.9640 6.7365 27.9900 7.8300 ;
      RECT 27.8560 6.7365 27.8820 7.8300 ;
      RECT 27.7480 6.7365 27.7740 7.8300 ;
      RECT 27.6400 6.7365 27.6660 7.8300 ;
      RECT 27.5320 6.7365 27.5580 7.8300 ;
      RECT 27.4240 6.7365 27.4500 7.8300 ;
      RECT 27.3160 6.7365 27.3420 7.8300 ;
      RECT 27.2080 6.7365 27.2340 7.8300 ;
      RECT 27.1000 6.7365 27.1260 7.8300 ;
      RECT 26.9920 6.7365 27.0180 7.8300 ;
      RECT 26.8840 6.7365 26.9100 7.8300 ;
      RECT 26.7760 6.7365 26.8020 7.8300 ;
      RECT 26.6680 6.7365 26.6940 7.8300 ;
      RECT 26.5600 6.7365 26.5860 7.8300 ;
      RECT 26.4520 6.7365 26.4780 7.8300 ;
      RECT 26.3440 6.7365 26.3700 7.8300 ;
      RECT 26.2360 6.7365 26.2620 7.8300 ;
      RECT 26.1280 6.7365 26.1540 7.8300 ;
      RECT 26.0200 6.7365 26.0460 7.8300 ;
      RECT 25.9120 6.7365 25.9380 7.8300 ;
      RECT 25.8040 6.7365 25.8300 7.8300 ;
      RECT 25.6960 6.7365 25.7220 7.8300 ;
      RECT 25.5880 6.7365 25.6140 7.8300 ;
      RECT 25.4800 6.7365 25.5060 7.8300 ;
      RECT 25.3720 6.7365 25.3980 7.8300 ;
      RECT 25.2640 6.7365 25.2900 7.8300 ;
      RECT 25.1560 6.7365 25.1820 7.8300 ;
      RECT 25.0480 6.7365 25.0740 7.8300 ;
      RECT 24.9400 6.7365 24.9660 7.8300 ;
      RECT 24.8320 6.7365 24.8580 7.8300 ;
      RECT 24.7240 6.7365 24.7500 7.8300 ;
      RECT 24.6160 6.7365 24.6420 7.8300 ;
      RECT 24.5080 6.7365 24.5340 7.8300 ;
      RECT 24.4000 6.7365 24.4260 7.8300 ;
      RECT 24.2920 6.7365 24.3180 7.8300 ;
      RECT 24.1840 6.7365 24.2100 7.8300 ;
      RECT 24.0760 6.7365 24.1020 7.8300 ;
      RECT 23.9680 6.7365 23.9940 7.8300 ;
      RECT 23.8600 6.7365 23.8860 7.8300 ;
      RECT 23.7520 6.7365 23.7780 7.8300 ;
      RECT 23.6440 6.7365 23.6700 7.8300 ;
      RECT 23.5360 6.7365 23.5620 7.8300 ;
      RECT 23.4280 6.7365 23.4540 7.8300 ;
      RECT 23.3200 6.7365 23.3460 7.8300 ;
      RECT 23.2120 6.7365 23.2380 7.8300 ;
      RECT 23.1040 6.7365 23.1300 7.8300 ;
      RECT 22.9960 6.7365 23.0220 7.8300 ;
      RECT 22.8880 6.7365 22.9140 7.8300 ;
      RECT 22.7800 6.7365 22.8060 7.8300 ;
      RECT 22.6720 6.7365 22.6980 7.8300 ;
      RECT 22.5640 6.7365 22.5900 7.8300 ;
      RECT 22.4560 6.7365 22.4820 7.8300 ;
      RECT 22.3480 6.7365 22.3740 7.8300 ;
      RECT 22.2400 6.7365 22.2660 7.8300 ;
      RECT 22.1320 6.7365 22.1580 7.8300 ;
      RECT 22.0240 6.7365 22.0500 7.8300 ;
      RECT 21.9160 6.7365 21.9420 7.8300 ;
      RECT 21.8080 6.7365 21.8340 7.8300 ;
      RECT 21.7000 6.7365 21.7260 7.8300 ;
      RECT 21.5920 6.7365 21.6180 7.8300 ;
      RECT 21.4840 6.7365 21.5100 7.8300 ;
      RECT 21.3760 6.7365 21.4020 7.8300 ;
      RECT 21.2680 6.7365 21.2940 7.8300 ;
      RECT 21.1600 6.7365 21.1860 7.8300 ;
      RECT 21.0520 6.7365 21.0780 7.8300 ;
      RECT 20.9440 6.7365 20.9700 7.8300 ;
      RECT 20.8360 6.7365 20.8620 7.8300 ;
      RECT 20.7280 6.7365 20.7540 7.8300 ;
      RECT 20.6200 6.7365 20.6460 7.8300 ;
      RECT 20.5120 6.7365 20.5380 7.8300 ;
      RECT 20.4040 6.7365 20.4300 7.8300 ;
      RECT 20.2960 6.7365 20.3220 7.8300 ;
      RECT 20.1880 6.7365 20.2140 7.8300 ;
      RECT 20.0800 6.7365 20.1060 7.8300 ;
      RECT 19.9720 6.7365 19.9980 7.8300 ;
      RECT 19.8640 6.7365 19.8900 7.8300 ;
      RECT 19.7560 6.7365 19.7820 7.8300 ;
      RECT 19.6480 6.7365 19.6740 7.8300 ;
      RECT 19.5400 6.7365 19.5660 7.8300 ;
      RECT 19.4320 6.7365 19.4580 7.8300 ;
      RECT 19.3240 6.7365 19.3500 7.8300 ;
      RECT 19.2160 6.7365 19.2420 7.8300 ;
      RECT 19.1080 6.7365 19.1340 7.8300 ;
      RECT 19.0000 6.7365 19.0260 7.8300 ;
      RECT 18.8920 6.7365 18.9180 7.8300 ;
      RECT 18.7840 6.7365 18.8100 7.8300 ;
      RECT 18.6760 6.7365 18.7020 7.8300 ;
      RECT 18.5680 6.7365 18.5940 7.8300 ;
      RECT 18.4600 6.7365 18.4860 7.8300 ;
      RECT 18.3520 6.7365 18.3780 7.8300 ;
      RECT 18.2440 6.7365 18.2700 7.8300 ;
      RECT 18.1360 6.7365 18.1620 7.8300 ;
      RECT 18.0280 6.7365 18.0540 7.8300 ;
      RECT 17.9200 6.7365 17.9460 7.8300 ;
      RECT 17.8120 6.7365 17.8380 7.8300 ;
      RECT 17.7040 6.7365 17.7300 7.8300 ;
      RECT 17.5960 6.7365 17.6220 7.8300 ;
      RECT 17.4880 6.7365 17.5140 7.8300 ;
      RECT 17.3800 6.7365 17.4060 7.8300 ;
      RECT 17.2720 6.7365 17.2980 7.8300 ;
      RECT 17.1640 6.7365 17.1900 7.8300 ;
      RECT 17.0560 6.7365 17.0820 7.8300 ;
      RECT 16.9480 6.7365 16.9740 7.8300 ;
      RECT 16.8400 6.7365 16.8660 7.8300 ;
      RECT 16.7320 6.7365 16.7580 7.8300 ;
      RECT 16.6240 6.7365 16.6500 7.8300 ;
      RECT 16.5160 6.7365 16.5420 7.8300 ;
      RECT 16.4080 6.7365 16.4340 7.8300 ;
      RECT 16.3000 6.7365 16.3260 7.8300 ;
      RECT 16.0870 6.7365 16.1640 7.8300 ;
      RECT 14.1940 6.7365 14.2710 7.8300 ;
      RECT 14.0320 6.7365 14.0580 7.8300 ;
      RECT 13.9240 6.7365 13.9500 7.8300 ;
      RECT 13.8160 6.7365 13.8420 7.8300 ;
      RECT 13.7080 6.7365 13.7340 7.8300 ;
      RECT 13.6000 6.7365 13.6260 7.8300 ;
      RECT 13.4920 6.7365 13.5180 7.8300 ;
      RECT 13.3840 6.7365 13.4100 7.8300 ;
      RECT 13.2760 6.7365 13.3020 7.8300 ;
      RECT 13.1680 6.7365 13.1940 7.8300 ;
      RECT 13.0600 6.7365 13.0860 7.8300 ;
      RECT 12.9520 6.7365 12.9780 7.8300 ;
      RECT 12.8440 6.7365 12.8700 7.8300 ;
      RECT 12.7360 6.7365 12.7620 7.8300 ;
      RECT 12.6280 6.7365 12.6540 7.8300 ;
      RECT 12.5200 6.7365 12.5460 7.8300 ;
      RECT 12.4120 6.7365 12.4380 7.8300 ;
      RECT 12.3040 6.7365 12.3300 7.8300 ;
      RECT 12.1960 6.7365 12.2220 7.8300 ;
      RECT 12.0880 6.7365 12.1140 7.8300 ;
      RECT 11.9800 6.7365 12.0060 7.8300 ;
      RECT 11.8720 6.7365 11.8980 7.8300 ;
      RECT 11.7640 6.7365 11.7900 7.8300 ;
      RECT 11.6560 6.7365 11.6820 7.8300 ;
      RECT 11.5480 6.7365 11.5740 7.8300 ;
      RECT 11.4400 6.7365 11.4660 7.8300 ;
      RECT 11.3320 6.7365 11.3580 7.8300 ;
      RECT 11.2240 6.7365 11.2500 7.8300 ;
      RECT 11.1160 6.7365 11.1420 7.8300 ;
      RECT 11.0080 6.7365 11.0340 7.8300 ;
      RECT 10.9000 6.7365 10.9260 7.8300 ;
      RECT 10.7920 6.7365 10.8180 7.8300 ;
      RECT 10.6840 6.7365 10.7100 7.8300 ;
      RECT 10.5760 6.7365 10.6020 7.8300 ;
      RECT 10.4680 6.7365 10.4940 7.8300 ;
      RECT 10.3600 6.7365 10.3860 7.8300 ;
      RECT 10.2520 6.7365 10.2780 7.8300 ;
      RECT 10.1440 6.7365 10.1700 7.8300 ;
      RECT 10.0360 6.7365 10.0620 7.8300 ;
      RECT 9.9280 6.7365 9.9540 7.8300 ;
      RECT 9.8200 6.7365 9.8460 7.8300 ;
      RECT 9.7120 6.7365 9.7380 7.8300 ;
      RECT 9.6040 6.7365 9.6300 7.8300 ;
      RECT 9.4960 6.7365 9.5220 7.8300 ;
      RECT 9.3880 6.7365 9.4140 7.8300 ;
      RECT 9.2800 6.7365 9.3060 7.8300 ;
      RECT 9.1720 6.7365 9.1980 7.8300 ;
      RECT 9.0640 6.7365 9.0900 7.8300 ;
      RECT 8.9560 6.7365 8.9820 7.8300 ;
      RECT 8.8480 6.7365 8.8740 7.8300 ;
      RECT 8.7400 6.7365 8.7660 7.8300 ;
      RECT 8.6320 6.7365 8.6580 7.8300 ;
      RECT 8.5240 6.7365 8.5500 7.8300 ;
      RECT 8.4160 6.7365 8.4420 7.8300 ;
      RECT 8.3080 6.7365 8.3340 7.8300 ;
      RECT 8.2000 6.7365 8.2260 7.8300 ;
      RECT 8.0920 6.7365 8.1180 7.8300 ;
      RECT 7.9840 6.7365 8.0100 7.8300 ;
      RECT 7.8760 6.7365 7.9020 7.8300 ;
      RECT 7.7680 6.7365 7.7940 7.8300 ;
      RECT 7.6600 6.7365 7.6860 7.8300 ;
      RECT 7.5520 6.7365 7.5780 7.8300 ;
      RECT 7.4440 6.7365 7.4700 7.8300 ;
      RECT 7.3360 6.7365 7.3620 7.8300 ;
      RECT 7.2280 6.7365 7.2540 7.8300 ;
      RECT 7.1200 6.7365 7.1460 7.8300 ;
      RECT 7.0120 6.7365 7.0380 7.8300 ;
      RECT 6.9040 6.7365 6.9300 7.8300 ;
      RECT 6.7960 6.7365 6.8220 7.8300 ;
      RECT 6.6880 6.7365 6.7140 7.8300 ;
      RECT 6.5800 6.7365 6.6060 7.8300 ;
      RECT 6.4720 6.7365 6.4980 7.8300 ;
      RECT 6.3640 6.7365 6.3900 7.8300 ;
      RECT 6.2560 6.7365 6.2820 7.8300 ;
      RECT 6.1480 6.7365 6.1740 7.8300 ;
      RECT 6.0400 6.7365 6.0660 7.8300 ;
      RECT 5.9320 6.7365 5.9580 7.8300 ;
      RECT 5.8240 6.7365 5.8500 7.8300 ;
      RECT 5.7160 6.7365 5.7420 7.8300 ;
      RECT 5.6080 6.7365 5.6340 7.8300 ;
      RECT 5.5000 6.7365 5.5260 7.8300 ;
      RECT 5.3920 6.7365 5.4180 7.8300 ;
      RECT 5.2840 6.7365 5.3100 7.8300 ;
      RECT 5.1760 6.7365 5.2020 7.8300 ;
      RECT 5.0680 6.7365 5.0940 7.8300 ;
      RECT 4.9600 6.7365 4.9860 7.8300 ;
      RECT 4.8520 6.7365 4.8780 7.8300 ;
      RECT 4.7440 6.7365 4.7700 7.8300 ;
      RECT 4.6360 6.7365 4.6620 7.8300 ;
      RECT 4.5280 6.7365 4.5540 7.8300 ;
      RECT 4.4200 6.7365 4.4460 7.8300 ;
      RECT 4.3120 6.7365 4.3380 7.8300 ;
      RECT 4.2040 6.7365 4.2300 7.8300 ;
      RECT 4.0960 6.7365 4.1220 7.8300 ;
      RECT 3.9880 6.7365 4.0140 7.8300 ;
      RECT 3.8800 6.7365 3.9060 7.8300 ;
      RECT 3.7720 6.7365 3.7980 7.8300 ;
      RECT 3.6640 6.7365 3.6900 7.8300 ;
      RECT 3.5560 6.7365 3.5820 7.8300 ;
      RECT 3.4480 6.7365 3.4740 7.8300 ;
      RECT 3.3400 6.7365 3.3660 7.8300 ;
      RECT 3.2320 6.7365 3.2580 7.8300 ;
      RECT 3.1240 6.7365 3.1500 7.8300 ;
      RECT 3.0160 6.7365 3.0420 7.8300 ;
      RECT 2.9080 6.7365 2.9340 7.8300 ;
      RECT 2.8000 6.7365 2.8260 7.8300 ;
      RECT 2.6920 6.7365 2.7180 7.8300 ;
      RECT 2.5840 6.7365 2.6100 7.8300 ;
      RECT 2.4760 6.7365 2.5020 7.8300 ;
      RECT 2.3680 6.7365 2.3940 7.8300 ;
      RECT 2.2600 6.7365 2.2860 7.8300 ;
      RECT 2.1520 6.7365 2.1780 7.8300 ;
      RECT 2.0440 6.7365 2.0700 7.8300 ;
      RECT 1.9360 6.7365 1.9620 7.8300 ;
      RECT 1.8280 6.7365 1.8540 7.8300 ;
      RECT 1.7200 6.7365 1.7460 7.8300 ;
      RECT 1.6120 6.7365 1.6380 7.8300 ;
      RECT 1.5040 6.7365 1.5300 7.8300 ;
      RECT 1.3960 6.7365 1.4220 7.8300 ;
      RECT 1.2880 6.7365 1.3140 7.8300 ;
      RECT 1.1800 6.7365 1.2060 7.8300 ;
      RECT 1.0720 6.7365 1.0980 7.8300 ;
      RECT 0.9640 6.7365 0.9900 7.8300 ;
      RECT 0.8560 6.7365 0.8820 7.8300 ;
      RECT 0.7480 6.7365 0.7740 7.8300 ;
      RECT 0.6400 6.7365 0.6660 7.8300 ;
      RECT 0.5320 6.7365 0.5580 7.8300 ;
      RECT 0.4240 6.7365 0.4500 7.8300 ;
      RECT 0.3160 6.7365 0.3420 7.8300 ;
      RECT 0.2080 6.7365 0.2340 7.8300 ;
      RECT 0.0050 6.7365 0.0900 7.8300 ;
      RECT 15.5530 7.8165 15.6810 8.9100 ;
      RECT 15.5390 8.4820 15.6810 8.8045 ;
      RECT 15.3190 8.2090 15.4530 8.9100 ;
      RECT 15.2960 8.5440 15.4530 8.8020 ;
      RECT 15.3190 7.8165 15.4170 8.9100 ;
      RECT 15.3190 7.9375 15.4310 8.1770 ;
      RECT 15.3190 7.8165 15.4530 7.9055 ;
      RECT 15.0940 8.2670 15.2280 8.9100 ;
      RECT 15.0940 7.8165 15.1920 8.9100 ;
      RECT 14.6770 7.8165 14.7600 8.9100 ;
      RECT 14.6770 7.9050 14.7740 8.8405 ;
      RECT 30.2680 7.8165 30.3530 8.9100 ;
      RECT 30.1240 7.8165 30.1500 8.9100 ;
      RECT 30.0160 7.8165 30.0420 8.9100 ;
      RECT 29.9080 7.8165 29.9340 8.9100 ;
      RECT 29.8000 7.8165 29.8260 8.9100 ;
      RECT 29.6920 7.8165 29.7180 8.9100 ;
      RECT 29.5840 7.8165 29.6100 8.9100 ;
      RECT 29.4760 7.8165 29.5020 8.9100 ;
      RECT 29.3680 7.8165 29.3940 8.9100 ;
      RECT 29.2600 7.8165 29.2860 8.9100 ;
      RECT 29.1520 7.8165 29.1780 8.9100 ;
      RECT 29.0440 7.8165 29.0700 8.9100 ;
      RECT 28.9360 7.8165 28.9620 8.9100 ;
      RECT 28.8280 7.8165 28.8540 8.9100 ;
      RECT 28.7200 7.8165 28.7460 8.9100 ;
      RECT 28.6120 7.8165 28.6380 8.9100 ;
      RECT 28.5040 7.8165 28.5300 8.9100 ;
      RECT 28.3960 7.8165 28.4220 8.9100 ;
      RECT 28.2880 7.8165 28.3140 8.9100 ;
      RECT 28.1800 7.8165 28.2060 8.9100 ;
      RECT 28.0720 7.8165 28.0980 8.9100 ;
      RECT 27.9640 7.8165 27.9900 8.9100 ;
      RECT 27.8560 7.8165 27.8820 8.9100 ;
      RECT 27.7480 7.8165 27.7740 8.9100 ;
      RECT 27.6400 7.8165 27.6660 8.9100 ;
      RECT 27.5320 7.8165 27.5580 8.9100 ;
      RECT 27.4240 7.8165 27.4500 8.9100 ;
      RECT 27.3160 7.8165 27.3420 8.9100 ;
      RECT 27.2080 7.8165 27.2340 8.9100 ;
      RECT 27.1000 7.8165 27.1260 8.9100 ;
      RECT 26.9920 7.8165 27.0180 8.9100 ;
      RECT 26.8840 7.8165 26.9100 8.9100 ;
      RECT 26.7760 7.8165 26.8020 8.9100 ;
      RECT 26.6680 7.8165 26.6940 8.9100 ;
      RECT 26.5600 7.8165 26.5860 8.9100 ;
      RECT 26.4520 7.8165 26.4780 8.9100 ;
      RECT 26.3440 7.8165 26.3700 8.9100 ;
      RECT 26.2360 7.8165 26.2620 8.9100 ;
      RECT 26.1280 7.8165 26.1540 8.9100 ;
      RECT 26.0200 7.8165 26.0460 8.9100 ;
      RECT 25.9120 7.8165 25.9380 8.9100 ;
      RECT 25.8040 7.8165 25.8300 8.9100 ;
      RECT 25.6960 7.8165 25.7220 8.9100 ;
      RECT 25.5880 7.8165 25.6140 8.9100 ;
      RECT 25.4800 7.8165 25.5060 8.9100 ;
      RECT 25.3720 7.8165 25.3980 8.9100 ;
      RECT 25.2640 7.8165 25.2900 8.9100 ;
      RECT 25.1560 7.8165 25.1820 8.9100 ;
      RECT 25.0480 7.8165 25.0740 8.9100 ;
      RECT 24.9400 7.8165 24.9660 8.9100 ;
      RECT 24.8320 7.8165 24.8580 8.9100 ;
      RECT 24.7240 7.8165 24.7500 8.9100 ;
      RECT 24.6160 7.8165 24.6420 8.9100 ;
      RECT 24.5080 7.8165 24.5340 8.9100 ;
      RECT 24.4000 7.8165 24.4260 8.9100 ;
      RECT 24.2920 7.8165 24.3180 8.9100 ;
      RECT 24.1840 7.8165 24.2100 8.9100 ;
      RECT 24.0760 7.8165 24.1020 8.9100 ;
      RECT 23.9680 7.8165 23.9940 8.9100 ;
      RECT 23.8600 7.8165 23.8860 8.9100 ;
      RECT 23.7520 7.8165 23.7780 8.9100 ;
      RECT 23.6440 7.8165 23.6700 8.9100 ;
      RECT 23.5360 7.8165 23.5620 8.9100 ;
      RECT 23.4280 7.8165 23.4540 8.9100 ;
      RECT 23.3200 7.8165 23.3460 8.9100 ;
      RECT 23.2120 7.8165 23.2380 8.9100 ;
      RECT 23.1040 7.8165 23.1300 8.9100 ;
      RECT 22.9960 7.8165 23.0220 8.9100 ;
      RECT 22.8880 7.8165 22.9140 8.9100 ;
      RECT 22.7800 7.8165 22.8060 8.9100 ;
      RECT 22.6720 7.8165 22.6980 8.9100 ;
      RECT 22.5640 7.8165 22.5900 8.9100 ;
      RECT 22.4560 7.8165 22.4820 8.9100 ;
      RECT 22.3480 7.8165 22.3740 8.9100 ;
      RECT 22.2400 7.8165 22.2660 8.9100 ;
      RECT 22.1320 7.8165 22.1580 8.9100 ;
      RECT 22.0240 7.8165 22.0500 8.9100 ;
      RECT 21.9160 7.8165 21.9420 8.9100 ;
      RECT 21.8080 7.8165 21.8340 8.9100 ;
      RECT 21.7000 7.8165 21.7260 8.9100 ;
      RECT 21.5920 7.8165 21.6180 8.9100 ;
      RECT 21.4840 7.8165 21.5100 8.9100 ;
      RECT 21.3760 7.8165 21.4020 8.9100 ;
      RECT 21.2680 7.8165 21.2940 8.9100 ;
      RECT 21.1600 7.8165 21.1860 8.9100 ;
      RECT 21.0520 7.8165 21.0780 8.9100 ;
      RECT 20.9440 7.8165 20.9700 8.9100 ;
      RECT 20.8360 7.8165 20.8620 8.9100 ;
      RECT 20.7280 7.8165 20.7540 8.9100 ;
      RECT 20.6200 7.8165 20.6460 8.9100 ;
      RECT 20.5120 7.8165 20.5380 8.9100 ;
      RECT 20.4040 7.8165 20.4300 8.9100 ;
      RECT 20.2960 7.8165 20.3220 8.9100 ;
      RECT 20.1880 7.8165 20.2140 8.9100 ;
      RECT 20.0800 7.8165 20.1060 8.9100 ;
      RECT 19.9720 7.8165 19.9980 8.9100 ;
      RECT 19.8640 7.8165 19.8900 8.9100 ;
      RECT 19.7560 7.8165 19.7820 8.9100 ;
      RECT 19.6480 7.8165 19.6740 8.9100 ;
      RECT 19.5400 7.8165 19.5660 8.9100 ;
      RECT 19.4320 7.8165 19.4580 8.9100 ;
      RECT 19.3240 7.8165 19.3500 8.9100 ;
      RECT 19.2160 7.8165 19.2420 8.9100 ;
      RECT 19.1080 7.8165 19.1340 8.9100 ;
      RECT 19.0000 7.8165 19.0260 8.9100 ;
      RECT 18.8920 7.8165 18.9180 8.9100 ;
      RECT 18.7840 7.8165 18.8100 8.9100 ;
      RECT 18.6760 7.8165 18.7020 8.9100 ;
      RECT 18.5680 7.8165 18.5940 8.9100 ;
      RECT 18.4600 7.8165 18.4860 8.9100 ;
      RECT 18.3520 7.8165 18.3780 8.9100 ;
      RECT 18.2440 7.8165 18.2700 8.9100 ;
      RECT 18.1360 7.8165 18.1620 8.9100 ;
      RECT 18.0280 7.8165 18.0540 8.9100 ;
      RECT 17.9200 7.8165 17.9460 8.9100 ;
      RECT 17.8120 7.8165 17.8380 8.9100 ;
      RECT 17.7040 7.8165 17.7300 8.9100 ;
      RECT 17.5960 7.8165 17.6220 8.9100 ;
      RECT 17.4880 7.8165 17.5140 8.9100 ;
      RECT 17.3800 7.8165 17.4060 8.9100 ;
      RECT 17.2720 7.8165 17.2980 8.9100 ;
      RECT 17.1640 7.8165 17.1900 8.9100 ;
      RECT 17.0560 7.8165 17.0820 8.9100 ;
      RECT 16.9480 7.8165 16.9740 8.9100 ;
      RECT 16.8400 7.8165 16.8660 8.9100 ;
      RECT 16.7320 7.8165 16.7580 8.9100 ;
      RECT 16.6240 7.8165 16.6500 8.9100 ;
      RECT 16.5160 7.8165 16.5420 8.9100 ;
      RECT 16.4080 7.8165 16.4340 8.9100 ;
      RECT 16.3000 7.8165 16.3260 8.9100 ;
      RECT 16.0870 7.8165 16.1640 8.9100 ;
      RECT 14.1940 7.8165 14.2710 8.9100 ;
      RECT 14.0320 7.8165 14.0580 8.9100 ;
      RECT 13.9240 7.8165 13.9500 8.9100 ;
      RECT 13.8160 7.8165 13.8420 8.9100 ;
      RECT 13.7080 7.8165 13.7340 8.9100 ;
      RECT 13.6000 7.8165 13.6260 8.9100 ;
      RECT 13.4920 7.8165 13.5180 8.9100 ;
      RECT 13.3840 7.8165 13.4100 8.9100 ;
      RECT 13.2760 7.8165 13.3020 8.9100 ;
      RECT 13.1680 7.8165 13.1940 8.9100 ;
      RECT 13.0600 7.8165 13.0860 8.9100 ;
      RECT 12.9520 7.8165 12.9780 8.9100 ;
      RECT 12.8440 7.8165 12.8700 8.9100 ;
      RECT 12.7360 7.8165 12.7620 8.9100 ;
      RECT 12.6280 7.8165 12.6540 8.9100 ;
      RECT 12.5200 7.8165 12.5460 8.9100 ;
      RECT 12.4120 7.8165 12.4380 8.9100 ;
      RECT 12.3040 7.8165 12.3300 8.9100 ;
      RECT 12.1960 7.8165 12.2220 8.9100 ;
      RECT 12.0880 7.8165 12.1140 8.9100 ;
      RECT 11.9800 7.8165 12.0060 8.9100 ;
      RECT 11.8720 7.8165 11.8980 8.9100 ;
      RECT 11.7640 7.8165 11.7900 8.9100 ;
      RECT 11.6560 7.8165 11.6820 8.9100 ;
      RECT 11.5480 7.8165 11.5740 8.9100 ;
      RECT 11.4400 7.8165 11.4660 8.9100 ;
      RECT 11.3320 7.8165 11.3580 8.9100 ;
      RECT 11.2240 7.8165 11.2500 8.9100 ;
      RECT 11.1160 7.8165 11.1420 8.9100 ;
      RECT 11.0080 7.8165 11.0340 8.9100 ;
      RECT 10.9000 7.8165 10.9260 8.9100 ;
      RECT 10.7920 7.8165 10.8180 8.9100 ;
      RECT 10.6840 7.8165 10.7100 8.9100 ;
      RECT 10.5760 7.8165 10.6020 8.9100 ;
      RECT 10.4680 7.8165 10.4940 8.9100 ;
      RECT 10.3600 7.8165 10.3860 8.9100 ;
      RECT 10.2520 7.8165 10.2780 8.9100 ;
      RECT 10.1440 7.8165 10.1700 8.9100 ;
      RECT 10.0360 7.8165 10.0620 8.9100 ;
      RECT 9.9280 7.8165 9.9540 8.9100 ;
      RECT 9.8200 7.8165 9.8460 8.9100 ;
      RECT 9.7120 7.8165 9.7380 8.9100 ;
      RECT 9.6040 7.8165 9.6300 8.9100 ;
      RECT 9.4960 7.8165 9.5220 8.9100 ;
      RECT 9.3880 7.8165 9.4140 8.9100 ;
      RECT 9.2800 7.8165 9.3060 8.9100 ;
      RECT 9.1720 7.8165 9.1980 8.9100 ;
      RECT 9.0640 7.8165 9.0900 8.9100 ;
      RECT 8.9560 7.8165 8.9820 8.9100 ;
      RECT 8.8480 7.8165 8.8740 8.9100 ;
      RECT 8.7400 7.8165 8.7660 8.9100 ;
      RECT 8.6320 7.8165 8.6580 8.9100 ;
      RECT 8.5240 7.8165 8.5500 8.9100 ;
      RECT 8.4160 7.8165 8.4420 8.9100 ;
      RECT 8.3080 7.8165 8.3340 8.9100 ;
      RECT 8.2000 7.8165 8.2260 8.9100 ;
      RECT 8.0920 7.8165 8.1180 8.9100 ;
      RECT 7.9840 7.8165 8.0100 8.9100 ;
      RECT 7.8760 7.8165 7.9020 8.9100 ;
      RECT 7.7680 7.8165 7.7940 8.9100 ;
      RECT 7.6600 7.8165 7.6860 8.9100 ;
      RECT 7.5520 7.8165 7.5780 8.9100 ;
      RECT 7.4440 7.8165 7.4700 8.9100 ;
      RECT 7.3360 7.8165 7.3620 8.9100 ;
      RECT 7.2280 7.8165 7.2540 8.9100 ;
      RECT 7.1200 7.8165 7.1460 8.9100 ;
      RECT 7.0120 7.8165 7.0380 8.9100 ;
      RECT 6.9040 7.8165 6.9300 8.9100 ;
      RECT 6.7960 7.8165 6.8220 8.9100 ;
      RECT 6.6880 7.8165 6.7140 8.9100 ;
      RECT 6.5800 7.8165 6.6060 8.9100 ;
      RECT 6.4720 7.8165 6.4980 8.9100 ;
      RECT 6.3640 7.8165 6.3900 8.9100 ;
      RECT 6.2560 7.8165 6.2820 8.9100 ;
      RECT 6.1480 7.8165 6.1740 8.9100 ;
      RECT 6.0400 7.8165 6.0660 8.9100 ;
      RECT 5.9320 7.8165 5.9580 8.9100 ;
      RECT 5.8240 7.8165 5.8500 8.9100 ;
      RECT 5.7160 7.8165 5.7420 8.9100 ;
      RECT 5.6080 7.8165 5.6340 8.9100 ;
      RECT 5.5000 7.8165 5.5260 8.9100 ;
      RECT 5.3920 7.8165 5.4180 8.9100 ;
      RECT 5.2840 7.8165 5.3100 8.9100 ;
      RECT 5.1760 7.8165 5.2020 8.9100 ;
      RECT 5.0680 7.8165 5.0940 8.9100 ;
      RECT 4.9600 7.8165 4.9860 8.9100 ;
      RECT 4.8520 7.8165 4.8780 8.9100 ;
      RECT 4.7440 7.8165 4.7700 8.9100 ;
      RECT 4.6360 7.8165 4.6620 8.9100 ;
      RECT 4.5280 7.8165 4.5540 8.9100 ;
      RECT 4.4200 7.8165 4.4460 8.9100 ;
      RECT 4.3120 7.8165 4.3380 8.9100 ;
      RECT 4.2040 7.8165 4.2300 8.9100 ;
      RECT 4.0960 7.8165 4.1220 8.9100 ;
      RECT 3.9880 7.8165 4.0140 8.9100 ;
      RECT 3.8800 7.8165 3.9060 8.9100 ;
      RECT 3.7720 7.8165 3.7980 8.9100 ;
      RECT 3.6640 7.8165 3.6900 8.9100 ;
      RECT 3.5560 7.8165 3.5820 8.9100 ;
      RECT 3.4480 7.8165 3.4740 8.9100 ;
      RECT 3.3400 7.8165 3.3660 8.9100 ;
      RECT 3.2320 7.8165 3.2580 8.9100 ;
      RECT 3.1240 7.8165 3.1500 8.9100 ;
      RECT 3.0160 7.8165 3.0420 8.9100 ;
      RECT 2.9080 7.8165 2.9340 8.9100 ;
      RECT 2.8000 7.8165 2.8260 8.9100 ;
      RECT 2.6920 7.8165 2.7180 8.9100 ;
      RECT 2.5840 7.8165 2.6100 8.9100 ;
      RECT 2.4760 7.8165 2.5020 8.9100 ;
      RECT 2.3680 7.8165 2.3940 8.9100 ;
      RECT 2.2600 7.8165 2.2860 8.9100 ;
      RECT 2.1520 7.8165 2.1780 8.9100 ;
      RECT 2.0440 7.8165 2.0700 8.9100 ;
      RECT 1.9360 7.8165 1.9620 8.9100 ;
      RECT 1.8280 7.8165 1.8540 8.9100 ;
      RECT 1.7200 7.8165 1.7460 8.9100 ;
      RECT 1.6120 7.8165 1.6380 8.9100 ;
      RECT 1.5040 7.8165 1.5300 8.9100 ;
      RECT 1.3960 7.8165 1.4220 8.9100 ;
      RECT 1.2880 7.8165 1.3140 8.9100 ;
      RECT 1.1800 7.8165 1.2060 8.9100 ;
      RECT 1.0720 7.8165 1.0980 8.9100 ;
      RECT 0.9640 7.8165 0.9900 8.9100 ;
      RECT 0.8560 7.8165 0.8820 8.9100 ;
      RECT 0.7480 7.8165 0.7740 8.9100 ;
      RECT 0.6400 7.8165 0.6660 8.9100 ;
      RECT 0.5320 7.8165 0.5580 8.9100 ;
      RECT 0.4240 7.8165 0.4500 8.9100 ;
      RECT 0.3160 7.8165 0.3420 8.9100 ;
      RECT 0.2080 7.8165 0.2340 8.9100 ;
      RECT 0.0050 7.8165 0.0900 8.9100 ;
      RECT 15.5530 8.8965 15.6810 9.9900 ;
      RECT 15.5390 9.5620 15.6810 9.8845 ;
      RECT 15.3190 9.2890 15.4530 9.9900 ;
      RECT 15.2960 9.6240 15.4530 9.8820 ;
      RECT 15.3190 8.8965 15.4170 9.9900 ;
      RECT 15.3190 9.0175 15.4310 9.2570 ;
      RECT 15.3190 8.8965 15.4530 8.9855 ;
      RECT 15.0940 9.3470 15.2280 9.9900 ;
      RECT 15.0940 8.8965 15.1920 9.9900 ;
      RECT 14.6770 8.8965 14.7600 9.9900 ;
      RECT 14.6770 8.9850 14.7740 9.9205 ;
      RECT 30.2680 8.8965 30.3530 9.9900 ;
      RECT 30.1240 8.8965 30.1500 9.9900 ;
      RECT 30.0160 8.8965 30.0420 9.9900 ;
      RECT 29.9080 8.8965 29.9340 9.9900 ;
      RECT 29.8000 8.8965 29.8260 9.9900 ;
      RECT 29.6920 8.8965 29.7180 9.9900 ;
      RECT 29.5840 8.8965 29.6100 9.9900 ;
      RECT 29.4760 8.8965 29.5020 9.9900 ;
      RECT 29.3680 8.8965 29.3940 9.9900 ;
      RECT 29.2600 8.8965 29.2860 9.9900 ;
      RECT 29.1520 8.8965 29.1780 9.9900 ;
      RECT 29.0440 8.8965 29.0700 9.9900 ;
      RECT 28.9360 8.8965 28.9620 9.9900 ;
      RECT 28.8280 8.8965 28.8540 9.9900 ;
      RECT 28.7200 8.8965 28.7460 9.9900 ;
      RECT 28.6120 8.8965 28.6380 9.9900 ;
      RECT 28.5040 8.8965 28.5300 9.9900 ;
      RECT 28.3960 8.8965 28.4220 9.9900 ;
      RECT 28.2880 8.8965 28.3140 9.9900 ;
      RECT 28.1800 8.8965 28.2060 9.9900 ;
      RECT 28.0720 8.8965 28.0980 9.9900 ;
      RECT 27.9640 8.8965 27.9900 9.9900 ;
      RECT 27.8560 8.8965 27.8820 9.9900 ;
      RECT 27.7480 8.8965 27.7740 9.9900 ;
      RECT 27.6400 8.8965 27.6660 9.9900 ;
      RECT 27.5320 8.8965 27.5580 9.9900 ;
      RECT 27.4240 8.8965 27.4500 9.9900 ;
      RECT 27.3160 8.8965 27.3420 9.9900 ;
      RECT 27.2080 8.8965 27.2340 9.9900 ;
      RECT 27.1000 8.8965 27.1260 9.9900 ;
      RECT 26.9920 8.8965 27.0180 9.9900 ;
      RECT 26.8840 8.8965 26.9100 9.9900 ;
      RECT 26.7760 8.8965 26.8020 9.9900 ;
      RECT 26.6680 8.8965 26.6940 9.9900 ;
      RECT 26.5600 8.8965 26.5860 9.9900 ;
      RECT 26.4520 8.8965 26.4780 9.9900 ;
      RECT 26.3440 8.8965 26.3700 9.9900 ;
      RECT 26.2360 8.8965 26.2620 9.9900 ;
      RECT 26.1280 8.8965 26.1540 9.9900 ;
      RECT 26.0200 8.8965 26.0460 9.9900 ;
      RECT 25.9120 8.8965 25.9380 9.9900 ;
      RECT 25.8040 8.8965 25.8300 9.9900 ;
      RECT 25.6960 8.8965 25.7220 9.9900 ;
      RECT 25.5880 8.8965 25.6140 9.9900 ;
      RECT 25.4800 8.8965 25.5060 9.9900 ;
      RECT 25.3720 8.8965 25.3980 9.9900 ;
      RECT 25.2640 8.8965 25.2900 9.9900 ;
      RECT 25.1560 8.8965 25.1820 9.9900 ;
      RECT 25.0480 8.8965 25.0740 9.9900 ;
      RECT 24.9400 8.8965 24.9660 9.9900 ;
      RECT 24.8320 8.8965 24.8580 9.9900 ;
      RECT 24.7240 8.8965 24.7500 9.9900 ;
      RECT 24.6160 8.8965 24.6420 9.9900 ;
      RECT 24.5080 8.8965 24.5340 9.9900 ;
      RECT 24.4000 8.8965 24.4260 9.9900 ;
      RECT 24.2920 8.8965 24.3180 9.9900 ;
      RECT 24.1840 8.8965 24.2100 9.9900 ;
      RECT 24.0760 8.8965 24.1020 9.9900 ;
      RECT 23.9680 8.8965 23.9940 9.9900 ;
      RECT 23.8600 8.8965 23.8860 9.9900 ;
      RECT 23.7520 8.8965 23.7780 9.9900 ;
      RECT 23.6440 8.8965 23.6700 9.9900 ;
      RECT 23.5360 8.8965 23.5620 9.9900 ;
      RECT 23.4280 8.8965 23.4540 9.9900 ;
      RECT 23.3200 8.8965 23.3460 9.9900 ;
      RECT 23.2120 8.8965 23.2380 9.9900 ;
      RECT 23.1040 8.8965 23.1300 9.9900 ;
      RECT 22.9960 8.8965 23.0220 9.9900 ;
      RECT 22.8880 8.8965 22.9140 9.9900 ;
      RECT 22.7800 8.8965 22.8060 9.9900 ;
      RECT 22.6720 8.8965 22.6980 9.9900 ;
      RECT 22.5640 8.8965 22.5900 9.9900 ;
      RECT 22.4560 8.8965 22.4820 9.9900 ;
      RECT 22.3480 8.8965 22.3740 9.9900 ;
      RECT 22.2400 8.8965 22.2660 9.9900 ;
      RECT 22.1320 8.8965 22.1580 9.9900 ;
      RECT 22.0240 8.8965 22.0500 9.9900 ;
      RECT 21.9160 8.8965 21.9420 9.9900 ;
      RECT 21.8080 8.8965 21.8340 9.9900 ;
      RECT 21.7000 8.8965 21.7260 9.9900 ;
      RECT 21.5920 8.8965 21.6180 9.9900 ;
      RECT 21.4840 8.8965 21.5100 9.9900 ;
      RECT 21.3760 8.8965 21.4020 9.9900 ;
      RECT 21.2680 8.8965 21.2940 9.9900 ;
      RECT 21.1600 8.8965 21.1860 9.9900 ;
      RECT 21.0520 8.8965 21.0780 9.9900 ;
      RECT 20.9440 8.8965 20.9700 9.9900 ;
      RECT 20.8360 8.8965 20.8620 9.9900 ;
      RECT 20.7280 8.8965 20.7540 9.9900 ;
      RECT 20.6200 8.8965 20.6460 9.9900 ;
      RECT 20.5120 8.8965 20.5380 9.9900 ;
      RECT 20.4040 8.8965 20.4300 9.9900 ;
      RECT 20.2960 8.8965 20.3220 9.9900 ;
      RECT 20.1880 8.8965 20.2140 9.9900 ;
      RECT 20.0800 8.8965 20.1060 9.9900 ;
      RECT 19.9720 8.8965 19.9980 9.9900 ;
      RECT 19.8640 8.8965 19.8900 9.9900 ;
      RECT 19.7560 8.8965 19.7820 9.9900 ;
      RECT 19.6480 8.8965 19.6740 9.9900 ;
      RECT 19.5400 8.8965 19.5660 9.9900 ;
      RECT 19.4320 8.8965 19.4580 9.9900 ;
      RECT 19.3240 8.8965 19.3500 9.9900 ;
      RECT 19.2160 8.8965 19.2420 9.9900 ;
      RECT 19.1080 8.8965 19.1340 9.9900 ;
      RECT 19.0000 8.8965 19.0260 9.9900 ;
      RECT 18.8920 8.8965 18.9180 9.9900 ;
      RECT 18.7840 8.8965 18.8100 9.9900 ;
      RECT 18.6760 8.8965 18.7020 9.9900 ;
      RECT 18.5680 8.8965 18.5940 9.9900 ;
      RECT 18.4600 8.8965 18.4860 9.9900 ;
      RECT 18.3520 8.8965 18.3780 9.9900 ;
      RECT 18.2440 8.8965 18.2700 9.9900 ;
      RECT 18.1360 8.8965 18.1620 9.9900 ;
      RECT 18.0280 8.8965 18.0540 9.9900 ;
      RECT 17.9200 8.8965 17.9460 9.9900 ;
      RECT 17.8120 8.8965 17.8380 9.9900 ;
      RECT 17.7040 8.8965 17.7300 9.9900 ;
      RECT 17.5960 8.8965 17.6220 9.9900 ;
      RECT 17.4880 8.8965 17.5140 9.9900 ;
      RECT 17.3800 8.8965 17.4060 9.9900 ;
      RECT 17.2720 8.8965 17.2980 9.9900 ;
      RECT 17.1640 8.8965 17.1900 9.9900 ;
      RECT 17.0560 8.8965 17.0820 9.9900 ;
      RECT 16.9480 8.8965 16.9740 9.9900 ;
      RECT 16.8400 8.8965 16.8660 9.9900 ;
      RECT 16.7320 8.8965 16.7580 9.9900 ;
      RECT 16.6240 8.8965 16.6500 9.9900 ;
      RECT 16.5160 8.8965 16.5420 9.9900 ;
      RECT 16.4080 8.8965 16.4340 9.9900 ;
      RECT 16.3000 8.8965 16.3260 9.9900 ;
      RECT 16.0870 8.8965 16.1640 9.9900 ;
      RECT 14.1940 8.8965 14.2710 9.9900 ;
      RECT 14.0320 8.8965 14.0580 9.9900 ;
      RECT 13.9240 8.8965 13.9500 9.9900 ;
      RECT 13.8160 8.8965 13.8420 9.9900 ;
      RECT 13.7080 8.8965 13.7340 9.9900 ;
      RECT 13.6000 8.8965 13.6260 9.9900 ;
      RECT 13.4920 8.8965 13.5180 9.9900 ;
      RECT 13.3840 8.8965 13.4100 9.9900 ;
      RECT 13.2760 8.8965 13.3020 9.9900 ;
      RECT 13.1680 8.8965 13.1940 9.9900 ;
      RECT 13.0600 8.8965 13.0860 9.9900 ;
      RECT 12.9520 8.8965 12.9780 9.9900 ;
      RECT 12.8440 8.8965 12.8700 9.9900 ;
      RECT 12.7360 8.8965 12.7620 9.9900 ;
      RECT 12.6280 8.8965 12.6540 9.9900 ;
      RECT 12.5200 8.8965 12.5460 9.9900 ;
      RECT 12.4120 8.8965 12.4380 9.9900 ;
      RECT 12.3040 8.8965 12.3300 9.9900 ;
      RECT 12.1960 8.8965 12.2220 9.9900 ;
      RECT 12.0880 8.8965 12.1140 9.9900 ;
      RECT 11.9800 8.8965 12.0060 9.9900 ;
      RECT 11.8720 8.8965 11.8980 9.9900 ;
      RECT 11.7640 8.8965 11.7900 9.9900 ;
      RECT 11.6560 8.8965 11.6820 9.9900 ;
      RECT 11.5480 8.8965 11.5740 9.9900 ;
      RECT 11.4400 8.8965 11.4660 9.9900 ;
      RECT 11.3320 8.8965 11.3580 9.9900 ;
      RECT 11.2240 8.8965 11.2500 9.9900 ;
      RECT 11.1160 8.8965 11.1420 9.9900 ;
      RECT 11.0080 8.8965 11.0340 9.9900 ;
      RECT 10.9000 8.8965 10.9260 9.9900 ;
      RECT 10.7920 8.8965 10.8180 9.9900 ;
      RECT 10.6840 8.8965 10.7100 9.9900 ;
      RECT 10.5760 8.8965 10.6020 9.9900 ;
      RECT 10.4680 8.8965 10.4940 9.9900 ;
      RECT 10.3600 8.8965 10.3860 9.9900 ;
      RECT 10.2520 8.8965 10.2780 9.9900 ;
      RECT 10.1440 8.8965 10.1700 9.9900 ;
      RECT 10.0360 8.8965 10.0620 9.9900 ;
      RECT 9.9280 8.8965 9.9540 9.9900 ;
      RECT 9.8200 8.8965 9.8460 9.9900 ;
      RECT 9.7120 8.8965 9.7380 9.9900 ;
      RECT 9.6040 8.8965 9.6300 9.9900 ;
      RECT 9.4960 8.8965 9.5220 9.9900 ;
      RECT 9.3880 8.8965 9.4140 9.9900 ;
      RECT 9.2800 8.8965 9.3060 9.9900 ;
      RECT 9.1720 8.8965 9.1980 9.9900 ;
      RECT 9.0640 8.8965 9.0900 9.9900 ;
      RECT 8.9560 8.8965 8.9820 9.9900 ;
      RECT 8.8480 8.8965 8.8740 9.9900 ;
      RECT 8.7400 8.8965 8.7660 9.9900 ;
      RECT 8.6320 8.8965 8.6580 9.9900 ;
      RECT 8.5240 8.8965 8.5500 9.9900 ;
      RECT 8.4160 8.8965 8.4420 9.9900 ;
      RECT 8.3080 8.8965 8.3340 9.9900 ;
      RECT 8.2000 8.8965 8.2260 9.9900 ;
      RECT 8.0920 8.8965 8.1180 9.9900 ;
      RECT 7.9840 8.8965 8.0100 9.9900 ;
      RECT 7.8760 8.8965 7.9020 9.9900 ;
      RECT 7.7680 8.8965 7.7940 9.9900 ;
      RECT 7.6600 8.8965 7.6860 9.9900 ;
      RECT 7.5520 8.8965 7.5780 9.9900 ;
      RECT 7.4440 8.8965 7.4700 9.9900 ;
      RECT 7.3360 8.8965 7.3620 9.9900 ;
      RECT 7.2280 8.8965 7.2540 9.9900 ;
      RECT 7.1200 8.8965 7.1460 9.9900 ;
      RECT 7.0120 8.8965 7.0380 9.9900 ;
      RECT 6.9040 8.8965 6.9300 9.9900 ;
      RECT 6.7960 8.8965 6.8220 9.9900 ;
      RECT 6.6880 8.8965 6.7140 9.9900 ;
      RECT 6.5800 8.8965 6.6060 9.9900 ;
      RECT 6.4720 8.8965 6.4980 9.9900 ;
      RECT 6.3640 8.8965 6.3900 9.9900 ;
      RECT 6.2560 8.8965 6.2820 9.9900 ;
      RECT 6.1480 8.8965 6.1740 9.9900 ;
      RECT 6.0400 8.8965 6.0660 9.9900 ;
      RECT 5.9320 8.8965 5.9580 9.9900 ;
      RECT 5.8240 8.8965 5.8500 9.9900 ;
      RECT 5.7160 8.8965 5.7420 9.9900 ;
      RECT 5.6080 8.8965 5.6340 9.9900 ;
      RECT 5.5000 8.8965 5.5260 9.9900 ;
      RECT 5.3920 8.8965 5.4180 9.9900 ;
      RECT 5.2840 8.8965 5.3100 9.9900 ;
      RECT 5.1760 8.8965 5.2020 9.9900 ;
      RECT 5.0680 8.8965 5.0940 9.9900 ;
      RECT 4.9600 8.8965 4.9860 9.9900 ;
      RECT 4.8520 8.8965 4.8780 9.9900 ;
      RECT 4.7440 8.8965 4.7700 9.9900 ;
      RECT 4.6360 8.8965 4.6620 9.9900 ;
      RECT 4.5280 8.8965 4.5540 9.9900 ;
      RECT 4.4200 8.8965 4.4460 9.9900 ;
      RECT 4.3120 8.8965 4.3380 9.9900 ;
      RECT 4.2040 8.8965 4.2300 9.9900 ;
      RECT 4.0960 8.8965 4.1220 9.9900 ;
      RECT 3.9880 8.8965 4.0140 9.9900 ;
      RECT 3.8800 8.8965 3.9060 9.9900 ;
      RECT 3.7720 8.8965 3.7980 9.9900 ;
      RECT 3.6640 8.8965 3.6900 9.9900 ;
      RECT 3.5560 8.8965 3.5820 9.9900 ;
      RECT 3.4480 8.8965 3.4740 9.9900 ;
      RECT 3.3400 8.8965 3.3660 9.9900 ;
      RECT 3.2320 8.8965 3.2580 9.9900 ;
      RECT 3.1240 8.8965 3.1500 9.9900 ;
      RECT 3.0160 8.8965 3.0420 9.9900 ;
      RECT 2.9080 8.8965 2.9340 9.9900 ;
      RECT 2.8000 8.8965 2.8260 9.9900 ;
      RECT 2.6920 8.8965 2.7180 9.9900 ;
      RECT 2.5840 8.8965 2.6100 9.9900 ;
      RECT 2.4760 8.8965 2.5020 9.9900 ;
      RECT 2.3680 8.8965 2.3940 9.9900 ;
      RECT 2.2600 8.8965 2.2860 9.9900 ;
      RECT 2.1520 8.8965 2.1780 9.9900 ;
      RECT 2.0440 8.8965 2.0700 9.9900 ;
      RECT 1.9360 8.8965 1.9620 9.9900 ;
      RECT 1.8280 8.8965 1.8540 9.9900 ;
      RECT 1.7200 8.8965 1.7460 9.9900 ;
      RECT 1.6120 8.8965 1.6380 9.9900 ;
      RECT 1.5040 8.8965 1.5300 9.9900 ;
      RECT 1.3960 8.8965 1.4220 9.9900 ;
      RECT 1.2880 8.8965 1.3140 9.9900 ;
      RECT 1.1800 8.8965 1.2060 9.9900 ;
      RECT 1.0720 8.8965 1.0980 9.9900 ;
      RECT 0.9640 8.8965 0.9900 9.9900 ;
      RECT 0.8560 8.8965 0.8820 9.9900 ;
      RECT 0.7480 8.8965 0.7740 9.9900 ;
      RECT 0.6400 8.8965 0.6660 9.9900 ;
      RECT 0.5320 8.8965 0.5580 9.9900 ;
      RECT 0.4240 8.8965 0.4500 9.9900 ;
      RECT 0.3160 8.8965 0.3420 9.9900 ;
      RECT 0.2080 8.8965 0.2340 9.9900 ;
      RECT 0.0050 8.8965 0.0900 9.9900 ;
      RECT 15.5530 9.9765 15.6810 11.0700 ;
      RECT 15.5390 10.6420 15.6810 10.9645 ;
      RECT 15.3190 10.3690 15.4530 11.0700 ;
      RECT 15.2960 10.7040 15.4530 10.9620 ;
      RECT 15.3190 9.9765 15.4170 11.0700 ;
      RECT 15.3190 10.0975 15.4310 10.3370 ;
      RECT 15.3190 9.9765 15.4530 10.0655 ;
      RECT 15.0940 10.4270 15.2280 11.0700 ;
      RECT 15.0940 9.9765 15.1920 11.0700 ;
      RECT 14.6770 9.9765 14.7600 11.0700 ;
      RECT 14.6770 10.0650 14.7740 11.0005 ;
      RECT 30.2680 9.9765 30.3530 11.0700 ;
      RECT 30.1240 9.9765 30.1500 11.0700 ;
      RECT 30.0160 9.9765 30.0420 11.0700 ;
      RECT 29.9080 9.9765 29.9340 11.0700 ;
      RECT 29.8000 9.9765 29.8260 11.0700 ;
      RECT 29.6920 9.9765 29.7180 11.0700 ;
      RECT 29.5840 9.9765 29.6100 11.0700 ;
      RECT 29.4760 9.9765 29.5020 11.0700 ;
      RECT 29.3680 9.9765 29.3940 11.0700 ;
      RECT 29.2600 9.9765 29.2860 11.0700 ;
      RECT 29.1520 9.9765 29.1780 11.0700 ;
      RECT 29.0440 9.9765 29.0700 11.0700 ;
      RECT 28.9360 9.9765 28.9620 11.0700 ;
      RECT 28.8280 9.9765 28.8540 11.0700 ;
      RECT 28.7200 9.9765 28.7460 11.0700 ;
      RECT 28.6120 9.9765 28.6380 11.0700 ;
      RECT 28.5040 9.9765 28.5300 11.0700 ;
      RECT 28.3960 9.9765 28.4220 11.0700 ;
      RECT 28.2880 9.9765 28.3140 11.0700 ;
      RECT 28.1800 9.9765 28.2060 11.0700 ;
      RECT 28.0720 9.9765 28.0980 11.0700 ;
      RECT 27.9640 9.9765 27.9900 11.0700 ;
      RECT 27.8560 9.9765 27.8820 11.0700 ;
      RECT 27.7480 9.9765 27.7740 11.0700 ;
      RECT 27.6400 9.9765 27.6660 11.0700 ;
      RECT 27.5320 9.9765 27.5580 11.0700 ;
      RECT 27.4240 9.9765 27.4500 11.0700 ;
      RECT 27.3160 9.9765 27.3420 11.0700 ;
      RECT 27.2080 9.9765 27.2340 11.0700 ;
      RECT 27.1000 9.9765 27.1260 11.0700 ;
      RECT 26.9920 9.9765 27.0180 11.0700 ;
      RECT 26.8840 9.9765 26.9100 11.0700 ;
      RECT 26.7760 9.9765 26.8020 11.0700 ;
      RECT 26.6680 9.9765 26.6940 11.0700 ;
      RECT 26.5600 9.9765 26.5860 11.0700 ;
      RECT 26.4520 9.9765 26.4780 11.0700 ;
      RECT 26.3440 9.9765 26.3700 11.0700 ;
      RECT 26.2360 9.9765 26.2620 11.0700 ;
      RECT 26.1280 9.9765 26.1540 11.0700 ;
      RECT 26.0200 9.9765 26.0460 11.0700 ;
      RECT 25.9120 9.9765 25.9380 11.0700 ;
      RECT 25.8040 9.9765 25.8300 11.0700 ;
      RECT 25.6960 9.9765 25.7220 11.0700 ;
      RECT 25.5880 9.9765 25.6140 11.0700 ;
      RECT 25.4800 9.9765 25.5060 11.0700 ;
      RECT 25.3720 9.9765 25.3980 11.0700 ;
      RECT 25.2640 9.9765 25.2900 11.0700 ;
      RECT 25.1560 9.9765 25.1820 11.0700 ;
      RECT 25.0480 9.9765 25.0740 11.0700 ;
      RECT 24.9400 9.9765 24.9660 11.0700 ;
      RECT 24.8320 9.9765 24.8580 11.0700 ;
      RECT 24.7240 9.9765 24.7500 11.0700 ;
      RECT 24.6160 9.9765 24.6420 11.0700 ;
      RECT 24.5080 9.9765 24.5340 11.0700 ;
      RECT 24.4000 9.9765 24.4260 11.0700 ;
      RECT 24.2920 9.9765 24.3180 11.0700 ;
      RECT 24.1840 9.9765 24.2100 11.0700 ;
      RECT 24.0760 9.9765 24.1020 11.0700 ;
      RECT 23.9680 9.9765 23.9940 11.0700 ;
      RECT 23.8600 9.9765 23.8860 11.0700 ;
      RECT 23.7520 9.9765 23.7780 11.0700 ;
      RECT 23.6440 9.9765 23.6700 11.0700 ;
      RECT 23.5360 9.9765 23.5620 11.0700 ;
      RECT 23.4280 9.9765 23.4540 11.0700 ;
      RECT 23.3200 9.9765 23.3460 11.0700 ;
      RECT 23.2120 9.9765 23.2380 11.0700 ;
      RECT 23.1040 9.9765 23.1300 11.0700 ;
      RECT 22.9960 9.9765 23.0220 11.0700 ;
      RECT 22.8880 9.9765 22.9140 11.0700 ;
      RECT 22.7800 9.9765 22.8060 11.0700 ;
      RECT 22.6720 9.9765 22.6980 11.0700 ;
      RECT 22.5640 9.9765 22.5900 11.0700 ;
      RECT 22.4560 9.9765 22.4820 11.0700 ;
      RECT 22.3480 9.9765 22.3740 11.0700 ;
      RECT 22.2400 9.9765 22.2660 11.0700 ;
      RECT 22.1320 9.9765 22.1580 11.0700 ;
      RECT 22.0240 9.9765 22.0500 11.0700 ;
      RECT 21.9160 9.9765 21.9420 11.0700 ;
      RECT 21.8080 9.9765 21.8340 11.0700 ;
      RECT 21.7000 9.9765 21.7260 11.0700 ;
      RECT 21.5920 9.9765 21.6180 11.0700 ;
      RECT 21.4840 9.9765 21.5100 11.0700 ;
      RECT 21.3760 9.9765 21.4020 11.0700 ;
      RECT 21.2680 9.9765 21.2940 11.0700 ;
      RECT 21.1600 9.9765 21.1860 11.0700 ;
      RECT 21.0520 9.9765 21.0780 11.0700 ;
      RECT 20.9440 9.9765 20.9700 11.0700 ;
      RECT 20.8360 9.9765 20.8620 11.0700 ;
      RECT 20.7280 9.9765 20.7540 11.0700 ;
      RECT 20.6200 9.9765 20.6460 11.0700 ;
      RECT 20.5120 9.9765 20.5380 11.0700 ;
      RECT 20.4040 9.9765 20.4300 11.0700 ;
      RECT 20.2960 9.9765 20.3220 11.0700 ;
      RECT 20.1880 9.9765 20.2140 11.0700 ;
      RECT 20.0800 9.9765 20.1060 11.0700 ;
      RECT 19.9720 9.9765 19.9980 11.0700 ;
      RECT 19.8640 9.9765 19.8900 11.0700 ;
      RECT 19.7560 9.9765 19.7820 11.0700 ;
      RECT 19.6480 9.9765 19.6740 11.0700 ;
      RECT 19.5400 9.9765 19.5660 11.0700 ;
      RECT 19.4320 9.9765 19.4580 11.0700 ;
      RECT 19.3240 9.9765 19.3500 11.0700 ;
      RECT 19.2160 9.9765 19.2420 11.0700 ;
      RECT 19.1080 9.9765 19.1340 11.0700 ;
      RECT 19.0000 9.9765 19.0260 11.0700 ;
      RECT 18.8920 9.9765 18.9180 11.0700 ;
      RECT 18.7840 9.9765 18.8100 11.0700 ;
      RECT 18.6760 9.9765 18.7020 11.0700 ;
      RECT 18.5680 9.9765 18.5940 11.0700 ;
      RECT 18.4600 9.9765 18.4860 11.0700 ;
      RECT 18.3520 9.9765 18.3780 11.0700 ;
      RECT 18.2440 9.9765 18.2700 11.0700 ;
      RECT 18.1360 9.9765 18.1620 11.0700 ;
      RECT 18.0280 9.9765 18.0540 11.0700 ;
      RECT 17.9200 9.9765 17.9460 11.0700 ;
      RECT 17.8120 9.9765 17.8380 11.0700 ;
      RECT 17.7040 9.9765 17.7300 11.0700 ;
      RECT 17.5960 9.9765 17.6220 11.0700 ;
      RECT 17.4880 9.9765 17.5140 11.0700 ;
      RECT 17.3800 9.9765 17.4060 11.0700 ;
      RECT 17.2720 9.9765 17.2980 11.0700 ;
      RECT 17.1640 9.9765 17.1900 11.0700 ;
      RECT 17.0560 9.9765 17.0820 11.0700 ;
      RECT 16.9480 9.9765 16.9740 11.0700 ;
      RECT 16.8400 9.9765 16.8660 11.0700 ;
      RECT 16.7320 9.9765 16.7580 11.0700 ;
      RECT 16.6240 9.9765 16.6500 11.0700 ;
      RECT 16.5160 9.9765 16.5420 11.0700 ;
      RECT 16.4080 9.9765 16.4340 11.0700 ;
      RECT 16.3000 9.9765 16.3260 11.0700 ;
      RECT 16.0870 9.9765 16.1640 11.0700 ;
      RECT 14.1940 9.9765 14.2710 11.0700 ;
      RECT 14.0320 9.9765 14.0580 11.0700 ;
      RECT 13.9240 9.9765 13.9500 11.0700 ;
      RECT 13.8160 9.9765 13.8420 11.0700 ;
      RECT 13.7080 9.9765 13.7340 11.0700 ;
      RECT 13.6000 9.9765 13.6260 11.0700 ;
      RECT 13.4920 9.9765 13.5180 11.0700 ;
      RECT 13.3840 9.9765 13.4100 11.0700 ;
      RECT 13.2760 9.9765 13.3020 11.0700 ;
      RECT 13.1680 9.9765 13.1940 11.0700 ;
      RECT 13.0600 9.9765 13.0860 11.0700 ;
      RECT 12.9520 9.9765 12.9780 11.0700 ;
      RECT 12.8440 9.9765 12.8700 11.0700 ;
      RECT 12.7360 9.9765 12.7620 11.0700 ;
      RECT 12.6280 9.9765 12.6540 11.0700 ;
      RECT 12.5200 9.9765 12.5460 11.0700 ;
      RECT 12.4120 9.9765 12.4380 11.0700 ;
      RECT 12.3040 9.9765 12.3300 11.0700 ;
      RECT 12.1960 9.9765 12.2220 11.0700 ;
      RECT 12.0880 9.9765 12.1140 11.0700 ;
      RECT 11.9800 9.9765 12.0060 11.0700 ;
      RECT 11.8720 9.9765 11.8980 11.0700 ;
      RECT 11.7640 9.9765 11.7900 11.0700 ;
      RECT 11.6560 9.9765 11.6820 11.0700 ;
      RECT 11.5480 9.9765 11.5740 11.0700 ;
      RECT 11.4400 9.9765 11.4660 11.0700 ;
      RECT 11.3320 9.9765 11.3580 11.0700 ;
      RECT 11.2240 9.9765 11.2500 11.0700 ;
      RECT 11.1160 9.9765 11.1420 11.0700 ;
      RECT 11.0080 9.9765 11.0340 11.0700 ;
      RECT 10.9000 9.9765 10.9260 11.0700 ;
      RECT 10.7920 9.9765 10.8180 11.0700 ;
      RECT 10.6840 9.9765 10.7100 11.0700 ;
      RECT 10.5760 9.9765 10.6020 11.0700 ;
      RECT 10.4680 9.9765 10.4940 11.0700 ;
      RECT 10.3600 9.9765 10.3860 11.0700 ;
      RECT 10.2520 9.9765 10.2780 11.0700 ;
      RECT 10.1440 9.9765 10.1700 11.0700 ;
      RECT 10.0360 9.9765 10.0620 11.0700 ;
      RECT 9.9280 9.9765 9.9540 11.0700 ;
      RECT 9.8200 9.9765 9.8460 11.0700 ;
      RECT 9.7120 9.9765 9.7380 11.0700 ;
      RECT 9.6040 9.9765 9.6300 11.0700 ;
      RECT 9.4960 9.9765 9.5220 11.0700 ;
      RECT 9.3880 9.9765 9.4140 11.0700 ;
      RECT 9.2800 9.9765 9.3060 11.0700 ;
      RECT 9.1720 9.9765 9.1980 11.0700 ;
      RECT 9.0640 9.9765 9.0900 11.0700 ;
      RECT 8.9560 9.9765 8.9820 11.0700 ;
      RECT 8.8480 9.9765 8.8740 11.0700 ;
      RECT 8.7400 9.9765 8.7660 11.0700 ;
      RECT 8.6320 9.9765 8.6580 11.0700 ;
      RECT 8.5240 9.9765 8.5500 11.0700 ;
      RECT 8.4160 9.9765 8.4420 11.0700 ;
      RECT 8.3080 9.9765 8.3340 11.0700 ;
      RECT 8.2000 9.9765 8.2260 11.0700 ;
      RECT 8.0920 9.9765 8.1180 11.0700 ;
      RECT 7.9840 9.9765 8.0100 11.0700 ;
      RECT 7.8760 9.9765 7.9020 11.0700 ;
      RECT 7.7680 9.9765 7.7940 11.0700 ;
      RECT 7.6600 9.9765 7.6860 11.0700 ;
      RECT 7.5520 9.9765 7.5780 11.0700 ;
      RECT 7.4440 9.9765 7.4700 11.0700 ;
      RECT 7.3360 9.9765 7.3620 11.0700 ;
      RECT 7.2280 9.9765 7.2540 11.0700 ;
      RECT 7.1200 9.9765 7.1460 11.0700 ;
      RECT 7.0120 9.9765 7.0380 11.0700 ;
      RECT 6.9040 9.9765 6.9300 11.0700 ;
      RECT 6.7960 9.9765 6.8220 11.0700 ;
      RECT 6.6880 9.9765 6.7140 11.0700 ;
      RECT 6.5800 9.9765 6.6060 11.0700 ;
      RECT 6.4720 9.9765 6.4980 11.0700 ;
      RECT 6.3640 9.9765 6.3900 11.0700 ;
      RECT 6.2560 9.9765 6.2820 11.0700 ;
      RECT 6.1480 9.9765 6.1740 11.0700 ;
      RECT 6.0400 9.9765 6.0660 11.0700 ;
      RECT 5.9320 9.9765 5.9580 11.0700 ;
      RECT 5.8240 9.9765 5.8500 11.0700 ;
      RECT 5.7160 9.9765 5.7420 11.0700 ;
      RECT 5.6080 9.9765 5.6340 11.0700 ;
      RECT 5.5000 9.9765 5.5260 11.0700 ;
      RECT 5.3920 9.9765 5.4180 11.0700 ;
      RECT 5.2840 9.9765 5.3100 11.0700 ;
      RECT 5.1760 9.9765 5.2020 11.0700 ;
      RECT 5.0680 9.9765 5.0940 11.0700 ;
      RECT 4.9600 9.9765 4.9860 11.0700 ;
      RECT 4.8520 9.9765 4.8780 11.0700 ;
      RECT 4.7440 9.9765 4.7700 11.0700 ;
      RECT 4.6360 9.9765 4.6620 11.0700 ;
      RECT 4.5280 9.9765 4.5540 11.0700 ;
      RECT 4.4200 9.9765 4.4460 11.0700 ;
      RECT 4.3120 9.9765 4.3380 11.0700 ;
      RECT 4.2040 9.9765 4.2300 11.0700 ;
      RECT 4.0960 9.9765 4.1220 11.0700 ;
      RECT 3.9880 9.9765 4.0140 11.0700 ;
      RECT 3.8800 9.9765 3.9060 11.0700 ;
      RECT 3.7720 9.9765 3.7980 11.0700 ;
      RECT 3.6640 9.9765 3.6900 11.0700 ;
      RECT 3.5560 9.9765 3.5820 11.0700 ;
      RECT 3.4480 9.9765 3.4740 11.0700 ;
      RECT 3.3400 9.9765 3.3660 11.0700 ;
      RECT 3.2320 9.9765 3.2580 11.0700 ;
      RECT 3.1240 9.9765 3.1500 11.0700 ;
      RECT 3.0160 9.9765 3.0420 11.0700 ;
      RECT 2.9080 9.9765 2.9340 11.0700 ;
      RECT 2.8000 9.9765 2.8260 11.0700 ;
      RECT 2.6920 9.9765 2.7180 11.0700 ;
      RECT 2.5840 9.9765 2.6100 11.0700 ;
      RECT 2.4760 9.9765 2.5020 11.0700 ;
      RECT 2.3680 9.9765 2.3940 11.0700 ;
      RECT 2.2600 9.9765 2.2860 11.0700 ;
      RECT 2.1520 9.9765 2.1780 11.0700 ;
      RECT 2.0440 9.9765 2.0700 11.0700 ;
      RECT 1.9360 9.9765 1.9620 11.0700 ;
      RECT 1.8280 9.9765 1.8540 11.0700 ;
      RECT 1.7200 9.9765 1.7460 11.0700 ;
      RECT 1.6120 9.9765 1.6380 11.0700 ;
      RECT 1.5040 9.9765 1.5300 11.0700 ;
      RECT 1.3960 9.9765 1.4220 11.0700 ;
      RECT 1.2880 9.9765 1.3140 11.0700 ;
      RECT 1.1800 9.9765 1.2060 11.0700 ;
      RECT 1.0720 9.9765 1.0980 11.0700 ;
      RECT 0.9640 9.9765 0.9900 11.0700 ;
      RECT 0.8560 9.9765 0.8820 11.0700 ;
      RECT 0.7480 9.9765 0.7740 11.0700 ;
      RECT 0.6400 9.9765 0.6660 11.0700 ;
      RECT 0.5320 9.9765 0.5580 11.0700 ;
      RECT 0.4240 9.9765 0.4500 11.0700 ;
      RECT 0.3160 9.9765 0.3420 11.0700 ;
      RECT 0.2080 9.9765 0.2340 11.0700 ;
      RECT 0.0050 9.9765 0.0900 11.0700 ;
      RECT 15.5530 11.0565 15.6810 12.1500 ;
      RECT 15.5390 11.7220 15.6810 12.0445 ;
      RECT 15.3190 11.4490 15.4530 12.1500 ;
      RECT 15.2960 11.7840 15.4530 12.0420 ;
      RECT 15.3190 11.0565 15.4170 12.1500 ;
      RECT 15.3190 11.1775 15.4310 11.4170 ;
      RECT 15.3190 11.0565 15.4530 11.1455 ;
      RECT 15.0940 11.5070 15.2280 12.1500 ;
      RECT 15.0940 11.0565 15.1920 12.1500 ;
      RECT 14.6770 11.0565 14.7600 12.1500 ;
      RECT 14.6770 11.1450 14.7740 12.0805 ;
      RECT 30.2680 11.0565 30.3530 12.1500 ;
      RECT 30.1240 11.0565 30.1500 12.1500 ;
      RECT 30.0160 11.0565 30.0420 12.1500 ;
      RECT 29.9080 11.0565 29.9340 12.1500 ;
      RECT 29.8000 11.0565 29.8260 12.1500 ;
      RECT 29.6920 11.0565 29.7180 12.1500 ;
      RECT 29.5840 11.0565 29.6100 12.1500 ;
      RECT 29.4760 11.0565 29.5020 12.1500 ;
      RECT 29.3680 11.0565 29.3940 12.1500 ;
      RECT 29.2600 11.0565 29.2860 12.1500 ;
      RECT 29.1520 11.0565 29.1780 12.1500 ;
      RECT 29.0440 11.0565 29.0700 12.1500 ;
      RECT 28.9360 11.0565 28.9620 12.1500 ;
      RECT 28.8280 11.0565 28.8540 12.1500 ;
      RECT 28.7200 11.0565 28.7460 12.1500 ;
      RECT 28.6120 11.0565 28.6380 12.1500 ;
      RECT 28.5040 11.0565 28.5300 12.1500 ;
      RECT 28.3960 11.0565 28.4220 12.1500 ;
      RECT 28.2880 11.0565 28.3140 12.1500 ;
      RECT 28.1800 11.0565 28.2060 12.1500 ;
      RECT 28.0720 11.0565 28.0980 12.1500 ;
      RECT 27.9640 11.0565 27.9900 12.1500 ;
      RECT 27.8560 11.0565 27.8820 12.1500 ;
      RECT 27.7480 11.0565 27.7740 12.1500 ;
      RECT 27.6400 11.0565 27.6660 12.1500 ;
      RECT 27.5320 11.0565 27.5580 12.1500 ;
      RECT 27.4240 11.0565 27.4500 12.1500 ;
      RECT 27.3160 11.0565 27.3420 12.1500 ;
      RECT 27.2080 11.0565 27.2340 12.1500 ;
      RECT 27.1000 11.0565 27.1260 12.1500 ;
      RECT 26.9920 11.0565 27.0180 12.1500 ;
      RECT 26.8840 11.0565 26.9100 12.1500 ;
      RECT 26.7760 11.0565 26.8020 12.1500 ;
      RECT 26.6680 11.0565 26.6940 12.1500 ;
      RECT 26.5600 11.0565 26.5860 12.1500 ;
      RECT 26.4520 11.0565 26.4780 12.1500 ;
      RECT 26.3440 11.0565 26.3700 12.1500 ;
      RECT 26.2360 11.0565 26.2620 12.1500 ;
      RECT 26.1280 11.0565 26.1540 12.1500 ;
      RECT 26.0200 11.0565 26.0460 12.1500 ;
      RECT 25.9120 11.0565 25.9380 12.1500 ;
      RECT 25.8040 11.0565 25.8300 12.1500 ;
      RECT 25.6960 11.0565 25.7220 12.1500 ;
      RECT 25.5880 11.0565 25.6140 12.1500 ;
      RECT 25.4800 11.0565 25.5060 12.1500 ;
      RECT 25.3720 11.0565 25.3980 12.1500 ;
      RECT 25.2640 11.0565 25.2900 12.1500 ;
      RECT 25.1560 11.0565 25.1820 12.1500 ;
      RECT 25.0480 11.0565 25.0740 12.1500 ;
      RECT 24.9400 11.0565 24.9660 12.1500 ;
      RECT 24.8320 11.0565 24.8580 12.1500 ;
      RECT 24.7240 11.0565 24.7500 12.1500 ;
      RECT 24.6160 11.0565 24.6420 12.1500 ;
      RECT 24.5080 11.0565 24.5340 12.1500 ;
      RECT 24.4000 11.0565 24.4260 12.1500 ;
      RECT 24.2920 11.0565 24.3180 12.1500 ;
      RECT 24.1840 11.0565 24.2100 12.1500 ;
      RECT 24.0760 11.0565 24.1020 12.1500 ;
      RECT 23.9680 11.0565 23.9940 12.1500 ;
      RECT 23.8600 11.0565 23.8860 12.1500 ;
      RECT 23.7520 11.0565 23.7780 12.1500 ;
      RECT 23.6440 11.0565 23.6700 12.1500 ;
      RECT 23.5360 11.0565 23.5620 12.1500 ;
      RECT 23.4280 11.0565 23.4540 12.1500 ;
      RECT 23.3200 11.0565 23.3460 12.1500 ;
      RECT 23.2120 11.0565 23.2380 12.1500 ;
      RECT 23.1040 11.0565 23.1300 12.1500 ;
      RECT 22.9960 11.0565 23.0220 12.1500 ;
      RECT 22.8880 11.0565 22.9140 12.1500 ;
      RECT 22.7800 11.0565 22.8060 12.1500 ;
      RECT 22.6720 11.0565 22.6980 12.1500 ;
      RECT 22.5640 11.0565 22.5900 12.1500 ;
      RECT 22.4560 11.0565 22.4820 12.1500 ;
      RECT 22.3480 11.0565 22.3740 12.1500 ;
      RECT 22.2400 11.0565 22.2660 12.1500 ;
      RECT 22.1320 11.0565 22.1580 12.1500 ;
      RECT 22.0240 11.0565 22.0500 12.1500 ;
      RECT 21.9160 11.0565 21.9420 12.1500 ;
      RECT 21.8080 11.0565 21.8340 12.1500 ;
      RECT 21.7000 11.0565 21.7260 12.1500 ;
      RECT 21.5920 11.0565 21.6180 12.1500 ;
      RECT 21.4840 11.0565 21.5100 12.1500 ;
      RECT 21.3760 11.0565 21.4020 12.1500 ;
      RECT 21.2680 11.0565 21.2940 12.1500 ;
      RECT 21.1600 11.0565 21.1860 12.1500 ;
      RECT 21.0520 11.0565 21.0780 12.1500 ;
      RECT 20.9440 11.0565 20.9700 12.1500 ;
      RECT 20.8360 11.0565 20.8620 12.1500 ;
      RECT 20.7280 11.0565 20.7540 12.1500 ;
      RECT 20.6200 11.0565 20.6460 12.1500 ;
      RECT 20.5120 11.0565 20.5380 12.1500 ;
      RECT 20.4040 11.0565 20.4300 12.1500 ;
      RECT 20.2960 11.0565 20.3220 12.1500 ;
      RECT 20.1880 11.0565 20.2140 12.1500 ;
      RECT 20.0800 11.0565 20.1060 12.1500 ;
      RECT 19.9720 11.0565 19.9980 12.1500 ;
      RECT 19.8640 11.0565 19.8900 12.1500 ;
      RECT 19.7560 11.0565 19.7820 12.1500 ;
      RECT 19.6480 11.0565 19.6740 12.1500 ;
      RECT 19.5400 11.0565 19.5660 12.1500 ;
      RECT 19.4320 11.0565 19.4580 12.1500 ;
      RECT 19.3240 11.0565 19.3500 12.1500 ;
      RECT 19.2160 11.0565 19.2420 12.1500 ;
      RECT 19.1080 11.0565 19.1340 12.1500 ;
      RECT 19.0000 11.0565 19.0260 12.1500 ;
      RECT 18.8920 11.0565 18.9180 12.1500 ;
      RECT 18.7840 11.0565 18.8100 12.1500 ;
      RECT 18.6760 11.0565 18.7020 12.1500 ;
      RECT 18.5680 11.0565 18.5940 12.1500 ;
      RECT 18.4600 11.0565 18.4860 12.1500 ;
      RECT 18.3520 11.0565 18.3780 12.1500 ;
      RECT 18.2440 11.0565 18.2700 12.1500 ;
      RECT 18.1360 11.0565 18.1620 12.1500 ;
      RECT 18.0280 11.0565 18.0540 12.1500 ;
      RECT 17.9200 11.0565 17.9460 12.1500 ;
      RECT 17.8120 11.0565 17.8380 12.1500 ;
      RECT 17.7040 11.0565 17.7300 12.1500 ;
      RECT 17.5960 11.0565 17.6220 12.1500 ;
      RECT 17.4880 11.0565 17.5140 12.1500 ;
      RECT 17.3800 11.0565 17.4060 12.1500 ;
      RECT 17.2720 11.0565 17.2980 12.1500 ;
      RECT 17.1640 11.0565 17.1900 12.1500 ;
      RECT 17.0560 11.0565 17.0820 12.1500 ;
      RECT 16.9480 11.0565 16.9740 12.1500 ;
      RECT 16.8400 11.0565 16.8660 12.1500 ;
      RECT 16.7320 11.0565 16.7580 12.1500 ;
      RECT 16.6240 11.0565 16.6500 12.1500 ;
      RECT 16.5160 11.0565 16.5420 12.1500 ;
      RECT 16.4080 11.0565 16.4340 12.1500 ;
      RECT 16.3000 11.0565 16.3260 12.1500 ;
      RECT 16.0870 11.0565 16.1640 12.1500 ;
      RECT 14.1940 11.0565 14.2710 12.1500 ;
      RECT 14.0320 11.0565 14.0580 12.1500 ;
      RECT 13.9240 11.0565 13.9500 12.1500 ;
      RECT 13.8160 11.0565 13.8420 12.1500 ;
      RECT 13.7080 11.0565 13.7340 12.1500 ;
      RECT 13.6000 11.0565 13.6260 12.1500 ;
      RECT 13.4920 11.0565 13.5180 12.1500 ;
      RECT 13.3840 11.0565 13.4100 12.1500 ;
      RECT 13.2760 11.0565 13.3020 12.1500 ;
      RECT 13.1680 11.0565 13.1940 12.1500 ;
      RECT 13.0600 11.0565 13.0860 12.1500 ;
      RECT 12.9520 11.0565 12.9780 12.1500 ;
      RECT 12.8440 11.0565 12.8700 12.1500 ;
      RECT 12.7360 11.0565 12.7620 12.1500 ;
      RECT 12.6280 11.0565 12.6540 12.1500 ;
      RECT 12.5200 11.0565 12.5460 12.1500 ;
      RECT 12.4120 11.0565 12.4380 12.1500 ;
      RECT 12.3040 11.0565 12.3300 12.1500 ;
      RECT 12.1960 11.0565 12.2220 12.1500 ;
      RECT 12.0880 11.0565 12.1140 12.1500 ;
      RECT 11.9800 11.0565 12.0060 12.1500 ;
      RECT 11.8720 11.0565 11.8980 12.1500 ;
      RECT 11.7640 11.0565 11.7900 12.1500 ;
      RECT 11.6560 11.0565 11.6820 12.1500 ;
      RECT 11.5480 11.0565 11.5740 12.1500 ;
      RECT 11.4400 11.0565 11.4660 12.1500 ;
      RECT 11.3320 11.0565 11.3580 12.1500 ;
      RECT 11.2240 11.0565 11.2500 12.1500 ;
      RECT 11.1160 11.0565 11.1420 12.1500 ;
      RECT 11.0080 11.0565 11.0340 12.1500 ;
      RECT 10.9000 11.0565 10.9260 12.1500 ;
      RECT 10.7920 11.0565 10.8180 12.1500 ;
      RECT 10.6840 11.0565 10.7100 12.1500 ;
      RECT 10.5760 11.0565 10.6020 12.1500 ;
      RECT 10.4680 11.0565 10.4940 12.1500 ;
      RECT 10.3600 11.0565 10.3860 12.1500 ;
      RECT 10.2520 11.0565 10.2780 12.1500 ;
      RECT 10.1440 11.0565 10.1700 12.1500 ;
      RECT 10.0360 11.0565 10.0620 12.1500 ;
      RECT 9.9280 11.0565 9.9540 12.1500 ;
      RECT 9.8200 11.0565 9.8460 12.1500 ;
      RECT 9.7120 11.0565 9.7380 12.1500 ;
      RECT 9.6040 11.0565 9.6300 12.1500 ;
      RECT 9.4960 11.0565 9.5220 12.1500 ;
      RECT 9.3880 11.0565 9.4140 12.1500 ;
      RECT 9.2800 11.0565 9.3060 12.1500 ;
      RECT 9.1720 11.0565 9.1980 12.1500 ;
      RECT 9.0640 11.0565 9.0900 12.1500 ;
      RECT 8.9560 11.0565 8.9820 12.1500 ;
      RECT 8.8480 11.0565 8.8740 12.1500 ;
      RECT 8.7400 11.0565 8.7660 12.1500 ;
      RECT 8.6320 11.0565 8.6580 12.1500 ;
      RECT 8.5240 11.0565 8.5500 12.1500 ;
      RECT 8.4160 11.0565 8.4420 12.1500 ;
      RECT 8.3080 11.0565 8.3340 12.1500 ;
      RECT 8.2000 11.0565 8.2260 12.1500 ;
      RECT 8.0920 11.0565 8.1180 12.1500 ;
      RECT 7.9840 11.0565 8.0100 12.1500 ;
      RECT 7.8760 11.0565 7.9020 12.1500 ;
      RECT 7.7680 11.0565 7.7940 12.1500 ;
      RECT 7.6600 11.0565 7.6860 12.1500 ;
      RECT 7.5520 11.0565 7.5780 12.1500 ;
      RECT 7.4440 11.0565 7.4700 12.1500 ;
      RECT 7.3360 11.0565 7.3620 12.1500 ;
      RECT 7.2280 11.0565 7.2540 12.1500 ;
      RECT 7.1200 11.0565 7.1460 12.1500 ;
      RECT 7.0120 11.0565 7.0380 12.1500 ;
      RECT 6.9040 11.0565 6.9300 12.1500 ;
      RECT 6.7960 11.0565 6.8220 12.1500 ;
      RECT 6.6880 11.0565 6.7140 12.1500 ;
      RECT 6.5800 11.0565 6.6060 12.1500 ;
      RECT 6.4720 11.0565 6.4980 12.1500 ;
      RECT 6.3640 11.0565 6.3900 12.1500 ;
      RECT 6.2560 11.0565 6.2820 12.1500 ;
      RECT 6.1480 11.0565 6.1740 12.1500 ;
      RECT 6.0400 11.0565 6.0660 12.1500 ;
      RECT 5.9320 11.0565 5.9580 12.1500 ;
      RECT 5.8240 11.0565 5.8500 12.1500 ;
      RECT 5.7160 11.0565 5.7420 12.1500 ;
      RECT 5.6080 11.0565 5.6340 12.1500 ;
      RECT 5.5000 11.0565 5.5260 12.1500 ;
      RECT 5.3920 11.0565 5.4180 12.1500 ;
      RECT 5.2840 11.0565 5.3100 12.1500 ;
      RECT 5.1760 11.0565 5.2020 12.1500 ;
      RECT 5.0680 11.0565 5.0940 12.1500 ;
      RECT 4.9600 11.0565 4.9860 12.1500 ;
      RECT 4.8520 11.0565 4.8780 12.1500 ;
      RECT 4.7440 11.0565 4.7700 12.1500 ;
      RECT 4.6360 11.0565 4.6620 12.1500 ;
      RECT 4.5280 11.0565 4.5540 12.1500 ;
      RECT 4.4200 11.0565 4.4460 12.1500 ;
      RECT 4.3120 11.0565 4.3380 12.1500 ;
      RECT 4.2040 11.0565 4.2300 12.1500 ;
      RECT 4.0960 11.0565 4.1220 12.1500 ;
      RECT 3.9880 11.0565 4.0140 12.1500 ;
      RECT 3.8800 11.0565 3.9060 12.1500 ;
      RECT 3.7720 11.0565 3.7980 12.1500 ;
      RECT 3.6640 11.0565 3.6900 12.1500 ;
      RECT 3.5560 11.0565 3.5820 12.1500 ;
      RECT 3.4480 11.0565 3.4740 12.1500 ;
      RECT 3.3400 11.0565 3.3660 12.1500 ;
      RECT 3.2320 11.0565 3.2580 12.1500 ;
      RECT 3.1240 11.0565 3.1500 12.1500 ;
      RECT 3.0160 11.0565 3.0420 12.1500 ;
      RECT 2.9080 11.0565 2.9340 12.1500 ;
      RECT 2.8000 11.0565 2.8260 12.1500 ;
      RECT 2.6920 11.0565 2.7180 12.1500 ;
      RECT 2.5840 11.0565 2.6100 12.1500 ;
      RECT 2.4760 11.0565 2.5020 12.1500 ;
      RECT 2.3680 11.0565 2.3940 12.1500 ;
      RECT 2.2600 11.0565 2.2860 12.1500 ;
      RECT 2.1520 11.0565 2.1780 12.1500 ;
      RECT 2.0440 11.0565 2.0700 12.1500 ;
      RECT 1.9360 11.0565 1.9620 12.1500 ;
      RECT 1.8280 11.0565 1.8540 12.1500 ;
      RECT 1.7200 11.0565 1.7460 12.1500 ;
      RECT 1.6120 11.0565 1.6380 12.1500 ;
      RECT 1.5040 11.0565 1.5300 12.1500 ;
      RECT 1.3960 11.0565 1.4220 12.1500 ;
      RECT 1.2880 11.0565 1.3140 12.1500 ;
      RECT 1.1800 11.0565 1.2060 12.1500 ;
      RECT 1.0720 11.0565 1.0980 12.1500 ;
      RECT 0.9640 11.0565 0.9900 12.1500 ;
      RECT 0.8560 11.0565 0.8820 12.1500 ;
      RECT 0.7480 11.0565 0.7740 12.1500 ;
      RECT 0.6400 11.0565 0.6660 12.1500 ;
      RECT 0.5320 11.0565 0.5580 12.1500 ;
      RECT 0.4240 11.0565 0.4500 12.1500 ;
      RECT 0.3160 11.0565 0.3420 12.1500 ;
      RECT 0.2080 11.0565 0.2340 12.1500 ;
      RECT 0.0050 11.0565 0.0900 12.1500 ;
      RECT 15.5530 12.1365 15.6810 13.2300 ;
      RECT 15.5390 12.8020 15.6810 13.1245 ;
      RECT 15.3190 12.5290 15.4530 13.2300 ;
      RECT 15.2960 12.8640 15.4530 13.1220 ;
      RECT 15.3190 12.1365 15.4170 13.2300 ;
      RECT 15.3190 12.2575 15.4310 12.4970 ;
      RECT 15.3190 12.1365 15.4530 12.2255 ;
      RECT 15.0940 12.5870 15.2280 13.2300 ;
      RECT 15.0940 12.1365 15.1920 13.2300 ;
      RECT 14.6770 12.1365 14.7600 13.2300 ;
      RECT 14.6770 12.2250 14.7740 13.1605 ;
      RECT 30.2680 12.1365 30.3530 13.2300 ;
      RECT 30.1240 12.1365 30.1500 13.2300 ;
      RECT 30.0160 12.1365 30.0420 13.2300 ;
      RECT 29.9080 12.1365 29.9340 13.2300 ;
      RECT 29.8000 12.1365 29.8260 13.2300 ;
      RECT 29.6920 12.1365 29.7180 13.2300 ;
      RECT 29.5840 12.1365 29.6100 13.2300 ;
      RECT 29.4760 12.1365 29.5020 13.2300 ;
      RECT 29.3680 12.1365 29.3940 13.2300 ;
      RECT 29.2600 12.1365 29.2860 13.2300 ;
      RECT 29.1520 12.1365 29.1780 13.2300 ;
      RECT 29.0440 12.1365 29.0700 13.2300 ;
      RECT 28.9360 12.1365 28.9620 13.2300 ;
      RECT 28.8280 12.1365 28.8540 13.2300 ;
      RECT 28.7200 12.1365 28.7460 13.2300 ;
      RECT 28.6120 12.1365 28.6380 13.2300 ;
      RECT 28.5040 12.1365 28.5300 13.2300 ;
      RECT 28.3960 12.1365 28.4220 13.2300 ;
      RECT 28.2880 12.1365 28.3140 13.2300 ;
      RECT 28.1800 12.1365 28.2060 13.2300 ;
      RECT 28.0720 12.1365 28.0980 13.2300 ;
      RECT 27.9640 12.1365 27.9900 13.2300 ;
      RECT 27.8560 12.1365 27.8820 13.2300 ;
      RECT 27.7480 12.1365 27.7740 13.2300 ;
      RECT 27.6400 12.1365 27.6660 13.2300 ;
      RECT 27.5320 12.1365 27.5580 13.2300 ;
      RECT 27.4240 12.1365 27.4500 13.2300 ;
      RECT 27.3160 12.1365 27.3420 13.2300 ;
      RECT 27.2080 12.1365 27.2340 13.2300 ;
      RECT 27.1000 12.1365 27.1260 13.2300 ;
      RECT 26.9920 12.1365 27.0180 13.2300 ;
      RECT 26.8840 12.1365 26.9100 13.2300 ;
      RECT 26.7760 12.1365 26.8020 13.2300 ;
      RECT 26.6680 12.1365 26.6940 13.2300 ;
      RECT 26.5600 12.1365 26.5860 13.2300 ;
      RECT 26.4520 12.1365 26.4780 13.2300 ;
      RECT 26.3440 12.1365 26.3700 13.2300 ;
      RECT 26.2360 12.1365 26.2620 13.2300 ;
      RECT 26.1280 12.1365 26.1540 13.2300 ;
      RECT 26.0200 12.1365 26.0460 13.2300 ;
      RECT 25.9120 12.1365 25.9380 13.2300 ;
      RECT 25.8040 12.1365 25.8300 13.2300 ;
      RECT 25.6960 12.1365 25.7220 13.2300 ;
      RECT 25.5880 12.1365 25.6140 13.2300 ;
      RECT 25.4800 12.1365 25.5060 13.2300 ;
      RECT 25.3720 12.1365 25.3980 13.2300 ;
      RECT 25.2640 12.1365 25.2900 13.2300 ;
      RECT 25.1560 12.1365 25.1820 13.2300 ;
      RECT 25.0480 12.1365 25.0740 13.2300 ;
      RECT 24.9400 12.1365 24.9660 13.2300 ;
      RECT 24.8320 12.1365 24.8580 13.2300 ;
      RECT 24.7240 12.1365 24.7500 13.2300 ;
      RECT 24.6160 12.1365 24.6420 13.2300 ;
      RECT 24.5080 12.1365 24.5340 13.2300 ;
      RECT 24.4000 12.1365 24.4260 13.2300 ;
      RECT 24.2920 12.1365 24.3180 13.2300 ;
      RECT 24.1840 12.1365 24.2100 13.2300 ;
      RECT 24.0760 12.1365 24.1020 13.2300 ;
      RECT 23.9680 12.1365 23.9940 13.2300 ;
      RECT 23.8600 12.1365 23.8860 13.2300 ;
      RECT 23.7520 12.1365 23.7780 13.2300 ;
      RECT 23.6440 12.1365 23.6700 13.2300 ;
      RECT 23.5360 12.1365 23.5620 13.2300 ;
      RECT 23.4280 12.1365 23.4540 13.2300 ;
      RECT 23.3200 12.1365 23.3460 13.2300 ;
      RECT 23.2120 12.1365 23.2380 13.2300 ;
      RECT 23.1040 12.1365 23.1300 13.2300 ;
      RECT 22.9960 12.1365 23.0220 13.2300 ;
      RECT 22.8880 12.1365 22.9140 13.2300 ;
      RECT 22.7800 12.1365 22.8060 13.2300 ;
      RECT 22.6720 12.1365 22.6980 13.2300 ;
      RECT 22.5640 12.1365 22.5900 13.2300 ;
      RECT 22.4560 12.1365 22.4820 13.2300 ;
      RECT 22.3480 12.1365 22.3740 13.2300 ;
      RECT 22.2400 12.1365 22.2660 13.2300 ;
      RECT 22.1320 12.1365 22.1580 13.2300 ;
      RECT 22.0240 12.1365 22.0500 13.2300 ;
      RECT 21.9160 12.1365 21.9420 13.2300 ;
      RECT 21.8080 12.1365 21.8340 13.2300 ;
      RECT 21.7000 12.1365 21.7260 13.2300 ;
      RECT 21.5920 12.1365 21.6180 13.2300 ;
      RECT 21.4840 12.1365 21.5100 13.2300 ;
      RECT 21.3760 12.1365 21.4020 13.2300 ;
      RECT 21.2680 12.1365 21.2940 13.2300 ;
      RECT 21.1600 12.1365 21.1860 13.2300 ;
      RECT 21.0520 12.1365 21.0780 13.2300 ;
      RECT 20.9440 12.1365 20.9700 13.2300 ;
      RECT 20.8360 12.1365 20.8620 13.2300 ;
      RECT 20.7280 12.1365 20.7540 13.2300 ;
      RECT 20.6200 12.1365 20.6460 13.2300 ;
      RECT 20.5120 12.1365 20.5380 13.2300 ;
      RECT 20.4040 12.1365 20.4300 13.2300 ;
      RECT 20.2960 12.1365 20.3220 13.2300 ;
      RECT 20.1880 12.1365 20.2140 13.2300 ;
      RECT 20.0800 12.1365 20.1060 13.2300 ;
      RECT 19.9720 12.1365 19.9980 13.2300 ;
      RECT 19.8640 12.1365 19.8900 13.2300 ;
      RECT 19.7560 12.1365 19.7820 13.2300 ;
      RECT 19.6480 12.1365 19.6740 13.2300 ;
      RECT 19.5400 12.1365 19.5660 13.2300 ;
      RECT 19.4320 12.1365 19.4580 13.2300 ;
      RECT 19.3240 12.1365 19.3500 13.2300 ;
      RECT 19.2160 12.1365 19.2420 13.2300 ;
      RECT 19.1080 12.1365 19.1340 13.2300 ;
      RECT 19.0000 12.1365 19.0260 13.2300 ;
      RECT 18.8920 12.1365 18.9180 13.2300 ;
      RECT 18.7840 12.1365 18.8100 13.2300 ;
      RECT 18.6760 12.1365 18.7020 13.2300 ;
      RECT 18.5680 12.1365 18.5940 13.2300 ;
      RECT 18.4600 12.1365 18.4860 13.2300 ;
      RECT 18.3520 12.1365 18.3780 13.2300 ;
      RECT 18.2440 12.1365 18.2700 13.2300 ;
      RECT 18.1360 12.1365 18.1620 13.2300 ;
      RECT 18.0280 12.1365 18.0540 13.2300 ;
      RECT 17.9200 12.1365 17.9460 13.2300 ;
      RECT 17.8120 12.1365 17.8380 13.2300 ;
      RECT 17.7040 12.1365 17.7300 13.2300 ;
      RECT 17.5960 12.1365 17.6220 13.2300 ;
      RECT 17.4880 12.1365 17.5140 13.2300 ;
      RECT 17.3800 12.1365 17.4060 13.2300 ;
      RECT 17.2720 12.1365 17.2980 13.2300 ;
      RECT 17.1640 12.1365 17.1900 13.2300 ;
      RECT 17.0560 12.1365 17.0820 13.2300 ;
      RECT 16.9480 12.1365 16.9740 13.2300 ;
      RECT 16.8400 12.1365 16.8660 13.2300 ;
      RECT 16.7320 12.1365 16.7580 13.2300 ;
      RECT 16.6240 12.1365 16.6500 13.2300 ;
      RECT 16.5160 12.1365 16.5420 13.2300 ;
      RECT 16.4080 12.1365 16.4340 13.2300 ;
      RECT 16.3000 12.1365 16.3260 13.2300 ;
      RECT 16.0870 12.1365 16.1640 13.2300 ;
      RECT 14.1940 12.1365 14.2710 13.2300 ;
      RECT 14.0320 12.1365 14.0580 13.2300 ;
      RECT 13.9240 12.1365 13.9500 13.2300 ;
      RECT 13.8160 12.1365 13.8420 13.2300 ;
      RECT 13.7080 12.1365 13.7340 13.2300 ;
      RECT 13.6000 12.1365 13.6260 13.2300 ;
      RECT 13.4920 12.1365 13.5180 13.2300 ;
      RECT 13.3840 12.1365 13.4100 13.2300 ;
      RECT 13.2760 12.1365 13.3020 13.2300 ;
      RECT 13.1680 12.1365 13.1940 13.2300 ;
      RECT 13.0600 12.1365 13.0860 13.2300 ;
      RECT 12.9520 12.1365 12.9780 13.2300 ;
      RECT 12.8440 12.1365 12.8700 13.2300 ;
      RECT 12.7360 12.1365 12.7620 13.2300 ;
      RECT 12.6280 12.1365 12.6540 13.2300 ;
      RECT 12.5200 12.1365 12.5460 13.2300 ;
      RECT 12.4120 12.1365 12.4380 13.2300 ;
      RECT 12.3040 12.1365 12.3300 13.2300 ;
      RECT 12.1960 12.1365 12.2220 13.2300 ;
      RECT 12.0880 12.1365 12.1140 13.2300 ;
      RECT 11.9800 12.1365 12.0060 13.2300 ;
      RECT 11.8720 12.1365 11.8980 13.2300 ;
      RECT 11.7640 12.1365 11.7900 13.2300 ;
      RECT 11.6560 12.1365 11.6820 13.2300 ;
      RECT 11.5480 12.1365 11.5740 13.2300 ;
      RECT 11.4400 12.1365 11.4660 13.2300 ;
      RECT 11.3320 12.1365 11.3580 13.2300 ;
      RECT 11.2240 12.1365 11.2500 13.2300 ;
      RECT 11.1160 12.1365 11.1420 13.2300 ;
      RECT 11.0080 12.1365 11.0340 13.2300 ;
      RECT 10.9000 12.1365 10.9260 13.2300 ;
      RECT 10.7920 12.1365 10.8180 13.2300 ;
      RECT 10.6840 12.1365 10.7100 13.2300 ;
      RECT 10.5760 12.1365 10.6020 13.2300 ;
      RECT 10.4680 12.1365 10.4940 13.2300 ;
      RECT 10.3600 12.1365 10.3860 13.2300 ;
      RECT 10.2520 12.1365 10.2780 13.2300 ;
      RECT 10.1440 12.1365 10.1700 13.2300 ;
      RECT 10.0360 12.1365 10.0620 13.2300 ;
      RECT 9.9280 12.1365 9.9540 13.2300 ;
      RECT 9.8200 12.1365 9.8460 13.2300 ;
      RECT 9.7120 12.1365 9.7380 13.2300 ;
      RECT 9.6040 12.1365 9.6300 13.2300 ;
      RECT 9.4960 12.1365 9.5220 13.2300 ;
      RECT 9.3880 12.1365 9.4140 13.2300 ;
      RECT 9.2800 12.1365 9.3060 13.2300 ;
      RECT 9.1720 12.1365 9.1980 13.2300 ;
      RECT 9.0640 12.1365 9.0900 13.2300 ;
      RECT 8.9560 12.1365 8.9820 13.2300 ;
      RECT 8.8480 12.1365 8.8740 13.2300 ;
      RECT 8.7400 12.1365 8.7660 13.2300 ;
      RECT 8.6320 12.1365 8.6580 13.2300 ;
      RECT 8.5240 12.1365 8.5500 13.2300 ;
      RECT 8.4160 12.1365 8.4420 13.2300 ;
      RECT 8.3080 12.1365 8.3340 13.2300 ;
      RECT 8.2000 12.1365 8.2260 13.2300 ;
      RECT 8.0920 12.1365 8.1180 13.2300 ;
      RECT 7.9840 12.1365 8.0100 13.2300 ;
      RECT 7.8760 12.1365 7.9020 13.2300 ;
      RECT 7.7680 12.1365 7.7940 13.2300 ;
      RECT 7.6600 12.1365 7.6860 13.2300 ;
      RECT 7.5520 12.1365 7.5780 13.2300 ;
      RECT 7.4440 12.1365 7.4700 13.2300 ;
      RECT 7.3360 12.1365 7.3620 13.2300 ;
      RECT 7.2280 12.1365 7.2540 13.2300 ;
      RECT 7.1200 12.1365 7.1460 13.2300 ;
      RECT 7.0120 12.1365 7.0380 13.2300 ;
      RECT 6.9040 12.1365 6.9300 13.2300 ;
      RECT 6.7960 12.1365 6.8220 13.2300 ;
      RECT 6.6880 12.1365 6.7140 13.2300 ;
      RECT 6.5800 12.1365 6.6060 13.2300 ;
      RECT 6.4720 12.1365 6.4980 13.2300 ;
      RECT 6.3640 12.1365 6.3900 13.2300 ;
      RECT 6.2560 12.1365 6.2820 13.2300 ;
      RECT 6.1480 12.1365 6.1740 13.2300 ;
      RECT 6.0400 12.1365 6.0660 13.2300 ;
      RECT 5.9320 12.1365 5.9580 13.2300 ;
      RECT 5.8240 12.1365 5.8500 13.2300 ;
      RECT 5.7160 12.1365 5.7420 13.2300 ;
      RECT 5.6080 12.1365 5.6340 13.2300 ;
      RECT 5.5000 12.1365 5.5260 13.2300 ;
      RECT 5.3920 12.1365 5.4180 13.2300 ;
      RECT 5.2840 12.1365 5.3100 13.2300 ;
      RECT 5.1760 12.1365 5.2020 13.2300 ;
      RECT 5.0680 12.1365 5.0940 13.2300 ;
      RECT 4.9600 12.1365 4.9860 13.2300 ;
      RECT 4.8520 12.1365 4.8780 13.2300 ;
      RECT 4.7440 12.1365 4.7700 13.2300 ;
      RECT 4.6360 12.1365 4.6620 13.2300 ;
      RECT 4.5280 12.1365 4.5540 13.2300 ;
      RECT 4.4200 12.1365 4.4460 13.2300 ;
      RECT 4.3120 12.1365 4.3380 13.2300 ;
      RECT 4.2040 12.1365 4.2300 13.2300 ;
      RECT 4.0960 12.1365 4.1220 13.2300 ;
      RECT 3.9880 12.1365 4.0140 13.2300 ;
      RECT 3.8800 12.1365 3.9060 13.2300 ;
      RECT 3.7720 12.1365 3.7980 13.2300 ;
      RECT 3.6640 12.1365 3.6900 13.2300 ;
      RECT 3.5560 12.1365 3.5820 13.2300 ;
      RECT 3.4480 12.1365 3.4740 13.2300 ;
      RECT 3.3400 12.1365 3.3660 13.2300 ;
      RECT 3.2320 12.1365 3.2580 13.2300 ;
      RECT 3.1240 12.1365 3.1500 13.2300 ;
      RECT 3.0160 12.1365 3.0420 13.2300 ;
      RECT 2.9080 12.1365 2.9340 13.2300 ;
      RECT 2.8000 12.1365 2.8260 13.2300 ;
      RECT 2.6920 12.1365 2.7180 13.2300 ;
      RECT 2.5840 12.1365 2.6100 13.2300 ;
      RECT 2.4760 12.1365 2.5020 13.2300 ;
      RECT 2.3680 12.1365 2.3940 13.2300 ;
      RECT 2.2600 12.1365 2.2860 13.2300 ;
      RECT 2.1520 12.1365 2.1780 13.2300 ;
      RECT 2.0440 12.1365 2.0700 13.2300 ;
      RECT 1.9360 12.1365 1.9620 13.2300 ;
      RECT 1.8280 12.1365 1.8540 13.2300 ;
      RECT 1.7200 12.1365 1.7460 13.2300 ;
      RECT 1.6120 12.1365 1.6380 13.2300 ;
      RECT 1.5040 12.1365 1.5300 13.2300 ;
      RECT 1.3960 12.1365 1.4220 13.2300 ;
      RECT 1.2880 12.1365 1.3140 13.2300 ;
      RECT 1.1800 12.1365 1.2060 13.2300 ;
      RECT 1.0720 12.1365 1.0980 13.2300 ;
      RECT 0.9640 12.1365 0.9900 13.2300 ;
      RECT 0.8560 12.1365 0.8820 13.2300 ;
      RECT 0.7480 12.1365 0.7740 13.2300 ;
      RECT 0.6400 12.1365 0.6660 13.2300 ;
      RECT 0.5320 12.1365 0.5580 13.2300 ;
      RECT 0.4240 12.1365 0.4500 13.2300 ;
      RECT 0.3160 12.1365 0.3420 13.2300 ;
      RECT 0.2080 12.1365 0.2340 13.2300 ;
      RECT 0.0050 12.1365 0.0900 13.2300 ;
      RECT 15.5530 13.2165 15.6810 14.3100 ;
      RECT 15.5390 13.8820 15.6810 14.2045 ;
      RECT 15.3190 13.6090 15.4530 14.3100 ;
      RECT 15.2960 13.9440 15.4530 14.2020 ;
      RECT 15.3190 13.2165 15.4170 14.3100 ;
      RECT 15.3190 13.3375 15.4310 13.5770 ;
      RECT 15.3190 13.2165 15.4530 13.3055 ;
      RECT 15.0940 13.6670 15.2280 14.3100 ;
      RECT 15.0940 13.2165 15.1920 14.3100 ;
      RECT 14.6770 13.2165 14.7600 14.3100 ;
      RECT 14.6770 13.3050 14.7740 14.2405 ;
      RECT 30.2680 13.2165 30.3530 14.3100 ;
      RECT 30.1240 13.2165 30.1500 14.3100 ;
      RECT 30.0160 13.2165 30.0420 14.3100 ;
      RECT 29.9080 13.2165 29.9340 14.3100 ;
      RECT 29.8000 13.2165 29.8260 14.3100 ;
      RECT 29.6920 13.2165 29.7180 14.3100 ;
      RECT 29.5840 13.2165 29.6100 14.3100 ;
      RECT 29.4760 13.2165 29.5020 14.3100 ;
      RECT 29.3680 13.2165 29.3940 14.3100 ;
      RECT 29.2600 13.2165 29.2860 14.3100 ;
      RECT 29.1520 13.2165 29.1780 14.3100 ;
      RECT 29.0440 13.2165 29.0700 14.3100 ;
      RECT 28.9360 13.2165 28.9620 14.3100 ;
      RECT 28.8280 13.2165 28.8540 14.3100 ;
      RECT 28.7200 13.2165 28.7460 14.3100 ;
      RECT 28.6120 13.2165 28.6380 14.3100 ;
      RECT 28.5040 13.2165 28.5300 14.3100 ;
      RECT 28.3960 13.2165 28.4220 14.3100 ;
      RECT 28.2880 13.2165 28.3140 14.3100 ;
      RECT 28.1800 13.2165 28.2060 14.3100 ;
      RECT 28.0720 13.2165 28.0980 14.3100 ;
      RECT 27.9640 13.2165 27.9900 14.3100 ;
      RECT 27.8560 13.2165 27.8820 14.3100 ;
      RECT 27.7480 13.2165 27.7740 14.3100 ;
      RECT 27.6400 13.2165 27.6660 14.3100 ;
      RECT 27.5320 13.2165 27.5580 14.3100 ;
      RECT 27.4240 13.2165 27.4500 14.3100 ;
      RECT 27.3160 13.2165 27.3420 14.3100 ;
      RECT 27.2080 13.2165 27.2340 14.3100 ;
      RECT 27.1000 13.2165 27.1260 14.3100 ;
      RECT 26.9920 13.2165 27.0180 14.3100 ;
      RECT 26.8840 13.2165 26.9100 14.3100 ;
      RECT 26.7760 13.2165 26.8020 14.3100 ;
      RECT 26.6680 13.2165 26.6940 14.3100 ;
      RECT 26.5600 13.2165 26.5860 14.3100 ;
      RECT 26.4520 13.2165 26.4780 14.3100 ;
      RECT 26.3440 13.2165 26.3700 14.3100 ;
      RECT 26.2360 13.2165 26.2620 14.3100 ;
      RECT 26.1280 13.2165 26.1540 14.3100 ;
      RECT 26.0200 13.2165 26.0460 14.3100 ;
      RECT 25.9120 13.2165 25.9380 14.3100 ;
      RECT 25.8040 13.2165 25.8300 14.3100 ;
      RECT 25.6960 13.2165 25.7220 14.3100 ;
      RECT 25.5880 13.2165 25.6140 14.3100 ;
      RECT 25.4800 13.2165 25.5060 14.3100 ;
      RECT 25.3720 13.2165 25.3980 14.3100 ;
      RECT 25.2640 13.2165 25.2900 14.3100 ;
      RECT 25.1560 13.2165 25.1820 14.3100 ;
      RECT 25.0480 13.2165 25.0740 14.3100 ;
      RECT 24.9400 13.2165 24.9660 14.3100 ;
      RECT 24.8320 13.2165 24.8580 14.3100 ;
      RECT 24.7240 13.2165 24.7500 14.3100 ;
      RECT 24.6160 13.2165 24.6420 14.3100 ;
      RECT 24.5080 13.2165 24.5340 14.3100 ;
      RECT 24.4000 13.2165 24.4260 14.3100 ;
      RECT 24.2920 13.2165 24.3180 14.3100 ;
      RECT 24.1840 13.2165 24.2100 14.3100 ;
      RECT 24.0760 13.2165 24.1020 14.3100 ;
      RECT 23.9680 13.2165 23.9940 14.3100 ;
      RECT 23.8600 13.2165 23.8860 14.3100 ;
      RECT 23.7520 13.2165 23.7780 14.3100 ;
      RECT 23.6440 13.2165 23.6700 14.3100 ;
      RECT 23.5360 13.2165 23.5620 14.3100 ;
      RECT 23.4280 13.2165 23.4540 14.3100 ;
      RECT 23.3200 13.2165 23.3460 14.3100 ;
      RECT 23.2120 13.2165 23.2380 14.3100 ;
      RECT 23.1040 13.2165 23.1300 14.3100 ;
      RECT 22.9960 13.2165 23.0220 14.3100 ;
      RECT 22.8880 13.2165 22.9140 14.3100 ;
      RECT 22.7800 13.2165 22.8060 14.3100 ;
      RECT 22.6720 13.2165 22.6980 14.3100 ;
      RECT 22.5640 13.2165 22.5900 14.3100 ;
      RECT 22.4560 13.2165 22.4820 14.3100 ;
      RECT 22.3480 13.2165 22.3740 14.3100 ;
      RECT 22.2400 13.2165 22.2660 14.3100 ;
      RECT 22.1320 13.2165 22.1580 14.3100 ;
      RECT 22.0240 13.2165 22.0500 14.3100 ;
      RECT 21.9160 13.2165 21.9420 14.3100 ;
      RECT 21.8080 13.2165 21.8340 14.3100 ;
      RECT 21.7000 13.2165 21.7260 14.3100 ;
      RECT 21.5920 13.2165 21.6180 14.3100 ;
      RECT 21.4840 13.2165 21.5100 14.3100 ;
      RECT 21.3760 13.2165 21.4020 14.3100 ;
      RECT 21.2680 13.2165 21.2940 14.3100 ;
      RECT 21.1600 13.2165 21.1860 14.3100 ;
      RECT 21.0520 13.2165 21.0780 14.3100 ;
      RECT 20.9440 13.2165 20.9700 14.3100 ;
      RECT 20.8360 13.2165 20.8620 14.3100 ;
      RECT 20.7280 13.2165 20.7540 14.3100 ;
      RECT 20.6200 13.2165 20.6460 14.3100 ;
      RECT 20.5120 13.2165 20.5380 14.3100 ;
      RECT 20.4040 13.2165 20.4300 14.3100 ;
      RECT 20.2960 13.2165 20.3220 14.3100 ;
      RECT 20.1880 13.2165 20.2140 14.3100 ;
      RECT 20.0800 13.2165 20.1060 14.3100 ;
      RECT 19.9720 13.2165 19.9980 14.3100 ;
      RECT 19.8640 13.2165 19.8900 14.3100 ;
      RECT 19.7560 13.2165 19.7820 14.3100 ;
      RECT 19.6480 13.2165 19.6740 14.3100 ;
      RECT 19.5400 13.2165 19.5660 14.3100 ;
      RECT 19.4320 13.2165 19.4580 14.3100 ;
      RECT 19.3240 13.2165 19.3500 14.3100 ;
      RECT 19.2160 13.2165 19.2420 14.3100 ;
      RECT 19.1080 13.2165 19.1340 14.3100 ;
      RECT 19.0000 13.2165 19.0260 14.3100 ;
      RECT 18.8920 13.2165 18.9180 14.3100 ;
      RECT 18.7840 13.2165 18.8100 14.3100 ;
      RECT 18.6760 13.2165 18.7020 14.3100 ;
      RECT 18.5680 13.2165 18.5940 14.3100 ;
      RECT 18.4600 13.2165 18.4860 14.3100 ;
      RECT 18.3520 13.2165 18.3780 14.3100 ;
      RECT 18.2440 13.2165 18.2700 14.3100 ;
      RECT 18.1360 13.2165 18.1620 14.3100 ;
      RECT 18.0280 13.2165 18.0540 14.3100 ;
      RECT 17.9200 13.2165 17.9460 14.3100 ;
      RECT 17.8120 13.2165 17.8380 14.3100 ;
      RECT 17.7040 13.2165 17.7300 14.3100 ;
      RECT 17.5960 13.2165 17.6220 14.3100 ;
      RECT 17.4880 13.2165 17.5140 14.3100 ;
      RECT 17.3800 13.2165 17.4060 14.3100 ;
      RECT 17.2720 13.2165 17.2980 14.3100 ;
      RECT 17.1640 13.2165 17.1900 14.3100 ;
      RECT 17.0560 13.2165 17.0820 14.3100 ;
      RECT 16.9480 13.2165 16.9740 14.3100 ;
      RECT 16.8400 13.2165 16.8660 14.3100 ;
      RECT 16.7320 13.2165 16.7580 14.3100 ;
      RECT 16.6240 13.2165 16.6500 14.3100 ;
      RECT 16.5160 13.2165 16.5420 14.3100 ;
      RECT 16.4080 13.2165 16.4340 14.3100 ;
      RECT 16.3000 13.2165 16.3260 14.3100 ;
      RECT 16.0870 13.2165 16.1640 14.3100 ;
      RECT 14.1940 13.2165 14.2710 14.3100 ;
      RECT 14.0320 13.2165 14.0580 14.3100 ;
      RECT 13.9240 13.2165 13.9500 14.3100 ;
      RECT 13.8160 13.2165 13.8420 14.3100 ;
      RECT 13.7080 13.2165 13.7340 14.3100 ;
      RECT 13.6000 13.2165 13.6260 14.3100 ;
      RECT 13.4920 13.2165 13.5180 14.3100 ;
      RECT 13.3840 13.2165 13.4100 14.3100 ;
      RECT 13.2760 13.2165 13.3020 14.3100 ;
      RECT 13.1680 13.2165 13.1940 14.3100 ;
      RECT 13.0600 13.2165 13.0860 14.3100 ;
      RECT 12.9520 13.2165 12.9780 14.3100 ;
      RECT 12.8440 13.2165 12.8700 14.3100 ;
      RECT 12.7360 13.2165 12.7620 14.3100 ;
      RECT 12.6280 13.2165 12.6540 14.3100 ;
      RECT 12.5200 13.2165 12.5460 14.3100 ;
      RECT 12.4120 13.2165 12.4380 14.3100 ;
      RECT 12.3040 13.2165 12.3300 14.3100 ;
      RECT 12.1960 13.2165 12.2220 14.3100 ;
      RECT 12.0880 13.2165 12.1140 14.3100 ;
      RECT 11.9800 13.2165 12.0060 14.3100 ;
      RECT 11.8720 13.2165 11.8980 14.3100 ;
      RECT 11.7640 13.2165 11.7900 14.3100 ;
      RECT 11.6560 13.2165 11.6820 14.3100 ;
      RECT 11.5480 13.2165 11.5740 14.3100 ;
      RECT 11.4400 13.2165 11.4660 14.3100 ;
      RECT 11.3320 13.2165 11.3580 14.3100 ;
      RECT 11.2240 13.2165 11.2500 14.3100 ;
      RECT 11.1160 13.2165 11.1420 14.3100 ;
      RECT 11.0080 13.2165 11.0340 14.3100 ;
      RECT 10.9000 13.2165 10.9260 14.3100 ;
      RECT 10.7920 13.2165 10.8180 14.3100 ;
      RECT 10.6840 13.2165 10.7100 14.3100 ;
      RECT 10.5760 13.2165 10.6020 14.3100 ;
      RECT 10.4680 13.2165 10.4940 14.3100 ;
      RECT 10.3600 13.2165 10.3860 14.3100 ;
      RECT 10.2520 13.2165 10.2780 14.3100 ;
      RECT 10.1440 13.2165 10.1700 14.3100 ;
      RECT 10.0360 13.2165 10.0620 14.3100 ;
      RECT 9.9280 13.2165 9.9540 14.3100 ;
      RECT 9.8200 13.2165 9.8460 14.3100 ;
      RECT 9.7120 13.2165 9.7380 14.3100 ;
      RECT 9.6040 13.2165 9.6300 14.3100 ;
      RECT 9.4960 13.2165 9.5220 14.3100 ;
      RECT 9.3880 13.2165 9.4140 14.3100 ;
      RECT 9.2800 13.2165 9.3060 14.3100 ;
      RECT 9.1720 13.2165 9.1980 14.3100 ;
      RECT 9.0640 13.2165 9.0900 14.3100 ;
      RECT 8.9560 13.2165 8.9820 14.3100 ;
      RECT 8.8480 13.2165 8.8740 14.3100 ;
      RECT 8.7400 13.2165 8.7660 14.3100 ;
      RECT 8.6320 13.2165 8.6580 14.3100 ;
      RECT 8.5240 13.2165 8.5500 14.3100 ;
      RECT 8.4160 13.2165 8.4420 14.3100 ;
      RECT 8.3080 13.2165 8.3340 14.3100 ;
      RECT 8.2000 13.2165 8.2260 14.3100 ;
      RECT 8.0920 13.2165 8.1180 14.3100 ;
      RECT 7.9840 13.2165 8.0100 14.3100 ;
      RECT 7.8760 13.2165 7.9020 14.3100 ;
      RECT 7.7680 13.2165 7.7940 14.3100 ;
      RECT 7.6600 13.2165 7.6860 14.3100 ;
      RECT 7.5520 13.2165 7.5780 14.3100 ;
      RECT 7.4440 13.2165 7.4700 14.3100 ;
      RECT 7.3360 13.2165 7.3620 14.3100 ;
      RECT 7.2280 13.2165 7.2540 14.3100 ;
      RECT 7.1200 13.2165 7.1460 14.3100 ;
      RECT 7.0120 13.2165 7.0380 14.3100 ;
      RECT 6.9040 13.2165 6.9300 14.3100 ;
      RECT 6.7960 13.2165 6.8220 14.3100 ;
      RECT 6.6880 13.2165 6.7140 14.3100 ;
      RECT 6.5800 13.2165 6.6060 14.3100 ;
      RECT 6.4720 13.2165 6.4980 14.3100 ;
      RECT 6.3640 13.2165 6.3900 14.3100 ;
      RECT 6.2560 13.2165 6.2820 14.3100 ;
      RECT 6.1480 13.2165 6.1740 14.3100 ;
      RECT 6.0400 13.2165 6.0660 14.3100 ;
      RECT 5.9320 13.2165 5.9580 14.3100 ;
      RECT 5.8240 13.2165 5.8500 14.3100 ;
      RECT 5.7160 13.2165 5.7420 14.3100 ;
      RECT 5.6080 13.2165 5.6340 14.3100 ;
      RECT 5.5000 13.2165 5.5260 14.3100 ;
      RECT 5.3920 13.2165 5.4180 14.3100 ;
      RECT 5.2840 13.2165 5.3100 14.3100 ;
      RECT 5.1760 13.2165 5.2020 14.3100 ;
      RECT 5.0680 13.2165 5.0940 14.3100 ;
      RECT 4.9600 13.2165 4.9860 14.3100 ;
      RECT 4.8520 13.2165 4.8780 14.3100 ;
      RECT 4.7440 13.2165 4.7700 14.3100 ;
      RECT 4.6360 13.2165 4.6620 14.3100 ;
      RECT 4.5280 13.2165 4.5540 14.3100 ;
      RECT 4.4200 13.2165 4.4460 14.3100 ;
      RECT 4.3120 13.2165 4.3380 14.3100 ;
      RECT 4.2040 13.2165 4.2300 14.3100 ;
      RECT 4.0960 13.2165 4.1220 14.3100 ;
      RECT 3.9880 13.2165 4.0140 14.3100 ;
      RECT 3.8800 13.2165 3.9060 14.3100 ;
      RECT 3.7720 13.2165 3.7980 14.3100 ;
      RECT 3.6640 13.2165 3.6900 14.3100 ;
      RECT 3.5560 13.2165 3.5820 14.3100 ;
      RECT 3.4480 13.2165 3.4740 14.3100 ;
      RECT 3.3400 13.2165 3.3660 14.3100 ;
      RECT 3.2320 13.2165 3.2580 14.3100 ;
      RECT 3.1240 13.2165 3.1500 14.3100 ;
      RECT 3.0160 13.2165 3.0420 14.3100 ;
      RECT 2.9080 13.2165 2.9340 14.3100 ;
      RECT 2.8000 13.2165 2.8260 14.3100 ;
      RECT 2.6920 13.2165 2.7180 14.3100 ;
      RECT 2.5840 13.2165 2.6100 14.3100 ;
      RECT 2.4760 13.2165 2.5020 14.3100 ;
      RECT 2.3680 13.2165 2.3940 14.3100 ;
      RECT 2.2600 13.2165 2.2860 14.3100 ;
      RECT 2.1520 13.2165 2.1780 14.3100 ;
      RECT 2.0440 13.2165 2.0700 14.3100 ;
      RECT 1.9360 13.2165 1.9620 14.3100 ;
      RECT 1.8280 13.2165 1.8540 14.3100 ;
      RECT 1.7200 13.2165 1.7460 14.3100 ;
      RECT 1.6120 13.2165 1.6380 14.3100 ;
      RECT 1.5040 13.2165 1.5300 14.3100 ;
      RECT 1.3960 13.2165 1.4220 14.3100 ;
      RECT 1.2880 13.2165 1.3140 14.3100 ;
      RECT 1.1800 13.2165 1.2060 14.3100 ;
      RECT 1.0720 13.2165 1.0980 14.3100 ;
      RECT 0.9640 13.2165 0.9900 14.3100 ;
      RECT 0.8560 13.2165 0.8820 14.3100 ;
      RECT 0.7480 13.2165 0.7740 14.3100 ;
      RECT 0.6400 13.2165 0.6660 14.3100 ;
      RECT 0.5320 13.2165 0.5580 14.3100 ;
      RECT 0.4240 13.2165 0.4500 14.3100 ;
      RECT 0.3160 13.2165 0.3420 14.3100 ;
      RECT 0.2080 13.2165 0.2340 14.3100 ;
      RECT 0.0050 13.2165 0.0900 14.3100 ;
      RECT 15.5530 14.2965 15.6810 15.3900 ;
      RECT 15.5390 14.9620 15.6810 15.2845 ;
      RECT 15.3190 14.6890 15.4530 15.3900 ;
      RECT 15.2960 15.0240 15.4530 15.2820 ;
      RECT 15.3190 14.2965 15.4170 15.3900 ;
      RECT 15.3190 14.4175 15.4310 14.6570 ;
      RECT 15.3190 14.2965 15.4530 14.3855 ;
      RECT 15.0940 14.7470 15.2280 15.3900 ;
      RECT 15.0940 14.2965 15.1920 15.3900 ;
      RECT 14.6770 14.2965 14.7600 15.3900 ;
      RECT 14.6770 14.3850 14.7740 15.3205 ;
      RECT 30.2680 14.2965 30.3530 15.3900 ;
      RECT 30.1240 14.2965 30.1500 15.3900 ;
      RECT 30.0160 14.2965 30.0420 15.3900 ;
      RECT 29.9080 14.2965 29.9340 15.3900 ;
      RECT 29.8000 14.2965 29.8260 15.3900 ;
      RECT 29.6920 14.2965 29.7180 15.3900 ;
      RECT 29.5840 14.2965 29.6100 15.3900 ;
      RECT 29.4760 14.2965 29.5020 15.3900 ;
      RECT 29.3680 14.2965 29.3940 15.3900 ;
      RECT 29.2600 14.2965 29.2860 15.3900 ;
      RECT 29.1520 14.2965 29.1780 15.3900 ;
      RECT 29.0440 14.2965 29.0700 15.3900 ;
      RECT 28.9360 14.2965 28.9620 15.3900 ;
      RECT 28.8280 14.2965 28.8540 15.3900 ;
      RECT 28.7200 14.2965 28.7460 15.3900 ;
      RECT 28.6120 14.2965 28.6380 15.3900 ;
      RECT 28.5040 14.2965 28.5300 15.3900 ;
      RECT 28.3960 14.2965 28.4220 15.3900 ;
      RECT 28.2880 14.2965 28.3140 15.3900 ;
      RECT 28.1800 14.2965 28.2060 15.3900 ;
      RECT 28.0720 14.2965 28.0980 15.3900 ;
      RECT 27.9640 14.2965 27.9900 15.3900 ;
      RECT 27.8560 14.2965 27.8820 15.3900 ;
      RECT 27.7480 14.2965 27.7740 15.3900 ;
      RECT 27.6400 14.2965 27.6660 15.3900 ;
      RECT 27.5320 14.2965 27.5580 15.3900 ;
      RECT 27.4240 14.2965 27.4500 15.3900 ;
      RECT 27.3160 14.2965 27.3420 15.3900 ;
      RECT 27.2080 14.2965 27.2340 15.3900 ;
      RECT 27.1000 14.2965 27.1260 15.3900 ;
      RECT 26.9920 14.2965 27.0180 15.3900 ;
      RECT 26.8840 14.2965 26.9100 15.3900 ;
      RECT 26.7760 14.2965 26.8020 15.3900 ;
      RECT 26.6680 14.2965 26.6940 15.3900 ;
      RECT 26.5600 14.2965 26.5860 15.3900 ;
      RECT 26.4520 14.2965 26.4780 15.3900 ;
      RECT 26.3440 14.2965 26.3700 15.3900 ;
      RECT 26.2360 14.2965 26.2620 15.3900 ;
      RECT 26.1280 14.2965 26.1540 15.3900 ;
      RECT 26.0200 14.2965 26.0460 15.3900 ;
      RECT 25.9120 14.2965 25.9380 15.3900 ;
      RECT 25.8040 14.2965 25.8300 15.3900 ;
      RECT 25.6960 14.2965 25.7220 15.3900 ;
      RECT 25.5880 14.2965 25.6140 15.3900 ;
      RECT 25.4800 14.2965 25.5060 15.3900 ;
      RECT 25.3720 14.2965 25.3980 15.3900 ;
      RECT 25.2640 14.2965 25.2900 15.3900 ;
      RECT 25.1560 14.2965 25.1820 15.3900 ;
      RECT 25.0480 14.2965 25.0740 15.3900 ;
      RECT 24.9400 14.2965 24.9660 15.3900 ;
      RECT 24.8320 14.2965 24.8580 15.3900 ;
      RECT 24.7240 14.2965 24.7500 15.3900 ;
      RECT 24.6160 14.2965 24.6420 15.3900 ;
      RECT 24.5080 14.2965 24.5340 15.3900 ;
      RECT 24.4000 14.2965 24.4260 15.3900 ;
      RECT 24.2920 14.2965 24.3180 15.3900 ;
      RECT 24.1840 14.2965 24.2100 15.3900 ;
      RECT 24.0760 14.2965 24.1020 15.3900 ;
      RECT 23.9680 14.2965 23.9940 15.3900 ;
      RECT 23.8600 14.2965 23.8860 15.3900 ;
      RECT 23.7520 14.2965 23.7780 15.3900 ;
      RECT 23.6440 14.2965 23.6700 15.3900 ;
      RECT 23.5360 14.2965 23.5620 15.3900 ;
      RECT 23.4280 14.2965 23.4540 15.3900 ;
      RECT 23.3200 14.2965 23.3460 15.3900 ;
      RECT 23.2120 14.2965 23.2380 15.3900 ;
      RECT 23.1040 14.2965 23.1300 15.3900 ;
      RECT 22.9960 14.2965 23.0220 15.3900 ;
      RECT 22.8880 14.2965 22.9140 15.3900 ;
      RECT 22.7800 14.2965 22.8060 15.3900 ;
      RECT 22.6720 14.2965 22.6980 15.3900 ;
      RECT 22.5640 14.2965 22.5900 15.3900 ;
      RECT 22.4560 14.2965 22.4820 15.3900 ;
      RECT 22.3480 14.2965 22.3740 15.3900 ;
      RECT 22.2400 14.2965 22.2660 15.3900 ;
      RECT 22.1320 14.2965 22.1580 15.3900 ;
      RECT 22.0240 14.2965 22.0500 15.3900 ;
      RECT 21.9160 14.2965 21.9420 15.3900 ;
      RECT 21.8080 14.2965 21.8340 15.3900 ;
      RECT 21.7000 14.2965 21.7260 15.3900 ;
      RECT 21.5920 14.2965 21.6180 15.3900 ;
      RECT 21.4840 14.2965 21.5100 15.3900 ;
      RECT 21.3760 14.2965 21.4020 15.3900 ;
      RECT 21.2680 14.2965 21.2940 15.3900 ;
      RECT 21.1600 14.2965 21.1860 15.3900 ;
      RECT 21.0520 14.2965 21.0780 15.3900 ;
      RECT 20.9440 14.2965 20.9700 15.3900 ;
      RECT 20.8360 14.2965 20.8620 15.3900 ;
      RECT 20.7280 14.2965 20.7540 15.3900 ;
      RECT 20.6200 14.2965 20.6460 15.3900 ;
      RECT 20.5120 14.2965 20.5380 15.3900 ;
      RECT 20.4040 14.2965 20.4300 15.3900 ;
      RECT 20.2960 14.2965 20.3220 15.3900 ;
      RECT 20.1880 14.2965 20.2140 15.3900 ;
      RECT 20.0800 14.2965 20.1060 15.3900 ;
      RECT 19.9720 14.2965 19.9980 15.3900 ;
      RECT 19.8640 14.2965 19.8900 15.3900 ;
      RECT 19.7560 14.2965 19.7820 15.3900 ;
      RECT 19.6480 14.2965 19.6740 15.3900 ;
      RECT 19.5400 14.2965 19.5660 15.3900 ;
      RECT 19.4320 14.2965 19.4580 15.3900 ;
      RECT 19.3240 14.2965 19.3500 15.3900 ;
      RECT 19.2160 14.2965 19.2420 15.3900 ;
      RECT 19.1080 14.2965 19.1340 15.3900 ;
      RECT 19.0000 14.2965 19.0260 15.3900 ;
      RECT 18.8920 14.2965 18.9180 15.3900 ;
      RECT 18.7840 14.2965 18.8100 15.3900 ;
      RECT 18.6760 14.2965 18.7020 15.3900 ;
      RECT 18.5680 14.2965 18.5940 15.3900 ;
      RECT 18.4600 14.2965 18.4860 15.3900 ;
      RECT 18.3520 14.2965 18.3780 15.3900 ;
      RECT 18.2440 14.2965 18.2700 15.3900 ;
      RECT 18.1360 14.2965 18.1620 15.3900 ;
      RECT 18.0280 14.2965 18.0540 15.3900 ;
      RECT 17.9200 14.2965 17.9460 15.3900 ;
      RECT 17.8120 14.2965 17.8380 15.3900 ;
      RECT 17.7040 14.2965 17.7300 15.3900 ;
      RECT 17.5960 14.2965 17.6220 15.3900 ;
      RECT 17.4880 14.2965 17.5140 15.3900 ;
      RECT 17.3800 14.2965 17.4060 15.3900 ;
      RECT 17.2720 14.2965 17.2980 15.3900 ;
      RECT 17.1640 14.2965 17.1900 15.3900 ;
      RECT 17.0560 14.2965 17.0820 15.3900 ;
      RECT 16.9480 14.2965 16.9740 15.3900 ;
      RECT 16.8400 14.2965 16.8660 15.3900 ;
      RECT 16.7320 14.2965 16.7580 15.3900 ;
      RECT 16.6240 14.2965 16.6500 15.3900 ;
      RECT 16.5160 14.2965 16.5420 15.3900 ;
      RECT 16.4080 14.2965 16.4340 15.3900 ;
      RECT 16.3000 14.2965 16.3260 15.3900 ;
      RECT 16.0870 14.2965 16.1640 15.3900 ;
      RECT 14.1940 14.2965 14.2710 15.3900 ;
      RECT 14.0320 14.2965 14.0580 15.3900 ;
      RECT 13.9240 14.2965 13.9500 15.3900 ;
      RECT 13.8160 14.2965 13.8420 15.3900 ;
      RECT 13.7080 14.2965 13.7340 15.3900 ;
      RECT 13.6000 14.2965 13.6260 15.3900 ;
      RECT 13.4920 14.2965 13.5180 15.3900 ;
      RECT 13.3840 14.2965 13.4100 15.3900 ;
      RECT 13.2760 14.2965 13.3020 15.3900 ;
      RECT 13.1680 14.2965 13.1940 15.3900 ;
      RECT 13.0600 14.2965 13.0860 15.3900 ;
      RECT 12.9520 14.2965 12.9780 15.3900 ;
      RECT 12.8440 14.2965 12.8700 15.3900 ;
      RECT 12.7360 14.2965 12.7620 15.3900 ;
      RECT 12.6280 14.2965 12.6540 15.3900 ;
      RECT 12.5200 14.2965 12.5460 15.3900 ;
      RECT 12.4120 14.2965 12.4380 15.3900 ;
      RECT 12.3040 14.2965 12.3300 15.3900 ;
      RECT 12.1960 14.2965 12.2220 15.3900 ;
      RECT 12.0880 14.2965 12.1140 15.3900 ;
      RECT 11.9800 14.2965 12.0060 15.3900 ;
      RECT 11.8720 14.2965 11.8980 15.3900 ;
      RECT 11.7640 14.2965 11.7900 15.3900 ;
      RECT 11.6560 14.2965 11.6820 15.3900 ;
      RECT 11.5480 14.2965 11.5740 15.3900 ;
      RECT 11.4400 14.2965 11.4660 15.3900 ;
      RECT 11.3320 14.2965 11.3580 15.3900 ;
      RECT 11.2240 14.2965 11.2500 15.3900 ;
      RECT 11.1160 14.2965 11.1420 15.3900 ;
      RECT 11.0080 14.2965 11.0340 15.3900 ;
      RECT 10.9000 14.2965 10.9260 15.3900 ;
      RECT 10.7920 14.2965 10.8180 15.3900 ;
      RECT 10.6840 14.2965 10.7100 15.3900 ;
      RECT 10.5760 14.2965 10.6020 15.3900 ;
      RECT 10.4680 14.2965 10.4940 15.3900 ;
      RECT 10.3600 14.2965 10.3860 15.3900 ;
      RECT 10.2520 14.2965 10.2780 15.3900 ;
      RECT 10.1440 14.2965 10.1700 15.3900 ;
      RECT 10.0360 14.2965 10.0620 15.3900 ;
      RECT 9.9280 14.2965 9.9540 15.3900 ;
      RECT 9.8200 14.2965 9.8460 15.3900 ;
      RECT 9.7120 14.2965 9.7380 15.3900 ;
      RECT 9.6040 14.2965 9.6300 15.3900 ;
      RECT 9.4960 14.2965 9.5220 15.3900 ;
      RECT 9.3880 14.2965 9.4140 15.3900 ;
      RECT 9.2800 14.2965 9.3060 15.3900 ;
      RECT 9.1720 14.2965 9.1980 15.3900 ;
      RECT 9.0640 14.2965 9.0900 15.3900 ;
      RECT 8.9560 14.2965 8.9820 15.3900 ;
      RECT 8.8480 14.2965 8.8740 15.3900 ;
      RECT 8.7400 14.2965 8.7660 15.3900 ;
      RECT 8.6320 14.2965 8.6580 15.3900 ;
      RECT 8.5240 14.2965 8.5500 15.3900 ;
      RECT 8.4160 14.2965 8.4420 15.3900 ;
      RECT 8.3080 14.2965 8.3340 15.3900 ;
      RECT 8.2000 14.2965 8.2260 15.3900 ;
      RECT 8.0920 14.2965 8.1180 15.3900 ;
      RECT 7.9840 14.2965 8.0100 15.3900 ;
      RECT 7.8760 14.2965 7.9020 15.3900 ;
      RECT 7.7680 14.2965 7.7940 15.3900 ;
      RECT 7.6600 14.2965 7.6860 15.3900 ;
      RECT 7.5520 14.2965 7.5780 15.3900 ;
      RECT 7.4440 14.2965 7.4700 15.3900 ;
      RECT 7.3360 14.2965 7.3620 15.3900 ;
      RECT 7.2280 14.2965 7.2540 15.3900 ;
      RECT 7.1200 14.2965 7.1460 15.3900 ;
      RECT 7.0120 14.2965 7.0380 15.3900 ;
      RECT 6.9040 14.2965 6.9300 15.3900 ;
      RECT 6.7960 14.2965 6.8220 15.3900 ;
      RECT 6.6880 14.2965 6.7140 15.3900 ;
      RECT 6.5800 14.2965 6.6060 15.3900 ;
      RECT 6.4720 14.2965 6.4980 15.3900 ;
      RECT 6.3640 14.2965 6.3900 15.3900 ;
      RECT 6.2560 14.2965 6.2820 15.3900 ;
      RECT 6.1480 14.2965 6.1740 15.3900 ;
      RECT 6.0400 14.2965 6.0660 15.3900 ;
      RECT 5.9320 14.2965 5.9580 15.3900 ;
      RECT 5.8240 14.2965 5.8500 15.3900 ;
      RECT 5.7160 14.2965 5.7420 15.3900 ;
      RECT 5.6080 14.2965 5.6340 15.3900 ;
      RECT 5.5000 14.2965 5.5260 15.3900 ;
      RECT 5.3920 14.2965 5.4180 15.3900 ;
      RECT 5.2840 14.2965 5.3100 15.3900 ;
      RECT 5.1760 14.2965 5.2020 15.3900 ;
      RECT 5.0680 14.2965 5.0940 15.3900 ;
      RECT 4.9600 14.2965 4.9860 15.3900 ;
      RECT 4.8520 14.2965 4.8780 15.3900 ;
      RECT 4.7440 14.2965 4.7700 15.3900 ;
      RECT 4.6360 14.2965 4.6620 15.3900 ;
      RECT 4.5280 14.2965 4.5540 15.3900 ;
      RECT 4.4200 14.2965 4.4460 15.3900 ;
      RECT 4.3120 14.2965 4.3380 15.3900 ;
      RECT 4.2040 14.2965 4.2300 15.3900 ;
      RECT 4.0960 14.2965 4.1220 15.3900 ;
      RECT 3.9880 14.2965 4.0140 15.3900 ;
      RECT 3.8800 14.2965 3.9060 15.3900 ;
      RECT 3.7720 14.2965 3.7980 15.3900 ;
      RECT 3.6640 14.2965 3.6900 15.3900 ;
      RECT 3.5560 14.2965 3.5820 15.3900 ;
      RECT 3.4480 14.2965 3.4740 15.3900 ;
      RECT 3.3400 14.2965 3.3660 15.3900 ;
      RECT 3.2320 14.2965 3.2580 15.3900 ;
      RECT 3.1240 14.2965 3.1500 15.3900 ;
      RECT 3.0160 14.2965 3.0420 15.3900 ;
      RECT 2.9080 14.2965 2.9340 15.3900 ;
      RECT 2.8000 14.2965 2.8260 15.3900 ;
      RECT 2.6920 14.2965 2.7180 15.3900 ;
      RECT 2.5840 14.2965 2.6100 15.3900 ;
      RECT 2.4760 14.2965 2.5020 15.3900 ;
      RECT 2.3680 14.2965 2.3940 15.3900 ;
      RECT 2.2600 14.2965 2.2860 15.3900 ;
      RECT 2.1520 14.2965 2.1780 15.3900 ;
      RECT 2.0440 14.2965 2.0700 15.3900 ;
      RECT 1.9360 14.2965 1.9620 15.3900 ;
      RECT 1.8280 14.2965 1.8540 15.3900 ;
      RECT 1.7200 14.2965 1.7460 15.3900 ;
      RECT 1.6120 14.2965 1.6380 15.3900 ;
      RECT 1.5040 14.2965 1.5300 15.3900 ;
      RECT 1.3960 14.2965 1.4220 15.3900 ;
      RECT 1.2880 14.2965 1.3140 15.3900 ;
      RECT 1.1800 14.2965 1.2060 15.3900 ;
      RECT 1.0720 14.2965 1.0980 15.3900 ;
      RECT 0.9640 14.2965 0.9900 15.3900 ;
      RECT 0.8560 14.2965 0.8820 15.3900 ;
      RECT 0.7480 14.2965 0.7740 15.3900 ;
      RECT 0.6400 14.2965 0.6660 15.3900 ;
      RECT 0.5320 14.2965 0.5580 15.3900 ;
      RECT 0.4240 14.2965 0.4500 15.3900 ;
      RECT 0.3160 14.2965 0.3420 15.3900 ;
      RECT 0.2080 14.2965 0.2340 15.3900 ;
      RECT 0.0050 14.2965 0.0900 15.3900 ;
      RECT 15.5530 15.3765 15.6810 16.4700 ;
      RECT 15.5390 16.0420 15.6810 16.3645 ;
      RECT 15.3190 15.7690 15.4530 16.4700 ;
      RECT 15.2960 16.1040 15.4530 16.3620 ;
      RECT 15.3190 15.3765 15.4170 16.4700 ;
      RECT 15.3190 15.4975 15.4310 15.7370 ;
      RECT 15.3190 15.3765 15.4530 15.4655 ;
      RECT 15.0940 15.8270 15.2280 16.4700 ;
      RECT 15.0940 15.3765 15.1920 16.4700 ;
      RECT 14.6770 15.3765 14.7600 16.4700 ;
      RECT 14.6770 15.4650 14.7740 16.4005 ;
      RECT 30.2680 15.3765 30.3530 16.4700 ;
      RECT 30.1240 15.3765 30.1500 16.4700 ;
      RECT 30.0160 15.3765 30.0420 16.4700 ;
      RECT 29.9080 15.3765 29.9340 16.4700 ;
      RECT 29.8000 15.3765 29.8260 16.4700 ;
      RECT 29.6920 15.3765 29.7180 16.4700 ;
      RECT 29.5840 15.3765 29.6100 16.4700 ;
      RECT 29.4760 15.3765 29.5020 16.4700 ;
      RECT 29.3680 15.3765 29.3940 16.4700 ;
      RECT 29.2600 15.3765 29.2860 16.4700 ;
      RECT 29.1520 15.3765 29.1780 16.4700 ;
      RECT 29.0440 15.3765 29.0700 16.4700 ;
      RECT 28.9360 15.3765 28.9620 16.4700 ;
      RECT 28.8280 15.3765 28.8540 16.4700 ;
      RECT 28.7200 15.3765 28.7460 16.4700 ;
      RECT 28.6120 15.3765 28.6380 16.4700 ;
      RECT 28.5040 15.3765 28.5300 16.4700 ;
      RECT 28.3960 15.3765 28.4220 16.4700 ;
      RECT 28.2880 15.3765 28.3140 16.4700 ;
      RECT 28.1800 15.3765 28.2060 16.4700 ;
      RECT 28.0720 15.3765 28.0980 16.4700 ;
      RECT 27.9640 15.3765 27.9900 16.4700 ;
      RECT 27.8560 15.3765 27.8820 16.4700 ;
      RECT 27.7480 15.3765 27.7740 16.4700 ;
      RECT 27.6400 15.3765 27.6660 16.4700 ;
      RECT 27.5320 15.3765 27.5580 16.4700 ;
      RECT 27.4240 15.3765 27.4500 16.4700 ;
      RECT 27.3160 15.3765 27.3420 16.4700 ;
      RECT 27.2080 15.3765 27.2340 16.4700 ;
      RECT 27.1000 15.3765 27.1260 16.4700 ;
      RECT 26.9920 15.3765 27.0180 16.4700 ;
      RECT 26.8840 15.3765 26.9100 16.4700 ;
      RECT 26.7760 15.3765 26.8020 16.4700 ;
      RECT 26.6680 15.3765 26.6940 16.4700 ;
      RECT 26.5600 15.3765 26.5860 16.4700 ;
      RECT 26.4520 15.3765 26.4780 16.4700 ;
      RECT 26.3440 15.3765 26.3700 16.4700 ;
      RECT 26.2360 15.3765 26.2620 16.4700 ;
      RECT 26.1280 15.3765 26.1540 16.4700 ;
      RECT 26.0200 15.3765 26.0460 16.4700 ;
      RECT 25.9120 15.3765 25.9380 16.4700 ;
      RECT 25.8040 15.3765 25.8300 16.4700 ;
      RECT 25.6960 15.3765 25.7220 16.4700 ;
      RECT 25.5880 15.3765 25.6140 16.4700 ;
      RECT 25.4800 15.3765 25.5060 16.4700 ;
      RECT 25.3720 15.3765 25.3980 16.4700 ;
      RECT 25.2640 15.3765 25.2900 16.4700 ;
      RECT 25.1560 15.3765 25.1820 16.4700 ;
      RECT 25.0480 15.3765 25.0740 16.4700 ;
      RECT 24.9400 15.3765 24.9660 16.4700 ;
      RECT 24.8320 15.3765 24.8580 16.4700 ;
      RECT 24.7240 15.3765 24.7500 16.4700 ;
      RECT 24.6160 15.3765 24.6420 16.4700 ;
      RECT 24.5080 15.3765 24.5340 16.4700 ;
      RECT 24.4000 15.3765 24.4260 16.4700 ;
      RECT 24.2920 15.3765 24.3180 16.4700 ;
      RECT 24.1840 15.3765 24.2100 16.4700 ;
      RECT 24.0760 15.3765 24.1020 16.4700 ;
      RECT 23.9680 15.3765 23.9940 16.4700 ;
      RECT 23.8600 15.3765 23.8860 16.4700 ;
      RECT 23.7520 15.3765 23.7780 16.4700 ;
      RECT 23.6440 15.3765 23.6700 16.4700 ;
      RECT 23.5360 15.3765 23.5620 16.4700 ;
      RECT 23.4280 15.3765 23.4540 16.4700 ;
      RECT 23.3200 15.3765 23.3460 16.4700 ;
      RECT 23.2120 15.3765 23.2380 16.4700 ;
      RECT 23.1040 15.3765 23.1300 16.4700 ;
      RECT 22.9960 15.3765 23.0220 16.4700 ;
      RECT 22.8880 15.3765 22.9140 16.4700 ;
      RECT 22.7800 15.3765 22.8060 16.4700 ;
      RECT 22.6720 15.3765 22.6980 16.4700 ;
      RECT 22.5640 15.3765 22.5900 16.4700 ;
      RECT 22.4560 15.3765 22.4820 16.4700 ;
      RECT 22.3480 15.3765 22.3740 16.4700 ;
      RECT 22.2400 15.3765 22.2660 16.4700 ;
      RECT 22.1320 15.3765 22.1580 16.4700 ;
      RECT 22.0240 15.3765 22.0500 16.4700 ;
      RECT 21.9160 15.3765 21.9420 16.4700 ;
      RECT 21.8080 15.3765 21.8340 16.4700 ;
      RECT 21.7000 15.3765 21.7260 16.4700 ;
      RECT 21.5920 15.3765 21.6180 16.4700 ;
      RECT 21.4840 15.3765 21.5100 16.4700 ;
      RECT 21.3760 15.3765 21.4020 16.4700 ;
      RECT 21.2680 15.3765 21.2940 16.4700 ;
      RECT 21.1600 15.3765 21.1860 16.4700 ;
      RECT 21.0520 15.3765 21.0780 16.4700 ;
      RECT 20.9440 15.3765 20.9700 16.4700 ;
      RECT 20.8360 15.3765 20.8620 16.4700 ;
      RECT 20.7280 15.3765 20.7540 16.4700 ;
      RECT 20.6200 15.3765 20.6460 16.4700 ;
      RECT 20.5120 15.3765 20.5380 16.4700 ;
      RECT 20.4040 15.3765 20.4300 16.4700 ;
      RECT 20.2960 15.3765 20.3220 16.4700 ;
      RECT 20.1880 15.3765 20.2140 16.4700 ;
      RECT 20.0800 15.3765 20.1060 16.4700 ;
      RECT 19.9720 15.3765 19.9980 16.4700 ;
      RECT 19.8640 15.3765 19.8900 16.4700 ;
      RECT 19.7560 15.3765 19.7820 16.4700 ;
      RECT 19.6480 15.3765 19.6740 16.4700 ;
      RECT 19.5400 15.3765 19.5660 16.4700 ;
      RECT 19.4320 15.3765 19.4580 16.4700 ;
      RECT 19.3240 15.3765 19.3500 16.4700 ;
      RECT 19.2160 15.3765 19.2420 16.4700 ;
      RECT 19.1080 15.3765 19.1340 16.4700 ;
      RECT 19.0000 15.3765 19.0260 16.4700 ;
      RECT 18.8920 15.3765 18.9180 16.4700 ;
      RECT 18.7840 15.3765 18.8100 16.4700 ;
      RECT 18.6760 15.3765 18.7020 16.4700 ;
      RECT 18.5680 15.3765 18.5940 16.4700 ;
      RECT 18.4600 15.3765 18.4860 16.4700 ;
      RECT 18.3520 15.3765 18.3780 16.4700 ;
      RECT 18.2440 15.3765 18.2700 16.4700 ;
      RECT 18.1360 15.3765 18.1620 16.4700 ;
      RECT 18.0280 15.3765 18.0540 16.4700 ;
      RECT 17.9200 15.3765 17.9460 16.4700 ;
      RECT 17.8120 15.3765 17.8380 16.4700 ;
      RECT 17.7040 15.3765 17.7300 16.4700 ;
      RECT 17.5960 15.3765 17.6220 16.4700 ;
      RECT 17.4880 15.3765 17.5140 16.4700 ;
      RECT 17.3800 15.3765 17.4060 16.4700 ;
      RECT 17.2720 15.3765 17.2980 16.4700 ;
      RECT 17.1640 15.3765 17.1900 16.4700 ;
      RECT 17.0560 15.3765 17.0820 16.4700 ;
      RECT 16.9480 15.3765 16.9740 16.4700 ;
      RECT 16.8400 15.3765 16.8660 16.4700 ;
      RECT 16.7320 15.3765 16.7580 16.4700 ;
      RECT 16.6240 15.3765 16.6500 16.4700 ;
      RECT 16.5160 15.3765 16.5420 16.4700 ;
      RECT 16.4080 15.3765 16.4340 16.4700 ;
      RECT 16.3000 15.3765 16.3260 16.4700 ;
      RECT 16.0870 15.3765 16.1640 16.4700 ;
      RECT 14.1940 15.3765 14.2710 16.4700 ;
      RECT 14.0320 15.3765 14.0580 16.4700 ;
      RECT 13.9240 15.3765 13.9500 16.4700 ;
      RECT 13.8160 15.3765 13.8420 16.4700 ;
      RECT 13.7080 15.3765 13.7340 16.4700 ;
      RECT 13.6000 15.3765 13.6260 16.4700 ;
      RECT 13.4920 15.3765 13.5180 16.4700 ;
      RECT 13.3840 15.3765 13.4100 16.4700 ;
      RECT 13.2760 15.3765 13.3020 16.4700 ;
      RECT 13.1680 15.3765 13.1940 16.4700 ;
      RECT 13.0600 15.3765 13.0860 16.4700 ;
      RECT 12.9520 15.3765 12.9780 16.4700 ;
      RECT 12.8440 15.3765 12.8700 16.4700 ;
      RECT 12.7360 15.3765 12.7620 16.4700 ;
      RECT 12.6280 15.3765 12.6540 16.4700 ;
      RECT 12.5200 15.3765 12.5460 16.4700 ;
      RECT 12.4120 15.3765 12.4380 16.4700 ;
      RECT 12.3040 15.3765 12.3300 16.4700 ;
      RECT 12.1960 15.3765 12.2220 16.4700 ;
      RECT 12.0880 15.3765 12.1140 16.4700 ;
      RECT 11.9800 15.3765 12.0060 16.4700 ;
      RECT 11.8720 15.3765 11.8980 16.4700 ;
      RECT 11.7640 15.3765 11.7900 16.4700 ;
      RECT 11.6560 15.3765 11.6820 16.4700 ;
      RECT 11.5480 15.3765 11.5740 16.4700 ;
      RECT 11.4400 15.3765 11.4660 16.4700 ;
      RECT 11.3320 15.3765 11.3580 16.4700 ;
      RECT 11.2240 15.3765 11.2500 16.4700 ;
      RECT 11.1160 15.3765 11.1420 16.4700 ;
      RECT 11.0080 15.3765 11.0340 16.4700 ;
      RECT 10.9000 15.3765 10.9260 16.4700 ;
      RECT 10.7920 15.3765 10.8180 16.4700 ;
      RECT 10.6840 15.3765 10.7100 16.4700 ;
      RECT 10.5760 15.3765 10.6020 16.4700 ;
      RECT 10.4680 15.3765 10.4940 16.4700 ;
      RECT 10.3600 15.3765 10.3860 16.4700 ;
      RECT 10.2520 15.3765 10.2780 16.4700 ;
      RECT 10.1440 15.3765 10.1700 16.4700 ;
      RECT 10.0360 15.3765 10.0620 16.4700 ;
      RECT 9.9280 15.3765 9.9540 16.4700 ;
      RECT 9.8200 15.3765 9.8460 16.4700 ;
      RECT 9.7120 15.3765 9.7380 16.4700 ;
      RECT 9.6040 15.3765 9.6300 16.4700 ;
      RECT 9.4960 15.3765 9.5220 16.4700 ;
      RECT 9.3880 15.3765 9.4140 16.4700 ;
      RECT 9.2800 15.3765 9.3060 16.4700 ;
      RECT 9.1720 15.3765 9.1980 16.4700 ;
      RECT 9.0640 15.3765 9.0900 16.4700 ;
      RECT 8.9560 15.3765 8.9820 16.4700 ;
      RECT 8.8480 15.3765 8.8740 16.4700 ;
      RECT 8.7400 15.3765 8.7660 16.4700 ;
      RECT 8.6320 15.3765 8.6580 16.4700 ;
      RECT 8.5240 15.3765 8.5500 16.4700 ;
      RECT 8.4160 15.3765 8.4420 16.4700 ;
      RECT 8.3080 15.3765 8.3340 16.4700 ;
      RECT 8.2000 15.3765 8.2260 16.4700 ;
      RECT 8.0920 15.3765 8.1180 16.4700 ;
      RECT 7.9840 15.3765 8.0100 16.4700 ;
      RECT 7.8760 15.3765 7.9020 16.4700 ;
      RECT 7.7680 15.3765 7.7940 16.4700 ;
      RECT 7.6600 15.3765 7.6860 16.4700 ;
      RECT 7.5520 15.3765 7.5780 16.4700 ;
      RECT 7.4440 15.3765 7.4700 16.4700 ;
      RECT 7.3360 15.3765 7.3620 16.4700 ;
      RECT 7.2280 15.3765 7.2540 16.4700 ;
      RECT 7.1200 15.3765 7.1460 16.4700 ;
      RECT 7.0120 15.3765 7.0380 16.4700 ;
      RECT 6.9040 15.3765 6.9300 16.4700 ;
      RECT 6.7960 15.3765 6.8220 16.4700 ;
      RECT 6.6880 15.3765 6.7140 16.4700 ;
      RECT 6.5800 15.3765 6.6060 16.4700 ;
      RECT 6.4720 15.3765 6.4980 16.4700 ;
      RECT 6.3640 15.3765 6.3900 16.4700 ;
      RECT 6.2560 15.3765 6.2820 16.4700 ;
      RECT 6.1480 15.3765 6.1740 16.4700 ;
      RECT 6.0400 15.3765 6.0660 16.4700 ;
      RECT 5.9320 15.3765 5.9580 16.4700 ;
      RECT 5.8240 15.3765 5.8500 16.4700 ;
      RECT 5.7160 15.3765 5.7420 16.4700 ;
      RECT 5.6080 15.3765 5.6340 16.4700 ;
      RECT 5.5000 15.3765 5.5260 16.4700 ;
      RECT 5.3920 15.3765 5.4180 16.4700 ;
      RECT 5.2840 15.3765 5.3100 16.4700 ;
      RECT 5.1760 15.3765 5.2020 16.4700 ;
      RECT 5.0680 15.3765 5.0940 16.4700 ;
      RECT 4.9600 15.3765 4.9860 16.4700 ;
      RECT 4.8520 15.3765 4.8780 16.4700 ;
      RECT 4.7440 15.3765 4.7700 16.4700 ;
      RECT 4.6360 15.3765 4.6620 16.4700 ;
      RECT 4.5280 15.3765 4.5540 16.4700 ;
      RECT 4.4200 15.3765 4.4460 16.4700 ;
      RECT 4.3120 15.3765 4.3380 16.4700 ;
      RECT 4.2040 15.3765 4.2300 16.4700 ;
      RECT 4.0960 15.3765 4.1220 16.4700 ;
      RECT 3.9880 15.3765 4.0140 16.4700 ;
      RECT 3.8800 15.3765 3.9060 16.4700 ;
      RECT 3.7720 15.3765 3.7980 16.4700 ;
      RECT 3.6640 15.3765 3.6900 16.4700 ;
      RECT 3.5560 15.3765 3.5820 16.4700 ;
      RECT 3.4480 15.3765 3.4740 16.4700 ;
      RECT 3.3400 15.3765 3.3660 16.4700 ;
      RECT 3.2320 15.3765 3.2580 16.4700 ;
      RECT 3.1240 15.3765 3.1500 16.4700 ;
      RECT 3.0160 15.3765 3.0420 16.4700 ;
      RECT 2.9080 15.3765 2.9340 16.4700 ;
      RECT 2.8000 15.3765 2.8260 16.4700 ;
      RECT 2.6920 15.3765 2.7180 16.4700 ;
      RECT 2.5840 15.3765 2.6100 16.4700 ;
      RECT 2.4760 15.3765 2.5020 16.4700 ;
      RECT 2.3680 15.3765 2.3940 16.4700 ;
      RECT 2.2600 15.3765 2.2860 16.4700 ;
      RECT 2.1520 15.3765 2.1780 16.4700 ;
      RECT 2.0440 15.3765 2.0700 16.4700 ;
      RECT 1.9360 15.3765 1.9620 16.4700 ;
      RECT 1.8280 15.3765 1.8540 16.4700 ;
      RECT 1.7200 15.3765 1.7460 16.4700 ;
      RECT 1.6120 15.3765 1.6380 16.4700 ;
      RECT 1.5040 15.3765 1.5300 16.4700 ;
      RECT 1.3960 15.3765 1.4220 16.4700 ;
      RECT 1.2880 15.3765 1.3140 16.4700 ;
      RECT 1.1800 15.3765 1.2060 16.4700 ;
      RECT 1.0720 15.3765 1.0980 16.4700 ;
      RECT 0.9640 15.3765 0.9900 16.4700 ;
      RECT 0.8560 15.3765 0.8820 16.4700 ;
      RECT 0.7480 15.3765 0.7740 16.4700 ;
      RECT 0.6400 15.3765 0.6660 16.4700 ;
      RECT 0.5320 15.3765 0.5580 16.4700 ;
      RECT 0.4240 15.3765 0.4500 16.4700 ;
      RECT 0.3160 15.3765 0.3420 16.4700 ;
      RECT 0.2080 15.3765 0.2340 16.4700 ;
      RECT 0.0050 15.3765 0.0900 16.4700 ;
      RECT 15.5530 16.4565 15.6810 17.5500 ;
      RECT 15.5390 17.1220 15.6810 17.4445 ;
      RECT 15.3190 16.8490 15.4530 17.5500 ;
      RECT 15.2960 17.1840 15.4530 17.4420 ;
      RECT 15.3190 16.4565 15.4170 17.5500 ;
      RECT 15.3190 16.5775 15.4310 16.8170 ;
      RECT 15.3190 16.4565 15.4530 16.5455 ;
      RECT 15.0940 16.9070 15.2280 17.5500 ;
      RECT 15.0940 16.4565 15.1920 17.5500 ;
      RECT 14.6770 16.4565 14.7600 17.5500 ;
      RECT 14.6770 16.5450 14.7740 17.4805 ;
      RECT 30.2680 16.4565 30.3530 17.5500 ;
      RECT 30.1240 16.4565 30.1500 17.5500 ;
      RECT 30.0160 16.4565 30.0420 17.5500 ;
      RECT 29.9080 16.4565 29.9340 17.5500 ;
      RECT 29.8000 16.4565 29.8260 17.5500 ;
      RECT 29.6920 16.4565 29.7180 17.5500 ;
      RECT 29.5840 16.4565 29.6100 17.5500 ;
      RECT 29.4760 16.4565 29.5020 17.5500 ;
      RECT 29.3680 16.4565 29.3940 17.5500 ;
      RECT 29.2600 16.4565 29.2860 17.5500 ;
      RECT 29.1520 16.4565 29.1780 17.5500 ;
      RECT 29.0440 16.4565 29.0700 17.5500 ;
      RECT 28.9360 16.4565 28.9620 17.5500 ;
      RECT 28.8280 16.4565 28.8540 17.5500 ;
      RECT 28.7200 16.4565 28.7460 17.5500 ;
      RECT 28.6120 16.4565 28.6380 17.5500 ;
      RECT 28.5040 16.4565 28.5300 17.5500 ;
      RECT 28.3960 16.4565 28.4220 17.5500 ;
      RECT 28.2880 16.4565 28.3140 17.5500 ;
      RECT 28.1800 16.4565 28.2060 17.5500 ;
      RECT 28.0720 16.4565 28.0980 17.5500 ;
      RECT 27.9640 16.4565 27.9900 17.5500 ;
      RECT 27.8560 16.4565 27.8820 17.5500 ;
      RECT 27.7480 16.4565 27.7740 17.5500 ;
      RECT 27.6400 16.4565 27.6660 17.5500 ;
      RECT 27.5320 16.4565 27.5580 17.5500 ;
      RECT 27.4240 16.4565 27.4500 17.5500 ;
      RECT 27.3160 16.4565 27.3420 17.5500 ;
      RECT 27.2080 16.4565 27.2340 17.5500 ;
      RECT 27.1000 16.4565 27.1260 17.5500 ;
      RECT 26.9920 16.4565 27.0180 17.5500 ;
      RECT 26.8840 16.4565 26.9100 17.5500 ;
      RECT 26.7760 16.4565 26.8020 17.5500 ;
      RECT 26.6680 16.4565 26.6940 17.5500 ;
      RECT 26.5600 16.4565 26.5860 17.5500 ;
      RECT 26.4520 16.4565 26.4780 17.5500 ;
      RECT 26.3440 16.4565 26.3700 17.5500 ;
      RECT 26.2360 16.4565 26.2620 17.5500 ;
      RECT 26.1280 16.4565 26.1540 17.5500 ;
      RECT 26.0200 16.4565 26.0460 17.5500 ;
      RECT 25.9120 16.4565 25.9380 17.5500 ;
      RECT 25.8040 16.4565 25.8300 17.5500 ;
      RECT 25.6960 16.4565 25.7220 17.5500 ;
      RECT 25.5880 16.4565 25.6140 17.5500 ;
      RECT 25.4800 16.4565 25.5060 17.5500 ;
      RECT 25.3720 16.4565 25.3980 17.5500 ;
      RECT 25.2640 16.4565 25.2900 17.5500 ;
      RECT 25.1560 16.4565 25.1820 17.5500 ;
      RECT 25.0480 16.4565 25.0740 17.5500 ;
      RECT 24.9400 16.4565 24.9660 17.5500 ;
      RECT 24.8320 16.4565 24.8580 17.5500 ;
      RECT 24.7240 16.4565 24.7500 17.5500 ;
      RECT 24.6160 16.4565 24.6420 17.5500 ;
      RECT 24.5080 16.4565 24.5340 17.5500 ;
      RECT 24.4000 16.4565 24.4260 17.5500 ;
      RECT 24.2920 16.4565 24.3180 17.5500 ;
      RECT 24.1840 16.4565 24.2100 17.5500 ;
      RECT 24.0760 16.4565 24.1020 17.5500 ;
      RECT 23.9680 16.4565 23.9940 17.5500 ;
      RECT 23.8600 16.4565 23.8860 17.5500 ;
      RECT 23.7520 16.4565 23.7780 17.5500 ;
      RECT 23.6440 16.4565 23.6700 17.5500 ;
      RECT 23.5360 16.4565 23.5620 17.5500 ;
      RECT 23.4280 16.4565 23.4540 17.5500 ;
      RECT 23.3200 16.4565 23.3460 17.5500 ;
      RECT 23.2120 16.4565 23.2380 17.5500 ;
      RECT 23.1040 16.4565 23.1300 17.5500 ;
      RECT 22.9960 16.4565 23.0220 17.5500 ;
      RECT 22.8880 16.4565 22.9140 17.5500 ;
      RECT 22.7800 16.4565 22.8060 17.5500 ;
      RECT 22.6720 16.4565 22.6980 17.5500 ;
      RECT 22.5640 16.4565 22.5900 17.5500 ;
      RECT 22.4560 16.4565 22.4820 17.5500 ;
      RECT 22.3480 16.4565 22.3740 17.5500 ;
      RECT 22.2400 16.4565 22.2660 17.5500 ;
      RECT 22.1320 16.4565 22.1580 17.5500 ;
      RECT 22.0240 16.4565 22.0500 17.5500 ;
      RECT 21.9160 16.4565 21.9420 17.5500 ;
      RECT 21.8080 16.4565 21.8340 17.5500 ;
      RECT 21.7000 16.4565 21.7260 17.5500 ;
      RECT 21.5920 16.4565 21.6180 17.5500 ;
      RECT 21.4840 16.4565 21.5100 17.5500 ;
      RECT 21.3760 16.4565 21.4020 17.5500 ;
      RECT 21.2680 16.4565 21.2940 17.5500 ;
      RECT 21.1600 16.4565 21.1860 17.5500 ;
      RECT 21.0520 16.4565 21.0780 17.5500 ;
      RECT 20.9440 16.4565 20.9700 17.5500 ;
      RECT 20.8360 16.4565 20.8620 17.5500 ;
      RECT 20.7280 16.4565 20.7540 17.5500 ;
      RECT 20.6200 16.4565 20.6460 17.5500 ;
      RECT 20.5120 16.4565 20.5380 17.5500 ;
      RECT 20.4040 16.4565 20.4300 17.5500 ;
      RECT 20.2960 16.4565 20.3220 17.5500 ;
      RECT 20.1880 16.4565 20.2140 17.5500 ;
      RECT 20.0800 16.4565 20.1060 17.5500 ;
      RECT 19.9720 16.4565 19.9980 17.5500 ;
      RECT 19.8640 16.4565 19.8900 17.5500 ;
      RECT 19.7560 16.4565 19.7820 17.5500 ;
      RECT 19.6480 16.4565 19.6740 17.5500 ;
      RECT 19.5400 16.4565 19.5660 17.5500 ;
      RECT 19.4320 16.4565 19.4580 17.5500 ;
      RECT 19.3240 16.4565 19.3500 17.5500 ;
      RECT 19.2160 16.4565 19.2420 17.5500 ;
      RECT 19.1080 16.4565 19.1340 17.5500 ;
      RECT 19.0000 16.4565 19.0260 17.5500 ;
      RECT 18.8920 16.4565 18.9180 17.5500 ;
      RECT 18.7840 16.4565 18.8100 17.5500 ;
      RECT 18.6760 16.4565 18.7020 17.5500 ;
      RECT 18.5680 16.4565 18.5940 17.5500 ;
      RECT 18.4600 16.4565 18.4860 17.5500 ;
      RECT 18.3520 16.4565 18.3780 17.5500 ;
      RECT 18.2440 16.4565 18.2700 17.5500 ;
      RECT 18.1360 16.4565 18.1620 17.5500 ;
      RECT 18.0280 16.4565 18.0540 17.5500 ;
      RECT 17.9200 16.4565 17.9460 17.5500 ;
      RECT 17.8120 16.4565 17.8380 17.5500 ;
      RECT 17.7040 16.4565 17.7300 17.5500 ;
      RECT 17.5960 16.4565 17.6220 17.5500 ;
      RECT 17.4880 16.4565 17.5140 17.5500 ;
      RECT 17.3800 16.4565 17.4060 17.5500 ;
      RECT 17.2720 16.4565 17.2980 17.5500 ;
      RECT 17.1640 16.4565 17.1900 17.5500 ;
      RECT 17.0560 16.4565 17.0820 17.5500 ;
      RECT 16.9480 16.4565 16.9740 17.5500 ;
      RECT 16.8400 16.4565 16.8660 17.5500 ;
      RECT 16.7320 16.4565 16.7580 17.5500 ;
      RECT 16.6240 16.4565 16.6500 17.5500 ;
      RECT 16.5160 16.4565 16.5420 17.5500 ;
      RECT 16.4080 16.4565 16.4340 17.5500 ;
      RECT 16.3000 16.4565 16.3260 17.5500 ;
      RECT 16.0870 16.4565 16.1640 17.5500 ;
      RECT 14.1940 16.4565 14.2710 17.5500 ;
      RECT 14.0320 16.4565 14.0580 17.5500 ;
      RECT 13.9240 16.4565 13.9500 17.5500 ;
      RECT 13.8160 16.4565 13.8420 17.5500 ;
      RECT 13.7080 16.4565 13.7340 17.5500 ;
      RECT 13.6000 16.4565 13.6260 17.5500 ;
      RECT 13.4920 16.4565 13.5180 17.5500 ;
      RECT 13.3840 16.4565 13.4100 17.5500 ;
      RECT 13.2760 16.4565 13.3020 17.5500 ;
      RECT 13.1680 16.4565 13.1940 17.5500 ;
      RECT 13.0600 16.4565 13.0860 17.5500 ;
      RECT 12.9520 16.4565 12.9780 17.5500 ;
      RECT 12.8440 16.4565 12.8700 17.5500 ;
      RECT 12.7360 16.4565 12.7620 17.5500 ;
      RECT 12.6280 16.4565 12.6540 17.5500 ;
      RECT 12.5200 16.4565 12.5460 17.5500 ;
      RECT 12.4120 16.4565 12.4380 17.5500 ;
      RECT 12.3040 16.4565 12.3300 17.5500 ;
      RECT 12.1960 16.4565 12.2220 17.5500 ;
      RECT 12.0880 16.4565 12.1140 17.5500 ;
      RECT 11.9800 16.4565 12.0060 17.5500 ;
      RECT 11.8720 16.4565 11.8980 17.5500 ;
      RECT 11.7640 16.4565 11.7900 17.5500 ;
      RECT 11.6560 16.4565 11.6820 17.5500 ;
      RECT 11.5480 16.4565 11.5740 17.5500 ;
      RECT 11.4400 16.4565 11.4660 17.5500 ;
      RECT 11.3320 16.4565 11.3580 17.5500 ;
      RECT 11.2240 16.4565 11.2500 17.5500 ;
      RECT 11.1160 16.4565 11.1420 17.5500 ;
      RECT 11.0080 16.4565 11.0340 17.5500 ;
      RECT 10.9000 16.4565 10.9260 17.5500 ;
      RECT 10.7920 16.4565 10.8180 17.5500 ;
      RECT 10.6840 16.4565 10.7100 17.5500 ;
      RECT 10.5760 16.4565 10.6020 17.5500 ;
      RECT 10.4680 16.4565 10.4940 17.5500 ;
      RECT 10.3600 16.4565 10.3860 17.5500 ;
      RECT 10.2520 16.4565 10.2780 17.5500 ;
      RECT 10.1440 16.4565 10.1700 17.5500 ;
      RECT 10.0360 16.4565 10.0620 17.5500 ;
      RECT 9.9280 16.4565 9.9540 17.5500 ;
      RECT 9.8200 16.4565 9.8460 17.5500 ;
      RECT 9.7120 16.4565 9.7380 17.5500 ;
      RECT 9.6040 16.4565 9.6300 17.5500 ;
      RECT 9.4960 16.4565 9.5220 17.5500 ;
      RECT 9.3880 16.4565 9.4140 17.5500 ;
      RECT 9.2800 16.4565 9.3060 17.5500 ;
      RECT 9.1720 16.4565 9.1980 17.5500 ;
      RECT 9.0640 16.4565 9.0900 17.5500 ;
      RECT 8.9560 16.4565 8.9820 17.5500 ;
      RECT 8.8480 16.4565 8.8740 17.5500 ;
      RECT 8.7400 16.4565 8.7660 17.5500 ;
      RECT 8.6320 16.4565 8.6580 17.5500 ;
      RECT 8.5240 16.4565 8.5500 17.5500 ;
      RECT 8.4160 16.4565 8.4420 17.5500 ;
      RECT 8.3080 16.4565 8.3340 17.5500 ;
      RECT 8.2000 16.4565 8.2260 17.5500 ;
      RECT 8.0920 16.4565 8.1180 17.5500 ;
      RECT 7.9840 16.4565 8.0100 17.5500 ;
      RECT 7.8760 16.4565 7.9020 17.5500 ;
      RECT 7.7680 16.4565 7.7940 17.5500 ;
      RECT 7.6600 16.4565 7.6860 17.5500 ;
      RECT 7.5520 16.4565 7.5780 17.5500 ;
      RECT 7.4440 16.4565 7.4700 17.5500 ;
      RECT 7.3360 16.4565 7.3620 17.5500 ;
      RECT 7.2280 16.4565 7.2540 17.5500 ;
      RECT 7.1200 16.4565 7.1460 17.5500 ;
      RECT 7.0120 16.4565 7.0380 17.5500 ;
      RECT 6.9040 16.4565 6.9300 17.5500 ;
      RECT 6.7960 16.4565 6.8220 17.5500 ;
      RECT 6.6880 16.4565 6.7140 17.5500 ;
      RECT 6.5800 16.4565 6.6060 17.5500 ;
      RECT 6.4720 16.4565 6.4980 17.5500 ;
      RECT 6.3640 16.4565 6.3900 17.5500 ;
      RECT 6.2560 16.4565 6.2820 17.5500 ;
      RECT 6.1480 16.4565 6.1740 17.5500 ;
      RECT 6.0400 16.4565 6.0660 17.5500 ;
      RECT 5.9320 16.4565 5.9580 17.5500 ;
      RECT 5.8240 16.4565 5.8500 17.5500 ;
      RECT 5.7160 16.4565 5.7420 17.5500 ;
      RECT 5.6080 16.4565 5.6340 17.5500 ;
      RECT 5.5000 16.4565 5.5260 17.5500 ;
      RECT 5.3920 16.4565 5.4180 17.5500 ;
      RECT 5.2840 16.4565 5.3100 17.5500 ;
      RECT 5.1760 16.4565 5.2020 17.5500 ;
      RECT 5.0680 16.4565 5.0940 17.5500 ;
      RECT 4.9600 16.4565 4.9860 17.5500 ;
      RECT 4.8520 16.4565 4.8780 17.5500 ;
      RECT 4.7440 16.4565 4.7700 17.5500 ;
      RECT 4.6360 16.4565 4.6620 17.5500 ;
      RECT 4.5280 16.4565 4.5540 17.5500 ;
      RECT 4.4200 16.4565 4.4460 17.5500 ;
      RECT 4.3120 16.4565 4.3380 17.5500 ;
      RECT 4.2040 16.4565 4.2300 17.5500 ;
      RECT 4.0960 16.4565 4.1220 17.5500 ;
      RECT 3.9880 16.4565 4.0140 17.5500 ;
      RECT 3.8800 16.4565 3.9060 17.5500 ;
      RECT 3.7720 16.4565 3.7980 17.5500 ;
      RECT 3.6640 16.4565 3.6900 17.5500 ;
      RECT 3.5560 16.4565 3.5820 17.5500 ;
      RECT 3.4480 16.4565 3.4740 17.5500 ;
      RECT 3.3400 16.4565 3.3660 17.5500 ;
      RECT 3.2320 16.4565 3.2580 17.5500 ;
      RECT 3.1240 16.4565 3.1500 17.5500 ;
      RECT 3.0160 16.4565 3.0420 17.5500 ;
      RECT 2.9080 16.4565 2.9340 17.5500 ;
      RECT 2.8000 16.4565 2.8260 17.5500 ;
      RECT 2.6920 16.4565 2.7180 17.5500 ;
      RECT 2.5840 16.4565 2.6100 17.5500 ;
      RECT 2.4760 16.4565 2.5020 17.5500 ;
      RECT 2.3680 16.4565 2.3940 17.5500 ;
      RECT 2.2600 16.4565 2.2860 17.5500 ;
      RECT 2.1520 16.4565 2.1780 17.5500 ;
      RECT 2.0440 16.4565 2.0700 17.5500 ;
      RECT 1.9360 16.4565 1.9620 17.5500 ;
      RECT 1.8280 16.4565 1.8540 17.5500 ;
      RECT 1.7200 16.4565 1.7460 17.5500 ;
      RECT 1.6120 16.4565 1.6380 17.5500 ;
      RECT 1.5040 16.4565 1.5300 17.5500 ;
      RECT 1.3960 16.4565 1.4220 17.5500 ;
      RECT 1.2880 16.4565 1.3140 17.5500 ;
      RECT 1.1800 16.4565 1.2060 17.5500 ;
      RECT 1.0720 16.4565 1.0980 17.5500 ;
      RECT 0.9640 16.4565 0.9900 17.5500 ;
      RECT 0.8560 16.4565 0.8820 17.5500 ;
      RECT 0.7480 16.4565 0.7740 17.5500 ;
      RECT 0.6400 16.4565 0.6660 17.5500 ;
      RECT 0.5320 16.4565 0.5580 17.5500 ;
      RECT 0.4240 16.4565 0.4500 17.5500 ;
      RECT 0.3160 16.4565 0.3420 17.5500 ;
      RECT 0.2080 16.4565 0.2340 17.5500 ;
      RECT 0.0050 16.4565 0.0900 17.5500 ;
      RECT 15.5530 17.5365 15.6810 18.6300 ;
      RECT 15.5390 18.2020 15.6810 18.5245 ;
      RECT 15.3190 17.9290 15.4530 18.6300 ;
      RECT 15.2960 18.2640 15.4530 18.5220 ;
      RECT 15.3190 17.5365 15.4170 18.6300 ;
      RECT 15.3190 17.6575 15.4310 17.8970 ;
      RECT 15.3190 17.5365 15.4530 17.6255 ;
      RECT 15.0940 17.9870 15.2280 18.6300 ;
      RECT 15.0940 17.5365 15.1920 18.6300 ;
      RECT 14.6770 17.5365 14.7600 18.6300 ;
      RECT 14.6770 17.6250 14.7740 18.5605 ;
      RECT 30.2680 17.5365 30.3530 18.6300 ;
      RECT 30.1240 17.5365 30.1500 18.6300 ;
      RECT 30.0160 17.5365 30.0420 18.6300 ;
      RECT 29.9080 17.5365 29.9340 18.6300 ;
      RECT 29.8000 17.5365 29.8260 18.6300 ;
      RECT 29.6920 17.5365 29.7180 18.6300 ;
      RECT 29.5840 17.5365 29.6100 18.6300 ;
      RECT 29.4760 17.5365 29.5020 18.6300 ;
      RECT 29.3680 17.5365 29.3940 18.6300 ;
      RECT 29.2600 17.5365 29.2860 18.6300 ;
      RECT 29.1520 17.5365 29.1780 18.6300 ;
      RECT 29.0440 17.5365 29.0700 18.6300 ;
      RECT 28.9360 17.5365 28.9620 18.6300 ;
      RECT 28.8280 17.5365 28.8540 18.6300 ;
      RECT 28.7200 17.5365 28.7460 18.6300 ;
      RECT 28.6120 17.5365 28.6380 18.6300 ;
      RECT 28.5040 17.5365 28.5300 18.6300 ;
      RECT 28.3960 17.5365 28.4220 18.6300 ;
      RECT 28.2880 17.5365 28.3140 18.6300 ;
      RECT 28.1800 17.5365 28.2060 18.6300 ;
      RECT 28.0720 17.5365 28.0980 18.6300 ;
      RECT 27.9640 17.5365 27.9900 18.6300 ;
      RECT 27.8560 17.5365 27.8820 18.6300 ;
      RECT 27.7480 17.5365 27.7740 18.6300 ;
      RECT 27.6400 17.5365 27.6660 18.6300 ;
      RECT 27.5320 17.5365 27.5580 18.6300 ;
      RECT 27.4240 17.5365 27.4500 18.6300 ;
      RECT 27.3160 17.5365 27.3420 18.6300 ;
      RECT 27.2080 17.5365 27.2340 18.6300 ;
      RECT 27.1000 17.5365 27.1260 18.6300 ;
      RECT 26.9920 17.5365 27.0180 18.6300 ;
      RECT 26.8840 17.5365 26.9100 18.6300 ;
      RECT 26.7760 17.5365 26.8020 18.6300 ;
      RECT 26.6680 17.5365 26.6940 18.6300 ;
      RECT 26.5600 17.5365 26.5860 18.6300 ;
      RECT 26.4520 17.5365 26.4780 18.6300 ;
      RECT 26.3440 17.5365 26.3700 18.6300 ;
      RECT 26.2360 17.5365 26.2620 18.6300 ;
      RECT 26.1280 17.5365 26.1540 18.6300 ;
      RECT 26.0200 17.5365 26.0460 18.6300 ;
      RECT 25.9120 17.5365 25.9380 18.6300 ;
      RECT 25.8040 17.5365 25.8300 18.6300 ;
      RECT 25.6960 17.5365 25.7220 18.6300 ;
      RECT 25.5880 17.5365 25.6140 18.6300 ;
      RECT 25.4800 17.5365 25.5060 18.6300 ;
      RECT 25.3720 17.5365 25.3980 18.6300 ;
      RECT 25.2640 17.5365 25.2900 18.6300 ;
      RECT 25.1560 17.5365 25.1820 18.6300 ;
      RECT 25.0480 17.5365 25.0740 18.6300 ;
      RECT 24.9400 17.5365 24.9660 18.6300 ;
      RECT 24.8320 17.5365 24.8580 18.6300 ;
      RECT 24.7240 17.5365 24.7500 18.6300 ;
      RECT 24.6160 17.5365 24.6420 18.6300 ;
      RECT 24.5080 17.5365 24.5340 18.6300 ;
      RECT 24.4000 17.5365 24.4260 18.6300 ;
      RECT 24.2920 17.5365 24.3180 18.6300 ;
      RECT 24.1840 17.5365 24.2100 18.6300 ;
      RECT 24.0760 17.5365 24.1020 18.6300 ;
      RECT 23.9680 17.5365 23.9940 18.6300 ;
      RECT 23.8600 17.5365 23.8860 18.6300 ;
      RECT 23.7520 17.5365 23.7780 18.6300 ;
      RECT 23.6440 17.5365 23.6700 18.6300 ;
      RECT 23.5360 17.5365 23.5620 18.6300 ;
      RECT 23.4280 17.5365 23.4540 18.6300 ;
      RECT 23.3200 17.5365 23.3460 18.6300 ;
      RECT 23.2120 17.5365 23.2380 18.6300 ;
      RECT 23.1040 17.5365 23.1300 18.6300 ;
      RECT 22.9960 17.5365 23.0220 18.6300 ;
      RECT 22.8880 17.5365 22.9140 18.6300 ;
      RECT 22.7800 17.5365 22.8060 18.6300 ;
      RECT 22.6720 17.5365 22.6980 18.6300 ;
      RECT 22.5640 17.5365 22.5900 18.6300 ;
      RECT 22.4560 17.5365 22.4820 18.6300 ;
      RECT 22.3480 17.5365 22.3740 18.6300 ;
      RECT 22.2400 17.5365 22.2660 18.6300 ;
      RECT 22.1320 17.5365 22.1580 18.6300 ;
      RECT 22.0240 17.5365 22.0500 18.6300 ;
      RECT 21.9160 17.5365 21.9420 18.6300 ;
      RECT 21.8080 17.5365 21.8340 18.6300 ;
      RECT 21.7000 17.5365 21.7260 18.6300 ;
      RECT 21.5920 17.5365 21.6180 18.6300 ;
      RECT 21.4840 17.5365 21.5100 18.6300 ;
      RECT 21.3760 17.5365 21.4020 18.6300 ;
      RECT 21.2680 17.5365 21.2940 18.6300 ;
      RECT 21.1600 17.5365 21.1860 18.6300 ;
      RECT 21.0520 17.5365 21.0780 18.6300 ;
      RECT 20.9440 17.5365 20.9700 18.6300 ;
      RECT 20.8360 17.5365 20.8620 18.6300 ;
      RECT 20.7280 17.5365 20.7540 18.6300 ;
      RECT 20.6200 17.5365 20.6460 18.6300 ;
      RECT 20.5120 17.5365 20.5380 18.6300 ;
      RECT 20.4040 17.5365 20.4300 18.6300 ;
      RECT 20.2960 17.5365 20.3220 18.6300 ;
      RECT 20.1880 17.5365 20.2140 18.6300 ;
      RECT 20.0800 17.5365 20.1060 18.6300 ;
      RECT 19.9720 17.5365 19.9980 18.6300 ;
      RECT 19.8640 17.5365 19.8900 18.6300 ;
      RECT 19.7560 17.5365 19.7820 18.6300 ;
      RECT 19.6480 17.5365 19.6740 18.6300 ;
      RECT 19.5400 17.5365 19.5660 18.6300 ;
      RECT 19.4320 17.5365 19.4580 18.6300 ;
      RECT 19.3240 17.5365 19.3500 18.6300 ;
      RECT 19.2160 17.5365 19.2420 18.6300 ;
      RECT 19.1080 17.5365 19.1340 18.6300 ;
      RECT 19.0000 17.5365 19.0260 18.6300 ;
      RECT 18.8920 17.5365 18.9180 18.6300 ;
      RECT 18.7840 17.5365 18.8100 18.6300 ;
      RECT 18.6760 17.5365 18.7020 18.6300 ;
      RECT 18.5680 17.5365 18.5940 18.6300 ;
      RECT 18.4600 17.5365 18.4860 18.6300 ;
      RECT 18.3520 17.5365 18.3780 18.6300 ;
      RECT 18.2440 17.5365 18.2700 18.6300 ;
      RECT 18.1360 17.5365 18.1620 18.6300 ;
      RECT 18.0280 17.5365 18.0540 18.6300 ;
      RECT 17.9200 17.5365 17.9460 18.6300 ;
      RECT 17.8120 17.5365 17.8380 18.6300 ;
      RECT 17.7040 17.5365 17.7300 18.6300 ;
      RECT 17.5960 17.5365 17.6220 18.6300 ;
      RECT 17.4880 17.5365 17.5140 18.6300 ;
      RECT 17.3800 17.5365 17.4060 18.6300 ;
      RECT 17.2720 17.5365 17.2980 18.6300 ;
      RECT 17.1640 17.5365 17.1900 18.6300 ;
      RECT 17.0560 17.5365 17.0820 18.6300 ;
      RECT 16.9480 17.5365 16.9740 18.6300 ;
      RECT 16.8400 17.5365 16.8660 18.6300 ;
      RECT 16.7320 17.5365 16.7580 18.6300 ;
      RECT 16.6240 17.5365 16.6500 18.6300 ;
      RECT 16.5160 17.5365 16.5420 18.6300 ;
      RECT 16.4080 17.5365 16.4340 18.6300 ;
      RECT 16.3000 17.5365 16.3260 18.6300 ;
      RECT 16.0870 17.5365 16.1640 18.6300 ;
      RECT 14.1940 17.5365 14.2710 18.6300 ;
      RECT 14.0320 17.5365 14.0580 18.6300 ;
      RECT 13.9240 17.5365 13.9500 18.6300 ;
      RECT 13.8160 17.5365 13.8420 18.6300 ;
      RECT 13.7080 17.5365 13.7340 18.6300 ;
      RECT 13.6000 17.5365 13.6260 18.6300 ;
      RECT 13.4920 17.5365 13.5180 18.6300 ;
      RECT 13.3840 17.5365 13.4100 18.6300 ;
      RECT 13.2760 17.5365 13.3020 18.6300 ;
      RECT 13.1680 17.5365 13.1940 18.6300 ;
      RECT 13.0600 17.5365 13.0860 18.6300 ;
      RECT 12.9520 17.5365 12.9780 18.6300 ;
      RECT 12.8440 17.5365 12.8700 18.6300 ;
      RECT 12.7360 17.5365 12.7620 18.6300 ;
      RECT 12.6280 17.5365 12.6540 18.6300 ;
      RECT 12.5200 17.5365 12.5460 18.6300 ;
      RECT 12.4120 17.5365 12.4380 18.6300 ;
      RECT 12.3040 17.5365 12.3300 18.6300 ;
      RECT 12.1960 17.5365 12.2220 18.6300 ;
      RECT 12.0880 17.5365 12.1140 18.6300 ;
      RECT 11.9800 17.5365 12.0060 18.6300 ;
      RECT 11.8720 17.5365 11.8980 18.6300 ;
      RECT 11.7640 17.5365 11.7900 18.6300 ;
      RECT 11.6560 17.5365 11.6820 18.6300 ;
      RECT 11.5480 17.5365 11.5740 18.6300 ;
      RECT 11.4400 17.5365 11.4660 18.6300 ;
      RECT 11.3320 17.5365 11.3580 18.6300 ;
      RECT 11.2240 17.5365 11.2500 18.6300 ;
      RECT 11.1160 17.5365 11.1420 18.6300 ;
      RECT 11.0080 17.5365 11.0340 18.6300 ;
      RECT 10.9000 17.5365 10.9260 18.6300 ;
      RECT 10.7920 17.5365 10.8180 18.6300 ;
      RECT 10.6840 17.5365 10.7100 18.6300 ;
      RECT 10.5760 17.5365 10.6020 18.6300 ;
      RECT 10.4680 17.5365 10.4940 18.6300 ;
      RECT 10.3600 17.5365 10.3860 18.6300 ;
      RECT 10.2520 17.5365 10.2780 18.6300 ;
      RECT 10.1440 17.5365 10.1700 18.6300 ;
      RECT 10.0360 17.5365 10.0620 18.6300 ;
      RECT 9.9280 17.5365 9.9540 18.6300 ;
      RECT 9.8200 17.5365 9.8460 18.6300 ;
      RECT 9.7120 17.5365 9.7380 18.6300 ;
      RECT 9.6040 17.5365 9.6300 18.6300 ;
      RECT 9.4960 17.5365 9.5220 18.6300 ;
      RECT 9.3880 17.5365 9.4140 18.6300 ;
      RECT 9.2800 17.5365 9.3060 18.6300 ;
      RECT 9.1720 17.5365 9.1980 18.6300 ;
      RECT 9.0640 17.5365 9.0900 18.6300 ;
      RECT 8.9560 17.5365 8.9820 18.6300 ;
      RECT 8.8480 17.5365 8.8740 18.6300 ;
      RECT 8.7400 17.5365 8.7660 18.6300 ;
      RECT 8.6320 17.5365 8.6580 18.6300 ;
      RECT 8.5240 17.5365 8.5500 18.6300 ;
      RECT 8.4160 17.5365 8.4420 18.6300 ;
      RECT 8.3080 17.5365 8.3340 18.6300 ;
      RECT 8.2000 17.5365 8.2260 18.6300 ;
      RECT 8.0920 17.5365 8.1180 18.6300 ;
      RECT 7.9840 17.5365 8.0100 18.6300 ;
      RECT 7.8760 17.5365 7.9020 18.6300 ;
      RECT 7.7680 17.5365 7.7940 18.6300 ;
      RECT 7.6600 17.5365 7.6860 18.6300 ;
      RECT 7.5520 17.5365 7.5780 18.6300 ;
      RECT 7.4440 17.5365 7.4700 18.6300 ;
      RECT 7.3360 17.5365 7.3620 18.6300 ;
      RECT 7.2280 17.5365 7.2540 18.6300 ;
      RECT 7.1200 17.5365 7.1460 18.6300 ;
      RECT 7.0120 17.5365 7.0380 18.6300 ;
      RECT 6.9040 17.5365 6.9300 18.6300 ;
      RECT 6.7960 17.5365 6.8220 18.6300 ;
      RECT 6.6880 17.5365 6.7140 18.6300 ;
      RECT 6.5800 17.5365 6.6060 18.6300 ;
      RECT 6.4720 17.5365 6.4980 18.6300 ;
      RECT 6.3640 17.5365 6.3900 18.6300 ;
      RECT 6.2560 17.5365 6.2820 18.6300 ;
      RECT 6.1480 17.5365 6.1740 18.6300 ;
      RECT 6.0400 17.5365 6.0660 18.6300 ;
      RECT 5.9320 17.5365 5.9580 18.6300 ;
      RECT 5.8240 17.5365 5.8500 18.6300 ;
      RECT 5.7160 17.5365 5.7420 18.6300 ;
      RECT 5.6080 17.5365 5.6340 18.6300 ;
      RECT 5.5000 17.5365 5.5260 18.6300 ;
      RECT 5.3920 17.5365 5.4180 18.6300 ;
      RECT 5.2840 17.5365 5.3100 18.6300 ;
      RECT 5.1760 17.5365 5.2020 18.6300 ;
      RECT 5.0680 17.5365 5.0940 18.6300 ;
      RECT 4.9600 17.5365 4.9860 18.6300 ;
      RECT 4.8520 17.5365 4.8780 18.6300 ;
      RECT 4.7440 17.5365 4.7700 18.6300 ;
      RECT 4.6360 17.5365 4.6620 18.6300 ;
      RECT 4.5280 17.5365 4.5540 18.6300 ;
      RECT 4.4200 17.5365 4.4460 18.6300 ;
      RECT 4.3120 17.5365 4.3380 18.6300 ;
      RECT 4.2040 17.5365 4.2300 18.6300 ;
      RECT 4.0960 17.5365 4.1220 18.6300 ;
      RECT 3.9880 17.5365 4.0140 18.6300 ;
      RECT 3.8800 17.5365 3.9060 18.6300 ;
      RECT 3.7720 17.5365 3.7980 18.6300 ;
      RECT 3.6640 17.5365 3.6900 18.6300 ;
      RECT 3.5560 17.5365 3.5820 18.6300 ;
      RECT 3.4480 17.5365 3.4740 18.6300 ;
      RECT 3.3400 17.5365 3.3660 18.6300 ;
      RECT 3.2320 17.5365 3.2580 18.6300 ;
      RECT 3.1240 17.5365 3.1500 18.6300 ;
      RECT 3.0160 17.5365 3.0420 18.6300 ;
      RECT 2.9080 17.5365 2.9340 18.6300 ;
      RECT 2.8000 17.5365 2.8260 18.6300 ;
      RECT 2.6920 17.5365 2.7180 18.6300 ;
      RECT 2.5840 17.5365 2.6100 18.6300 ;
      RECT 2.4760 17.5365 2.5020 18.6300 ;
      RECT 2.3680 17.5365 2.3940 18.6300 ;
      RECT 2.2600 17.5365 2.2860 18.6300 ;
      RECT 2.1520 17.5365 2.1780 18.6300 ;
      RECT 2.0440 17.5365 2.0700 18.6300 ;
      RECT 1.9360 17.5365 1.9620 18.6300 ;
      RECT 1.8280 17.5365 1.8540 18.6300 ;
      RECT 1.7200 17.5365 1.7460 18.6300 ;
      RECT 1.6120 17.5365 1.6380 18.6300 ;
      RECT 1.5040 17.5365 1.5300 18.6300 ;
      RECT 1.3960 17.5365 1.4220 18.6300 ;
      RECT 1.2880 17.5365 1.3140 18.6300 ;
      RECT 1.1800 17.5365 1.2060 18.6300 ;
      RECT 1.0720 17.5365 1.0980 18.6300 ;
      RECT 0.9640 17.5365 0.9900 18.6300 ;
      RECT 0.8560 17.5365 0.8820 18.6300 ;
      RECT 0.7480 17.5365 0.7740 18.6300 ;
      RECT 0.6400 17.5365 0.6660 18.6300 ;
      RECT 0.5320 17.5365 0.5580 18.6300 ;
      RECT 0.4240 17.5365 0.4500 18.6300 ;
      RECT 0.3160 17.5365 0.3420 18.6300 ;
      RECT 0.2080 17.5365 0.2340 18.6300 ;
      RECT 0.0050 17.5365 0.0900 18.6300 ;
      RECT 15.5530 18.6165 15.6810 19.7100 ;
      RECT 15.5390 19.2820 15.6810 19.6045 ;
      RECT 15.3190 19.0090 15.4530 19.7100 ;
      RECT 15.2960 19.3440 15.4530 19.6020 ;
      RECT 15.3190 18.6165 15.4170 19.7100 ;
      RECT 15.3190 18.7375 15.4310 18.9770 ;
      RECT 15.3190 18.6165 15.4530 18.7055 ;
      RECT 15.0940 19.0670 15.2280 19.7100 ;
      RECT 15.0940 18.6165 15.1920 19.7100 ;
      RECT 14.6770 18.6165 14.7600 19.7100 ;
      RECT 14.6770 18.7050 14.7740 19.6405 ;
      RECT 30.2680 18.6165 30.3530 19.7100 ;
      RECT 30.1240 18.6165 30.1500 19.7100 ;
      RECT 30.0160 18.6165 30.0420 19.7100 ;
      RECT 29.9080 18.6165 29.9340 19.7100 ;
      RECT 29.8000 18.6165 29.8260 19.7100 ;
      RECT 29.6920 18.6165 29.7180 19.7100 ;
      RECT 29.5840 18.6165 29.6100 19.7100 ;
      RECT 29.4760 18.6165 29.5020 19.7100 ;
      RECT 29.3680 18.6165 29.3940 19.7100 ;
      RECT 29.2600 18.6165 29.2860 19.7100 ;
      RECT 29.1520 18.6165 29.1780 19.7100 ;
      RECT 29.0440 18.6165 29.0700 19.7100 ;
      RECT 28.9360 18.6165 28.9620 19.7100 ;
      RECT 28.8280 18.6165 28.8540 19.7100 ;
      RECT 28.7200 18.6165 28.7460 19.7100 ;
      RECT 28.6120 18.6165 28.6380 19.7100 ;
      RECT 28.5040 18.6165 28.5300 19.7100 ;
      RECT 28.3960 18.6165 28.4220 19.7100 ;
      RECT 28.2880 18.6165 28.3140 19.7100 ;
      RECT 28.1800 18.6165 28.2060 19.7100 ;
      RECT 28.0720 18.6165 28.0980 19.7100 ;
      RECT 27.9640 18.6165 27.9900 19.7100 ;
      RECT 27.8560 18.6165 27.8820 19.7100 ;
      RECT 27.7480 18.6165 27.7740 19.7100 ;
      RECT 27.6400 18.6165 27.6660 19.7100 ;
      RECT 27.5320 18.6165 27.5580 19.7100 ;
      RECT 27.4240 18.6165 27.4500 19.7100 ;
      RECT 27.3160 18.6165 27.3420 19.7100 ;
      RECT 27.2080 18.6165 27.2340 19.7100 ;
      RECT 27.1000 18.6165 27.1260 19.7100 ;
      RECT 26.9920 18.6165 27.0180 19.7100 ;
      RECT 26.8840 18.6165 26.9100 19.7100 ;
      RECT 26.7760 18.6165 26.8020 19.7100 ;
      RECT 26.6680 18.6165 26.6940 19.7100 ;
      RECT 26.5600 18.6165 26.5860 19.7100 ;
      RECT 26.4520 18.6165 26.4780 19.7100 ;
      RECT 26.3440 18.6165 26.3700 19.7100 ;
      RECT 26.2360 18.6165 26.2620 19.7100 ;
      RECT 26.1280 18.6165 26.1540 19.7100 ;
      RECT 26.0200 18.6165 26.0460 19.7100 ;
      RECT 25.9120 18.6165 25.9380 19.7100 ;
      RECT 25.8040 18.6165 25.8300 19.7100 ;
      RECT 25.6960 18.6165 25.7220 19.7100 ;
      RECT 25.5880 18.6165 25.6140 19.7100 ;
      RECT 25.4800 18.6165 25.5060 19.7100 ;
      RECT 25.3720 18.6165 25.3980 19.7100 ;
      RECT 25.2640 18.6165 25.2900 19.7100 ;
      RECT 25.1560 18.6165 25.1820 19.7100 ;
      RECT 25.0480 18.6165 25.0740 19.7100 ;
      RECT 24.9400 18.6165 24.9660 19.7100 ;
      RECT 24.8320 18.6165 24.8580 19.7100 ;
      RECT 24.7240 18.6165 24.7500 19.7100 ;
      RECT 24.6160 18.6165 24.6420 19.7100 ;
      RECT 24.5080 18.6165 24.5340 19.7100 ;
      RECT 24.4000 18.6165 24.4260 19.7100 ;
      RECT 24.2920 18.6165 24.3180 19.7100 ;
      RECT 24.1840 18.6165 24.2100 19.7100 ;
      RECT 24.0760 18.6165 24.1020 19.7100 ;
      RECT 23.9680 18.6165 23.9940 19.7100 ;
      RECT 23.8600 18.6165 23.8860 19.7100 ;
      RECT 23.7520 18.6165 23.7780 19.7100 ;
      RECT 23.6440 18.6165 23.6700 19.7100 ;
      RECT 23.5360 18.6165 23.5620 19.7100 ;
      RECT 23.4280 18.6165 23.4540 19.7100 ;
      RECT 23.3200 18.6165 23.3460 19.7100 ;
      RECT 23.2120 18.6165 23.2380 19.7100 ;
      RECT 23.1040 18.6165 23.1300 19.7100 ;
      RECT 22.9960 18.6165 23.0220 19.7100 ;
      RECT 22.8880 18.6165 22.9140 19.7100 ;
      RECT 22.7800 18.6165 22.8060 19.7100 ;
      RECT 22.6720 18.6165 22.6980 19.7100 ;
      RECT 22.5640 18.6165 22.5900 19.7100 ;
      RECT 22.4560 18.6165 22.4820 19.7100 ;
      RECT 22.3480 18.6165 22.3740 19.7100 ;
      RECT 22.2400 18.6165 22.2660 19.7100 ;
      RECT 22.1320 18.6165 22.1580 19.7100 ;
      RECT 22.0240 18.6165 22.0500 19.7100 ;
      RECT 21.9160 18.6165 21.9420 19.7100 ;
      RECT 21.8080 18.6165 21.8340 19.7100 ;
      RECT 21.7000 18.6165 21.7260 19.7100 ;
      RECT 21.5920 18.6165 21.6180 19.7100 ;
      RECT 21.4840 18.6165 21.5100 19.7100 ;
      RECT 21.3760 18.6165 21.4020 19.7100 ;
      RECT 21.2680 18.6165 21.2940 19.7100 ;
      RECT 21.1600 18.6165 21.1860 19.7100 ;
      RECT 21.0520 18.6165 21.0780 19.7100 ;
      RECT 20.9440 18.6165 20.9700 19.7100 ;
      RECT 20.8360 18.6165 20.8620 19.7100 ;
      RECT 20.7280 18.6165 20.7540 19.7100 ;
      RECT 20.6200 18.6165 20.6460 19.7100 ;
      RECT 20.5120 18.6165 20.5380 19.7100 ;
      RECT 20.4040 18.6165 20.4300 19.7100 ;
      RECT 20.2960 18.6165 20.3220 19.7100 ;
      RECT 20.1880 18.6165 20.2140 19.7100 ;
      RECT 20.0800 18.6165 20.1060 19.7100 ;
      RECT 19.9720 18.6165 19.9980 19.7100 ;
      RECT 19.8640 18.6165 19.8900 19.7100 ;
      RECT 19.7560 18.6165 19.7820 19.7100 ;
      RECT 19.6480 18.6165 19.6740 19.7100 ;
      RECT 19.5400 18.6165 19.5660 19.7100 ;
      RECT 19.4320 18.6165 19.4580 19.7100 ;
      RECT 19.3240 18.6165 19.3500 19.7100 ;
      RECT 19.2160 18.6165 19.2420 19.7100 ;
      RECT 19.1080 18.6165 19.1340 19.7100 ;
      RECT 19.0000 18.6165 19.0260 19.7100 ;
      RECT 18.8920 18.6165 18.9180 19.7100 ;
      RECT 18.7840 18.6165 18.8100 19.7100 ;
      RECT 18.6760 18.6165 18.7020 19.7100 ;
      RECT 18.5680 18.6165 18.5940 19.7100 ;
      RECT 18.4600 18.6165 18.4860 19.7100 ;
      RECT 18.3520 18.6165 18.3780 19.7100 ;
      RECT 18.2440 18.6165 18.2700 19.7100 ;
      RECT 18.1360 18.6165 18.1620 19.7100 ;
      RECT 18.0280 18.6165 18.0540 19.7100 ;
      RECT 17.9200 18.6165 17.9460 19.7100 ;
      RECT 17.8120 18.6165 17.8380 19.7100 ;
      RECT 17.7040 18.6165 17.7300 19.7100 ;
      RECT 17.5960 18.6165 17.6220 19.7100 ;
      RECT 17.4880 18.6165 17.5140 19.7100 ;
      RECT 17.3800 18.6165 17.4060 19.7100 ;
      RECT 17.2720 18.6165 17.2980 19.7100 ;
      RECT 17.1640 18.6165 17.1900 19.7100 ;
      RECT 17.0560 18.6165 17.0820 19.7100 ;
      RECT 16.9480 18.6165 16.9740 19.7100 ;
      RECT 16.8400 18.6165 16.8660 19.7100 ;
      RECT 16.7320 18.6165 16.7580 19.7100 ;
      RECT 16.6240 18.6165 16.6500 19.7100 ;
      RECT 16.5160 18.6165 16.5420 19.7100 ;
      RECT 16.4080 18.6165 16.4340 19.7100 ;
      RECT 16.3000 18.6165 16.3260 19.7100 ;
      RECT 16.0870 18.6165 16.1640 19.7100 ;
      RECT 14.1940 18.6165 14.2710 19.7100 ;
      RECT 14.0320 18.6165 14.0580 19.7100 ;
      RECT 13.9240 18.6165 13.9500 19.7100 ;
      RECT 13.8160 18.6165 13.8420 19.7100 ;
      RECT 13.7080 18.6165 13.7340 19.7100 ;
      RECT 13.6000 18.6165 13.6260 19.7100 ;
      RECT 13.4920 18.6165 13.5180 19.7100 ;
      RECT 13.3840 18.6165 13.4100 19.7100 ;
      RECT 13.2760 18.6165 13.3020 19.7100 ;
      RECT 13.1680 18.6165 13.1940 19.7100 ;
      RECT 13.0600 18.6165 13.0860 19.7100 ;
      RECT 12.9520 18.6165 12.9780 19.7100 ;
      RECT 12.8440 18.6165 12.8700 19.7100 ;
      RECT 12.7360 18.6165 12.7620 19.7100 ;
      RECT 12.6280 18.6165 12.6540 19.7100 ;
      RECT 12.5200 18.6165 12.5460 19.7100 ;
      RECT 12.4120 18.6165 12.4380 19.7100 ;
      RECT 12.3040 18.6165 12.3300 19.7100 ;
      RECT 12.1960 18.6165 12.2220 19.7100 ;
      RECT 12.0880 18.6165 12.1140 19.7100 ;
      RECT 11.9800 18.6165 12.0060 19.7100 ;
      RECT 11.8720 18.6165 11.8980 19.7100 ;
      RECT 11.7640 18.6165 11.7900 19.7100 ;
      RECT 11.6560 18.6165 11.6820 19.7100 ;
      RECT 11.5480 18.6165 11.5740 19.7100 ;
      RECT 11.4400 18.6165 11.4660 19.7100 ;
      RECT 11.3320 18.6165 11.3580 19.7100 ;
      RECT 11.2240 18.6165 11.2500 19.7100 ;
      RECT 11.1160 18.6165 11.1420 19.7100 ;
      RECT 11.0080 18.6165 11.0340 19.7100 ;
      RECT 10.9000 18.6165 10.9260 19.7100 ;
      RECT 10.7920 18.6165 10.8180 19.7100 ;
      RECT 10.6840 18.6165 10.7100 19.7100 ;
      RECT 10.5760 18.6165 10.6020 19.7100 ;
      RECT 10.4680 18.6165 10.4940 19.7100 ;
      RECT 10.3600 18.6165 10.3860 19.7100 ;
      RECT 10.2520 18.6165 10.2780 19.7100 ;
      RECT 10.1440 18.6165 10.1700 19.7100 ;
      RECT 10.0360 18.6165 10.0620 19.7100 ;
      RECT 9.9280 18.6165 9.9540 19.7100 ;
      RECT 9.8200 18.6165 9.8460 19.7100 ;
      RECT 9.7120 18.6165 9.7380 19.7100 ;
      RECT 9.6040 18.6165 9.6300 19.7100 ;
      RECT 9.4960 18.6165 9.5220 19.7100 ;
      RECT 9.3880 18.6165 9.4140 19.7100 ;
      RECT 9.2800 18.6165 9.3060 19.7100 ;
      RECT 9.1720 18.6165 9.1980 19.7100 ;
      RECT 9.0640 18.6165 9.0900 19.7100 ;
      RECT 8.9560 18.6165 8.9820 19.7100 ;
      RECT 8.8480 18.6165 8.8740 19.7100 ;
      RECT 8.7400 18.6165 8.7660 19.7100 ;
      RECT 8.6320 18.6165 8.6580 19.7100 ;
      RECT 8.5240 18.6165 8.5500 19.7100 ;
      RECT 8.4160 18.6165 8.4420 19.7100 ;
      RECT 8.3080 18.6165 8.3340 19.7100 ;
      RECT 8.2000 18.6165 8.2260 19.7100 ;
      RECT 8.0920 18.6165 8.1180 19.7100 ;
      RECT 7.9840 18.6165 8.0100 19.7100 ;
      RECT 7.8760 18.6165 7.9020 19.7100 ;
      RECT 7.7680 18.6165 7.7940 19.7100 ;
      RECT 7.6600 18.6165 7.6860 19.7100 ;
      RECT 7.5520 18.6165 7.5780 19.7100 ;
      RECT 7.4440 18.6165 7.4700 19.7100 ;
      RECT 7.3360 18.6165 7.3620 19.7100 ;
      RECT 7.2280 18.6165 7.2540 19.7100 ;
      RECT 7.1200 18.6165 7.1460 19.7100 ;
      RECT 7.0120 18.6165 7.0380 19.7100 ;
      RECT 6.9040 18.6165 6.9300 19.7100 ;
      RECT 6.7960 18.6165 6.8220 19.7100 ;
      RECT 6.6880 18.6165 6.7140 19.7100 ;
      RECT 6.5800 18.6165 6.6060 19.7100 ;
      RECT 6.4720 18.6165 6.4980 19.7100 ;
      RECT 6.3640 18.6165 6.3900 19.7100 ;
      RECT 6.2560 18.6165 6.2820 19.7100 ;
      RECT 6.1480 18.6165 6.1740 19.7100 ;
      RECT 6.0400 18.6165 6.0660 19.7100 ;
      RECT 5.9320 18.6165 5.9580 19.7100 ;
      RECT 5.8240 18.6165 5.8500 19.7100 ;
      RECT 5.7160 18.6165 5.7420 19.7100 ;
      RECT 5.6080 18.6165 5.6340 19.7100 ;
      RECT 5.5000 18.6165 5.5260 19.7100 ;
      RECT 5.3920 18.6165 5.4180 19.7100 ;
      RECT 5.2840 18.6165 5.3100 19.7100 ;
      RECT 5.1760 18.6165 5.2020 19.7100 ;
      RECT 5.0680 18.6165 5.0940 19.7100 ;
      RECT 4.9600 18.6165 4.9860 19.7100 ;
      RECT 4.8520 18.6165 4.8780 19.7100 ;
      RECT 4.7440 18.6165 4.7700 19.7100 ;
      RECT 4.6360 18.6165 4.6620 19.7100 ;
      RECT 4.5280 18.6165 4.5540 19.7100 ;
      RECT 4.4200 18.6165 4.4460 19.7100 ;
      RECT 4.3120 18.6165 4.3380 19.7100 ;
      RECT 4.2040 18.6165 4.2300 19.7100 ;
      RECT 4.0960 18.6165 4.1220 19.7100 ;
      RECT 3.9880 18.6165 4.0140 19.7100 ;
      RECT 3.8800 18.6165 3.9060 19.7100 ;
      RECT 3.7720 18.6165 3.7980 19.7100 ;
      RECT 3.6640 18.6165 3.6900 19.7100 ;
      RECT 3.5560 18.6165 3.5820 19.7100 ;
      RECT 3.4480 18.6165 3.4740 19.7100 ;
      RECT 3.3400 18.6165 3.3660 19.7100 ;
      RECT 3.2320 18.6165 3.2580 19.7100 ;
      RECT 3.1240 18.6165 3.1500 19.7100 ;
      RECT 3.0160 18.6165 3.0420 19.7100 ;
      RECT 2.9080 18.6165 2.9340 19.7100 ;
      RECT 2.8000 18.6165 2.8260 19.7100 ;
      RECT 2.6920 18.6165 2.7180 19.7100 ;
      RECT 2.5840 18.6165 2.6100 19.7100 ;
      RECT 2.4760 18.6165 2.5020 19.7100 ;
      RECT 2.3680 18.6165 2.3940 19.7100 ;
      RECT 2.2600 18.6165 2.2860 19.7100 ;
      RECT 2.1520 18.6165 2.1780 19.7100 ;
      RECT 2.0440 18.6165 2.0700 19.7100 ;
      RECT 1.9360 18.6165 1.9620 19.7100 ;
      RECT 1.8280 18.6165 1.8540 19.7100 ;
      RECT 1.7200 18.6165 1.7460 19.7100 ;
      RECT 1.6120 18.6165 1.6380 19.7100 ;
      RECT 1.5040 18.6165 1.5300 19.7100 ;
      RECT 1.3960 18.6165 1.4220 19.7100 ;
      RECT 1.2880 18.6165 1.3140 19.7100 ;
      RECT 1.1800 18.6165 1.2060 19.7100 ;
      RECT 1.0720 18.6165 1.0980 19.7100 ;
      RECT 0.9640 18.6165 0.9900 19.7100 ;
      RECT 0.8560 18.6165 0.8820 19.7100 ;
      RECT 0.7480 18.6165 0.7740 19.7100 ;
      RECT 0.6400 18.6165 0.6660 19.7100 ;
      RECT 0.5320 18.6165 0.5580 19.7100 ;
      RECT 0.4240 18.6165 0.4500 19.7100 ;
      RECT 0.3160 18.6165 0.3420 19.7100 ;
      RECT 0.2080 18.6165 0.2340 19.7100 ;
      RECT 0.0050 18.6165 0.0900 19.7100 ;
      RECT 15.5530 19.6965 15.6810 20.7900 ;
      RECT 15.5390 20.3620 15.6810 20.6845 ;
      RECT 15.3190 20.0890 15.4530 20.7900 ;
      RECT 15.2960 20.4240 15.4530 20.6820 ;
      RECT 15.3190 19.6965 15.4170 20.7900 ;
      RECT 15.3190 19.8175 15.4310 20.0570 ;
      RECT 15.3190 19.6965 15.4530 19.7855 ;
      RECT 15.0940 20.1470 15.2280 20.7900 ;
      RECT 15.0940 19.6965 15.1920 20.7900 ;
      RECT 14.6770 19.6965 14.7600 20.7900 ;
      RECT 14.6770 19.7850 14.7740 20.7205 ;
      RECT 30.2680 19.6965 30.3530 20.7900 ;
      RECT 30.1240 19.6965 30.1500 20.7900 ;
      RECT 30.0160 19.6965 30.0420 20.7900 ;
      RECT 29.9080 19.6965 29.9340 20.7900 ;
      RECT 29.8000 19.6965 29.8260 20.7900 ;
      RECT 29.6920 19.6965 29.7180 20.7900 ;
      RECT 29.5840 19.6965 29.6100 20.7900 ;
      RECT 29.4760 19.6965 29.5020 20.7900 ;
      RECT 29.3680 19.6965 29.3940 20.7900 ;
      RECT 29.2600 19.6965 29.2860 20.7900 ;
      RECT 29.1520 19.6965 29.1780 20.7900 ;
      RECT 29.0440 19.6965 29.0700 20.7900 ;
      RECT 28.9360 19.6965 28.9620 20.7900 ;
      RECT 28.8280 19.6965 28.8540 20.7900 ;
      RECT 28.7200 19.6965 28.7460 20.7900 ;
      RECT 28.6120 19.6965 28.6380 20.7900 ;
      RECT 28.5040 19.6965 28.5300 20.7900 ;
      RECT 28.3960 19.6965 28.4220 20.7900 ;
      RECT 28.2880 19.6965 28.3140 20.7900 ;
      RECT 28.1800 19.6965 28.2060 20.7900 ;
      RECT 28.0720 19.6965 28.0980 20.7900 ;
      RECT 27.9640 19.6965 27.9900 20.7900 ;
      RECT 27.8560 19.6965 27.8820 20.7900 ;
      RECT 27.7480 19.6965 27.7740 20.7900 ;
      RECT 27.6400 19.6965 27.6660 20.7900 ;
      RECT 27.5320 19.6965 27.5580 20.7900 ;
      RECT 27.4240 19.6965 27.4500 20.7900 ;
      RECT 27.3160 19.6965 27.3420 20.7900 ;
      RECT 27.2080 19.6965 27.2340 20.7900 ;
      RECT 27.1000 19.6965 27.1260 20.7900 ;
      RECT 26.9920 19.6965 27.0180 20.7900 ;
      RECT 26.8840 19.6965 26.9100 20.7900 ;
      RECT 26.7760 19.6965 26.8020 20.7900 ;
      RECT 26.6680 19.6965 26.6940 20.7900 ;
      RECT 26.5600 19.6965 26.5860 20.7900 ;
      RECT 26.4520 19.6965 26.4780 20.7900 ;
      RECT 26.3440 19.6965 26.3700 20.7900 ;
      RECT 26.2360 19.6965 26.2620 20.7900 ;
      RECT 26.1280 19.6965 26.1540 20.7900 ;
      RECT 26.0200 19.6965 26.0460 20.7900 ;
      RECT 25.9120 19.6965 25.9380 20.7900 ;
      RECT 25.8040 19.6965 25.8300 20.7900 ;
      RECT 25.6960 19.6965 25.7220 20.7900 ;
      RECT 25.5880 19.6965 25.6140 20.7900 ;
      RECT 25.4800 19.6965 25.5060 20.7900 ;
      RECT 25.3720 19.6965 25.3980 20.7900 ;
      RECT 25.2640 19.6965 25.2900 20.7900 ;
      RECT 25.1560 19.6965 25.1820 20.7900 ;
      RECT 25.0480 19.6965 25.0740 20.7900 ;
      RECT 24.9400 19.6965 24.9660 20.7900 ;
      RECT 24.8320 19.6965 24.8580 20.7900 ;
      RECT 24.7240 19.6965 24.7500 20.7900 ;
      RECT 24.6160 19.6965 24.6420 20.7900 ;
      RECT 24.5080 19.6965 24.5340 20.7900 ;
      RECT 24.4000 19.6965 24.4260 20.7900 ;
      RECT 24.2920 19.6965 24.3180 20.7900 ;
      RECT 24.1840 19.6965 24.2100 20.7900 ;
      RECT 24.0760 19.6965 24.1020 20.7900 ;
      RECT 23.9680 19.6965 23.9940 20.7900 ;
      RECT 23.8600 19.6965 23.8860 20.7900 ;
      RECT 23.7520 19.6965 23.7780 20.7900 ;
      RECT 23.6440 19.6965 23.6700 20.7900 ;
      RECT 23.5360 19.6965 23.5620 20.7900 ;
      RECT 23.4280 19.6965 23.4540 20.7900 ;
      RECT 23.3200 19.6965 23.3460 20.7900 ;
      RECT 23.2120 19.6965 23.2380 20.7900 ;
      RECT 23.1040 19.6965 23.1300 20.7900 ;
      RECT 22.9960 19.6965 23.0220 20.7900 ;
      RECT 22.8880 19.6965 22.9140 20.7900 ;
      RECT 22.7800 19.6965 22.8060 20.7900 ;
      RECT 22.6720 19.6965 22.6980 20.7900 ;
      RECT 22.5640 19.6965 22.5900 20.7900 ;
      RECT 22.4560 19.6965 22.4820 20.7900 ;
      RECT 22.3480 19.6965 22.3740 20.7900 ;
      RECT 22.2400 19.6965 22.2660 20.7900 ;
      RECT 22.1320 19.6965 22.1580 20.7900 ;
      RECT 22.0240 19.6965 22.0500 20.7900 ;
      RECT 21.9160 19.6965 21.9420 20.7900 ;
      RECT 21.8080 19.6965 21.8340 20.7900 ;
      RECT 21.7000 19.6965 21.7260 20.7900 ;
      RECT 21.5920 19.6965 21.6180 20.7900 ;
      RECT 21.4840 19.6965 21.5100 20.7900 ;
      RECT 21.3760 19.6965 21.4020 20.7900 ;
      RECT 21.2680 19.6965 21.2940 20.7900 ;
      RECT 21.1600 19.6965 21.1860 20.7900 ;
      RECT 21.0520 19.6965 21.0780 20.7900 ;
      RECT 20.9440 19.6965 20.9700 20.7900 ;
      RECT 20.8360 19.6965 20.8620 20.7900 ;
      RECT 20.7280 19.6965 20.7540 20.7900 ;
      RECT 20.6200 19.6965 20.6460 20.7900 ;
      RECT 20.5120 19.6965 20.5380 20.7900 ;
      RECT 20.4040 19.6965 20.4300 20.7900 ;
      RECT 20.2960 19.6965 20.3220 20.7900 ;
      RECT 20.1880 19.6965 20.2140 20.7900 ;
      RECT 20.0800 19.6965 20.1060 20.7900 ;
      RECT 19.9720 19.6965 19.9980 20.7900 ;
      RECT 19.8640 19.6965 19.8900 20.7900 ;
      RECT 19.7560 19.6965 19.7820 20.7900 ;
      RECT 19.6480 19.6965 19.6740 20.7900 ;
      RECT 19.5400 19.6965 19.5660 20.7900 ;
      RECT 19.4320 19.6965 19.4580 20.7900 ;
      RECT 19.3240 19.6965 19.3500 20.7900 ;
      RECT 19.2160 19.6965 19.2420 20.7900 ;
      RECT 19.1080 19.6965 19.1340 20.7900 ;
      RECT 19.0000 19.6965 19.0260 20.7900 ;
      RECT 18.8920 19.6965 18.9180 20.7900 ;
      RECT 18.7840 19.6965 18.8100 20.7900 ;
      RECT 18.6760 19.6965 18.7020 20.7900 ;
      RECT 18.5680 19.6965 18.5940 20.7900 ;
      RECT 18.4600 19.6965 18.4860 20.7900 ;
      RECT 18.3520 19.6965 18.3780 20.7900 ;
      RECT 18.2440 19.6965 18.2700 20.7900 ;
      RECT 18.1360 19.6965 18.1620 20.7900 ;
      RECT 18.0280 19.6965 18.0540 20.7900 ;
      RECT 17.9200 19.6965 17.9460 20.7900 ;
      RECT 17.8120 19.6965 17.8380 20.7900 ;
      RECT 17.7040 19.6965 17.7300 20.7900 ;
      RECT 17.5960 19.6965 17.6220 20.7900 ;
      RECT 17.4880 19.6965 17.5140 20.7900 ;
      RECT 17.3800 19.6965 17.4060 20.7900 ;
      RECT 17.2720 19.6965 17.2980 20.7900 ;
      RECT 17.1640 19.6965 17.1900 20.7900 ;
      RECT 17.0560 19.6965 17.0820 20.7900 ;
      RECT 16.9480 19.6965 16.9740 20.7900 ;
      RECT 16.8400 19.6965 16.8660 20.7900 ;
      RECT 16.7320 19.6965 16.7580 20.7900 ;
      RECT 16.6240 19.6965 16.6500 20.7900 ;
      RECT 16.5160 19.6965 16.5420 20.7900 ;
      RECT 16.4080 19.6965 16.4340 20.7900 ;
      RECT 16.3000 19.6965 16.3260 20.7900 ;
      RECT 16.0870 19.6965 16.1640 20.7900 ;
      RECT 14.1940 19.6965 14.2710 20.7900 ;
      RECT 14.0320 19.6965 14.0580 20.7900 ;
      RECT 13.9240 19.6965 13.9500 20.7900 ;
      RECT 13.8160 19.6965 13.8420 20.7900 ;
      RECT 13.7080 19.6965 13.7340 20.7900 ;
      RECT 13.6000 19.6965 13.6260 20.7900 ;
      RECT 13.4920 19.6965 13.5180 20.7900 ;
      RECT 13.3840 19.6965 13.4100 20.7900 ;
      RECT 13.2760 19.6965 13.3020 20.7900 ;
      RECT 13.1680 19.6965 13.1940 20.7900 ;
      RECT 13.0600 19.6965 13.0860 20.7900 ;
      RECT 12.9520 19.6965 12.9780 20.7900 ;
      RECT 12.8440 19.6965 12.8700 20.7900 ;
      RECT 12.7360 19.6965 12.7620 20.7900 ;
      RECT 12.6280 19.6965 12.6540 20.7900 ;
      RECT 12.5200 19.6965 12.5460 20.7900 ;
      RECT 12.4120 19.6965 12.4380 20.7900 ;
      RECT 12.3040 19.6965 12.3300 20.7900 ;
      RECT 12.1960 19.6965 12.2220 20.7900 ;
      RECT 12.0880 19.6965 12.1140 20.7900 ;
      RECT 11.9800 19.6965 12.0060 20.7900 ;
      RECT 11.8720 19.6965 11.8980 20.7900 ;
      RECT 11.7640 19.6965 11.7900 20.7900 ;
      RECT 11.6560 19.6965 11.6820 20.7900 ;
      RECT 11.5480 19.6965 11.5740 20.7900 ;
      RECT 11.4400 19.6965 11.4660 20.7900 ;
      RECT 11.3320 19.6965 11.3580 20.7900 ;
      RECT 11.2240 19.6965 11.2500 20.7900 ;
      RECT 11.1160 19.6965 11.1420 20.7900 ;
      RECT 11.0080 19.6965 11.0340 20.7900 ;
      RECT 10.9000 19.6965 10.9260 20.7900 ;
      RECT 10.7920 19.6965 10.8180 20.7900 ;
      RECT 10.6840 19.6965 10.7100 20.7900 ;
      RECT 10.5760 19.6965 10.6020 20.7900 ;
      RECT 10.4680 19.6965 10.4940 20.7900 ;
      RECT 10.3600 19.6965 10.3860 20.7900 ;
      RECT 10.2520 19.6965 10.2780 20.7900 ;
      RECT 10.1440 19.6965 10.1700 20.7900 ;
      RECT 10.0360 19.6965 10.0620 20.7900 ;
      RECT 9.9280 19.6965 9.9540 20.7900 ;
      RECT 9.8200 19.6965 9.8460 20.7900 ;
      RECT 9.7120 19.6965 9.7380 20.7900 ;
      RECT 9.6040 19.6965 9.6300 20.7900 ;
      RECT 9.4960 19.6965 9.5220 20.7900 ;
      RECT 9.3880 19.6965 9.4140 20.7900 ;
      RECT 9.2800 19.6965 9.3060 20.7900 ;
      RECT 9.1720 19.6965 9.1980 20.7900 ;
      RECT 9.0640 19.6965 9.0900 20.7900 ;
      RECT 8.9560 19.6965 8.9820 20.7900 ;
      RECT 8.8480 19.6965 8.8740 20.7900 ;
      RECT 8.7400 19.6965 8.7660 20.7900 ;
      RECT 8.6320 19.6965 8.6580 20.7900 ;
      RECT 8.5240 19.6965 8.5500 20.7900 ;
      RECT 8.4160 19.6965 8.4420 20.7900 ;
      RECT 8.3080 19.6965 8.3340 20.7900 ;
      RECT 8.2000 19.6965 8.2260 20.7900 ;
      RECT 8.0920 19.6965 8.1180 20.7900 ;
      RECT 7.9840 19.6965 8.0100 20.7900 ;
      RECT 7.8760 19.6965 7.9020 20.7900 ;
      RECT 7.7680 19.6965 7.7940 20.7900 ;
      RECT 7.6600 19.6965 7.6860 20.7900 ;
      RECT 7.5520 19.6965 7.5780 20.7900 ;
      RECT 7.4440 19.6965 7.4700 20.7900 ;
      RECT 7.3360 19.6965 7.3620 20.7900 ;
      RECT 7.2280 19.6965 7.2540 20.7900 ;
      RECT 7.1200 19.6965 7.1460 20.7900 ;
      RECT 7.0120 19.6965 7.0380 20.7900 ;
      RECT 6.9040 19.6965 6.9300 20.7900 ;
      RECT 6.7960 19.6965 6.8220 20.7900 ;
      RECT 6.6880 19.6965 6.7140 20.7900 ;
      RECT 6.5800 19.6965 6.6060 20.7900 ;
      RECT 6.4720 19.6965 6.4980 20.7900 ;
      RECT 6.3640 19.6965 6.3900 20.7900 ;
      RECT 6.2560 19.6965 6.2820 20.7900 ;
      RECT 6.1480 19.6965 6.1740 20.7900 ;
      RECT 6.0400 19.6965 6.0660 20.7900 ;
      RECT 5.9320 19.6965 5.9580 20.7900 ;
      RECT 5.8240 19.6965 5.8500 20.7900 ;
      RECT 5.7160 19.6965 5.7420 20.7900 ;
      RECT 5.6080 19.6965 5.6340 20.7900 ;
      RECT 5.5000 19.6965 5.5260 20.7900 ;
      RECT 5.3920 19.6965 5.4180 20.7900 ;
      RECT 5.2840 19.6965 5.3100 20.7900 ;
      RECT 5.1760 19.6965 5.2020 20.7900 ;
      RECT 5.0680 19.6965 5.0940 20.7900 ;
      RECT 4.9600 19.6965 4.9860 20.7900 ;
      RECT 4.8520 19.6965 4.8780 20.7900 ;
      RECT 4.7440 19.6965 4.7700 20.7900 ;
      RECT 4.6360 19.6965 4.6620 20.7900 ;
      RECT 4.5280 19.6965 4.5540 20.7900 ;
      RECT 4.4200 19.6965 4.4460 20.7900 ;
      RECT 4.3120 19.6965 4.3380 20.7900 ;
      RECT 4.2040 19.6965 4.2300 20.7900 ;
      RECT 4.0960 19.6965 4.1220 20.7900 ;
      RECT 3.9880 19.6965 4.0140 20.7900 ;
      RECT 3.8800 19.6965 3.9060 20.7900 ;
      RECT 3.7720 19.6965 3.7980 20.7900 ;
      RECT 3.6640 19.6965 3.6900 20.7900 ;
      RECT 3.5560 19.6965 3.5820 20.7900 ;
      RECT 3.4480 19.6965 3.4740 20.7900 ;
      RECT 3.3400 19.6965 3.3660 20.7900 ;
      RECT 3.2320 19.6965 3.2580 20.7900 ;
      RECT 3.1240 19.6965 3.1500 20.7900 ;
      RECT 3.0160 19.6965 3.0420 20.7900 ;
      RECT 2.9080 19.6965 2.9340 20.7900 ;
      RECT 2.8000 19.6965 2.8260 20.7900 ;
      RECT 2.6920 19.6965 2.7180 20.7900 ;
      RECT 2.5840 19.6965 2.6100 20.7900 ;
      RECT 2.4760 19.6965 2.5020 20.7900 ;
      RECT 2.3680 19.6965 2.3940 20.7900 ;
      RECT 2.2600 19.6965 2.2860 20.7900 ;
      RECT 2.1520 19.6965 2.1780 20.7900 ;
      RECT 2.0440 19.6965 2.0700 20.7900 ;
      RECT 1.9360 19.6965 1.9620 20.7900 ;
      RECT 1.8280 19.6965 1.8540 20.7900 ;
      RECT 1.7200 19.6965 1.7460 20.7900 ;
      RECT 1.6120 19.6965 1.6380 20.7900 ;
      RECT 1.5040 19.6965 1.5300 20.7900 ;
      RECT 1.3960 19.6965 1.4220 20.7900 ;
      RECT 1.2880 19.6965 1.3140 20.7900 ;
      RECT 1.1800 19.6965 1.2060 20.7900 ;
      RECT 1.0720 19.6965 1.0980 20.7900 ;
      RECT 0.9640 19.6965 0.9900 20.7900 ;
      RECT 0.8560 19.6965 0.8820 20.7900 ;
      RECT 0.7480 19.6965 0.7740 20.7900 ;
      RECT 0.6400 19.6965 0.6660 20.7900 ;
      RECT 0.5320 19.6965 0.5580 20.7900 ;
      RECT 0.4240 19.6965 0.4500 20.7900 ;
      RECT 0.3160 19.6965 0.3420 20.7900 ;
      RECT 0.2080 19.6965 0.2340 20.7900 ;
      RECT 0.0050 19.6965 0.0900 20.7900 ;
      RECT 15.5530 20.7765 15.6810 21.8700 ;
      RECT 15.5390 21.4420 15.6810 21.7645 ;
      RECT 15.3190 21.1690 15.4530 21.8700 ;
      RECT 15.2960 21.5040 15.4530 21.7620 ;
      RECT 15.3190 20.7765 15.4170 21.8700 ;
      RECT 15.3190 20.8975 15.4310 21.1370 ;
      RECT 15.3190 20.7765 15.4530 20.8655 ;
      RECT 15.0940 21.2270 15.2280 21.8700 ;
      RECT 15.0940 20.7765 15.1920 21.8700 ;
      RECT 14.6770 20.7765 14.7600 21.8700 ;
      RECT 14.6770 20.8650 14.7740 21.8005 ;
      RECT 30.2680 20.7765 30.3530 21.8700 ;
      RECT 30.1240 20.7765 30.1500 21.8700 ;
      RECT 30.0160 20.7765 30.0420 21.8700 ;
      RECT 29.9080 20.7765 29.9340 21.8700 ;
      RECT 29.8000 20.7765 29.8260 21.8700 ;
      RECT 29.6920 20.7765 29.7180 21.8700 ;
      RECT 29.5840 20.7765 29.6100 21.8700 ;
      RECT 29.4760 20.7765 29.5020 21.8700 ;
      RECT 29.3680 20.7765 29.3940 21.8700 ;
      RECT 29.2600 20.7765 29.2860 21.8700 ;
      RECT 29.1520 20.7765 29.1780 21.8700 ;
      RECT 29.0440 20.7765 29.0700 21.8700 ;
      RECT 28.9360 20.7765 28.9620 21.8700 ;
      RECT 28.8280 20.7765 28.8540 21.8700 ;
      RECT 28.7200 20.7765 28.7460 21.8700 ;
      RECT 28.6120 20.7765 28.6380 21.8700 ;
      RECT 28.5040 20.7765 28.5300 21.8700 ;
      RECT 28.3960 20.7765 28.4220 21.8700 ;
      RECT 28.2880 20.7765 28.3140 21.8700 ;
      RECT 28.1800 20.7765 28.2060 21.8700 ;
      RECT 28.0720 20.7765 28.0980 21.8700 ;
      RECT 27.9640 20.7765 27.9900 21.8700 ;
      RECT 27.8560 20.7765 27.8820 21.8700 ;
      RECT 27.7480 20.7765 27.7740 21.8700 ;
      RECT 27.6400 20.7765 27.6660 21.8700 ;
      RECT 27.5320 20.7765 27.5580 21.8700 ;
      RECT 27.4240 20.7765 27.4500 21.8700 ;
      RECT 27.3160 20.7765 27.3420 21.8700 ;
      RECT 27.2080 20.7765 27.2340 21.8700 ;
      RECT 27.1000 20.7765 27.1260 21.8700 ;
      RECT 26.9920 20.7765 27.0180 21.8700 ;
      RECT 26.8840 20.7765 26.9100 21.8700 ;
      RECT 26.7760 20.7765 26.8020 21.8700 ;
      RECT 26.6680 20.7765 26.6940 21.8700 ;
      RECT 26.5600 20.7765 26.5860 21.8700 ;
      RECT 26.4520 20.7765 26.4780 21.8700 ;
      RECT 26.3440 20.7765 26.3700 21.8700 ;
      RECT 26.2360 20.7765 26.2620 21.8700 ;
      RECT 26.1280 20.7765 26.1540 21.8700 ;
      RECT 26.0200 20.7765 26.0460 21.8700 ;
      RECT 25.9120 20.7765 25.9380 21.8700 ;
      RECT 25.8040 20.7765 25.8300 21.8700 ;
      RECT 25.6960 20.7765 25.7220 21.8700 ;
      RECT 25.5880 20.7765 25.6140 21.8700 ;
      RECT 25.4800 20.7765 25.5060 21.8700 ;
      RECT 25.3720 20.7765 25.3980 21.8700 ;
      RECT 25.2640 20.7765 25.2900 21.8700 ;
      RECT 25.1560 20.7765 25.1820 21.8700 ;
      RECT 25.0480 20.7765 25.0740 21.8700 ;
      RECT 24.9400 20.7765 24.9660 21.8700 ;
      RECT 24.8320 20.7765 24.8580 21.8700 ;
      RECT 24.7240 20.7765 24.7500 21.8700 ;
      RECT 24.6160 20.7765 24.6420 21.8700 ;
      RECT 24.5080 20.7765 24.5340 21.8700 ;
      RECT 24.4000 20.7765 24.4260 21.8700 ;
      RECT 24.2920 20.7765 24.3180 21.8700 ;
      RECT 24.1840 20.7765 24.2100 21.8700 ;
      RECT 24.0760 20.7765 24.1020 21.8700 ;
      RECT 23.9680 20.7765 23.9940 21.8700 ;
      RECT 23.8600 20.7765 23.8860 21.8700 ;
      RECT 23.7520 20.7765 23.7780 21.8700 ;
      RECT 23.6440 20.7765 23.6700 21.8700 ;
      RECT 23.5360 20.7765 23.5620 21.8700 ;
      RECT 23.4280 20.7765 23.4540 21.8700 ;
      RECT 23.3200 20.7765 23.3460 21.8700 ;
      RECT 23.2120 20.7765 23.2380 21.8700 ;
      RECT 23.1040 20.7765 23.1300 21.8700 ;
      RECT 22.9960 20.7765 23.0220 21.8700 ;
      RECT 22.8880 20.7765 22.9140 21.8700 ;
      RECT 22.7800 20.7765 22.8060 21.8700 ;
      RECT 22.6720 20.7765 22.6980 21.8700 ;
      RECT 22.5640 20.7765 22.5900 21.8700 ;
      RECT 22.4560 20.7765 22.4820 21.8700 ;
      RECT 22.3480 20.7765 22.3740 21.8700 ;
      RECT 22.2400 20.7765 22.2660 21.8700 ;
      RECT 22.1320 20.7765 22.1580 21.8700 ;
      RECT 22.0240 20.7765 22.0500 21.8700 ;
      RECT 21.9160 20.7765 21.9420 21.8700 ;
      RECT 21.8080 20.7765 21.8340 21.8700 ;
      RECT 21.7000 20.7765 21.7260 21.8700 ;
      RECT 21.5920 20.7765 21.6180 21.8700 ;
      RECT 21.4840 20.7765 21.5100 21.8700 ;
      RECT 21.3760 20.7765 21.4020 21.8700 ;
      RECT 21.2680 20.7765 21.2940 21.8700 ;
      RECT 21.1600 20.7765 21.1860 21.8700 ;
      RECT 21.0520 20.7765 21.0780 21.8700 ;
      RECT 20.9440 20.7765 20.9700 21.8700 ;
      RECT 20.8360 20.7765 20.8620 21.8700 ;
      RECT 20.7280 20.7765 20.7540 21.8700 ;
      RECT 20.6200 20.7765 20.6460 21.8700 ;
      RECT 20.5120 20.7765 20.5380 21.8700 ;
      RECT 20.4040 20.7765 20.4300 21.8700 ;
      RECT 20.2960 20.7765 20.3220 21.8700 ;
      RECT 20.1880 20.7765 20.2140 21.8700 ;
      RECT 20.0800 20.7765 20.1060 21.8700 ;
      RECT 19.9720 20.7765 19.9980 21.8700 ;
      RECT 19.8640 20.7765 19.8900 21.8700 ;
      RECT 19.7560 20.7765 19.7820 21.8700 ;
      RECT 19.6480 20.7765 19.6740 21.8700 ;
      RECT 19.5400 20.7765 19.5660 21.8700 ;
      RECT 19.4320 20.7765 19.4580 21.8700 ;
      RECT 19.3240 20.7765 19.3500 21.8700 ;
      RECT 19.2160 20.7765 19.2420 21.8700 ;
      RECT 19.1080 20.7765 19.1340 21.8700 ;
      RECT 19.0000 20.7765 19.0260 21.8700 ;
      RECT 18.8920 20.7765 18.9180 21.8700 ;
      RECT 18.7840 20.7765 18.8100 21.8700 ;
      RECT 18.6760 20.7765 18.7020 21.8700 ;
      RECT 18.5680 20.7765 18.5940 21.8700 ;
      RECT 18.4600 20.7765 18.4860 21.8700 ;
      RECT 18.3520 20.7765 18.3780 21.8700 ;
      RECT 18.2440 20.7765 18.2700 21.8700 ;
      RECT 18.1360 20.7765 18.1620 21.8700 ;
      RECT 18.0280 20.7765 18.0540 21.8700 ;
      RECT 17.9200 20.7765 17.9460 21.8700 ;
      RECT 17.8120 20.7765 17.8380 21.8700 ;
      RECT 17.7040 20.7765 17.7300 21.8700 ;
      RECT 17.5960 20.7765 17.6220 21.8700 ;
      RECT 17.4880 20.7765 17.5140 21.8700 ;
      RECT 17.3800 20.7765 17.4060 21.8700 ;
      RECT 17.2720 20.7765 17.2980 21.8700 ;
      RECT 17.1640 20.7765 17.1900 21.8700 ;
      RECT 17.0560 20.7765 17.0820 21.8700 ;
      RECT 16.9480 20.7765 16.9740 21.8700 ;
      RECT 16.8400 20.7765 16.8660 21.8700 ;
      RECT 16.7320 20.7765 16.7580 21.8700 ;
      RECT 16.6240 20.7765 16.6500 21.8700 ;
      RECT 16.5160 20.7765 16.5420 21.8700 ;
      RECT 16.4080 20.7765 16.4340 21.8700 ;
      RECT 16.3000 20.7765 16.3260 21.8700 ;
      RECT 16.0870 20.7765 16.1640 21.8700 ;
      RECT 14.1940 20.7765 14.2710 21.8700 ;
      RECT 14.0320 20.7765 14.0580 21.8700 ;
      RECT 13.9240 20.7765 13.9500 21.8700 ;
      RECT 13.8160 20.7765 13.8420 21.8700 ;
      RECT 13.7080 20.7765 13.7340 21.8700 ;
      RECT 13.6000 20.7765 13.6260 21.8700 ;
      RECT 13.4920 20.7765 13.5180 21.8700 ;
      RECT 13.3840 20.7765 13.4100 21.8700 ;
      RECT 13.2760 20.7765 13.3020 21.8700 ;
      RECT 13.1680 20.7765 13.1940 21.8700 ;
      RECT 13.0600 20.7765 13.0860 21.8700 ;
      RECT 12.9520 20.7765 12.9780 21.8700 ;
      RECT 12.8440 20.7765 12.8700 21.8700 ;
      RECT 12.7360 20.7765 12.7620 21.8700 ;
      RECT 12.6280 20.7765 12.6540 21.8700 ;
      RECT 12.5200 20.7765 12.5460 21.8700 ;
      RECT 12.4120 20.7765 12.4380 21.8700 ;
      RECT 12.3040 20.7765 12.3300 21.8700 ;
      RECT 12.1960 20.7765 12.2220 21.8700 ;
      RECT 12.0880 20.7765 12.1140 21.8700 ;
      RECT 11.9800 20.7765 12.0060 21.8700 ;
      RECT 11.8720 20.7765 11.8980 21.8700 ;
      RECT 11.7640 20.7765 11.7900 21.8700 ;
      RECT 11.6560 20.7765 11.6820 21.8700 ;
      RECT 11.5480 20.7765 11.5740 21.8700 ;
      RECT 11.4400 20.7765 11.4660 21.8700 ;
      RECT 11.3320 20.7765 11.3580 21.8700 ;
      RECT 11.2240 20.7765 11.2500 21.8700 ;
      RECT 11.1160 20.7765 11.1420 21.8700 ;
      RECT 11.0080 20.7765 11.0340 21.8700 ;
      RECT 10.9000 20.7765 10.9260 21.8700 ;
      RECT 10.7920 20.7765 10.8180 21.8700 ;
      RECT 10.6840 20.7765 10.7100 21.8700 ;
      RECT 10.5760 20.7765 10.6020 21.8700 ;
      RECT 10.4680 20.7765 10.4940 21.8700 ;
      RECT 10.3600 20.7765 10.3860 21.8700 ;
      RECT 10.2520 20.7765 10.2780 21.8700 ;
      RECT 10.1440 20.7765 10.1700 21.8700 ;
      RECT 10.0360 20.7765 10.0620 21.8700 ;
      RECT 9.9280 20.7765 9.9540 21.8700 ;
      RECT 9.8200 20.7765 9.8460 21.8700 ;
      RECT 9.7120 20.7765 9.7380 21.8700 ;
      RECT 9.6040 20.7765 9.6300 21.8700 ;
      RECT 9.4960 20.7765 9.5220 21.8700 ;
      RECT 9.3880 20.7765 9.4140 21.8700 ;
      RECT 9.2800 20.7765 9.3060 21.8700 ;
      RECT 9.1720 20.7765 9.1980 21.8700 ;
      RECT 9.0640 20.7765 9.0900 21.8700 ;
      RECT 8.9560 20.7765 8.9820 21.8700 ;
      RECT 8.8480 20.7765 8.8740 21.8700 ;
      RECT 8.7400 20.7765 8.7660 21.8700 ;
      RECT 8.6320 20.7765 8.6580 21.8700 ;
      RECT 8.5240 20.7765 8.5500 21.8700 ;
      RECT 8.4160 20.7765 8.4420 21.8700 ;
      RECT 8.3080 20.7765 8.3340 21.8700 ;
      RECT 8.2000 20.7765 8.2260 21.8700 ;
      RECT 8.0920 20.7765 8.1180 21.8700 ;
      RECT 7.9840 20.7765 8.0100 21.8700 ;
      RECT 7.8760 20.7765 7.9020 21.8700 ;
      RECT 7.7680 20.7765 7.7940 21.8700 ;
      RECT 7.6600 20.7765 7.6860 21.8700 ;
      RECT 7.5520 20.7765 7.5780 21.8700 ;
      RECT 7.4440 20.7765 7.4700 21.8700 ;
      RECT 7.3360 20.7765 7.3620 21.8700 ;
      RECT 7.2280 20.7765 7.2540 21.8700 ;
      RECT 7.1200 20.7765 7.1460 21.8700 ;
      RECT 7.0120 20.7765 7.0380 21.8700 ;
      RECT 6.9040 20.7765 6.9300 21.8700 ;
      RECT 6.7960 20.7765 6.8220 21.8700 ;
      RECT 6.6880 20.7765 6.7140 21.8700 ;
      RECT 6.5800 20.7765 6.6060 21.8700 ;
      RECT 6.4720 20.7765 6.4980 21.8700 ;
      RECT 6.3640 20.7765 6.3900 21.8700 ;
      RECT 6.2560 20.7765 6.2820 21.8700 ;
      RECT 6.1480 20.7765 6.1740 21.8700 ;
      RECT 6.0400 20.7765 6.0660 21.8700 ;
      RECT 5.9320 20.7765 5.9580 21.8700 ;
      RECT 5.8240 20.7765 5.8500 21.8700 ;
      RECT 5.7160 20.7765 5.7420 21.8700 ;
      RECT 5.6080 20.7765 5.6340 21.8700 ;
      RECT 5.5000 20.7765 5.5260 21.8700 ;
      RECT 5.3920 20.7765 5.4180 21.8700 ;
      RECT 5.2840 20.7765 5.3100 21.8700 ;
      RECT 5.1760 20.7765 5.2020 21.8700 ;
      RECT 5.0680 20.7765 5.0940 21.8700 ;
      RECT 4.9600 20.7765 4.9860 21.8700 ;
      RECT 4.8520 20.7765 4.8780 21.8700 ;
      RECT 4.7440 20.7765 4.7700 21.8700 ;
      RECT 4.6360 20.7765 4.6620 21.8700 ;
      RECT 4.5280 20.7765 4.5540 21.8700 ;
      RECT 4.4200 20.7765 4.4460 21.8700 ;
      RECT 4.3120 20.7765 4.3380 21.8700 ;
      RECT 4.2040 20.7765 4.2300 21.8700 ;
      RECT 4.0960 20.7765 4.1220 21.8700 ;
      RECT 3.9880 20.7765 4.0140 21.8700 ;
      RECT 3.8800 20.7765 3.9060 21.8700 ;
      RECT 3.7720 20.7765 3.7980 21.8700 ;
      RECT 3.6640 20.7765 3.6900 21.8700 ;
      RECT 3.5560 20.7765 3.5820 21.8700 ;
      RECT 3.4480 20.7765 3.4740 21.8700 ;
      RECT 3.3400 20.7765 3.3660 21.8700 ;
      RECT 3.2320 20.7765 3.2580 21.8700 ;
      RECT 3.1240 20.7765 3.1500 21.8700 ;
      RECT 3.0160 20.7765 3.0420 21.8700 ;
      RECT 2.9080 20.7765 2.9340 21.8700 ;
      RECT 2.8000 20.7765 2.8260 21.8700 ;
      RECT 2.6920 20.7765 2.7180 21.8700 ;
      RECT 2.5840 20.7765 2.6100 21.8700 ;
      RECT 2.4760 20.7765 2.5020 21.8700 ;
      RECT 2.3680 20.7765 2.3940 21.8700 ;
      RECT 2.2600 20.7765 2.2860 21.8700 ;
      RECT 2.1520 20.7765 2.1780 21.8700 ;
      RECT 2.0440 20.7765 2.0700 21.8700 ;
      RECT 1.9360 20.7765 1.9620 21.8700 ;
      RECT 1.8280 20.7765 1.8540 21.8700 ;
      RECT 1.7200 20.7765 1.7460 21.8700 ;
      RECT 1.6120 20.7765 1.6380 21.8700 ;
      RECT 1.5040 20.7765 1.5300 21.8700 ;
      RECT 1.3960 20.7765 1.4220 21.8700 ;
      RECT 1.2880 20.7765 1.3140 21.8700 ;
      RECT 1.1800 20.7765 1.2060 21.8700 ;
      RECT 1.0720 20.7765 1.0980 21.8700 ;
      RECT 0.9640 20.7765 0.9900 21.8700 ;
      RECT 0.8560 20.7765 0.8820 21.8700 ;
      RECT 0.7480 20.7765 0.7740 21.8700 ;
      RECT 0.6400 20.7765 0.6660 21.8700 ;
      RECT 0.5320 20.7765 0.5580 21.8700 ;
      RECT 0.4240 20.7765 0.4500 21.8700 ;
      RECT 0.3160 20.7765 0.3420 21.8700 ;
      RECT 0.2080 20.7765 0.2340 21.8700 ;
      RECT 0.0050 20.7765 0.0900 21.8700 ;
      RECT 15.5530 21.8565 15.6810 22.9500 ;
      RECT 15.5390 22.5220 15.6810 22.8445 ;
      RECT 15.3190 22.2490 15.4530 22.9500 ;
      RECT 15.2960 22.5840 15.4530 22.8420 ;
      RECT 15.3190 21.8565 15.4170 22.9500 ;
      RECT 15.3190 21.9775 15.4310 22.2170 ;
      RECT 15.3190 21.8565 15.4530 21.9455 ;
      RECT 15.0940 22.3070 15.2280 22.9500 ;
      RECT 15.0940 21.8565 15.1920 22.9500 ;
      RECT 14.6770 21.8565 14.7600 22.9500 ;
      RECT 14.6770 21.9450 14.7740 22.8805 ;
      RECT 30.2680 21.8565 30.3530 22.9500 ;
      RECT 30.1240 21.8565 30.1500 22.9500 ;
      RECT 30.0160 21.8565 30.0420 22.9500 ;
      RECT 29.9080 21.8565 29.9340 22.9500 ;
      RECT 29.8000 21.8565 29.8260 22.9500 ;
      RECT 29.6920 21.8565 29.7180 22.9500 ;
      RECT 29.5840 21.8565 29.6100 22.9500 ;
      RECT 29.4760 21.8565 29.5020 22.9500 ;
      RECT 29.3680 21.8565 29.3940 22.9500 ;
      RECT 29.2600 21.8565 29.2860 22.9500 ;
      RECT 29.1520 21.8565 29.1780 22.9500 ;
      RECT 29.0440 21.8565 29.0700 22.9500 ;
      RECT 28.9360 21.8565 28.9620 22.9500 ;
      RECT 28.8280 21.8565 28.8540 22.9500 ;
      RECT 28.7200 21.8565 28.7460 22.9500 ;
      RECT 28.6120 21.8565 28.6380 22.9500 ;
      RECT 28.5040 21.8565 28.5300 22.9500 ;
      RECT 28.3960 21.8565 28.4220 22.9500 ;
      RECT 28.2880 21.8565 28.3140 22.9500 ;
      RECT 28.1800 21.8565 28.2060 22.9500 ;
      RECT 28.0720 21.8565 28.0980 22.9500 ;
      RECT 27.9640 21.8565 27.9900 22.9500 ;
      RECT 27.8560 21.8565 27.8820 22.9500 ;
      RECT 27.7480 21.8565 27.7740 22.9500 ;
      RECT 27.6400 21.8565 27.6660 22.9500 ;
      RECT 27.5320 21.8565 27.5580 22.9500 ;
      RECT 27.4240 21.8565 27.4500 22.9500 ;
      RECT 27.3160 21.8565 27.3420 22.9500 ;
      RECT 27.2080 21.8565 27.2340 22.9500 ;
      RECT 27.1000 21.8565 27.1260 22.9500 ;
      RECT 26.9920 21.8565 27.0180 22.9500 ;
      RECT 26.8840 21.8565 26.9100 22.9500 ;
      RECT 26.7760 21.8565 26.8020 22.9500 ;
      RECT 26.6680 21.8565 26.6940 22.9500 ;
      RECT 26.5600 21.8565 26.5860 22.9500 ;
      RECT 26.4520 21.8565 26.4780 22.9500 ;
      RECT 26.3440 21.8565 26.3700 22.9500 ;
      RECT 26.2360 21.8565 26.2620 22.9500 ;
      RECT 26.1280 21.8565 26.1540 22.9500 ;
      RECT 26.0200 21.8565 26.0460 22.9500 ;
      RECT 25.9120 21.8565 25.9380 22.9500 ;
      RECT 25.8040 21.8565 25.8300 22.9500 ;
      RECT 25.6960 21.8565 25.7220 22.9500 ;
      RECT 25.5880 21.8565 25.6140 22.9500 ;
      RECT 25.4800 21.8565 25.5060 22.9500 ;
      RECT 25.3720 21.8565 25.3980 22.9500 ;
      RECT 25.2640 21.8565 25.2900 22.9500 ;
      RECT 25.1560 21.8565 25.1820 22.9500 ;
      RECT 25.0480 21.8565 25.0740 22.9500 ;
      RECT 24.9400 21.8565 24.9660 22.9500 ;
      RECT 24.8320 21.8565 24.8580 22.9500 ;
      RECT 24.7240 21.8565 24.7500 22.9500 ;
      RECT 24.6160 21.8565 24.6420 22.9500 ;
      RECT 24.5080 21.8565 24.5340 22.9500 ;
      RECT 24.4000 21.8565 24.4260 22.9500 ;
      RECT 24.2920 21.8565 24.3180 22.9500 ;
      RECT 24.1840 21.8565 24.2100 22.9500 ;
      RECT 24.0760 21.8565 24.1020 22.9500 ;
      RECT 23.9680 21.8565 23.9940 22.9500 ;
      RECT 23.8600 21.8565 23.8860 22.9500 ;
      RECT 23.7520 21.8565 23.7780 22.9500 ;
      RECT 23.6440 21.8565 23.6700 22.9500 ;
      RECT 23.5360 21.8565 23.5620 22.9500 ;
      RECT 23.4280 21.8565 23.4540 22.9500 ;
      RECT 23.3200 21.8565 23.3460 22.9500 ;
      RECT 23.2120 21.8565 23.2380 22.9500 ;
      RECT 23.1040 21.8565 23.1300 22.9500 ;
      RECT 22.9960 21.8565 23.0220 22.9500 ;
      RECT 22.8880 21.8565 22.9140 22.9500 ;
      RECT 22.7800 21.8565 22.8060 22.9500 ;
      RECT 22.6720 21.8565 22.6980 22.9500 ;
      RECT 22.5640 21.8565 22.5900 22.9500 ;
      RECT 22.4560 21.8565 22.4820 22.9500 ;
      RECT 22.3480 21.8565 22.3740 22.9500 ;
      RECT 22.2400 21.8565 22.2660 22.9500 ;
      RECT 22.1320 21.8565 22.1580 22.9500 ;
      RECT 22.0240 21.8565 22.0500 22.9500 ;
      RECT 21.9160 21.8565 21.9420 22.9500 ;
      RECT 21.8080 21.8565 21.8340 22.9500 ;
      RECT 21.7000 21.8565 21.7260 22.9500 ;
      RECT 21.5920 21.8565 21.6180 22.9500 ;
      RECT 21.4840 21.8565 21.5100 22.9500 ;
      RECT 21.3760 21.8565 21.4020 22.9500 ;
      RECT 21.2680 21.8565 21.2940 22.9500 ;
      RECT 21.1600 21.8565 21.1860 22.9500 ;
      RECT 21.0520 21.8565 21.0780 22.9500 ;
      RECT 20.9440 21.8565 20.9700 22.9500 ;
      RECT 20.8360 21.8565 20.8620 22.9500 ;
      RECT 20.7280 21.8565 20.7540 22.9500 ;
      RECT 20.6200 21.8565 20.6460 22.9500 ;
      RECT 20.5120 21.8565 20.5380 22.9500 ;
      RECT 20.4040 21.8565 20.4300 22.9500 ;
      RECT 20.2960 21.8565 20.3220 22.9500 ;
      RECT 20.1880 21.8565 20.2140 22.9500 ;
      RECT 20.0800 21.8565 20.1060 22.9500 ;
      RECT 19.9720 21.8565 19.9980 22.9500 ;
      RECT 19.8640 21.8565 19.8900 22.9500 ;
      RECT 19.7560 21.8565 19.7820 22.9500 ;
      RECT 19.6480 21.8565 19.6740 22.9500 ;
      RECT 19.5400 21.8565 19.5660 22.9500 ;
      RECT 19.4320 21.8565 19.4580 22.9500 ;
      RECT 19.3240 21.8565 19.3500 22.9500 ;
      RECT 19.2160 21.8565 19.2420 22.9500 ;
      RECT 19.1080 21.8565 19.1340 22.9500 ;
      RECT 19.0000 21.8565 19.0260 22.9500 ;
      RECT 18.8920 21.8565 18.9180 22.9500 ;
      RECT 18.7840 21.8565 18.8100 22.9500 ;
      RECT 18.6760 21.8565 18.7020 22.9500 ;
      RECT 18.5680 21.8565 18.5940 22.9500 ;
      RECT 18.4600 21.8565 18.4860 22.9500 ;
      RECT 18.3520 21.8565 18.3780 22.9500 ;
      RECT 18.2440 21.8565 18.2700 22.9500 ;
      RECT 18.1360 21.8565 18.1620 22.9500 ;
      RECT 18.0280 21.8565 18.0540 22.9500 ;
      RECT 17.9200 21.8565 17.9460 22.9500 ;
      RECT 17.8120 21.8565 17.8380 22.9500 ;
      RECT 17.7040 21.8565 17.7300 22.9500 ;
      RECT 17.5960 21.8565 17.6220 22.9500 ;
      RECT 17.4880 21.8565 17.5140 22.9500 ;
      RECT 17.3800 21.8565 17.4060 22.9500 ;
      RECT 17.2720 21.8565 17.2980 22.9500 ;
      RECT 17.1640 21.8565 17.1900 22.9500 ;
      RECT 17.0560 21.8565 17.0820 22.9500 ;
      RECT 16.9480 21.8565 16.9740 22.9500 ;
      RECT 16.8400 21.8565 16.8660 22.9500 ;
      RECT 16.7320 21.8565 16.7580 22.9500 ;
      RECT 16.6240 21.8565 16.6500 22.9500 ;
      RECT 16.5160 21.8565 16.5420 22.9500 ;
      RECT 16.4080 21.8565 16.4340 22.9500 ;
      RECT 16.3000 21.8565 16.3260 22.9500 ;
      RECT 16.0870 21.8565 16.1640 22.9500 ;
      RECT 14.1940 21.8565 14.2710 22.9500 ;
      RECT 14.0320 21.8565 14.0580 22.9500 ;
      RECT 13.9240 21.8565 13.9500 22.9500 ;
      RECT 13.8160 21.8565 13.8420 22.9500 ;
      RECT 13.7080 21.8565 13.7340 22.9500 ;
      RECT 13.6000 21.8565 13.6260 22.9500 ;
      RECT 13.4920 21.8565 13.5180 22.9500 ;
      RECT 13.3840 21.8565 13.4100 22.9500 ;
      RECT 13.2760 21.8565 13.3020 22.9500 ;
      RECT 13.1680 21.8565 13.1940 22.9500 ;
      RECT 13.0600 21.8565 13.0860 22.9500 ;
      RECT 12.9520 21.8565 12.9780 22.9500 ;
      RECT 12.8440 21.8565 12.8700 22.9500 ;
      RECT 12.7360 21.8565 12.7620 22.9500 ;
      RECT 12.6280 21.8565 12.6540 22.9500 ;
      RECT 12.5200 21.8565 12.5460 22.9500 ;
      RECT 12.4120 21.8565 12.4380 22.9500 ;
      RECT 12.3040 21.8565 12.3300 22.9500 ;
      RECT 12.1960 21.8565 12.2220 22.9500 ;
      RECT 12.0880 21.8565 12.1140 22.9500 ;
      RECT 11.9800 21.8565 12.0060 22.9500 ;
      RECT 11.8720 21.8565 11.8980 22.9500 ;
      RECT 11.7640 21.8565 11.7900 22.9500 ;
      RECT 11.6560 21.8565 11.6820 22.9500 ;
      RECT 11.5480 21.8565 11.5740 22.9500 ;
      RECT 11.4400 21.8565 11.4660 22.9500 ;
      RECT 11.3320 21.8565 11.3580 22.9500 ;
      RECT 11.2240 21.8565 11.2500 22.9500 ;
      RECT 11.1160 21.8565 11.1420 22.9500 ;
      RECT 11.0080 21.8565 11.0340 22.9500 ;
      RECT 10.9000 21.8565 10.9260 22.9500 ;
      RECT 10.7920 21.8565 10.8180 22.9500 ;
      RECT 10.6840 21.8565 10.7100 22.9500 ;
      RECT 10.5760 21.8565 10.6020 22.9500 ;
      RECT 10.4680 21.8565 10.4940 22.9500 ;
      RECT 10.3600 21.8565 10.3860 22.9500 ;
      RECT 10.2520 21.8565 10.2780 22.9500 ;
      RECT 10.1440 21.8565 10.1700 22.9500 ;
      RECT 10.0360 21.8565 10.0620 22.9500 ;
      RECT 9.9280 21.8565 9.9540 22.9500 ;
      RECT 9.8200 21.8565 9.8460 22.9500 ;
      RECT 9.7120 21.8565 9.7380 22.9500 ;
      RECT 9.6040 21.8565 9.6300 22.9500 ;
      RECT 9.4960 21.8565 9.5220 22.9500 ;
      RECT 9.3880 21.8565 9.4140 22.9500 ;
      RECT 9.2800 21.8565 9.3060 22.9500 ;
      RECT 9.1720 21.8565 9.1980 22.9500 ;
      RECT 9.0640 21.8565 9.0900 22.9500 ;
      RECT 8.9560 21.8565 8.9820 22.9500 ;
      RECT 8.8480 21.8565 8.8740 22.9500 ;
      RECT 8.7400 21.8565 8.7660 22.9500 ;
      RECT 8.6320 21.8565 8.6580 22.9500 ;
      RECT 8.5240 21.8565 8.5500 22.9500 ;
      RECT 8.4160 21.8565 8.4420 22.9500 ;
      RECT 8.3080 21.8565 8.3340 22.9500 ;
      RECT 8.2000 21.8565 8.2260 22.9500 ;
      RECT 8.0920 21.8565 8.1180 22.9500 ;
      RECT 7.9840 21.8565 8.0100 22.9500 ;
      RECT 7.8760 21.8565 7.9020 22.9500 ;
      RECT 7.7680 21.8565 7.7940 22.9500 ;
      RECT 7.6600 21.8565 7.6860 22.9500 ;
      RECT 7.5520 21.8565 7.5780 22.9500 ;
      RECT 7.4440 21.8565 7.4700 22.9500 ;
      RECT 7.3360 21.8565 7.3620 22.9500 ;
      RECT 7.2280 21.8565 7.2540 22.9500 ;
      RECT 7.1200 21.8565 7.1460 22.9500 ;
      RECT 7.0120 21.8565 7.0380 22.9500 ;
      RECT 6.9040 21.8565 6.9300 22.9500 ;
      RECT 6.7960 21.8565 6.8220 22.9500 ;
      RECT 6.6880 21.8565 6.7140 22.9500 ;
      RECT 6.5800 21.8565 6.6060 22.9500 ;
      RECT 6.4720 21.8565 6.4980 22.9500 ;
      RECT 6.3640 21.8565 6.3900 22.9500 ;
      RECT 6.2560 21.8565 6.2820 22.9500 ;
      RECT 6.1480 21.8565 6.1740 22.9500 ;
      RECT 6.0400 21.8565 6.0660 22.9500 ;
      RECT 5.9320 21.8565 5.9580 22.9500 ;
      RECT 5.8240 21.8565 5.8500 22.9500 ;
      RECT 5.7160 21.8565 5.7420 22.9500 ;
      RECT 5.6080 21.8565 5.6340 22.9500 ;
      RECT 5.5000 21.8565 5.5260 22.9500 ;
      RECT 5.3920 21.8565 5.4180 22.9500 ;
      RECT 5.2840 21.8565 5.3100 22.9500 ;
      RECT 5.1760 21.8565 5.2020 22.9500 ;
      RECT 5.0680 21.8565 5.0940 22.9500 ;
      RECT 4.9600 21.8565 4.9860 22.9500 ;
      RECT 4.8520 21.8565 4.8780 22.9500 ;
      RECT 4.7440 21.8565 4.7700 22.9500 ;
      RECT 4.6360 21.8565 4.6620 22.9500 ;
      RECT 4.5280 21.8565 4.5540 22.9500 ;
      RECT 4.4200 21.8565 4.4460 22.9500 ;
      RECT 4.3120 21.8565 4.3380 22.9500 ;
      RECT 4.2040 21.8565 4.2300 22.9500 ;
      RECT 4.0960 21.8565 4.1220 22.9500 ;
      RECT 3.9880 21.8565 4.0140 22.9500 ;
      RECT 3.8800 21.8565 3.9060 22.9500 ;
      RECT 3.7720 21.8565 3.7980 22.9500 ;
      RECT 3.6640 21.8565 3.6900 22.9500 ;
      RECT 3.5560 21.8565 3.5820 22.9500 ;
      RECT 3.4480 21.8565 3.4740 22.9500 ;
      RECT 3.3400 21.8565 3.3660 22.9500 ;
      RECT 3.2320 21.8565 3.2580 22.9500 ;
      RECT 3.1240 21.8565 3.1500 22.9500 ;
      RECT 3.0160 21.8565 3.0420 22.9500 ;
      RECT 2.9080 21.8565 2.9340 22.9500 ;
      RECT 2.8000 21.8565 2.8260 22.9500 ;
      RECT 2.6920 21.8565 2.7180 22.9500 ;
      RECT 2.5840 21.8565 2.6100 22.9500 ;
      RECT 2.4760 21.8565 2.5020 22.9500 ;
      RECT 2.3680 21.8565 2.3940 22.9500 ;
      RECT 2.2600 21.8565 2.2860 22.9500 ;
      RECT 2.1520 21.8565 2.1780 22.9500 ;
      RECT 2.0440 21.8565 2.0700 22.9500 ;
      RECT 1.9360 21.8565 1.9620 22.9500 ;
      RECT 1.8280 21.8565 1.8540 22.9500 ;
      RECT 1.7200 21.8565 1.7460 22.9500 ;
      RECT 1.6120 21.8565 1.6380 22.9500 ;
      RECT 1.5040 21.8565 1.5300 22.9500 ;
      RECT 1.3960 21.8565 1.4220 22.9500 ;
      RECT 1.2880 21.8565 1.3140 22.9500 ;
      RECT 1.1800 21.8565 1.2060 22.9500 ;
      RECT 1.0720 21.8565 1.0980 22.9500 ;
      RECT 0.9640 21.8565 0.9900 22.9500 ;
      RECT 0.8560 21.8565 0.8820 22.9500 ;
      RECT 0.7480 21.8565 0.7740 22.9500 ;
      RECT 0.6400 21.8565 0.6660 22.9500 ;
      RECT 0.5320 21.8565 0.5580 22.9500 ;
      RECT 0.4240 21.8565 0.4500 22.9500 ;
      RECT 0.3160 21.8565 0.3420 22.9500 ;
      RECT 0.2080 21.8565 0.2340 22.9500 ;
      RECT 0.0050 21.8565 0.0900 22.9500 ;
      RECT 15.5530 22.9365 15.6810 24.0300 ;
      RECT 15.5390 23.6020 15.6810 23.9245 ;
      RECT 15.3190 23.3290 15.4530 24.0300 ;
      RECT 15.2960 23.6640 15.4530 23.9220 ;
      RECT 15.3190 22.9365 15.4170 24.0300 ;
      RECT 15.3190 23.0575 15.4310 23.2970 ;
      RECT 15.3190 22.9365 15.4530 23.0255 ;
      RECT 15.0940 23.3870 15.2280 24.0300 ;
      RECT 15.0940 22.9365 15.1920 24.0300 ;
      RECT 14.6770 22.9365 14.7600 24.0300 ;
      RECT 14.6770 23.0250 14.7740 23.9605 ;
      RECT 30.2680 22.9365 30.3530 24.0300 ;
      RECT 30.1240 22.9365 30.1500 24.0300 ;
      RECT 30.0160 22.9365 30.0420 24.0300 ;
      RECT 29.9080 22.9365 29.9340 24.0300 ;
      RECT 29.8000 22.9365 29.8260 24.0300 ;
      RECT 29.6920 22.9365 29.7180 24.0300 ;
      RECT 29.5840 22.9365 29.6100 24.0300 ;
      RECT 29.4760 22.9365 29.5020 24.0300 ;
      RECT 29.3680 22.9365 29.3940 24.0300 ;
      RECT 29.2600 22.9365 29.2860 24.0300 ;
      RECT 29.1520 22.9365 29.1780 24.0300 ;
      RECT 29.0440 22.9365 29.0700 24.0300 ;
      RECT 28.9360 22.9365 28.9620 24.0300 ;
      RECT 28.8280 22.9365 28.8540 24.0300 ;
      RECT 28.7200 22.9365 28.7460 24.0300 ;
      RECT 28.6120 22.9365 28.6380 24.0300 ;
      RECT 28.5040 22.9365 28.5300 24.0300 ;
      RECT 28.3960 22.9365 28.4220 24.0300 ;
      RECT 28.2880 22.9365 28.3140 24.0300 ;
      RECT 28.1800 22.9365 28.2060 24.0300 ;
      RECT 28.0720 22.9365 28.0980 24.0300 ;
      RECT 27.9640 22.9365 27.9900 24.0300 ;
      RECT 27.8560 22.9365 27.8820 24.0300 ;
      RECT 27.7480 22.9365 27.7740 24.0300 ;
      RECT 27.6400 22.9365 27.6660 24.0300 ;
      RECT 27.5320 22.9365 27.5580 24.0300 ;
      RECT 27.4240 22.9365 27.4500 24.0300 ;
      RECT 27.3160 22.9365 27.3420 24.0300 ;
      RECT 27.2080 22.9365 27.2340 24.0300 ;
      RECT 27.1000 22.9365 27.1260 24.0300 ;
      RECT 26.9920 22.9365 27.0180 24.0300 ;
      RECT 26.8840 22.9365 26.9100 24.0300 ;
      RECT 26.7760 22.9365 26.8020 24.0300 ;
      RECT 26.6680 22.9365 26.6940 24.0300 ;
      RECT 26.5600 22.9365 26.5860 24.0300 ;
      RECT 26.4520 22.9365 26.4780 24.0300 ;
      RECT 26.3440 22.9365 26.3700 24.0300 ;
      RECT 26.2360 22.9365 26.2620 24.0300 ;
      RECT 26.1280 22.9365 26.1540 24.0300 ;
      RECT 26.0200 22.9365 26.0460 24.0300 ;
      RECT 25.9120 22.9365 25.9380 24.0300 ;
      RECT 25.8040 22.9365 25.8300 24.0300 ;
      RECT 25.6960 22.9365 25.7220 24.0300 ;
      RECT 25.5880 22.9365 25.6140 24.0300 ;
      RECT 25.4800 22.9365 25.5060 24.0300 ;
      RECT 25.3720 22.9365 25.3980 24.0300 ;
      RECT 25.2640 22.9365 25.2900 24.0300 ;
      RECT 25.1560 22.9365 25.1820 24.0300 ;
      RECT 25.0480 22.9365 25.0740 24.0300 ;
      RECT 24.9400 22.9365 24.9660 24.0300 ;
      RECT 24.8320 22.9365 24.8580 24.0300 ;
      RECT 24.7240 22.9365 24.7500 24.0300 ;
      RECT 24.6160 22.9365 24.6420 24.0300 ;
      RECT 24.5080 22.9365 24.5340 24.0300 ;
      RECT 24.4000 22.9365 24.4260 24.0300 ;
      RECT 24.2920 22.9365 24.3180 24.0300 ;
      RECT 24.1840 22.9365 24.2100 24.0300 ;
      RECT 24.0760 22.9365 24.1020 24.0300 ;
      RECT 23.9680 22.9365 23.9940 24.0300 ;
      RECT 23.8600 22.9365 23.8860 24.0300 ;
      RECT 23.7520 22.9365 23.7780 24.0300 ;
      RECT 23.6440 22.9365 23.6700 24.0300 ;
      RECT 23.5360 22.9365 23.5620 24.0300 ;
      RECT 23.4280 22.9365 23.4540 24.0300 ;
      RECT 23.3200 22.9365 23.3460 24.0300 ;
      RECT 23.2120 22.9365 23.2380 24.0300 ;
      RECT 23.1040 22.9365 23.1300 24.0300 ;
      RECT 22.9960 22.9365 23.0220 24.0300 ;
      RECT 22.8880 22.9365 22.9140 24.0300 ;
      RECT 22.7800 22.9365 22.8060 24.0300 ;
      RECT 22.6720 22.9365 22.6980 24.0300 ;
      RECT 22.5640 22.9365 22.5900 24.0300 ;
      RECT 22.4560 22.9365 22.4820 24.0300 ;
      RECT 22.3480 22.9365 22.3740 24.0300 ;
      RECT 22.2400 22.9365 22.2660 24.0300 ;
      RECT 22.1320 22.9365 22.1580 24.0300 ;
      RECT 22.0240 22.9365 22.0500 24.0300 ;
      RECT 21.9160 22.9365 21.9420 24.0300 ;
      RECT 21.8080 22.9365 21.8340 24.0300 ;
      RECT 21.7000 22.9365 21.7260 24.0300 ;
      RECT 21.5920 22.9365 21.6180 24.0300 ;
      RECT 21.4840 22.9365 21.5100 24.0300 ;
      RECT 21.3760 22.9365 21.4020 24.0300 ;
      RECT 21.2680 22.9365 21.2940 24.0300 ;
      RECT 21.1600 22.9365 21.1860 24.0300 ;
      RECT 21.0520 22.9365 21.0780 24.0300 ;
      RECT 20.9440 22.9365 20.9700 24.0300 ;
      RECT 20.8360 22.9365 20.8620 24.0300 ;
      RECT 20.7280 22.9365 20.7540 24.0300 ;
      RECT 20.6200 22.9365 20.6460 24.0300 ;
      RECT 20.5120 22.9365 20.5380 24.0300 ;
      RECT 20.4040 22.9365 20.4300 24.0300 ;
      RECT 20.2960 22.9365 20.3220 24.0300 ;
      RECT 20.1880 22.9365 20.2140 24.0300 ;
      RECT 20.0800 22.9365 20.1060 24.0300 ;
      RECT 19.9720 22.9365 19.9980 24.0300 ;
      RECT 19.8640 22.9365 19.8900 24.0300 ;
      RECT 19.7560 22.9365 19.7820 24.0300 ;
      RECT 19.6480 22.9365 19.6740 24.0300 ;
      RECT 19.5400 22.9365 19.5660 24.0300 ;
      RECT 19.4320 22.9365 19.4580 24.0300 ;
      RECT 19.3240 22.9365 19.3500 24.0300 ;
      RECT 19.2160 22.9365 19.2420 24.0300 ;
      RECT 19.1080 22.9365 19.1340 24.0300 ;
      RECT 19.0000 22.9365 19.0260 24.0300 ;
      RECT 18.8920 22.9365 18.9180 24.0300 ;
      RECT 18.7840 22.9365 18.8100 24.0300 ;
      RECT 18.6760 22.9365 18.7020 24.0300 ;
      RECT 18.5680 22.9365 18.5940 24.0300 ;
      RECT 18.4600 22.9365 18.4860 24.0300 ;
      RECT 18.3520 22.9365 18.3780 24.0300 ;
      RECT 18.2440 22.9365 18.2700 24.0300 ;
      RECT 18.1360 22.9365 18.1620 24.0300 ;
      RECT 18.0280 22.9365 18.0540 24.0300 ;
      RECT 17.9200 22.9365 17.9460 24.0300 ;
      RECT 17.8120 22.9365 17.8380 24.0300 ;
      RECT 17.7040 22.9365 17.7300 24.0300 ;
      RECT 17.5960 22.9365 17.6220 24.0300 ;
      RECT 17.4880 22.9365 17.5140 24.0300 ;
      RECT 17.3800 22.9365 17.4060 24.0300 ;
      RECT 17.2720 22.9365 17.2980 24.0300 ;
      RECT 17.1640 22.9365 17.1900 24.0300 ;
      RECT 17.0560 22.9365 17.0820 24.0300 ;
      RECT 16.9480 22.9365 16.9740 24.0300 ;
      RECT 16.8400 22.9365 16.8660 24.0300 ;
      RECT 16.7320 22.9365 16.7580 24.0300 ;
      RECT 16.6240 22.9365 16.6500 24.0300 ;
      RECT 16.5160 22.9365 16.5420 24.0300 ;
      RECT 16.4080 22.9365 16.4340 24.0300 ;
      RECT 16.3000 22.9365 16.3260 24.0300 ;
      RECT 16.0870 22.9365 16.1640 24.0300 ;
      RECT 14.1940 22.9365 14.2710 24.0300 ;
      RECT 14.0320 22.9365 14.0580 24.0300 ;
      RECT 13.9240 22.9365 13.9500 24.0300 ;
      RECT 13.8160 22.9365 13.8420 24.0300 ;
      RECT 13.7080 22.9365 13.7340 24.0300 ;
      RECT 13.6000 22.9365 13.6260 24.0300 ;
      RECT 13.4920 22.9365 13.5180 24.0300 ;
      RECT 13.3840 22.9365 13.4100 24.0300 ;
      RECT 13.2760 22.9365 13.3020 24.0300 ;
      RECT 13.1680 22.9365 13.1940 24.0300 ;
      RECT 13.0600 22.9365 13.0860 24.0300 ;
      RECT 12.9520 22.9365 12.9780 24.0300 ;
      RECT 12.8440 22.9365 12.8700 24.0300 ;
      RECT 12.7360 22.9365 12.7620 24.0300 ;
      RECT 12.6280 22.9365 12.6540 24.0300 ;
      RECT 12.5200 22.9365 12.5460 24.0300 ;
      RECT 12.4120 22.9365 12.4380 24.0300 ;
      RECT 12.3040 22.9365 12.3300 24.0300 ;
      RECT 12.1960 22.9365 12.2220 24.0300 ;
      RECT 12.0880 22.9365 12.1140 24.0300 ;
      RECT 11.9800 22.9365 12.0060 24.0300 ;
      RECT 11.8720 22.9365 11.8980 24.0300 ;
      RECT 11.7640 22.9365 11.7900 24.0300 ;
      RECT 11.6560 22.9365 11.6820 24.0300 ;
      RECT 11.5480 22.9365 11.5740 24.0300 ;
      RECT 11.4400 22.9365 11.4660 24.0300 ;
      RECT 11.3320 22.9365 11.3580 24.0300 ;
      RECT 11.2240 22.9365 11.2500 24.0300 ;
      RECT 11.1160 22.9365 11.1420 24.0300 ;
      RECT 11.0080 22.9365 11.0340 24.0300 ;
      RECT 10.9000 22.9365 10.9260 24.0300 ;
      RECT 10.7920 22.9365 10.8180 24.0300 ;
      RECT 10.6840 22.9365 10.7100 24.0300 ;
      RECT 10.5760 22.9365 10.6020 24.0300 ;
      RECT 10.4680 22.9365 10.4940 24.0300 ;
      RECT 10.3600 22.9365 10.3860 24.0300 ;
      RECT 10.2520 22.9365 10.2780 24.0300 ;
      RECT 10.1440 22.9365 10.1700 24.0300 ;
      RECT 10.0360 22.9365 10.0620 24.0300 ;
      RECT 9.9280 22.9365 9.9540 24.0300 ;
      RECT 9.8200 22.9365 9.8460 24.0300 ;
      RECT 9.7120 22.9365 9.7380 24.0300 ;
      RECT 9.6040 22.9365 9.6300 24.0300 ;
      RECT 9.4960 22.9365 9.5220 24.0300 ;
      RECT 9.3880 22.9365 9.4140 24.0300 ;
      RECT 9.2800 22.9365 9.3060 24.0300 ;
      RECT 9.1720 22.9365 9.1980 24.0300 ;
      RECT 9.0640 22.9365 9.0900 24.0300 ;
      RECT 8.9560 22.9365 8.9820 24.0300 ;
      RECT 8.8480 22.9365 8.8740 24.0300 ;
      RECT 8.7400 22.9365 8.7660 24.0300 ;
      RECT 8.6320 22.9365 8.6580 24.0300 ;
      RECT 8.5240 22.9365 8.5500 24.0300 ;
      RECT 8.4160 22.9365 8.4420 24.0300 ;
      RECT 8.3080 22.9365 8.3340 24.0300 ;
      RECT 8.2000 22.9365 8.2260 24.0300 ;
      RECT 8.0920 22.9365 8.1180 24.0300 ;
      RECT 7.9840 22.9365 8.0100 24.0300 ;
      RECT 7.8760 22.9365 7.9020 24.0300 ;
      RECT 7.7680 22.9365 7.7940 24.0300 ;
      RECT 7.6600 22.9365 7.6860 24.0300 ;
      RECT 7.5520 22.9365 7.5780 24.0300 ;
      RECT 7.4440 22.9365 7.4700 24.0300 ;
      RECT 7.3360 22.9365 7.3620 24.0300 ;
      RECT 7.2280 22.9365 7.2540 24.0300 ;
      RECT 7.1200 22.9365 7.1460 24.0300 ;
      RECT 7.0120 22.9365 7.0380 24.0300 ;
      RECT 6.9040 22.9365 6.9300 24.0300 ;
      RECT 6.7960 22.9365 6.8220 24.0300 ;
      RECT 6.6880 22.9365 6.7140 24.0300 ;
      RECT 6.5800 22.9365 6.6060 24.0300 ;
      RECT 6.4720 22.9365 6.4980 24.0300 ;
      RECT 6.3640 22.9365 6.3900 24.0300 ;
      RECT 6.2560 22.9365 6.2820 24.0300 ;
      RECT 6.1480 22.9365 6.1740 24.0300 ;
      RECT 6.0400 22.9365 6.0660 24.0300 ;
      RECT 5.9320 22.9365 5.9580 24.0300 ;
      RECT 5.8240 22.9365 5.8500 24.0300 ;
      RECT 5.7160 22.9365 5.7420 24.0300 ;
      RECT 5.6080 22.9365 5.6340 24.0300 ;
      RECT 5.5000 22.9365 5.5260 24.0300 ;
      RECT 5.3920 22.9365 5.4180 24.0300 ;
      RECT 5.2840 22.9365 5.3100 24.0300 ;
      RECT 5.1760 22.9365 5.2020 24.0300 ;
      RECT 5.0680 22.9365 5.0940 24.0300 ;
      RECT 4.9600 22.9365 4.9860 24.0300 ;
      RECT 4.8520 22.9365 4.8780 24.0300 ;
      RECT 4.7440 22.9365 4.7700 24.0300 ;
      RECT 4.6360 22.9365 4.6620 24.0300 ;
      RECT 4.5280 22.9365 4.5540 24.0300 ;
      RECT 4.4200 22.9365 4.4460 24.0300 ;
      RECT 4.3120 22.9365 4.3380 24.0300 ;
      RECT 4.2040 22.9365 4.2300 24.0300 ;
      RECT 4.0960 22.9365 4.1220 24.0300 ;
      RECT 3.9880 22.9365 4.0140 24.0300 ;
      RECT 3.8800 22.9365 3.9060 24.0300 ;
      RECT 3.7720 22.9365 3.7980 24.0300 ;
      RECT 3.6640 22.9365 3.6900 24.0300 ;
      RECT 3.5560 22.9365 3.5820 24.0300 ;
      RECT 3.4480 22.9365 3.4740 24.0300 ;
      RECT 3.3400 22.9365 3.3660 24.0300 ;
      RECT 3.2320 22.9365 3.2580 24.0300 ;
      RECT 3.1240 22.9365 3.1500 24.0300 ;
      RECT 3.0160 22.9365 3.0420 24.0300 ;
      RECT 2.9080 22.9365 2.9340 24.0300 ;
      RECT 2.8000 22.9365 2.8260 24.0300 ;
      RECT 2.6920 22.9365 2.7180 24.0300 ;
      RECT 2.5840 22.9365 2.6100 24.0300 ;
      RECT 2.4760 22.9365 2.5020 24.0300 ;
      RECT 2.3680 22.9365 2.3940 24.0300 ;
      RECT 2.2600 22.9365 2.2860 24.0300 ;
      RECT 2.1520 22.9365 2.1780 24.0300 ;
      RECT 2.0440 22.9365 2.0700 24.0300 ;
      RECT 1.9360 22.9365 1.9620 24.0300 ;
      RECT 1.8280 22.9365 1.8540 24.0300 ;
      RECT 1.7200 22.9365 1.7460 24.0300 ;
      RECT 1.6120 22.9365 1.6380 24.0300 ;
      RECT 1.5040 22.9365 1.5300 24.0300 ;
      RECT 1.3960 22.9365 1.4220 24.0300 ;
      RECT 1.2880 22.9365 1.3140 24.0300 ;
      RECT 1.1800 22.9365 1.2060 24.0300 ;
      RECT 1.0720 22.9365 1.0980 24.0300 ;
      RECT 0.9640 22.9365 0.9900 24.0300 ;
      RECT 0.8560 22.9365 0.8820 24.0300 ;
      RECT 0.7480 22.9365 0.7740 24.0300 ;
      RECT 0.6400 22.9365 0.6660 24.0300 ;
      RECT 0.5320 22.9365 0.5580 24.0300 ;
      RECT 0.4240 22.9365 0.4500 24.0300 ;
      RECT 0.3160 22.9365 0.3420 24.0300 ;
      RECT 0.2080 22.9365 0.2340 24.0300 ;
      RECT 0.0050 22.9365 0.0900 24.0300 ;
      RECT 15.5530 24.0165 15.6810 25.1100 ;
      RECT 15.5390 24.6820 15.6810 25.0045 ;
      RECT 15.3190 24.4090 15.4530 25.1100 ;
      RECT 15.2960 24.7440 15.4530 25.0020 ;
      RECT 15.3190 24.0165 15.4170 25.1100 ;
      RECT 15.3190 24.1375 15.4310 24.3770 ;
      RECT 15.3190 24.0165 15.4530 24.1055 ;
      RECT 15.0940 24.4670 15.2280 25.1100 ;
      RECT 15.0940 24.0165 15.1920 25.1100 ;
      RECT 14.6770 24.0165 14.7600 25.1100 ;
      RECT 14.6770 24.1050 14.7740 25.0405 ;
      RECT 30.2680 24.0165 30.3530 25.1100 ;
      RECT 30.1240 24.0165 30.1500 25.1100 ;
      RECT 30.0160 24.0165 30.0420 25.1100 ;
      RECT 29.9080 24.0165 29.9340 25.1100 ;
      RECT 29.8000 24.0165 29.8260 25.1100 ;
      RECT 29.6920 24.0165 29.7180 25.1100 ;
      RECT 29.5840 24.0165 29.6100 25.1100 ;
      RECT 29.4760 24.0165 29.5020 25.1100 ;
      RECT 29.3680 24.0165 29.3940 25.1100 ;
      RECT 29.2600 24.0165 29.2860 25.1100 ;
      RECT 29.1520 24.0165 29.1780 25.1100 ;
      RECT 29.0440 24.0165 29.0700 25.1100 ;
      RECT 28.9360 24.0165 28.9620 25.1100 ;
      RECT 28.8280 24.0165 28.8540 25.1100 ;
      RECT 28.7200 24.0165 28.7460 25.1100 ;
      RECT 28.6120 24.0165 28.6380 25.1100 ;
      RECT 28.5040 24.0165 28.5300 25.1100 ;
      RECT 28.3960 24.0165 28.4220 25.1100 ;
      RECT 28.2880 24.0165 28.3140 25.1100 ;
      RECT 28.1800 24.0165 28.2060 25.1100 ;
      RECT 28.0720 24.0165 28.0980 25.1100 ;
      RECT 27.9640 24.0165 27.9900 25.1100 ;
      RECT 27.8560 24.0165 27.8820 25.1100 ;
      RECT 27.7480 24.0165 27.7740 25.1100 ;
      RECT 27.6400 24.0165 27.6660 25.1100 ;
      RECT 27.5320 24.0165 27.5580 25.1100 ;
      RECT 27.4240 24.0165 27.4500 25.1100 ;
      RECT 27.3160 24.0165 27.3420 25.1100 ;
      RECT 27.2080 24.0165 27.2340 25.1100 ;
      RECT 27.1000 24.0165 27.1260 25.1100 ;
      RECT 26.9920 24.0165 27.0180 25.1100 ;
      RECT 26.8840 24.0165 26.9100 25.1100 ;
      RECT 26.7760 24.0165 26.8020 25.1100 ;
      RECT 26.6680 24.0165 26.6940 25.1100 ;
      RECT 26.5600 24.0165 26.5860 25.1100 ;
      RECT 26.4520 24.0165 26.4780 25.1100 ;
      RECT 26.3440 24.0165 26.3700 25.1100 ;
      RECT 26.2360 24.0165 26.2620 25.1100 ;
      RECT 26.1280 24.0165 26.1540 25.1100 ;
      RECT 26.0200 24.0165 26.0460 25.1100 ;
      RECT 25.9120 24.0165 25.9380 25.1100 ;
      RECT 25.8040 24.0165 25.8300 25.1100 ;
      RECT 25.6960 24.0165 25.7220 25.1100 ;
      RECT 25.5880 24.0165 25.6140 25.1100 ;
      RECT 25.4800 24.0165 25.5060 25.1100 ;
      RECT 25.3720 24.0165 25.3980 25.1100 ;
      RECT 25.2640 24.0165 25.2900 25.1100 ;
      RECT 25.1560 24.0165 25.1820 25.1100 ;
      RECT 25.0480 24.0165 25.0740 25.1100 ;
      RECT 24.9400 24.0165 24.9660 25.1100 ;
      RECT 24.8320 24.0165 24.8580 25.1100 ;
      RECT 24.7240 24.0165 24.7500 25.1100 ;
      RECT 24.6160 24.0165 24.6420 25.1100 ;
      RECT 24.5080 24.0165 24.5340 25.1100 ;
      RECT 24.4000 24.0165 24.4260 25.1100 ;
      RECT 24.2920 24.0165 24.3180 25.1100 ;
      RECT 24.1840 24.0165 24.2100 25.1100 ;
      RECT 24.0760 24.0165 24.1020 25.1100 ;
      RECT 23.9680 24.0165 23.9940 25.1100 ;
      RECT 23.8600 24.0165 23.8860 25.1100 ;
      RECT 23.7520 24.0165 23.7780 25.1100 ;
      RECT 23.6440 24.0165 23.6700 25.1100 ;
      RECT 23.5360 24.0165 23.5620 25.1100 ;
      RECT 23.4280 24.0165 23.4540 25.1100 ;
      RECT 23.3200 24.0165 23.3460 25.1100 ;
      RECT 23.2120 24.0165 23.2380 25.1100 ;
      RECT 23.1040 24.0165 23.1300 25.1100 ;
      RECT 22.9960 24.0165 23.0220 25.1100 ;
      RECT 22.8880 24.0165 22.9140 25.1100 ;
      RECT 22.7800 24.0165 22.8060 25.1100 ;
      RECT 22.6720 24.0165 22.6980 25.1100 ;
      RECT 22.5640 24.0165 22.5900 25.1100 ;
      RECT 22.4560 24.0165 22.4820 25.1100 ;
      RECT 22.3480 24.0165 22.3740 25.1100 ;
      RECT 22.2400 24.0165 22.2660 25.1100 ;
      RECT 22.1320 24.0165 22.1580 25.1100 ;
      RECT 22.0240 24.0165 22.0500 25.1100 ;
      RECT 21.9160 24.0165 21.9420 25.1100 ;
      RECT 21.8080 24.0165 21.8340 25.1100 ;
      RECT 21.7000 24.0165 21.7260 25.1100 ;
      RECT 21.5920 24.0165 21.6180 25.1100 ;
      RECT 21.4840 24.0165 21.5100 25.1100 ;
      RECT 21.3760 24.0165 21.4020 25.1100 ;
      RECT 21.2680 24.0165 21.2940 25.1100 ;
      RECT 21.1600 24.0165 21.1860 25.1100 ;
      RECT 21.0520 24.0165 21.0780 25.1100 ;
      RECT 20.9440 24.0165 20.9700 25.1100 ;
      RECT 20.8360 24.0165 20.8620 25.1100 ;
      RECT 20.7280 24.0165 20.7540 25.1100 ;
      RECT 20.6200 24.0165 20.6460 25.1100 ;
      RECT 20.5120 24.0165 20.5380 25.1100 ;
      RECT 20.4040 24.0165 20.4300 25.1100 ;
      RECT 20.2960 24.0165 20.3220 25.1100 ;
      RECT 20.1880 24.0165 20.2140 25.1100 ;
      RECT 20.0800 24.0165 20.1060 25.1100 ;
      RECT 19.9720 24.0165 19.9980 25.1100 ;
      RECT 19.8640 24.0165 19.8900 25.1100 ;
      RECT 19.7560 24.0165 19.7820 25.1100 ;
      RECT 19.6480 24.0165 19.6740 25.1100 ;
      RECT 19.5400 24.0165 19.5660 25.1100 ;
      RECT 19.4320 24.0165 19.4580 25.1100 ;
      RECT 19.3240 24.0165 19.3500 25.1100 ;
      RECT 19.2160 24.0165 19.2420 25.1100 ;
      RECT 19.1080 24.0165 19.1340 25.1100 ;
      RECT 19.0000 24.0165 19.0260 25.1100 ;
      RECT 18.8920 24.0165 18.9180 25.1100 ;
      RECT 18.7840 24.0165 18.8100 25.1100 ;
      RECT 18.6760 24.0165 18.7020 25.1100 ;
      RECT 18.5680 24.0165 18.5940 25.1100 ;
      RECT 18.4600 24.0165 18.4860 25.1100 ;
      RECT 18.3520 24.0165 18.3780 25.1100 ;
      RECT 18.2440 24.0165 18.2700 25.1100 ;
      RECT 18.1360 24.0165 18.1620 25.1100 ;
      RECT 18.0280 24.0165 18.0540 25.1100 ;
      RECT 17.9200 24.0165 17.9460 25.1100 ;
      RECT 17.8120 24.0165 17.8380 25.1100 ;
      RECT 17.7040 24.0165 17.7300 25.1100 ;
      RECT 17.5960 24.0165 17.6220 25.1100 ;
      RECT 17.4880 24.0165 17.5140 25.1100 ;
      RECT 17.3800 24.0165 17.4060 25.1100 ;
      RECT 17.2720 24.0165 17.2980 25.1100 ;
      RECT 17.1640 24.0165 17.1900 25.1100 ;
      RECT 17.0560 24.0165 17.0820 25.1100 ;
      RECT 16.9480 24.0165 16.9740 25.1100 ;
      RECT 16.8400 24.0165 16.8660 25.1100 ;
      RECT 16.7320 24.0165 16.7580 25.1100 ;
      RECT 16.6240 24.0165 16.6500 25.1100 ;
      RECT 16.5160 24.0165 16.5420 25.1100 ;
      RECT 16.4080 24.0165 16.4340 25.1100 ;
      RECT 16.3000 24.0165 16.3260 25.1100 ;
      RECT 16.0870 24.0165 16.1640 25.1100 ;
      RECT 14.1940 24.0165 14.2710 25.1100 ;
      RECT 14.0320 24.0165 14.0580 25.1100 ;
      RECT 13.9240 24.0165 13.9500 25.1100 ;
      RECT 13.8160 24.0165 13.8420 25.1100 ;
      RECT 13.7080 24.0165 13.7340 25.1100 ;
      RECT 13.6000 24.0165 13.6260 25.1100 ;
      RECT 13.4920 24.0165 13.5180 25.1100 ;
      RECT 13.3840 24.0165 13.4100 25.1100 ;
      RECT 13.2760 24.0165 13.3020 25.1100 ;
      RECT 13.1680 24.0165 13.1940 25.1100 ;
      RECT 13.0600 24.0165 13.0860 25.1100 ;
      RECT 12.9520 24.0165 12.9780 25.1100 ;
      RECT 12.8440 24.0165 12.8700 25.1100 ;
      RECT 12.7360 24.0165 12.7620 25.1100 ;
      RECT 12.6280 24.0165 12.6540 25.1100 ;
      RECT 12.5200 24.0165 12.5460 25.1100 ;
      RECT 12.4120 24.0165 12.4380 25.1100 ;
      RECT 12.3040 24.0165 12.3300 25.1100 ;
      RECT 12.1960 24.0165 12.2220 25.1100 ;
      RECT 12.0880 24.0165 12.1140 25.1100 ;
      RECT 11.9800 24.0165 12.0060 25.1100 ;
      RECT 11.8720 24.0165 11.8980 25.1100 ;
      RECT 11.7640 24.0165 11.7900 25.1100 ;
      RECT 11.6560 24.0165 11.6820 25.1100 ;
      RECT 11.5480 24.0165 11.5740 25.1100 ;
      RECT 11.4400 24.0165 11.4660 25.1100 ;
      RECT 11.3320 24.0165 11.3580 25.1100 ;
      RECT 11.2240 24.0165 11.2500 25.1100 ;
      RECT 11.1160 24.0165 11.1420 25.1100 ;
      RECT 11.0080 24.0165 11.0340 25.1100 ;
      RECT 10.9000 24.0165 10.9260 25.1100 ;
      RECT 10.7920 24.0165 10.8180 25.1100 ;
      RECT 10.6840 24.0165 10.7100 25.1100 ;
      RECT 10.5760 24.0165 10.6020 25.1100 ;
      RECT 10.4680 24.0165 10.4940 25.1100 ;
      RECT 10.3600 24.0165 10.3860 25.1100 ;
      RECT 10.2520 24.0165 10.2780 25.1100 ;
      RECT 10.1440 24.0165 10.1700 25.1100 ;
      RECT 10.0360 24.0165 10.0620 25.1100 ;
      RECT 9.9280 24.0165 9.9540 25.1100 ;
      RECT 9.8200 24.0165 9.8460 25.1100 ;
      RECT 9.7120 24.0165 9.7380 25.1100 ;
      RECT 9.6040 24.0165 9.6300 25.1100 ;
      RECT 9.4960 24.0165 9.5220 25.1100 ;
      RECT 9.3880 24.0165 9.4140 25.1100 ;
      RECT 9.2800 24.0165 9.3060 25.1100 ;
      RECT 9.1720 24.0165 9.1980 25.1100 ;
      RECT 9.0640 24.0165 9.0900 25.1100 ;
      RECT 8.9560 24.0165 8.9820 25.1100 ;
      RECT 8.8480 24.0165 8.8740 25.1100 ;
      RECT 8.7400 24.0165 8.7660 25.1100 ;
      RECT 8.6320 24.0165 8.6580 25.1100 ;
      RECT 8.5240 24.0165 8.5500 25.1100 ;
      RECT 8.4160 24.0165 8.4420 25.1100 ;
      RECT 8.3080 24.0165 8.3340 25.1100 ;
      RECT 8.2000 24.0165 8.2260 25.1100 ;
      RECT 8.0920 24.0165 8.1180 25.1100 ;
      RECT 7.9840 24.0165 8.0100 25.1100 ;
      RECT 7.8760 24.0165 7.9020 25.1100 ;
      RECT 7.7680 24.0165 7.7940 25.1100 ;
      RECT 7.6600 24.0165 7.6860 25.1100 ;
      RECT 7.5520 24.0165 7.5780 25.1100 ;
      RECT 7.4440 24.0165 7.4700 25.1100 ;
      RECT 7.3360 24.0165 7.3620 25.1100 ;
      RECT 7.2280 24.0165 7.2540 25.1100 ;
      RECT 7.1200 24.0165 7.1460 25.1100 ;
      RECT 7.0120 24.0165 7.0380 25.1100 ;
      RECT 6.9040 24.0165 6.9300 25.1100 ;
      RECT 6.7960 24.0165 6.8220 25.1100 ;
      RECT 6.6880 24.0165 6.7140 25.1100 ;
      RECT 6.5800 24.0165 6.6060 25.1100 ;
      RECT 6.4720 24.0165 6.4980 25.1100 ;
      RECT 6.3640 24.0165 6.3900 25.1100 ;
      RECT 6.2560 24.0165 6.2820 25.1100 ;
      RECT 6.1480 24.0165 6.1740 25.1100 ;
      RECT 6.0400 24.0165 6.0660 25.1100 ;
      RECT 5.9320 24.0165 5.9580 25.1100 ;
      RECT 5.8240 24.0165 5.8500 25.1100 ;
      RECT 5.7160 24.0165 5.7420 25.1100 ;
      RECT 5.6080 24.0165 5.6340 25.1100 ;
      RECT 5.5000 24.0165 5.5260 25.1100 ;
      RECT 5.3920 24.0165 5.4180 25.1100 ;
      RECT 5.2840 24.0165 5.3100 25.1100 ;
      RECT 5.1760 24.0165 5.2020 25.1100 ;
      RECT 5.0680 24.0165 5.0940 25.1100 ;
      RECT 4.9600 24.0165 4.9860 25.1100 ;
      RECT 4.8520 24.0165 4.8780 25.1100 ;
      RECT 4.7440 24.0165 4.7700 25.1100 ;
      RECT 4.6360 24.0165 4.6620 25.1100 ;
      RECT 4.5280 24.0165 4.5540 25.1100 ;
      RECT 4.4200 24.0165 4.4460 25.1100 ;
      RECT 4.3120 24.0165 4.3380 25.1100 ;
      RECT 4.2040 24.0165 4.2300 25.1100 ;
      RECT 4.0960 24.0165 4.1220 25.1100 ;
      RECT 3.9880 24.0165 4.0140 25.1100 ;
      RECT 3.8800 24.0165 3.9060 25.1100 ;
      RECT 3.7720 24.0165 3.7980 25.1100 ;
      RECT 3.6640 24.0165 3.6900 25.1100 ;
      RECT 3.5560 24.0165 3.5820 25.1100 ;
      RECT 3.4480 24.0165 3.4740 25.1100 ;
      RECT 3.3400 24.0165 3.3660 25.1100 ;
      RECT 3.2320 24.0165 3.2580 25.1100 ;
      RECT 3.1240 24.0165 3.1500 25.1100 ;
      RECT 3.0160 24.0165 3.0420 25.1100 ;
      RECT 2.9080 24.0165 2.9340 25.1100 ;
      RECT 2.8000 24.0165 2.8260 25.1100 ;
      RECT 2.6920 24.0165 2.7180 25.1100 ;
      RECT 2.5840 24.0165 2.6100 25.1100 ;
      RECT 2.4760 24.0165 2.5020 25.1100 ;
      RECT 2.3680 24.0165 2.3940 25.1100 ;
      RECT 2.2600 24.0165 2.2860 25.1100 ;
      RECT 2.1520 24.0165 2.1780 25.1100 ;
      RECT 2.0440 24.0165 2.0700 25.1100 ;
      RECT 1.9360 24.0165 1.9620 25.1100 ;
      RECT 1.8280 24.0165 1.8540 25.1100 ;
      RECT 1.7200 24.0165 1.7460 25.1100 ;
      RECT 1.6120 24.0165 1.6380 25.1100 ;
      RECT 1.5040 24.0165 1.5300 25.1100 ;
      RECT 1.3960 24.0165 1.4220 25.1100 ;
      RECT 1.2880 24.0165 1.3140 25.1100 ;
      RECT 1.1800 24.0165 1.2060 25.1100 ;
      RECT 1.0720 24.0165 1.0980 25.1100 ;
      RECT 0.9640 24.0165 0.9900 25.1100 ;
      RECT 0.8560 24.0165 0.8820 25.1100 ;
      RECT 0.7480 24.0165 0.7740 25.1100 ;
      RECT 0.6400 24.0165 0.6660 25.1100 ;
      RECT 0.5320 24.0165 0.5580 25.1100 ;
      RECT 0.4240 24.0165 0.4500 25.1100 ;
      RECT 0.3160 24.0165 0.3420 25.1100 ;
      RECT 0.2080 24.0165 0.2340 25.1100 ;
      RECT 0.0050 24.0165 0.0900 25.1100 ;
      RECT 15.5530 25.0965 15.6810 26.1900 ;
      RECT 15.5390 25.7620 15.6810 26.0845 ;
      RECT 15.3190 25.4890 15.4530 26.1900 ;
      RECT 15.2960 25.8240 15.4530 26.0820 ;
      RECT 15.3190 25.0965 15.4170 26.1900 ;
      RECT 15.3190 25.2175 15.4310 25.4570 ;
      RECT 15.3190 25.0965 15.4530 25.1855 ;
      RECT 15.0940 25.5470 15.2280 26.1900 ;
      RECT 15.0940 25.0965 15.1920 26.1900 ;
      RECT 14.6770 25.0965 14.7600 26.1900 ;
      RECT 14.6770 25.1850 14.7740 26.1205 ;
      RECT 30.2680 25.0965 30.3530 26.1900 ;
      RECT 30.1240 25.0965 30.1500 26.1900 ;
      RECT 30.0160 25.0965 30.0420 26.1900 ;
      RECT 29.9080 25.0965 29.9340 26.1900 ;
      RECT 29.8000 25.0965 29.8260 26.1900 ;
      RECT 29.6920 25.0965 29.7180 26.1900 ;
      RECT 29.5840 25.0965 29.6100 26.1900 ;
      RECT 29.4760 25.0965 29.5020 26.1900 ;
      RECT 29.3680 25.0965 29.3940 26.1900 ;
      RECT 29.2600 25.0965 29.2860 26.1900 ;
      RECT 29.1520 25.0965 29.1780 26.1900 ;
      RECT 29.0440 25.0965 29.0700 26.1900 ;
      RECT 28.9360 25.0965 28.9620 26.1900 ;
      RECT 28.8280 25.0965 28.8540 26.1900 ;
      RECT 28.7200 25.0965 28.7460 26.1900 ;
      RECT 28.6120 25.0965 28.6380 26.1900 ;
      RECT 28.5040 25.0965 28.5300 26.1900 ;
      RECT 28.3960 25.0965 28.4220 26.1900 ;
      RECT 28.2880 25.0965 28.3140 26.1900 ;
      RECT 28.1800 25.0965 28.2060 26.1900 ;
      RECT 28.0720 25.0965 28.0980 26.1900 ;
      RECT 27.9640 25.0965 27.9900 26.1900 ;
      RECT 27.8560 25.0965 27.8820 26.1900 ;
      RECT 27.7480 25.0965 27.7740 26.1900 ;
      RECT 27.6400 25.0965 27.6660 26.1900 ;
      RECT 27.5320 25.0965 27.5580 26.1900 ;
      RECT 27.4240 25.0965 27.4500 26.1900 ;
      RECT 27.3160 25.0965 27.3420 26.1900 ;
      RECT 27.2080 25.0965 27.2340 26.1900 ;
      RECT 27.1000 25.0965 27.1260 26.1900 ;
      RECT 26.9920 25.0965 27.0180 26.1900 ;
      RECT 26.8840 25.0965 26.9100 26.1900 ;
      RECT 26.7760 25.0965 26.8020 26.1900 ;
      RECT 26.6680 25.0965 26.6940 26.1900 ;
      RECT 26.5600 25.0965 26.5860 26.1900 ;
      RECT 26.4520 25.0965 26.4780 26.1900 ;
      RECT 26.3440 25.0965 26.3700 26.1900 ;
      RECT 26.2360 25.0965 26.2620 26.1900 ;
      RECT 26.1280 25.0965 26.1540 26.1900 ;
      RECT 26.0200 25.0965 26.0460 26.1900 ;
      RECT 25.9120 25.0965 25.9380 26.1900 ;
      RECT 25.8040 25.0965 25.8300 26.1900 ;
      RECT 25.6960 25.0965 25.7220 26.1900 ;
      RECT 25.5880 25.0965 25.6140 26.1900 ;
      RECT 25.4800 25.0965 25.5060 26.1900 ;
      RECT 25.3720 25.0965 25.3980 26.1900 ;
      RECT 25.2640 25.0965 25.2900 26.1900 ;
      RECT 25.1560 25.0965 25.1820 26.1900 ;
      RECT 25.0480 25.0965 25.0740 26.1900 ;
      RECT 24.9400 25.0965 24.9660 26.1900 ;
      RECT 24.8320 25.0965 24.8580 26.1900 ;
      RECT 24.7240 25.0965 24.7500 26.1900 ;
      RECT 24.6160 25.0965 24.6420 26.1900 ;
      RECT 24.5080 25.0965 24.5340 26.1900 ;
      RECT 24.4000 25.0965 24.4260 26.1900 ;
      RECT 24.2920 25.0965 24.3180 26.1900 ;
      RECT 24.1840 25.0965 24.2100 26.1900 ;
      RECT 24.0760 25.0965 24.1020 26.1900 ;
      RECT 23.9680 25.0965 23.9940 26.1900 ;
      RECT 23.8600 25.0965 23.8860 26.1900 ;
      RECT 23.7520 25.0965 23.7780 26.1900 ;
      RECT 23.6440 25.0965 23.6700 26.1900 ;
      RECT 23.5360 25.0965 23.5620 26.1900 ;
      RECT 23.4280 25.0965 23.4540 26.1900 ;
      RECT 23.3200 25.0965 23.3460 26.1900 ;
      RECT 23.2120 25.0965 23.2380 26.1900 ;
      RECT 23.1040 25.0965 23.1300 26.1900 ;
      RECT 22.9960 25.0965 23.0220 26.1900 ;
      RECT 22.8880 25.0965 22.9140 26.1900 ;
      RECT 22.7800 25.0965 22.8060 26.1900 ;
      RECT 22.6720 25.0965 22.6980 26.1900 ;
      RECT 22.5640 25.0965 22.5900 26.1900 ;
      RECT 22.4560 25.0965 22.4820 26.1900 ;
      RECT 22.3480 25.0965 22.3740 26.1900 ;
      RECT 22.2400 25.0965 22.2660 26.1900 ;
      RECT 22.1320 25.0965 22.1580 26.1900 ;
      RECT 22.0240 25.0965 22.0500 26.1900 ;
      RECT 21.9160 25.0965 21.9420 26.1900 ;
      RECT 21.8080 25.0965 21.8340 26.1900 ;
      RECT 21.7000 25.0965 21.7260 26.1900 ;
      RECT 21.5920 25.0965 21.6180 26.1900 ;
      RECT 21.4840 25.0965 21.5100 26.1900 ;
      RECT 21.3760 25.0965 21.4020 26.1900 ;
      RECT 21.2680 25.0965 21.2940 26.1900 ;
      RECT 21.1600 25.0965 21.1860 26.1900 ;
      RECT 21.0520 25.0965 21.0780 26.1900 ;
      RECT 20.9440 25.0965 20.9700 26.1900 ;
      RECT 20.8360 25.0965 20.8620 26.1900 ;
      RECT 20.7280 25.0965 20.7540 26.1900 ;
      RECT 20.6200 25.0965 20.6460 26.1900 ;
      RECT 20.5120 25.0965 20.5380 26.1900 ;
      RECT 20.4040 25.0965 20.4300 26.1900 ;
      RECT 20.2960 25.0965 20.3220 26.1900 ;
      RECT 20.1880 25.0965 20.2140 26.1900 ;
      RECT 20.0800 25.0965 20.1060 26.1900 ;
      RECT 19.9720 25.0965 19.9980 26.1900 ;
      RECT 19.8640 25.0965 19.8900 26.1900 ;
      RECT 19.7560 25.0965 19.7820 26.1900 ;
      RECT 19.6480 25.0965 19.6740 26.1900 ;
      RECT 19.5400 25.0965 19.5660 26.1900 ;
      RECT 19.4320 25.0965 19.4580 26.1900 ;
      RECT 19.3240 25.0965 19.3500 26.1900 ;
      RECT 19.2160 25.0965 19.2420 26.1900 ;
      RECT 19.1080 25.0965 19.1340 26.1900 ;
      RECT 19.0000 25.0965 19.0260 26.1900 ;
      RECT 18.8920 25.0965 18.9180 26.1900 ;
      RECT 18.7840 25.0965 18.8100 26.1900 ;
      RECT 18.6760 25.0965 18.7020 26.1900 ;
      RECT 18.5680 25.0965 18.5940 26.1900 ;
      RECT 18.4600 25.0965 18.4860 26.1900 ;
      RECT 18.3520 25.0965 18.3780 26.1900 ;
      RECT 18.2440 25.0965 18.2700 26.1900 ;
      RECT 18.1360 25.0965 18.1620 26.1900 ;
      RECT 18.0280 25.0965 18.0540 26.1900 ;
      RECT 17.9200 25.0965 17.9460 26.1900 ;
      RECT 17.8120 25.0965 17.8380 26.1900 ;
      RECT 17.7040 25.0965 17.7300 26.1900 ;
      RECT 17.5960 25.0965 17.6220 26.1900 ;
      RECT 17.4880 25.0965 17.5140 26.1900 ;
      RECT 17.3800 25.0965 17.4060 26.1900 ;
      RECT 17.2720 25.0965 17.2980 26.1900 ;
      RECT 17.1640 25.0965 17.1900 26.1900 ;
      RECT 17.0560 25.0965 17.0820 26.1900 ;
      RECT 16.9480 25.0965 16.9740 26.1900 ;
      RECT 16.8400 25.0965 16.8660 26.1900 ;
      RECT 16.7320 25.0965 16.7580 26.1900 ;
      RECT 16.6240 25.0965 16.6500 26.1900 ;
      RECT 16.5160 25.0965 16.5420 26.1900 ;
      RECT 16.4080 25.0965 16.4340 26.1900 ;
      RECT 16.3000 25.0965 16.3260 26.1900 ;
      RECT 16.0870 25.0965 16.1640 26.1900 ;
      RECT 14.1940 25.0965 14.2710 26.1900 ;
      RECT 14.0320 25.0965 14.0580 26.1900 ;
      RECT 13.9240 25.0965 13.9500 26.1900 ;
      RECT 13.8160 25.0965 13.8420 26.1900 ;
      RECT 13.7080 25.0965 13.7340 26.1900 ;
      RECT 13.6000 25.0965 13.6260 26.1900 ;
      RECT 13.4920 25.0965 13.5180 26.1900 ;
      RECT 13.3840 25.0965 13.4100 26.1900 ;
      RECT 13.2760 25.0965 13.3020 26.1900 ;
      RECT 13.1680 25.0965 13.1940 26.1900 ;
      RECT 13.0600 25.0965 13.0860 26.1900 ;
      RECT 12.9520 25.0965 12.9780 26.1900 ;
      RECT 12.8440 25.0965 12.8700 26.1900 ;
      RECT 12.7360 25.0965 12.7620 26.1900 ;
      RECT 12.6280 25.0965 12.6540 26.1900 ;
      RECT 12.5200 25.0965 12.5460 26.1900 ;
      RECT 12.4120 25.0965 12.4380 26.1900 ;
      RECT 12.3040 25.0965 12.3300 26.1900 ;
      RECT 12.1960 25.0965 12.2220 26.1900 ;
      RECT 12.0880 25.0965 12.1140 26.1900 ;
      RECT 11.9800 25.0965 12.0060 26.1900 ;
      RECT 11.8720 25.0965 11.8980 26.1900 ;
      RECT 11.7640 25.0965 11.7900 26.1900 ;
      RECT 11.6560 25.0965 11.6820 26.1900 ;
      RECT 11.5480 25.0965 11.5740 26.1900 ;
      RECT 11.4400 25.0965 11.4660 26.1900 ;
      RECT 11.3320 25.0965 11.3580 26.1900 ;
      RECT 11.2240 25.0965 11.2500 26.1900 ;
      RECT 11.1160 25.0965 11.1420 26.1900 ;
      RECT 11.0080 25.0965 11.0340 26.1900 ;
      RECT 10.9000 25.0965 10.9260 26.1900 ;
      RECT 10.7920 25.0965 10.8180 26.1900 ;
      RECT 10.6840 25.0965 10.7100 26.1900 ;
      RECT 10.5760 25.0965 10.6020 26.1900 ;
      RECT 10.4680 25.0965 10.4940 26.1900 ;
      RECT 10.3600 25.0965 10.3860 26.1900 ;
      RECT 10.2520 25.0965 10.2780 26.1900 ;
      RECT 10.1440 25.0965 10.1700 26.1900 ;
      RECT 10.0360 25.0965 10.0620 26.1900 ;
      RECT 9.9280 25.0965 9.9540 26.1900 ;
      RECT 9.8200 25.0965 9.8460 26.1900 ;
      RECT 9.7120 25.0965 9.7380 26.1900 ;
      RECT 9.6040 25.0965 9.6300 26.1900 ;
      RECT 9.4960 25.0965 9.5220 26.1900 ;
      RECT 9.3880 25.0965 9.4140 26.1900 ;
      RECT 9.2800 25.0965 9.3060 26.1900 ;
      RECT 9.1720 25.0965 9.1980 26.1900 ;
      RECT 9.0640 25.0965 9.0900 26.1900 ;
      RECT 8.9560 25.0965 8.9820 26.1900 ;
      RECT 8.8480 25.0965 8.8740 26.1900 ;
      RECT 8.7400 25.0965 8.7660 26.1900 ;
      RECT 8.6320 25.0965 8.6580 26.1900 ;
      RECT 8.5240 25.0965 8.5500 26.1900 ;
      RECT 8.4160 25.0965 8.4420 26.1900 ;
      RECT 8.3080 25.0965 8.3340 26.1900 ;
      RECT 8.2000 25.0965 8.2260 26.1900 ;
      RECT 8.0920 25.0965 8.1180 26.1900 ;
      RECT 7.9840 25.0965 8.0100 26.1900 ;
      RECT 7.8760 25.0965 7.9020 26.1900 ;
      RECT 7.7680 25.0965 7.7940 26.1900 ;
      RECT 7.6600 25.0965 7.6860 26.1900 ;
      RECT 7.5520 25.0965 7.5780 26.1900 ;
      RECT 7.4440 25.0965 7.4700 26.1900 ;
      RECT 7.3360 25.0965 7.3620 26.1900 ;
      RECT 7.2280 25.0965 7.2540 26.1900 ;
      RECT 7.1200 25.0965 7.1460 26.1900 ;
      RECT 7.0120 25.0965 7.0380 26.1900 ;
      RECT 6.9040 25.0965 6.9300 26.1900 ;
      RECT 6.7960 25.0965 6.8220 26.1900 ;
      RECT 6.6880 25.0965 6.7140 26.1900 ;
      RECT 6.5800 25.0965 6.6060 26.1900 ;
      RECT 6.4720 25.0965 6.4980 26.1900 ;
      RECT 6.3640 25.0965 6.3900 26.1900 ;
      RECT 6.2560 25.0965 6.2820 26.1900 ;
      RECT 6.1480 25.0965 6.1740 26.1900 ;
      RECT 6.0400 25.0965 6.0660 26.1900 ;
      RECT 5.9320 25.0965 5.9580 26.1900 ;
      RECT 5.8240 25.0965 5.8500 26.1900 ;
      RECT 5.7160 25.0965 5.7420 26.1900 ;
      RECT 5.6080 25.0965 5.6340 26.1900 ;
      RECT 5.5000 25.0965 5.5260 26.1900 ;
      RECT 5.3920 25.0965 5.4180 26.1900 ;
      RECT 5.2840 25.0965 5.3100 26.1900 ;
      RECT 5.1760 25.0965 5.2020 26.1900 ;
      RECT 5.0680 25.0965 5.0940 26.1900 ;
      RECT 4.9600 25.0965 4.9860 26.1900 ;
      RECT 4.8520 25.0965 4.8780 26.1900 ;
      RECT 4.7440 25.0965 4.7700 26.1900 ;
      RECT 4.6360 25.0965 4.6620 26.1900 ;
      RECT 4.5280 25.0965 4.5540 26.1900 ;
      RECT 4.4200 25.0965 4.4460 26.1900 ;
      RECT 4.3120 25.0965 4.3380 26.1900 ;
      RECT 4.2040 25.0965 4.2300 26.1900 ;
      RECT 4.0960 25.0965 4.1220 26.1900 ;
      RECT 3.9880 25.0965 4.0140 26.1900 ;
      RECT 3.8800 25.0965 3.9060 26.1900 ;
      RECT 3.7720 25.0965 3.7980 26.1900 ;
      RECT 3.6640 25.0965 3.6900 26.1900 ;
      RECT 3.5560 25.0965 3.5820 26.1900 ;
      RECT 3.4480 25.0965 3.4740 26.1900 ;
      RECT 3.3400 25.0965 3.3660 26.1900 ;
      RECT 3.2320 25.0965 3.2580 26.1900 ;
      RECT 3.1240 25.0965 3.1500 26.1900 ;
      RECT 3.0160 25.0965 3.0420 26.1900 ;
      RECT 2.9080 25.0965 2.9340 26.1900 ;
      RECT 2.8000 25.0965 2.8260 26.1900 ;
      RECT 2.6920 25.0965 2.7180 26.1900 ;
      RECT 2.5840 25.0965 2.6100 26.1900 ;
      RECT 2.4760 25.0965 2.5020 26.1900 ;
      RECT 2.3680 25.0965 2.3940 26.1900 ;
      RECT 2.2600 25.0965 2.2860 26.1900 ;
      RECT 2.1520 25.0965 2.1780 26.1900 ;
      RECT 2.0440 25.0965 2.0700 26.1900 ;
      RECT 1.9360 25.0965 1.9620 26.1900 ;
      RECT 1.8280 25.0965 1.8540 26.1900 ;
      RECT 1.7200 25.0965 1.7460 26.1900 ;
      RECT 1.6120 25.0965 1.6380 26.1900 ;
      RECT 1.5040 25.0965 1.5300 26.1900 ;
      RECT 1.3960 25.0965 1.4220 26.1900 ;
      RECT 1.2880 25.0965 1.3140 26.1900 ;
      RECT 1.1800 25.0965 1.2060 26.1900 ;
      RECT 1.0720 25.0965 1.0980 26.1900 ;
      RECT 0.9640 25.0965 0.9900 26.1900 ;
      RECT 0.8560 25.0965 0.8820 26.1900 ;
      RECT 0.7480 25.0965 0.7740 26.1900 ;
      RECT 0.6400 25.0965 0.6660 26.1900 ;
      RECT 0.5320 25.0965 0.5580 26.1900 ;
      RECT 0.4240 25.0965 0.4500 26.1900 ;
      RECT 0.3160 25.0965 0.3420 26.1900 ;
      RECT 0.2080 25.0965 0.2340 26.1900 ;
      RECT 0.0050 25.0965 0.0900 26.1900 ;
      RECT 15.5530 26.1765 15.6810 27.2700 ;
      RECT 15.5390 26.8420 15.6810 27.1645 ;
      RECT 15.3190 26.5690 15.4530 27.2700 ;
      RECT 15.2960 26.9040 15.4530 27.1620 ;
      RECT 15.3190 26.1765 15.4170 27.2700 ;
      RECT 15.3190 26.2975 15.4310 26.5370 ;
      RECT 15.3190 26.1765 15.4530 26.2655 ;
      RECT 15.0940 26.6270 15.2280 27.2700 ;
      RECT 15.0940 26.1765 15.1920 27.2700 ;
      RECT 14.6770 26.1765 14.7600 27.2700 ;
      RECT 14.6770 26.2650 14.7740 27.2005 ;
      RECT 30.2680 26.1765 30.3530 27.2700 ;
      RECT 30.1240 26.1765 30.1500 27.2700 ;
      RECT 30.0160 26.1765 30.0420 27.2700 ;
      RECT 29.9080 26.1765 29.9340 27.2700 ;
      RECT 29.8000 26.1765 29.8260 27.2700 ;
      RECT 29.6920 26.1765 29.7180 27.2700 ;
      RECT 29.5840 26.1765 29.6100 27.2700 ;
      RECT 29.4760 26.1765 29.5020 27.2700 ;
      RECT 29.3680 26.1765 29.3940 27.2700 ;
      RECT 29.2600 26.1765 29.2860 27.2700 ;
      RECT 29.1520 26.1765 29.1780 27.2700 ;
      RECT 29.0440 26.1765 29.0700 27.2700 ;
      RECT 28.9360 26.1765 28.9620 27.2700 ;
      RECT 28.8280 26.1765 28.8540 27.2700 ;
      RECT 28.7200 26.1765 28.7460 27.2700 ;
      RECT 28.6120 26.1765 28.6380 27.2700 ;
      RECT 28.5040 26.1765 28.5300 27.2700 ;
      RECT 28.3960 26.1765 28.4220 27.2700 ;
      RECT 28.2880 26.1765 28.3140 27.2700 ;
      RECT 28.1800 26.1765 28.2060 27.2700 ;
      RECT 28.0720 26.1765 28.0980 27.2700 ;
      RECT 27.9640 26.1765 27.9900 27.2700 ;
      RECT 27.8560 26.1765 27.8820 27.2700 ;
      RECT 27.7480 26.1765 27.7740 27.2700 ;
      RECT 27.6400 26.1765 27.6660 27.2700 ;
      RECT 27.5320 26.1765 27.5580 27.2700 ;
      RECT 27.4240 26.1765 27.4500 27.2700 ;
      RECT 27.3160 26.1765 27.3420 27.2700 ;
      RECT 27.2080 26.1765 27.2340 27.2700 ;
      RECT 27.1000 26.1765 27.1260 27.2700 ;
      RECT 26.9920 26.1765 27.0180 27.2700 ;
      RECT 26.8840 26.1765 26.9100 27.2700 ;
      RECT 26.7760 26.1765 26.8020 27.2700 ;
      RECT 26.6680 26.1765 26.6940 27.2700 ;
      RECT 26.5600 26.1765 26.5860 27.2700 ;
      RECT 26.4520 26.1765 26.4780 27.2700 ;
      RECT 26.3440 26.1765 26.3700 27.2700 ;
      RECT 26.2360 26.1765 26.2620 27.2700 ;
      RECT 26.1280 26.1765 26.1540 27.2700 ;
      RECT 26.0200 26.1765 26.0460 27.2700 ;
      RECT 25.9120 26.1765 25.9380 27.2700 ;
      RECT 25.8040 26.1765 25.8300 27.2700 ;
      RECT 25.6960 26.1765 25.7220 27.2700 ;
      RECT 25.5880 26.1765 25.6140 27.2700 ;
      RECT 25.4800 26.1765 25.5060 27.2700 ;
      RECT 25.3720 26.1765 25.3980 27.2700 ;
      RECT 25.2640 26.1765 25.2900 27.2700 ;
      RECT 25.1560 26.1765 25.1820 27.2700 ;
      RECT 25.0480 26.1765 25.0740 27.2700 ;
      RECT 24.9400 26.1765 24.9660 27.2700 ;
      RECT 24.8320 26.1765 24.8580 27.2700 ;
      RECT 24.7240 26.1765 24.7500 27.2700 ;
      RECT 24.6160 26.1765 24.6420 27.2700 ;
      RECT 24.5080 26.1765 24.5340 27.2700 ;
      RECT 24.4000 26.1765 24.4260 27.2700 ;
      RECT 24.2920 26.1765 24.3180 27.2700 ;
      RECT 24.1840 26.1765 24.2100 27.2700 ;
      RECT 24.0760 26.1765 24.1020 27.2700 ;
      RECT 23.9680 26.1765 23.9940 27.2700 ;
      RECT 23.8600 26.1765 23.8860 27.2700 ;
      RECT 23.7520 26.1765 23.7780 27.2700 ;
      RECT 23.6440 26.1765 23.6700 27.2700 ;
      RECT 23.5360 26.1765 23.5620 27.2700 ;
      RECT 23.4280 26.1765 23.4540 27.2700 ;
      RECT 23.3200 26.1765 23.3460 27.2700 ;
      RECT 23.2120 26.1765 23.2380 27.2700 ;
      RECT 23.1040 26.1765 23.1300 27.2700 ;
      RECT 22.9960 26.1765 23.0220 27.2700 ;
      RECT 22.8880 26.1765 22.9140 27.2700 ;
      RECT 22.7800 26.1765 22.8060 27.2700 ;
      RECT 22.6720 26.1765 22.6980 27.2700 ;
      RECT 22.5640 26.1765 22.5900 27.2700 ;
      RECT 22.4560 26.1765 22.4820 27.2700 ;
      RECT 22.3480 26.1765 22.3740 27.2700 ;
      RECT 22.2400 26.1765 22.2660 27.2700 ;
      RECT 22.1320 26.1765 22.1580 27.2700 ;
      RECT 22.0240 26.1765 22.0500 27.2700 ;
      RECT 21.9160 26.1765 21.9420 27.2700 ;
      RECT 21.8080 26.1765 21.8340 27.2700 ;
      RECT 21.7000 26.1765 21.7260 27.2700 ;
      RECT 21.5920 26.1765 21.6180 27.2700 ;
      RECT 21.4840 26.1765 21.5100 27.2700 ;
      RECT 21.3760 26.1765 21.4020 27.2700 ;
      RECT 21.2680 26.1765 21.2940 27.2700 ;
      RECT 21.1600 26.1765 21.1860 27.2700 ;
      RECT 21.0520 26.1765 21.0780 27.2700 ;
      RECT 20.9440 26.1765 20.9700 27.2700 ;
      RECT 20.8360 26.1765 20.8620 27.2700 ;
      RECT 20.7280 26.1765 20.7540 27.2700 ;
      RECT 20.6200 26.1765 20.6460 27.2700 ;
      RECT 20.5120 26.1765 20.5380 27.2700 ;
      RECT 20.4040 26.1765 20.4300 27.2700 ;
      RECT 20.2960 26.1765 20.3220 27.2700 ;
      RECT 20.1880 26.1765 20.2140 27.2700 ;
      RECT 20.0800 26.1765 20.1060 27.2700 ;
      RECT 19.9720 26.1765 19.9980 27.2700 ;
      RECT 19.8640 26.1765 19.8900 27.2700 ;
      RECT 19.7560 26.1765 19.7820 27.2700 ;
      RECT 19.6480 26.1765 19.6740 27.2700 ;
      RECT 19.5400 26.1765 19.5660 27.2700 ;
      RECT 19.4320 26.1765 19.4580 27.2700 ;
      RECT 19.3240 26.1765 19.3500 27.2700 ;
      RECT 19.2160 26.1765 19.2420 27.2700 ;
      RECT 19.1080 26.1765 19.1340 27.2700 ;
      RECT 19.0000 26.1765 19.0260 27.2700 ;
      RECT 18.8920 26.1765 18.9180 27.2700 ;
      RECT 18.7840 26.1765 18.8100 27.2700 ;
      RECT 18.6760 26.1765 18.7020 27.2700 ;
      RECT 18.5680 26.1765 18.5940 27.2700 ;
      RECT 18.4600 26.1765 18.4860 27.2700 ;
      RECT 18.3520 26.1765 18.3780 27.2700 ;
      RECT 18.2440 26.1765 18.2700 27.2700 ;
      RECT 18.1360 26.1765 18.1620 27.2700 ;
      RECT 18.0280 26.1765 18.0540 27.2700 ;
      RECT 17.9200 26.1765 17.9460 27.2700 ;
      RECT 17.8120 26.1765 17.8380 27.2700 ;
      RECT 17.7040 26.1765 17.7300 27.2700 ;
      RECT 17.5960 26.1765 17.6220 27.2700 ;
      RECT 17.4880 26.1765 17.5140 27.2700 ;
      RECT 17.3800 26.1765 17.4060 27.2700 ;
      RECT 17.2720 26.1765 17.2980 27.2700 ;
      RECT 17.1640 26.1765 17.1900 27.2700 ;
      RECT 17.0560 26.1765 17.0820 27.2700 ;
      RECT 16.9480 26.1765 16.9740 27.2700 ;
      RECT 16.8400 26.1765 16.8660 27.2700 ;
      RECT 16.7320 26.1765 16.7580 27.2700 ;
      RECT 16.6240 26.1765 16.6500 27.2700 ;
      RECT 16.5160 26.1765 16.5420 27.2700 ;
      RECT 16.4080 26.1765 16.4340 27.2700 ;
      RECT 16.3000 26.1765 16.3260 27.2700 ;
      RECT 16.0870 26.1765 16.1640 27.2700 ;
      RECT 14.1940 26.1765 14.2710 27.2700 ;
      RECT 14.0320 26.1765 14.0580 27.2700 ;
      RECT 13.9240 26.1765 13.9500 27.2700 ;
      RECT 13.8160 26.1765 13.8420 27.2700 ;
      RECT 13.7080 26.1765 13.7340 27.2700 ;
      RECT 13.6000 26.1765 13.6260 27.2700 ;
      RECT 13.4920 26.1765 13.5180 27.2700 ;
      RECT 13.3840 26.1765 13.4100 27.2700 ;
      RECT 13.2760 26.1765 13.3020 27.2700 ;
      RECT 13.1680 26.1765 13.1940 27.2700 ;
      RECT 13.0600 26.1765 13.0860 27.2700 ;
      RECT 12.9520 26.1765 12.9780 27.2700 ;
      RECT 12.8440 26.1765 12.8700 27.2700 ;
      RECT 12.7360 26.1765 12.7620 27.2700 ;
      RECT 12.6280 26.1765 12.6540 27.2700 ;
      RECT 12.5200 26.1765 12.5460 27.2700 ;
      RECT 12.4120 26.1765 12.4380 27.2700 ;
      RECT 12.3040 26.1765 12.3300 27.2700 ;
      RECT 12.1960 26.1765 12.2220 27.2700 ;
      RECT 12.0880 26.1765 12.1140 27.2700 ;
      RECT 11.9800 26.1765 12.0060 27.2700 ;
      RECT 11.8720 26.1765 11.8980 27.2700 ;
      RECT 11.7640 26.1765 11.7900 27.2700 ;
      RECT 11.6560 26.1765 11.6820 27.2700 ;
      RECT 11.5480 26.1765 11.5740 27.2700 ;
      RECT 11.4400 26.1765 11.4660 27.2700 ;
      RECT 11.3320 26.1765 11.3580 27.2700 ;
      RECT 11.2240 26.1765 11.2500 27.2700 ;
      RECT 11.1160 26.1765 11.1420 27.2700 ;
      RECT 11.0080 26.1765 11.0340 27.2700 ;
      RECT 10.9000 26.1765 10.9260 27.2700 ;
      RECT 10.7920 26.1765 10.8180 27.2700 ;
      RECT 10.6840 26.1765 10.7100 27.2700 ;
      RECT 10.5760 26.1765 10.6020 27.2700 ;
      RECT 10.4680 26.1765 10.4940 27.2700 ;
      RECT 10.3600 26.1765 10.3860 27.2700 ;
      RECT 10.2520 26.1765 10.2780 27.2700 ;
      RECT 10.1440 26.1765 10.1700 27.2700 ;
      RECT 10.0360 26.1765 10.0620 27.2700 ;
      RECT 9.9280 26.1765 9.9540 27.2700 ;
      RECT 9.8200 26.1765 9.8460 27.2700 ;
      RECT 9.7120 26.1765 9.7380 27.2700 ;
      RECT 9.6040 26.1765 9.6300 27.2700 ;
      RECT 9.4960 26.1765 9.5220 27.2700 ;
      RECT 9.3880 26.1765 9.4140 27.2700 ;
      RECT 9.2800 26.1765 9.3060 27.2700 ;
      RECT 9.1720 26.1765 9.1980 27.2700 ;
      RECT 9.0640 26.1765 9.0900 27.2700 ;
      RECT 8.9560 26.1765 8.9820 27.2700 ;
      RECT 8.8480 26.1765 8.8740 27.2700 ;
      RECT 8.7400 26.1765 8.7660 27.2700 ;
      RECT 8.6320 26.1765 8.6580 27.2700 ;
      RECT 8.5240 26.1765 8.5500 27.2700 ;
      RECT 8.4160 26.1765 8.4420 27.2700 ;
      RECT 8.3080 26.1765 8.3340 27.2700 ;
      RECT 8.2000 26.1765 8.2260 27.2700 ;
      RECT 8.0920 26.1765 8.1180 27.2700 ;
      RECT 7.9840 26.1765 8.0100 27.2700 ;
      RECT 7.8760 26.1765 7.9020 27.2700 ;
      RECT 7.7680 26.1765 7.7940 27.2700 ;
      RECT 7.6600 26.1765 7.6860 27.2700 ;
      RECT 7.5520 26.1765 7.5780 27.2700 ;
      RECT 7.4440 26.1765 7.4700 27.2700 ;
      RECT 7.3360 26.1765 7.3620 27.2700 ;
      RECT 7.2280 26.1765 7.2540 27.2700 ;
      RECT 7.1200 26.1765 7.1460 27.2700 ;
      RECT 7.0120 26.1765 7.0380 27.2700 ;
      RECT 6.9040 26.1765 6.9300 27.2700 ;
      RECT 6.7960 26.1765 6.8220 27.2700 ;
      RECT 6.6880 26.1765 6.7140 27.2700 ;
      RECT 6.5800 26.1765 6.6060 27.2700 ;
      RECT 6.4720 26.1765 6.4980 27.2700 ;
      RECT 6.3640 26.1765 6.3900 27.2700 ;
      RECT 6.2560 26.1765 6.2820 27.2700 ;
      RECT 6.1480 26.1765 6.1740 27.2700 ;
      RECT 6.0400 26.1765 6.0660 27.2700 ;
      RECT 5.9320 26.1765 5.9580 27.2700 ;
      RECT 5.8240 26.1765 5.8500 27.2700 ;
      RECT 5.7160 26.1765 5.7420 27.2700 ;
      RECT 5.6080 26.1765 5.6340 27.2700 ;
      RECT 5.5000 26.1765 5.5260 27.2700 ;
      RECT 5.3920 26.1765 5.4180 27.2700 ;
      RECT 5.2840 26.1765 5.3100 27.2700 ;
      RECT 5.1760 26.1765 5.2020 27.2700 ;
      RECT 5.0680 26.1765 5.0940 27.2700 ;
      RECT 4.9600 26.1765 4.9860 27.2700 ;
      RECT 4.8520 26.1765 4.8780 27.2700 ;
      RECT 4.7440 26.1765 4.7700 27.2700 ;
      RECT 4.6360 26.1765 4.6620 27.2700 ;
      RECT 4.5280 26.1765 4.5540 27.2700 ;
      RECT 4.4200 26.1765 4.4460 27.2700 ;
      RECT 4.3120 26.1765 4.3380 27.2700 ;
      RECT 4.2040 26.1765 4.2300 27.2700 ;
      RECT 4.0960 26.1765 4.1220 27.2700 ;
      RECT 3.9880 26.1765 4.0140 27.2700 ;
      RECT 3.8800 26.1765 3.9060 27.2700 ;
      RECT 3.7720 26.1765 3.7980 27.2700 ;
      RECT 3.6640 26.1765 3.6900 27.2700 ;
      RECT 3.5560 26.1765 3.5820 27.2700 ;
      RECT 3.4480 26.1765 3.4740 27.2700 ;
      RECT 3.3400 26.1765 3.3660 27.2700 ;
      RECT 3.2320 26.1765 3.2580 27.2700 ;
      RECT 3.1240 26.1765 3.1500 27.2700 ;
      RECT 3.0160 26.1765 3.0420 27.2700 ;
      RECT 2.9080 26.1765 2.9340 27.2700 ;
      RECT 2.8000 26.1765 2.8260 27.2700 ;
      RECT 2.6920 26.1765 2.7180 27.2700 ;
      RECT 2.5840 26.1765 2.6100 27.2700 ;
      RECT 2.4760 26.1765 2.5020 27.2700 ;
      RECT 2.3680 26.1765 2.3940 27.2700 ;
      RECT 2.2600 26.1765 2.2860 27.2700 ;
      RECT 2.1520 26.1765 2.1780 27.2700 ;
      RECT 2.0440 26.1765 2.0700 27.2700 ;
      RECT 1.9360 26.1765 1.9620 27.2700 ;
      RECT 1.8280 26.1765 1.8540 27.2700 ;
      RECT 1.7200 26.1765 1.7460 27.2700 ;
      RECT 1.6120 26.1765 1.6380 27.2700 ;
      RECT 1.5040 26.1765 1.5300 27.2700 ;
      RECT 1.3960 26.1765 1.4220 27.2700 ;
      RECT 1.2880 26.1765 1.3140 27.2700 ;
      RECT 1.1800 26.1765 1.2060 27.2700 ;
      RECT 1.0720 26.1765 1.0980 27.2700 ;
      RECT 0.9640 26.1765 0.9900 27.2700 ;
      RECT 0.8560 26.1765 0.8820 27.2700 ;
      RECT 0.7480 26.1765 0.7740 27.2700 ;
      RECT 0.6400 26.1765 0.6660 27.2700 ;
      RECT 0.5320 26.1765 0.5580 27.2700 ;
      RECT 0.4240 26.1765 0.4500 27.2700 ;
      RECT 0.3160 26.1765 0.3420 27.2700 ;
      RECT 0.2080 26.1765 0.2340 27.2700 ;
      RECT 0.0050 26.1765 0.0900 27.2700 ;
      RECT 15.5530 27.2565 15.6810 28.3500 ;
      RECT 15.5390 27.9220 15.6810 28.2445 ;
      RECT 15.3190 27.6490 15.4530 28.3500 ;
      RECT 15.2960 27.9840 15.4530 28.2420 ;
      RECT 15.3190 27.2565 15.4170 28.3500 ;
      RECT 15.3190 27.3775 15.4310 27.6170 ;
      RECT 15.3190 27.2565 15.4530 27.3455 ;
      RECT 15.0940 27.7070 15.2280 28.3500 ;
      RECT 15.0940 27.2565 15.1920 28.3500 ;
      RECT 14.6770 27.2565 14.7600 28.3500 ;
      RECT 14.6770 27.3450 14.7740 28.2805 ;
      RECT 30.2680 27.2565 30.3530 28.3500 ;
      RECT 30.1240 27.2565 30.1500 28.3500 ;
      RECT 30.0160 27.2565 30.0420 28.3500 ;
      RECT 29.9080 27.2565 29.9340 28.3500 ;
      RECT 29.8000 27.2565 29.8260 28.3500 ;
      RECT 29.6920 27.2565 29.7180 28.3500 ;
      RECT 29.5840 27.2565 29.6100 28.3500 ;
      RECT 29.4760 27.2565 29.5020 28.3500 ;
      RECT 29.3680 27.2565 29.3940 28.3500 ;
      RECT 29.2600 27.2565 29.2860 28.3500 ;
      RECT 29.1520 27.2565 29.1780 28.3500 ;
      RECT 29.0440 27.2565 29.0700 28.3500 ;
      RECT 28.9360 27.2565 28.9620 28.3500 ;
      RECT 28.8280 27.2565 28.8540 28.3500 ;
      RECT 28.7200 27.2565 28.7460 28.3500 ;
      RECT 28.6120 27.2565 28.6380 28.3500 ;
      RECT 28.5040 27.2565 28.5300 28.3500 ;
      RECT 28.3960 27.2565 28.4220 28.3500 ;
      RECT 28.2880 27.2565 28.3140 28.3500 ;
      RECT 28.1800 27.2565 28.2060 28.3500 ;
      RECT 28.0720 27.2565 28.0980 28.3500 ;
      RECT 27.9640 27.2565 27.9900 28.3500 ;
      RECT 27.8560 27.2565 27.8820 28.3500 ;
      RECT 27.7480 27.2565 27.7740 28.3500 ;
      RECT 27.6400 27.2565 27.6660 28.3500 ;
      RECT 27.5320 27.2565 27.5580 28.3500 ;
      RECT 27.4240 27.2565 27.4500 28.3500 ;
      RECT 27.3160 27.2565 27.3420 28.3500 ;
      RECT 27.2080 27.2565 27.2340 28.3500 ;
      RECT 27.1000 27.2565 27.1260 28.3500 ;
      RECT 26.9920 27.2565 27.0180 28.3500 ;
      RECT 26.8840 27.2565 26.9100 28.3500 ;
      RECT 26.7760 27.2565 26.8020 28.3500 ;
      RECT 26.6680 27.2565 26.6940 28.3500 ;
      RECT 26.5600 27.2565 26.5860 28.3500 ;
      RECT 26.4520 27.2565 26.4780 28.3500 ;
      RECT 26.3440 27.2565 26.3700 28.3500 ;
      RECT 26.2360 27.2565 26.2620 28.3500 ;
      RECT 26.1280 27.2565 26.1540 28.3500 ;
      RECT 26.0200 27.2565 26.0460 28.3500 ;
      RECT 25.9120 27.2565 25.9380 28.3500 ;
      RECT 25.8040 27.2565 25.8300 28.3500 ;
      RECT 25.6960 27.2565 25.7220 28.3500 ;
      RECT 25.5880 27.2565 25.6140 28.3500 ;
      RECT 25.4800 27.2565 25.5060 28.3500 ;
      RECT 25.3720 27.2565 25.3980 28.3500 ;
      RECT 25.2640 27.2565 25.2900 28.3500 ;
      RECT 25.1560 27.2565 25.1820 28.3500 ;
      RECT 25.0480 27.2565 25.0740 28.3500 ;
      RECT 24.9400 27.2565 24.9660 28.3500 ;
      RECT 24.8320 27.2565 24.8580 28.3500 ;
      RECT 24.7240 27.2565 24.7500 28.3500 ;
      RECT 24.6160 27.2565 24.6420 28.3500 ;
      RECT 24.5080 27.2565 24.5340 28.3500 ;
      RECT 24.4000 27.2565 24.4260 28.3500 ;
      RECT 24.2920 27.2565 24.3180 28.3500 ;
      RECT 24.1840 27.2565 24.2100 28.3500 ;
      RECT 24.0760 27.2565 24.1020 28.3500 ;
      RECT 23.9680 27.2565 23.9940 28.3500 ;
      RECT 23.8600 27.2565 23.8860 28.3500 ;
      RECT 23.7520 27.2565 23.7780 28.3500 ;
      RECT 23.6440 27.2565 23.6700 28.3500 ;
      RECT 23.5360 27.2565 23.5620 28.3500 ;
      RECT 23.4280 27.2565 23.4540 28.3500 ;
      RECT 23.3200 27.2565 23.3460 28.3500 ;
      RECT 23.2120 27.2565 23.2380 28.3500 ;
      RECT 23.1040 27.2565 23.1300 28.3500 ;
      RECT 22.9960 27.2565 23.0220 28.3500 ;
      RECT 22.8880 27.2565 22.9140 28.3500 ;
      RECT 22.7800 27.2565 22.8060 28.3500 ;
      RECT 22.6720 27.2565 22.6980 28.3500 ;
      RECT 22.5640 27.2565 22.5900 28.3500 ;
      RECT 22.4560 27.2565 22.4820 28.3500 ;
      RECT 22.3480 27.2565 22.3740 28.3500 ;
      RECT 22.2400 27.2565 22.2660 28.3500 ;
      RECT 22.1320 27.2565 22.1580 28.3500 ;
      RECT 22.0240 27.2565 22.0500 28.3500 ;
      RECT 21.9160 27.2565 21.9420 28.3500 ;
      RECT 21.8080 27.2565 21.8340 28.3500 ;
      RECT 21.7000 27.2565 21.7260 28.3500 ;
      RECT 21.5920 27.2565 21.6180 28.3500 ;
      RECT 21.4840 27.2565 21.5100 28.3500 ;
      RECT 21.3760 27.2565 21.4020 28.3500 ;
      RECT 21.2680 27.2565 21.2940 28.3500 ;
      RECT 21.1600 27.2565 21.1860 28.3500 ;
      RECT 21.0520 27.2565 21.0780 28.3500 ;
      RECT 20.9440 27.2565 20.9700 28.3500 ;
      RECT 20.8360 27.2565 20.8620 28.3500 ;
      RECT 20.7280 27.2565 20.7540 28.3500 ;
      RECT 20.6200 27.2565 20.6460 28.3500 ;
      RECT 20.5120 27.2565 20.5380 28.3500 ;
      RECT 20.4040 27.2565 20.4300 28.3500 ;
      RECT 20.2960 27.2565 20.3220 28.3500 ;
      RECT 20.1880 27.2565 20.2140 28.3500 ;
      RECT 20.0800 27.2565 20.1060 28.3500 ;
      RECT 19.9720 27.2565 19.9980 28.3500 ;
      RECT 19.8640 27.2565 19.8900 28.3500 ;
      RECT 19.7560 27.2565 19.7820 28.3500 ;
      RECT 19.6480 27.2565 19.6740 28.3500 ;
      RECT 19.5400 27.2565 19.5660 28.3500 ;
      RECT 19.4320 27.2565 19.4580 28.3500 ;
      RECT 19.3240 27.2565 19.3500 28.3500 ;
      RECT 19.2160 27.2565 19.2420 28.3500 ;
      RECT 19.1080 27.2565 19.1340 28.3500 ;
      RECT 19.0000 27.2565 19.0260 28.3500 ;
      RECT 18.8920 27.2565 18.9180 28.3500 ;
      RECT 18.7840 27.2565 18.8100 28.3500 ;
      RECT 18.6760 27.2565 18.7020 28.3500 ;
      RECT 18.5680 27.2565 18.5940 28.3500 ;
      RECT 18.4600 27.2565 18.4860 28.3500 ;
      RECT 18.3520 27.2565 18.3780 28.3500 ;
      RECT 18.2440 27.2565 18.2700 28.3500 ;
      RECT 18.1360 27.2565 18.1620 28.3500 ;
      RECT 18.0280 27.2565 18.0540 28.3500 ;
      RECT 17.9200 27.2565 17.9460 28.3500 ;
      RECT 17.8120 27.2565 17.8380 28.3500 ;
      RECT 17.7040 27.2565 17.7300 28.3500 ;
      RECT 17.5960 27.2565 17.6220 28.3500 ;
      RECT 17.4880 27.2565 17.5140 28.3500 ;
      RECT 17.3800 27.2565 17.4060 28.3500 ;
      RECT 17.2720 27.2565 17.2980 28.3500 ;
      RECT 17.1640 27.2565 17.1900 28.3500 ;
      RECT 17.0560 27.2565 17.0820 28.3500 ;
      RECT 16.9480 27.2565 16.9740 28.3500 ;
      RECT 16.8400 27.2565 16.8660 28.3500 ;
      RECT 16.7320 27.2565 16.7580 28.3500 ;
      RECT 16.6240 27.2565 16.6500 28.3500 ;
      RECT 16.5160 27.2565 16.5420 28.3500 ;
      RECT 16.4080 27.2565 16.4340 28.3500 ;
      RECT 16.3000 27.2565 16.3260 28.3500 ;
      RECT 16.0870 27.2565 16.1640 28.3500 ;
      RECT 14.1940 27.2565 14.2710 28.3500 ;
      RECT 14.0320 27.2565 14.0580 28.3500 ;
      RECT 13.9240 27.2565 13.9500 28.3500 ;
      RECT 13.8160 27.2565 13.8420 28.3500 ;
      RECT 13.7080 27.2565 13.7340 28.3500 ;
      RECT 13.6000 27.2565 13.6260 28.3500 ;
      RECT 13.4920 27.2565 13.5180 28.3500 ;
      RECT 13.3840 27.2565 13.4100 28.3500 ;
      RECT 13.2760 27.2565 13.3020 28.3500 ;
      RECT 13.1680 27.2565 13.1940 28.3500 ;
      RECT 13.0600 27.2565 13.0860 28.3500 ;
      RECT 12.9520 27.2565 12.9780 28.3500 ;
      RECT 12.8440 27.2565 12.8700 28.3500 ;
      RECT 12.7360 27.2565 12.7620 28.3500 ;
      RECT 12.6280 27.2565 12.6540 28.3500 ;
      RECT 12.5200 27.2565 12.5460 28.3500 ;
      RECT 12.4120 27.2565 12.4380 28.3500 ;
      RECT 12.3040 27.2565 12.3300 28.3500 ;
      RECT 12.1960 27.2565 12.2220 28.3500 ;
      RECT 12.0880 27.2565 12.1140 28.3500 ;
      RECT 11.9800 27.2565 12.0060 28.3500 ;
      RECT 11.8720 27.2565 11.8980 28.3500 ;
      RECT 11.7640 27.2565 11.7900 28.3500 ;
      RECT 11.6560 27.2565 11.6820 28.3500 ;
      RECT 11.5480 27.2565 11.5740 28.3500 ;
      RECT 11.4400 27.2565 11.4660 28.3500 ;
      RECT 11.3320 27.2565 11.3580 28.3500 ;
      RECT 11.2240 27.2565 11.2500 28.3500 ;
      RECT 11.1160 27.2565 11.1420 28.3500 ;
      RECT 11.0080 27.2565 11.0340 28.3500 ;
      RECT 10.9000 27.2565 10.9260 28.3500 ;
      RECT 10.7920 27.2565 10.8180 28.3500 ;
      RECT 10.6840 27.2565 10.7100 28.3500 ;
      RECT 10.5760 27.2565 10.6020 28.3500 ;
      RECT 10.4680 27.2565 10.4940 28.3500 ;
      RECT 10.3600 27.2565 10.3860 28.3500 ;
      RECT 10.2520 27.2565 10.2780 28.3500 ;
      RECT 10.1440 27.2565 10.1700 28.3500 ;
      RECT 10.0360 27.2565 10.0620 28.3500 ;
      RECT 9.9280 27.2565 9.9540 28.3500 ;
      RECT 9.8200 27.2565 9.8460 28.3500 ;
      RECT 9.7120 27.2565 9.7380 28.3500 ;
      RECT 9.6040 27.2565 9.6300 28.3500 ;
      RECT 9.4960 27.2565 9.5220 28.3500 ;
      RECT 9.3880 27.2565 9.4140 28.3500 ;
      RECT 9.2800 27.2565 9.3060 28.3500 ;
      RECT 9.1720 27.2565 9.1980 28.3500 ;
      RECT 9.0640 27.2565 9.0900 28.3500 ;
      RECT 8.9560 27.2565 8.9820 28.3500 ;
      RECT 8.8480 27.2565 8.8740 28.3500 ;
      RECT 8.7400 27.2565 8.7660 28.3500 ;
      RECT 8.6320 27.2565 8.6580 28.3500 ;
      RECT 8.5240 27.2565 8.5500 28.3500 ;
      RECT 8.4160 27.2565 8.4420 28.3500 ;
      RECT 8.3080 27.2565 8.3340 28.3500 ;
      RECT 8.2000 27.2565 8.2260 28.3500 ;
      RECT 8.0920 27.2565 8.1180 28.3500 ;
      RECT 7.9840 27.2565 8.0100 28.3500 ;
      RECT 7.8760 27.2565 7.9020 28.3500 ;
      RECT 7.7680 27.2565 7.7940 28.3500 ;
      RECT 7.6600 27.2565 7.6860 28.3500 ;
      RECT 7.5520 27.2565 7.5780 28.3500 ;
      RECT 7.4440 27.2565 7.4700 28.3500 ;
      RECT 7.3360 27.2565 7.3620 28.3500 ;
      RECT 7.2280 27.2565 7.2540 28.3500 ;
      RECT 7.1200 27.2565 7.1460 28.3500 ;
      RECT 7.0120 27.2565 7.0380 28.3500 ;
      RECT 6.9040 27.2565 6.9300 28.3500 ;
      RECT 6.7960 27.2565 6.8220 28.3500 ;
      RECT 6.6880 27.2565 6.7140 28.3500 ;
      RECT 6.5800 27.2565 6.6060 28.3500 ;
      RECT 6.4720 27.2565 6.4980 28.3500 ;
      RECT 6.3640 27.2565 6.3900 28.3500 ;
      RECT 6.2560 27.2565 6.2820 28.3500 ;
      RECT 6.1480 27.2565 6.1740 28.3500 ;
      RECT 6.0400 27.2565 6.0660 28.3500 ;
      RECT 5.9320 27.2565 5.9580 28.3500 ;
      RECT 5.8240 27.2565 5.8500 28.3500 ;
      RECT 5.7160 27.2565 5.7420 28.3500 ;
      RECT 5.6080 27.2565 5.6340 28.3500 ;
      RECT 5.5000 27.2565 5.5260 28.3500 ;
      RECT 5.3920 27.2565 5.4180 28.3500 ;
      RECT 5.2840 27.2565 5.3100 28.3500 ;
      RECT 5.1760 27.2565 5.2020 28.3500 ;
      RECT 5.0680 27.2565 5.0940 28.3500 ;
      RECT 4.9600 27.2565 4.9860 28.3500 ;
      RECT 4.8520 27.2565 4.8780 28.3500 ;
      RECT 4.7440 27.2565 4.7700 28.3500 ;
      RECT 4.6360 27.2565 4.6620 28.3500 ;
      RECT 4.5280 27.2565 4.5540 28.3500 ;
      RECT 4.4200 27.2565 4.4460 28.3500 ;
      RECT 4.3120 27.2565 4.3380 28.3500 ;
      RECT 4.2040 27.2565 4.2300 28.3500 ;
      RECT 4.0960 27.2565 4.1220 28.3500 ;
      RECT 3.9880 27.2565 4.0140 28.3500 ;
      RECT 3.8800 27.2565 3.9060 28.3500 ;
      RECT 3.7720 27.2565 3.7980 28.3500 ;
      RECT 3.6640 27.2565 3.6900 28.3500 ;
      RECT 3.5560 27.2565 3.5820 28.3500 ;
      RECT 3.4480 27.2565 3.4740 28.3500 ;
      RECT 3.3400 27.2565 3.3660 28.3500 ;
      RECT 3.2320 27.2565 3.2580 28.3500 ;
      RECT 3.1240 27.2565 3.1500 28.3500 ;
      RECT 3.0160 27.2565 3.0420 28.3500 ;
      RECT 2.9080 27.2565 2.9340 28.3500 ;
      RECT 2.8000 27.2565 2.8260 28.3500 ;
      RECT 2.6920 27.2565 2.7180 28.3500 ;
      RECT 2.5840 27.2565 2.6100 28.3500 ;
      RECT 2.4760 27.2565 2.5020 28.3500 ;
      RECT 2.3680 27.2565 2.3940 28.3500 ;
      RECT 2.2600 27.2565 2.2860 28.3500 ;
      RECT 2.1520 27.2565 2.1780 28.3500 ;
      RECT 2.0440 27.2565 2.0700 28.3500 ;
      RECT 1.9360 27.2565 1.9620 28.3500 ;
      RECT 1.8280 27.2565 1.8540 28.3500 ;
      RECT 1.7200 27.2565 1.7460 28.3500 ;
      RECT 1.6120 27.2565 1.6380 28.3500 ;
      RECT 1.5040 27.2565 1.5300 28.3500 ;
      RECT 1.3960 27.2565 1.4220 28.3500 ;
      RECT 1.2880 27.2565 1.3140 28.3500 ;
      RECT 1.1800 27.2565 1.2060 28.3500 ;
      RECT 1.0720 27.2565 1.0980 28.3500 ;
      RECT 0.9640 27.2565 0.9900 28.3500 ;
      RECT 0.8560 27.2565 0.8820 28.3500 ;
      RECT 0.7480 27.2565 0.7740 28.3500 ;
      RECT 0.6400 27.2565 0.6660 28.3500 ;
      RECT 0.5320 27.2565 0.5580 28.3500 ;
      RECT 0.4240 27.2565 0.4500 28.3500 ;
      RECT 0.3160 27.2565 0.3420 28.3500 ;
      RECT 0.2080 27.2565 0.2340 28.3500 ;
      RECT 0.0050 27.2565 0.0900 28.3500 ;
      RECT 15.5530 28.3365 15.6810 29.4300 ;
      RECT 15.5390 29.0020 15.6810 29.3245 ;
      RECT 15.3190 28.7290 15.4530 29.4300 ;
      RECT 15.2960 29.0640 15.4530 29.3220 ;
      RECT 15.3190 28.3365 15.4170 29.4300 ;
      RECT 15.3190 28.4575 15.4310 28.6970 ;
      RECT 15.3190 28.3365 15.4530 28.4255 ;
      RECT 15.0940 28.7870 15.2280 29.4300 ;
      RECT 15.0940 28.3365 15.1920 29.4300 ;
      RECT 14.6770 28.3365 14.7600 29.4300 ;
      RECT 14.6770 28.4250 14.7740 29.3605 ;
      RECT 30.2680 28.3365 30.3530 29.4300 ;
      RECT 30.1240 28.3365 30.1500 29.4300 ;
      RECT 30.0160 28.3365 30.0420 29.4300 ;
      RECT 29.9080 28.3365 29.9340 29.4300 ;
      RECT 29.8000 28.3365 29.8260 29.4300 ;
      RECT 29.6920 28.3365 29.7180 29.4300 ;
      RECT 29.5840 28.3365 29.6100 29.4300 ;
      RECT 29.4760 28.3365 29.5020 29.4300 ;
      RECT 29.3680 28.3365 29.3940 29.4300 ;
      RECT 29.2600 28.3365 29.2860 29.4300 ;
      RECT 29.1520 28.3365 29.1780 29.4300 ;
      RECT 29.0440 28.3365 29.0700 29.4300 ;
      RECT 28.9360 28.3365 28.9620 29.4300 ;
      RECT 28.8280 28.3365 28.8540 29.4300 ;
      RECT 28.7200 28.3365 28.7460 29.4300 ;
      RECT 28.6120 28.3365 28.6380 29.4300 ;
      RECT 28.5040 28.3365 28.5300 29.4300 ;
      RECT 28.3960 28.3365 28.4220 29.4300 ;
      RECT 28.2880 28.3365 28.3140 29.4300 ;
      RECT 28.1800 28.3365 28.2060 29.4300 ;
      RECT 28.0720 28.3365 28.0980 29.4300 ;
      RECT 27.9640 28.3365 27.9900 29.4300 ;
      RECT 27.8560 28.3365 27.8820 29.4300 ;
      RECT 27.7480 28.3365 27.7740 29.4300 ;
      RECT 27.6400 28.3365 27.6660 29.4300 ;
      RECT 27.5320 28.3365 27.5580 29.4300 ;
      RECT 27.4240 28.3365 27.4500 29.4300 ;
      RECT 27.3160 28.3365 27.3420 29.4300 ;
      RECT 27.2080 28.3365 27.2340 29.4300 ;
      RECT 27.1000 28.3365 27.1260 29.4300 ;
      RECT 26.9920 28.3365 27.0180 29.4300 ;
      RECT 26.8840 28.3365 26.9100 29.4300 ;
      RECT 26.7760 28.3365 26.8020 29.4300 ;
      RECT 26.6680 28.3365 26.6940 29.4300 ;
      RECT 26.5600 28.3365 26.5860 29.4300 ;
      RECT 26.4520 28.3365 26.4780 29.4300 ;
      RECT 26.3440 28.3365 26.3700 29.4300 ;
      RECT 26.2360 28.3365 26.2620 29.4300 ;
      RECT 26.1280 28.3365 26.1540 29.4300 ;
      RECT 26.0200 28.3365 26.0460 29.4300 ;
      RECT 25.9120 28.3365 25.9380 29.4300 ;
      RECT 25.8040 28.3365 25.8300 29.4300 ;
      RECT 25.6960 28.3365 25.7220 29.4300 ;
      RECT 25.5880 28.3365 25.6140 29.4300 ;
      RECT 25.4800 28.3365 25.5060 29.4300 ;
      RECT 25.3720 28.3365 25.3980 29.4300 ;
      RECT 25.2640 28.3365 25.2900 29.4300 ;
      RECT 25.1560 28.3365 25.1820 29.4300 ;
      RECT 25.0480 28.3365 25.0740 29.4300 ;
      RECT 24.9400 28.3365 24.9660 29.4300 ;
      RECT 24.8320 28.3365 24.8580 29.4300 ;
      RECT 24.7240 28.3365 24.7500 29.4300 ;
      RECT 24.6160 28.3365 24.6420 29.4300 ;
      RECT 24.5080 28.3365 24.5340 29.4300 ;
      RECT 24.4000 28.3365 24.4260 29.4300 ;
      RECT 24.2920 28.3365 24.3180 29.4300 ;
      RECT 24.1840 28.3365 24.2100 29.4300 ;
      RECT 24.0760 28.3365 24.1020 29.4300 ;
      RECT 23.9680 28.3365 23.9940 29.4300 ;
      RECT 23.8600 28.3365 23.8860 29.4300 ;
      RECT 23.7520 28.3365 23.7780 29.4300 ;
      RECT 23.6440 28.3365 23.6700 29.4300 ;
      RECT 23.5360 28.3365 23.5620 29.4300 ;
      RECT 23.4280 28.3365 23.4540 29.4300 ;
      RECT 23.3200 28.3365 23.3460 29.4300 ;
      RECT 23.2120 28.3365 23.2380 29.4300 ;
      RECT 23.1040 28.3365 23.1300 29.4300 ;
      RECT 22.9960 28.3365 23.0220 29.4300 ;
      RECT 22.8880 28.3365 22.9140 29.4300 ;
      RECT 22.7800 28.3365 22.8060 29.4300 ;
      RECT 22.6720 28.3365 22.6980 29.4300 ;
      RECT 22.5640 28.3365 22.5900 29.4300 ;
      RECT 22.4560 28.3365 22.4820 29.4300 ;
      RECT 22.3480 28.3365 22.3740 29.4300 ;
      RECT 22.2400 28.3365 22.2660 29.4300 ;
      RECT 22.1320 28.3365 22.1580 29.4300 ;
      RECT 22.0240 28.3365 22.0500 29.4300 ;
      RECT 21.9160 28.3365 21.9420 29.4300 ;
      RECT 21.8080 28.3365 21.8340 29.4300 ;
      RECT 21.7000 28.3365 21.7260 29.4300 ;
      RECT 21.5920 28.3365 21.6180 29.4300 ;
      RECT 21.4840 28.3365 21.5100 29.4300 ;
      RECT 21.3760 28.3365 21.4020 29.4300 ;
      RECT 21.2680 28.3365 21.2940 29.4300 ;
      RECT 21.1600 28.3365 21.1860 29.4300 ;
      RECT 21.0520 28.3365 21.0780 29.4300 ;
      RECT 20.9440 28.3365 20.9700 29.4300 ;
      RECT 20.8360 28.3365 20.8620 29.4300 ;
      RECT 20.7280 28.3365 20.7540 29.4300 ;
      RECT 20.6200 28.3365 20.6460 29.4300 ;
      RECT 20.5120 28.3365 20.5380 29.4300 ;
      RECT 20.4040 28.3365 20.4300 29.4300 ;
      RECT 20.2960 28.3365 20.3220 29.4300 ;
      RECT 20.1880 28.3365 20.2140 29.4300 ;
      RECT 20.0800 28.3365 20.1060 29.4300 ;
      RECT 19.9720 28.3365 19.9980 29.4300 ;
      RECT 19.8640 28.3365 19.8900 29.4300 ;
      RECT 19.7560 28.3365 19.7820 29.4300 ;
      RECT 19.6480 28.3365 19.6740 29.4300 ;
      RECT 19.5400 28.3365 19.5660 29.4300 ;
      RECT 19.4320 28.3365 19.4580 29.4300 ;
      RECT 19.3240 28.3365 19.3500 29.4300 ;
      RECT 19.2160 28.3365 19.2420 29.4300 ;
      RECT 19.1080 28.3365 19.1340 29.4300 ;
      RECT 19.0000 28.3365 19.0260 29.4300 ;
      RECT 18.8920 28.3365 18.9180 29.4300 ;
      RECT 18.7840 28.3365 18.8100 29.4300 ;
      RECT 18.6760 28.3365 18.7020 29.4300 ;
      RECT 18.5680 28.3365 18.5940 29.4300 ;
      RECT 18.4600 28.3365 18.4860 29.4300 ;
      RECT 18.3520 28.3365 18.3780 29.4300 ;
      RECT 18.2440 28.3365 18.2700 29.4300 ;
      RECT 18.1360 28.3365 18.1620 29.4300 ;
      RECT 18.0280 28.3365 18.0540 29.4300 ;
      RECT 17.9200 28.3365 17.9460 29.4300 ;
      RECT 17.8120 28.3365 17.8380 29.4300 ;
      RECT 17.7040 28.3365 17.7300 29.4300 ;
      RECT 17.5960 28.3365 17.6220 29.4300 ;
      RECT 17.4880 28.3365 17.5140 29.4300 ;
      RECT 17.3800 28.3365 17.4060 29.4300 ;
      RECT 17.2720 28.3365 17.2980 29.4300 ;
      RECT 17.1640 28.3365 17.1900 29.4300 ;
      RECT 17.0560 28.3365 17.0820 29.4300 ;
      RECT 16.9480 28.3365 16.9740 29.4300 ;
      RECT 16.8400 28.3365 16.8660 29.4300 ;
      RECT 16.7320 28.3365 16.7580 29.4300 ;
      RECT 16.6240 28.3365 16.6500 29.4300 ;
      RECT 16.5160 28.3365 16.5420 29.4300 ;
      RECT 16.4080 28.3365 16.4340 29.4300 ;
      RECT 16.3000 28.3365 16.3260 29.4300 ;
      RECT 16.0870 28.3365 16.1640 29.4300 ;
      RECT 14.1940 28.3365 14.2710 29.4300 ;
      RECT 14.0320 28.3365 14.0580 29.4300 ;
      RECT 13.9240 28.3365 13.9500 29.4300 ;
      RECT 13.8160 28.3365 13.8420 29.4300 ;
      RECT 13.7080 28.3365 13.7340 29.4300 ;
      RECT 13.6000 28.3365 13.6260 29.4300 ;
      RECT 13.4920 28.3365 13.5180 29.4300 ;
      RECT 13.3840 28.3365 13.4100 29.4300 ;
      RECT 13.2760 28.3365 13.3020 29.4300 ;
      RECT 13.1680 28.3365 13.1940 29.4300 ;
      RECT 13.0600 28.3365 13.0860 29.4300 ;
      RECT 12.9520 28.3365 12.9780 29.4300 ;
      RECT 12.8440 28.3365 12.8700 29.4300 ;
      RECT 12.7360 28.3365 12.7620 29.4300 ;
      RECT 12.6280 28.3365 12.6540 29.4300 ;
      RECT 12.5200 28.3365 12.5460 29.4300 ;
      RECT 12.4120 28.3365 12.4380 29.4300 ;
      RECT 12.3040 28.3365 12.3300 29.4300 ;
      RECT 12.1960 28.3365 12.2220 29.4300 ;
      RECT 12.0880 28.3365 12.1140 29.4300 ;
      RECT 11.9800 28.3365 12.0060 29.4300 ;
      RECT 11.8720 28.3365 11.8980 29.4300 ;
      RECT 11.7640 28.3365 11.7900 29.4300 ;
      RECT 11.6560 28.3365 11.6820 29.4300 ;
      RECT 11.5480 28.3365 11.5740 29.4300 ;
      RECT 11.4400 28.3365 11.4660 29.4300 ;
      RECT 11.3320 28.3365 11.3580 29.4300 ;
      RECT 11.2240 28.3365 11.2500 29.4300 ;
      RECT 11.1160 28.3365 11.1420 29.4300 ;
      RECT 11.0080 28.3365 11.0340 29.4300 ;
      RECT 10.9000 28.3365 10.9260 29.4300 ;
      RECT 10.7920 28.3365 10.8180 29.4300 ;
      RECT 10.6840 28.3365 10.7100 29.4300 ;
      RECT 10.5760 28.3365 10.6020 29.4300 ;
      RECT 10.4680 28.3365 10.4940 29.4300 ;
      RECT 10.3600 28.3365 10.3860 29.4300 ;
      RECT 10.2520 28.3365 10.2780 29.4300 ;
      RECT 10.1440 28.3365 10.1700 29.4300 ;
      RECT 10.0360 28.3365 10.0620 29.4300 ;
      RECT 9.9280 28.3365 9.9540 29.4300 ;
      RECT 9.8200 28.3365 9.8460 29.4300 ;
      RECT 9.7120 28.3365 9.7380 29.4300 ;
      RECT 9.6040 28.3365 9.6300 29.4300 ;
      RECT 9.4960 28.3365 9.5220 29.4300 ;
      RECT 9.3880 28.3365 9.4140 29.4300 ;
      RECT 9.2800 28.3365 9.3060 29.4300 ;
      RECT 9.1720 28.3365 9.1980 29.4300 ;
      RECT 9.0640 28.3365 9.0900 29.4300 ;
      RECT 8.9560 28.3365 8.9820 29.4300 ;
      RECT 8.8480 28.3365 8.8740 29.4300 ;
      RECT 8.7400 28.3365 8.7660 29.4300 ;
      RECT 8.6320 28.3365 8.6580 29.4300 ;
      RECT 8.5240 28.3365 8.5500 29.4300 ;
      RECT 8.4160 28.3365 8.4420 29.4300 ;
      RECT 8.3080 28.3365 8.3340 29.4300 ;
      RECT 8.2000 28.3365 8.2260 29.4300 ;
      RECT 8.0920 28.3365 8.1180 29.4300 ;
      RECT 7.9840 28.3365 8.0100 29.4300 ;
      RECT 7.8760 28.3365 7.9020 29.4300 ;
      RECT 7.7680 28.3365 7.7940 29.4300 ;
      RECT 7.6600 28.3365 7.6860 29.4300 ;
      RECT 7.5520 28.3365 7.5780 29.4300 ;
      RECT 7.4440 28.3365 7.4700 29.4300 ;
      RECT 7.3360 28.3365 7.3620 29.4300 ;
      RECT 7.2280 28.3365 7.2540 29.4300 ;
      RECT 7.1200 28.3365 7.1460 29.4300 ;
      RECT 7.0120 28.3365 7.0380 29.4300 ;
      RECT 6.9040 28.3365 6.9300 29.4300 ;
      RECT 6.7960 28.3365 6.8220 29.4300 ;
      RECT 6.6880 28.3365 6.7140 29.4300 ;
      RECT 6.5800 28.3365 6.6060 29.4300 ;
      RECT 6.4720 28.3365 6.4980 29.4300 ;
      RECT 6.3640 28.3365 6.3900 29.4300 ;
      RECT 6.2560 28.3365 6.2820 29.4300 ;
      RECT 6.1480 28.3365 6.1740 29.4300 ;
      RECT 6.0400 28.3365 6.0660 29.4300 ;
      RECT 5.9320 28.3365 5.9580 29.4300 ;
      RECT 5.8240 28.3365 5.8500 29.4300 ;
      RECT 5.7160 28.3365 5.7420 29.4300 ;
      RECT 5.6080 28.3365 5.6340 29.4300 ;
      RECT 5.5000 28.3365 5.5260 29.4300 ;
      RECT 5.3920 28.3365 5.4180 29.4300 ;
      RECT 5.2840 28.3365 5.3100 29.4300 ;
      RECT 5.1760 28.3365 5.2020 29.4300 ;
      RECT 5.0680 28.3365 5.0940 29.4300 ;
      RECT 4.9600 28.3365 4.9860 29.4300 ;
      RECT 4.8520 28.3365 4.8780 29.4300 ;
      RECT 4.7440 28.3365 4.7700 29.4300 ;
      RECT 4.6360 28.3365 4.6620 29.4300 ;
      RECT 4.5280 28.3365 4.5540 29.4300 ;
      RECT 4.4200 28.3365 4.4460 29.4300 ;
      RECT 4.3120 28.3365 4.3380 29.4300 ;
      RECT 4.2040 28.3365 4.2300 29.4300 ;
      RECT 4.0960 28.3365 4.1220 29.4300 ;
      RECT 3.9880 28.3365 4.0140 29.4300 ;
      RECT 3.8800 28.3365 3.9060 29.4300 ;
      RECT 3.7720 28.3365 3.7980 29.4300 ;
      RECT 3.6640 28.3365 3.6900 29.4300 ;
      RECT 3.5560 28.3365 3.5820 29.4300 ;
      RECT 3.4480 28.3365 3.4740 29.4300 ;
      RECT 3.3400 28.3365 3.3660 29.4300 ;
      RECT 3.2320 28.3365 3.2580 29.4300 ;
      RECT 3.1240 28.3365 3.1500 29.4300 ;
      RECT 3.0160 28.3365 3.0420 29.4300 ;
      RECT 2.9080 28.3365 2.9340 29.4300 ;
      RECT 2.8000 28.3365 2.8260 29.4300 ;
      RECT 2.6920 28.3365 2.7180 29.4300 ;
      RECT 2.5840 28.3365 2.6100 29.4300 ;
      RECT 2.4760 28.3365 2.5020 29.4300 ;
      RECT 2.3680 28.3365 2.3940 29.4300 ;
      RECT 2.2600 28.3365 2.2860 29.4300 ;
      RECT 2.1520 28.3365 2.1780 29.4300 ;
      RECT 2.0440 28.3365 2.0700 29.4300 ;
      RECT 1.9360 28.3365 1.9620 29.4300 ;
      RECT 1.8280 28.3365 1.8540 29.4300 ;
      RECT 1.7200 28.3365 1.7460 29.4300 ;
      RECT 1.6120 28.3365 1.6380 29.4300 ;
      RECT 1.5040 28.3365 1.5300 29.4300 ;
      RECT 1.3960 28.3365 1.4220 29.4300 ;
      RECT 1.2880 28.3365 1.3140 29.4300 ;
      RECT 1.1800 28.3365 1.2060 29.4300 ;
      RECT 1.0720 28.3365 1.0980 29.4300 ;
      RECT 0.9640 28.3365 0.9900 29.4300 ;
      RECT 0.8560 28.3365 0.8820 29.4300 ;
      RECT 0.7480 28.3365 0.7740 29.4300 ;
      RECT 0.6400 28.3365 0.6660 29.4300 ;
      RECT 0.5320 28.3365 0.5580 29.4300 ;
      RECT 0.4240 28.3365 0.4500 29.4300 ;
      RECT 0.3160 28.3365 0.3420 29.4300 ;
      RECT 0.2080 28.3365 0.2340 29.4300 ;
      RECT 0.0050 28.3365 0.0900 29.4300 ;
      RECT 15.5530 29.4165 15.6810 30.5100 ;
      RECT 15.5390 30.0820 15.6810 30.4045 ;
      RECT 15.3190 29.8090 15.4530 30.5100 ;
      RECT 15.2960 30.1440 15.4530 30.4020 ;
      RECT 15.3190 29.4165 15.4170 30.5100 ;
      RECT 15.3190 29.5375 15.4310 29.7770 ;
      RECT 15.3190 29.4165 15.4530 29.5055 ;
      RECT 15.0940 29.8670 15.2280 30.5100 ;
      RECT 15.0940 29.4165 15.1920 30.5100 ;
      RECT 14.6770 29.4165 14.7600 30.5100 ;
      RECT 14.6770 29.5050 14.7740 30.4405 ;
      RECT 30.2680 29.4165 30.3530 30.5100 ;
      RECT 30.1240 29.4165 30.1500 30.5100 ;
      RECT 30.0160 29.4165 30.0420 30.5100 ;
      RECT 29.9080 29.4165 29.9340 30.5100 ;
      RECT 29.8000 29.4165 29.8260 30.5100 ;
      RECT 29.6920 29.4165 29.7180 30.5100 ;
      RECT 29.5840 29.4165 29.6100 30.5100 ;
      RECT 29.4760 29.4165 29.5020 30.5100 ;
      RECT 29.3680 29.4165 29.3940 30.5100 ;
      RECT 29.2600 29.4165 29.2860 30.5100 ;
      RECT 29.1520 29.4165 29.1780 30.5100 ;
      RECT 29.0440 29.4165 29.0700 30.5100 ;
      RECT 28.9360 29.4165 28.9620 30.5100 ;
      RECT 28.8280 29.4165 28.8540 30.5100 ;
      RECT 28.7200 29.4165 28.7460 30.5100 ;
      RECT 28.6120 29.4165 28.6380 30.5100 ;
      RECT 28.5040 29.4165 28.5300 30.5100 ;
      RECT 28.3960 29.4165 28.4220 30.5100 ;
      RECT 28.2880 29.4165 28.3140 30.5100 ;
      RECT 28.1800 29.4165 28.2060 30.5100 ;
      RECT 28.0720 29.4165 28.0980 30.5100 ;
      RECT 27.9640 29.4165 27.9900 30.5100 ;
      RECT 27.8560 29.4165 27.8820 30.5100 ;
      RECT 27.7480 29.4165 27.7740 30.5100 ;
      RECT 27.6400 29.4165 27.6660 30.5100 ;
      RECT 27.5320 29.4165 27.5580 30.5100 ;
      RECT 27.4240 29.4165 27.4500 30.5100 ;
      RECT 27.3160 29.4165 27.3420 30.5100 ;
      RECT 27.2080 29.4165 27.2340 30.5100 ;
      RECT 27.1000 29.4165 27.1260 30.5100 ;
      RECT 26.9920 29.4165 27.0180 30.5100 ;
      RECT 26.8840 29.4165 26.9100 30.5100 ;
      RECT 26.7760 29.4165 26.8020 30.5100 ;
      RECT 26.6680 29.4165 26.6940 30.5100 ;
      RECT 26.5600 29.4165 26.5860 30.5100 ;
      RECT 26.4520 29.4165 26.4780 30.5100 ;
      RECT 26.3440 29.4165 26.3700 30.5100 ;
      RECT 26.2360 29.4165 26.2620 30.5100 ;
      RECT 26.1280 29.4165 26.1540 30.5100 ;
      RECT 26.0200 29.4165 26.0460 30.5100 ;
      RECT 25.9120 29.4165 25.9380 30.5100 ;
      RECT 25.8040 29.4165 25.8300 30.5100 ;
      RECT 25.6960 29.4165 25.7220 30.5100 ;
      RECT 25.5880 29.4165 25.6140 30.5100 ;
      RECT 25.4800 29.4165 25.5060 30.5100 ;
      RECT 25.3720 29.4165 25.3980 30.5100 ;
      RECT 25.2640 29.4165 25.2900 30.5100 ;
      RECT 25.1560 29.4165 25.1820 30.5100 ;
      RECT 25.0480 29.4165 25.0740 30.5100 ;
      RECT 24.9400 29.4165 24.9660 30.5100 ;
      RECT 24.8320 29.4165 24.8580 30.5100 ;
      RECT 24.7240 29.4165 24.7500 30.5100 ;
      RECT 24.6160 29.4165 24.6420 30.5100 ;
      RECT 24.5080 29.4165 24.5340 30.5100 ;
      RECT 24.4000 29.4165 24.4260 30.5100 ;
      RECT 24.2920 29.4165 24.3180 30.5100 ;
      RECT 24.1840 29.4165 24.2100 30.5100 ;
      RECT 24.0760 29.4165 24.1020 30.5100 ;
      RECT 23.9680 29.4165 23.9940 30.5100 ;
      RECT 23.8600 29.4165 23.8860 30.5100 ;
      RECT 23.7520 29.4165 23.7780 30.5100 ;
      RECT 23.6440 29.4165 23.6700 30.5100 ;
      RECT 23.5360 29.4165 23.5620 30.5100 ;
      RECT 23.4280 29.4165 23.4540 30.5100 ;
      RECT 23.3200 29.4165 23.3460 30.5100 ;
      RECT 23.2120 29.4165 23.2380 30.5100 ;
      RECT 23.1040 29.4165 23.1300 30.5100 ;
      RECT 22.9960 29.4165 23.0220 30.5100 ;
      RECT 22.8880 29.4165 22.9140 30.5100 ;
      RECT 22.7800 29.4165 22.8060 30.5100 ;
      RECT 22.6720 29.4165 22.6980 30.5100 ;
      RECT 22.5640 29.4165 22.5900 30.5100 ;
      RECT 22.4560 29.4165 22.4820 30.5100 ;
      RECT 22.3480 29.4165 22.3740 30.5100 ;
      RECT 22.2400 29.4165 22.2660 30.5100 ;
      RECT 22.1320 29.4165 22.1580 30.5100 ;
      RECT 22.0240 29.4165 22.0500 30.5100 ;
      RECT 21.9160 29.4165 21.9420 30.5100 ;
      RECT 21.8080 29.4165 21.8340 30.5100 ;
      RECT 21.7000 29.4165 21.7260 30.5100 ;
      RECT 21.5920 29.4165 21.6180 30.5100 ;
      RECT 21.4840 29.4165 21.5100 30.5100 ;
      RECT 21.3760 29.4165 21.4020 30.5100 ;
      RECT 21.2680 29.4165 21.2940 30.5100 ;
      RECT 21.1600 29.4165 21.1860 30.5100 ;
      RECT 21.0520 29.4165 21.0780 30.5100 ;
      RECT 20.9440 29.4165 20.9700 30.5100 ;
      RECT 20.8360 29.4165 20.8620 30.5100 ;
      RECT 20.7280 29.4165 20.7540 30.5100 ;
      RECT 20.6200 29.4165 20.6460 30.5100 ;
      RECT 20.5120 29.4165 20.5380 30.5100 ;
      RECT 20.4040 29.4165 20.4300 30.5100 ;
      RECT 20.2960 29.4165 20.3220 30.5100 ;
      RECT 20.1880 29.4165 20.2140 30.5100 ;
      RECT 20.0800 29.4165 20.1060 30.5100 ;
      RECT 19.9720 29.4165 19.9980 30.5100 ;
      RECT 19.8640 29.4165 19.8900 30.5100 ;
      RECT 19.7560 29.4165 19.7820 30.5100 ;
      RECT 19.6480 29.4165 19.6740 30.5100 ;
      RECT 19.5400 29.4165 19.5660 30.5100 ;
      RECT 19.4320 29.4165 19.4580 30.5100 ;
      RECT 19.3240 29.4165 19.3500 30.5100 ;
      RECT 19.2160 29.4165 19.2420 30.5100 ;
      RECT 19.1080 29.4165 19.1340 30.5100 ;
      RECT 19.0000 29.4165 19.0260 30.5100 ;
      RECT 18.8920 29.4165 18.9180 30.5100 ;
      RECT 18.7840 29.4165 18.8100 30.5100 ;
      RECT 18.6760 29.4165 18.7020 30.5100 ;
      RECT 18.5680 29.4165 18.5940 30.5100 ;
      RECT 18.4600 29.4165 18.4860 30.5100 ;
      RECT 18.3520 29.4165 18.3780 30.5100 ;
      RECT 18.2440 29.4165 18.2700 30.5100 ;
      RECT 18.1360 29.4165 18.1620 30.5100 ;
      RECT 18.0280 29.4165 18.0540 30.5100 ;
      RECT 17.9200 29.4165 17.9460 30.5100 ;
      RECT 17.8120 29.4165 17.8380 30.5100 ;
      RECT 17.7040 29.4165 17.7300 30.5100 ;
      RECT 17.5960 29.4165 17.6220 30.5100 ;
      RECT 17.4880 29.4165 17.5140 30.5100 ;
      RECT 17.3800 29.4165 17.4060 30.5100 ;
      RECT 17.2720 29.4165 17.2980 30.5100 ;
      RECT 17.1640 29.4165 17.1900 30.5100 ;
      RECT 17.0560 29.4165 17.0820 30.5100 ;
      RECT 16.9480 29.4165 16.9740 30.5100 ;
      RECT 16.8400 29.4165 16.8660 30.5100 ;
      RECT 16.7320 29.4165 16.7580 30.5100 ;
      RECT 16.6240 29.4165 16.6500 30.5100 ;
      RECT 16.5160 29.4165 16.5420 30.5100 ;
      RECT 16.4080 29.4165 16.4340 30.5100 ;
      RECT 16.3000 29.4165 16.3260 30.5100 ;
      RECT 16.0870 29.4165 16.1640 30.5100 ;
      RECT 14.1940 29.4165 14.2710 30.5100 ;
      RECT 14.0320 29.4165 14.0580 30.5100 ;
      RECT 13.9240 29.4165 13.9500 30.5100 ;
      RECT 13.8160 29.4165 13.8420 30.5100 ;
      RECT 13.7080 29.4165 13.7340 30.5100 ;
      RECT 13.6000 29.4165 13.6260 30.5100 ;
      RECT 13.4920 29.4165 13.5180 30.5100 ;
      RECT 13.3840 29.4165 13.4100 30.5100 ;
      RECT 13.2760 29.4165 13.3020 30.5100 ;
      RECT 13.1680 29.4165 13.1940 30.5100 ;
      RECT 13.0600 29.4165 13.0860 30.5100 ;
      RECT 12.9520 29.4165 12.9780 30.5100 ;
      RECT 12.8440 29.4165 12.8700 30.5100 ;
      RECT 12.7360 29.4165 12.7620 30.5100 ;
      RECT 12.6280 29.4165 12.6540 30.5100 ;
      RECT 12.5200 29.4165 12.5460 30.5100 ;
      RECT 12.4120 29.4165 12.4380 30.5100 ;
      RECT 12.3040 29.4165 12.3300 30.5100 ;
      RECT 12.1960 29.4165 12.2220 30.5100 ;
      RECT 12.0880 29.4165 12.1140 30.5100 ;
      RECT 11.9800 29.4165 12.0060 30.5100 ;
      RECT 11.8720 29.4165 11.8980 30.5100 ;
      RECT 11.7640 29.4165 11.7900 30.5100 ;
      RECT 11.6560 29.4165 11.6820 30.5100 ;
      RECT 11.5480 29.4165 11.5740 30.5100 ;
      RECT 11.4400 29.4165 11.4660 30.5100 ;
      RECT 11.3320 29.4165 11.3580 30.5100 ;
      RECT 11.2240 29.4165 11.2500 30.5100 ;
      RECT 11.1160 29.4165 11.1420 30.5100 ;
      RECT 11.0080 29.4165 11.0340 30.5100 ;
      RECT 10.9000 29.4165 10.9260 30.5100 ;
      RECT 10.7920 29.4165 10.8180 30.5100 ;
      RECT 10.6840 29.4165 10.7100 30.5100 ;
      RECT 10.5760 29.4165 10.6020 30.5100 ;
      RECT 10.4680 29.4165 10.4940 30.5100 ;
      RECT 10.3600 29.4165 10.3860 30.5100 ;
      RECT 10.2520 29.4165 10.2780 30.5100 ;
      RECT 10.1440 29.4165 10.1700 30.5100 ;
      RECT 10.0360 29.4165 10.0620 30.5100 ;
      RECT 9.9280 29.4165 9.9540 30.5100 ;
      RECT 9.8200 29.4165 9.8460 30.5100 ;
      RECT 9.7120 29.4165 9.7380 30.5100 ;
      RECT 9.6040 29.4165 9.6300 30.5100 ;
      RECT 9.4960 29.4165 9.5220 30.5100 ;
      RECT 9.3880 29.4165 9.4140 30.5100 ;
      RECT 9.2800 29.4165 9.3060 30.5100 ;
      RECT 9.1720 29.4165 9.1980 30.5100 ;
      RECT 9.0640 29.4165 9.0900 30.5100 ;
      RECT 8.9560 29.4165 8.9820 30.5100 ;
      RECT 8.8480 29.4165 8.8740 30.5100 ;
      RECT 8.7400 29.4165 8.7660 30.5100 ;
      RECT 8.6320 29.4165 8.6580 30.5100 ;
      RECT 8.5240 29.4165 8.5500 30.5100 ;
      RECT 8.4160 29.4165 8.4420 30.5100 ;
      RECT 8.3080 29.4165 8.3340 30.5100 ;
      RECT 8.2000 29.4165 8.2260 30.5100 ;
      RECT 8.0920 29.4165 8.1180 30.5100 ;
      RECT 7.9840 29.4165 8.0100 30.5100 ;
      RECT 7.8760 29.4165 7.9020 30.5100 ;
      RECT 7.7680 29.4165 7.7940 30.5100 ;
      RECT 7.6600 29.4165 7.6860 30.5100 ;
      RECT 7.5520 29.4165 7.5780 30.5100 ;
      RECT 7.4440 29.4165 7.4700 30.5100 ;
      RECT 7.3360 29.4165 7.3620 30.5100 ;
      RECT 7.2280 29.4165 7.2540 30.5100 ;
      RECT 7.1200 29.4165 7.1460 30.5100 ;
      RECT 7.0120 29.4165 7.0380 30.5100 ;
      RECT 6.9040 29.4165 6.9300 30.5100 ;
      RECT 6.7960 29.4165 6.8220 30.5100 ;
      RECT 6.6880 29.4165 6.7140 30.5100 ;
      RECT 6.5800 29.4165 6.6060 30.5100 ;
      RECT 6.4720 29.4165 6.4980 30.5100 ;
      RECT 6.3640 29.4165 6.3900 30.5100 ;
      RECT 6.2560 29.4165 6.2820 30.5100 ;
      RECT 6.1480 29.4165 6.1740 30.5100 ;
      RECT 6.0400 29.4165 6.0660 30.5100 ;
      RECT 5.9320 29.4165 5.9580 30.5100 ;
      RECT 5.8240 29.4165 5.8500 30.5100 ;
      RECT 5.7160 29.4165 5.7420 30.5100 ;
      RECT 5.6080 29.4165 5.6340 30.5100 ;
      RECT 5.5000 29.4165 5.5260 30.5100 ;
      RECT 5.3920 29.4165 5.4180 30.5100 ;
      RECT 5.2840 29.4165 5.3100 30.5100 ;
      RECT 5.1760 29.4165 5.2020 30.5100 ;
      RECT 5.0680 29.4165 5.0940 30.5100 ;
      RECT 4.9600 29.4165 4.9860 30.5100 ;
      RECT 4.8520 29.4165 4.8780 30.5100 ;
      RECT 4.7440 29.4165 4.7700 30.5100 ;
      RECT 4.6360 29.4165 4.6620 30.5100 ;
      RECT 4.5280 29.4165 4.5540 30.5100 ;
      RECT 4.4200 29.4165 4.4460 30.5100 ;
      RECT 4.3120 29.4165 4.3380 30.5100 ;
      RECT 4.2040 29.4165 4.2300 30.5100 ;
      RECT 4.0960 29.4165 4.1220 30.5100 ;
      RECT 3.9880 29.4165 4.0140 30.5100 ;
      RECT 3.8800 29.4165 3.9060 30.5100 ;
      RECT 3.7720 29.4165 3.7980 30.5100 ;
      RECT 3.6640 29.4165 3.6900 30.5100 ;
      RECT 3.5560 29.4165 3.5820 30.5100 ;
      RECT 3.4480 29.4165 3.4740 30.5100 ;
      RECT 3.3400 29.4165 3.3660 30.5100 ;
      RECT 3.2320 29.4165 3.2580 30.5100 ;
      RECT 3.1240 29.4165 3.1500 30.5100 ;
      RECT 3.0160 29.4165 3.0420 30.5100 ;
      RECT 2.9080 29.4165 2.9340 30.5100 ;
      RECT 2.8000 29.4165 2.8260 30.5100 ;
      RECT 2.6920 29.4165 2.7180 30.5100 ;
      RECT 2.5840 29.4165 2.6100 30.5100 ;
      RECT 2.4760 29.4165 2.5020 30.5100 ;
      RECT 2.3680 29.4165 2.3940 30.5100 ;
      RECT 2.2600 29.4165 2.2860 30.5100 ;
      RECT 2.1520 29.4165 2.1780 30.5100 ;
      RECT 2.0440 29.4165 2.0700 30.5100 ;
      RECT 1.9360 29.4165 1.9620 30.5100 ;
      RECT 1.8280 29.4165 1.8540 30.5100 ;
      RECT 1.7200 29.4165 1.7460 30.5100 ;
      RECT 1.6120 29.4165 1.6380 30.5100 ;
      RECT 1.5040 29.4165 1.5300 30.5100 ;
      RECT 1.3960 29.4165 1.4220 30.5100 ;
      RECT 1.2880 29.4165 1.3140 30.5100 ;
      RECT 1.1800 29.4165 1.2060 30.5100 ;
      RECT 1.0720 29.4165 1.0980 30.5100 ;
      RECT 0.9640 29.4165 0.9900 30.5100 ;
      RECT 0.8560 29.4165 0.8820 30.5100 ;
      RECT 0.7480 29.4165 0.7740 30.5100 ;
      RECT 0.6400 29.4165 0.6660 30.5100 ;
      RECT 0.5320 29.4165 0.5580 30.5100 ;
      RECT 0.4240 29.4165 0.4500 30.5100 ;
      RECT 0.3160 29.4165 0.3420 30.5100 ;
      RECT 0.2080 29.4165 0.2340 30.5100 ;
      RECT 0.0050 29.4165 0.0900 30.5100 ;
      RECT 15.5530 30.4965 15.6810 31.5900 ;
      RECT 15.5390 31.1620 15.6810 31.4845 ;
      RECT 15.3190 30.8890 15.4530 31.5900 ;
      RECT 15.2960 31.2240 15.4530 31.4820 ;
      RECT 15.3190 30.4965 15.4170 31.5900 ;
      RECT 15.3190 30.6175 15.4310 30.8570 ;
      RECT 15.3190 30.4965 15.4530 30.5855 ;
      RECT 15.0940 30.9470 15.2280 31.5900 ;
      RECT 15.0940 30.4965 15.1920 31.5900 ;
      RECT 14.6770 30.4965 14.7600 31.5900 ;
      RECT 14.6770 30.5850 14.7740 31.5205 ;
      RECT 30.2680 30.4965 30.3530 31.5900 ;
      RECT 30.1240 30.4965 30.1500 31.5900 ;
      RECT 30.0160 30.4965 30.0420 31.5900 ;
      RECT 29.9080 30.4965 29.9340 31.5900 ;
      RECT 29.8000 30.4965 29.8260 31.5900 ;
      RECT 29.6920 30.4965 29.7180 31.5900 ;
      RECT 29.5840 30.4965 29.6100 31.5900 ;
      RECT 29.4760 30.4965 29.5020 31.5900 ;
      RECT 29.3680 30.4965 29.3940 31.5900 ;
      RECT 29.2600 30.4965 29.2860 31.5900 ;
      RECT 29.1520 30.4965 29.1780 31.5900 ;
      RECT 29.0440 30.4965 29.0700 31.5900 ;
      RECT 28.9360 30.4965 28.9620 31.5900 ;
      RECT 28.8280 30.4965 28.8540 31.5900 ;
      RECT 28.7200 30.4965 28.7460 31.5900 ;
      RECT 28.6120 30.4965 28.6380 31.5900 ;
      RECT 28.5040 30.4965 28.5300 31.5900 ;
      RECT 28.3960 30.4965 28.4220 31.5900 ;
      RECT 28.2880 30.4965 28.3140 31.5900 ;
      RECT 28.1800 30.4965 28.2060 31.5900 ;
      RECT 28.0720 30.4965 28.0980 31.5900 ;
      RECT 27.9640 30.4965 27.9900 31.5900 ;
      RECT 27.8560 30.4965 27.8820 31.5900 ;
      RECT 27.7480 30.4965 27.7740 31.5900 ;
      RECT 27.6400 30.4965 27.6660 31.5900 ;
      RECT 27.5320 30.4965 27.5580 31.5900 ;
      RECT 27.4240 30.4965 27.4500 31.5900 ;
      RECT 27.3160 30.4965 27.3420 31.5900 ;
      RECT 27.2080 30.4965 27.2340 31.5900 ;
      RECT 27.1000 30.4965 27.1260 31.5900 ;
      RECT 26.9920 30.4965 27.0180 31.5900 ;
      RECT 26.8840 30.4965 26.9100 31.5900 ;
      RECT 26.7760 30.4965 26.8020 31.5900 ;
      RECT 26.6680 30.4965 26.6940 31.5900 ;
      RECT 26.5600 30.4965 26.5860 31.5900 ;
      RECT 26.4520 30.4965 26.4780 31.5900 ;
      RECT 26.3440 30.4965 26.3700 31.5900 ;
      RECT 26.2360 30.4965 26.2620 31.5900 ;
      RECT 26.1280 30.4965 26.1540 31.5900 ;
      RECT 26.0200 30.4965 26.0460 31.5900 ;
      RECT 25.9120 30.4965 25.9380 31.5900 ;
      RECT 25.8040 30.4965 25.8300 31.5900 ;
      RECT 25.6960 30.4965 25.7220 31.5900 ;
      RECT 25.5880 30.4965 25.6140 31.5900 ;
      RECT 25.4800 30.4965 25.5060 31.5900 ;
      RECT 25.3720 30.4965 25.3980 31.5900 ;
      RECT 25.2640 30.4965 25.2900 31.5900 ;
      RECT 25.1560 30.4965 25.1820 31.5900 ;
      RECT 25.0480 30.4965 25.0740 31.5900 ;
      RECT 24.9400 30.4965 24.9660 31.5900 ;
      RECT 24.8320 30.4965 24.8580 31.5900 ;
      RECT 24.7240 30.4965 24.7500 31.5900 ;
      RECT 24.6160 30.4965 24.6420 31.5900 ;
      RECT 24.5080 30.4965 24.5340 31.5900 ;
      RECT 24.4000 30.4965 24.4260 31.5900 ;
      RECT 24.2920 30.4965 24.3180 31.5900 ;
      RECT 24.1840 30.4965 24.2100 31.5900 ;
      RECT 24.0760 30.4965 24.1020 31.5900 ;
      RECT 23.9680 30.4965 23.9940 31.5900 ;
      RECT 23.8600 30.4965 23.8860 31.5900 ;
      RECT 23.7520 30.4965 23.7780 31.5900 ;
      RECT 23.6440 30.4965 23.6700 31.5900 ;
      RECT 23.5360 30.4965 23.5620 31.5900 ;
      RECT 23.4280 30.4965 23.4540 31.5900 ;
      RECT 23.3200 30.4965 23.3460 31.5900 ;
      RECT 23.2120 30.4965 23.2380 31.5900 ;
      RECT 23.1040 30.4965 23.1300 31.5900 ;
      RECT 22.9960 30.4965 23.0220 31.5900 ;
      RECT 22.8880 30.4965 22.9140 31.5900 ;
      RECT 22.7800 30.4965 22.8060 31.5900 ;
      RECT 22.6720 30.4965 22.6980 31.5900 ;
      RECT 22.5640 30.4965 22.5900 31.5900 ;
      RECT 22.4560 30.4965 22.4820 31.5900 ;
      RECT 22.3480 30.4965 22.3740 31.5900 ;
      RECT 22.2400 30.4965 22.2660 31.5900 ;
      RECT 22.1320 30.4965 22.1580 31.5900 ;
      RECT 22.0240 30.4965 22.0500 31.5900 ;
      RECT 21.9160 30.4965 21.9420 31.5900 ;
      RECT 21.8080 30.4965 21.8340 31.5900 ;
      RECT 21.7000 30.4965 21.7260 31.5900 ;
      RECT 21.5920 30.4965 21.6180 31.5900 ;
      RECT 21.4840 30.4965 21.5100 31.5900 ;
      RECT 21.3760 30.4965 21.4020 31.5900 ;
      RECT 21.2680 30.4965 21.2940 31.5900 ;
      RECT 21.1600 30.4965 21.1860 31.5900 ;
      RECT 21.0520 30.4965 21.0780 31.5900 ;
      RECT 20.9440 30.4965 20.9700 31.5900 ;
      RECT 20.8360 30.4965 20.8620 31.5900 ;
      RECT 20.7280 30.4965 20.7540 31.5900 ;
      RECT 20.6200 30.4965 20.6460 31.5900 ;
      RECT 20.5120 30.4965 20.5380 31.5900 ;
      RECT 20.4040 30.4965 20.4300 31.5900 ;
      RECT 20.2960 30.4965 20.3220 31.5900 ;
      RECT 20.1880 30.4965 20.2140 31.5900 ;
      RECT 20.0800 30.4965 20.1060 31.5900 ;
      RECT 19.9720 30.4965 19.9980 31.5900 ;
      RECT 19.8640 30.4965 19.8900 31.5900 ;
      RECT 19.7560 30.4965 19.7820 31.5900 ;
      RECT 19.6480 30.4965 19.6740 31.5900 ;
      RECT 19.5400 30.4965 19.5660 31.5900 ;
      RECT 19.4320 30.4965 19.4580 31.5900 ;
      RECT 19.3240 30.4965 19.3500 31.5900 ;
      RECT 19.2160 30.4965 19.2420 31.5900 ;
      RECT 19.1080 30.4965 19.1340 31.5900 ;
      RECT 19.0000 30.4965 19.0260 31.5900 ;
      RECT 18.8920 30.4965 18.9180 31.5900 ;
      RECT 18.7840 30.4965 18.8100 31.5900 ;
      RECT 18.6760 30.4965 18.7020 31.5900 ;
      RECT 18.5680 30.4965 18.5940 31.5900 ;
      RECT 18.4600 30.4965 18.4860 31.5900 ;
      RECT 18.3520 30.4965 18.3780 31.5900 ;
      RECT 18.2440 30.4965 18.2700 31.5900 ;
      RECT 18.1360 30.4965 18.1620 31.5900 ;
      RECT 18.0280 30.4965 18.0540 31.5900 ;
      RECT 17.9200 30.4965 17.9460 31.5900 ;
      RECT 17.8120 30.4965 17.8380 31.5900 ;
      RECT 17.7040 30.4965 17.7300 31.5900 ;
      RECT 17.5960 30.4965 17.6220 31.5900 ;
      RECT 17.4880 30.4965 17.5140 31.5900 ;
      RECT 17.3800 30.4965 17.4060 31.5900 ;
      RECT 17.2720 30.4965 17.2980 31.5900 ;
      RECT 17.1640 30.4965 17.1900 31.5900 ;
      RECT 17.0560 30.4965 17.0820 31.5900 ;
      RECT 16.9480 30.4965 16.9740 31.5900 ;
      RECT 16.8400 30.4965 16.8660 31.5900 ;
      RECT 16.7320 30.4965 16.7580 31.5900 ;
      RECT 16.6240 30.4965 16.6500 31.5900 ;
      RECT 16.5160 30.4965 16.5420 31.5900 ;
      RECT 16.4080 30.4965 16.4340 31.5900 ;
      RECT 16.3000 30.4965 16.3260 31.5900 ;
      RECT 16.0870 30.4965 16.1640 31.5900 ;
      RECT 14.1940 30.4965 14.2710 31.5900 ;
      RECT 14.0320 30.4965 14.0580 31.5900 ;
      RECT 13.9240 30.4965 13.9500 31.5900 ;
      RECT 13.8160 30.4965 13.8420 31.5900 ;
      RECT 13.7080 30.4965 13.7340 31.5900 ;
      RECT 13.6000 30.4965 13.6260 31.5900 ;
      RECT 13.4920 30.4965 13.5180 31.5900 ;
      RECT 13.3840 30.4965 13.4100 31.5900 ;
      RECT 13.2760 30.4965 13.3020 31.5900 ;
      RECT 13.1680 30.4965 13.1940 31.5900 ;
      RECT 13.0600 30.4965 13.0860 31.5900 ;
      RECT 12.9520 30.4965 12.9780 31.5900 ;
      RECT 12.8440 30.4965 12.8700 31.5900 ;
      RECT 12.7360 30.4965 12.7620 31.5900 ;
      RECT 12.6280 30.4965 12.6540 31.5900 ;
      RECT 12.5200 30.4965 12.5460 31.5900 ;
      RECT 12.4120 30.4965 12.4380 31.5900 ;
      RECT 12.3040 30.4965 12.3300 31.5900 ;
      RECT 12.1960 30.4965 12.2220 31.5900 ;
      RECT 12.0880 30.4965 12.1140 31.5900 ;
      RECT 11.9800 30.4965 12.0060 31.5900 ;
      RECT 11.8720 30.4965 11.8980 31.5900 ;
      RECT 11.7640 30.4965 11.7900 31.5900 ;
      RECT 11.6560 30.4965 11.6820 31.5900 ;
      RECT 11.5480 30.4965 11.5740 31.5900 ;
      RECT 11.4400 30.4965 11.4660 31.5900 ;
      RECT 11.3320 30.4965 11.3580 31.5900 ;
      RECT 11.2240 30.4965 11.2500 31.5900 ;
      RECT 11.1160 30.4965 11.1420 31.5900 ;
      RECT 11.0080 30.4965 11.0340 31.5900 ;
      RECT 10.9000 30.4965 10.9260 31.5900 ;
      RECT 10.7920 30.4965 10.8180 31.5900 ;
      RECT 10.6840 30.4965 10.7100 31.5900 ;
      RECT 10.5760 30.4965 10.6020 31.5900 ;
      RECT 10.4680 30.4965 10.4940 31.5900 ;
      RECT 10.3600 30.4965 10.3860 31.5900 ;
      RECT 10.2520 30.4965 10.2780 31.5900 ;
      RECT 10.1440 30.4965 10.1700 31.5900 ;
      RECT 10.0360 30.4965 10.0620 31.5900 ;
      RECT 9.9280 30.4965 9.9540 31.5900 ;
      RECT 9.8200 30.4965 9.8460 31.5900 ;
      RECT 9.7120 30.4965 9.7380 31.5900 ;
      RECT 9.6040 30.4965 9.6300 31.5900 ;
      RECT 9.4960 30.4965 9.5220 31.5900 ;
      RECT 9.3880 30.4965 9.4140 31.5900 ;
      RECT 9.2800 30.4965 9.3060 31.5900 ;
      RECT 9.1720 30.4965 9.1980 31.5900 ;
      RECT 9.0640 30.4965 9.0900 31.5900 ;
      RECT 8.9560 30.4965 8.9820 31.5900 ;
      RECT 8.8480 30.4965 8.8740 31.5900 ;
      RECT 8.7400 30.4965 8.7660 31.5900 ;
      RECT 8.6320 30.4965 8.6580 31.5900 ;
      RECT 8.5240 30.4965 8.5500 31.5900 ;
      RECT 8.4160 30.4965 8.4420 31.5900 ;
      RECT 8.3080 30.4965 8.3340 31.5900 ;
      RECT 8.2000 30.4965 8.2260 31.5900 ;
      RECT 8.0920 30.4965 8.1180 31.5900 ;
      RECT 7.9840 30.4965 8.0100 31.5900 ;
      RECT 7.8760 30.4965 7.9020 31.5900 ;
      RECT 7.7680 30.4965 7.7940 31.5900 ;
      RECT 7.6600 30.4965 7.6860 31.5900 ;
      RECT 7.5520 30.4965 7.5780 31.5900 ;
      RECT 7.4440 30.4965 7.4700 31.5900 ;
      RECT 7.3360 30.4965 7.3620 31.5900 ;
      RECT 7.2280 30.4965 7.2540 31.5900 ;
      RECT 7.1200 30.4965 7.1460 31.5900 ;
      RECT 7.0120 30.4965 7.0380 31.5900 ;
      RECT 6.9040 30.4965 6.9300 31.5900 ;
      RECT 6.7960 30.4965 6.8220 31.5900 ;
      RECT 6.6880 30.4965 6.7140 31.5900 ;
      RECT 6.5800 30.4965 6.6060 31.5900 ;
      RECT 6.4720 30.4965 6.4980 31.5900 ;
      RECT 6.3640 30.4965 6.3900 31.5900 ;
      RECT 6.2560 30.4965 6.2820 31.5900 ;
      RECT 6.1480 30.4965 6.1740 31.5900 ;
      RECT 6.0400 30.4965 6.0660 31.5900 ;
      RECT 5.9320 30.4965 5.9580 31.5900 ;
      RECT 5.8240 30.4965 5.8500 31.5900 ;
      RECT 5.7160 30.4965 5.7420 31.5900 ;
      RECT 5.6080 30.4965 5.6340 31.5900 ;
      RECT 5.5000 30.4965 5.5260 31.5900 ;
      RECT 5.3920 30.4965 5.4180 31.5900 ;
      RECT 5.2840 30.4965 5.3100 31.5900 ;
      RECT 5.1760 30.4965 5.2020 31.5900 ;
      RECT 5.0680 30.4965 5.0940 31.5900 ;
      RECT 4.9600 30.4965 4.9860 31.5900 ;
      RECT 4.8520 30.4965 4.8780 31.5900 ;
      RECT 4.7440 30.4965 4.7700 31.5900 ;
      RECT 4.6360 30.4965 4.6620 31.5900 ;
      RECT 4.5280 30.4965 4.5540 31.5900 ;
      RECT 4.4200 30.4965 4.4460 31.5900 ;
      RECT 4.3120 30.4965 4.3380 31.5900 ;
      RECT 4.2040 30.4965 4.2300 31.5900 ;
      RECT 4.0960 30.4965 4.1220 31.5900 ;
      RECT 3.9880 30.4965 4.0140 31.5900 ;
      RECT 3.8800 30.4965 3.9060 31.5900 ;
      RECT 3.7720 30.4965 3.7980 31.5900 ;
      RECT 3.6640 30.4965 3.6900 31.5900 ;
      RECT 3.5560 30.4965 3.5820 31.5900 ;
      RECT 3.4480 30.4965 3.4740 31.5900 ;
      RECT 3.3400 30.4965 3.3660 31.5900 ;
      RECT 3.2320 30.4965 3.2580 31.5900 ;
      RECT 3.1240 30.4965 3.1500 31.5900 ;
      RECT 3.0160 30.4965 3.0420 31.5900 ;
      RECT 2.9080 30.4965 2.9340 31.5900 ;
      RECT 2.8000 30.4965 2.8260 31.5900 ;
      RECT 2.6920 30.4965 2.7180 31.5900 ;
      RECT 2.5840 30.4965 2.6100 31.5900 ;
      RECT 2.4760 30.4965 2.5020 31.5900 ;
      RECT 2.3680 30.4965 2.3940 31.5900 ;
      RECT 2.2600 30.4965 2.2860 31.5900 ;
      RECT 2.1520 30.4965 2.1780 31.5900 ;
      RECT 2.0440 30.4965 2.0700 31.5900 ;
      RECT 1.9360 30.4965 1.9620 31.5900 ;
      RECT 1.8280 30.4965 1.8540 31.5900 ;
      RECT 1.7200 30.4965 1.7460 31.5900 ;
      RECT 1.6120 30.4965 1.6380 31.5900 ;
      RECT 1.5040 30.4965 1.5300 31.5900 ;
      RECT 1.3960 30.4965 1.4220 31.5900 ;
      RECT 1.2880 30.4965 1.3140 31.5900 ;
      RECT 1.1800 30.4965 1.2060 31.5900 ;
      RECT 1.0720 30.4965 1.0980 31.5900 ;
      RECT 0.9640 30.4965 0.9900 31.5900 ;
      RECT 0.8560 30.4965 0.8820 31.5900 ;
      RECT 0.7480 30.4965 0.7740 31.5900 ;
      RECT 0.6400 30.4965 0.6660 31.5900 ;
      RECT 0.5320 30.4965 0.5580 31.5900 ;
      RECT 0.4240 30.4965 0.4500 31.5900 ;
      RECT 0.3160 30.4965 0.3420 31.5900 ;
      RECT 0.2080 30.4965 0.2340 31.5900 ;
      RECT 0.0050 30.4965 0.0900 31.5900 ;
      RECT 15.5530 31.5765 15.6810 32.6700 ;
      RECT 15.5390 32.2420 15.6810 32.5645 ;
      RECT 15.3190 31.9690 15.4530 32.6700 ;
      RECT 15.2960 32.3040 15.4530 32.5620 ;
      RECT 15.3190 31.5765 15.4170 32.6700 ;
      RECT 15.3190 31.6975 15.4310 31.9370 ;
      RECT 15.3190 31.5765 15.4530 31.6655 ;
      RECT 15.0940 32.0270 15.2280 32.6700 ;
      RECT 15.0940 31.5765 15.1920 32.6700 ;
      RECT 14.6770 31.5765 14.7600 32.6700 ;
      RECT 14.6770 31.6650 14.7740 32.6005 ;
      RECT 30.2680 31.5765 30.3530 32.6700 ;
      RECT 30.1240 31.5765 30.1500 32.6700 ;
      RECT 30.0160 31.5765 30.0420 32.6700 ;
      RECT 29.9080 31.5765 29.9340 32.6700 ;
      RECT 29.8000 31.5765 29.8260 32.6700 ;
      RECT 29.6920 31.5765 29.7180 32.6700 ;
      RECT 29.5840 31.5765 29.6100 32.6700 ;
      RECT 29.4760 31.5765 29.5020 32.6700 ;
      RECT 29.3680 31.5765 29.3940 32.6700 ;
      RECT 29.2600 31.5765 29.2860 32.6700 ;
      RECT 29.1520 31.5765 29.1780 32.6700 ;
      RECT 29.0440 31.5765 29.0700 32.6700 ;
      RECT 28.9360 31.5765 28.9620 32.6700 ;
      RECT 28.8280 31.5765 28.8540 32.6700 ;
      RECT 28.7200 31.5765 28.7460 32.6700 ;
      RECT 28.6120 31.5765 28.6380 32.6700 ;
      RECT 28.5040 31.5765 28.5300 32.6700 ;
      RECT 28.3960 31.5765 28.4220 32.6700 ;
      RECT 28.2880 31.5765 28.3140 32.6700 ;
      RECT 28.1800 31.5765 28.2060 32.6700 ;
      RECT 28.0720 31.5765 28.0980 32.6700 ;
      RECT 27.9640 31.5765 27.9900 32.6700 ;
      RECT 27.8560 31.5765 27.8820 32.6700 ;
      RECT 27.7480 31.5765 27.7740 32.6700 ;
      RECT 27.6400 31.5765 27.6660 32.6700 ;
      RECT 27.5320 31.5765 27.5580 32.6700 ;
      RECT 27.4240 31.5765 27.4500 32.6700 ;
      RECT 27.3160 31.5765 27.3420 32.6700 ;
      RECT 27.2080 31.5765 27.2340 32.6700 ;
      RECT 27.1000 31.5765 27.1260 32.6700 ;
      RECT 26.9920 31.5765 27.0180 32.6700 ;
      RECT 26.8840 31.5765 26.9100 32.6700 ;
      RECT 26.7760 31.5765 26.8020 32.6700 ;
      RECT 26.6680 31.5765 26.6940 32.6700 ;
      RECT 26.5600 31.5765 26.5860 32.6700 ;
      RECT 26.4520 31.5765 26.4780 32.6700 ;
      RECT 26.3440 31.5765 26.3700 32.6700 ;
      RECT 26.2360 31.5765 26.2620 32.6700 ;
      RECT 26.1280 31.5765 26.1540 32.6700 ;
      RECT 26.0200 31.5765 26.0460 32.6700 ;
      RECT 25.9120 31.5765 25.9380 32.6700 ;
      RECT 25.8040 31.5765 25.8300 32.6700 ;
      RECT 25.6960 31.5765 25.7220 32.6700 ;
      RECT 25.5880 31.5765 25.6140 32.6700 ;
      RECT 25.4800 31.5765 25.5060 32.6700 ;
      RECT 25.3720 31.5765 25.3980 32.6700 ;
      RECT 25.2640 31.5765 25.2900 32.6700 ;
      RECT 25.1560 31.5765 25.1820 32.6700 ;
      RECT 25.0480 31.5765 25.0740 32.6700 ;
      RECT 24.9400 31.5765 24.9660 32.6700 ;
      RECT 24.8320 31.5765 24.8580 32.6700 ;
      RECT 24.7240 31.5765 24.7500 32.6700 ;
      RECT 24.6160 31.5765 24.6420 32.6700 ;
      RECT 24.5080 31.5765 24.5340 32.6700 ;
      RECT 24.4000 31.5765 24.4260 32.6700 ;
      RECT 24.2920 31.5765 24.3180 32.6700 ;
      RECT 24.1840 31.5765 24.2100 32.6700 ;
      RECT 24.0760 31.5765 24.1020 32.6700 ;
      RECT 23.9680 31.5765 23.9940 32.6700 ;
      RECT 23.8600 31.5765 23.8860 32.6700 ;
      RECT 23.7520 31.5765 23.7780 32.6700 ;
      RECT 23.6440 31.5765 23.6700 32.6700 ;
      RECT 23.5360 31.5765 23.5620 32.6700 ;
      RECT 23.4280 31.5765 23.4540 32.6700 ;
      RECT 23.3200 31.5765 23.3460 32.6700 ;
      RECT 23.2120 31.5765 23.2380 32.6700 ;
      RECT 23.1040 31.5765 23.1300 32.6700 ;
      RECT 22.9960 31.5765 23.0220 32.6700 ;
      RECT 22.8880 31.5765 22.9140 32.6700 ;
      RECT 22.7800 31.5765 22.8060 32.6700 ;
      RECT 22.6720 31.5765 22.6980 32.6700 ;
      RECT 22.5640 31.5765 22.5900 32.6700 ;
      RECT 22.4560 31.5765 22.4820 32.6700 ;
      RECT 22.3480 31.5765 22.3740 32.6700 ;
      RECT 22.2400 31.5765 22.2660 32.6700 ;
      RECT 22.1320 31.5765 22.1580 32.6700 ;
      RECT 22.0240 31.5765 22.0500 32.6700 ;
      RECT 21.9160 31.5765 21.9420 32.6700 ;
      RECT 21.8080 31.5765 21.8340 32.6700 ;
      RECT 21.7000 31.5765 21.7260 32.6700 ;
      RECT 21.5920 31.5765 21.6180 32.6700 ;
      RECT 21.4840 31.5765 21.5100 32.6700 ;
      RECT 21.3760 31.5765 21.4020 32.6700 ;
      RECT 21.2680 31.5765 21.2940 32.6700 ;
      RECT 21.1600 31.5765 21.1860 32.6700 ;
      RECT 21.0520 31.5765 21.0780 32.6700 ;
      RECT 20.9440 31.5765 20.9700 32.6700 ;
      RECT 20.8360 31.5765 20.8620 32.6700 ;
      RECT 20.7280 31.5765 20.7540 32.6700 ;
      RECT 20.6200 31.5765 20.6460 32.6700 ;
      RECT 20.5120 31.5765 20.5380 32.6700 ;
      RECT 20.4040 31.5765 20.4300 32.6700 ;
      RECT 20.2960 31.5765 20.3220 32.6700 ;
      RECT 20.1880 31.5765 20.2140 32.6700 ;
      RECT 20.0800 31.5765 20.1060 32.6700 ;
      RECT 19.9720 31.5765 19.9980 32.6700 ;
      RECT 19.8640 31.5765 19.8900 32.6700 ;
      RECT 19.7560 31.5765 19.7820 32.6700 ;
      RECT 19.6480 31.5765 19.6740 32.6700 ;
      RECT 19.5400 31.5765 19.5660 32.6700 ;
      RECT 19.4320 31.5765 19.4580 32.6700 ;
      RECT 19.3240 31.5765 19.3500 32.6700 ;
      RECT 19.2160 31.5765 19.2420 32.6700 ;
      RECT 19.1080 31.5765 19.1340 32.6700 ;
      RECT 19.0000 31.5765 19.0260 32.6700 ;
      RECT 18.8920 31.5765 18.9180 32.6700 ;
      RECT 18.7840 31.5765 18.8100 32.6700 ;
      RECT 18.6760 31.5765 18.7020 32.6700 ;
      RECT 18.5680 31.5765 18.5940 32.6700 ;
      RECT 18.4600 31.5765 18.4860 32.6700 ;
      RECT 18.3520 31.5765 18.3780 32.6700 ;
      RECT 18.2440 31.5765 18.2700 32.6700 ;
      RECT 18.1360 31.5765 18.1620 32.6700 ;
      RECT 18.0280 31.5765 18.0540 32.6700 ;
      RECT 17.9200 31.5765 17.9460 32.6700 ;
      RECT 17.8120 31.5765 17.8380 32.6700 ;
      RECT 17.7040 31.5765 17.7300 32.6700 ;
      RECT 17.5960 31.5765 17.6220 32.6700 ;
      RECT 17.4880 31.5765 17.5140 32.6700 ;
      RECT 17.3800 31.5765 17.4060 32.6700 ;
      RECT 17.2720 31.5765 17.2980 32.6700 ;
      RECT 17.1640 31.5765 17.1900 32.6700 ;
      RECT 17.0560 31.5765 17.0820 32.6700 ;
      RECT 16.9480 31.5765 16.9740 32.6700 ;
      RECT 16.8400 31.5765 16.8660 32.6700 ;
      RECT 16.7320 31.5765 16.7580 32.6700 ;
      RECT 16.6240 31.5765 16.6500 32.6700 ;
      RECT 16.5160 31.5765 16.5420 32.6700 ;
      RECT 16.4080 31.5765 16.4340 32.6700 ;
      RECT 16.3000 31.5765 16.3260 32.6700 ;
      RECT 16.0870 31.5765 16.1640 32.6700 ;
      RECT 14.1940 31.5765 14.2710 32.6700 ;
      RECT 14.0320 31.5765 14.0580 32.6700 ;
      RECT 13.9240 31.5765 13.9500 32.6700 ;
      RECT 13.8160 31.5765 13.8420 32.6700 ;
      RECT 13.7080 31.5765 13.7340 32.6700 ;
      RECT 13.6000 31.5765 13.6260 32.6700 ;
      RECT 13.4920 31.5765 13.5180 32.6700 ;
      RECT 13.3840 31.5765 13.4100 32.6700 ;
      RECT 13.2760 31.5765 13.3020 32.6700 ;
      RECT 13.1680 31.5765 13.1940 32.6700 ;
      RECT 13.0600 31.5765 13.0860 32.6700 ;
      RECT 12.9520 31.5765 12.9780 32.6700 ;
      RECT 12.8440 31.5765 12.8700 32.6700 ;
      RECT 12.7360 31.5765 12.7620 32.6700 ;
      RECT 12.6280 31.5765 12.6540 32.6700 ;
      RECT 12.5200 31.5765 12.5460 32.6700 ;
      RECT 12.4120 31.5765 12.4380 32.6700 ;
      RECT 12.3040 31.5765 12.3300 32.6700 ;
      RECT 12.1960 31.5765 12.2220 32.6700 ;
      RECT 12.0880 31.5765 12.1140 32.6700 ;
      RECT 11.9800 31.5765 12.0060 32.6700 ;
      RECT 11.8720 31.5765 11.8980 32.6700 ;
      RECT 11.7640 31.5765 11.7900 32.6700 ;
      RECT 11.6560 31.5765 11.6820 32.6700 ;
      RECT 11.5480 31.5765 11.5740 32.6700 ;
      RECT 11.4400 31.5765 11.4660 32.6700 ;
      RECT 11.3320 31.5765 11.3580 32.6700 ;
      RECT 11.2240 31.5765 11.2500 32.6700 ;
      RECT 11.1160 31.5765 11.1420 32.6700 ;
      RECT 11.0080 31.5765 11.0340 32.6700 ;
      RECT 10.9000 31.5765 10.9260 32.6700 ;
      RECT 10.7920 31.5765 10.8180 32.6700 ;
      RECT 10.6840 31.5765 10.7100 32.6700 ;
      RECT 10.5760 31.5765 10.6020 32.6700 ;
      RECT 10.4680 31.5765 10.4940 32.6700 ;
      RECT 10.3600 31.5765 10.3860 32.6700 ;
      RECT 10.2520 31.5765 10.2780 32.6700 ;
      RECT 10.1440 31.5765 10.1700 32.6700 ;
      RECT 10.0360 31.5765 10.0620 32.6700 ;
      RECT 9.9280 31.5765 9.9540 32.6700 ;
      RECT 9.8200 31.5765 9.8460 32.6700 ;
      RECT 9.7120 31.5765 9.7380 32.6700 ;
      RECT 9.6040 31.5765 9.6300 32.6700 ;
      RECT 9.4960 31.5765 9.5220 32.6700 ;
      RECT 9.3880 31.5765 9.4140 32.6700 ;
      RECT 9.2800 31.5765 9.3060 32.6700 ;
      RECT 9.1720 31.5765 9.1980 32.6700 ;
      RECT 9.0640 31.5765 9.0900 32.6700 ;
      RECT 8.9560 31.5765 8.9820 32.6700 ;
      RECT 8.8480 31.5765 8.8740 32.6700 ;
      RECT 8.7400 31.5765 8.7660 32.6700 ;
      RECT 8.6320 31.5765 8.6580 32.6700 ;
      RECT 8.5240 31.5765 8.5500 32.6700 ;
      RECT 8.4160 31.5765 8.4420 32.6700 ;
      RECT 8.3080 31.5765 8.3340 32.6700 ;
      RECT 8.2000 31.5765 8.2260 32.6700 ;
      RECT 8.0920 31.5765 8.1180 32.6700 ;
      RECT 7.9840 31.5765 8.0100 32.6700 ;
      RECT 7.8760 31.5765 7.9020 32.6700 ;
      RECT 7.7680 31.5765 7.7940 32.6700 ;
      RECT 7.6600 31.5765 7.6860 32.6700 ;
      RECT 7.5520 31.5765 7.5780 32.6700 ;
      RECT 7.4440 31.5765 7.4700 32.6700 ;
      RECT 7.3360 31.5765 7.3620 32.6700 ;
      RECT 7.2280 31.5765 7.2540 32.6700 ;
      RECT 7.1200 31.5765 7.1460 32.6700 ;
      RECT 7.0120 31.5765 7.0380 32.6700 ;
      RECT 6.9040 31.5765 6.9300 32.6700 ;
      RECT 6.7960 31.5765 6.8220 32.6700 ;
      RECT 6.6880 31.5765 6.7140 32.6700 ;
      RECT 6.5800 31.5765 6.6060 32.6700 ;
      RECT 6.4720 31.5765 6.4980 32.6700 ;
      RECT 6.3640 31.5765 6.3900 32.6700 ;
      RECT 6.2560 31.5765 6.2820 32.6700 ;
      RECT 6.1480 31.5765 6.1740 32.6700 ;
      RECT 6.0400 31.5765 6.0660 32.6700 ;
      RECT 5.9320 31.5765 5.9580 32.6700 ;
      RECT 5.8240 31.5765 5.8500 32.6700 ;
      RECT 5.7160 31.5765 5.7420 32.6700 ;
      RECT 5.6080 31.5765 5.6340 32.6700 ;
      RECT 5.5000 31.5765 5.5260 32.6700 ;
      RECT 5.3920 31.5765 5.4180 32.6700 ;
      RECT 5.2840 31.5765 5.3100 32.6700 ;
      RECT 5.1760 31.5765 5.2020 32.6700 ;
      RECT 5.0680 31.5765 5.0940 32.6700 ;
      RECT 4.9600 31.5765 4.9860 32.6700 ;
      RECT 4.8520 31.5765 4.8780 32.6700 ;
      RECT 4.7440 31.5765 4.7700 32.6700 ;
      RECT 4.6360 31.5765 4.6620 32.6700 ;
      RECT 4.5280 31.5765 4.5540 32.6700 ;
      RECT 4.4200 31.5765 4.4460 32.6700 ;
      RECT 4.3120 31.5765 4.3380 32.6700 ;
      RECT 4.2040 31.5765 4.2300 32.6700 ;
      RECT 4.0960 31.5765 4.1220 32.6700 ;
      RECT 3.9880 31.5765 4.0140 32.6700 ;
      RECT 3.8800 31.5765 3.9060 32.6700 ;
      RECT 3.7720 31.5765 3.7980 32.6700 ;
      RECT 3.6640 31.5765 3.6900 32.6700 ;
      RECT 3.5560 31.5765 3.5820 32.6700 ;
      RECT 3.4480 31.5765 3.4740 32.6700 ;
      RECT 3.3400 31.5765 3.3660 32.6700 ;
      RECT 3.2320 31.5765 3.2580 32.6700 ;
      RECT 3.1240 31.5765 3.1500 32.6700 ;
      RECT 3.0160 31.5765 3.0420 32.6700 ;
      RECT 2.9080 31.5765 2.9340 32.6700 ;
      RECT 2.8000 31.5765 2.8260 32.6700 ;
      RECT 2.6920 31.5765 2.7180 32.6700 ;
      RECT 2.5840 31.5765 2.6100 32.6700 ;
      RECT 2.4760 31.5765 2.5020 32.6700 ;
      RECT 2.3680 31.5765 2.3940 32.6700 ;
      RECT 2.2600 31.5765 2.2860 32.6700 ;
      RECT 2.1520 31.5765 2.1780 32.6700 ;
      RECT 2.0440 31.5765 2.0700 32.6700 ;
      RECT 1.9360 31.5765 1.9620 32.6700 ;
      RECT 1.8280 31.5765 1.8540 32.6700 ;
      RECT 1.7200 31.5765 1.7460 32.6700 ;
      RECT 1.6120 31.5765 1.6380 32.6700 ;
      RECT 1.5040 31.5765 1.5300 32.6700 ;
      RECT 1.3960 31.5765 1.4220 32.6700 ;
      RECT 1.2880 31.5765 1.3140 32.6700 ;
      RECT 1.1800 31.5765 1.2060 32.6700 ;
      RECT 1.0720 31.5765 1.0980 32.6700 ;
      RECT 0.9640 31.5765 0.9900 32.6700 ;
      RECT 0.8560 31.5765 0.8820 32.6700 ;
      RECT 0.7480 31.5765 0.7740 32.6700 ;
      RECT 0.6400 31.5765 0.6660 32.6700 ;
      RECT 0.5320 31.5765 0.5580 32.6700 ;
      RECT 0.4240 31.5765 0.4500 32.6700 ;
      RECT 0.3160 31.5765 0.3420 32.6700 ;
      RECT 0.2080 31.5765 0.2340 32.6700 ;
      RECT 0.0050 31.5765 0.0900 32.6700 ;
      RECT 15.5530 32.6565 15.6810 33.7500 ;
      RECT 15.5390 33.3220 15.6810 33.6445 ;
      RECT 15.3190 33.0490 15.4530 33.7500 ;
      RECT 15.2960 33.3840 15.4530 33.6420 ;
      RECT 15.3190 32.6565 15.4170 33.7500 ;
      RECT 15.3190 32.7775 15.4310 33.0170 ;
      RECT 15.3190 32.6565 15.4530 32.7455 ;
      RECT 15.0940 33.1070 15.2280 33.7500 ;
      RECT 15.0940 32.6565 15.1920 33.7500 ;
      RECT 14.6770 32.6565 14.7600 33.7500 ;
      RECT 14.6770 32.7450 14.7740 33.6805 ;
      RECT 30.2680 32.6565 30.3530 33.7500 ;
      RECT 30.1240 32.6565 30.1500 33.7500 ;
      RECT 30.0160 32.6565 30.0420 33.7500 ;
      RECT 29.9080 32.6565 29.9340 33.7500 ;
      RECT 29.8000 32.6565 29.8260 33.7500 ;
      RECT 29.6920 32.6565 29.7180 33.7500 ;
      RECT 29.5840 32.6565 29.6100 33.7500 ;
      RECT 29.4760 32.6565 29.5020 33.7500 ;
      RECT 29.3680 32.6565 29.3940 33.7500 ;
      RECT 29.2600 32.6565 29.2860 33.7500 ;
      RECT 29.1520 32.6565 29.1780 33.7500 ;
      RECT 29.0440 32.6565 29.0700 33.7500 ;
      RECT 28.9360 32.6565 28.9620 33.7500 ;
      RECT 28.8280 32.6565 28.8540 33.7500 ;
      RECT 28.7200 32.6565 28.7460 33.7500 ;
      RECT 28.6120 32.6565 28.6380 33.7500 ;
      RECT 28.5040 32.6565 28.5300 33.7500 ;
      RECT 28.3960 32.6565 28.4220 33.7500 ;
      RECT 28.2880 32.6565 28.3140 33.7500 ;
      RECT 28.1800 32.6565 28.2060 33.7500 ;
      RECT 28.0720 32.6565 28.0980 33.7500 ;
      RECT 27.9640 32.6565 27.9900 33.7500 ;
      RECT 27.8560 32.6565 27.8820 33.7500 ;
      RECT 27.7480 32.6565 27.7740 33.7500 ;
      RECT 27.6400 32.6565 27.6660 33.7500 ;
      RECT 27.5320 32.6565 27.5580 33.7500 ;
      RECT 27.4240 32.6565 27.4500 33.7500 ;
      RECT 27.3160 32.6565 27.3420 33.7500 ;
      RECT 27.2080 32.6565 27.2340 33.7500 ;
      RECT 27.1000 32.6565 27.1260 33.7500 ;
      RECT 26.9920 32.6565 27.0180 33.7500 ;
      RECT 26.8840 32.6565 26.9100 33.7500 ;
      RECT 26.7760 32.6565 26.8020 33.7500 ;
      RECT 26.6680 32.6565 26.6940 33.7500 ;
      RECT 26.5600 32.6565 26.5860 33.7500 ;
      RECT 26.4520 32.6565 26.4780 33.7500 ;
      RECT 26.3440 32.6565 26.3700 33.7500 ;
      RECT 26.2360 32.6565 26.2620 33.7500 ;
      RECT 26.1280 32.6565 26.1540 33.7500 ;
      RECT 26.0200 32.6565 26.0460 33.7500 ;
      RECT 25.9120 32.6565 25.9380 33.7500 ;
      RECT 25.8040 32.6565 25.8300 33.7500 ;
      RECT 25.6960 32.6565 25.7220 33.7500 ;
      RECT 25.5880 32.6565 25.6140 33.7500 ;
      RECT 25.4800 32.6565 25.5060 33.7500 ;
      RECT 25.3720 32.6565 25.3980 33.7500 ;
      RECT 25.2640 32.6565 25.2900 33.7500 ;
      RECT 25.1560 32.6565 25.1820 33.7500 ;
      RECT 25.0480 32.6565 25.0740 33.7500 ;
      RECT 24.9400 32.6565 24.9660 33.7500 ;
      RECT 24.8320 32.6565 24.8580 33.7500 ;
      RECT 24.7240 32.6565 24.7500 33.7500 ;
      RECT 24.6160 32.6565 24.6420 33.7500 ;
      RECT 24.5080 32.6565 24.5340 33.7500 ;
      RECT 24.4000 32.6565 24.4260 33.7500 ;
      RECT 24.2920 32.6565 24.3180 33.7500 ;
      RECT 24.1840 32.6565 24.2100 33.7500 ;
      RECT 24.0760 32.6565 24.1020 33.7500 ;
      RECT 23.9680 32.6565 23.9940 33.7500 ;
      RECT 23.8600 32.6565 23.8860 33.7500 ;
      RECT 23.7520 32.6565 23.7780 33.7500 ;
      RECT 23.6440 32.6565 23.6700 33.7500 ;
      RECT 23.5360 32.6565 23.5620 33.7500 ;
      RECT 23.4280 32.6565 23.4540 33.7500 ;
      RECT 23.3200 32.6565 23.3460 33.7500 ;
      RECT 23.2120 32.6565 23.2380 33.7500 ;
      RECT 23.1040 32.6565 23.1300 33.7500 ;
      RECT 22.9960 32.6565 23.0220 33.7500 ;
      RECT 22.8880 32.6565 22.9140 33.7500 ;
      RECT 22.7800 32.6565 22.8060 33.7500 ;
      RECT 22.6720 32.6565 22.6980 33.7500 ;
      RECT 22.5640 32.6565 22.5900 33.7500 ;
      RECT 22.4560 32.6565 22.4820 33.7500 ;
      RECT 22.3480 32.6565 22.3740 33.7500 ;
      RECT 22.2400 32.6565 22.2660 33.7500 ;
      RECT 22.1320 32.6565 22.1580 33.7500 ;
      RECT 22.0240 32.6565 22.0500 33.7500 ;
      RECT 21.9160 32.6565 21.9420 33.7500 ;
      RECT 21.8080 32.6565 21.8340 33.7500 ;
      RECT 21.7000 32.6565 21.7260 33.7500 ;
      RECT 21.5920 32.6565 21.6180 33.7500 ;
      RECT 21.4840 32.6565 21.5100 33.7500 ;
      RECT 21.3760 32.6565 21.4020 33.7500 ;
      RECT 21.2680 32.6565 21.2940 33.7500 ;
      RECT 21.1600 32.6565 21.1860 33.7500 ;
      RECT 21.0520 32.6565 21.0780 33.7500 ;
      RECT 20.9440 32.6565 20.9700 33.7500 ;
      RECT 20.8360 32.6565 20.8620 33.7500 ;
      RECT 20.7280 32.6565 20.7540 33.7500 ;
      RECT 20.6200 32.6565 20.6460 33.7500 ;
      RECT 20.5120 32.6565 20.5380 33.7500 ;
      RECT 20.4040 32.6565 20.4300 33.7500 ;
      RECT 20.2960 32.6565 20.3220 33.7500 ;
      RECT 20.1880 32.6565 20.2140 33.7500 ;
      RECT 20.0800 32.6565 20.1060 33.7500 ;
      RECT 19.9720 32.6565 19.9980 33.7500 ;
      RECT 19.8640 32.6565 19.8900 33.7500 ;
      RECT 19.7560 32.6565 19.7820 33.7500 ;
      RECT 19.6480 32.6565 19.6740 33.7500 ;
      RECT 19.5400 32.6565 19.5660 33.7500 ;
      RECT 19.4320 32.6565 19.4580 33.7500 ;
      RECT 19.3240 32.6565 19.3500 33.7500 ;
      RECT 19.2160 32.6565 19.2420 33.7500 ;
      RECT 19.1080 32.6565 19.1340 33.7500 ;
      RECT 19.0000 32.6565 19.0260 33.7500 ;
      RECT 18.8920 32.6565 18.9180 33.7500 ;
      RECT 18.7840 32.6565 18.8100 33.7500 ;
      RECT 18.6760 32.6565 18.7020 33.7500 ;
      RECT 18.5680 32.6565 18.5940 33.7500 ;
      RECT 18.4600 32.6565 18.4860 33.7500 ;
      RECT 18.3520 32.6565 18.3780 33.7500 ;
      RECT 18.2440 32.6565 18.2700 33.7500 ;
      RECT 18.1360 32.6565 18.1620 33.7500 ;
      RECT 18.0280 32.6565 18.0540 33.7500 ;
      RECT 17.9200 32.6565 17.9460 33.7500 ;
      RECT 17.8120 32.6565 17.8380 33.7500 ;
      RECT 17.7040 32.6565 17.7300 33.7500 ;
      RECT 17.5960 32.6565 17.6220 33.7500 ;
      RECT 17.4880 32.6565 17.5140 33.7500 ;
      RECT 17.3800 32.6565 17.4060 33.7500 ;
      RECT 17.2720 32.6565 17.2980 33.7500 ;
      RECT 17.1640 32.6565 17.1900 33.7500 ;
      RECT 17.0560 32.6565 17.0820 33.7500 ;
      RECT 16.9480 32.6565 16.9740 33.7500 ;
      RECT 16.8400 32.6565 16.8660 33.7500 ;
      RECT 16.7320 32.6565 16.7580 33.7500 ;
      RECT 16.6240 32.6565 16.6500 33.7500 ;
      RECT 16.5160 32.6565 16.5420 33.7500 ;
      RECT 16.4080 32.6565 16.4340 33.7500 ;
      RECT 16.3000 32.6565 16.3260 33.7500 ;
      RECT 16.0870 32.6565 16.1640 33.7500 ;
      RECT 14.1940 32.6565 14.2710 33.7500 ;
      RECT 14.0320 32.6565 14.0580 33.7500 ;
      RECT 13.9240 32.6565 13.9500 33.7500 ;
      RECT 13.8160 32.6565 13.8420 33.7500 ;
      RECT 13.7080 32.6565 13.7340 33.7500 ;
      RECT 13.6000 32.6565 13.6260 33.7500 ;
      RECT 13.4920 32.6565 13.5180 33.7500 ;
      RECT 13.3840 32.6565 13.4100 33.7500 ;
      RECT 13.2760 32.6565 13.3020 33.7500 ;
      RECT 13.1680 32.6565 13.1940 33.7500 ;
      RECT 13.0600 32.6565 13.0860 33.7500 ;
      RECT 12.9520 32.6565 12.9780 33.7500 ;
      RECT 12.8440 32.6565 12.8700 33.7500 ;
      RECT 12.7360 32.6565 12.7620 33.7500 ;
      RECT 12.6280 32.6565 12.6540 33.7500 ;
      RECT 12.5200 32.6565 12.5460 33.7500 ;
      RECT 12.4120 32.6565 12.4380 33.7500 ;
      RECT 12.3040 32.6565 12.3300 33.7500 ;
      RECT 12.1960 32.6565 12.2220 33.7500 ;
      RECT 12.0880 32.6565 12.1140 33.7500 ;
      RECT 11.9800 32.6565 12.0060 33.7500 ;
      RECT 11.8720 32.6565 11.8980 33.7500 ;
      RECT 11.7640 32.6565 11.7900 33.7500 ;
      RECT 11.6560 32.6565 11.6820 33.7500 ;
      RECT 11.5480 32.6565 11.5740 33.7500 ;
      RECT 11.4400 32.6565 11.4660 33.7500 ;
      RECT 11.3320 32.6565 11.3580 33.7500 ;
      RECT 11.2240 32.6565 11.2500 33.7500 ;
      RECT 11.1160 32.6565 11.1420 33.7500 ;
      RECT 11.0080 32.6565 11.0340 33.7500 ;
      RECT 10.9000 32.6565 10.9260 33.7500 ;
      RECT 10.7920 32.6565 10.8180 33.7500 ;
      RECT 10.6840 32.6565 10.7100 33.7500 ;
      RECT 10.5760 32.6565 10.6020 33.7500 ;
      RECT 10.4680 32.6565 10.4940 33.7500 ;
      RECT 10.3600 32.6565 10.3860 33.7500 ;
      RECT 10.2520 32.6565 10.2780 33.7500 ;
      RECT 10.1440 32.6565 10.1700 33.7500 ;
      RECT 10.0360 32.6565 10.0620 33.7500 ;
      RECT 9.9280 32.6565 9.9540 33.7500 ;
      RECT 9.8200 32.6565 9.8460 33.7500 ;
      RECT 9.7120 32.6565 9.7380 33.7500 ;
      RECT 9.6040 32.6565 9.6300 33.7500 ;
      RECT 9.4960 32.6565 9.5220 33.7500 ;
      RECT 9.3880 32.6565 9.4140 33.7500 ;
      RECT 9.2800 32.6565 9.3060 33.7500 ;
      RECT 9.1720 32.6565 9.1980 33.7500 ;
      RECT 9.0640 32.6565 9.0900 33.7500 ;
      RECT 8.9560 32.6565 8.9820 33.7500 ;
      RECT 8.8480 32.6565 8.8740 33.7500 ;
      RECT 8.7400 32.6565 8.7660 33.7500 ;
      RECT 8.6320 32.6565 8.6580 33.7500 ;
      RECT 8.5240 32.6565 8.5500 33.7500 ;
      RECT 8.4160 32.6565 8.4420 33.7500 ;
      RECT 8.3080 32.6565 8.3340 33.7500 ;
      RECT 8.2000 32.6565 8.2260 33.7500 ;
      RECT 8.0920 32.6565 8.1180 33.7500 ;
      RECT 7.9840 32.6565 8.0100 33.7500 ;
      RECT 7.8760 32.6565 7.9020 33.7500 ;
      RECT 7.7680 32.6565 7.7940 33.7500 ;
      RECT 7.6600 32.6565 7.6860 33.7500 ;
      RECT 7.5520 32.6565 7.5780 33.7500 ;
      RECT 7.4440 32.6565 7.4700 33.7500 ;
      RECT 7.3360 32.6565 7.3620 33.7500 ;
      RECT 7.2280 32.6565 7.2540 33.7500 ;
      RECT 7.1200 32.6565 7.1460 33.7500 ;
      RECT 7.0120 32.6565 7.0380 33.7500 ;
      RECT 6.9040 32.6565 6.9300 33.7500 ;
      RECT 6.7960 32.6565 6.8220 33.7500 ;
      RECT 6.6880 32.6565 6.7140 33.7500 ;
      RECT 6.5800 32.6565 6.6060 33.7500 ;
      RECT 6.4720 32.6565 6.4980 33.7500 ;
      RECT 6.3640 32.6565 6.3900 33.7500 ;
      RECT 6.2560 32.6565 6.2820 33.7500 ;
      RECT 6.1480 32.6565 6.1740 33.7500 ;
      RECT 6.0400 32.6565 6.0660 33.7500 ;
      RECT 5.9320 32.6565 5.9580 33.7500 ;
      RECT 5.8240 32.6565 5.8500 33.7500 ;
      RECT 5.7160 32.6565 5.7420 33.7500 ;
      RECT 5.6080 32.6565 5.6340 33.7500 ;
      RECT 5.5000 32.6565 5.5260 33.7500 ;
      RECT 5.3920 32.6565 5.4180 33.7500 ;
      RECT 5.2840 32.6565 5.3100 33.7500 ;
      RECT 5.1760 32.6565 5.2020 33.7500 ;
      RECT 5.0680 32.6565 5.0940 33.7500 ;
      RECT 4.9600 32.6565 4.9860 33.7500 ;
      RECT 4.8520 32.6565 4.8780 33.7500 ;
      RECT 4.7440 32.6565 4.7700 33.7500 ;
      RECT 4.6360 32.6565 4.6620 33.7500 ;
      RECT 4.5280 32.6565 4.5540 33.7500 ;
      RECT 4.4200 32.6565 4.4460 33.7500 ;
      RECT 4.3120 32.6565 4.3380 33.7500 ;
      RECT 4.2040 32.6565 4.2300 33.7500 ;
      RECT 4.0960 32.6565 4.1220 33.7500 ;
      RECT 3.9880 32.6565 4.0140 33.7500 ;
      RECT 3.8800 32.6565 3.9060 33.7500 ;
      RECT 3.7720 32.6565 3.7980 33.7500 ;
      RECT 3.6640 32.6565 3.6900 33.7500 ;
      RECT 3.5560 32.6565 3.5820 33.7500 ;
      RECT 3.4480 32.6565 3.4740 33.7500 ;
      RECT 3.3400 32.6565 3.3660 33.7500 ;
      RECT 3.2320 32.6565 3.2580 33.7500 ;
      RECT 3.1240 32.6565 3.1500 33.7500 ;
      RECT 3.0160 32.6565 3.0420 33.7500 ;
      RECT 2.9080 32.6565 2.9340 33.7500 ;
      RECT 2.8000 32.6565 2.8260 33.7500 ;
      RECT 2.6920 32.6565 2.7180 33.7500 ;
      RECT 2.5840 32.6565 2.6100 33.7500 ;
      RECT 2.4760 32.6565 2.5020 33.7500 ;
      RECT 2.3680 32.6565 2.3940 33.7500 ;
      RECT 2.2600 32.6565 2.2860 33.7500 ;
      RECT 2.1520 32.6565 2.1780 33.7500 ;
      RECT 2.0440 32.6565 2.0700 33.7500 ;
      RECT 1.9360 32.6565 1.9620 33.7500 ;
      RECT 1.8280 32.6565 1.8540 33.7500 ;
      RECT 1.7200 32.6565 1.7460 33.7500 ;
      RECT 1.6120 32.6565 1.6380 33.7500 ;
      RECT 1.5040 32.6565 1.5300 33.7500 ;
      RECT 1.3960 32.6565 1.4220 33.7500 ;
      RECT 1.2880 32.6565 1.3140 33.7500 ;
      RECT 1.1800 32.6565 1.2060 33.7500 ;
      RECT 1.0720 32.6565 1.0980 33.7500 ;
      RECT 0.9640 32.6565 0.9900 33.7500 ;
      RECT 0.8560 32.6565 0.8820 33.7500 ;
      RECT 0.7480 32.6565 0.7740 33.7500 ;
      RECT 0.6400 32.6565 0.6660 33.7500 ;
      RECT 0.5320 32.6565 0.5580 33.7500 ;
      RECT 0.4240 32.6565 0.4500 33.7500 ;
      RECT 0.3160 32.6565 0.3420 33.7500 ;
      RECT 0.2080 32.6565 0.2340 33.7500 ;
      RECT 0.0050 32.6565 0.0900 33.7500 ;
      RECT 15.5530 33.7365 15.6810 34.8300 ;
      RECT 15.5390 34.4020 15.6810 34.7245 ;
      RECT 15.3190 34.1290 15.4530 34.8300 ;
      RECT 15.2960 34.4640 15.4530 34.7220 ;
      RECT 15.3190 33.7365 15.4170 34.8300 ;
      RECT 15.3190 33.8575 15.4310 34.0970 ;
      RECT 15.3190 33.7365 15.4530 33.8255 ;
      RECT 15.0940 34.1870 15.2280 34.8300 ;
      RECT 15.0940 33.7365 15.1920 34.8300 ;
      RECT 14.6770 33.7365 14.7600 34.8300 ;
      RECT 14.6770 33.8250 14.7740 34.7605 ;
      RECT 30.2680 33.7365 30.3530 34.8300 ;
      RECT 30.1240 33.7365 30.1500 34.8300 ;
      RECT 30.0160 33.7365 30.0420 34.8300 ;
      RECT 29.9080 33.7365 29.9340 34.8300 ;
      RECT 29.8000 33.7365 29.8260 34.8300 ;
      RECT 29.6920 33.7365 29.7180 34.8300 ;
      RECT 29.5840 33.7365 29.6100 34.8300 ;
      RECT 29.4760 33.7365 29.5020 34.8300 ;
      RECT 29.3680 33.7365 29.3940 34.8300 ;
      RECT 29.2600 33.7365 29.2860 34.8300 ;
      RECT 29.1520 33.7365 29.1780 34.8300 ;
      RECT 29.0440 33.7365 29.0700 34.8300 ;
      RECT 28.9360 33.7365 28.9620 34.8300 ;
      RECT 28.8280 33.7365 28.8540 34.8300 ;
      RECT 28.7200 33.7365 28.7460 34.8300 ;
      RECT 28.6120 33.7365 28.6380 34.8300 ;
      RECT 28.5040 33.7365 28.5300 34.8300 ;
      RECT 28.3960 33.7365 28.4220 34.8300 ;
      RECT 28.2880 33.7365 28.3140 34.8300 ;
      RECT 28.1800 33.7365 28.2060 34.8300 ;
      RECT 28.0720 33.7365 28.0980 34.8300 ;
      RECT 27.9640 33.7365 27.9900 34.8300 ;
      RECT 27.8560 33.7365 27.8820 34.8300 ;
      RECT 27.7480 33.7365 27.7740 34.8300 ;
      RECT 27.6400 33.7365 27.6660 34.8300 ;
      RECT 27.5320 33.7365 27.5580 34.8300 ;
      RECT 27.4240 33.7365 27.4500 34.8300 ;
      RECT 27.3160 33.7365 27.3420 34.8300 ;
      RECT 27.2080 33.7365 27.2340 34.8300 ;
      RECT 27.1000 33.7365 27.1260 34.8300 ;
      RECT 26.9920 33.7365 27.0180 34.8300 ;
      RECT 26.8840 33.7365 26.9100 34.8300 ;
      RECT 26.7760 33.7365 26.8020 34.8300 ;
      RECT 26.6680 33.7365 26.6940 34.8300 ;
      RECT 26.5600 33.7365 26.5860 34.8300 ;
      RECT 26.4520 33.7365 26.4780 34.8300 ;
      RECT 26.3440 33.7365 26.3700 34.8300 ;
      RECT 26.2360 33.7365 26.2620 34.8300 ;
      RECT 26.1280 33.7365 26.1540 34.8300 ;
      RECT 26.0200 33.7365 26.0460 34.8300 ;
      RECT 25.9120 33.7365 25.9380 34.8300 ;
      RECT 25.8040 33.7365 25.8300 34.8300 ;
      RECT 25.6960 33.7365 25.7220 34.8300 ;
      RECT 25.5880 33.7365 25.6140 34.8300 ;
      RECT 25.4800 33.7365 25.5060 34.8300 ;
      RECT 25.3720 33.7365 25.3980 34.8300 ;
      RECT 25.2640 33.7365 25.2900 34.8300 ;
      RECT 25.1560 33.7365 25.1820 34.8300 ;
      RECT 25.0480 33.7365 25.0740 34.8300 ;
      RECT 24.9400 33.7365 24.9660 34.8300 ;
      RECT 24.8320 33.7365 24.8580 34.8300 ;
      RECT 24.7240 33.7365 24.7500 34.8300 ;
      RECT 24.6160 33.7365 24.6420 34.8300 ;
      RECT 24.5080 33.7365 24.5340 34.8300 ;
      RECT 24.4000 33.7365 24.4260 34.8300 ;
      RECT 24.2920 33.7365 24.3180 34.8300 ;
      RECT 24.1840 33.7365 24.2100 34.8300 ;
      RECT 24.0760 33.7365 24.1020 34.8300 ;
      RECT 23.9680 33.7365 23.9940 34.8300 ;
      RECT 23.8600 33.7365 23.8860 34.8300 ;
      RECT 23.7520 33.7365 23.7780 34.8300 ;
      RECT 23.6440 33.7365 23.6700 34.8300 ;
      RECT 23.5360 33.7365 23.5620 34.8300 ;
      RECT 23.4280 33.7365 23.4540 34.8300 ;
      RECT 23.3200 33.7365 23.3460 34.8300 ;
      RECT 23.2120 33.7365 23.2380 34.8300 ;
      RECT 23.1040 33.7365 23.1300 34.8300 ;
      RECT 22.9960 33.7365 23.0220 34.8300 ;
      RECT 22.8880 33.7365 22.9140 34.8300 ;
      RECT 22.7800 33.7365 22.8060 34.8300 ;
      RECT 22.6720 33.7365 22.6980 34.8300 ;
      RECT 22.5640 33.7365 22.5900 34.8300 ;
      RECT 22.4560 33.7365 22.4820 34.8300 ;
      RECT 22.3480 33.7365 22.3740 34.8300 ;
      RECT 22.2400 33.7365 22.2660 34.8300 ;
      RECT 22.1320 33.7365 22.1580 34.8300 ;
      RECT 22.0240 33.7365 22.0500 34.8300 ;
      RECT 21.9160 33.7365 21.9420 34.8300 ;
      RECT 21.8080 33.7365 21.8340 34.8300 ;
      RECT 21.7000 33.7365 21.7260 34.8300 ;
      RECT 21.5920 33.7365 21.6180 34.8300 ;
      RECT 21.4840 33.7365 21.5100 34.8300 ;
      RECT 21.3760 33.7365 21.4020 34.8300 ;
      RECT 21.2680 33.7365 21.2940 34.8300 ;
      RECT 21.1600 33.7365 21.1860 34.8300 ;
      RECT 21.0520 33.7365 21.0780 34.8300 ;
      RECT 20.9440 33.7365 20.9700 34.8300 ;
      RECT 20.8360 33.7365 20.8620 34.8300 ;
      RECT 20.7280 33.7365 20.7540 34.8300 ;
      RECT 20.6200 33.7365 20.6460 34.8300 ;
      RECT 20.5120 33.7365 20.5380 34.8300 ;
      RECT 20.4040 33.7365 20.4300 34.8300 ;
      RECT 20.2960 33.7365 20.3220 34.8300 ;
      RECT 20.1880 33.7365 20.2140 34.8300 ;
      RECT 20.0800 33.7365 20.1060 34.8300 ;
      RECT 19.9720 33.7365 19.9980 34.8300 ;
      RECT 19.8640 33.7365 19.8900 34.8300 ;
      RECT 19.7560 33.7365 19.7820 34.8300 ;
      RECT 19.6480 33.7365 19.6740 34.8300 ;
      RECT 19.5400 33.7365 19.5660 34.8300 ;
      RECT 19.4320 33.7365 19.4580 34.8300 ;
      RECT 19.3240 33.7365 19.3500 34.8300 ;
      RECT 19.2160 33.7365 19.2420 34.8300 ;
      RECT 19.1080 33.7365 19.1340 34.8300 ;
      RECT 19.0000 33.7365 19.0260 34.8300 ;
      RECT 18.8920 33.7365 18.9180 34.8300 ;
      RECT 18.7840 33.7365 18.8100 34.8300 ;
      RECT 18.6760 33.7365 18.7020 34.8300 ;
      RECT 18.5680 33.7365 18.5940 34.8300 ;
      RECT 18.4600 33.7365 18.4860 34.8300 ;
      RECT 18.3520 33.7365 18.3780 34.8300 ;
      RECT 18.2440 33.7365 18.2700 34.8300 ;
      RECT 18.1360 33.7365 18.1620 34.8300 ;
      RECT 18.0280 33.7365 18.0540 34.8300 ;
      RECT 17.9200 33.7365 17.9460 34.8300 ;
      RECT 17.8120 33.7365 17.8380 34.8300 ;
      RECT 17.7040 33.7365 17.7300 34.8300 ;
      RECT 17.5960 33.7365 17.6220 34.8300 ;
      RECT 17.4880 33.7365 17.5140 34.8300 ;
      RECT 17.3800 33.7365 17.4060 34.8300 ;
      RECT 17.2720 33.7365 17.2980 34.8300 ;
      RECT 17.1640 33.7365 17.1900 34.8300 ;
      RECT 17.0560 33.7365 17.0820 34.8300 ;
      RECT 16.9480 33.7365 16.9740 34.8300 ;
      RECT 16.8400 33.7365 16.8660 34.8300 ;
      RECT 16.7320 33.7365 16.7580 34.8300 ;
      RECT 16.6240 33.7365 16.6500 34.8300 ;
      RECT 16.5160 33.7365 16.5420 34.8300 ;
      RECT 16.4080 33.7365 16.4340 34.8300 ;
      RECT 16.3000 33.7365 16.3260 34.8300 ;
      RECT 16.0870 33.7365 16.1640 34.8300 ;
      RECT 14.1940 33.7365 14.2710 34.8300 ;
      RECT 14.0320 33.7365 14.0580 34.8300 ;
      RECT 13.9240 33.7365 13.9500 34.8300 ;
      RECT 13.8160 33.7365 13.8420 34.8300 ;
      RECT 13.7080 33.7365 13.7340 34.8300 ;
      RECT 13.6000 33.7365 13.6260 34.8300 ;
      RECT 13.4920 33.7365 13.5180 34.8300 ;
      RECT 13.3840 33.7365 13.4100 34.8300 ;
      RECT 13.2760 33.7365 13.3020 34.8300 ;
      RECT 13.1680 33.7365 13.1940 34.8300 ;
      RECT 13.0600 33.7365 13.0860 34.8300 ;
      RECT 12.9520 33.7365 12.9780 34.8300 ;
      RECT 12.8440 33.7365 12.8700 34.8300 ;
      RECT 12.7360 33.7365 12.7620 34.8300 ;
      RECT 12.6280 33.7365 12.6540 34.8300 ;
      RECT 12.5200 33.7365 12.5460 34.8300 ;
      RECT 12.4120 33.7365 12.4380 34.8300 ;
      RECT 12.3040 33.7365 12.3300 34.8300 ;
      RECT 12.1960 33.7365 12.2220 34.8300 ;
      RECT 12.0880 33.7365 12.1140 34.8300 ;
      RECT 11.9800 33.7365 12.0060 34.8300 ;
      RECT 11.8720 33.7365 11.8980 34.8300 ;
      RECT 11.7640 33.7365 11.7900 34.8300 ;
      RECT 11.6560 33.7365 11.6820 34.8300 ;
      RECT 11.5480 33.7365 11.5740 34.8300 ;
      RECT 11.4400 33.7365 11.4660 34.8300 ;
      RECT 11.3320 33.7365 11.3580 34.8300 ;
      RECT 11.2240 33.7365 11.2500 34.8300 ;
      RECT 11.1160 33.7365 11.1420 34.8300 ;
      RECT 11.0080 33.7365 11.0340 34.8300 ;
      RECT 10.9000 33.7365 10.9260 34.8300 ;
      RECT 10.7920 33.7365 10.8180 34.8300 ;
      RECT 10.6840 33.7365 10.7100 34.8300 ;
      RECT 10.5760 33.7365 10.6020 34.8300 ;
      RECT 10.4680 33.7365 10.4940 34.8300 ;
      RECT 10.3600 33.7365 10.3860 34.8300 ;
      RECT 10.2520 33.7365 10.2780 34.8300 ;
      RECT 10.1440 33.7365 10.1700 34.8300 ;
      RECT 10.0360 33.7365 10.0620 34.8300 ;
      RECT 9.9280 33.7365 9.9540 34.8300 ;
      RECT 9.8200 33.7365 9.8460 34.8300 ;
      RECT 9.7120 33.7365 9.7380 34.8300 ;
      RECT 9.6040 33.7365 9.6300 34.8300 ;
      RECT 9.4960 33.7365 9.5220 34.8300 ;
      RECT 9.3880 33.7365 9.4140 34.8300 ;
      RECT 9.2800 33.7365 9.3060 34.8300 ;
      RECT 9.1720 33.7365 9.1980 34.8300 ;
      RECT 9.0640 33.7365 9.0900 34.8300 ;
      RECT 8.9560 33.7365 8.9820 34.8300 ;
      RECT 8.8480 33.7365 8.8740 34.8300 ;
      RECT 8.7400 33.7365 8.7660 34.8300 ;
      RECT 8.6320 33.7365 8.6580 34.8300 ;
      RECT 8.5240 33.7365 8.5500 34.8300 ;
      RECT 8.4160 33.7365 8.4420 34.8300 ;
      RECT 8.3080 33.7365 8.3340 34.8300 ;
      RECT 8.2000 33.7365 8.2260 34.8300 ;
      RECT 8.0920 33.7365 8.1180 34.8300 ;
      RECT 7.9840 33.7365 8.0100 34.8300 ;
      RECT 7.8760 33.7365 7.9020 34.8300 ;
      RECT 7.7680 33.7365 7.7940 34.8300 ;
      RECT 7.6600 33.7365 7.6860 34.8300 ;
      RECT 7.5520 33.7365 7.5780 34.8300 ;
      RECT 7.4440 33.7365 7.4700 34.8300 ;
      RECT 7.3360 33.7365 7.3620 34.8300 ;
      RECT 7.2280 33.7365 7.2540 34.8300 ;
      RECT 7.1200 33.7365 7.1460 34.8300 ;
      RECT 7.0120 33.7365 7.0380 34.8300 ;
      RECT 6.9040 33.7365 6.9300 34.8300 ;
      RECT 6.7960 33.7365 6.8220 34.8300 ;
      RECT 6.6880 33.7365 6.7140 34.8300 ;
      RECT 6.5800 33.7365 6.6060 34.8300 ;
      RECT 6.4720 33.7365 6.4980 34.8300 ;
      RECT 6.3640 33.7365 6.3900 34.8300 ;
      RECT 6.2560 33.7365 6.2820 34.8300 ;
      RECT 6.1480 33.7365 6.1740 34.8300 ;
      RECT 6.0400 33.7365 6.0660 34.8300 ;
      RECT 5.9320 33.7365 5.9580 34.8300 ;
      RECT 5.8240 33.7365 5.8500 34.8300 ;
      RECT 5.7160 33.7365 5.7420 34.8300 ;
      RECT 5.6080 33.7365 5.6340 34.8300 ;
      RECT 5.5000 33.7365 5.5260 34.8300 ;
      RECT 5.3920 33.7365 5.4180 34.8300 ;
      RECT 5.2840 33.7365 5.3100 34.8300 ;
      RECT 5.1760 33.7365 5.2020 34.8300 ;
      RECT 5.0680 33.7365 5.0940 34.8300 ;
      RECT 4.9600 33.7365 4.9860 34.8300 ;
      RECT 4.8520 33.7365 4.8780 34.8300 ;
      RECT 4.7440 33.7365 4.7700 34.8300 ;
      RECT 4.6360 33.7365 4.6620 34.8300 ;
      RECT 4.5280 33.7365 4.5540 34.8300 ;
      RECT 4.4200 33.7365 4.4460 34.8300 ;
      RECT 4.3120 33.7365 4.3380 34.8300 ;
      RECT 4.2040 33.7365 4.2300 34.8300 ;
      RECT 4.0960 33.7365 4.1220 34.8300 ;
      RECT 3.9880 33.7365 4.0140 34.8300 ;
      RECT 3.8800 33.7365 3.9060 34.8300 ;
      RECT 3.7720 33.7365 3.7980 34.8300 ;
      RECT 3.6640 33.7365 3.6900 34.8300 ;
      RECT 3.5560 33.7365 3.5820 34.8300 ;
      RECT 3.4480 33.7365 3.4740 34.8300 ;
      RECT 3.3400 33.7365 3.3660 34.8300 ;
      RECT 3.2320 33.7365 3.2580 34.8300 ;
      RECT 3.1240 33.7365 3.1500 34.8300 ;
      RECT 3.0160 33.7365 3.0420 34.8300 ;
      RECT 2.9080 33.7365 2.9340 34.8300 ;
      RECT 2.8000 33.7365 2.8260 34.8300 ;
      RECT 2.6920 33.7365 2.7180 34.8300 ;
      RECT 2.5840 33.7365 2.6100 34.8300 ;
      RECT 2.4760 33.7365 2.5020 34.8300 ;
      RECT 2.3680 33.7365 2.3940 34.8300 ;
      RECT 2.2600 33.7365 2.2860 34.8300 ;
      RECT 2.1520 33.7365 2.1780 34.8300 ;
      RECT 2.0440 33.7365 2.0700 34.8300 ;
      RECT 1.9360 33.7365 1.9620 34.8300 ;
      RECT 1.8280 33.7365 1.8540 34.8300 ;
      RECT 1.7200 33.7365 1.7460 34.8300 ;
      RECT 1.6120 33.7365 1.6380 34.8300 ;
      RECT 1.5040 33.7365 1.5300 34.8300 ;
      RECT 1.3960 33.7365 1.4220 34.8300 ;
      RECT 1.2880 33.7365 1.3140 34.8300 ;
      RECT 1.1800 33.7365 1.2060 34.8300 ;
      RECT 1.0720 33.7365 1.0980 34.8300 ;
      RECT 0.9640 33.7365 0.9900 34.8300 ;
      RECT 0.8560 33.7365 0.8820 34.8300 ;
      RECT 0.7480 33.7365 0.7740 34.8300 ;
      RECT 0.6400 33.7365 0.6660 34.8300 ;
      RECT 0.5320 33.7365 0.5580 34.8300 ;
      RECT 0.4240 33.7365 0.4500 34.8300 ;
      RECT 0.3160 33.7365 0.3420 34.8300 ;
      RECT 0.2080 33.7365 0.2340 34.8300 ;
      RECT 0.0050 33.7365 0.0900 34.8300 ;
      RECT 14.1350 43.0660 30.3480 43.5070 ;
      RECT 17.7530 34.8535 30.3480 43.5070 ;
      RECT 16.2950 36.3575 30.3480 43.5070 ;
      RECT 17.5370 36.1625 30.3480 43.5070 ;
      RECT 14.1350 42.7655 16.2130 43.5070 ;
      RECT 15.5570 36.2585 16.2130 43.5070 ;
      RECT 14.1350 36.4655 15.2590 43.5070 ;
      RECT 15.1970 34.8535 15.2590 43.5070 ;
      RECT 15.5430 41.4995 16.2130 42.6075 ;
      RECT 16.2810 38.6465 30.3480 42.2395 ;
      RECT 14.1350 41.7335 15.2730 41.9955 ;
      RECT 15.5430 38.9615 16.2130 41.2935 ;
      RECT 14.1350 39.3395 15.2730 40.6455 ;
      RECT 14.1350 36.6755 15.2730 39.2955 ;
      RECT 15.5430 36.1355 16.1590 37.9215 ;
      RECT 14.1890 36.4055 15.2730 36.5955 ;
      RECT 14.1890 35.6195 15.2590 43.5070 ;
      RECT 14.4050 35.5385 15.2590 43.5070 ;
      RECT 14.1890 36.1355 15.2730 36.3615 ;
      RECT 16.4570 36.1655 30.3480 43.5070 ;
      RECT 16.2950 34.8535 16.3750 43.5070 ;
      RECT 14.1350 35.5385 14.3230 36.3525 ;
      RECT 16.2950 34.8535 16.5910 36.2565 ;
      RECT 16.2950 35.9705 17.4550 36.2565 ;
      RECT 17.5370 34.8535 17.6710 43.5070 ;
      RECT 15.5570 35.9705 16.1590 43.5070 ;
      RECT 15.8810 34.8535 16.2130 36.1035 ;
      RECT 16.2950 35.9705 17.6710 36.0645 ;
      RECT 17.3210 34.8535 30.3480 36.0615 ;
      RECT 14.1350 35.9915 15.2730 36.0555 ;
      RECT 17.1050 35.5865 30.3480 36.0615 ;
      RECT 16.2950 35.6195 17.0230 36.2565 ;
      RECT 15.5570 35.6195 15.7990 43.5070 ;
      RECT 14.4050 35.5955 15.2730 35.8575 ;
      RECT 15.5930 34.8535 16.2130 35.7615 ;
      RECT 16.8890 34.8535 17.2390 35.7255 ;
      RECT 16.2950 35.5385 16.8070 36.2565 ;
      RECT 16.6730 34.8535 16.8070 43.5070 ;
      RECT 14.4050 34.8535 15.1150 43.5070 ;
      RECT 14.2250 34.8535 14.3230 43.5070 ;
      RECT 16.6730 34.8535 17.2390 35.4885 ;
      RECT 15.5570 34.8535 16.2130 35.4885 ;
      RECT 14.2250 34.8535 15.1150 35.4885 ;
      RECT 16.6730 34.8535 30.3480 35.4855 ;
      RECT 15.5430 35.3255 16.2130 35.4795 ;
      RECT 16.2950 34.8535 30.3480 35.2215 ;
      RECT 14.1350 34.8535 15.2590 35.2215 ;
      RECT 14.1350 34.8535 16.2130 35.0185 ;
      RECT 17.7570 34.6635 17.7750 43.5070 ;
      RECT 17.6490 34.6635 17.6670 43.5070 ;
      RECT 17.5410 34.6635 17.5590 43.5070 ;
      RECT 17.4330 34.6635 17.4510 43.5070 ;
      RECT 17.3250 34.6635 17.3430 43.5070 ;
      RECT 17.2170 34.6635 17.2350 43.5070 ;
      RECT 17.1090 34.6635 17.1270 43.5070 ;
      RECT 17.0010 34.6635 17.0190 43.5070 ;
      RECT 16.8930 34.6635 16.9110 43.5070 ;
      RECT 16.7850 34.6635 16.8030 43.5070 ;
      RECT 16.6770 34.6635 16.6950 43.5070 ;
      RECT 16.5690 34.6635 16.5870 43.5070 ;
      RECT 16.4610 34.6635 16.4790 43.5070 ;
      RECT 16.3530 34.6635 16.3710 43.5070 ;
      RECT 0.0000 36.1625 14.0170 43.5070 ;
      RECT 0.0000 38.9515 14.0310 39.0345 ;
      RECT 13.7570 34.8535 14.0530 38.6130 ;
      RECT 12.8930 35.7815 13.6750 43.5070 ;
      RECT 0.0000 34.8535 12.8110 43.5070 ;
      RECT 13.5410 34.8535 14.0530 36.0615 ;
      RECT 0.0000 35.5865 13.4590 36.0615 ;
      RECT 13.3250 34.8535 13.4590 43.5070 ;
      RECT 13.1090 35.5385 13.4590 43.5070 ;
      RECT 0.0000 34.8535 13.0270 36.0615 ;
      RECT 13.1090 34.8535 13.2430 43.5070 ;
      RECT 13.3250 34.8535 14.0530 35.4885 ;
      RECT 0.0000 34.8535 13.2430 35.4855 ;
      RECT 0.0000 34.8535 14.0530 35.2215 ;
      RECT 13.3290 34.8270 13.3470 43.5070 ;
      RECT 13.2210 34.8270 13.2390 43.5070 ;
        RECT 15.5530 42.9435 15.6810 44.0370 ;
        RECT 15.5390 43.6090 15.6810 43.9315 ;
        RECT 15.3190 43.3360 15.4530 44.0370 ;
        RECT 15.2960 43.6710 15.4530 43.9290 ;
        RECT 15.3190 42.9435 15.4170 44.0370 ;
        RECT 15.3190 43.0645 15.4310 43.3040 ;
        RECT 15.3190 42.9435 15.4530 43.0325 ;
        RECT 15.0940 43.3940 15.2280 44.0370 ;
        RECT 15.0940 42.9435 15.1920 44.0370 ;
        RECT 14.6770 42.9435 14.7600 44.0370 ;
        RECT 14.6770 43.0320 14.7740 43.9675 ;
        RECT 30.2680 42.9435 30.3530 44.0370 ;
        RECT 30.1240 42.9435 30.1500 44.0370 ;
        RECT 30.0160 42.9435 30.0420 44.0370 ;
        RECT 29.9080 42.9435 29.9340 44.0370 ;
        RECT 29.8000 42.9435 29.8260 44.0370 ;
        RECT 29.6920 42.9435 29.7180 44.0370 ;
        RECT 29.5840 42.9435 29.6100 44.0370 ;
        RECT 29.4760 42.9435 29.5020 44.0370 ;
        RECT 29.3680 42.9435 29.3940 44.0370 ;
        RECT 29.2600 42.9435 29.2860 44.0370 ;
        RECT 29.1520 42.9435 29.1780 44.0370 ;
        RECT 29.0440 42.9435 29.0700 44.0370 ;
        RECT 28.9360 42.9435 28.9620 44.0370 ;
        RECT 28.8280 42.9435 28.8540 44.0370 ;
        RECT 28.7200 42.9435 28.7460 44.0370 ;
        RECT 28.6120 42.9435 28.6380 44.0370 ;
        RECT 28.5040 42.9435 28.5300 44.0370 ;
        RECT 28.3960 42.9435 28.4220 44.0370 ;
        RECT 28.2880 42.9435 28.3140 44.0370 ;
        RECT 28.1800 42.9435 28.2060 44.0370 ;
        RECT 28.0720 42.9435 28.0980 44.0370 ;
        RECT 27.9640 42.9435 27.9900 44.0370 ;
        RECT 27.8560 42.9435 27.8820 44.0370 ;
        RECT 27.7480 42.9435 27.7740 44.0370 ;
        RECT 27.6400 42.9435 27.6660 44.0370 ;
        RECT 27.5320 42.9435 27.5580 44.0370 ;
        RECT 27.4240 42.9435 27.4500 44.0370 ;
        RECT 27.3160 42.9435 27.3420 44.0370 ;
        RECT 27.2080 42.9435 27.2340 44.0370 ;
        RECT 27.1000 42.9435 27.1260 44.0370 ;
        RECT 26.9920 42.9435 27.0180 44.0370 ;
        RECT 26.8840 42.9435 26.9100 44.0370 ;
        RECT 26.7760 42.9435 26.8020 44.0370 ;
        RECT 26.6680 42.9435 26.6940 44.0370 ;
        RECT 26.5600 42.9435 26.5860 44.0370 ;
        RECT 26.4520 42.9435 26.4780 44.0370 ;
        RECT 26.3440 42.9435 26.3700 44.0370 ;
        RECT 26.2360 42.9435 26.2620 44.0370 ;
        RECT 26.1280 42.9435 26.1540 44.0370 ;
        RECT 26.0200 42.9435 26.0460 44.0370 ;
        RECT 25.9120 42.9435 25.9380 44.0370 ;
        RECT 25.8040 42.9435 25.8300 44.0370 ;
        RECT 25.6960 42.9435 25.7220 44.0370 ;
        RECT 25.5880 42.9435 25.6140 44.0370 ;
        RECT 25.4800 42.9435 25.5060 44.0370 ;
        RECT 25.3720 42.9435 25.3980 44.0370 ;
        RECT 25.2640 42.9435 25.2900 44.0370 ;
        RECT 25.1560 42.9435 25.1820 44.0370 ;
        RECT 25.0480 42.9435 25.0740 44.0370 ;
        RECT 24.9400 42.9435 24.9660 44.0370 ;
        RECT 24.8320 42.9435 24.8580 44.0370 ;
        RECT 24.7240 42.9435 24.7500 44.0370 ;
        RECT 24.6160 42.9435 24.6420 44.0370 ;
        RECT 24.5080 42.9435 24.5340 44.0370 ;
        RECT 24.4000 42.9435 24.4260 44.0370 ;
        RECT 24.2920 42.9435 24.3180 44.0370 ;
        RECT 24.1840 42.9435 24.2100 44.0370 ;
        RECT 24.0760 42.9435 24.1020 44.0370 ;
        RECT 23.9680 42.9435 23.9940 44.0370 ;
        RECT 23.8600 42.9435 23.8860 44.0370 ;
        RECT 23.7520 42.9435 23.7780 44.0370 ;
        RECT 23.6440 42.9435 23.6700 44.0370 ;
        RECT 23.5360 42.9435 23.5620 44.0370 ;
        RECT 23.4280 42.9435 23.4540 44.0370 ;
        RECT 23.3200 42.9435 23.3460 44.0370 ;
        RECT 23.2120 42.9435 23.2380 44.0370 ;
        RECT 23.1040 42.9435 23.1300 44.0370 ;
        RECT 22.9960 42.9435 23.0220 44.0370 ;
        RECT 22.8880 42.9435 22.9140 44.0370 ;
        RECT 22.7800 42.9435 22.8060 44.0370 ;
        RECT 22.6720 42.9435 22.6980 44.0370 ;
        RECT 22.5640 42.9435 22.5900 44.0370 ;
        RECT 22.4560 42.9435 22.4820 44.0370 ;
        RECT 22.3480 42.9435 22.3740 44.0370 ;
        RECT 22.2400 42.9435 22.2660 44.0370 ;
        RECT 22.1320 42.9435 22.1580 44.0370 ;
        RECT 22.0240 42.9435 22.0500 44.0370 ;
        RECT 21.9160 42.9435 21.9420 44.0370 ;
        RECT 21.8080 42.9435 21.8340 44.0370 ;
        RECT 21.7000 42.9435 21.7260 44.0370 ;
        RECT 21.5920 42.9435 21.6180 44.0370 ;
        RECT 21.4840 42.9435 21.5100 44.0370 ;
        RECT 21.3760 42.9435 21.4020 44.0370 ;
        RECT 21.2680 42.9435 21.2940 44.0370 ;
        RECT 21.1600 42.9435 21.1860 44.0370 ;
        RECT 21.0520 42.9435 21.0780 44.0370 ;
        RECT 20.9440 42.9435 20.9700 44.0370 ;
        RECT 20.8360 42.9435 20.8620 44.0370 ;
        RECT 20.7280 42.9435 20.7540 44.0370 ;
        RECT 20.6200 42.9435 20.6460 44.0370 ;
        RECT 20.5120 42.9435 20.5380 44.0370 ;
        RECT 20.4040 42.9435 20.4300 44.0370 ;
        RECT 20.2960 42.9435 20.3220 44.0370 ;
        RECT 20.1880 42.9435 20.2140 44.0370 ;
        RECT 20.0800 42.9435 20.1060 44.0370 ;
        RECT 19.9720 42.9435 19.9980 44.0370 ;
        RECT 19.8640 42.9435 19.8900 44.0370 ;
        RECT 19.7560 42.9435 19.7820 44.0370 ;
        RECT 19.6480 42.9435 19.6740 44.0370 ;
        RECT 19.5400 42.9435 19.5660 44.0370 ;
        RECT 19.4320 42.9435 19.4580 44.0370 ;
        RECT 19.3240 42.9435 19.3500 44.0370 ;
        RECT 19.2160 42.9435 19.2420 44.0370 ;
        RECT 19.1080 42.9435 19.1340 44.0370 ;
        RECT 19.0000 42.9435 19.0260 44.0370 ;
        RECT 18.8920 42.9435 18.9180 44.0370 ;
        RECT 18.7840 42.9435 18.8100 44.0370 ;
        RECT 18.6760 42.9435 18.7020 44.0370 ;
        RECT 18.5680 42.9435 18.5940 44.0370 ;
        RECT 18.4600 42.9435 18.4860 44.0370 ;
        RECT 18.3520 42.9435 18.3780 44.0370 ;
        RECT 18.2440 42.9435 18.2700 44.0370 ;
        RECT 18.1360 42.9435 18.1620 44.0370 ;
        RECT 18.0280 42.9435 18.0540 44.0370 ;
        RECT 17.9200 42.9435 17.9460 44.0370 ;
        RECT 17.8120 42.9435 17.8380 44.0370 ;
        RECT 17.7040 42.9435 17.7300 44.0370 ;
        RECT 17.5960 42.9435 17.6220 44.0370 ;
        RECT 17.4880 42.9435 17.5140 44.0370 ;
        RECT 17.3800 42.9435 17.4060 44.0370 ;
        RECT 17.2720 42.9435 17.2980 44.0370 ;
        RECT 17.1640 42.9435 17.1900 44.0370 ;
        RECT 17.0560 42.9435 17.0820 44.0370 ;
        RECT 16.9480 42.9435 16.9740 44.0370 ;
        RECT 16.8400 42.9435 16.8660 44.0370 ;
        RECT 16.7320 42.9435 16.7580 44.0370 ;
        RECT 16.6240 42.9435 16.6500 44.0370 ;
        RECT 16.5160 42.9435 16.5420 44.0370 ;
        RECT 16.4080 42.9435 16.4340 44.0370 ;
        RECT 16.3000 42.9435 16.3260 44.0370 ;
        RECT 16.0870 42.9435 16.1640 44.0370 ;
        RECT 14.1940 42.9435 14.2710 44.0370 ;
        RECT 14.0320 42.9435 14.0580 44.0370 ;
        RECT 13.9240 42.9435 13.9500 44.0370 ;
        RECT 13.8160 42.9435 13.8420 44.0370 ;
        RECT 13.7080 42.9435 13.7340 44.0370 ;
        RECT 13.6000 42.9435 13.6260 44.0370 ;
        RECT 13.4920 42.9435 13.5180 44.0370 ;
        RECT 13.3840 42.9435 13.4100 44.0370 ;
        RECT 13.2760 42.9435 13.3020 44.0370 ;
        RECT 13.1680 42.9435 13.1940 44.0370 ;
        RECT 13.0600 42.9435 13.0860 44.0370 ;
        RECT 12.9520 42.9435 12.9780 44.0370 ;
        RECT 12.8440 42.9435 12.8700 44.0370 ;
        RECT 12.7360 42.9435 12.7620 44.0370 ;
        RECT 12.6280 42.9435 12.6540 44.0370 ;
        RECT 12.5200 42.9435 12.5460 44.0370 ;
        RECT 12.4120 42.9435 12.4380 44.0370 ;
        RECT 12.3040 42.9435 12.3300 44.0370 ;
        RECT 12.1960 42.9435 12.2220 44.0370 ;
        RECT 12.0880 42.9435 12.1140 44.0370 ;
        RECT 11.9800 42.9435 12.0060 44.0370 ;
        RECT 11.8720 42.9435 11.8980 44.0370 ;
        RECT 11.7640 42.9435 11.7900 44.0370 ;
        RECT 11.6560 42.9435 11.6820 44.0370 ;
        RECT 11.5480 42.9435 11.5740 44.0370 ;
        RECT 11.4400 42.9435 11.4660 44.0370 ;
        RECT 11.3320 42.9435 11.3580 44.0370 ;
        RECT 11.2240 42.9435 11.2500 44.0370 ;
        RECT 11.1160 42.9435 11.1420 44.0370 ;
        RECT 11.0080 42.9435 11.0340 44.0370 ;
        RECT 10.9000 42.9435 10.9260 44.0370 ;
        RECT 10.7920 42.9435 10.8180 44.0370 ;
        RECT 10.6840 42.9435 10.7100 44.0370 ;
        RECT 10.5760 42.9435 10.6020 44.0370 ;
        RECT 10.4680 42.9435 10.4940 44.0370 ;
        RECT 10.3600 42.9435 10.3860 44.0370 ;
        RECT 10.2520 42.9435 10.2780 44.0370 ;
        RECT 10.1440 42.9435 10.1700 44.0370 ;
        RECT 10.0360 42.9435 10.0620 44.0370 ;
        RECT 9.9280 42.9435 9.9540 44.0370 ;
        RECT 9.8200 42.9435 9.8460 44.0370 ;
        RECT 9.7120 42.9435 9.7380 44.0370 ;
        RECT 9.6040 42.9435 9.6300 44.0370 ;
        RECT 9.4960 42.9435 9.5220 44.0370 ;
        RECT 9.3880 42.9435 9.4140 44.0370 ;
        RECT 9.2800 42.9435 9.3060 44.0370 ;
        RECT 9.1720 42.9435 9.1980 44.0370 ;
        RECT 9.0640 42.9435 9.0900 44.0370 ;
        RECT 8.9560 42.9435 8.9820 44.0370 ;
        RECT 8.8480 42.9435 8.8740 44.0370 ;
        RECT 8.7400 42.9435 8.7660 44.0370 ;
        RECT 8.6320 42.9435 8.6580 44.0370 ;
        RECT 8.5240 42.9435 8.5500 44.0370 ;
        RECT 8.4160 42.9435 8.4420 44.0370 ;
        RECT 8.3080 42.9435 8.3340 44.0370 ;
        RECT 8.2000 42.9435 8.2260 44.0370 ;
        RECT 8.0920 42.9435 8.1180 44.0370 ;
        RECT 7.9840 42.9435 8.0100 44.0370 ;
        RECT 7.8760 42.9435 7.9020 44.0370 ;
        RECT 7.7680 42.9435 7.7940 44.0370 ;
        RECT 7.6600 42.9435 7.6860 44.0370 ;
        RECT 7.5520 42.9435 7.5780 44.0370 ;
        RECT 7.4440 42.9435 7.4700 44.0370 ;
        RECT 7.3360 42.9435 7.3620 44.0370 ;
        RECT 7.2280 42.9435 7.2540 44.0370 ;
        RECT 7.1200 42.9435 7.1460 44.0370 ;
        RECT 7.0120 42.9435 7.0380 44.0370 ;
        RECT 6.9040 42.9435 6.9300 44.0370 ;
        RECT 6.7960 42.9435 6.8220 44.0370 ;
        RECT 6.6880 42.9435 6.7140 44.0370 ;
        RECT 6.5800 42.9435 6.6060 44.0370 ;
        RECT 6.4720 42.9435 6.4980 44.0370 ;
        RECT 6.3640 42.9435 6.3900 44.0370 ;
        RECT 6.2560 42.9435 6.2820 44.0370 ;
        RECT 6.1480 42.9435 6.1740 44.0370 ;
        RECT 6.0400 42.9435 6.0660 44.0370 ;
        RECT 5.9320 42.9435 5.9580 44.0370 ;
        RECT 5.8240 42.9435 5.8500 44.0370 ;
        RECT 5.7160 42.9435 5.7420 44.0370 ;
        RECT 5.6080 42.9435 5.6340 44.0370 ;
        RECT 5.5000 42.9435 5.5260 44.0370 ;
        RECT 5.3920 42.9435 5.4180 44.0370 ;
        RECT 5.2840 42.9435 5.3100 44.0370 ;
        RECT 5.1760 42.9435 5.2020 44.0370 ;
        RECT 5.0680 42.9435 5.0940 44.0370 ;
        RECT 4.9600 42.9435 4.9860 44.0370 ;
        RECT 4.8520 42.9435 4.8780 44.0370 ;
        RECT 4.7440 42.9435 4.7700 44.0370 ;
        RECT 4.6360 42.9435 4.6620 44.0370 ;
        RECT 4.5280 42.9435 4.5540 44.0370 ;
        RECT 4.4200 42.9435 4.4460 44.0370 ;
        RECT 4.3120 42.9435 4.3380 44.0370 ;
        RECT 4.2040 42.9435 4.2300 44.0370 ;
        RECT 4.0960 42.9435 4.1220 44.0370 ;
        RECT 3.9880 42.9435 4.0140 44.0370 ;
        RECT 3.8800 42.9435 3.9060 44.0370 ;
        RECT 3.7720 42.9435 3.7980 44.0370 ;
        RECT 3.6640 42.9435 3.6900 44.0370 ;
        RECT 3.5560 42.9435 3.5820 44.0370 ;
        RECT 3.4480 42.9435 3.4740 44.0370 ;
        RECT 3.3400 42.9435 3.3660 44.0370 ;
        RECT 3.2320 42.9435 3.2580 44.0370 ;
        RECT 3.1240 42.9435 3.1500 44.0370 ;
        RECT 3.0160 42.9435 3.0420 44.0370 ;
        RECT 2.9080 42.9435 2.9340 44.0370 ;
        RECT 2.8000 42.9435 2.8260 44.0370 ;
        RECT 2.6920 42.9435 2.7180 44.0370 ;
        RECT 2.5840 42.9435 2.6100 44.0370 ;
        RECT 2.4760 42.9435 2.5020 44.0370 ;
        RECT 2.3680 42.9435 2.3940 44.0370 ;
        RECT 2.2600 42.9435 2.2860 44.0370 ;
        RECT 2.1520 42.9435 2.1780 44.0370 ;
        RECT 2.0440 42.9435 2.0700 44.0370 ;
        RECT 1.9360 42.9435 1.9620 44.0370 ;
        RECT 1.8280 42.9435 1.8540 44.0370 ;
        RECT 1.7200 42.9435 1.7460 44.0370 ;
        RECT 1.6120 42.9435 1.6380 44.0370 ;
        RECT 1.5040 42.9435 1.5300 44.0370 ;
        RECT 1.3960 42.9435 1.4220 44.0370 ;
        RECT 1.2880 42.9435 1.3140 44.0370 ;
        RECT 1.1800 42.9435 1.2060 44.0370 ;
        RECT 1.0720 42.9435 1.0980 44.0370 ;
        RECT 0.9640 42.9435 0.9900 44.0370 ;
        RECT 0.8560 42.9435 0.8820 44.0370 ;
        RECT 0.7480 42.9435 0.7740 44.0370 ;
        RECT 0.6400 42.9435 0.6660 44.0370 ;
        RECT 0.5320 42.9435 0.5580 44.0370 ;
        RECT 0.4240 42.9435 0.4500 44.0370 ;
        RECT 0.3160 42.9435 0.3420 44.0370 ;
        RECT 0.2080 42.9435 0.2340 44.0370 ;
        RECT 0.0050 42.9435 0.0900 44.0370 ;
        RECT 15.5530 44.0235 15.6810 45.1170 ;
        RECT 15.5390 44.6890 15.6810 45.0115 ;
        RECT 15.3190 44.4160 15.4530 45.1170 ;
        RECT 15.2960 44.7510 15.4530 45.0090 ;
        RECT 15.3190 44.0235 15.4170 45.1170 ;
        RECT 15.3190 44.1445 15.4310 44.3840 ;
        RECT 15.3190 44.0235 15.4530 44.1125 ;
        RECT 15.0940 44.4740 15.2280 45.1170 ;
        RECT 15.0940 44.0235 15.1920 45.1170 ;
        RECT 14.6770 44.0235 14.7600 45.1170 ;
        RECT 14.6770 44.1120 14.7740 45.0475 ;
        RECT 30.2680 44.0235 30.3530 45.1170 ;
        RECT 30.1240 44.0235 30.1500 45.1170 ;
        RECT 30.0160 44.0235 30.0420 45.1170 ;
        RECT 29.9080 44.0235 29.9340 45.1170 ;
        RECT 29.8000 44.0235 29.8260 45.1170 ;
        RECT 29.6920 44.0235 29.7180 45.1170 ;
        RECT 29.5840 44.0235 29.6100 45.1170 ;
        RECT 29.4760 44.0235 29.5020 45.1170 ;
        RECT 29.3680 44.0235 29.3940 45.1170 ;
        RECT 29.2600 44.0235 29.2860 45.1170 ;
        RECT 29.1520 44.0235 29.1780 45.1170 ;
        RECT 29.0440 44.0235 29.0700 45.1170 ;
        RECT 28.9360 44.0235 28.9620 45.1170 ;
        RECT 28.8280 44.0235 28.8540 45.1170 ;
        RECT 28.7200 44.0235 28.7460 45.1170 ;
        RECT 28.6120 44.0235 28.6380 45.1170 ;
        RECT 28.5040 44.0235 28.5300 45.1170 ;
        RECT 28.3960 44.0235 28.4220 45.1170 ;
        RECT 28.2880 44.0235 28.3140 45.1170 ;
        RECT 28.1800 44.0235 28.2060 45.1170 ;
        RECT 28.0720 44.0235 28.0980 45.1170 ;
        RECT 27.9640 44.0235 27.9900 45.1170 ;
        RECT 27.8560 44.0235 27.8820 45.1170 ;
        RECT 27.7480 44.0235 27.7740 45.1170 ;
        RECT 27.6400 44.0235 27.6660 45.1170 ;
        RECT 27.5320 44.0235 27.5580 45.1170 ;
        RECT 27.4240 44.0235 27.4500 45.1170 ;
        RECT 27.3160 44.0235 27.3420 45.1170 ;
        RECT 27.2080 44.0235 27.2340 45.1170 ;
        RECT 27.1000 44.0235 27.1260 45.1170 ;
        RECT 26.9920 44.0235 27.0180 45.1170 ;
        RECT 26.8840 44.0235 26.9100 45.1170 ;
        RECT 26.7760 44.0235 26.8020 45.1170 ;
        RECT 26.6680 44.0235 26.6940 45.1170 ;
        RECT 26.5600 44.0235 26.5860 45.1170 ;
        RECT 26.4520 44.0235 26.4780 45.1170 ;
        RECT 26.3440 44.0235 26.3700 45.1170 ;
        RECT 26.2360 44.0235 26.2620 45.1170 ;
        RECT 26.1280 44.0235 26.1540 45.1170 ;
        RECT 26.0200 44.0235 26.0460 45.1170 ;
        RECT 25.9120 44.0235 25.9380 45.1170 ;
        RECT 25.8040 44.0235 25.8300 45.1170 ;
        RECT 25.6960 44.0235 25.7220 45.1170 ;
        RECT 25.5880 44.0235 25.6140 45.1170 ;
        RECT 25.4800 44.0235 25.5060 45.1170 ;
        RECT 25.3720 44.0235 25.3980 45.1170 ;
        RECT 25.2640 44.0235 25.2900 45.1170 ;
        RECT 25.1560 44.0235 25.1820 45.1170 ;
        RECT 25.0480 44.0235 25.0740 45.1170 ;
        RECT 24.9400 44.0235 24.9660 45.1170 ;
        RECT 24.8320 44.0235 24.8580 45.1170 ;
        RECT 24.7240 44.0235 24.7500 45.1170 ;
        RECT 24.6160 44.0235 24.6420 45.1170 ;
        RECT 24.5080 44.0235 24.5340 45.1170 ;
        RECT 24.4000 44.0235 24.4260 45.1170 ;
        RECT 24.2920 44.0235 24.3180 45.1170 ;
        RECT 24.1840 44.0235 24.2100 45.1170 ;
        RECT 24.0760 44.0235 24.1020 45.1170 ;
        RECT 23.9680 44.0235 23.9940 45.1170 ;
        RECT 23.8600 44.0235 23.8860 45.1170 ;
        RECT 23.7520 44.0235 23.7780 45.1170 ;
        RECT 23.6440 44.0235 23.6700 45.1170 ;
        RECT 23.5360 44.0235 23.5620 45.1170 ;
        RECT 23.4280 44.0235 23.4540 45.1170 ;
        RECT 23.3200 44.0235 23.3460 45.1170 ;
        RECT 23.2120 44.0235 23.2380 45.1170 ;
        RECT 23.1040 44.0235 23.1300 45.1170 ;
        RECT 22.9960 44.0235 23.0220 45.1170 ;
        RECT 22.8880 44.0235 22.9140 45.1170 ;
        RECT 22.7800 44.0235 22.8060 45.1170 ;
        RECT 22.6720 44.0235 22.6980 45.1170 ;
        RECT 22.5640 44.0235 22.5900 45.1170 ;
        RECT 22.4560 44.0235 22.4820 45.1170 ;
        RECT 22.3480 44.0235 22.3740 45.1170 ;
        RECT 22.2400 44.0235 22.2660 45.1170 ;
        RECT 22.1320 44.0235 22.1580 45.1170 ;
        RECT 22.0240 44.0235 22.0500 45.1170 ;
        RECT 21.9160 44.0235 21.9420 45.1170 ;
        RECT 21.8080 44.0235 21.8340 45.1170 ;
        RECT 21.7000 44.0235 21.7260 45.1170 ;
        RECT 21.5920 44.0235 21.6180 45.1170 ;
        RECT 21.4840 44.0235 21.5100 45.1170 ;
        RECT 21.3760 44.0235 21.4020 45.1170 ;
        RECT 21.2680 44.0235 21.2940 45.1170 ;
        RECT 21.1600 44.0235 21.1860 45.1170 ;
        RECT 21.0520 44.0235 21.0780 45.1170 ;
        RECT 20.9440 44.0235 20.9700 45.1170 ;
        RECT 20.8360 44.0235 20.8620 45.1170 ;
        RECT 20.7280 44.0235 20.7540 45.1170 ;
        RECT 20.6200 44.0235 20.6460 45.1170 ;
        RECT 20.5120 44.0235 20.5380 45.1170 ;
        RECT 20.4040 44.0235 20.4300 45.1170 ;
        RECT 20.2960 44.0235 20.3220 45.1170 ;
        RECT 20.1880 44.0235 20.2140 45.1170 ;
        RECT 20.0800 44.0235 20.1060 45.1170 ;
        RECT 19.9720 44.0235 19.9980 45.1170 ;
        RECT 19.8640 44.0235 19.8900 45.1170 ;
        RECT 19.7560 44.0235 19.7820 45.1170 ;
        RECT 19.6480 44.0235 19.6740 45.1170 ;
        RECT 19.5400 44.0235 19.5660 45.1170 ;
        RECT 19.4320 44.0235 19.4580 45.1170 ;
        RECT 19.3240 44.0235 19.3500 45.1170 ;
        RECT 19.2160 44.0235 19.2420 45.1170 ;
        RECT 19.1080 44.0235 19.1340 45.1170 ;
        RECT 19.0000 44.0235 19.0260 45.1170 ;
        RECT 18.8920 44.0235 18.9180 45.1170 ;
        RECT 18.7840 44.0235 18.8100 45.1170 ;
        RECT 18.6760 44.0235 18.7020 45.1170 ;
        RECT 18.5680 44.0235 18.5940 45.1170 ;
        RECT 18.4600 44.0235 18.4860 45.1170 ;
        RECT 18.3520 44.0235 18.3780 45.1170 ;
        RECT 18.2440 44.0235 18.2700 45.1170 ;
        RECT 18.1360 44.0235 18.1620 45.1170 ;
        RECT 18.0280 44.0235 18.0540 45.1170 ;
        RECT 17.9200 44.0235 17.9460 45.1170 ;
        RECT 17.8120 44.0235 17.8380 45.1170 ;
        RECT 17.7040 44.0235 17.7300 45.1170 ;
        RECT 17.5960 44.0235 17.6220 45.1170 ;
        RECT 17.4880 44.0235 17.5140 45.1170 ;
        RECT 17.3800 44.0235 17.4060 45.1170 ;
        RECT 17.2720 44.0235 17.2980 45.1170 ;
        RECT 17.1640 44.0235 17.1900 45.1170 ;
        RECT 17.0560 44.0235 17.0820 45.1170 ;
        RECT 16.9480 44.0235 16.9740 45.1170 ;
        RECT 16.8400 44.0235 16.8660 45.1170 ;
        RECT 16.7320 44.0235 16.7580 45.1170 ;
        RECT 16.6240 44.0235 16.6500 45.1170 ;
        RECT 16.5160 44.0235 16.5420 45.1170 ;
        RECT 16.4080 44.0235 16.4340 45.1170 ;
        RECT 16.3000 44.0235 16.3260 45.1170 ;
        RECT 16.0870 44.0235 16.1640 45.1170 ;
        RECT 14.1940 44.0235 14.2710 45.1170 ;
        RECT 14.0320 44.0235 14.0580 45.1170 ;
        RECT 13.9240 44.0235 13.9500 45.1170 ;
        RECT 13.8160 44.0235 13.8420 45.1170 ;
        RECT 13.7080 44.0235 13.7340 45.1170 ;
        RECT 13.6000 44.0235 13.6260 45.1170 ;
        RECT 13.4920 44.0235 13.5180 45.1170 ;
        RECT 13.3840 44.0235 13.4100 45.1170 ;
        RECT 13.2760 44.0235 13.3020 45.1170 ;
        RECT 13.1680 44.0235 13.1940 45.1170 ;
        RECT 13.0600 44.0235 13.0860 45.1170 ;
        RECT 12.9520 44.0235 12.9780 45.1170 ;
        RECT 12.8440 44.0235 12.8700 45.1170 ;
        RECT 12.7360 44.0235 12.7620 45.1170 ;
        RECT 12.6280 44.0235 12.6540 45.1170 ;
        RECT 12.5200 44.0235 12.5460 45.1170 ;
        RECT 12.4120 44.0235 12.4380 45.1170 ;
        RECT 12.3040 44.0235 12.3300 45.1170 ;
        RECT 12.1960 44.0235 12.2220 45.1170 ;
        RECT 12.0880 44.0235 12.1140 45.1170 ;
        RECT 11.9800 44.0235 12.0060 45.1170 ;
        RECT 11.8720 44.0235 11.8980 45.1170 ;
        RECT 11.7640 44.0235 11.7900 45.1170 ;
        RECT 11.6560 44.0235 11.6820 45.1170 ;
        RECT 11.5480 44.0235 11.5740 45.1170 ;
        RECT 11.4400 44.0235 11.4660 45.1170 ;
        RECT 11.3320 44.0235 11.3580 45.1170 ;
        RECT 11.2240 44.0235 11.2500 45.1170 ;
        RECT 11.1160 44.0235 11.1420 45.1170 ;
        RECT 11.0080 44.0235 11.0340 45.1170 ;
        RECT 10.9000 44.0235 10.9260 45.1170 ;
        RECT 10.7920 44.0235 10.8180 45.1170 ;
        RECT 10.6840 44.0235 10.7100 45.1170 ;
        RECT 10.5760 44.0235 10.6020 45.1170 ;
        RECT 10.4680 44.0235 10.4940 45.1170 ;
        RECT 10.3600 44.0235 10.3860 45.1170 ;
        RECT 10.2520 44.0235 10.2780 45.1170 ;
        RECT 10.1440 44.0235 10.1700 45.1170 ;
        RECT 10.0360 44.0235 10.0620 45.1170 ;
        RECT 9.9280 44.0235 9.9540 45.1170 ;
        RECT 9.8200 44.0235 9.8460 45.1170 ;
        RECT 9.7120 44.0235 9.7380 45.1170 ;
        RECT 9.6040 44.0235 9.6300 45.1170 ;
        RECT 9.4960 44.0235 9.5220 45.1170 ;
        RECT 9.3880 44.0235 9.4140 45.1170 ;
        RECT 9.2800 44.0235 9.3060 45.1170 ;
        RECT 9.1720 44.0235 9.1980 45.1170 ;
        RECT 9.0640 44.0235 9.0900 45.1170 ;
        RECT 8.9560 44.0235 8.9820 45.1170 ;
        RECT 8.8480 44.0235 8.8740 45.1170 ;
        RECT 8.7400 44.0235 8.7660 45.1170 ;
        RECT 8.6320 44.0235 8.6580 45.1170 ;
        RECT 8.5240 44.0235 8.5500 45.1170 ;
        RECT 8.4160 44.0235 8.4420 45.1170 ;
        RECT 8.3080 44.0235 8.3340 45.1170 ;
        RECT 8.2000 44.0235 8.2260 45.1170 ;
        RECT 8.0920 44.0235 8.1180 45.1170 ;
        RECT 7.9840 44.0235 8.0100 45.1170 ;
        RECT 7.8760 44.0235 7.9020 45.1170 ;
        RECT 7.7680 44.0235 7.7940 45.1170 ;
        RECT 7.6600 44.0235 7.6860 45.1170 ;
        RECT 7.5520 44.0235 7.5780 45.1170 ;
        RECT 7.4440 44.0235 7.4700 45.1170 ;
        RECT 7.3360 44.0235 7.3620 45.1170 ;
        RECT 7.2280 44.0235 7.2540 45.1170 ;
        RECT 7.1200 44.0235 7.1460 45.1170 ;
        RECT 7.0120 44.0235 7.0380 45.1170 ;
        RECT 6.9040 44.0235 6.9300 45.1170 ;
        RECT 6.7960 44.0235 6.8220 45.1170 ;
        RECT 6.6880 44.0235 6.7140 45.1170 ;
        RECT 6.5800 44.0235 6.6060 45.1170 ;
        RECT 6.4720 44.0235 6.4980 45.1170 ;
        RECT 6.3640 44.0235 6.3900 45.1170 ;
        RECT 6.2560 44.0235 6.2820 45.1170 ;
        RECT 6.1480 44.0235 6.1740 45.1170 ;
        RECT 6.0400 44.0235 6.0660 45.1170 ;
        RECT 5.9320 44.0235 5.9580 45.1170 ;
        RECT 5.8240 44.0235 5.8500 45.1170 ;
        RECT 5.7160 44.0235 5.7420 45.1170 ;
        RECT 5.6080 44.0235 5.6340 45.1170 ;
        RECT 5.5000 44.0235 5.5260 45.1170 ;
        RECT 5.3920 44.0235 5.4180 45.1170 ;
        RECT 5.2840 44.0235 5.3100 45.1170 ;
        RECT 5.1760 44.0235 5.2020 45.1170 ;
        RECT 5.0680 44.0235 5.0940 45.1170 ;
        RECT 4.9600 44.0235 4.9860 45.1170 ;
        RECT 4.8520 44.0235 4.8780 45.1170 ;
        RECT 4.7440 44.0235 4.7700 45.1170 ;
        RECT 4.6360 44.0235 4.6620 45.1170 ;
        RECT 4.5280 44.0235 4.5540 45.1170 ;
        RECT 4.4200 44.0235 4.4460 45.1170 ;
        RECT 4.3120 44.0235 4.3380 45.1170 ;
        RECT 4.2040 44.0235 4.2300 45.1170 ;
        RECT 4.0960 44.0235 4.1220 45.1170 ;
        RECT 3.9880 44.0235 4.0140 45.1170 ;
        RECT 3.8800 44.0235 3.9060 45.1170 ;
        RECT 3.7720 44.0235 3.7980 45.1170 ;
        RECT 3.6640 44.0235 3.6900 45.1170 ;
        RECT 3.5560 44.0235 3.5820 45.1170 ;
        RECT 3.4480 44.0235 3.4740 45.1170 ;
        RECT 3.3400 44.0235 3.3660 45.1170 ;
        RECT 3.2320 44.0235 3.2580 45.1170 ;
        RECT 3.1240 44.0235 3.1500 45.1170 ;
        RECT 3.0160 44.0235 3.0420 45.1170 ;
        RECT 2.9080 44.0235 2.9340 45.1170 ;
        RECT 2.8000 44.0235 2.8260 45.1170 ;
        RECT 2.6920 44.0235 2.7180 45.1170 ;
        RECT 2.5840 44.0235 2.6100 45.1170 ;
        RECT 2.4760 44.0235 2.5020 45.1170 ;
        RECT 2.3680 44.0235 2.3940 45.1170 ;
        RECT 2.2600 44.0235 2.2860 45.1170 ;
        RECT 2.1520 44.0235 2.1780 45.1170 ;
        RECT 2.0440 44.0235 2.0700 45.1170 ;
        RECT 1.9360 44.0235 1.9620 45.1170 ;
        RECT 1.8280 44.0235 1.8540 45.1170 ;
        RECT 1.7200 44.0235 1.7460 45.1170 ;
        RECT 1.6120 44.0235 1.6380 45.1170 ;
        RECT 1.5040 44.0235 1.5300 45.1170 ;
        RECT 1.3960 44.0235 1.4220 45.1170 ;
        RECT 1.2880 44.0235 1.3140 45.1170 ;
        RECT 1.1800 44.0235 1.2060 45.1170 ;
        RECT 1.0720 44.0235 1.0980 45.1170 ;
        RECT 0.9640 44.0235 0.9900 45.1170 ;
        RECT 0.8560 44.0235 0.8820 45.1170 ;
        RECT 0.7480 44.0235 0.7740 45.1170 ;
        RECT 0.6400 44.0235 0.6660 45.1170 ;
        RECT 0.5320 44.0235 0.5580 45.1170 ;
        RECT 0.4240 44.0235 0.4500 45.1170 ;
        RECT 0.3160 44.0235 0.3420 45.1170 ;
        RECT 0.2080 44.0235 0.2340 45.1170 ;
        RECT 0.0050 44.0235 0.0900 45.1170 ;
        RECT 15.5530 45.1035 15.6810 46.1970 ;
        RECT 15.5390 45.7690 15.6810 46.0915 ;
        RECT 15.3190 45.4960 15.4530 46.1970 ;
        RECT 15.2960 45.8310 15.4530 46.0890 ;
        RECT 15.3190 45.1035 15.4170 46.1970 ;
        RECT 15.3190 45.2245 15.4310 45.4640 ;
        RECT 15.3190 45.1035 15.4530 45.1925 ;
        RECT 15.0940 45.5540 15.2280 46.1970 ;
        RECT 15.0940 45.1035 15.1920 46.1970 ;
        RECT 14.6770 45.1035 14.7600 46.1970 ;
        RECT 14.6770 45.1920 14.7740 46.1275 ;
        RECT 30.2680 45.1035 30.3530 46.1970 ;
        RECT 30.1240 45.1035 30.1500 46.1970 ;
        RECT 30.0160 45.1035 30.0420 46.1970 ;
        RECT 29.9080 45.1035 29.9340 46.1970 ;
        RECT 29.8000 45.1035 29.8260 46.1970 ;
        RECT 29.6920 45.1035 29.7180 46.1970 ;
        RECT 29.5840 45.1035 29.6100 46.1970 ;
        RECT 29.4760 45.1035 29.5020 46.1970 ;
        RECT 29.3680 45.1035 29.3940 46.1970 ;
        RECT 29.2600 45.1035 29.2860 46.1970 ;
        RECT 29.1520 45.1035 29.1780 46.1970 ;
        RECT 29.0440 45.1035 29.0700 46.1970 ;
        RECT 28.9360 45.1035 28.9620 46.1970 ;
        RECT 28.8280 45.1035 28.8540 46.1970 ;
        RECT 28.7200 45.1035 28.7460 46.1970 ;
        RECT 28.6120 45.1035 28.6380 46.1970 ;
        RECT 28.5040 45.1035 28.5300 46.1970 ;
        RECT 28.3960 45.1035 28.4220 46.1970 ;
        RECT 28.2880 45.1035 28.3140 46.1970 ;
        RECT 28.1800 45.1035 28.2060 46.1970 ;
        RECT 28.0720 45.1035 28.0980 46.1970 ;
        RECT 27.9640 45.1035 27.9900 46.1970 ;
        RECT 27.8560 45.1035 27.8820 46.1970 ;
        RECT 27.7480 45.1035 27.7740 46.1970 ;
        RECT 27.6400 45.1035 27.6660 46.1970 ;
        RECT 27.5320 45.1035 27.5580 46.1970 ;
        RECT 27.4240 45.1035 27.4500 46.1970 ;
        RECT 27.3160 45.1035 27.3420 46.1970 ;
        RECT 27.2080 45.1035 27.2340 46.1970 ;
        RECT 27.1000 45.1035 27.1260 46.1970 ;
        RECT 26.9920 45.1035 27.0180 46.1970 ;
        RECT 26.8840 45.1035 26.9100 46.1970 ;
        RECT 26.7760 45.1035 26.8020 46.1970 ;
        RECT 26.6680 45.1035 26.6940 46.1970 ;
        RECT 26.5600 45.1035 26.5860 46.1970 ;
        RECT 26.4520 45.1035 26.4780 46.1970 ;
        RECT 26.3440 45.1035 26.3700 46.1970 ;
        RECT 26.2360 45.1035 26.2620 46.1970 ;
        RECT 26.1280 45.1035 26.1540 46.1970 ;
        RECT 26.0200 45.1035 26.0460 46.1970 ;
        RECT 25.9120 45.1035 25.9380 46.1970 ;
        RECT 25.8040 45.1035 25.8300 46.1970 ;
        RECT 25.6960 45.1035 25.7220 46.1970 ;
        RECT 25.5880 45.1035 25.6140 46.1970 ;
        RECT 25.4800 45.1035 25.5060 46.1970 ;
        RECT 25.3720 45.1035 25.3980 46.1970 ;
        RECT 25.2640 45.1035 25.2900 46.1970 ;
        RECT 25.1560 45.1035 25.1820 46.1970 ;
        RECT 25.0480 45.1035 25.0740 46.1970 ;
        RECT 24.9400 45.1035 24.9660 46.1970 ;
        RECT 24.8320 45.1035 24.8580 46.1970 ;
        RECT 24.7240 45.1035 24.7500 46.1970 ;
        RECT 24.6160 45.1035 24.6420 46.1970 ;
        RECT 24.5080 45.1035 24.5340 46.1970 ;
        RECT 24.4000 45.1035 24.4260 46.1970 ;
        RECT 24.2920 45.1035 24.3180 46.1970 ;
        RECT 24.1840 45.1035 24.2100 46.1970 ;
        RECT 24.0760 45.1035 24.1020 46.1970 ;
        RECT 23.9680 45.1035 23.9940 46.1970 ;
        RECT 23.8600 45.1035 23.8860 46.1970 ;
        RECT 23.7520 45.1035 23.7780 46.1970 ;
        RECT 23.6440 45.1035 23.6700 46.1970 ;
        RECT 23.5360 45.1035 23.5620 46.1970 ;
        RECT 23.4280 45.1035 23.4540 46.1970 ;
        RECT 23.3200 45.1035 23.3460 46.1970 ;
        RECT 23.2120 45.1035 23.2380 46.1970 ;
        RECT 23.1040 45.1035 23.1300 46.1970 ;
        RECT 22.9960 45.1035 23.0220 46.1970 ;
        RECT 22.8880 45.1035 22.9140 46.1970 ;
        RECT 22.7800 45.1035 22.8060 46.1970 ;
        RECT 22.6720 45.1035 22.6980 46.1970 ;
        RECT 22.5640 45.1035 22.5900 46.1970 ;
        RECT 22.4560 45.1035 22.4820 46.1970 ;
        RECT 22.3480 45.1035 22.3740 46.1970 ;
        RECT 22.2400 45.1035 22.2660 46.1970 ;
        RECT 22.1320 45.1035 22.1580 46.1970 ;
        RECT 22.0240 45.1035 22.0500 46.1970 ;
        RECT 21.9160 45.1035 21.9420 46.1970 ;
        RECT 21.8080 45.1035 21.8340 46.1970 ;
        RECT 21.7000 45.1035 21.7260 46.1970 ;
        RECT 21.5920 45.1035 21.6180 46.1970 ;
        RECT 21.4840 45.1035 21.5100 46.1970 ;
        RECT 21.3760 45.1035 21.4020 46.1970 ;
        RECT 21.2680 45.1035 21.2940 46.1970 ;
        RECT 21.1600 45.1035 21.1860 46.1970 ;
        RECT 21.0520 45.1035 21.0780 46.1970 ;
        RECT 20.9440 45.1035 20.9700 46.1970 ;
        RECT 20.8360 45.1035 20.8620 46.1970 ;
        RECT 20.7280 45.1035 20.7540 46.1970 ;
        RECT 20.6200 45.1035 20.6460 46.1970 ;
        RECT 20.5120 45.1035 20.5380 46.1970 ;
        RECT 20.4040 45.1035 20.4300 46.1970 ;
        RECT 20.2960 45.1035 20.3220 46.1970 ;
        RECT 20.1880 45.1035 20.2140 46.1970 ;
        RECT 20.0800 45.1035 20.1060 46.1970 ;
        RECT 19.9720 45.1035 19.9980 46.1970 ;
        RECT 19.8640 45.1035 19.8900 46.1970 ;
        RECT 19.7560 45.1035 19.7820 46.1970 ;
        RECT 19.6480 45.1035 19.6740 46.1970 ;
        RECT 19.5400 45.1035 19.5660 46.1970 ;
        RECT 19.4320 45.1035 19.4580 46.1970 ;
        RECT 19.3240 45.1035 19.3500 46.1970 ;
        RECT 19.2160 45.1035 19.2420 46.1970 ;
        RECT 19.1080 45.1035 19.1340 46.1970 ;
        RECT 19.0000 45.1035 19.0260 46.1970 ;
        RECT 18.8920 45.1035 18.9180 46.1970 ;
        RECT 18.7840 45.1035 18.8100 46.1970 ;
        RECT 18.6760 45.1035 18.7020 46.1970 ;
        RECT 18.5680 45.1035 18.5940 46.1970 ;
        RECT 18.4600 45.1035 18.4860 46.1970 ;
        RECT 18.3520 45.1035 18.3780 46.1970 ;
        RECT 18.2440 45.1035 18.2700 46.1970 ;
        RECT 18.1360 45.1035 18.1620 46.1970 ;
        RECT 18.0280 45.1035 18.0540 46.1970 ;
        RECT 17.9200 45.1035 17.9460 46.1970 ;
        RECT 17.8120 45.1035 17.8380 46.1970 ;
        RECT 17.7040 45.1035 17.7300 46.1970 ;
        RECT 17.5960 45.1035 17.6220 46.1970 ;
        RECT 17.4880 45.1035 17.5140 46.1970 ;
        RECT 17.3800 45.1035 17.4060 46.1970 ;
        RECT 17.2720 45.1035 17.2980 46.1970 ;
        RECT 17.1640 45.1035 17.1900 46.1970 ;
        RECT 17.0560 45.1035 17.0820 46.1970 ;
        RECT 16.9480 45.1035 16.9740 46.1970 ;
        RECT 16.8400 45.1035 16.8660 46.1970 ;
        RECT 16.7320 45.1035 16.7580 46.1970 ;
        RECT 16.6240 45.1035 16.6500 46.1970 ;
        RECT 16.5160 45.1035 16.5420 46.1970 ;
        RECT 16.4080 45.1035 16.4340 46.1970 ;
        RECT 16.3000 45.1035 16.3260 46.1970 ;
        RECT 16.0870 45.1035 16.1640 46.1970 ;
        RECT 14.1940 45.1035 14.2710 46.1970 ;
        RECT 14.0320 45.1035 14.0580 46.1970 ;
        RECT 13.9240 45.1035 13.9500 46.1970 ;
        RECT 13.8160 45.1035 13.8420 46.1970 ;
        RECT 13.7080 45.1035 13.7340 46.1970 ;
        RECT 13.6000 45.1035 13.6260 46.1970 ;
        RECT 13.4920 45.1035 13.5180 46.1970 ;
        RECT 13.3840 45.1035 13.4100 46.1970 ;
        RECT 13.2760 45.1035 13.3020 46.1970 ;
        RECT 13.1680 45.1035 13.1940 46.1970 ;
        RECT 13.0600 45.1035 13.0860 46.1970 ;
        RECT 12.9520 45.1035 12.9780 46.1970 ;
        RECT 12.8440 45.1035 12.8700 46.1970 ;
        RECT 12.7360 45.1035 12.7620 46.1970 ;
        RECT 12.6280 45.1035 12.6540 46.1970 ;
        RECT 12.5200 45.1035 12.5460 46.1970 ;
        RECT 12.4120 45.1035 12.4380 46.1970 ;
        RECT 12.3040 45.1035 12.3300 46.1970 ;
        RECT 12.1960 45.1035 12.2220 46.1970 ;
        RECT 12.0880 45.1035 12.1140 46.1970 ;
        RECT 11.9800 45.1035 12.0060 46.1970 ;
        RECT 11.8720 45.1035 11.8980 46.1970 ;
        RECT 11.7640 45.1035 11.7900 46.1970 ;
        RECT 11.6560 45.1035 11.6820 46.1970 ;
        RECT 11.5480 45.1035 11.5740 46.1970 ;
        RECT 11.4400 45.1035 11.4660 46.1970 ;
        RECT 11.3320 45.1035 11.3580 46.1970 ;
        RECT 11.2240 45.1035 11.2500 46.1970 ;
        RECT 11.1160 45.1035 11.1420 46.1970 ;
        RECT 11.0080 45.1035 11.0340 46.1970 ;
        RECT 10.9000 45.1035 10.9260 46.1970 ;
        RECT 10.7920 45.1035 10.8180 46.1970 ;
        RECT 10.6840 45.1035 10.7100 46.1970 ;
        RECT 10.5760 45.1035 10.6020 46.1970 ;
        RECT 10.4680 45.1035 10.4940 46.1970 ;
        RECT 10.3600 45.1035 10.3860 46.1970 ;
        RECT 10.2520 45.1035 10.2780 46.1970 ;
        RECT 10.1440 45.1035 10.1700 46.1970 ;
        RECT 10.0360 45.1035 10.0620 46.1970 ;
        RECT 9.9280 45.1035 9.9540 46.1970 ;
        RECT 9.8200 45.1035 9.8460 46.1970 ;
        RECT 9.7120 45.1035 9.7380 46.1970 ;
        RECT 9.6040 45.1035 9.6300 46.1970 ;
        RECT 9.4960 45.1035 9.5220 46.1970 ;
        RECT 9.3880 45.1035 9.4140 46.1970 ;
        RECT 9.2800 45.1035 9.3060 46.1970 ;
        RECT 9.1720 45.1035 9.1980 46.1970 ;
        RECT 9.0640 45.1035 9.0900 46.1970 ;
        RECT 8.9560 45.1035 8.9820 46.1970 ;
        RECT 8.8480 45.1035 8.8740 46.1970 ;
        RECT 8.7400 45.1035 8.7660 46.1970 ;
        RECT 8.6320 45.1035 8.6580 46.1970 ;
        RECT 8.5240 45.1035 8.5500 46.1970 ;
        RECT 8.4160 45.1035 8.4420 46.1970 ;
        RECT 8.3080 45.1035 8.3340 46.1970 ;
        RECT 8.2000 45.1035 8.2260 46.1970 ;
        RECT 8.0920 45.1035 8.1180 46.1970 ;
        RECT 7.9840 45.1035 8.0100 46.1970 ;
        RECT 7.8760 45.1035 7.9020 46.1970 ;
        RECT 7.7680 45.1035 7.7940 46.1970 ;
        RECT 7.6600 45.1035 7.6860 46.1970 ;
        RECT 7.5520 45.1035 7.5780 46.1970 ;
        RECT 7.4440 45.1035 7.4700 46.1970 ;
        RECT 7.3360 45.1035 7.3620 46.1970 ;
        RECT 7.2280 45.1035 7.2540 46.1970 ;
        RECT 7.1200 45.1035 7.1460 46.1970 ;
        RECT 7.0120 45.1035 7.0380 46.1970 ;
        RECT 6.9040 45.1035 6.9300 46.1970 ;
        RECT 6.7960 45.1035 6.8220 46.1970 ;
        RECT 6.6880 45.1035 6.7140 46.1970 ;
        RECT 6.5800 45.1035 6.6060 46.1970 ;
        RECT 6.4720 45.1035 6.4980 46.1970 ;
        RECT 6.3640 45.1035 6.3900 46.1970 ;
        RECT 6.2560 45.1035 6.2820 46.1970 ;
        RECT 6.1480 45.1035 6.1740 46.1970 ;
        RECT 6.0400 45.1035 6.0660 46.1970 ;
        RECT 5.9320 45.1035 5.9580 46.1970 ;
        RECT 5.8240 45.1035 5.8500 46.1970 ;
        RECT 5.7160 45.1035 5.7420 46.1970 ;
        RECT 5.6080 45.1035 5.6340 46.1970 ;
        RECT 5.5000 45.1035 5.5260 46.1970 ;
        RECT 5.3920 45.1035 5.4180 46.1970 ;
        RECT 5.2840 45.1035 5.3100 46.1970 ;
        RECT 5.1760 45.1035 5.2020 46.1970 ;
        RECT 5.0680 45.1035 5.0940 46.1970 ;
        RECT 4.9600 45.1035 4.9860 46.1970 ;
        RECT 4.8520 45.1035 4.8780 46.1970 ;
        RECT 4.7440 45.1035 4.7700 46.1970 ;
        RECT 4.6360 45.1035 4.6620 46.1970 ;
        RECT 4.5280 45.1035 4.5540 46.1970 ;
        RECT 4.4200 45.1035 4.4460 46.1970 ;
        RECT 4.3120 45.1035 4.3380 46.1970 ;
        RECT 4.2040 45.1035 4.2300 46.1970 ;
        RECT 4.0960 45.1035 4.1220 46.1970 ;
        RECT 3.9880 45.1035 4.0140 46.1970 ;
        RECT 3.8800 45.1035 3.9060 46.1970 ;
        RECT 3.7720 45.1035 3.7980 46.1970 ;
        RECT 3.6640 45.1035 3.6900 46.1970 ;
        RECT 3.5560 45.1035 3.5820 46.1970 ;
        RECT 3.4480 45.1035 3.4740 46.1970 ;
        RECT 3.3400 45.1035 3.3660 46.1970 ;
        RECT 3.2320 45.1035 3.2580 46.1970 ;
        RECT 3.1240 45.1035 3.1500 46.1970 ;
        RECT 3.0160 45.1035 3.0420 46.1970 ;
        RECT 2.9080 45.1035 2.9340 46.1970 ;
        RECT 2.8000 45.1035 2.8260 46.1970 ;
        RECT 2.6920 45.1035 2.7180 46.1970 ;
        RECT 2.5840 45.1035 2.6100 46.1970 ;
        RECT 2.4760 45.1035 2.5020 46.1970 ;
        RECT 2.3680 45.1035 2.3940 46.1970 ;
        RECT 2.2600 45.1035 2.2860 46.1970 ;
        RECT 2.1520 45.1035 2.1780 46.1970 ;
        RECT 2.0440 45.1035 2.0700 46.1970 ;
        RECT 1.9360 45.1035 1.9620 46.1970 ;
        RECT 1.8280 45.1035 1.8540 46.1970 ;
        RECT 1.7200 45.1035 1.7460 46.1970 ;
        RECT 1.6120 45.1035 1.6380 46.1970 ;
        RECT 1.5040 45.1035 1.5300 46.1970 ;
        RECT 1.3960 45.1035 1.4220 46.1970 ;
        RECT 1.2880 45.1035 1.3140 46.1970 ;
        RECT 1.1800 45.1035 1.2060 46.1970 ;
        RECT 1.0720 45.1035 1.0980 46.1970 ;
        RECT 0.9640 45.1035 0.9900 46.1970 ;
        RECT 0.8560 45.1035 0.8820 46.1970 ;
        RECT 0.7480 45.1035 0.7740 46.1970 ;
        RECT 0.6400 45.1035 0.6660 46.1970 ;
        RECT 0.5320 45.1035 0.5580 46.1970 ;
        RECT 0.4240 45.1035 0.4500 46.1970 ;
        RECT 0.3160 45.1035 0.3420 46.1970 ;
        RECT 0.2080 45.1035 0.2340 46.1970 ;
        RECT 0.0050 45.1035 0.0900 46.1970 ;
        RECT 15.5530 46.1835 15.6810 47.2770 ;
        RECT 15.5390 46.8490 15.6810 47.1715 ;
        RECT 15.3190 46.5760 15.4530 47.2770 ;
        RECT 15.2960 46.9110 15.4530 47.1690 ;
        RECT 15.3190 46.1835 15.4170 47.2770 ;
        RECT 15.3190 46.3045 15.4310 46.5440 ;
        RECT 15.3190 46.1835 15.4530 46.2725 ;
        RECT 15.0940 46.6340 15.2280 47.2770 ;
        RECT 15.0940 46.1835 15.1920 47.2770 ;
        RECT 14.6770 46.1835 14.7600 47.2770 ;
        RECT 14.6770 46.2720 14.7740 47.2075 ;
        RECT 30.2680 46.1835 30.3530 47.2770 ;
        RECT 30.1240 46.1835 30.1500 47.2770 ;
        RECT 30.0160 46.1835 30.0420 47.2770 ;
        RECT 29.9080 46.1835 29.9340 47.2770 ;
        RECT 29.8000 46.1835 29.8260 47.2770 ;
        RECT 29.6920 46.1835 29.7180 47.2770 ;
        RECT 29.5840 46.1835 29.6100 47.2770 ;
        RECT 29.4760 46.1835 29.5020 47.2770 ;
        RECT 29.3680 46.1835 29.3940 47.2770 ;
        RECT 29.2600 46.1835 29.2860 47.2770 ;
        RECT 29.1520 46.1835 29.1780 47.2770 ;
        RECT 29.0440 46.1835 29.0700 47.2770 ;
        RECT 28.9360 46.1835 28.9620 47.2770 ;
        RECT 28.8280 46.1835 28.8540 47.2770 ;
        RECT 28.7200 46.1835 28.7460 47.2770 ;
        RECT 28.6120 46.1835 28.6380 47.2770 ;
        RECT 28.5040 46.1835 28.5300 47.2770 ;
        RECT 28.3960 46.1835 28.4220 47.2770 ;
        RECT 28.2880 46.1835 28.3140 47.2770 ;
        RECT 28.1800 46.1835 28.2060 47.2770 ;
        RECT 28.0720 46.1835 28.0980 47.2770 ;
        RECT 27.9640 46.1835 27.9900 47.2770 ;
        RECT 27.8560 46.1835 27.8820 47.2770 ;
        RECT 27.7480 46.1835 27.7740 47.2770 ;
        RECT 27.6400 46.1835 27.6660 47.2770 ;
        RECT 27.5320 46.1835 27.5580 47.2770 ;
        RECT 27.4240 46.1835 27.4500 47.2770 ;
        RECT 27.3160 46.1835 27.3420 47.2770 ;
        RECT 27.2080 46.1835 27.2340 47.2770 ;
        RECT 27.1000 46.1835 27.1260 47.2770 ;
        RECT 26.9920 46.1835 27.0180 47.2770 ;
        RECT 26.8840 46.1835 26.9100 47.2770 ;
        RECT 26.7760 46.1835 26.8020 47.2770 ;
        RECT 26.6680 46.1835 26.6940 47.2770 ;
        RECT 26.5600 46.1835 26.5860 47.2770 ;
        RECT 26.4520 46.1835 26.4780 47.2770 ;
        RECT 26.3440 46.1835 26.3700 47.2770 ;
        RECT 26.2360 46.1835 26.2620 47.2770 ;
        RECT 26.1280 46.1835 26.1540 47.2770 ;
        RECT 26.0200 46.1835 26.0460 47.2770 ;
        RECT 25.9120 46.1835 25.9380 47.2770 ;
        RECT 25.8040 46.1835 25.8300 47.2770 ;
        RECT 25.6960 46.1835 25.7220 47.2770 ;
        RECT 25.5880 46.1835 25.6140 47.2770 ;
        RECT 25.4800 46.1835 25.5060 47.2770 ;
        RECT 25.3720 46.1835 25.3980 47.2770 ;
        RECT 25.2640 46.1835 25.2900 47.2770 ;
        RECT 25.1560 46.1835 25.1820 47.2770 ;
        RECT 25.0480 46.1835 25.0740 47.2770 ;
        RECT 24.9400 46.1835 24.9660 47.2770 ;
        RECT 24.8320 46.1835 24.8580 47.2770 ;
        RECT 24.7240 46.1835 24.7500 47.2770 ;
        RECT 24.6160 46.1835 24.6420 47.2770 ;
        RECT 24.5080 46.1835 24.5340 47.2770 ;
        RECT 24.4000 46.1835 24.4260 47.2770 ;
        RECT 24.2920 46.1835 24.3180 47.2770 ;
        RECT 24.1840 46.1835 24.2100 47.2770 ;
        RECT 24.0760 46.1835 24.1020 47.2770 ;
        RECT 23.9680 46.1835 23.9940 47.2770 ;
        RECT 23.8600 46.1835 23.8860 47.2770 ;
        RECT 23.7520 46.1835 23.7780 47.2770 ;
        RECT 23.6440 46.1835 23.6700 47.2770 ;
        RECT 23.5360 46.1835 23.5620 47.2770 ;
        RECT 23.4280 46.1835 23.4540 47.2770 ;
        RECT 23.3200 46.1835 23.3460 47.2770 ;
        RECT 23.2120 46.1835 23.2380 47.2770 ;
        RECT 23.1040 46.1835 23.1300 47.2770 ;
        RECT 22.9960 46.1835 23.0220 47.2770 ;
        RECT 22.8880 46.1835 22.9140 47.2770 ;
        RECT 22.7800 46.1835 22.8060 47.2770 ;
        RECT 22.6720 46.1835 22.6980 47.2770 ;
        RECT 22.5640 46.1835 22.5900 47.2770 ;
        RECT 22.4560 46.1835 22.4820 47.2770 ;
        RECT 22.3480 46.1835 22.3740 47.2770 ;
        RECT 22.2400 46.1835 22.2660 47.2770 ;
        RECT 22.1320 46.1835 22.1580 47.2770 ;
        RECT 22.0240 46.1835 22.0500 47.2770 ;
        RECT 21.9160 46.1835 21.9420 47.2770 ;
        RECT 21.8080 46.1835 21.8340 47.2770 ;
        RECT 21.7000 46.1835 21.7260 47.2770 ;
        RECT 21.5920 46.1835 21.6180 47.2770 ;
        RECT 21.4840 46.1835 21.5100 47.2770 ;
        RECT 21.3760 46.1835 21.4020 47.2770 ;
        RECT 21.2680 46.1835 21.2940 47.2770 ;
        RECT 21.1600 46.1835 21.1860 47.2770 ;
        RECT 21.0520 46.1835 21.0780 47.2770 ;
        RECT 20.9440 46.1835 20.9700 47.2770 ;
        RECT 20.8360 46.1835 20.8620 47.2770 ;
        RECT 20.7280 46.1835 20.7540 47.2770 ;
        RECT 20.6200 46.1835 20.6460 47.2770 ;
        RECT 20.5120 46.1835 20.5380 47.2770 ;
        RECT 20.4040 46.1835 20.4300 47.2770 ;
        RECT 20.2960 46.1835 20.3220 47.2770 ;
        RECT 20.1880 46.1835 20.2140 47.2770 ;
        RECT 20.0800 46.1835 20.1060 47.2770 ;
        RECT 19.9720 46.1835 19.9980 47.2770 ;
        RECT 19.8640 46.1835 19.8900 47.2770 ;
        RECT 19.7560 46.1835 19.7820 47.2770 ;
        RECT 19.6480 46.1835 19.6740 47.2770 ;
        RECT 19.5400 46.1835 19.5660 47.2770 ;
        RECT 19.4320 46.1835 19.4580 47.2770 ;
        RECT 19.3240 46.1835 19.3500 47.2770 ;
        RECT 19.2160 46.1835 19.2420 47.2770 ;
        RECT 19.1080 46.1835 19.1340 47.2770 ;
        RECT 19.0000 46.1835 19.0260 47.2770 ;
        RECT 18.8920 46.1835 18.9180 47.2770 ;
        RECT 18.7840 46.1835 18.8100 47.2770 ;
        RECT 18.6760 46.1835 18.7020 47.2770 ;
        RECT 18.5680 46.1835 18.5940 47.2770 ;
        RECT 18.4600 46.1835 18.4860 47.2770 ;
        RECT 18.3520 46.1835 18.3780 47.2770 ;
        RECT 18.2440 46.1835 18.2700 47.2770 ;
        RECT 18.1360 46.1835 18.1620 47.2770 ;
        RECT 18.0280 46.1835 18.0540 47.2770 ;
        RECT 17.9200 46.1835 17.9460 47.2770 ;
        RECT 17.8120 46.1835 17.8380 47.2770 ;
        RECT 17.7040 46.1835 17.7300 47.2770 ;
        RECT 17.5960 46.1835 17.6220 47.2770 ;
        RECT 17.4880 46.1835 17.5140 47.2770 ;
        RECT 17.3800 46.1835 17.4060 47.2770 ;
        RECT 17.2720 46.1835 17.2980 47.2770 ;
        RECT 17.1640 46.1835 17.1900 47.2770 ;
        RECT 17.0560 46.1835 17.0820 47.2770 ;
        RECT 16.9480 46.1835 16.9740 47.2770 ;
        RECT 16.8400 46.1835 16.8660 47.2770 ;
        RECT 16.7320 46.1835 16.7580 47.2770 ;
        RECT 16.6240 46.1835 16.6500 47.2770 ;
        RECT 16.5160 46.1835 16.5420 47.2770 ;
        RECT 16.4080 46.1835 16.4340 47.2770 ;
        RECT 16.3000 46.1835 16.3260 47.2770 ;
        RECT 16.0870 46.1835 16.1640 47.2770 ;
        RECT 14.1940 46.1835 14.2710 47.2770 ;
        RECT 14.0320 46.1835 14.0580 47.2770 ;
        RECT 13.9240 46.1835 13.9500 47.2770 ;
        RECT 13.8160 46.1835 13.8420 47.2770 ;
        RECT 13.7080 46.1835 13.7340 47.2770 ;
        RECT 13.6000 46.1835 13.6260 47.2770 ;
        RECT 13.4920 46.1835 13.5180 47.2770 ;
        RECT 13.3840 46.1835 13.4100 47.2770 ;
        RECT 13.2760 46.1835 13.3020 47.2770 ;
        RECT 13.1680 46.1835 13.1940 47.2770 ;
        RECT 13.0600 46.1835 13.0860 47.2770 ;
        RECT 12.9520 46.1835 12.9780 47.2770 ;
        RECT 12.8440 46.1835 12.8700 47.2770 ;
        RECT 12.7360 46.1835 12.7620 47.2770 ;
        RECT 12.6280 46.1835 12.6540 47.2770 ;
        RECT 12.5200 46.1835 12.5460 47.2770 ;
        RECT 12.4120 46.1835 12.4380 47.2770 ;
        RECT 12.3040 46.1835 12.3300 47.2770 ;
        RECT 12.1960 46.1835 12.2220 47.2770 ;
        RECT 12.0880 46.1835 12.1140 47.2770 ;
        RECT 11.9800 46.1835 12.0060 47.2770 ;
        RECT 11.8720 46.1835 11.8980 47.2770 ;
        RECT 11.7640 46.1835 11.7900 47.2770 ;
        RECT 11.6560 46.1835 11.6820 47.2770 ;
        RECT 11.5480 46.1835 11.5740 47.2770 ;
        RECT 11.4400 46.1835 11.4660 47.2770 ;
        RECT 11.3320 46.1835 11.3580 47.2770 ;
        RECT 11.2240 46.1835 11.2500 47.2770 ;
        RECT 11.1160 46.1835 11.1420 47.2770 ;
        RECT 11.0080 46.1835 11.0340 47.2770 ;
        RECT 10.9000 46.1835 10.9260 47.2770 ;
        RECT 10.7920 46.1835 10.8180 47.2770 ;
        RECT 10.6840 46.1835 10.7100 47.2770 ;
        RECT 10.5760 46.1835 10.6020 47.2770 ;
        RECT 10.4680 46.1835 10.4940 47.2770 ;
        RECT 10.3600 46.1835 10.3860 47.2770 ;
        RECT 10.2520 46.1835 10.2780 47.2770 ;
        RECT 10.1440 46.1835 10.1700 47.2770 ;
        RECT 10.0360 46.1835 10.0620 47.2770 ;
        RECT 9.9280 46.1835 9.9540 47.2770 ;
        RECT 9.8200 46.1835 9.8460 47.2770 ;
        RECT 9.7120 46.1835 9.7380 47.2770 ;
        RECT 9.6040 46.1835 9.6300 47.2770 ;
        RECT 9.4960 46.1835 9.5220 47.2770 ;
        RECT 9.3880 46.1835 9.4140 47.2770 ;
        RECT 9.2800 46.1835 9.3060 47.2770 ;
        RECT 9.1720 46.1835 9.1980 47.2770 ;
        RECT 9.0640 46.1835 9.0900 47.2770 ;
        RECT 8.9560 46.1835 8.9820 47.2770 ;
        RECT 8.8480 46.1835 8.8740 47.2770 ;
        RECT 8.7400 46.1835 8.7660 47.2770 ;
        RECT 8.6320 46.1835 8.6580 47.2770 ;
        RECT 8.5240 46.1835 8.5500 47.2770 ;
        RECT 8.4160 46.1835 8.4420 47.2770 ;
        RECT 8.3080 46.1835 8.3340 47.2770 ;
        RECT 8.2000 46.1835 8.2260 47.2770 ;
        RECT 8.0920 46.1835 8.1180 47.2770 ;
        RECT 7.9840 46.1835 8.0100 47.2770 ;
        RECT 7.8760 46.1835 7.9020 47.2770 ;
        RECT 7.7680 46.1835 7.7940 47.2770 ;
        RECT 7.6600 46.1835 7.6860 47.2770 ;
        RECT 7.5520 46.1835 7.5780 47.2770 ;
        RECT 7.4440 46.1835 7.4700 47.2770 ;
        RECT 7.3360 46.1835 7.3620 47.2770 ;
        RECT 7.2280 46.1835 7.2540 47.2770 ;
        RECT 7.1200 46.1835 7.1460 47.2770 ;
        RECT 7.0120 46.1835 7.0380 47.2770 ;
        RECT 6.9040 46.1835 6.9300 47.2770 ;
        RECT 6.7960 46.1835 6.8220 47.2770 ;
        RECT 6.6880 46.1835 6.7140 47.2770 ;
        RECT 6.5800 46.1835 6.6060 47.2770 ;
        RECT 6.4720 46.1835 6.4980 47.2770 ;
        RECT 6.3640 46.1835 6.3900 47.2770 ;
        RECT 6.2560 46.1835 6.2820 47.2770 ;
        RECT 6.1480 46.1835 6.1740 47.2770 ;
        RECT 6.0400 46.1835 6.0660 47.2770 ;
        RECT 5.9320 46.1835 5.9580 47.2770 ;
        RECT 5.8240 46.1835 5.8500 47.2770 ;
        RECT 5.7160 46.1835 5.7420 47.2770 ;
        RECT 5.6080 46.1835 5.6340 47.2770 ;
        RECT 5.5000 46.1835 5.5260 47.2770 ;
        RECT 5.3920 46.1835 5.4180 47.2770 ;
        RECT 5.2840 46.1835 5.3100 47.2770 ;
        RECT 5.1760 46.1835 5.2020 47.2770 ;
        RECT 5.0680 46.1835 5.0940 47.2770 ;
        RECT 4.9600 46.1835 4.9860 47.2770 ;
        RECT 4.8520 46.1835 4.8780 47.2770 ;
        RECT 4.7440 46.1835 4.7700 47.2770 ;
        RECT 4.6360 46.1835 4.6620 47.2770 ;
        RECT 4.5280 46.1835 4.5540 47.2770 ;
        RECT 4.4200 46.1835 4.4460 47.2770 ;
        RECT 4.3120 46.1835 4.3380 47.2770 ;
        RECT 4.2040 46.1835 4.2300 47.2770 ;
        RECT 4.0960 46.1835 4.1220 47.2770 ;
        RECT 3.9880 46.1835 4.0140 47.2770 ;
        RECT 3.8800 46.1835 3.9060 47.2770 ;
        RECT 3.7720 46.1835 3.7980 47.2770 ;
        RECT 3.6640 46.1835 3.6900 47.2770 ;
        RECT 3.5560 46.1835 3.5820 47.2770 ;
        RECT 3.4480 46.1835 3.4740 47.2770 ;
        RECT 3.3400 46.1835 3.3660 47.2770 ;
        RECT 3.2320 46.1835 3.2580 47.2770 ;
        RECT 3.1240 46.1835 3.1500 47.2770 ;
        RECT 3.0160 46.1835 3.0420 47.2770 ;
        RECT 2.9080 46.1835 2.9340 47.2770 ;
        RECT 2.8000 46.1835 2.8260 47.2770 ;
        RECT 2.6920 46.1835 2.7180 47.2770 ;
        RECT 2.5840 46.1835 2.6100 47.2770 ;
        RECT 2.4760 46.1835 2.5020 47.2770 ;
        RECT 2.3680 46.1835 2.3940 47.2770 ;
        RECT 2.2600 46.1835 2.2860 47.2770 ;
        RECT 2.1520 46.1835 2.1780 47.2770 ;
        RECT 2.0440 46.1835 2.0700 47.2770 ;
        RECT 1.9360 46.1835 1.9620 47.2770 ;
        RECT 1.8280 46.1835 1.8540 47.2770 ;
        RECT 1.7200 46.1835 1.7460 47.2770 ;
        RECT 1.6120 46.1835 1.6380 47.2770 ;
        RECT 1.5040 46.1835 1.5300 47.2770 ;
        RECT 1.3960 46.1835 1.4220 47.2770 ;
        RECT 1.2880 46.1835 1.3140 47.2770 ;
        RECT 1.1800 46.1835 1.2060 47.2770 ;
        RECT 1.0720 46.1835 1.0980 47.2770 ;
        RECT 0.9640 46.1835 0.9900 47.2770 ;
        RECT 0.8560 46.1835 0.8820 47.2770 ;
        RECT 0.7480 46.1835 0.7740 47.2770 ;
        RECT 0.6400 46.1835 0.6660 47.2770 ;
        RECT 0.5320 46.1835 0.5580 47.2770 ;
        RECT 0.4240 46.1835 0.4500 47.2770 ;
        RECT 0.3160 46.1835 0.3420 47.2770 ;
        RECT 0.2080 46.1835 0.2340 47.2770 ;
        RECT 0.0050 46.1835 0.0900 47.2770 ;
        RECT 15.5530 47.2635 15.6810 48.3570 ;
        RECT 15.5390 47.9290 15.6810 48.2515 ;
        RECT 15.3190 47.6560 15.4530 48.3570 ;
        RECT 15.2960 47.9910 15.4530 48.2490 ;
        RECT 15.3190 47.2635 15.4170 48.3570 ;
        RECT 15.3190 47.3845 15.4310 47.6240 ;
        RECT 15.3190 47.2635 15.4530 47.3525 ;
        RECT 15.0940 47.7140 15.2280 48.3570 ;
        RECT 15.0940 47.2635 15.1920 48.3570 ;
        RECT 14.6770 47.2635 14.7600 48.3570 ;
        RECT 14.6770 47.3520 14.7740 48.2875 ;
        RECT 30.2680 47.2635 30.3530 48.3570 ;
        RECT 30.1240 47.2635 30.1500 48.3570 ;
        RECT 30.0160 47.2635 30.0420 48.3570 ;
        RECT 29.9080 47.2635 29.9340 48.3570 ;
        RECT 29.8000 47.2635 29.8260 48.3570 ;
        RECT 29.6920 47.2635 29.7180 48.3570 ;
        RECT 29.5840 47.2635 29.6100 48.3570 ;
        RECT 29.4760 47.2635 29.5020 48.3570 ;
        RECT 29.3680 47.2635 29.3940 48.3570 ;
        RECT 29.2600 47.2635 29.2860 48.3570 ;
        RECT 29.1520 47.2635 29.1780 48.3570 ;
        RECT 29.0440 47.2635 29.0700 48.3570 ;
        RECT 28.9360 47.2635 28.9620 48.3570 ;
        RECT 28.8280 47.2635 28.8540 48.3570 ;
        RECT 28.7200 47.2635 28.7460 48.3570 ;
        RECT 28.6120 47.2635 28.6380 48.3570 ;
        RECT 28.5040 47.2635 28.5300 48.3570 ;
        RECT 28.3960 47.2635 28.4220 48.3570 ;
        RECT 28.2880 47.2635 28.3140 48.3570 ;
        RECT 28.1800 47.2635 28.2060 48.3570 ;
        RECT 28.0720 47.2635 28.0980 48.3570 ;
        RECT 27.9640 47.2635 27.9900 48.3570 ;
        RECT 27.8560 47.2635 27.8820 48.3570 ;
        RECT 27.7480 47.2635 27.7740 48.3570 ;
        RECT 27.6400 47.2635 27.6660 48.3570 ;
        RECT 27.5320 47.2635 27.5580 48.3570 ;
        RECT 27.4240 47.2635 27.4500 48.3570 ;
        RECT 27.3160 47.2635 27.3420 48.3570 ;
        RECT 27.2080 47.2635 27.2340 48.3570 ;
        RECT 27.1000 47.2635 27.1260 48.3570 ;
        RECT 26.9920 47.2635 27.0180 48.3570 ;
        RECT 26.8840 47.2635 26.9100 48.3570 ;
        RECT 26.7760 47.2635 26.8020 48.3570 ;
        RECT 26.6680 47.2635 26.6940 48.3570 ;
        RECT 26.5600 47.2635 26.5860 48.3570 ;
        RECT 26.4520 47.2635 26.4780 48.3570 ;
        RECT 26.3440 47.2635 26.3700 48.3570 ;
        RECT 26.2360 47.2635 26.2620 48.3570 ;
        RECT 26.1280 47.2635 26.1540 48.3570 ;
        RECT 26.0200 47.2635 26.0460 48.3570 ;
        RECT 25.9120 47.2635 25.9380 48.3570 ;
        RECT 25.8040 47.2635 25.8300 48.3570 ;
        RECT 25.6960 47.2635 25.7220 48.3570 ;
        RECT 25.5880 47.2635 25.6140 48.3570 ;
        RECT 25.4800 47.2635 25.5060 48.3570 ;
        RECT 25.3720 47.2635 25.3980 48.3570 ;
        RECT 25.2640 47.2635 25.2900 48.3570 ;
        RECT 25.1560 47.2635 25.1820 48.3570 ;
        RECT 25.0480 47.2635 25.0740 48.3570 ;
        RECT 24.9400 47.2635 24.9660 48.3570 ;
        RECT 24.8320 47.2635 24.8580 48.3570 ;
        RECT 24.7240 47.2635 24.7500 48.3570 ;
        RECT 24.6160 47.2635 24.6420 48.3570 ;
        RECT 24.5080 47.2635 24.5340 48.3570 ;
        RECT 24.4000 47.2635 24.4260 48.3570 ;
        RECT 24.2920 47.2635 24.3180 48.3570 ;
        RECT 24.1840 47.2635 24.2100 48.3570 ;
        RECT 24.0760 47.2635 24.1020 48.3570 ;
        RECT 23.9680 47.2635 23.9940 48.3570 ;
        RECT 23.8600 47.2635 23.8860 48.3570 ;
        RECT 23.7520 47.2635 23.7780 48.3570 ;
        RECT 23.6440 47.2635 23.6700 48.3570 ;
        RECT 23.5360 47.2635 23.5620 48.3570 ;
        RECT 23.4280 47.2635 23.4540 48.3570 ;
        RECT 23.3200 47.2635 23.3460 48.3570 ;
        RECT 23.2120 47.2635 23.2380 48.3570 ;
        RECT 23.1040 47.2635 23.1300 48.3570 ;
        RECT 22.9960 47.2635 23.0220 48.3570 ;
        RECT 22.8880 47.2635 22.9140 48.3570 ;
        RECT 22.7800 47.2635 22.8060 48.3570 ;
        RECT 22.6720 47.2635 22.6980 48.3570 ;
        RECT 22.5640 47.2635 22.5900 48.3570 ;
        RECT 22.4560 47.2635 22.4820 48.3570 ;
        RECT 22.3480 47.2635 22.3740 48.3570 ;
        RECT 22.2400 47.2635 22.2660 48.3570 ;
        RECT 22.1320 47.2635 22.1580 48.3570 ;
        RECT 22.0240 47.2635 22.0500 48.3570 ;
        RECT 21.9160 47.2635 21.9420 48.3570 ;
        RECT 21.8080 47.2635 21.8340 48.3570 ;
        RECT 21.7000 47.2635 21.7260 48.3570 ;
        RECT 21.5920 47.2635 21.6180 48.3570 ;
        RECT 21.4840 47.2635 21.5100 48.3570 ;
        RECT 21.3760 47.2635 21.4020 48.3570 ;
        RECT 21.2680 47.2635 21.2940 48.3570 ;
        RECT 21.1600 47.2635 21.1860 48.3570 ;
        RECT 21.0520 47.2635 21.0780 48.3570 ;
        RECT 20.9440 47.2635 20.9700 48.3570 ;
        RECT 20.8360 47.2635 20.8620 48.3570 ;
        RECT 20.7280 47.2635 20.7540 48.3570 ;
        RECT 20.6200 47.2635 20.6460 48.3570 ;
        RECT 20.5120 47.2635 20.5380 48.3570 ;
        RECT 20.4040 47.2635 20.4300 48.3570 ;
        RECT 20.2960 47.2635 20.3220 48.3570 ;
        RECT 20.1880 47.2635 20.2140 48.3570 ;
        RECT 20.0800 47.2635 20.1060 48.3570 ;
        RECT 19.9720 47.2635 19.9980 48.3570 ;
        RECT 19.8640 47.2635 19.8900 48.3570 ;
        RECT 19.7560 47.2635 19.7820 48.3570 ;
        RECT 19.6480 47.2635 19.6740 48.3570 ;
        RECT 19.5400 47.2635 19.5660 48.3570 ;
        RECT 19.4320 47.2635 19.4580 48.3570 ;
        RECT 19.3240 47.2635 19.3500 48.3570 ;
        RECT 19.2160 47.2635 19.2420 48.3570 ;
        RECT 19.1080 47.2635 19.1340 48.3570 ;
        RECT 19.0000 47.2635 19.0260 48.3570 ;
        RECT 18.8920 47.2635 18.9180 48.3570 ;
        RECT 18.7840 47.2635 18.8100 48.3570 ;
        RECT 18.6760 47.2635 18.7020 48.3570 ;
        RECT 18.5680 47.2635 18.5940 48.3570 ;
        RECT 18.4600 47.2635 18.4860 48.3570 ;
        RECT 18.3520 47.2635 18.3780 48.3570 ;
        RECT 18.2440 47.2635 18.2700 48.3570 ;
        RECT 18.1360 47.2635 18.1620 48.3570 ;
        RECT 18.0280 47.2635 18.0540 48.3570 ;
        RECT 17.9200 47.2635 17.9460 48.3570 ;
        RECT 17.8120 47.2635 17.8380 48.3570 ;
        RECT 17.7040 47.2635 17.7300 48.3570 ;
        RECT 17.5960 47.2635 17.6220 48.3570 ;
        RECT 17.4880 47.2635 17.5140 48.3570 ;
        RECT 17.3800 47.2635 17.4060 48.3570 ;
        RECT 17.2720 47.2635 17.2980 48.3570 ;
        RECT 17.1640 47.2635 17.1900 48.3570 ;
        RECT 17.0560 47.2635 17.0820 48.3570 ;
        RECT 16.9480 47.2635 16.9740 48.3570 ;
        RECT 16.8400 47.2635 16.8660 48.3570 ;
        RECT 16.7320 47.2635 16.7580 48.3570 ;
        RECT 16.6240 47.2635 16.6500 48.3570 ;
        RECT 16.5160 47.2635 16.5420 48.3570 ;
        RECT 16.4080 47.2635 16.4340 48.3570 ;
        RECT 16.3000 47.2635 16.3260 48.3570 ;
        RECT 16.0870 47.2635 16.1640 48.3570 ;
        RECT 14.1940 47.2635 14.2710 48.3570 ;
        RECT 14.0320 47.2635 14.0580 48.3570 ;
        RECT 13.9240 47.2635 13.9500 48.3570 ;
        RECT 13.8160 47.2635 13.8420 48.3570 ;
        RECT 13.7080 47.2635 13.7340 48.3570 ;
        RECT 13.6000 47.2635 13.6260 48.3570 ;
        RECT 13.4920 47.2635 13.5180 48.3570 ;
        RECT 13.3840 47.2635 13.4100 48.3570 ;
        RECT 13.2760 47.2635 13.3020 48.3570 ;
        RECT 13.1680 47.2635 13.1940 48.3570 ;
        RECT 13.0600 47.2635 13.0860 48.3570 ;
        RECT 12.9520 47.2635 12.9780 48.3570 ;
        RECT 12.8440 47.2635 12.8700 48.3570 ;
        RECT 12.7360 47.2635 12.7620 48.3570 ;
        RECT 12.6280 47.2635 12.6540 48.3570 ;
        RECT 12.5200 47.2635 12.5460 48.3570 ;
        RECT 12.4120 47.2635 12.4380 48.3570 ;
        RECT 12.3040 47.2635 12.3300 48.3570 ;
        RECT 12.1960 47.2635 12.2220 48.3570 ;
        RECT 12.0880 47.2635 12.1140 48.3570 ;
        RECT 11.9800 47.2635 12.0060 48.3570 ;
        RECT 11.8720 47.2635 11.8980 48.3570 ;
        RECT 11.7640 47.2635 11.7900 48.3570 ;
        RECT 11.6560 47.2635 11.6820 48.3570 ;
        RECT 11.5480 47.2635 11.5740 48.3570 ;
        RECT 11.4400 47.2635 11.4660 48.3570 ;
        RECT 11.3320 47.2635 11.3580 48.3570 ;
        RECT 11.2240 47.2635 11.2500 48.3570 ;
        RECT 11.1160 47.2635 11.1420 48.3570 ;
        RECT 11.0080 47.2635 11.0340 48.3570 ;
        RECT 10.9000 47.2635 10.9260 48.3570 ;
        RECT 10.7920 47.2635 10.8180 48.3570 ;
        RECT 10.6840 47.2635 10.7100 48.3570 ;
        RECT 10.5760 47.2635 10.6020 48.3570 ;
        RECT 10.4680 47.2635 10.4940 48.3570 ;
        RECT 10.3600 47.2635 10.3860 48.3570 ;
        RECT 10.2520 47.2635 10.2780 48.3570 ;
        RECT 10.1440 47.2635 10.1700 48.3570 ;
        RECT 10.0360 47.2635 10.0620 48.3570 ;
        RECT 9.9280 47.2635 9.9540 48.3570 ;
        RECT 9.8200 47.2635 9.8460 48.3570 ;
        RECT 9.7120 47.2635 9.7380 48.3570 ;
        RECT 9.6040 47.2635 9.6300 48.3570 ;
        RECT 9.4960 47.2635 9.5220 48.3570 ;
        RECT 9.3880 47.2635 9.4140 48.3570 ;
        RECT 9.2800 47.2635 9.3060 48.3570 ;
        RECT 9.1720 47.2635 9.1980 48.3570 ;
        RECT 9.0640 47.2635 9.0900 48.3570 ;
        RECT 8.9560 47.2635 8.9820 48.3570 ;
        RECT 8.8480 47.2635 8.8740 48.3570 ;
        RECT 8.7400 47.2635 8.7660 48.3570 ;
        RECT 8.6320 47.2635 8.6580 48.3570 ;
        RECT 8.5240 47.2635 8.5500 48.3570 ;
        RECT 8.4160 47.2635 8.4420 48.3570 ;
        RECT 8.3080 47.2635 8.3340 48.3570 ;
        RECT 8.2000 47.2635 8.2260 48.3570 ;
        RECT 8.0920 47.2635 8.1180 48.3570 ;
        RECT 7.9840 47.2635 8.0100 48.3570 ;
        RECT 7.8760 47.2635 7.9020 48.3570 ;
        RECT 7.7680 47.2635 7.7940 48.3570 ;
        RECT 7.6600 47.2635 7.6860 48.3570 ;
        RECT 7.5520 47.2635 7.5780 48.3570 ;
        RECT 7.4440 47.2635 7.4700 48.3570 ;
        RECT 7.3360 47.2635 7.3620 48.3570 ;
        RECT 7.2280 47.2635 7.2540 48.3570 ;
        RECT 7.1200 47.2635 7.1460 48.3570 ;
        RECT 7.0120 47.2635 7.0380 48.3570 ;
        RECT 6.9040 47.2635 6.9300 48.3570 ;
        RECT 6.7960 47.2635 6.8220 48.3570 ;
        RECT 6.6880 47.2635 6.7140 48.3570 ;
        RECT 6.5800 47.2635 6.6060 48.3570 ;
        RECT 6.4720 47.2635 6.4980 48.3570 ;
        RECT 6.3640 47.2635 6.3900 48.3570 ;
        RECT 6.2560 47.2635 6.2820 48.3570 ;
        RECT 6.1480 47.2635 6.1740 48.3570 ;
        RECT 6.0400 47.2635 6.0660 48.3570 ;
        RECT 5.9320 47.2635 5.9580 48.3570 ;
        RECT 5.8240 47.2635 5.8500 48.3570 ;
        RECT 5.7160 47.2635 5.7420 48.3570 ;
        RECT 5.6080 47.2635 5.6340 48.3570 ;
        RECT 5.5000 47.2635 5.5260 48.3570 ;
        RECT 5.3920 47.2635 5.4180 48.3570 ;
        RECT 5.2840 47.2635 5.3100 48.3570 ;
        RECT 5.1760 47.2635 5.2020 48.3570 ;
        RECT 5.0680 47.2635 5.0940 48.3570 ;
        RECT 4.9600 47.2635 4.9860 48.3570 ;
        RECT 4.8520 47.2635 4.8780 48.3570 ;
        RECT 4.7440 47.2635 4.7700 48.3570 ;
        RECT 4.6360 47.2635 4.6620 48.3570 ;
        RECT 4.5280 47.2635 4.5540 48.3570 ;
        RECT 4.4200 47.2635 4.4460 48.3570 ;
        RECT 4.3120 47.2635 4.3380 48.3570 ;
        RECT 4.2040 47.2635 4.2300 48.3570 ;
        RECT 4.0960 47.2635 4.1220 48.3570 ;
        RECT 3.9880 47.2635 4.0140 48.3570 ;
        RECT 3.8800 47.2635 3.9060 48.3570 ;
        RECT 3.7720 47.2635 3.7980 48.3570 ;
        RECT 3.6640 47.2635 3.6900 48.3570 ;
        RECT 3.5560 47.2635 3.5820 48.3570 ;
        RECT 3.4480 47.2635 3.4740 48.3570 ;
        RECT 3.3400 47.2635 3.3660 48.3570 ;
        RECT 3.2320 47.2635 3.2580 48.3570 ;
        RECT 3.1240 47.2635 3.1500 48.3570 ;
        RECT 3.0160 47.2635 3.0420 48.3570 ;
        RECT 2.9080 47.2635 2.9340 48.3570 ;
        RECT 2.8000 47.2635 2.8260 48.3570 ;
        RECT 2.6920 47.2635 2.7180 48.3570 ;
        RECT 2.5840 47.2635 2.6100 48.3570 ;
        RECT 2.4760 47.2635 2.5020 48.3570 ;
        RECT 2.3680 47.2635 2.3940 48.3570 ;
        RECT 2.2600 47.2635 2.2860 48.3570 ;
        RECT 2.1520 47.2635 2.1780 48.3570 ;
        RECT 2.0440 47.2635 2.0700 48.3570 ;
        RECT 1.9360 47.2635 1.9620 48.3570 ;
        RECT 1.8280 47.2635 1.8540 48.3570 ;
        RECT 1.7200 47.2635 1.7460 48.3570 ;
        RECT 1.6120 47.2635 1.6380 48.3570 ;
        RECT 1.5040 47.2635 1.5300 48.3570 ;
        RECT 1.3960 47.2635 1.4220 48.3570 ;
        RECT 1.2880 47.2635 1.3140 48.3570 ;
        RECT 1.1800 47.2635 1.2060 48.3570 ;
        RECT 1.0720 47.2635 1.0980 48.3570 ;
        RECT 0.9640 47.2635 0.9900 48.3570 ;
        RECT 0.8560 47.2635 0.8820 48.3570 ;
        RECT 0.7480 47.2635 0.7740 48.3570 ;
        RECT 0.6400 47.2635 0.6660 48.3570 ;
        RECT 0.5320 47.2635 0.5580 48.3570 ;
        RECT 0.4240 47.2635 0.4500 48.3570 ;
        RECT 0.3160 47.2635 0.3420 48.3570 ;
        RECT 0.2080 47.2635 0.2340 48.3570 ;
        RECT 0.0050 47.2635 0.0900 48.3570 ;
        RECT 15.5530 48.3435 15.6810 49.4370 ;
        RECT 15.5390 49.0090 15.6810 49.3315 ;
        RECT 15.3190 48.7360 15.4530 49.4370 ;
        RECT 15.2960 49.0710 15.4530 49.3290 ;
        RECT 15.3190 48.3435 15.4170 49.4370 ;
        RECT 15.3190 48.4645 15.4310 48.7040 ;
        RECT 15.3190 48.3435 15.4530 48.4325 ;
        RECT 15.0940 48.7940 15.2280 49.4370 ;
        RECT 15.0940 48.3435 15.1920 49.4370 ;
        RECT 14.6770 48.3435 14.7600 49.4370 ;
        RECT 14.6770 48.4320 14.7740 49.3675 ;
        RECT 30.2680 48.3435 30.3530 49.4370 ;
        RECT 30.1240 48.3435 30.1500 49.4370 ;
        RECT 30.0160 48.3435 30.0420 49.4370 ;
        RECT 29.9080 48.3435 29.9340 49.4370 ;
        RECT 29.8000 48.3435 29.8260 49.4370 ;
        RECT 29.6920 48.3435 29.7180 49.4370 ;
        RECT 29.5840 48.3435 29.6100 49.4370 ;
        RECT 29.4760 48.3435 29.5020 49.4370 ;
        RECT 29.3680 48.3435 29.3940 49.4370 ;
        RECT 29.2600 48.3435 29.2860 49.4370 ;
        RECT 29.1520 48.3435 29.1780 49.4370 ;
        RECT 29.0440 48.3435 29.0700 49.4370 ;
        RECT 28.9360 48.3435 28.9620 49.4370 ;
        RECT 28.8280 48.3435 28.8540 49.4370 ;
        RECT 28.7200 48.3435 28.7460 49.4370 ;
        RECT 28.6120 48.3435 28.6380 49.4370 ;
        RECT 28.5040 48.3435 28.5300 49.4370 ;
        RECT 28.3960 48.3435 28.4220 49.4370 ;
        RECT 28.2880 48.3435 28.3140 49.4370 ;
        RECT 28.1800 48.3435 28.2060 49.4370 ;
        RECT 28.0720 48.3435 28.0980 49.4370 ;
        RECT 27.9640 48.3435 27.9900 49.4370 ;
        RECT 27.8560 48.3435 27.8820 49.4370 ;
        RECT 27.7480 48.3435 27.7740 49.4370 ;
        RECT 27.6400 48.3435 27.6660 49.4370 ;
        RECT 27.5320 48.3435 27.5580 49.4370 ;
        RECT 27.4240 48.3435 27.4500 49.4370 ;
        RECT 27.3160 48.3435 27.3420 49.4370 ;
        RECT 27.2080 48.3435 27.2340 49.4370 ;
        RECT 27.1000 48.3435 27.1260 49.4370 ;
        RECT 26.9920 48.3435 27.0180 49.4370 ;
        RECT 26.8840 48.3435 26.9100 49.4370 ;
        RECT 26.7760 48.3435 26.8020 49.4370 ;
        RECT 26.6680 48.3435 26.6940 49.4370 ;
        RECT 26.5600 48.3435 26.5860 49.4370 ;
        RECT 26.4520 48.3435 26.4780 49.4370 ;
        RECT 26.3440 48.3435 26.3700 49.4370 ;
        RECT 26.2360 48.3435 26.2620 49.4370 ;
        RECT 26.1280 48.3435 26.1540 49.4370 ;
        RECT 26.0200 48.3435 26.0460 49.4370 ;
        RECT 25.9120 48.3435 25.9380 49.4370 ;
        RECT 25.8040 48.3435 25.8300 49.4370 ;
        RECT 25.6960 48.3435 25.7220 49.4370 ;
        RECT 25.5880 48.3435 25.6140 49.4370 ;
        RECT 25.4800 48.3435 25.5060 49.4370 ;
        RECT 25.3720 48.3435 25.3980 49.4370 ;
        RECT 25.2640 48.3435 25.2900 49.4370 ;
        RECT 25.1560 48.3435 25.1820 49.4370 ;
        RECT 25.0480 48.3435 25.0740 49.4370 ;
        RECT 24.9400 48.3435 24.9660 49.4370 ;
        RECT 24.8320 48.3435 24.8580 49.4370 ;
        RECT 24.7240 48.3435 24.7500 49.4370 ;
        RECT 24.6160 48.3435 24.6420 49.4370 ;
        RECT 24.5080 48.3435 24.5340 49.4370 ;
        RECT 24.4000 48.3435 24.4260 49.4370 ;
        RECT 24.2920 48.3435 24.3180 49.4370 ;
        RECT 24.1840 48.3435 24.2100 49.4370 ;
        RECT 24.0760 48.3435 24.1020 49.4370 ;
        RECT 23.9680 48.3435 23.9940 49.4370 ;
        RECT 23.8600 48.3435 23.8860 49.4370 ;
        RECT 23.7520 48.3435 23.7780 49.4370 ;
        RECT 23.6440 48.3435 23.6700 49.4370 ;
        RECT 23.5360 48.3435 23.5620 49.4370 ;
        RECT 23.4280 48.3435 23.4540 49.4370 ;
        RECT 23.3200 48.3435 23.3460 49.4370 ;
        RECT 23.2120 48.3435 23.2380 49.4370 ;
        RECT 23.1040 48.3435 23.1300 49.4370 ;
        RECT 22.9960 48.3435 23.0220 49.4370 ;
        RECT 22.8880 48.3435 22.9140 49.4370 ;
        RECT 22.7800 48.3435 22.8060 49.4370 ;
        RECT 22.6720 48.3435 22.6980 49.4370 ;
        RECT 22.5640 48.3435 22.5900 49.4370 ;
        RECT 22.4560 48.3435 22.4820 49.4370 ;
        RECT 22.3480 48.3435 22.3740 49.4370 ;
        RECT 22.2400 48.3435 22.2660 49.4370 ;
        RECT 22.1320 48.3435 22.1580 49.4370 ;
        RECT 22.0240 48.3435 22.0500 49.4370 ;
        RECT 21.9160 48.3435 21.9420 49.4370 ;
        RECT 21.8080 48.3435 21.8340 49.4370 ;
        RECT 21.7000 48.3435 21.7260 49.4370 ;
        RECT 21.5920 48.3435 21.6180 49.4370 ;
        RECT 21.4840 48.3435 21.5100 49.4370 ;
        RECT 21.3760 48.3435 21.4020 49.4370 ;
        RECT 21.2680 48.3435 21.2940 49.4370 ;
        RECT 21.1600 48.3435 21.1860 49.4370 ;
        RECT 21.0520 48.3435 21.0780 49.4370 ;
        RECT 20.9440 48.3435 20.9700 49.4370 ;
        RECT 20.8360 48.3435 20.8620 49.4370 ;
        RECT 20.7280 48.3435 20.7540 49.4370 ;
        RECT 20.6200 48.3435 20.6460 49.4370 ;
        RECT 20.5120 48.3435 20.5380 49.4370 ;
        RECT 20.4040 48.3435 20.4300 49.4370 ;
        RECT 20.2960 48.3435 20.3220 49.4370 ;
        RECT 20.1880 48.3435 20.2140 49.4370 ;
        RECT 20.0800 48.3435 20.1060 49.4370 ;
        RECT 19.9720 48.3435 19.9980 49.4370 ;
        RECT 19.8640 48.3435 19.8900 49.4370 ;
        RECT 19.7560 48.3435 19.7820 49.4370 ;
        RECT 19.6480 48.3435 19.6740 49.4370 ;
        RECT 19.5400 48.3435 19.5660 49.4370 ;
        RECT 19.4320 48.3435 19.4580 49.4370 ;
        RECT 19.3240 48.3435 19.3500 49.4370 ;
        RECT 19.2160 48.3435 19.2420 49.4370 ;
        RECT 19.1080 48.3435 19.1340 49.4370 ;
        RECT 19.0000 48.3435 19.0260 49.4370 ;
        RECT 18.8920 48.3435 18.9180 49.4370 ;
        RECT 18.7840 48.3435 18.8100 49.4370 ;
        RECT 18.6760 48.3435 18.7020 49.4370 ;
        RECT 18.5680 48.3435 18.5940 49.4370 ;
        RECT 18.4600 48.3435 18.4860 49.4370 ;
        RECT 18.3520 48.3435 18.3780 49.4370 ;
        RECT 18.2440 48.3435 18.2700 49.4370 ;
        RECT 18.1360 48.3435 18.1620 49.4370 ;
        RECT 18.0280 48.3435 18.0540 49.4370 ;
        RECT 17.9200 48.3435 17.9460 49.4370 ;
        RECT 17.8120 48.3435 17.8380 49.4370 ;
        RECT 17.7040 48.3435 17.7300 49.4370 ;
        RECT 17.5960 48.3435 17.6220 49.4370 ;
        RECT 17.4880 48.3435 17.5140 49.4370 ;
        RECT 17.3800 48.3435 17.4060 49.4370 ;
        RECT 17.2720 48.3435 17.2980 49.4370 ;
        RECT 17.1640 48.3435 17.1900 49.4370 ;
        RECT 17.0560 48.3435 17.0820 49.4370 ;
        RECT 16.9480 48.3435 16.9740 49.4370 ;
        RECT 16.8400 48.3435 16.8660 49.4370 ;
        RECT 16.7320 48.3435 16.7580 49.4370 ;
        RECT 16.6240 48.3435 16.6500 49.4370 ;
        RECT 16.5160 48.3435 16.5420 49.4370 ;
        RECT 16.4080 48.3435 16.4340 49.4370 ;
        RECT 16.3000 48.3435 16.3260 49.4370 ;
        RECT 16.0870 48.3435 16.1640 49.4370 ;
        RECT 14.1940 48.3435 14.2710 49.4370 ;
        RECT 14.0320 48.3435 14.0580 49.4370 ;
        RECT 13.9240 48.3435 13.9500 49.4370 ;
        RECT 13.8160 48.3435 13.8420 49.4370 ;
        RECT 13.7080 48.3435 13.7340 49.4370 ;
        RECT 13.6000 48.3435 13.6260 49.4370 ;
        RECT 13.4920 48.3435 13.5180 49.4370 ;
        RECT 13.3840 48.3435 13.4100 49.4370 ;
        RECT 13.2760 48.3435 13.3020 49.4370 ;
        RECT 13.1680 48.3435 13.1940 49.4370 ;
        RECT 13.0600 48.3435 13.0860 49.4370 ;
        RECT 12.9520 48.3435 12.9780 49.4370 ;
        RECT 12.8440 48.3435 12.8700 49.4370 ;
        RECT 12.7360 48.3435 12.7620 49.4370 ;
        RECT 12.6280 48.3435 12.6540 49.4370 ;
        RECT 12.5200 48.3435 12.5460 49.4370 ;
        RECT 12.4120 48.3435 12.4380 49.4370 ;
        RECT 12.3040 48.3435 12.3300 49.4370 ;
        RECT 12.1960 48.3435 12.2220 49.4370 ;
        RECT 12.0880 48.3435 12.1140 49.4370 ;
        RECT 11.9800 48.3435 12.0060 49.4370 ;
        RECT 11.8720 48.3435 11.8980 49.4370 ;
        RECT 11.7640 48.3435 11.7900 49.4370 ;
        RECT 11.6560 48.3435 11.6820 49.4370 ;
        RECT 11.5480 48.3435 11.5740 49.4370 ;
        RECT 11.4400 48.3435 11.4660 49.4370 ;
        RECT 11.3320 48.3435 11.3580 49.4370 ;
        RECT 11.2240 48.3435 11.2500 49.4370 ;
        RECT 11.1160 48.3435 11.1420 49.4370 ;
        RECT 11.0080 48.3435 11.0340 49.4370 ;
        RECT 10.9000 48.3435 10.9260 49.4370 ;
        RECT 10.7920 48.3435 10.8180 49.4370 ;
        RECT 10.6840 48.3435 10.7100 49.4370 ;
        RECT 10.5760 48.3435 10.6020 49.4370 ;
        RECT 10.4680 48.3435 10.4940 49.4370 ;
        RECT 10.3600 48.3435 10.3860 49.4370 ;
        RECT 10.2520 48.3435 10.2780 49.4370 ;
        RECT 10.1440 48.3435 10.1700 49.4370 ;
        RECT 10.0360 48.3435 10.0620 49.4370 ;
        RECT 9.9280 48.3435 9.9540 49.4370 ;
        RECT 9.8200 48.3435 9.8460 49.4370 ;
        RECT 9.7120 48.3435 9.7380 49.4370 ;
        RECT 9.6040 48.3435 9.6300 49.4370 ;
        RECT 9.4960 48.3435 9.5220 49.4370 ;
        RECT 9.3880 48.3435 9.4140 49.4370 ;
        RECT 9.2800 48.3435 9.3060 49.4370 ;
        RECT 9.1720 48.3435 9.1980 49.4370 ;
        RECT 9.0640 48.3435 9.0900 49.4370 ;
        RECT 8.9560 48.3435 8.9820 49.4370 ;
        RECT 8.8480 48.3435 8.8740 49.4370 ;
        RECT 8.7400 48.3435 8.7660 49.4370 ;
        RECT 8.6320 48.3435 8.6580 49.4370 ;
        RECT 8.5240 48.3435 8.5500 49.4370 ;
        RECT 8.4160 48.3435 8.4420 49.4370 ;
        RECT 8.3080 48.3435 8.3340 49.4370 ;
        RECT 8.2000 48.3435 8.2260 49.4370 ;
        RECT 8.0920 48.3435 8.1180 49.4370 ;
        RECT 7.9840 48.3435 8.0100 49.4370 ;
        RECT 7.8760 48.3435 7.9020 49.4370 ;
        RECT 7.7680 48.3435 7.7940 49.4370 ;
        RECT 7.6600 48.3435 7.6860 49.4370 ;
        RECT 7.5520 48.3435 7.5780 49.4370 ;
        RECT 7.4440 48.3435 7.4700 49.4370 ;
        RECT 7.3360 48.3435 7.3620 49.4370 ;
        RECT 7.2280 48.3435 7.2540 49.4370 ;
        RECT 7.1200 48.3435 7.1460 49.4370 ;
        RECT 7.0120 48.3435 7.0380 49.4370 ;
        RECT 6.9040 48.3435 6.9300 49.4370 ;
        RECT 6.7960 48.3435 6.8220 49.4370 ;
        RECT 6.6880 48.3435 6.7140 49.4370 ;
        RECT 6.5800 48.3435 6.6060 49.4370 ;
        RECT 6.4720 48.3435 6.4980 49.4370 ;
        RECT 6.3640 48.3435 6.3900 49.4370 ;
        RECT 6.2560 48.3435 6.2820 49.4370 ;
        RECT 6.1480 48.3435 6.1740 49.4370 ;
        RECT 6.0400 48.3435 6.0660 49.4370 ;
        RECT 5.9320 48.3435 5.9580 49.4370 ;
        RECT 5.8240 48.3435 5.8500 49.4370 ;
        RECT 5.7160 48.3435 5.7420 49.4370 ;
        RECT 5.6080 48.3435 5.6340 49.4370 ;
        RECT 5.5000 48.3435 5.5260 49.4370 ;
        RECT 5.3920 48.3435 5.4180 49.4370 ;
        RECT 5.2840 48.3435 5.3100 49.4370 ;
        RECT 5.1760 48.3435 5.2020 49.4370 ;
        RECT 5.0680 48.3435 5.0940 49.4370 ;
        RECT 4.9600 48.3435 4.9860 49.4370 ;
        RECT 4.8520 48.3435 4.8780 49.4370 ;
        RECT 4.7440 48.3435 4.7700 49.4370 ;
        RECT 4.6360 48.3435 4.6620 49.4370 ;
        RECT 4.5280 48.3435 4.5540 49.4370 ;
        RECT 4.4200 48.3435 4.4460 49.4370 ;
        RECT 4.3120 48.3435 4.3380 49.4370 ;
        RECT 4.2040 48.3435 4.2300 49.4370 ;
        RECT 4.0960 48.3435 4.1220 49.4370 ;
        RECT 3.9880 48.3435 4.0140 49.4370 ;
        RECT 3.8800 48.3435 3.9060 49.4370 ;
        RECT 3.7720 48.3435 3.7980 49.4370 ;
        RECT 3.6640 48.3435 3.6900 49.4370 ;
        RECT 3.5560 48.3435 3.5820 49.4370 ;
        RECT 3.4480 48.3435 3.4740 49.4370 ;
        RECT 3.3400 48.3435 3.3660 49.4370 ;
        RECT 3.2320 48.3435 3.2580 49.4370 ;
        RECT 3.1240 48.3435 3.1500 49.4370 ;
        RECT 3.0160 48.3435 3.0420 49.4370 ;
        RECT 2.9080 48.3435 2.9340 49.4370 ;
        RECT 2.8000 48.3435 2.8260 49.4370 ;
        RECT 2.6920 48.3435 2.7180 49.4370 ;
        RECT 2.5840 48.3435 2.6100 49.4370 ;
        RECT 2.4760 48.3435 2.5020 49.4370 ;
        RECT 2.3680 48.3435 2.3940 49.4370 ;
        RECT 2.2600 48.3435 2.2860 49.4370 ;
        RECT 2.1520 48.3435 2.1780 49.4370 ;
        RECT 2.0440 48.3435 2.0700 49.4370 ;
        RECT 1.9360 48.3435 1.9620 49.4370 ;
        RECT 1.8280 48.3435 1.8540 49.4370 ;
        RECT 1.7200 48.3435 1.7460 49.4370 ;
        RECT 1.6120 48.3435 1.6380 49.4370 ;
        RECT 1.5040 48.3435 1.5300 49.4370 ;
        RECT 1.3960 48.3435 1.4220 49.4370 ;
        RECT 1.2880 48.3435 1.3140 49.4370 ;
        RECT 1.1800 48.3435 1.2060 49.4370 ;
        RECT 1.0720 48.3435 1.0980 49.4370 ;
        RECT 0.9640 48.3435 0.9900 49.4370 ;
        RECT 0.8560 48.3435 0.8820 49.4370 ;
        RECT 0.7480 48.3435 0.7740 49.4370 ;
        RECT 0.6400 48.3435 0.6660 49.4370 ;
        RECT 0.5320 48.3435 0.5580 49.4370 ;
        RECT 0.4240 48.3435 0.4500 49.4370 ;
        RECT 0.3160 48.3435 0.3420 49.4370 ;
        RECT 0.2080 48.3435 0.2340 49.4370 ;
        RECT 0.0050 48.3435 0.0900 49.4370 ;
        RECT 15.5530 49.4235 15.6810 50.5170 ;
        RECT 15.5390 50.0890 15.6810 50.4115 ;
        RECT 15.3190 49.8160 15.4530 50.5170 ;
        RECT 15.2960 50.1510 15.4530 50.4090 ;
        RECT 15.3190 49.4235 15.4170 50.5170 ;
        RECT 15.3190 49.5445 15.4310 49.7840 ;
        RECT 15.3190 49.4235 15.4530 49.5125 ;
        RECT 15.0940 49.8740 15.2280 50.5170 ;
        RECT 15.0940 49.4235 15.1920 50.5170 ;
        RECT 14.6770 49.4235 14.7600 50.5170 ;
        RECT 14.6770 49.5120 14.7740 50.4475 ;
        RECT 30.2680 49.4235 30.3530 50.5170 ;
        RECT 30.1240 49.4235 30.1500 50.5170 ;
        RECT 30.0160 49.4235 30.0420 50.5170 ;
        RECT 29.9080 49.4235 29.9340 50.5170 ;
        RECT 29.8000 49.4235 29.8260 50.5170 ;
        RECT 29.6920 49.4235 29.7180 50.5170 ;
        RECT 29.5840 49.4235 29.6100 50.5170 ;
        RECT 29.4760 49.4235 29.5020 50.5170 ;
        RECT 29.3680 49.4235 29.3940 50.5170 ;
        RECT 29.2600 49.4235 29.2860 50.5170 ;
        RECT 29.1520 49.4235 29.1780 50.5170 ;
        RECT 29.0440 49.4235 29.0700 50.5170 ;
        RECT 28.9360 49.4235 28.9620 50.5170 ;
        RECT 28.8280 49.4235 28.8540 50.5170 ;
        RECT 28.7200 49.4235 28.7460 50.5170 ;
        RECT 28.6120 49.4235 28.6380 50.5170 ;
        RECT 28.5040 49.4235 28.5300 50.5170 ;
        RECT 28.3960 49.4235 28.4220 50.5170 ;
        RECT 28.2880 49.4235 28.3140 50.5170 ;
        RECT 28.1800 49.4235 28.2060 50.5170 ;
        RECT 28.0720 49.4235 28.0980 50.5170 ;
        RECT 27.9640 49.4235 27.9900 50.5170 ;
        RECT 27.8560 49.4235 27.8820 50.5170 ;
        RECT 27.7480 49.4235 27.7740 50.5170 ;
        RECT 27.6400 49.4235 27.6660 50.5170 ;
        RECT 27.5320 49.4235 27.5580 50.5170 ;
        RECT 27.4240 49.4235 27.4500 50.5170 ;
        RECT 27.3160 49.4235 27.3420 50.5170 ;
        RECT 27.2080 49.4235 27.2340 50.5170 ;
        RECT 27.1000 49.4235 27.1260 50.5170 ;
        RECT 26.9920 49.4235 27.0180 50.5170 ;
        RECT 26.8840 49.4235 26.9100 50.5170 ;
        RECT 26.7760 49.4235 26.8020 50.5170 ;
        RECT 26.6680 49.4235 26.6940 50.5170 ;
        RECT 26.5600 49.4235 26.5860 50.5170 ;
        RECT 26.4520 49.4235 26.4780 50.5170 ;
        RECT 26.3440 49.4235 26.3700 50.5170 ;
        RECT 26.2360 49.4235 26.2620 50.5170 ;
        RECT 26.1280 49.4235 26.1540 50.5170 ;
        RECT 26.0200 49.4235 26.0460 50.5170 ;
        RECT 25.9120 49.4235 25.9380 50.5170 ;
        RECT 25.8040 49.4235 25.8300 50.5170 ;
        RECT 25.6960 49.4235 25.7220 50.5170 ;
        RECT 25.5880 49.4235 25.6140 50.5170 ;
        RECT 25.4800 49.4235 25.5060 50.5170 ;
        RECT 25.3720 49.4235 25.3980 50.5170 ;
        RECT 25.2640 49.4235 25.2900 50.5170 ;
        RECT 25.1560 49.4235 25.1820 50.5170 ;
        RECT 25.0480 49.4235 25.0740 50.5170 ;
        RECT 24.9400 49.4235 24.9660 50.5170 ;
        RECT 24.8320 49.4235 24.8580 50.5170 ;
        RECT 24.7240 49.4235 24.7500 50.5170 ;
        RECT 24.6160 49.4235 24.6420 50.5170 ;
        RECT 24.5080 49.4235 24.5340 50.5170 ;
        RECT 24.4000 49.4235 24.4260 50.5170 ;
        RECT 24.2920 49.4235 24.3180 50.5170 ;
        RECT 24.1840 49.4235 24.2100 50.5170 ;
        RECT 24.0760 49.4235 24.1020 50.5170 ;
        RECT 23.9680 49.4235 23.9940 50.5170 ;
        RECT 23.8600 49.4235 23.8860 50.5170 ;
        RECT 23.7520 49.4235 23.7780 50.5170 ;
        RECT 23.6440 49.4235 23.6700 50.5170 ;
        RECT 23.5360 49.4235 23.5620 50.5170 ;
        RECT 23.4280 49.4235 23.4540 50.5170 ;
        RECT 23.3200 49.4235 23.3460 50.5170 ;
        RECT 23.2120 49.4235 23.2380 50.5170 ;
        RECT 23.1040 49.4235 23.1300 50.5170 ;
        RECT 22.9960 49.4235 23.0220 50.5170 ;
        RECT 22.8880 49.4235 22.9140 50.5170 ;
        RECT 22.7800 49.4235 22.8060 50.5170 ;
        RECT 22.6720 49.4235 22.6980 50.5170 ;
        RECT 22.5640 49.4235 22.5900 50.5170 ;
        RECT 22.4560 49.4235 22.4820 50.5170 ;
        RECT 22.3480 49.4235 22.3740 50.5170 ;
        RECT 22.2400 49.4235 22.2660 50.5170 ;
        RECT 22.1320 49.4235 22.1580 50.5170 ;
        RECT 22.0240 49.4235 22.0500 50.5170 ;
        RECT 21.9160 49.4235 21.9420 50.5170 ;
        RECT 21.8080 49.4235 21.8340 50.5170 ;
        RECT 21.7000 49.4235 21.7260 50.5170 ;
        RECT 21.5920 49.4235 21.6180 50.5170 ;
        RECT 21.4840 49.4235 21.5100 50.5170 ;
        RECT 21.3760 49.4235 21.4020 50.5170 ;
        RECT 21.2680 49.4235 21.2940 50.5170 ;
        RECT 21.1600 49.4235 21.1860 50.5170 ;
        RECT 21.0520 49.4235 21.0780 50.5170 ;
        RECT 20.9440 49.4235 20.9700 50.5170 ;
        RECT 20.8360 49.4235 20.8620 50.5170 ;
        RECT 20.7280 49.4235 20.7540 50.5170 ;
        RECT 20.6200 49.4235 20.6460 50.5170 ;
        RECT 20.5120 49.4235 20.5380 50.5170 ;
        RECT 20.4040 49.4235 20.4300 50.5170 ;
        RECT 20.2960 49.4235 20.3220 50.5170 ;
        RECT 20.1880 49.4235 20.2140 50.5170 ;
        RECT 20.0800 49.4235 20.1060 50.5170 ;
        RECT 19.9720 49.4235 19.9980 50.5170 ;
        RECT 19.8640 49.4235 19.8900 50.5170 ;
        RECT 19.7560 49.4235 19.7820 50.5170 ;
        RECT 19.6480 49.4235 19.6740 50.5170 ;
        RECT 19.5400 49.4235 19.5660 50.5170 ;
        RECT 19.4320 49.4235 19.4580 50.5170 ;
        RECT 19.3240 49.4235 19.3500 50.5170 ;
        RECT 19.2160 49.4235 19.2420 50.5170 ;
        RECT 19.1080 49.4235 19.1340 50.5170 ;
        RECT 19.0000 49.4235 19.0260 50.5170 ;
        RECT 18.8920 49.4235 18.9180 50.5170 ;
        RECT 18.7840 49.4235 18.8100 50.5170 ;
        RECT 18.6760 49.4235 18.7020 50.5170 ;
        RECT 18.5680 49.4235 18.5940 50.5170 ;
        RECT 18.4600 49.4235 18.4860 50.5170 ;
        RECT 18.3520 49.4235 18.3780 50.5170 ;
        RECT 18.2440 49.4235 18.2700 50.5170 ;
        RECT 18.1360 49.4235 18.1620 50.5170 ;
        RECT 18.0280 49.4235 18.0540 50.5170 ;
        RECT 17.9200 49.4235 17.9460 50.5170 ;
        RECT 17.8120 49.4235 17.8380 50.5170 ;
        RECT 17.7040 49.4235 17.7300 50.5170 ;
        RECT 17.5960 49.4235 17.6220 50.5170 ;
        RECT 17.4880 49.4235 17.5140 50.5170 ;
        RECT 17.3800 49.4235 17.4060 50.5170 ;
        RECT 17.2720 49.4235 17.2980 50.5170 ;
        RECT 17.1640 49.4235 17.1900 50.5170 ;
        RECT 17.0560 49.4235 17.0820 50.5170 ;
        RECT 16.9480 49.4235 16.9740 50.5170 ;
        RECT 16.8400 49.4235 16.8660 50.5170 ;
        RECT 16.7320 49.4235 16.7580 50.5170 ;
        RECT 16.6240 49.4235 16.6500 50.5170 ;
        RECT 16.5160 49.4235 16.5420 50.5170 ;
        RECT 16.4080 49.4235 16.4340 50.5170 ;
        RECT 16.3000 49.4235 16.3260 50.5170 ;
        RECT 16.0870 49.4235 16.1640 50.5170 ;
        RECT 14.1940 49.4235 14.2710 50.5170 ;
        RECT 14.0320 49.4235 14.0580 50.5170 ;
        RECT 13.9240 49.4235 13.9500 50.5170 ;
        RECT 13.8160 49.4235 13.8420 50.5170 ;
        RECT 13.7080 49.4235 13.7340 50.5170 ;
        RECT 13.6000 49.4235 13.6260 50.5170 ;
        RECT 13.4920 49.4235 13.5180 50.5170 ;
        RECT 13.3840 49.4235 13.4100 50.5170 ;
        RECT 13.2760 49.4235 13.3020 50.5170 ;
        RECT 13.1680 49.4235 13.1940 50.5170 ;
        RECT 13.0600 49.4235 13.0860 50.5170 ;
        RECT 12.9520 49.4235 12.9780 50.5170 ;
        RECT 12.8440 49.4235 12.8700 50.5170 ;
        RECT 12.7360 49.4235 12.7620 50.5170 ;
        RECT 12.6280 49.4235 12.6540 50.5170 ;
        RECT 12.5200 49.4235 12.5460 50.5170 ;
        RECT 12.4120 49.4235 12.4380 50.5170 ;
        RECT 12.3040 49.4235 12.3300 50.5170 ;
        RECT 12.1960 49.4235 12.2220 50.5170 ;
        RECT 12.0880 49.4235 12.1140 50.5170 ;
        RECT 11.9800 49.4235 12.0060 50.5170 ;
        RECT 11.8720 49.4235 11.8980 50.5170 ;
        RECT 11.7640 49.4235 11.7900 50.5170 ;
        RECT 11.6560 49.4235 11.6820 50.5170 ;
        RECT 11.5480 49.4235 11.5740 50.5170 ;
        RECT 11.4400 49.4235 11.4660 50.5170 ;
        RECT 11.3320 49.4235 11.3580 50.5170 ;
        RECT 11.2240 49.4235 11.2500 50.5170 ;
        RECT 11.1160 49.4235 11.1420 50.5170 ;
        RECT 11.0080 49.4235 11.0340 50.5170 ;
        RECT 10.9000 49.4235 10.9260 50.5170 ;
        RECT 10.7920 49.4235 10.8180 50.5170 ;
        RECT 10.6840 49.4235 10.7100 50.5170 ;
        RECT 10.5760 49.4235 10.6020 50.5170 ;
        RECT 10.4680 49.4235 10.4940 50.5170 ;
        RECT 10.3600 49.4235 10.3860 50.5170 ;
        RECT 10.2520 49.4235 10.2780 50.5170 ;
        RECT 10.1440 49.4235 10.1700 50.5170 ;
        RECT 10.0360 49.4235 10.0620 50.5170 ;
        RECT 9.9280 49.4235 9.9540 50.5170 ;
        RECT 9.8200 49.4235 9.8460 50.5170 ;
        RECT 9.7120 49.4235 9.7380 50.5170 ;
        RECT 9.6040 49.4235 9.6300 50.5170 ;
        RECT 9.4960 49.4235 9.5220 50.5170 ;
        RECT 9.3880 49.4235 9.4140 50.5170 ;
        RECT 9.2800 49.4235 9.3060 50.5170 ;
        RECT 9.1720 49.4235 9.1980 50.5170 ;
        RECT 9.0640 49.4235 9.0900 50.5170 ;
        RECT 8.9560 49.4235 8.9820 50.5170 ;
        RECT 8.8480 49.4235 8.8740 50.5170 ;
        RECT 8.7400 49.4235 8.7660 50.5170 ;
        RECT 8.6320 49.4235 8.6580 50.5170 ;
        RECT 8.5240 49.4235 8.5500 50.5170 ;
        RECT 8.4160 49.4235 8.4420 50.5170 ;
        RECT 8.3080 49.4235 8.3340 50.5170 ;
        RECT 8.2000 49.4235 8.2260 50.5170 ;
        RECT 8.0920 49.4235 8.1180 50.5170 ;
        RECT 7.9840 49.4235 8.0100 50.5170 ;
        RECT 7.8760 49.4235 7.9020 50.5170 ;
        RECT 7.7680 49.4235 7.7940 50.5170 ;
        RECT 7.6600 49.4235 7.6860 50.5170 ;
        RECT 7.5520 49.4235 7.5780 50.5170 ;
        RECT 7.4440 49.4235 7.4700 50.5170 ;
        RECT 7.3360 49.4235 7.3620 50.5170 ;
        RECT 7.2280 49.4235 7.2540 50.5170 ;
        RECT 7.1200 49.4235 7.1460 50.5170 ;
        RECT 7.0120 49.4235 7.0380 50.5170 ;
        RECT 6.9040 49.4235 6.9300 50.5170 ;
        RECT 6.7960 49.4235 6.8220 50.5170 ;
        RECT 6.6880 49.4235 6.7140 50.5170 ;
        RECT 6.5800 49.4235 6.6060 50.5170 ;
        RECT 6.4720 49.4235 6.4980 50.5170 ;
        RECT 6.3640 49.4235 6.3900 50.5170 ;
        RECT 6.2560 49.4235 6.2820 50.5170 ;
        RECT 6.1480 49.4235 6.1740 50.5170 ;
        RECT 6.0400 49.4235 6.0660 50.5170 ;
        RECT 5.9320 49.4235 5.9580 50.5170 ;
        RECT 5.8240 49.4235 5.8500 50.5170 ;
        RECT 5.7160 49.4235 5.7420 50.5170 ;
        RECT 5.6080 49.4235 5.6340 50.5170 ;
        RECT 5.5000 49.4235 5.5260 50.5170 ;
        RECT 5.3920 49.4235 5.4180 50.5170 ;
        RECT 5.2840 49.4235 5.3100 50.5170 ;
        RECT 5.1760 49.4235 5.2020 50.5170 ;
        RECT 5.0680 49.4235 5.0940 50.5170 ;
        RECT 4.9600 49.4235 4.9860 50.5170 ;
        RECT 4.8520 49.4235 4.8780 50.5170 ;
        RECT 4.7440 49.4235 4.7700 50.5170 ;
        RECT 4.6360 49.4235 4.6620 50.5170 ;
        RECT 4.5280 49.4235 4.5540 50.5170 ;
        RECT 4.4200 49.4235 4.4460 50.5170 ;
        RECT 4.3120 49.4235 4.3380 50.5170 ;
        RECT 4.2040 49.4235 4.2300 50.5170 ;
        RECT 4.0960 49.4235 4.1220 50.5170 ;
        RECT 3.9880 49.4235 4.0140 50.5170 ;
        RECT 3.8800 49.4235 3.9060 50.5170 ;
        RECT 3.7720 49.4235 3.7980 50.5170 ;
        RECT 3.6640 49.4235 3.6900 50.5170 ;
        RECT 3.5560 49.4235 3.5820 50.5170 ;
        RECT 3.4480 49.4235 3.4740 50.5170 ;
        RECT 3.3400 49.4235 3.3660 50.5170 ;
        RECT 3.2320 49.4235 3.2580 50.5170 ;
        RECT 3.1240 49.4235 3.1500 50.5170 ;
        RECT 3.0160 49.4235 3.0420 50.5170 ;
        RECT 2.9080 49.4235 2.9340 50.5170 ;
        RECT 2.8000 49.4235 2.8260 50.5170 ;
        RECT 2.6920 49.4235 2.7180 50.5170 ;
        RECT 2.5840 49.4235 2.6100 50.5170 ;
        RECT 2.4760 49.4235 2.5020 50.5170 ;
        RECT 2.3680 49.4235 2.3940 50.5170 ;
        RECT 2.2600 49.4235 2.2860 50.5170 ;
        RECT 2.1520 49.4235 2.1780 50.5170 ;
        RECT 2.0440 49.4235 2.0700 50.5170 ;
        RECT 1.9360 49.4235 1.9620 50.5170 ;
        RECT 1.8280 49.4235 1.8540 50.5170 ;
        RECT 1.7200 49.4235 1.7460 50.5170 ;
        RECT 1.6120 49.4235 1.6380 50.5170 ;
        RECT 1.5040 49.4235 1.5300 50.5170 ;
        RECT 1.3960 49.4235 1.4220 50.5170 ;
        RECT 1.2880 49.4235 1.3140 50.5170 ;
        RECT 1.1800 49.4235 1.2060 50.5170 ;
        RECT 1.0720 49.4235 1.0980 50.5170 ;
        RECT 0.9640 49.4235 0.9900 50.5170 ;
        RECT 0.8560 49.4235 0.8820 50.5170 ;
        RECT 0.7480 49.4235 0.7740 50.5170 ;
        RECT 0.6400 49.4235 0.6660 50.5170 ;
        RECT 0.5320 49.4235 0.5580 50.5170 ;
        RECT 0.4240 49.4235 0.4500 50.5170 ;
        RECT 0.3160 49.4235 0.3420 50.5170 ;
        RECT 0.2080 49.4235 0.2340 50.5170 ;
        RECT 0.0050 49.4235 0.0900 50.5170 ;
        RECT 15.5530 50.5035 15.6810 51.5970 ;
        RECT 15.5390 51.1690 15.6810 51.4915 ;
        RECT 15.3190 50.8960 15.4530 51.5970 ;
        RECT 15.2960 51.2310 15.4530 51.4890 ;
        RECT 15.3190 50.5035 15.4170 51.5970 ;
        RECT 15.3190 50.6245 15.4310 50.8640 ;
        RECT 15.3190 50.5035 15.4530 50.5925 ;
        RECT 15.0940 50.9540 15.2280 51.5970 ;
        RECT 15.0940 50.5035 15.1920 51.5970 ;
        RECT 14.6770 50.5035 14.7600 51.5970 ;
        RECT 14.6770 50.5920 14.7740 51.5275 ;
        RECT 30.2680 50.5035 30.3530 51.5970 ;
        RECT 30.1240 50.5035 30.1500 51.5970 ;
        RECT 30.0160 50.5035 30.0420 51.5970 ;
        RECT 29.9080 50.5035 29.9340 51.5970 ;
        RECT 29.8000 50.5035 29.8260 51.5970 ;
        RECT 29.6920 50.5035 29.7180 51.5970 ;
        RECT 29.5840 50.5035 29.6100 51.5970 ;
        RECT 29.4760 50.5035 29.5020 51.5970 ;
        RECT 29.3680 50.5035 29.3940 51.5970 ;
        RECT 29.2600 50.5035 29.2860 51.5970 ;
        RECT 29.1520 50.5035 29.1780 51.5970 ;
        RECT 29.0440 50.5035 29.0700 51.5970 ;
        RECT 28.9360 50.5035 28.9620 51.5970 ;
        RECT 28.8280 50.5035 28.8540 51.5970 ;
        RECT 28.7200 50.5035 28.7460 51.5970 ;
        RECT 28.6120 50.5035 28.6380 51.5970 ;
        RECT 28.5040 50.5035 28.5300 51.5970 ;
        RECT 28.3960 50.5035 28.4220 51.5970 ;
        RECT 28.2880 50.5035 28.3140 51.5970 ;
        RECT 28.1800 50.5035 28.2060 51.5970 ;
        RECT 28.0720 50.5035 28.0980 51.5970 ;
        RECT 27.9640 50.5035 27.9900 51.5970 ;
        RECT 27.8560 50.5035 27.8820 51.5970 ;
        RECT 27.7480 50.5035 27.7740 51.5970 ;
        RECT 27.6400 50.5035 27.6660 51.5970 ;
        RECT 27.5320 50.5035 27.5580 51.5970 ;
        RECT 27.4240 50.5035 27.4500 51.5970 ;
        RECT 27.3160 50.5035 27.3420 51.5970 ;
        RECT 27.2080 50.5035 27.2340 51.5970 ;
        RECT 27.1000 50.5035 27.1260 51.5970 ;
        RECT 26.9920 50.5035 27.0180 51.5970 ;
        RECT 26.8840 50.5035 26.9100 51.5970 ;
        RECT 26.7760 50.5035 26.8020 51.5970 ;
        RECT 26.6680 50.5035 26.6940 51.5970 ;
        RECT 26.5600 50.5035 26.5860 51.5970 ;
        RECT 26.4520 50.5035 26.4780 51.5970 ;
        RECT 26.3440 50.5035 26.3700 51.5970 ;
        RECT 26.2360 50.5035 26.2620 51.5970 ;
        RECT 26.1280 50.5035 26.1540 51.5970 ;
        RECT 26.0200 50.5035 26.0460 51.5970 ;
        RECT 25.9120 50.5035 25.9380 51.5970 ;
        RECT 25.8040 50.5035 25.8300 51.5970 ;
        RECT 25.6960 50.5035 25.7220 51.5970 ;
        RECT 25.5880 50.5035 25.6140 51.5970 ;
        RECT 25.4800 50.5035 25.5060 51.5970 ;
        RECT 25.3720 50.5035 25.3980 51.5970 ;
        RECT 25.2640 50.5035 25.2900 51.5970 ;
        RECT 25.1560 50.5035 25.1820 51.5970 ;
        RECT 25.0480 50.5035 25.0740 51.5970 ;
        RECT 24.9400 50.5035 24.9660 51.5970 ;
        RECT 24.8320 50.5035 24.8580 51.5970 ;
        RECT 24.7240 50.5035 24.7500 51.5970 ;
        RECT 24.6160 50.5035 24.6420 51.5970 ;
        RECT 24.5080 50.5035 24.5340 51.5970 ;
        RECT 24.4000 50.5035 24.4260 51.5970 ;
        RECT 24.2920 50.5035 24.3180 51.5970 ;
        RECT 24.1840 50.5035 24.2100 51.5970 ;
        RECT 24.0760 50.5035 24.1020 51.5970 ;
        RECT 23.9680 50.5035 23.9940 51.5970 ;
        RECT 23.8600 50.5035 23.8860 51.5970 ;
        RECT 23.7520 50.5035 23.7780 51.5970 ;
        RECT 23.6440 50.5035 23.6700 51.5970 ;
        RECT 23.5360 50.5035 23.5620 51.5970 ;
        RECT 23.4280 50.5035 23.4540 51.5970 ;
        RECT 23.3200 50.5035 23.3460 51.5970 ;
        RECT 23.2120 50.5035 23.2380 51.5970 ;
        RECT 23.1040 50.5035 23.1300 51.5970 ;
        RECT 22.9960 50.5035 23.0220 51.5970 ;
        RECT 22.8880 50.5035 22.9140 51.5970 ;
        RECT 22.7800 50.5035 22.8060 51.5970 ;
        RECT 22.6720 50.5035 22.6980 51.5970 ;
        RECT 22.5640 50.5035 22.5900 51.5970 ;
        RECT 22.4560 50.5035 22.4820 51.5970 ;
        RECT 22.3480 50.5035 22.3740 51.5970 ;
        RECT 22.2400 50.5035 22.2660 51.5970 ;
        RECT 22.1320 50.5035 22.1580 51.5970 ;
        RECT 22.0240 50.5035 22.0500 51.5970 ;
        RECT 21.9160 50.5035 21.9420 51.5970 ;
        RECT 21.8080 50.5035 21.8340 51.5970 ;
        RECT 21.7000 50.5035 21.7260 51.5970 ;
        RECT 21.5920 50.5035 21.6180 51.5970 ;
        RECT 21.4840 50.5035 21.5100 51.5970 ;
        RECT 21.3760 50.5035 21.4020 51.5970 ;
        RECT 21.2680 50.5035 21.2940 51.5970 ;
        RECT 21.1600 50.5035 21.1860 51.5970 ;
        RECT 21.0520 50.5035 21.0780 51.5970 ;
        RECT 20.9440 50.5035 20.9700 51.5970 ;
        RECT 20.8360 50.5035 20.8620 51.5970 ;
        RECT 20.7280 50.5035 20.7540 51.5970 ;
        RECT 20.6200 50.5035 20.6460 51.5970 ;
        RECT 20.5120 50.5035 20.5380 51.5970 ;
        RECT 20.4040 50.5035 20.4300 51.5970 ;
        RECT 20.2960 50.5035 20.3220 51.5970 ;
        RECT 20.1880 50.5035 20.2140 51.5970 ;
        RECT 20.0800 50.5035 20.1060 51.5970 ;
        RECT 19.9720 50.5035 19.9980 51.5970 ;
        RECT 19.8640 50.5035 19.8900 51.5970 ;
        RECT 19.7560 50.5035 19.7820 51.5970 ;
        RECT 19.6480 50.5035 19.6740 51.5970 ;
        RECT 19.5400 50.5035 19.5660 51.5970 ;
        RECT 19.4320 50.5035 19.4580 51.5970 ;
        RECT 19.3240 50.5035 19.3500 51.5970 ;
        RECT 19.2160 50.5035 19.2420 51.5970 ;
        RECT 19.1080 50.5035 19.1340 51.5970 ;
        RECT 19.0000 50.5035 19.0260 51.5970 ;
        RECT 18.8920 50.5035 18.9180 51.5970 ;
        RECT 18.7840 50.5035 18.8100 51.5970 ;
        RECT 18.6760 50.5035 18.7020 51.5970 ;
        RECT 18.5680 50.5035 18.5940 51.5970 ;
        RECT 18.4600 50.5035 18.4860 51.5970 ;
        RECT 18.3520 50.5035 18.3780 51.5970 ;
        RECT 18.2440 50.5035 18.2700 51.5970 ;
        RECT 18.1360 50.5035 18.1620 51.5970 ;
        RECT 18.0280 50.5035 18.0540 51.5970 ;
        RECT 17.9200 50.5035 17.9460 51.5970 ;
        RECT 17.8120 50.5035 17.8380 51.5970 ;
        RECT 17.7040 50.5035 17.7300 51.5970 ;
        RECT 17.5960 50.5035 17.6220 51.5970 ;
        RECT 17.4880 50.5035 17.5140 51.5970 ;
        RECT 17.3800 50.5035 17.4060 51.5970 ;
        RECT 17.2720 50.5035 17.2980 51.5970 ;
        RECT 17.1640 50.5035 17.1900 51.5970 ;
        RECT 17.0560 50.5035 17.0820 51.5970 ;
        RECT 16.9480 50.5035 16.9740 51.5970 ;
        RECT 16.8400 50.5035 16.8660 51.5970 ;
        RECT 16.7320 50.5035 16.7580 51.5970 ;
        RECT 16.6240 50.5035 16.6500 51.5970 ;
        RECT 16.5160 50.5035 16.5420 51.5970 ;
        RECT 16.4080 50.5035 16.4340 51.5970 ;
        RECT 16.3000 50.5035 16.3260 51.5970 ;
        RECT 16.0870 50.5035 16.1640 51.5970 ;
        RECT 14.1940 50.5035 14.2710 51.5970 ;
        RECT 14.0320 50.5035 14.0580 51.5970 ;
        RECT 13.9240 50.5035 13.9500 51.5970 ;
        RECT 13.8160 50.5035 13.8420 51.5970 ;
        RECT 13.7080 50.5035 13.7340 51.5970 ;
        RECT 13.6000 50.5035 13.6260 51.5970 ;
        RECT 13.4920 50.5035 13.5180 51.5970 ;
        RECT 13.3840 50.5035 13.4100 51.5970 ;
        RECT 13.2760 50.5035 13.3020 51.5970 ;
        RECT 13.1680 50.5035 13.1940 51.5970 ;
        RECT 13.0600 50.5035 13.0860 51.5970 ;
        RECT 12.9520 50.5035 12.9780 51.5970 ;
        RECT 12.8440 50.5035 12.8700 51.5970 ;
        RECT 12.7360 50.5035 12.7620 51.5970 ;
        RECT 12.6280 50.5035 12.6540 51.5970 ;
        RECT 12.5200 50.5035 12.5460 51.5970 ;
        RECT 12.4120 50.5035 12.4380 51.5970 ;
        RECT 12.3040 50.5035 12.3300 51.5970 ;
        RECT 12.1960 50.5035 12.2220 51.5970 ;
        RECT 12.0880 50.5035 12.1140 51.5970 ;
        RECT 11.9800 50.5035 12.0060 51.5970 ;
        RECT 11.8720 50.5035 11.8980 51.5970 ;
        RECT 11.7640 50.5035 11.7900 51.5970 ;
        RECT 11.6560 50.5035 11.6820 51.5970 ;
        RECT 11.5480 50.5035 11.5740 51.5970 ;
        RECT 11.4400 50.5035 11.4660 51.5970 ;
        RECT 11.3320 50.5035 11.3580 51.5970 ;
        RECT 11.2240 50.5035 11.2500 51.5970 ;
        RECT 11.1160 50.5035 11.1420 51.5970 ;
        RECT 11.0080 50.5035 11.0340 51.5970 ;
        RECT 10.9000 50.5035 10.9260 51.5970 ;
        RECT 10.7920 50.5035 10.8180 51.5970 ;
        RECT 10.6840 50.5035 10.7100 51.5970 ;
        RECT 10.5760 50.5035 10.6020 51.5970 ;
        RECT 10.4680 50.5035 10.4940 51.5970 ;
        RECT 10.3600 50.5035 10.3860 51.5970 ;
        RECT 10.2520 50.5035 10.2780 51.5970 ;
        RECT 10.1440 50.5035 10.1700 51.5970 ;
        RECT 10.0360 50.5035 10.0620 51.5970 ;
        RECT 9.9280 50.5035 9.9540 51.5970 ;
        RECT 9.8200 50.5035 9.8460 51.5970 ;
        RECT 9.7120 50.5035 9.7380 51.5970 ;
        RECT 9.6040 50.5035 9.6300 51.5970 ;
        RECT 9.4960 50.5035 9.5220 51.5970 ;
        RECT 9.3880 50.5035 9.4140 51.5970 ;
        RECT 9.2800 50.5035 9.3060 51.5970 ;
        RECT 9.1720 50.5035 9.1980 51.5970 ;
        RECT 9.0640 50.5035 9.0900 51.5970 ;
        RECT 8.9560 50.5035 8.9820 51.5970 ;
        RECT 8.8480 50.5035 8.8740 51.5970 ;
        RECT 8.7400 50.5035 8.7660 51.5970 ;
        RECT 8.6320 50.5035 8.6580 51.5970 ;
        RECT 8.5240 50.5035 8.5500 51.5970 ;
        RECT 8.4160 50.5035 8.4420 51.5970 ;
        RECT 8.3080 50.5035 8.3340 51.5970 ;
        RECT 8.2000 50.5035 8.2260 51.5970 ;
        RECT 8.0920 50.5035 8.1180 51.5970 ;
        RECT 7.9840 50.5035 8.0100 51.5970 ;
        RECT 7.8760 50.5035 7.9020 51.5970 ;
        RECT 7.7680 50.5035 7.7940 51.5970 ;
        RECT 7.6600 50.5035 7.6860 51.5970 ;
        RECT 7.5520 50.5035 7.5780 51.5970 ;
        RECT 7.4440 50.5035 7.4700 51.5970 ;
        RECT 7.3360 50.5035 7.3620 51.5970 ;
        RECT 7.2280 50.5035 7.2540 51.5970 ;
        RECT 7.1200 50.5035 7.1460 51.5970 ;
        RECT 7.0120 50.5035 7.0380 51.5970 ;
        RECT 6.9040 50.5035 6.9300 51.5970 ;
        RECT 6.7960 50.5035 6.8220 51.5970 ;
        RECT 6.6880 50.5035 6.7140 51.5970 ;
        RECT 6.5800 50.5035 6.6060 51.5970 ;
        RECT 6.4720 50.5035 6.4980 51.5970 ;
        RECT 6.3640 50.5035 6.3900 51.5970 ;
        RECT 6.2560 50.5035 6.2820 51.5970 ;
        RECT 6.1480 50.5035 6.1740 51.5970 ;
        RECT 6.0400 50.5035 6.0660 51.5970 ;
        RECT 5.9320 50.5035 5.9580 51.5970 ;
        RECT 5.8240 50.5035 5.8500 51.5970 ;
        RECT 5.7160 50.5035 5.7420 51.5970 ;
        RECT 5.6080 50.5035 5.6340 51.5970 ;
        RECT 5.5000 50.5035 5.5260 51.5970 ;
        RECT 5.3920 50.5035 5.4180 51.5970 ;
        RECT 5.2840 50.5035 5.3100 51.5970 ;
        RECT 5.1760 50.5035 5.2020 51.5970 ;
        RECT 5.0680 50.5035 5.0940 51.5970 ;
        RECT 4.9600 50.5035 4.9860 51.5970 ;
        RECT 4.8520 50.5035 4.8780 51.5970 ;
        RECT 4.7440 50.5035 4.7700 51.5970 ;
        RECT 4.6360 50.5035 4.6620 51.5970 ;
        RECT 4.5280 50.5035 4.5540 51.5970 ;
        RECT 4.4200 50.5035 4.4460 51.5970 ;
        RECT 4.3120 50.5035 4.3380 51.5970 ;
        RECT 4.2040 50.5035 4.2300 51.5970 ;
        RECT 4.0960 50.5035 4.1220 51.5970 ;
        RECT 3.9880 50.5035 4.0140 51.5970 ;
        RECT 3.8800 50.5035 3.9060 51.5970 ;
        RECT 3.7720 50.5035 3.7980 51.5970 ;
        RECT 3.6640 50.5035 3.6900 51.5970 ;
        RECT 3.5560 50.5035 3.5820 51.5970 ;
        RECT 3.4480 50.5035 3.4740 51.5970 ;
        RECT 3.3400 50.5035 3.3660 51.5970 ;
        RECT 3.2320 50.5035 3.2580 51.5970 ;
        RECT 3.1240 50.5035 3.1500 51.5970 ;
        RECT 3.0160 50.5035 3.0420 51.5970 ;
        RECT 2.9080 50.5035 2.9340 51.5970 ;
        RECT 2.8000 50.5035 2.8260 51.5970 ;
        RECT 2.6920 50.5035 2.7180 51.5970 ;
        RECT 2.5840 50.5035 2.6100 51.5970 ;
        RECT 2.4760 50.5035 2.5020 51.5970 ;
        RECT 2.3680 50.5035 2.3940 51.5970 ;
        RECT 2.2600 50.5035 2.2860 51.5970 ;
        RECT 2.1520 50.5035 2.1780 51.5970 ;
        RECT 2.0440 50.5035 2.0700 51.5970 ;
        RECT 1.9360 50.5035 1.9620 51.5970 ;
        RECT 1.8280 50.5035 1.8540 51.5970 ;
        RECT 1.7200 50.5035 1.7460 51.5970 ;
        RECT 1.6120 50.5035 1.6380 51.5970 ;
        RECT 1.5040 50.5035 1.5300 51.5970 ;
        RECT 1.3960 50.5035 1.4220 51.5970 ;
        RECT 1.2880 50.5035 1.3140 51.5970 ;
        RECT 1.1800 50.5035 1.2060 51.5970 ;
        RECT 1.0720 50.5035 1.0980 51.5970 ;
        RECT 0.9640 50.5035 0.9900 51.5970 ;
        RECT 0.8560 50.5035 0.8820 51.5970 ;
        RECT 0.7480 50.5035 0.7740 51.5970 ;
        RECT 0.6400 50.5035 0.6660 51.5970 ;
        RECT 0.5320 50.5035 0.5580 51.5970 ;
        RECT 0.4240 50.5035 0.4500 51.5970 ;
        RECT 0.3160 50.5035 0.3420 51.5970 ;
        RECT 0.2080 50.5035 0.2340 51.5970 ;
        RECT 0.0050 50.5035 0.0900 51.5970 ;
        RECT 15.5530 51.5835 15.6810 52.6770 ;
        RECT 15.5390 52.2490 15.6810 52.5715 ;
        RECT 15.3190 51.9760 15.4530 52.6770 ;
        RECT 15.2960 52.3110 15.4530 52.5690 ;
        RECT 15.3190 51.5835 15.4170 52.6770 ;
        RECT 15.3190 51.7045 15.4310 51.9440 ;
        RECT 15.3190 51.5835 15.4530 51.6725 ;
        RECT 15.0940 52.0340 15.2280 52.6770 ;
        RECT 15.0940 51.5835 15.1920 52.6770 ;
        RECT 14.6770 51.5835 14.7600 52.6770 ;
        RECT 14.6770 51.6720 14.7740 52.6075 ;
        RECT 30.2680 51.5835 30.3530 52.6770 ;
        RECT 30.1240 51.5835 30.1500 52.6770 ;
        RECT 30.0160 51.5835 30.0420 52.6770 ;
        RECT 29.9080 51.5835 29.9340 52.6770 ;
        RECT 29.8000 51.5835 29.8260 52.6770 ;
        RECT 29.6920 51.5835 29.7180 52.6770 ;
        RECT 29.5840 51.5835 29.6100 52.6770 ;
        RECT 29.4760 51.5835 29.5020 52.6770 ;
        RECT 29.3680 51.5835 29.3940 52.6770 ;
        RECT 29.2600 51.5835 29.2860 52.6770 ;
        RECT 29.1520 51.5835 29.1780 52.6770 ;
        RECT 29.0440 51.5835 29.0700 52.6770 ;
        RECT 28.9360 51.5835 28.9620 52.6770 ;
        RECT 28.8280 51.5835 28.8540 52.6770 ;
        RECT 28.7200 51.5835 28.7460 52.6770 ;
        RECT 28.6120 51.5835 28.6380 52.6770 ;
        RECT 28.5040 51.5835 28.5300 52.6770 ;
        RECT 28.3960 51.5835 28.4220 52.6770 ;
        RECT 28.2880 51.5835 28.3140 52.6770 ;
        RECT 28.1800 51.5835 28.2060 52.6770 ;
        RECT 28.0720 51.5835 28.0980 52.6770 ;
        RECT 27.9640 51.5835 27.9900 52.6770 ;
        RECT 27.8560 51.5835 27.8820 52.6770 ;
        RECT 27.7480 51.5835 27.7740 52.6770 ;
        RECT 27.6400 51.5835 27.6660 52.6770 ;
        RECT 27.5320 51.5835 27.5580 52.6770 ;
        RECT 27.4240 51.5835 27.4500 52.6770 ;
        RECT 27.3160 51.5835 27.3420 52.6770 ;
        RECT 27.2080 51.5835 27.2340 52.6770 ;
        RECT 27.1000 51.5835 27.1260 52.6770 ;
        RECT 26.9920 51.5835 27.0180 52.6770 ;
        RECT 26.8840 51.5835 26.9100 52.6770 ;
        RECT 26.7760 51.5835 26.8020 52.6770 ;
        RECT 26.6680 51.5835 26.6940 52.6770 ;
        RECT 26.5600 51.5835 26.5860 52.6770 ;
        RECT 26.4520 51.5835 26.4780 52.6770 ;
        RECT 26.3440 51.5835 26.3700 52.6770 ;
        RECT 26.2360 51.5835 26.2620 52.6770 ;
        RECT 26.1280 51.5835 26.1540 52.6770 ;
        RECT 26.0200 51.5835 26.0460 52.6770 ;
        RECT 25.9120 51.5835 25.9380 52.6770 ;
        RECT 25.8040 51.5835 25.8300 52.6770 ;
        RECT 25.6960 51.5835 25.7220 52.6770 ;
        RECT 25.5880 51.5835 25.6140 52.6770 ;
        RECT 25.4800 51.5835 25.5060 52.6770 ;
        RECT 25.3720 51.5835 25.3980 52.6770 ;
        RECT 25.2640 51.5835 25.2900 52.6770 ;
        RECT 25.1560 51.5835 25.1820 52.6770 ;
        RECT 25.0480 51.5835 25.0740 52.6770 ;
        RECT 24.9400 51.5835 24.9660 52.6770 ;
        RECT 24.8320 51.5835 24.8580 52.6770 ;
        RECT 24.7240 51.5835 24.7500 52.6770 ;
        RECT 24.6160 51.5835 24.6420 52.6770 ;
        RECT 24.5080 51.5835 24.5340 52.6770 ;
        RECT 24.4000 51.5835 24.4260 52.6770 ;
        RECT 24.2920 51.5835 24.3180 52.6770 ;
        RECT 24.1840 51.5835 24.2100 52.6770 ;
        RECT 24.0760 51.5835 24.1020 52.6770 ;
        RECT 23.9680 51.5835 23.9940 52.6770 ;
        RECT 23.8600 51.5835 23.8860 52.6770 ;
        RECT 23.7520 51.5835 23.7780 52.6770 ;
        RECT 23.6440 51.5835 23.6700 52.6770 ;
        RECT 23.5360 51.5835 23.5620 52.6770 ;
        RECT 23.4280 51.5835 23.4540 52.6770 ;
        RECT 23.3200 51.5835 23.3460 52.6770 ;
        RECT 23.2120 51.5835 23.2380 52.6770 ;
        RECT 23.1040 51.5835 23.1300 52.6770 ;
        RECT 22.9960 51.5835 23.0220 52.6770 ;
        RECT 22.8880 51.5835 22.9140 52.6770 ;
        RECT 22.7800 51.5835 22.8060 52.6770 ;
        RECT 22.6720 51.5835 22.6980 52.6770 ;
        RECT 22.5640 51.5835 22.5900 52.6770 ;
        RECT 22.4560 51.5835 22.4820 52.6770 ;
        RECT 22.3480 51.5835 22.3740 52.6770 ;
        RECT 22.2400 51.5835 22.2660 52.6770 ;
        RECT 22.1320 51.5835 22.1580 52.6770 ;
        RECT 22.0240 51.5835 22.0500 52.6770 ;
        RECT 21.9160 51.5835 21.9420 52.6770 ;
        RECT 21.8080 51.5835 21.8340 52.6770 ;
        RECT 21.7000 51.5835 21.7260 52.6770 ;
        RECT 21.5920 51.5835 21.6180 52.6770 ;
        RECT 21.4840 51.5835 21.5100 52.6770 ;
        RECT 21.3760 51.5835 21.4020 52.6770 ;
        RECT 21.2680 51.5835 21.2940 52.6770 ;
        RECT 21.1600 51.5835 21.1860 52.6770 ;
        RECT 21.0520 51.5835 21.0780 52.6770 ;
        RECT 20.9440 51.5835 20.9700 52.6770 ;
        RECT 20.8360 51.5835 20.8620 52.6770 ;
        RECT 20.7280 51.5835 20.7540 52.6770 ;
        RECT 20.6200 51.5835 20.6460 52.6770 ;
        RECT 20.5120 51.5835 20.5380 52.6770 ;
        RECT 20.4040 51.5835 20.4300 52.6770 ;
        RECT 20.2960 51.5835 20.3220 52.6770 ;
        RECT 20.1880 51.5835 20.2140 52.6770 ;
        RECT 20.0800 51.5835 20.1060 52.6770 ;
        RECT 19.9720 51.5835 19.9980 52.6770 ;
        RECT 19.8640 51.5835 19.8900 52.6770 ;
        RECT 19.7560 51.5835 19.7820 52.6770 ;
        RECT 19.6480 51.5835 19.6740 52.6770 ;
        RECT 19.5400 51.5835 19.5660 52.6770 ;
        RECT 19.4320 51.5835 19.4580 52.6770 ;
        RECT 19.3240 51.5835 19.3500 52.6770 ;
        RECT 19.2160 51.5835 19.2420 52.6770 ;
        RECT 19.1080 51.5835 19.1340 52.6770 ;
        RECT 19.0000 51.5835 19.0260 52.6770 ;
        RECT 18.8920 51.5835 18.9180 52.6770 ;
        RECT 18.7840 51.5835 18.8100 52.6770 ;
        RECT 18.6760 51.5835 18.7020 52.6770 ;
        RECT 18.5680 51.5835 18.5940 52.6770 ;
        RECT 18.4600 51.5835 18.4860 52.6770 ;
        RECT 18.3520 51.5835 18.3780 52.6770 ;
        RECT 18.2440 51.5835 18.2700 52.6770 ;
        RECT 18.1360 51.5835 18.1620 52.6770 ;
        RECT 18.0280 51.5835 18.0540 52.6770 ;
        RECT 17.9200 51.5835 17.9460 52.6770 ;
        RECT 17.8120 51.5835 17.8380 52.6770 ;
        RECT 17.7040 51.5835 17.7300 52.6770 ;
        RECT 17.5960 51.5835 17.6220 52.6770 ;
        RECT 17.4880 51.5835 17.5140 52.6770 ;
        RECT 17.3800 51.5835 17.4060 52.6770 ;
        RECT 17.2720 51.5835 17.2980 52.6770 ;
        RECT 17.1640 51.5835 17.1900 52.6770 ;
        RECT 17.0560 51.5835 17.0820 52.6770 ;
        RECT 16.9480 51.5835 16.9740 52.6770 ;
        RECT 16.8400 51.5835 16.8660 52.6770 ;
        RECT 16.7320 51.5835 16.7580 52.6770 ;
        RECT 16.6240 51.5835 16.6500 52.6770 ;
        RECT 16.5160 51.5835 16.5420 52.6770 ;
        RECT 16.4080 51.5835 16.4340 52.6770 ;
        RECT 16.3000 51.5835 16.3260 52.6770 ;
        RECT 16.0870 51.5835 16.1640 52.6770 ;
        RECT 14.1940 51.5835 14.2710 52.6770 ;
        RECT 14.0320 51.5835 14.0580 52.6770 ;
        RECT 13.9240 51.5835 13.9500 52.6770 ;
        RECT 13.8160 51.5835 13.8420 52.6770 ;
        RECT 13.7080 51.5835 13.7340 52.6770 ;
        RECT 13.6000 51.5835 13.6260 52.6770 ;
        RECT 13.4920 51.5835 13.5180 52.6770 ;
        RECT 13.3840 51.5835 13.4100 52.6770 ;
        RECT 13.2760 51.5835 13.3020 52.6770 ;
        RECT 13.1680 51.5835 13.1940 52.6770 ;
        RECT 13.0600 51.5835 13.0860 52.6770 ;
        RECT 12.9520 51.5835 12.9780 52.6770 ;
        RECT 12.8440 51.5835 12.8700 52.6770 ;
        RECT 12.7360 51.5835 12.7620 52.6770 ;
        RECT 12.6280 51.5835 12.6540 52.6770 ;
        RECT 12.5200 51.5835 12.5460 52.6770 ;
        RECT 12.4120 51.5835 12.4380 52.6770 ;
        RECT 12.3040 51.5835 12.3300 52.6770 ;
        RECT 12.1960 51.5835 12.2220 52.6770 ;
        RECT 12.0880 51.5835 12.1140 52.6770 ;
        RECT 11.9800 51.5835 12.0060 52.6770 ;
        RECT 11.8720 51.5835 11.8980 52.6770 ;
        RECT 11.7640 51.5835 11.7900 52.6770 ;
        RECT 11.6560 51.5835 11.6820 52.6770 ;
        RECT 11.5480 51.5835 11.5740 52.6770 ;
        RECT 11.4400 51.5835 11.4660 52.6770 ;
        RECT 11.3320 51.5835 11.3580 52.6770 ;
        RECT 11.2240 51.5835 11.2500 52.6770 ;
        RECT 11.1160 51.5835 11.1420 52.6770 ;
        RECT 11.0080 51.5835 11.0340 52.6770 ;
        RECT 10.9000 51.5835 10.9260 52.6770 ;
        RECT 10.7920 51.5835 10.8180 52.6770 ;
        RECT 10.6840 51.5835 10.7100 52.6770 ;
        RECT 10.5760 51.5835 10.6020 52.6770 ;
        RECT 10.4680 51.5835 10.4940 52.6770 ;
        RECT 10.3600 51.5835 10.3860 52.6770 ;
        RECT 10.2520 51.5835 10.2780 52.6770 ;
        RECT 10.1440 51.5835 10.1700 52.6770 ;
        RECT 10.0360 51.5835 10.0620 52.6770 ;
        RECT 9.9280 51.5835 9.9540 52.6770 ;
        RECT 9.8200 51.5835 9.8460 52.6770 ;
        RECT 9.7120 51.5835 9.7380 52.6770 ;
        RECT 9.6040 51.5835 9.6300 52.6770 ;
        RECT 9.4960 51.5835 9.5220 52.6770 ;
        RECT 9.3880 51.5835 9.4140 52.6770 ;
        RECT 9.2800 51.5835 9.3060 52.6770 ;
        RECT 9.1720 51.5835 9.1980 52.6770 ;
        RECT 9.0640 51.5835 9.0900 52.6770 ;
        RECT 8.9560 51.5835 8.9820 52.6770 ;
        RECT 8.8480 51.5835 8.8740 52.6770 ;
        RECT 8.7400 51.5835 8.7660 52.6770 ;
        RECT 8.6320 51.5835 8.6580 52.6770 ;
        RECT 8.5240 51.5835 8.5500 52.6770 ;
        RECT 8.4160 51.5835 8.4420 52.6770 ;
        RECT 8.3080 51.5835 8.3340 52.6770 ;
        RECT 8.2000 51.5835 8.2260 52.6770 ;
        RECT 8.0920 51.5835 8.1180 52.6770 ;
        RECT 7.9840 51.5835 8.0100 52.6770 ;
        RECT 7.8760 51.5835 7.9020 52.6770 ;
        RECT 7.7680 51.5835 7.7940 52.6770 ;
        RECT 7.6600 51.5835 7.6860 52.6770 ;
        RECT 7.5520 51.5835 7.5780 52.6770 ;
        RECT 7.4440 51.5835 7.4700 52.6770 ;
        RECT 7.3360 51.5835 7.3620 52.6770 ;
        RECT 7.2280 51.5835 7.2540 52.6770 ;
        RECT 7.1200 51.5835 7.1460 52.6770 ;
        RECT 7.0120 51.5835 7.0380 52.6770 ;
        RECT 6.9040 51.5835 6.9300 52.6770 ;
        RECT 6.7960 51.5835 6.8220 52.6770 ;
        RECT 6.6880 51.5835 6.7140 52.6770 ;
        RECT 6.5800 51.5835 6.6060 52.6770 ;
        RECT 6.4720 51.5835 6.4980 52.6770 ;
        RECT 6.3640 51.5835 6.3900 52.6770 ;
        RECT 6.2560 51.5835 6.2820 52.6770 ;
        RECT 6.1480 51.5835 6.1740 52.6770 ;
        RECT 6.0400 51.5835 6.0660 52.6770 ;
        RECT 5.9320 51.5835 5.9580 52.6770 ;
        RECT 5.8240 51.5835 5.8500 52.6770 ;
        RECT 5.7160 51.5835 5.7420 52.6770 ;
        RECT 5.6080 51.5835 5.6340 52.6770 ;
        RECT 5.5000 51.5835 5.5260 52.6770 ;
        RECT 5.3920 51.5835 5.4180 52.6770 ;
        RECT 5.2840 51.5835 5.3100 52.6770 ;
        RECT 5.1760 51.5835 5.2020 52.6770 ;
        RECT 5.0680 51.5835 5.0940 52.6770 ;
        RECT 4.9600 51.5835 4.9860 52.6770 ;
        RECT 4.8520 51.5835 4.8780 52.6770 ;
        RECT 4.7440 51.5835 4.7700 52.6770 ;
        RECT 4.6360 51.5835 4.6620 52.6770 ;
        RECT 4.5280 51.5835 4.5540 52.6770 ;
        RECT 4.4200 51.5835 4.4460 52.6770 ;
        RECT 4.3120 51.5835 4.3380 52.6770 ;
        RECT 4.2040 51.5835 4.2300 52.6770 ;
        RECT 4.0960 51.5835 4.1220 52.6770 ;
        RECT 3.9880 51.5835 4.0140 52.6770 ;
        RECT 3.8800 51.5835 3.9060 52.6770 ;
        RECT 3.7720 51.5835 3.7980 52.6770 ;
        RECT 3.6640 51.5835 3.6900 52.6770 ;
        RECT 3.5560 51.5835 3.5820 52.6770 ;
        RECT 3.4480 51.5835 3.4740 52.6770 ;
        RECT 3.3400 51.5835 3.3660 52.6770 ;
        RECT 3.2320 51.5835 3.2580 52.6770 ;
        RECT 3.1240 51.5835 3.1500 52.6770 ;
        RECT 3.0160 51.5835 3.0420 52.6770 ;
        RECT 2.9080 51.5835 2.9340 52.6770 ;
        RECT 2.8000 51.5835 2.8260 52.6770 ;
        RECT 2.6920 51.5835 2.7180 52.6770 ;
        RECT 2.5840 51.5835 2.6100 52.6770 ;
        RECT 2.4760 51.5835 2.5020 52.6770 ;
        RECT 2.3680 51.5835 2.3940 52.6770 ;
        RECT 2.2600 51.5835 2.2860 52.6770 ;
        RECT 2.1520 51.5835 2.1780 52.6770 ;
        RECT 2.0440 51.5835 2.0700 52.6770 ;
        RECT 1.9360 51.5835 1.9620 52.6770 ;
        RECT 1.8280 51.5835 1.8540 52.6770 ;
        RECT 1.7200 51.5835 1.7460 52.6770 ;
        RECT 1.6120 51.5835 1.6380 52.6770 ;
        RECT 1.5040 51.5835 1.5300 52.6770 ;
        RECT 1.3960 51.5835 1.4220 52.6770 ;
        RECT 1.2880 51.5835 1.3140 52.6770 ;
        RECT 1.1800 51.5835 1.2060 52.6770 ;
        RECT 1.0720 51.5835 1.0980 52.6770 ;
        RECT 0.9640 51.5835 0.9900 52.6770 ;
        RECT 0.8560 51.5835 0.8820 52.6770 ;
        RECT 0.7480 51.5835 0.7740 52.6770 ;
        RECT 0.6400 51.5835 0.6660 52.6770 ;
        RECT 0.5320 51.5835 0.5580 52.6770 ;
        RECT 0.4240 51.5835 0.4500 52.6770 ;
        RECT 0.3160 51.5835 0.3420 52.6770 ;
        RECT 0.2080 51.5835 0.2340 52.6770 ;
        RECT 0.0050 51.5835 0.0900 52.6770 ;
        RECT 15.5530 52.6635 15.6810 53.7570 ;
        RECT 15.5390 53.3290 15.6810 53.6515 ;
        RECT 15.3190 53.0560 15.4530 53.7570 ;
        RECT 15.2960 53.3910 15.4530 53.6490 ;
        RECT 15.3190 52.6635 15.4170 53.7570 ;
        RECT 15.3190 52.7845 15.4310 53.0240 ;
        RECT 15.3190 52.6635 15.4530 52.7525 ;
        RECT 15.0940 53.1140 15.2280 53.7570 ;
        RECT 15.0940 52.6635 15.1920 53.7570 ;
        RECT 14.6770 52.6635 14.7600 53.7570 ;
        RECT 14.6770 52.7520 14.7740 53.6875 ;
        RECT 30.2680 52.6635 30.3530 53.7570 ;
        RECT 30.1240 52.6635 30.1500 53.7570 ;
        RECT 30.0160 52.6635 30.0420 53.7570 ;
        RECT 29.9080 52.6635 29.9340 53.7570 ;
        RECT 29.8000 52.6635 29.8260 53.7570 ;
        RECT 29.6920 52.6635 29.7180 53.7570 ;
        RECT 29.5840 52.6635 29.6100 53.7570 ;
        RECT 29.4760 52.6635 29.5020 53.7570 ;
        RECT 29.3680 52.6635 29.3940 53.7570 ;
        RECT 29.2600 52.6635 29.2860 53.7570 ;
        RECT 29.1520 52.6635 29.1780 53.7570 ;
        RECT 29.0440 52.6635 29.0700 53.7570 ;
        RECT 28.9360 52.6635 28.9620 53.7570 ;
        RECT 28.8280 52.6635 28.8540 53.7570 ;
        RECT 28.7200 52.6635 28.7460 53.7570 ;
        RECT 28.6120 52.6635 28.6380 53.7570 ;
        RECT 28.5040 52.6635 28.5300 53.7570 ;
        RECT 28.3960 52.6635 28.4220 53.7570 ;
        RECT 28.2880 52.6635 28.3140 53.7570 ;
        RECT 28.1800 52.6635 28.2060 53.7570 ;
        RECT 28.0720 52.6635 28.0980 53.7570 ;
        RECT 27.9640 52.6635 27.9900 53.7570 ;
        RECT 27.8560 52.6635 27.8820 53.7570 ;
        RECT 27.7480 52.6635 27.7740 53.7570 ;
        RECT 27.6400 52.6635 27.6660 53.7570 ;
        RECT 27.5320 52.6635 27.5580 53.7570 ;
        RECT 27.4240 52.6635 27.4500 53.7570 ;
        RECT 27.3160 52.6635 27.3420 53.7570 ;
        RECT 27.2080 52.6635 27.2340 53.7570 ;
        RECT 27.1000 52.6635 27.1260 53.7570 ;
        RECT 26.9920 52.6635 27.0180 53.7570 ;
        RECT 26.8840 52.6635 26.9100 53.7570 ;
        RECT 26.7760 52.6635 26.8020 53.7570 ;
        RECT 26.6680 52.6635 26.6940 53.7570 ;
        RECT 26.5600 52.6635 26.5860 53.7570 ;
        RECT 26.4520 52.6635 26.4780 53.7570 ;
        RECT 26.3440 52.6635 26.3700 53.7570 ;
        RECT 26.2360 52.6635 26.2620 53.7570 ;
        RECT 26.1280 52.6635 26.1540 53.7570 ;
        RECT 26.0200 52.6635 26.0460 53.7570 ;
        RECT 25.9120 52.6635 25.9380 53.7570 ;
        RECT 25.8040 52.6635 25.8300 53.7570 ;
        RECT 25.6960 52.6635 25.7220 53.7570 ;
        RECT 25.5880 52.6635 25.6140 53.7570 ;
        RECT 25.4800 52.6635 25.5060 53.7570 ;
        RECT 25.3720 52.6635 25.3980 53.7570 ;
        RECT 25.2640 52.6635 25.2900 53.7570 ;
        RECT 25.1560 52.6635 25.1820 53.7570 ;
        RECT 25.0480 52.6635 25.0740 53.7570 ;
        RECT 24.9400 52.6635 24.9660 53.7570 ;
        RECT 24.8320 52.6635 24.8580 53.7570 ;
        RECT 24.7240 52.6635 24.7500 53.7570 ;
        RECT 24.6160 52.6635 24.6420 53.7570 ;
        RECT 24.5080 52.6635 24.5340 53.7570 ;
        RECT 24.4000 52.6635 24.4260 53.7570 ;
        RECT 24.2920 52.6635 24.3180 53.7570 ;
        RECT 24.1840 52.6635 24.2100 53.7570 ;
        RECT 24.0760 52.6635 24.1020 53.7570 ;
        RECT 23.9680 52.6635 23.9940 53.7570 ;
        RECT 23.8600 52.6635 23.8860 53.7570 ;
        RECT 23.7520 52.6635 23.7780 53.7570 ;
        RECT 23.6440 52.6635 23.6700 53.7570 ;
        RECT 23.5360 52.6635 23.5620 53.7570 ;
        RECT 23.4280 52.6635 23.4540 53.7570 ;
        RECT 23.3200 52.6635 23.3460 53.7570 ;
        RECT 23.2120 52.6635 23.2380 53.7570 ;
        RECT 23.1040 52.6635 23.1300 53.7570 ;
        RECT 22.9960 52.6635 23.0220 53.7570 ;
        RECT 22.8880 52.6635 22.9140 53.7570 ;
        RECT 22.7800 52.6635 22.8060 53.7570 ;
        RECT 22.6720 52.6635 22.6980 53.7570 ;
        RECT 22.5640 52.6635 22.5900 53.7570 ;
        RECT 22.4560 52.6635 22.4820 53.7570 ;
        RECT 22.3480 52.6635 22.3740 53.7570 ;
        RECT 22.2400 52.6635 22.2660 53.7570 ;
        RECT 22.1320 52.6635 22.1580 53.7570 ;
        RECT 22.0240 52.6635 22.0500 53.7570 ;
        RECT 21.9160 52.6635 21.9420 53.7570 ;
        RECT 21.8080 52.6635 21.8340 53.7570 ;
        RECT 21.7000 52.6635 21.7260 53.7570 ;
        RECT 21.5920 52.6635 21.6180 53.7570 ;
        RECT 21.4840 52.6635 21.5100 53.7570 ;
        RECT 21.3760 52.6635 21.4020 53.7570 ;
        RECT 21.2680 52.6635 21.2940 53.7570 ;
        RECT 21.1600 52.6635 21.1860 53.7570 ;
        RECT 21.0520 52.6635 21.0780 53.7570 ;
        RECT 20.9440 52.6635 20.9700 53.7570 ;
        RECT 20.8360 52.6635 20.8620 53.7570 ;
        RECT 20.7280 52.6635 20.7540 53.7570 ;
        RECT 20.6200 52.6635 20.6460 53.7570 ;
        RECT 20.5120 52.6635 20.5380 53.7570 ;
        RECT 20.4040 52.6635 20.4300 53.7570 ;
        RECT 20.2960 52.6635 20.3220 53.7570 ;
        RECT 20.1880 52.6635 20.2140 53.7570 ;
        RECT 20.0800 52.6635 20.1060 53.7570 ;
        RECT 19.9720 52.6635 19.9980 53.7570 ;
        RECT 19.8640 52.6635 19.8900 53.7570 ;
        RECT 19.7560 52.6635 19.7820 53.7570 ;
        RECT 19.6480 52.6635 19.6740 53.7570 ;
        RECT 19.5400 52.6635 19.5660 53.7570 ;
        RECT 19.4320 52.6635 19.4580 53.7570 ;
        RECT 19.3240 52.6635 19.3500 53.7570 ;
        RECT 19.2160 52.6635 19.2420 53.7570 ;
        RECT 19.1080 52.6635 19.1340 53.7570 ;
        RECT 19.0000 52.6635 19.0260 53.7570 ;
        RECT 18.8920 52.6635 18.9180 53.7570 ;
        RECT 18.7840 52.6635 18.8100 53.7570 ;
        RECT 18.6760 52.6635 18.7020 53.7570 ;
        RECT 18.5680 52.6635 18.5940 53.7570 ;
        RECT 18.4600 52.6635 18.4860 53.7570 ;
        RECT 18.3520 52.6635 18.3780 53.7570 ;
        RECT 18.2440 52.6635 18.2700 53.7570 ;
        RECT 18.1360 52.6635 18.1620 53.7570 ;
        RECT 18.0280 52.6635 18.0540 53.7570 ;
        RECT 17.9200 52.6635 17.9460 53.7570 ;
        RECT 17.8120 52.6635 17.8380 53.7570 ;
        RECT 17.7040 52.6635 17.7300 53.7570 ;
        RECT 17.5960 52.6635 17.6220 53.7570 ;
        RECT 17.4880 52.6635 17.5140 53.7570 ;
        RECT 17.3800 52.6635 17.4060 53.7570 ;
        RECT 17.2720 52.6635 17.2980 53.7570 ;
        RECT 17.1640 52.6635 17.1900 53.7570 ;
        RECT 17.0560 52.6635 17.0820 53.7570 ;
        RECT 16.9480 52.6635 16.9740 53.7570 ;
        RECT 16.8400 52.6635 16.8660 53.7570 ;
        RECT 16.7320 52.6635 16.7580 53.7570 ;
        RECT 16.6240 52.6635 16.6500 53.7570 ;
        RECT 16.5160 52.6635 16.5420 53.7570 ;
        RECT 16.4080 52.6635 16.4340 53.7570 ;
        RECT 16.3000 52.6635 16.3260 53.7570 ;
        RECT 16.0870 52.6635 16.1640 53.7570 ;
        RECT 14.1940 52.6635 14.2710 53.7570 ;
        RECT 14.0320 52.6635 14.0580 53.7570 ;
        RECT 13.9240 52.6635 13.9500 53.7570 ;
        RECT 13.8160 52.6635 13.8420 53.7570 ;
        RECT 13.7080 52.6635 13.7340 53.7570 ;
        RECT 13.6000 52.6635 13.6260 53.7570 ;
        RECT 13.4920 52.6635 13.5180 53.7570 ;
        RECT 13.3840 52.6635 13.4100 53.7570 ;
        RECT 13.2760 52.6635 13.3020 53.7570 ;
        RECT 13.1680 52.6635 13.1940 53.7570 ;
        RECT 13.0600 52.6635 13.0860 53.7570 ;
        RECT 12.9520 52.6635 12.9780 53.7570 ;
        RECT 12.8440 52.6635 12.8700 53.7570 ;
        RECT 12.7360 52.6635 12.7620 53.7570 ;
        RECT 12.6280 52.6635 12.6540 53.7570 ;
        RECT 12.5200 52.6635 12.5460 53.7570 ;
        RECT 12.4120 52.6635 12.4380 53.7570 ;
        RECT 12.3040 52.6635 12.3300 53.7570 ;
        RECT 12.1960 52.6635 12.2220 53.7570 ;
        RECT 12.0880 52.6635 12.1140 53.7570 ;
        RECT 11.9800 52.6635 12.0060 53.7570 ;
        RECT 11.8720 52.6635 11.8980 53.7570 ;
        RECT 11.7640 52.6635 11.7900 53.7570 ;
        RECT 11.6560 52.6635 11.6820 53.7570 ;
        RECT 11.5480 52.6635 11.5740 53.7570 ;
        RECT 11.4400 52.6635 11.4660 53.7570 ;
        RECT 11.3320 52.6635 11.3580 53.7570 ;
        RECT 11.2240 52.6635 11.2500 53.7570 ;
        RECT 11.1160 52.6635 11.1420 53.7570 ;
        RECT 11.0080 52.6635 11.0340 53.7570 ;
        RECT 10.9000 52.6635 10.9260 53.7570 ;
        RECT 10.7920 52.6635 10.8180 53.7570 ;
        RECT 10.6840 52.6635 10.7100 53.7570 ;
        RECT 10.5760 52.6635 10.6020 53.7570 ;
        RECT 10.4680 52.6635 10.4940 53.7570 ;
        RECT 10.3600 52.6635 10.3860 53.7570 ;
        RECT 10.2520 52.6635 10.2780 53.7570 ;
        RECT 10.1440 52.6635 10.1700 53.7570 ;
        RECT 10.0360 52.6635 10.0620 53.7570 ;
        RECT 9.9280 52.6635 9.9540 53.7570 ;
        RECT 9.8200 52.6635 9.8460 53.7570 ;
        RECT 9.7120 52.6635 9.7380 53.7570 ;
        RECT 9.6040 52.6635 9.6300 53.7570 ;
        RECT 9.4960 52.6635 9.5220 53.7570 ;
        RECT 9.3880 52.6635 9.4140 53.7570 ;
        RECT 9.2800 52.6635 9.3060 53.7570 ;
        RECT 9.1720 52.6635 9.1980 53.7570 ;
        RECT 9.0640 52.6635 9.0900 53.7570 ;
        RECT 8.9560 52.6635 8.9820 53.7570 ;
        RECT 8.8480 52.6635 8.8740 53.7570 ;
        RECT 8.7400 52.6635 8.7660 53.7570 ;
        RECT 8.6320 52.6635 8.6580 53.7570 ;
        RECT 8.5240 52.6635 8.5500 53.7570 ;
        RECT 8.4160 52.6635 8.4420 53.7570 ;
        RECT 8.3080 52.6635 8.3340 53.7570 ;
        RECT 8.2000 52.6635 8.2260 53.7570 ;
        RECT 8.0920 52.6635 8.1180 53.7570 ;
        RECT 7.9840 52.6635 8.0100 53.7570 ;
        RECT 7.8760 52.6635 7.9020 53.7570 ;
        RECT 7.7680 52.6635 7.7940 53.7570 ;
        RECT 7.6600 52.6635 7.6860 53.7570 ;
        RECT 7.5520 52.6635 7.5780 53.7570 ;
        RECT 7.4440 52.6635 7.4700 53.7570 ;
        RECT 7.3360 52.6635 7.3620 53.7570 ;
        RECT 7.2280 52.6635 7.2540 53.7570 ;
        RECT 7.1200 52.6635 7.1460 53.7570 ;
        RECT 7.0120 52.6635 7.0380 53.7570 ;
        RECT 6.9040 52.6635 6.9300 53.7570 ;
        RECT 6.7960 52.6635 6.8220 53.7570 ;
        RECT 6.6880 52.6635 6.7140 53.7570 ;
        RECT 6.5800 52.6635 6.6060 53.7570 ;
        RECT 6.4720 52.6635 6.4980 53.7570 ;
        RECT 6.3640 52.6635 6.3900 53.7570 ;
        RECT 6.2560 52.6635 6.2820 53.7570 ;
        RECT 6.1480 52.6635 6.1740 53.7570 ;
        RECT 6.0400 52.6635 6.0660 53.7570 ;
        RECT 5.9320 52.6635 5.9580 53.7570 ;
        RECT 5.8240 52.6635 5.8500 53.7570 ;
        RECT 5.7160 52.6635 5.7420 53.7570 ;
        RECT 5.6080 52.6635 5.6340 53.7570 ;
        RECT 5.5000 52.6635 5.5260 53.7570 ;
        RECT 5.3920 52.6635 5.4180 53.7570 ;
        RECT 5.2840 52.6635 5.3100 53.7570 ;
        RECT 5.1760 52.6635 5.2020 53.7570 ;
        RECT 5.0680 52.6635 5.0940 53.7570 ;
        RECT 4.9600 52.6635 4.9860 53.7570 ;
        RECT 4.8520 52.6635 4.8780 53.7570 ;
        RECT 4.7440 52.6635 4.7700 53.7570 ;
        RECT 4.6360 52.6635 4.6620 53.7570 ;
        RECT 4.5280 52.6635 4.5540 53.7570 ;
        RECT 4.4200 52.6635 4.4460 53.7570 ;
        RECT 4.3120 52.6635 4.3380 53.7570 ;
        RECT 4.2040 52.6635 4.2300 53.7570 ;
        RECT 4.0960 52.6635 4.1220 53.7570 ;
        RECT 3.9880 52.6635 4.0140 53.7570 ;
        RECT 3.8800 52.6635 3.9060 53.7570 ;
        RECT 3.7720 52.6635 3.7980 53.7570 ;
        RECT 3.6640 52.6635 3.6900 53.7570 ;
        RECT 3.5560 52.6635 3.5820 53.7570 ;
        RECT 3.4480 52.6635 3.4740 53.7570 ;
        RECT 3.3400 52.6635 3.3660 53.7570 ;
        RECT 3.2320 52.6635 3.2580 53.7570 ;
        RECT 3.1240 52.6635 3.1500 53.7570 ;
        RECT 3.0160 52.6635 3.0420 53.7570 ;
        RECT 2.9080 52.6635 2.9340 53.7570 ;
        RECT 2.8000 52.6635 2.8260 53.7570 ;
        RECT 2.6920 52.6635 2.7180 53.7570 ;
        RECT 2.5840 52.6635 2.6100 53.7570 ;
        RECT 2.4760 52.6635 2.5020 53.7570 ;
        RECT 2.3680 52.6635 2.3940 53.7570 ;
        RECT 2.2600 52.6635 2.2860 53.7570 ;
        RECT 2.1520 52.6635 2.1780 53.7570 ;
        RECT 2.0440 52.6635 2.0700 53.7570 ;
        RECT 1.9360 52.6635 1.9620 53.7570 ;
        RECT 1.8280 52.6635 1.8540 53.7570 ;
        RECT 1.7200 52.6635 1.7460 53.7570 ;
        RECT 1.6120 52.6635 1.6380 53.7570 ;
        RECT 1.5040 52.6635 1.5300 53.7570 ;
        RECT 1.3960 52.6635 1.4220 53.7570 ;
        RECT 1.2880 52.6635 1.3140 53.7570 ;
        RECT 1.1800 52.6635 1.2060 53.7570 ;
        RECT 1.0720 52.6635 1.0980 53.7570 ;
        RECT 0.9640 52.6635 0.9900 53.7570 ;
        RECT 0.8560 52.6635 0.8820 53.7570 ;
        RECT 0.7480 52.6635 0.7740 53.7570 ;
        RECT 0.6400 52.6635 0.6660 53.7570 ;
        RECT 0.5320 52.6635 0.5580 53.7570 ;
        RECT 0.4240 52.6635 0.4500 53.7570 ;
        RECT 0.3160 52.6635 0.3420 53.7570 ;
        RECT 0.2080 52.6635 0.2340 53.7570 ;
        RECT 0.0050 52.6635 0.0900 53.7570 ;
        RECT 15.5530 53.7435 15.6810 54.8370 ;
        RECT 15.5390 54.4090 15.6810 54.7315 ;
        RECT 15.3190 54.1360 15.4530 54.8370 ;
        RECT 15.2960 54.4710 15.4530 54.7290 ;
        RECT 15.3190 53.7435 15.4170 54.8370 ;
        RECT 15.3190 53.8645 15.4310 54.1040 ;
        RECT 15.3190 53.7435 15.4530 53.8325 ;
        RECT 15.0940 54.1940 15.2280 54.8370 ;
        RECT 15.0940 53.7435 15.1920 54.8370 ;
        RECT 14.6770 53.7435 14.7600 54.8370 ;
        RECT 14.6770 53.8320 14.7740 54.7675 ;
        RECT 30.2680 53.7435 30.3530 54.8370 ;
        RECT 30.1240 53.7435 30.1500 54.8370 ;
        RECT 30.0160 53.7435 30.0420 54.8370 ;
        RECT 29.9080 53.7435 29.9340 54.8370 ;
        RECT 29.8000 53.7435 29.8260 54.8370 ;
        RECT 29.6920 53.7435 29.7180 54.8370 ;
        RECT 29.5840 53.7435 29.6100 54.8370 ;
        RECT 29.4760 53.7435 29.5020 54.8370 ;
        RECT 29.3680 53.7435 29.3940 54.8370 ;
        RECT 29.2600 53.7435 29.2860 54.8370 ;
        RECT 29.1520 53.7435 29.1780 54.8370 ;
        RECT 29.0440 53.7435 29.0700 54.8370 ;
        RECT 28.9360 53.7435 28.9620 54.8370 ;
        RECT 28.8280 53.7435 28.8540 54.8370 ;
        RECT 28.7200 53.7435 28.7460 54.8370 ;
        RECT 28.6120 53.7435 28.6380 54.8370 ;
        RECT 28.5040 53.7435 28.5300 54.8370 ;
        RECT 28.3960 53.7435 28.4220 54.8370 ;
        RECT 28.2880 53.7435 28.3140 54.8370 ;
        RECT 28.1800 53.7435 28.2060 54.8370 ;
        RECT 28.0720 53.7435 28.0980 54.8370 ;
        RECT 27.9640 53.7435 27.9900 54.8370 ;
        RECT 27.8560 53.7435 27.8820 54.8370 ;
        RECT 27.7480 53.7435 27.7740 54.8370 ;
        RECT 27.6400 53.7435 27.6660 54.8370 ;
        RECT 27.5320 53.7435 27.5580 54.8370 ;
        RECT 27.4240 53.7435 27.4500 54.8370 ;
        RECT 27.3160 53.7435 27.3420 54.8370 ;
        RECT 27.2080 53.7435 27.2340 54.8370 ;
        RECT 27.1000 53.7435 27.1260 54.8370 ;
        RECT 26.9920 53.7435 27.0180 54.8370 ;
        RECT 26.8840 53.7435 26.9100 54.8370 ;
        RECT 26.7760 53.7435 26.8020 54.8370 ;
        RECT 26.6680 53.7435 26.6940 54.8370 ;
        RECT 26.5600 53.7435 26.5860 54.8370 ;
        RECT 26.4520 53.7435 26.4780 54.8370 ;
        RECT 26.3440 53.7435 26.3700 54.8370 ;
        RECT 26.2360 53.7435 26.2620 54.8370 ;
        RECT 26.1280 53.7435 26.1540 54.8370 ;
        RECT 26.0200 53.7435 26.0460 54.8370 ;
        RECT 25.9120 53.7435 25.9380 54.8370 ;
        RECT 25.8040 53.7435 25.8300 54.8370 ;
        RECT 25.6960 53.7435 25.7220 54.8370 ;
        RECT 25.5880 53.7435 25.6140 54.8370 ;
        RECT 25.4800 53.7435 25.5060 54.8370 ;
        RECT 25.3720 53.7435 25.3980 54.8370 ;
        RECT 25.2640 53.7435 25.2900 54.8370 ;
        RECT 25.1560 53.7435 25.1820 54.8370 ;
        RECT 25.0480 53.7435 25.0740 54.8370 ;
        RECT 24.9400 53.7435 24.9660 54.8370 ;
        RECT 24.8320 53.7435 24.8580 54.8370 ;
        RECT 24.7240 53.7435 24.7500 54.8370 ;
        RECT 24.6160 53.7435 24.6420 54.8370 ;
        RECT 24.5080 53.7435 24.5340 54.8370 ;
        RECT 24.4000 53.7435 24.4260 54.8370 ;
        RECT 24.2920 53.7435 24.3180 54.8370 ;
        RECT 24.1840 53.7435 24.2100 54.8370 ;
        RECT 24.0760 53.7435 24.1020 54.8370 ;
        RECT 23.9680 53.7435 23.9940 54.8370 ;
        RECT 23.8600 53.7435 23.8860 54.8370 ;
        RECT 23.7520 53.7435 23.7780 54.8370 ;
        RECT 23.6440 53.7435 23.6700 54.8370 ;
        RECT 23.5360 53.7435 23.5620 54.8370 ;
        RECT 23.4280 53.7435 23.4540 54.8370 ;
        RECT 23.3200 53.7435 23.3460 54.8370 ;
        RECT 23.2120 53.7435 23.2380 54.8370 ;
        RECT 23.1040 53.7435 23.1300 54.8370 ;
        RECT 22.9960 53.7435 23.0220 54.8370 ;
        RECT 22.8880 53.7435 22.9140 54.8370 ;
        RECT 22.7800 53.7435 22.8060 54.8370 ;
        RECT 22.6720 53.7435 22.6980 54.8370 ;
        RECT 22.5640 53.7435 22.5900 54.8370 ;
        RECT 22.4560 53.7435 22.4820 54.8370 ;
        RECT 22.3480 53.7435 22.3740 54.8370 ;
        RECT 22.2400 53.7435 22.2660 54.8370 ;
        RECT 22.1320 53.7435 22.1580 54.8370 ;
        RECT 22.0240 53.7435 22.0500 54.8370 ;
        RECT 21.9160 53.7435 21.9420 54.8370 ;
        RECT 21.8080 53.7435 21.8340 54.8370 ;
        RECT 21.7000 53.7435 21.7260 54.8370 ;
        RECT 21.5920 53.7435 21.6180 54.8370 ;
        RECT 21.4840 53.7435 21.5100 54.8370 ;
        RECT 21.3760 53.7435 21.4020 54.8370 ;
        RECT 21.2680 53.7435 21.2940 54.8370 ;
        RECT 21.1600 53.7435 21.1860 54.8370 ;
        RECT 21.0520 53.7435 21.0780 54.8370 ;
        RECT 20.9440 53.7435 20.9700 54.8370 ;
        RECT 20.8360 53.7435 20.8620 54.8370 ;
        RECT 20.7280 53.7435 20.7540 54.8370 ;
        RECT 20.6200 53.7435 20.6460 54.8370 ;
        RECT 20.5120 53.7435 20.5380 54.8370 ;
        RECT 20.4040 53.7435 20.4300 54.8370 ;
        RECT 20.2960 53.7435 20.3220 54.8370 ;
        RECT 20.1880 53.7435 20.2140 54.8370 ;
        RECT 20.0800 53.7435 20.1060 54.8370 ;
        RECT 19.9720 53.7435 19.9980 54.8370 ;
        RECT 19.8640 53.7435 19.8900 54.8370 ;
        RECT 19.7560 53.7435 19.7820 54.8370 ;
        RECT 19.6480 53.7435 19.6740 54.8370 ;
        RECT 19.5400 53.7435 19.5660 54.8370 ;
        RECT 19.4320 53.7435 19.4580 54.8370 ;
        RECT 19.3240 53.7435 19.3500 54.8370 ;
        RECT 19.2160 53.7435 19.2420 54.8370 ;
        RECT 19.1080 53.7435 19.1340 54.8370 ;
        RECT 19.0000 53.7435 19.0260 54.8370 ;
        RECT 18.8920 53.7435 18.9180 54.8370 ;
        RECT 18.7840 53.7435 18.8100 54.8370 ;
        RECT 18.6760 53.7435 18.7020 54.8370 ;
        RECT 18.5680 53.7435 18.5940 54.8370 ;
        RECT 18.4600 53.7435 18.4860 54.8370 ;
        RECT 18.3520 53.7435 18.3780 54.8370 ;
        RECT 18.2440 53.7435 18.2700 54.8370 ;
        RECT 18.1360 53.7435 18.1620 54.8370 ;
        RECT 18.0280 53.7435 18.0540 54.8370 ;
        RECT 17.9200 53.7435 17.9460 54.8370 ;
        RECT 17.8120 53.7435 17.8380 54.8370 ;
        RECT 17.7040 53.7435 17.7300 54.8370 ;
        RECT 17.5960 53.7435 17.6220 54.8370 ;
        RECT 17.4880 53.7435 17.5140 54.8370 ;
        RECT 17.3800 53.7435 17.4060 54.8370 ;
        RECT 17.2720 53.7435 17.2980 54.8370 ;
        RECT 17.1640 53.7435 17.1900 54.8370 ;
        RECT 17.0560 53.7435 17.0820 54.8370 ;
        RECT 16.9480 53.7435 16.9740 54.8370 ;
        RECT 16.8400 53.7435 16.8660 54.8370 ;
        RECT 16.7320 53.7435 16.7580 54.8370 ;
        RECT 16.6240 53.7435 16.6500 54.8370 ;
        RECT 16.5160 53.7435 16.5420 54.8370 ;
        RECT 16.4080 53.7435 16.4340 54.8370 ;
        RECT 16.3000 53.7435 16.3260 54.8370 ;
        RECT 16.0870 53.7435 16.1640 54.8370 ;
        RECT 14.1940 53.7435 14.2710 54.8370 ;
        RECT 14.0320 53.7435 14.0580 54.8370 ;
        RECT 13.9240 53.7435 13.9500 54.8370 ;
        RECT 13.8160 53.7435 13.8420 54.8370 ;
        RECT 13.7080 53.7435 13.7340 54.8370 ;
        RECT 13.6000 53.7435 13.6260 54.8370 ;
        RECT 13.4920 53.7435 13.5180 54.8370 ;
        RECT 13.3840 53.7435 13.4100 54.8370 ;
        RECT 13.2760 53.7435 13.3020 54.8370 ;
        RECT 13.1680 53.7435 13.1940 54.8370 ;
        RECT 13.0600 53.7435 13.0860 54.8370 ;
        RECT 12.9520 53.7435 12.9780 54.8370 ;
        RECT 12.8440 53.7435 12.8700 54.8370 ;
        RECT 12.7360 53.7435 12.7620 54.8370 ;
        RECT 12.6280 53.7435 12.6540 54.8370 ;
        RECT 12.5200 53.7435 12.5460 54.8370 ;
        RECT 12.4120 53.7435 12.4380 54.8370 ;
        RECT 12.3040 53.7435 12.3300 54.8370 ;
        RECT 12.1960 53.7435 12.2220 54.8370 ;
        RECT 12.0880 53.7435 12.1140 54.8370 ;
        RECT 11.9800 53.7435 12.0060 54.8370 ;
        RECT 11.8720 53.7435 11.8980 54.8370 ;
        RECT 11.7640 53.7435 11.7900 54.8370 ;
        RECT 11.6560 53.7435 11.6820 54.8370 ;
        RECT 11.5480 53.7435 11.5740 54.8370 ;
        RECT 11.4400 53.7435 11.4660 54.8370 ;
        RECT 11.3320 53.7435 11.3580 54.8370 ;
        RECT 11.2240 53.7435 11.2500 54.8370 ;
        RECT 11.1160 53.7435 11.1420 54.8370 ;
        RECT 11.0080 53.7435 11.0340 54.8370 ;
        RECT 10.9000 53.7435 10.9260 54.8370 ;
        RECT 10.7920 53.7435 10.8180 54.8370 ;
        RECT 10.6840 53.7435 10.7100 54.8370 ;
        RECT 10.5760 53.7435 10.6020 54.8370 ;
        RECT 10.4680 53.7435 10.4940 54.8370 ;
        RECT 10.3600 53.7435 10.3860 54.8370 ;
        RECT 10.2520 53.7435 10.2780 54.8370 ;
        RECT 10.1440 53.7435 10.1700 54.8370 ;
        RECT 10.0360 53.7435 10.0620 54.8370 ;
        RECT 9.9280 53.7435 9.9540 54.8370 ;
        RECT 9.8200 53.7435 9.8460 54.8370 ;
        RECT 9.7120 53.7435 9.7380 54.8370 ;
        RECT 9.6040 53.7435 9.6300 54.8370 ;
        RECT 9.4960 53.7435 9.5220 54.8370 ;
        RECT 9.3880 53.7435 9.4140 54.8370 ;
        RECT 9.2800 53.7435 9.3060 54.8370 ;
        RECT 9.1720 53.7435 9.1980 54.8370 ;
        RECT 9.0640 53.7435 9.0900 54.8370 ;
        RECT 8.9560 53.7435 8.9820 54.8370 ;
        RECT 8.8480 53.7435 8.8740 54.8370 ;
        RECT 8.7400 53.7435 8.7660 54.8370 ;
        RECT 8.6320 53.7435 8.6580 54.8370 ;
        RECT 8.5240 53.7435 8.5500 54.8370 ;
        RECT 8.4160 53.7435 8.4420 54.8370 ;
        RECT 8.3080 53.7435 8.3340 54.8370 ;
        RECT 8.2000 53.7435 8.2260 54.8370 ;
        RECT 8.0920 53.7435 8.1180 54.8370 ;
        RECT 7.9840 53.7435 8.0100 54.8370 ;
        RECT 7.8760 53.7435 7.9020 54.8370 ;
        RECT 7.7680 53.7435 7.7940 54.8370 ;
        RECT 7.6600 53.7435 7.6860 54.8370 ;
        RECT 7.5520 53.7435 7.5780 54.8370 ;
        RECT 7.4440 53.7435 7.4700 54.8370 ;
        RECT 7.3360 53.7435 7.3620 54.8370 ;
        RECT 7.2280 53.7435 7.2540 54.8370 ;
        RECT 7.1200 53.7435 7.1460 54.8370 ;
        RECT 7.0120 53.7435 7.0380 54.8370 ;
        RECT 6.9040 53.7435 6.9300 54.8370 ;
        RECT 6.7960 53.7435 6.8220 54.8370 ;
        RECT 6.6880 53.7435 6.7140 54.8370 ;
        RECT 6.5800 53.7435 6.6060 54.8370 ;
        RECT 6.4720 53.7435 6.4980 54.8370 ;
        RECT 6.3640 53.7435 6.3900 54.8370 ;
        RECT 6.2560 53.7435 6.2820 54.8370 ;
        RECT 6.1480 53.7435 6.1740 54.8370 ;
        RECT 6.0400 53.7435 6.0660 54.8370 ;
        RECT 5.9320 53.7435 5.9580 54.8370 ;
        RECT 5.8240 53.7435 5.8500 54.8370 ;
        RECT 5.7160 53.7435 5.7420 54.8370 ;
        RECT 5.6080 53.7435 5.6340 54.8370 ;
        RECT 5.5000 53.7435 5.5260 54.8370 ;
        RECT 5.3920 53.7435 5.4180 54.8370 ;
        RECT 5.2840 53.7435 5.3100 54.8370 ;
        RECT 5.1760 53.7435 5.2020 54.8370 ;
        RECT 5.0680 53.7435 5.0940 54.8370 ;
        RECT 4.9600 53.7435 4.9860 54.8370 ;
        RECT 4.8520 53.7435 4.8780 54.8370 ;
        RECT 4.7440 53.7435 4.7700 54.8370 ;
        RECT 4.6360 53.7435 4.6620 54.8370 ;
        RECT 4.5280 53.7435 4.5540 54.8370 ;
        RECT 4.4200 53.7435 4.4460 54.8370 ;
        RECT 4.3120 53.7435 4.3380 54.8370 ;
        RECT 4.2040 53.7435 4.2300 54.8370 ;
        RECT 4.0960 53.7435 4.1220 54.8370 ;
        RECT 3.9880 53.7435 4.0140 54.8370 ;
        RECT 3.8800 53.7435 3.9060 54.8370 ;
        RECT 3.7720 53.7435 3.7980 54.8370 ;
        RECT 3.6640 53.7435 3.6900 54.8370 ;
        RECT 3.5560 53.7435 3.5820 54.8370 ;
        RECT 3.4480 53.7435 3.4740 54.8370 ;
        RECT 3.3400 53.7435 3.3660 54.8370 ;
        RECT 3.2320 53.7435 3.2580 54.8370 ;
        RECT 3.1240 53.7435 3.1500 54.8370 ;
        RECT 3.0160 53.7435 3.0420 54.8370 ;
        RECT 2.9080 53.7435 2.9340 54.8370 ;
        RECT 2.8000 53.7435 2.8260 54.8370 ;
        RECT 2.6920 53.7435 2.7180 54.8370 ;
        RECT 2.5840 53.7435 2.6100 54.8370 ;
        RECT 2.4760 53.7435 2.5020 54.8370 ;
        RECT 2.3680 53.7435 2.3940 54.8370 ;
        RECT 2.2600 53.7435 2.2860 54.8370 ;
        RECT 2.1520 53.7435 2.1780 54.8370 ;
        RECT 2.0440 53.7435 2.0700 54.8370 ;
        RECT 1.9360 53.7435 1.9620 54.8370 ;
        RECT 1.8280 53.7435 1.8540 54.8370 ;
        RECT 1.7200 53.7435 1.7460 54.8370 ;
        RECT 1.6120 53.7435 1.6380 54.8370 ;
        RECT 1.5040 53.7435 1.5300 54.8370 ;
        RECT 1.3960 53.7435 1.4220 54.8370 ;
        RECT 1.2880 53.7435 1.3140 54.8370 ;
        RECT 1.1800 53.7435 1.2060 54.8370 ;
        RECT 1.0720 53.7435 1.0980 54.8370 ;
        RECT 0.9640 53.7435 0.9900 54.8370 ;
        RECT 0.8560 53.7435 0.8820 54.8370 ;
        RECT 0.7480 53.7435 0.7740 54.8370 ;
        RECT 0.6400 53.7435 0.6660 54.8370 ;
        RECT 0.5320 53.7435 0.5580 54.8370 ;
        RECT 0.4240 53.7435 0.4500 54.8370 ;
        RECT 0.3160 53.7435 0.3420 54.8370 ;
        RECT 0.2080 53.7435 0.2340 54.8370 ;
        RECT 0.0050 53.7435 0.0900 54.8370 ;
        RECT 15.5530 54.8235 15.6810 55.9170 ;
        RECT 15.5390 55.4890 15.6810 55.8115 ;
        RECT 15.3190 55.2160 15.4530 55.9170 ;
        RECT 15.2960 55.5510 15.4530 55.8090 ;
        RECT 15.3190 54.8235 15.4170 55.9170 ;
        RECT 15.3190 54.9445 15.4310 55.1840 ;
        RECT 15.3190 54.8235 15.4530 54.9125 ;
        RECT 15.0940 55.2740 15.2280 55.9170 ;
        RECT 15.0940 54.8235 15.1920 55.9170 ;
        RECT 14.6770 54.8235 14.7600 55.9170 ;
        RECT 14.6770 54.9120 14.7740 55.8475 ;
        RECT 30.2680 54.8235 30.3530 55.9170 ;
        RECT 30.1240 54.8235 30.1500 55.9170 ;
        RECT 30.0160 54.8235 30.0420 55.9170 ;
        RECT 29.9080 54.8235 29.9340 55.9170 ;
        RECT 29.8000 54.8235 29.8260 55.9170 ;
        RECT 29.6920 54.8235 29.7180 55.9170 ;
        RECT 29.5840 54.8235 29.6100 55.9170 ;
        RECT 29.4760 54.8235 29.5020 55.9170 ;
        RECT 29.3680 54.8235 29.3940 55.9170 ;
        RECT 29.2600 54.8235 29.2860 55.9170 ;
        RECT 29.1520 54.8235 29.1780 55.9170 ;
        RECT 29.0440 54.8235 29.0700 55.9170 ;
        RECT 28.9360 54.8235 28.9620 55.9170 ;
        RECT 28.8280 54.8235 28.8540 55.9170 ;
        RECT 28.7200 54.8235 28.7460 55.9170 ;
        RECT 28.6120 54.8235 28.6380 55.9170 ;
        RECT 28.5040 54.8235 28.5300 55.9170 ;
        RECT 28.3960 54.8235 28.4220 55.9170 ;
        RECT 28.2880 54.8235 28.3140 55.9170 ;
        RECT 28.1800 54.8235 28.2060 55.9170 ;
        RECT 28.0720 54.8235 28.0980 55.9170 ;
        RECT 27.9640 54.8235 27.9900 55.9170 ;
        RECT 27.8560 54.8235 27.8820 55.9170 ;
        RECT 27.7480 54.8235 27.7740 55.9170 ;
        RECT 27.6400 54.8235 27.6660 55.9170 ;
        RECT 27.5320 54.8235 27.5580 55.9170 ;
        RECT 27.4240 54.8235 27.4500 55.9170 ;
        RECT 27.3160 54.8235 27.3420 55.9170 ;
        RECT 27.2080 54.8235 27.2340 55.9170 ;
        RECT 27.1000 54.8235 27.1260 55.9170 ;
        RECT 26.9920 54.8235 27.0180 55.9170 ;
        RECT 26.8840 54.8235 26.9100 55.9170 ;
        RECT 26.7760 54.8235 26.8020 55.9170 ;
        RECT 26.6680 54.8235 26.6940 55.9170 ;
        RECT 26.5600 54.8235 26.5860 55.9170 ;
        RECT 26.4520 54.8235 26.4780 55.9170 ;
        RECT 26.3440 54.8235 26.3700 55.9170 ;
        RECT 26.2360 54.8235 26.2620 55.9170 ;
        RECT 26.1280 54.8235 26.1540 55.9170 ;
        RECT 26.0200 54.8235 26.0460 55.9170 ;
        RECT 25.9120 54.8235 25.9380 55.9170 ;
        RECT 25.8040 54.8235 25.8300 55.9170 ;
        RECT 25.6960 54.8235 25.7220 55.9170 ;
        RECT 25.5880 54.8235 25.6140 55.9170 ;
        RECT 25.4800 54.8235 25.5060 55.9170 ;
        RECT 25.3720 54.8235 25.3980 55.9170 ;
        RECT 25.2640 54.8235 25.2900 55.9170 ;
        RECT 25.1560 54.8235 25.1820 55.9170 ;
        RECT 25.0480 54.8235 25.0740 55.9170 ;
        RECT 24.9400 54.8235 24.9660 55.9170 ;
        RECT 24.8320 54.8235 24.8580 55.9170 ;
        RECT 24.7240 54.8235 24.7500 55.9170 ;
        RECT 24.6160 54.8235 24.6420 55.9170 ;
        RECT 24.5080 54.8235 24.5340 55.9170 ;
        RECT 24.4000 54.8235 24.4260 55.9170 ;
        RECT 24.2920 54.8235 24.3180 55.9170 ;
        RECT 24.1840 54.8235 24.2100 55.9170 ;
        RECT 24.0760 54.8235 24.1020 55.9170 ;
        RECT 23.9680 54.8235 23.9940 55.9170 ;
        RECT 23.8600 54.8235 23.8860 55.9170 ;
        RECT 23.7520 54.8235 23.7780 55.9170 ;
        RECT 23.6440 54.8235 23.6700 55.9170 ;
        RECT 23.5360 54.8235 23.5620 55.9170 ;
        RECT 23.4280 54.8235 23.4540 55.9170 ;
        RECT 23.3200 54.8235 23.3460 55.9170 ;
        RECT 23.2120 54.8235 23.2380 55.9170 ;
        RECT 23.1040 54.8235 23.1300 55.9170 ;
        RECT 22.9960 54.8235 23.0220 55.9170 ;
        RECT 22.8880 54.8235 22.9140 55.9170 ;
        RECT 22.7800 54.8235 22.8060 55.9170 ;
        RECT 22.6720 54.8235 22.6980 55.9170 ;
        RECT 22.5640 54.8235 22.5900 55.9170 ;
        RECT 22.4560 54.8235 22.4820 55.9170 ;
        RECT 22.3480 54.8235 22.3740 55.9170 ;
        RECT 22.2400 54.8235 22.2660 55.9170 ;
        RECT 22.1320 54.8235 22.1580 55.9170 ;
        RECT 22.0240 54.8235 22.0500 55.9170 ;
        RECT 21.9160 54.8235 21.9420 55.9170 ;
        RECT 21.8080 54.8235 21.8340 55.9170 ;
        RECT 21.7000 54.8235 21.7260 55.9170 ;
        RECT 21.5920 54.8235 21.6180 55.9170 ;
        RECT 21.4840 54.8235 21.5100 55.9170 ;
        RECT 21.3760 54.8235 21.4020 55.9170 ;
        RECT 21.2680 54.8235 21.2940 55.9170 ;
        RECT 21.1600 54.8235 21.1860 55.9170 ;
        RECT 21.0520 54.8235 21.0780 55.9170 ;
        RECT 20.9440 54.8235 20.9700 55.9170 ;
        RECT 20.8360 54.8235 20.8620 55.9170 ;
        RECT 20.7280 54.8235 20.7540 55.9170 ;
        RECT 20.6200 54.8235 20.6460 55.9170 ;
        RECT 20.5120 54.8235 20.5380 55.9170 ;
        RECT 20.4040 54.8235 20.4300 55.9170 ;
        RECT 20.2960 54.8235 20.3220 55.9170 ;
        RECT 20.1880 54.8235 20.2140 55.9170 ;
        RECT 20.0800 54.8235 20.1060 55.9170 ;
        RECT 19.9720 54.8235 19.9980 55.9170 ;
        RECT 19.8640 54.8235 19.8900 55.9170 ;
        RECT 19.7560 54.8235 19.7820 55.9170 ;
        RECT 19.6480 54.8235 19.6740 55.9170 ;
        RECT 19.5400 54.8235 19.5660 55.9170 ;
        RECT 19.4320 54.8235 19.4580 55.9170 ;
        RECT 19.3240 54.8235 19.3500 55.9170 ;
        RECT 19.2160 54.8235 19.2420 55.9170 ;
        RECT 19.1080 54.8235 19.1340 55.9170 ;
        RECT 19.0000 54.8235 19.0260 55.9170 ;
        RECT 18.8920 54.8235 18.9180 55.9170 ;
        RECT 18.7840 54.8235 18.8100 55.9170 ;
        RECT 18.6760 54.8235 18.7020 55.9170 ;
        RECT 18.5680 54.8235 18.5940 55.9170 ;
        RECT 18.4600 54.8235 18.4860 55.9170 ;
        RECT 18.3520 54.8235 18.3780 55.9170 ;
        RECT 18.2440 54.8235 18.2700 55.9170 ;
        RECT 18.1360 54.8235 18.1620 55.9170 ;
        RECT 18.0280 54.8235 18.0540 55.9170 ;
        RECT 17.9200 54.8235 17.9460 55.9170 ;
        RECT 17.8120 54.8235 17.8380 55.9170 ;
        RECT 17.7040 54.8235 17.7300 55.9170 ;
        RECT 17.5960 54.8235 17.6220 55.9170 ;
        RECT 17.4880 54.8235 17.5140 55.9170 ;
        RECT 17.3800 54.8235 17.4060 55.9170 ;
        RECT 17.2720 54.8235 17.2980 55.9170 ;
        RECT 17.1640 54.8235 17.1900 55.9170 ;
        RECT 17.0560 54.8235 17.0820 55.9170 ;
        RECT 16.9480 54.8235 16.9740 55.9170 ;
        RECT 16.8400 54.8235 16.8660 55.9170 ;
        RECT 16.7320 54.8235 16.7580 55.9170 ;
        RECT 16.6240 54.8235 16.6500 55.9170 ;
        RECT 16.5160 54.8235 16.5420 55.9170 ;
        RECT 16.4080 54.8235 16.4340 55.9170 ;
        RECT 16.3000 54.8235 16.3260 55.9170 ;
        RECT 16.0870 54.8235 16.1640 55.9170 ;
        RECT 14.1940 54.8235 14.2710 55.9170 ;
        RECT 14.0320 54.8235 14.0580 55.9170 ;
        RECT 13.9240 54.8235 13.9500 55.9170 ;
        RECT 13.8160 54.8235 13.8420 55.9170 ;
        RECT 13.7080 54.8235 13.7340 55.9170 ;
        RECT 13.6000 54.8235 13.6260 55.9170 ;
        RECT 13.4920 54.8235 13.5180 55.9170 ;
        RECT 13.3840 54.8235 13.4100 55.9170 ;
        RECT 13.2760 54.8235 13.3020 55.9170 ;
        RECT 13.1680 54.8235 13.1940 55.9170 ;
        RECT 13.0600 54.8235 13.0860 55.9170 ;
        RECT 12.9520 54.8235 12.9780 55.9170 ;
        RECT 12.8440 54.8235 12.8700 55.9170 ;
        RECT 12.7360 54.8235 12.7620 55.9170 ;
        RECT 12.6280 54.8235 12.6540 55.9170 ;
        RECT 12.5200 54.8235 12.5460 55.9170 ;
        RECT 12.4120 54.8235 12.4380 55.9170 ;
        RECT 12.3040 54.8235 12.3300 55.9170 ;
        RECT 12.1960 54.8235 12.2220 55.9170 ;
        RECT 12.0880 54.8235 12.1140 55.9170 ;
        RECT 11.9800 54.8235 12.0060 55.9170 ;
        RECT 11.8720 54.8235 11.8980 55.9170 ;
        RECT 11.7640 54.8235 11.7900 55.9170 ;
        RECT 11.6560 54.8235 11.6820 55.9170 ;
        RECT 11.5480 54.8235 11.5740 55.9170 ;
        RECT 11.4400 54.8235 11.4660 55.9170 ;
        RECT 11.3320 54.8235 11.3580 55.9170 ;
        RECT 11.2240 54.8235 11.2500 55.9170 ;
        RECT 11.1160 54.8235 11.1420 55.9170 ;
        RECT 11.0080 54.8235 11.0340 55.9170 ;
        RECT 10.9000 54.8235 10.9260 55.9170 ;
        RECT 10.7920 54.8235 10.8180 55.9170 ;
        RECT 10.6840 54.8235 10.7100 55.9170 ;
        RECT 10.5760 54.8235 10.6020 55.9170 ;
        RECT 10.4680 54.8235 10.4940 55.9170 ;
        RECT 10.3600 54.8235 10.3860 55.9170 ;
        RECT 10.2520 54.8235 10.2780 55.9170 ;
        RECT 10.1440 54.8235 10.1700 55.9170 ;
        RECT 10.0360 54.8235 10.0620 55.9170 ;
        RECT 9.9280 54.8235 9.9540 55.9170 ;
        RECT 9.8200 54.8235 9.8460 55.9170 ;
        RECT 9.7120 54.8235 9.7380 55.9170 ;
        RECT 9.6040 54.8235 9.6300 55.9170 ;
        RECT 9.4960 54.8235 9.5220 55.9170 ;
        RECT 9.3880 54.8235 9.4140 55.9170 ;
        RECT 9.2800 54.8235 9.3060 55.9170 ;
        RECT 9.1720 54.8235 9.1980 55.9170 ;
        RECT 9.0640 54.8235 9.0900 55.9170 ;
        RECT 8.9560 54.8235 8.9820 55.9170 ;
        RECT 8.8480 54.8235 8.8740 55.9170 ;
        RECT 8.7400 54.8235 8.7660 55.9170 ;
        RECT 8.6320 54.8235 8.6580 55.9170 ;
        RECT 8.5240 54.8235 8.5500 55.9170 ;
        RECT 8.4160 54.8235 8.4420 55.9170 ;
        RECT 8.3080 54.8235 8.3340 55.9170 ;
        RECT 8.2000 54.8235 8.2260 55.9170 ;
        RECT 8.0920 54.8235 8.1180 55.9170 ;
        RECT 7.9840 54.8235 8.0100 55.9170 ;
        RECT 7.8760 54.8235 7.9020 55.9170 ;
        RECT 7.7680 54.8235 7.7940 55.9170 ;
        RECT 7.6600 54.8235 7.6860 55.9170 ;
        RECT 7.5520 54.8235 7.5780 55.9170 ;
        RECT 7.4440 54.8235 7.4700 55.9170 ;
        RECT 7.3360 54.8235 7.3620 55.9170 ;
        RECT 7.2280 54.8235 7.2540 55.9170 ;
        RECT 7.1200 54.8235 7.1460 55.9170 ;
        RECT 7.0120 54.8235 7.0380 55.9170 ;
        RECT 6.9040 54.8235 6.9300 55.9170 ;
        RECT 6.7960 54.8235 6.8220 55.9170 ;
        RECT 6.6880 54.8235 6.7140 55.9170 ;
        RECT 6.5800 54.8235 6.6060 55.9170 ;
        RECT 6.4720 54.8235 6.4980 55.9170 ;
        RECT 6.3640 54.8235 6.3900 55.9170 ;
        RECT 6.2560 54.8235 6.2820 55.9170 ;
        RECT 6.1480 54.8235 6.1740 55.9170 ;
        RECT 6.0400 54.8235 6.0660 55.9170 ;
        RECT 5.9320 54.8235 5.9580 55.9170 ;
        RECT 5.8240 54.8235 5.8500 55.9170 ;
        RECT 5.7160 54.8235 5.7420 55.9170 ;
        RECT 5.6080 54.8235 5.6340 55.9170 ;
        RECT 5.5000 54.8235 5.5260 55.9170 ;
        RECT 5.3920 54.8235 5.4180 55.9170 ;
        RECT 5.2840 54.8235 5.3100 55.9170 ;
        RECT 5.1760 54.8235 5.2020 55.9170 ;
        RECT 5.0680 54.8235 5.0940 55.9170 ;
        RECT 4.9600 54.8235 4.9860 55.9170 ;
        RECT 4.8520 54.8235 4.8780 55.9170 ;
        RECT 4.7440 54.8235 4.7700 55.9170 ;
        RECT 4.6360 54.8235 4.6620 55.9170 ;
        RECT 4.5280 54.8235 4.5540 55.9170 ;
        RECT 4.4200 54.8235 4.4460 55.9170 ;
        RECT 4.3120 54.8235 4.3380 55.9170 ;
        RECT 4.2040 54.8235 4.2300 55.9170 ;
        RECT 4.0960 54.8235 4.1220 55.9170 ;
        RECT 3.9880 54.8235 4.0140 55.9170 ;
        RECT 3.8800 54.8235 3.9060 55.9170 ;
        RECT 3.7720 54.8235 3.7980 55.9170 ;
        RECT 3.6640 54.8235 3.6900 55.9170 ;
        RECT 3.5560 54.8235 3.5820 55.9170 ;
        RECT 3.4480 54.8235 3.4740 55.9170 ;
        RECT 3.3400 54.8235 3.3660 55.9170 ;
        RECT 3.2320 54.8235 3.2580 55.9170 ;
        RECT 3.1240 54.8235 3.1500 55.9170 ;
        RECT 3.0160 54.8235 3.0420 55.9170 ;
        RECT 2.9080 54.8235 2.9340 55.9170 ;
        RECT 2.8000 54.8235 2.8260 55.9170 ;
        RECT 2.6920 54.8235 2.7180 55.9170 ;
        RECT 2.5840 54.8235 2.6100 55.9170 ;
        RECT 2.4760 54.8235 2.5020 55.9170 ;
        RECT 2.3680 54.8235 2.3940 55.9170 ;
        RECT 2.2600 54.8235 2.2860 55.9170 ;
        RECT 2.1520 54.8235 2.1780 55.9170 ;
        RECT 2.0440 54.8235 2.0700 55.9170 ;
        RECT 1.9360 54.8235 1.9620 55.9170 ;
        RECT 1.8280 54.8235 1.8540 55.9170 ;
        RECT 1.7200 54.8235 1.7460 55.9170 ;
        RECT 1.6120 54.8235 1.6380 55.9170 ;
        RECT 1.5040 54.8235 1.5300 55.9170 ;
        RECT 1.3960 54.8235 1.4220 55.9170 ;
        RECT 1.2880 54.8235 1.3140 55.9170 ;
        RECT 1.1800 54.8235 1.2060 55.9170 ;
        RECT 1.0720 54.8235 1.0980 55.9170 ;
        RECT 0.9640 54.8235 0.9900 55.9170 ;
        RECT 0.8560 54.8235 0.8820 55.9170 ;
        RECT 0.7480 54.8235 0.7740 55.9170 ;
        RECT 0.6400 54.8235 0.6660 55.9170 ;
        RECT 0.5320 54.8235 0.5580 55.9170 ;
        RECT 0.4240 54.8235 0.4500 55.9170 ;
        RECT 0.3160 54.8235 0.3420 55.9170 ;
        RECT 0.2080 54.8235 0.2340 55.9170 ;
        RECT 0.0050 54.8235 0.0900 55.9170 ;
        RECT 15.5530 55.9035 15.6810 56.9970 ;
        RECT 15.5390 56.5690 15.6810 56.8915 ;
        RECT 15.3190 56.2960 15.4530 56.9970 ;
        RECT 15.2960 56.6310 15.4530 56.8890 ;
        RECT 15.3190 55.9035 15.4170 56.9970 ;
        RECT 15.3190 56.0245 15.4310 56.2640 ;
        RECT 15.3190 55.9035 15.4530 55.9925 ;
        RECT 15.0940 56.3540 15.2280 56.9970 ;
        RECT 15.0940 55.9035 15.1920 56.9970 ;
        RECT 14.6770 55.9035 14.7600 56.9970 ;
        RECT 14.6770 55.9920 14.7740 56.9275 ;
        RECT 30.2680 55.9035 30.3530 56.9970 ;
        RECT 30.1240 55.9035 30.1500 56.9970 ;
        RECT 30.0160 55.9035 30.0420 56.9970 ;
        RECT 29.9080 55.9035 29.9340 56.9970 ;
        RECT 29.8000 55.9035 29.8260 56.9970 ;
        RECT 29.6920 55.9035 29.7180 56.9970 ;
        RECT 29.5840 55.9035 29.6100 56.9970 ;
        RECT 29.4760 55.9035 29.5020 56.9970 ;
        RECT 29.3680 55.9035 29.3940 56.9970 ;
        RECT 29.2600 55.9035 29.2860 56.9970 ;
        RECT 29.1520 55.9035 29.1780 56.9970 ;
        RECT 29.0440 55.9035 29.0700 56.9970 ;
        RECT 28.9360 55.9035 28.9620 56.9970 ;
        RECT 28.8280 55.9035 28.8540 56.9970 ;
        RECT 28.7200 55.9035 28.7460 56.9970 ;
        RECT 28.6120 55.9035 28.6380 56.9970 ;
        RECT 28.5040 55.9035 28.5300 56.9970 ;
        RECT 28.3960 55.9035 28.4220 56.9970 ;
        RECT 28.2880 55.9035 28.3140 56.9970 ;
        RECT 28.1800 55.9035 28.2060 56.9970 ;
        RECT 28.0720 55.9035 28.0980 56.9970 ;
        RECT 27.9640 55.9035 27.9900 56.9970 ;
        RECT 27.8560 55.9035 27.8820 56.9970 ;
        RECT 27.7480 55.9035 27.7740 56.9970 ;
        RECT 27.6400 55.9035 27.6660 56.9970 ;
        RECT 27.5320 55.9035 27.5580 56.9970 ;
        RECT 27.4240 55.9035 27.4500 56.9970 ;
        RECT 27.3160 55.9035 27.3420 56.9970 ;
        RECT 27.2080 55.9035 27.2340 56.9970 ;
        RECT 27.1000 55.9035 27.1260 56.9970 ;
        RECT 26.9920 55.9035 27.0180 56.9970 ;
        RECT 26.8840 55.9035 26.9100 56.9970 ;
        RECT 26.7760 55.9035 26.8020 56.9970 ;
        RECT 26.6680 55.9035 26.6940 56.9970 ;
        RECT 26.5600 55.9035 26.5860 56.9970 ;
        RECT 26.4520 55.9035 26.4780 56.9970 ;
        RECT 26.3440 55.9035 26.3700 56.9970 ;
        RECT 26.2360 55.9035 26.2620 56.9970 ;
        RECT 26.1280 55.9035 26.1540 56.9970 ;
        RECT 26.0200 55.9035 26.0460 56.9970 ;
        RECT 25.9120 55.9035 25.9380 56.9970 ;
        RECT 25.8040 55.9035 25.8300 56.9970 ;
        RECT 25.6960 55.9035 25.7220 56.9970 ;
        RECT 25.5880 55.9035 25.6140 56.9970 ;
        RECT 25.4800 55.9035 25.5060 56.9970 ;
        RECT 25.3720 55.9035 25.3980 56.9970 ;
        RECT 25.2640 55.9035 25.2900 56.9970 ;
        RECT 25.1560 55.9035 25.1820 56.9970 ;
        RECT 25.0480 55.9035 25.0740 56.9970 ;
        RECT 24.9400 55.9035 24.9660 56.9970 ;
        RECT 24.8320 55.9035 24.8580 56.9970 ;
        RECT 24.7240 55.9035 24.7500 56.9970 ;
        RECT 24.6160 55.9035 24.6420 56.9970 ;
        RECT 24.5080 55.9035 24.5340 56.9970 ;
        RECT 24.4000 55.9035 24.4260 56.9970 ;
        RECT 24.2920 55.9035 24.3180 56.9970 ;
        RECT 24.1840 55.9035 24.2100 56.9970 ;
        RECT 24.0760 55.9035 24.1020 56.9970 ;
        RECT 23.9680 55.9035 23.9940 56.9970 ;
        RECT 23.8600 55.9035 23.8860 56.9970 ;
        RECT 23.7520 55.9035 23.7780 56.9970 ;
        RECT 23.6440 55.9035 23.6700 56.9970 ;
        RECT 23.5360 55.9035 23.5620 56.9970 ;
        RECT 23.4280 55.9035 23.4540 56.9970 ;
        RECT 23.3200 55.9035 23.3460 56.9970 ;
        RECT 23.2120 55.9035 23.2380 56.9970 ;
        RECT 23.1040 55.9035 23.1300 56.9970 ;
        RECT 22.9960 55.9035 23.0220 56.9970 ;
        RECT 22.8880 55.9035 22.9140 56.9970 ;
        RECT 22.7800 55.9035 22.8060 56.9970 ;
        RECT 22.6720 55.9035 22.6980 56.9970 ;
        RECT 22.5640 55.9035 22.5900 56.9970 ;
        RECT 22.4560 55.9035 22.4820 56.9970 ;
        RECT 22.3480 55.9035 22.3740 56.9970 ;
        RECT 22.2400 55.9035 22.2660 56.9970 ;
        RECT 22.1320 55.9035 22.1580 56.9970 ;
        RECT 22.0240 55.9035 22.0500 56.9970 ;
        RECT 21.9160 55.9035 21.9420 56.9970 ;
        RECT 21.8080 55.9035 21.8340 56.9970 ;
        RECT 21.7000 55.9035 21.7260 56.9970 ;
        RECT 21.5920 55.9035 21.6180 56.9970 ;
        RECT 21.4840 55.9035 21.5100 56.9970 ;
        RECT 21.3760 55.9035 21.4020 56.9970 ;
        RECT 21.2680 55.9035 21.2940 56.9970 ;
        RECT 21.1600 55.9035 21.1860 56.9970 ;
        RECT 21.0520 55.9035 21.0780 56.9970 ;
        RECT 20.9440 55.9035 20.9700 56.9970 ;
        RECT 20.8360 55.9035 20.8620 56.9970 ;
        RECT 20.7280 55.9035 20.7540 56.9970 ;
        RECT 20.6200 55.9035 20.6460 56.9970 ;
        RECT 20.5120 55.9035 20.5380 56.9970 ;
        RECT 20.4040 55.9035 20.4300 56.9970 ;
        RECT 20.2960 55.9035 20.3220 56.9970 ;
        RECT 20.1880 55.9035 20.2140 56.9970 ;
        RECT 20.0800 55.9035 20.1060 56.9970 ;
        RECT 19.9720 55.9035 19.9980 56.9970 ;
        RECT 19.8640 55.9035 19.8900 56.9970 ;
        RECT 19.7560 55.9035 19.7820 56.9970 ;
        RECT 19.6480 55.9035 19.6740 56.9970 ;
        RECT 19.5400 55.9035 19.5660 56.9970 ;
        RECT 19.4320 55.9035 19.4580 56.9970 ;
        RECT 19.3240 55.9035 19.3500 56.9970 ;
        RECT 19.2160 55.9035 19.2420 56.9970 ;
        RECT 19.1080 55.9035 19.1340 56.9970 ;
        RECT 19.0000 55.9035 19.0260 56.9970 ;
        RECT 18.8920 55.9035 18.9180 56.9970 ;
        RECT 18.7840 55.9035 18.8100 56.9970 ;
        RECT 18.6760 55.9035 18.7020 56.9970 ;
        RECT 18.5680 55.9035 18.5940 56.9970 ;
        RECT 18.4600 55.9035 18.4860 56.9970 ;
        RECT 18.3520 55.9035 18.3780 56.9970 ;
        RECT 18.2440 55.9035 18.2700 56.9970 ;
        RECT 18.1360 55.9035 18.1620 56.9970 ;
        RECT 18.0280 55.9035 18.0540 56.9970 ;
        RECT 17.9200 55.9035 17.9460 56.9970 ;
        RECT 17.8120 55.9035 17.8380 56.9970 ;
        RECT 17.7040 55.9035 17.7300 56.9970 ;
        RECT 17.5960 55.9035 17.6220 56.9970 ;
        RECT 17.4880 55.9035 17.5140 56.9970 ;
        RECT 17.3800 55.9035 17.4060 56.9970 ;
        RECT 17.2720 55.9035 17.2980 56.9970 ;
        RECT 17.1640 55.9035 17.1900 56.9970 ;
        RECT 17.0560 55.9035 17.0820 56.9970 ;
        RECT 16.9480 55.9035 16.9740 56.9970 ;
        RECT 16.8400 55.9035 16.8660 56.9970 ;
        RECT 16.7320 55.9035 16.7580 56.9970 ;
        RECT 16.6240 55.9035 16.6500 56.9970 ;
        RECT 16.5160 55.9035 16.5420 56.9970 ;
        RECT 16.4080 55.9035 16.4340 56.9970 ;
        RECT 16.3000 55.9035 16.3260 56.9970 ;
        RECT 16.0870 55.9035 16.1640 56.9970 ;
        RECT 14.1940 55.9035 14.2710 56.9970 ;
        RECT 14.0320 55.9035 14.0580 56.9970 ;
        RECT 13.9240 55.9035 13.9500 56.9970 ;
        RECT 13.8160 55.9035 13.8420 56.9970 ;
        RECT 13.7080 55.9035 13.7340 56.9970 ;
        RECT 13.6000 55.9035 13.6260 56.9970 ;
        RECT 13.4920 55.9035 13.5180 56.9970 ;
        RECT 13.3840 55.9035 13.4100 56.9970 ;
        RECT 13.2760 55.9035 13.3020 56.9970 ;
        RECT 13.1680 55.9035 13.1940 56.9970 ;
        RECT 13.0600 55.9035 13.0860 56.9970 ;
        RECT 12.9520 55.9035 12.9780 56.9970 ;
        RECT 12.8440 55.9035 12.8700 56.9970 ;
        RECT 12.7360 55.9035 12.7620 56.9970 ;
        RECT 12.6280 55.9035 12.6540 56.9970 ;
        RECT 12.5200 55.9035 12.5460 56.9970 ;
        RECT 12.4120 55.9035 12.4380 56.9970 ;
        RECT 12.3040 55.9035 12.3300 56.9970 ;
        RECT 12.1960 55.9035 12.2220 56.9970 ;
        RECT 12.0880 55.9035 12.1140 56.9970 ;
        RECT 11.9800 55.9035 12.0060 56.9970 ;
        RECT 11.8720 55.9035 11.8980 56.9970 ;
        RECT 11.7640 55.9035 11.7900 56.9970 ;
        RECT 11.6560 55.9035 11.6820 56.9970 ;
        RECT 11.5480 55.9035 11.5740 56.9970 ;
        RECT 11.4400 55.9035 11.4660 56.9970 ;
        RECT 11.3320 55.9035 11.3580 56.9970 ;
        RECT 11.2240 55.9035 11.2500 56.9970 ;
        RECT 11.1160 55.9035 11.1420 56.9970 ;
        RECT 11.0080 55.9035 11.0340 56.9970 ;
        RECT 10.9000 55.9035 10.9260 56.9970 ;
        RECT 10.7920 55.9035 10.8180 56.9970 ;
        RECT 10.6840 55.9035 10.7100 56.9970 ;
        RECT 10.5760 55.9035 10.6020 56.9970 ;
        RECT 10.4680 55.9035 10.4940 56.9970 ;
        RECT 10.3600 55.9035 10.3860 56.9970 ;
        RECT 10.2520 55.9035 10.2780 56.9970 ;
        RECT 10.1440 55.9035 10.1700 56.9970 ;
        RECT 10.0360 55.9035 10.0620 56.9970 ;
        RECT 9.9280 55.9035 9.9540 56.9970 ;
        RECT 9.8200 55.9035 9.8460 56.9970 ;
        RECT 9.7120 55.9035 9.7380 56.9970 ;
        RECT 9.6040 55.9035 9.6300 56.9970 ;
        RECT 9.4960 55.9035 9.5220 56.9970 ;
        RECT 9.3880 55.9035 9.4140 56.9970 ;
        RECT 9.2800 55.9035 9.3060 56.9970 ;
        RECT 9.1720 55.9035 9.1980 56.9970 ;
        RECT 9.0640 55.9035 9.0900 56.9970 ;
        RECT 8.9560 55.9035 8.9820 56.9970 ;
        RECT 8.8480 55.9035 8.8740 56.9970 ;
        RECT 8.7400 55.9035 8.7660 56.9970 ;
        RECT 8.6320 55.9035 8.6580 56.9970 ;
        RECT 8.5240 55.9035 8.5500 56.9970 ;
        RECT 8.4160 55.9035 8.4420 56.9970 ;
        RECT 8.3080 55.9035 8.3340 56.9970 ;
        RECT 8.2000 55.9035 8.2260 56.9970 ;
        RECT 8.0920 55.9035 8.1180 56.9970 ;
        RECT 7.9840 55.9035 8.0100 56.9970 ;
        RECT 7.8760 55.9035 7.9020 56.9970 ;
        RECT 7.7680 55.9035 7.7940 56.9970 ;
        RECT 7.6600 55.9035 7.6860 56.9970 ;
        RECT 7.5520 55.9035 7.5780 56.9970 ;
        RECT 7.4440 55.9035 7.4700 56.9970 ;
        RECT 7.3360 55.9035 7.3620 56.9970 ;
        RECT 7.2280 55.9035 7.2540 56.9970 ;
        RECT 7.1200 55.9035 7.1460 56.9970 ;
        RECT 7.0120 55.9035 7.0380 56.9970 ;
        RECT 6.9040 55.9035 6.9300 56.9970 ;
        RECT 6.7960 55.9035 6.8220 56.9970 ;
        RECT 6.6880 55.9035 6.7140 56.9970 ;
        RECT 6.5800 55.9035 6.6060 56.9970 ;
        RECT 6.4720 55.9035 6.4980 56.9970 ;
        RECT 6.3640 55.9035 6.3900 56.9970 ;
        RECT 6.2560 55.9035 6.2820 56.9970 ;
        RECT 6.1480 55.9035 6.1740 56.9970 ;
        RECT 6.0400 55.9035 6.0660 56.9970 ;
        RECT 5.9320 55.9035 5.9580 56.9970 ;
        RECT 5.8240 55.9035 5.8500 56.9970 ;
        RECT 5.7160 55.9035 5.7420 56.9970 ;
        RECT 5.6080 55.9035 5.6340 56.9970 ;
        RECT 5.5000 55.9035 5.5260 56.9970 ;
        RECT 5.3920 55.9035 5.4180 56.9970 ;
        RECT 5.2840 55.9035 5.3100 56.9970 ;
        RECT 5.1760 55.9035 5.2020 56.9970 ;
        RECT 5.0680 55.9035 5.0940 56.9970 ;
        RECT 4.9600 55.9035 4.9860 56.9970 ;
        RECT 4.8520 55.9035 4.8780 56.9970 ;
        RECT 4.7440 55.9035 4.7700 56.9970 ;
        RECT 4.6360 55.9035 4.6620 56.9970 ;
        RECT 4.5280 55.9035 4.5540 56.9970 ;
        RECT 4.4200 55.9035 4.4460 56.9970 ;
        RECT 4.3120 55.9035 4.3380 56.9970 ;
        RECT 4.2040 55.9035 4.2300 56.9970 ;
        RECT 4.0960 55.9035 4.1220 56.9970 ;
        RECT 3.9880 55.9035 4.0140 56.9970 ;
        RECT 3.8800 55.9035 3.9060 56.9970 ;
        RECT 3.7720 55.9035 3.7980 56.9970 ;
        RECT 3.6640 55.9035 3.6900 56.9970 ;
        RECT 3.5560 55.9035 3.5820 56.9970 ;
        RECT 3.4480 55.9035 3.4740 56.9970 ;
        RECT 3.3400 55.9035 3.3660 56.9970 ;
        RECT 3.2320 55.9035 3.2580 56.9970 ;
        RECT 3.1240 55.9035 3.1500 56.9970 ;
        RECT 3.0160 55.9035 3.0420 56.9970 ;
        RECT 2.9080 55.9035 2.9340 56.9970 ;
        RECT 2.8000 55.9035 2.8260 56.9970 ;
        RECT 2.6920 55.9035 2.7180 56.9970 ;
        RECT 2.5840 55.9035 2.6100 56.9970 ;
        RECT 2.4760 55.9035 2.5020 56.9970 ;
        RECT 2.3680 55.9035 2.3940 56.9970 ;
        RECT 2.2600 55.9035 2.2860 56.9970 ;
        RECT 2.1520 55.9035 2.1780 56.9970 ;
        RECT 2.0440 55.9035 2.0700 56.9970 ;
        RECT 1.9360 55.9035 1.9620 56.9970 ;
        RECT 1.8280 55.9035 1.8540 56.9970 ;
        RECT 1.7200 55.9035 1.7460 56.9970 ;
        RECT 1.6120 55.9035 1.6380 56.9970 ;
        RECT 1.5040 55.9035 1.5300 56.9970 ;
        RECT 1.3960 55.9035 1.4220 56.9970 ;
        RECT 1.2880 55.9035 1.3140 56.9970 ;
        RECT 1.1800 55.9035 1.2060 56.9970 ;
        RECT 1.0720 55.9035 1.0980 56.9970 ;
        RECT 0.9640 55.9035 0.9900 56.9970 ;
        RECT 0.8560 55.9035 0.8820 56.9970 ;
        RECT 0.7480 55.9035 0.7740 56.9970 ;
        RECT 0.6400 55.9035 0.6660 56.9970 ;
        RECT 0.5320 55.9035 0.5580 56.9970 ;
        RECT 0.4240 55.9035 0.4500 56.9970 ;
        RECT 0.3160 55.9035 0.3420 56.9970 ;
        RECT 0.2080 55.9035 0.2340 56.9970 ;
        RECT 0.0050 55.9035 0.0900 56.9970 ;
        RECT 15.5530 56.9835 15.6810 58.0770 ;
        RECT 15.5390 57.6490 15.6810 57.9715 ;
        RECT 15.3190 57.3760 15.4530 58.0770 ;
        RECT 15.2960 57.7110 15.4530 57.9690 ;
        RECT 15.3190 56.9835 15.4170 58.0770 ;
        RECT 15.3190 57.1045 15.4310 57.3440 ;
        RECT 15.3190 56.9835 15.4530 57.0725 ;
        RECT 15.0940 57.4340 15.2280 58.0770 ;
        RECT 15.0940 56.9835 15.1920 58.0770 ;
        RECT 14.6770 56.9835 14.7600 58.0770 ;
        RECT 14.6770 57.0720 14.7740 58.0075 ;
        RECT 30.2680 56.9835 30.3530 58.0770 ;
        RECT 30.1240 56.9835 30.1500 58.0770 ;
        RECT 30.0160 56.9835 30.0420 58.0770 ;
        RECT 29.9080 56.9835 29.9340 58.0770 ;
        RECT 29.8000 56.9835 29.8260 58.0770 ;
        RECT 29.6920 56.9835 29.7180 58.0770 ;
        RECT 29.5840 56.9835 29.6100 58.0770 ;
        RECT 29.4760 56.9835 29.5020 58.0770 ;
        RECT 29.3680 56.9835 29.3940 58.0770 ;
        RECT 29.2600 56.9835 29.2860 58.0770 ;
        RECT 29.1520 56.9835 29.1780 58.0770 ;
        RECT 29.0440 56.9835 29.0700 58.0770 ;
        RECT 28.9360 56.9835 28.9620 58.0770 ;
        RECT 28.8280 56.9835 28.8540 58.0770 ;
        RECT 28.7200 56.9835 28.7460 58.0770 ;
        RECT 28.6120 56.9835 28.6380 58.0770 ;
        RECT 28.5040 56.9835 28.5300 58.0770 ;
        RECT 28.3960 56.9835 28.4220 58.0770 ;
        RECT 28.2880 56.9835 28.3140 58.0770 ;
        RECT 28.1800 56.9835 28.2060 58.0770 ;
        RECT 28.0720 56.9835 28.0980 58.0770 ;
        RECT 27.9640 56.9835 27.9900 58.0770 ;
        RECT 27.8560 56.9835 27.8820 58.0770 ;
        RECT 27.7480 56.9835 27.7740 58.0770 ;
        RECT 27.6400 56.9835 27.6660 58.0770 ;
        RECT 27.5320 56.9835 27.5580 58.0770 ;
        RECT 27.4240 56.9835 27.4500 58.0770 ;
        RECT 27.3160 56.9835 27.3420 58.0770 ;
        RECT 27.2080 56.9835 27.2340 58.0770 ;
        RECT 27.1000 56.9835 27.1260 58.0770 ;
        RECT 26.9920 56.9835 27.0180 58.0770 ;
        RECT 26.8840 56.9835 26.9100 58.0770 ;
        RECT 26.7760 56.9835 26.8020 58.0770 ;
        RECT 26.6680 56.9835 26.6940 58.0770 ;
        RECT 26.5600 56.9835 26.5860 58.0770 ;
        RECT 26.4520 56.9835 26.4780 58.0770 ;
        RECT 26.3440 56.9835 26.3700 58.0770 ;
        RECT 26.2360 56.9835 26.2620 58.0770 ;
        RECT 26.1280 56.9835 26.1540 58.0770 ;
        RECT 26.0200 56.9835 26.0460 58.0770 ;
        RECT 25.9120 56.9835 25.9380 58.0770 ;
        RECT 25.8040 56.9835 25.8300 58.0770 ;
        RECT 25.6960 56.9835 25.7220 58.0770 ;
        RECT 25.5880 56.9835 25.6140 58.0770 ;
        RECT 25.4800 56.9835 25.5060 58.0770 ;
        RECT 25.3720 56.9835 25.3980 58.0770 ;
        RECT 25.2640 56.9835 25.2900 58.0770 ;
        RECT 25.1560 56.9835 25.1820 58.0770 ;
        RECT 25.0480 56.9835 25.0740 58.0770 ;
        RECT 24.9400 56.9835 24.9660 58.0770 ;
        RECT 24.8320 56.9835 24.8580 58.0770 ;
        RECT 24.7240 56.9835 24.7500 58.0770 ;
        RECT 24.6160 56.9835 24.6420 58.0770 ;
        RECT 24.5080 56.9835 24.5340 58.0770 ;
        RECT 24.4000 56.9835 24.4260 58.0770 ;
        RECT 24.2920 56.9835 24.3180 58.0770 ;
        RECT 24.1840 56.9835 24.2100 58.0770 ;
        RECT 24.0760 56.9835 24.1020 58.0770 ;
        RECT 23.9680 56.9835 23.9940 58.0770 ;
        RECT 23.8600 56.9835 23.8860 58.0770 ;
        RECT 23.7520 56.9835 23.7780 58.0770 ;
        RECT 23.6440 56.9835 23.6700 58.0770 ;
        RECT 23.5360 56.9835 23.5620 58.0770 ;
        RECT 23.4280 56.9835 23.4540 58.0770 ;
        RECT 23.3200 56.9835 23.3460 58.0770 ;
        RECT 23.2120 56.9835 23.2380 58.0770 ;
        RECT 23.1040 56.9835 23.1300 58.0770 ;
        RECT 22.9960 56.9835 23.0220 58.0770 ;
        RECT 22.8880 56.9835 22.9140 58.0770 ;
        RECT 22.7800 56.9835 22.8060 58.0770 ;
        RECT 22.6720 56.9835 22.6980 58.0770 ;
        RECT 22.5640 56.9835 22.5900 58.0770 ;
        RECT 22.4560 56.9835 22.4820 58.0770 ;
        RECT 22.3480 56.9835 22.3740 58.0770 ;
        RECT 22.2400 56.9835 22.2660 58.0770 ;
        RECT 22.1320 56.9835 22.1580 58.0770 ;
        RECT 22.0240 56.9835 22.0500 58.0770 ;
        RECT 21.9160 56.9835 21.9420 58.0770 ;
        RECT 21.8080 56.9835 21.8340 58.0770 ;
        RECT 21.7000 56.9835 21.7260 58.0770 ;
        RECT 21.5920 56.9835 21.6180 58.0770 ;
        RECT 21.4840 56.9835 21.5100 58.0770 ;
        RECT 21.3760 56.9835 21.4020 58.0770 ;
        RECT 21.2680 56.9835 21.2940 58.0770 ;
        RECT 21.1600 56.9835 21.1860 58.0770 ;
        RECT 21.0520 56.9835 21.0780 58.0770 ;
        RECT 20.9440 56.9835 20.9700 58.0770 ;
        RECT 20.8360 56.9835 20.8620 58.0770 ;
        RECT 20.7280 56.9835 20.7540 58.0770 ;
        RECT 20.6200 56.9835 20.6460 58.0770 ;
        RECT 20.5120 56.9835 20.5380 58.0770 ;
        RECT 20.4040 56.9835 20.4300 58.0770 ;
        RECT 20.2960 56.9835 20.3220 58.0770 ;
        RECT 20.1880 56.9835 20.2140 58.0770 ;
        RECT 20.0800 56.9835 20.1060 58.0770 ;
        RECT 19.9720 56.9835 19.9980 58.0770 ;
        RECT 19.8640 56.9835 19.8900 58.0770 ;
        RECT 19.7560 56.9835 19.7820 58.0770 ;
        RECT 19.6480 56.9835 19.6740 58.0770 ;
        RECT 19.5400 56.9835 19.5660 58.0770 ;
        RECT 19.4320 56.9835 19.4580 58.0770 ;
        RECT 19.3240 56.9835 19.3500 58.0770 ;
        RECT 19.2160 56.9835 19.2420 58.0770 ;
        RECT 19.1080 56.9835 19.1340 58.0770 ;
        RECT 19.0000 56.9835 19.0260 58.0770 ;
        RECT 18.8920 56.9835 18.9180 58.0770 ;
        RECT 18.7840 56.9835 18.8100 58.0770 ;
        RECT 18.6760 56.9835 18.7020 58.0770 ;
        RECT 18.5680 56.9835 18.5940 58.0770 ;
        RECT 18.4600 56.9835 18.4860 58.0770 ;
        RECT 18.3520 56.9835 18.3780 58.0770 ;
        RECT 18.2440 56.9835 18.2700 58.0770 ;
        RECT 18.1360 56.9835 18.1620 58.0770 ;
        RECT 18.0280 56.9835 18.0540 58.0770 ;
        RECT 17.9200 56.9835 17.9460 58.0770 ;
        RECT 17.8120 56.9835 17.8380 58.0770 ;
        RECT 17.7040 56.9835 17.7300 58.0770 ;
        RECT 17.5960 56.9835 17.6220 58.0770 ;
        RECT 17.4880 56.9835 17.5140 58.0770 ;
        RECT 17.3800 56.9835 17.4060 58.0770 ;
        RECT 17.2720 56.9835 17.2980 58.0770 ;
        RECT 17.1640 56.9835 17.1900 58.0770 ;
        RECT 17.0560 56.9835 17.0820 58.0770 ;
        RECT 16.9480 56.9835 16.9740 58.0770 ;
        RECT 16.8400 56.9835 16.8660 58.0770 ;
        RECT 16.7320 56.9835 16.7580 58.0770 ;
        RECT 16.6240 56.9835 16.6500 58.0770 ;
        RECT 16.5160 56.9835 16.5420 58.0770 ;
        RECT 16.4080 56.9835 16.4340 58.0770 ;
        RECT 16.3000 56.9835 16.3260 58.0770 ;
        RECT 16.0870 56.9835 16.1640 58.0770 ;
        RECT 14.1940 56.9835 14.2710 58.0770 ;
        RECT 14.0320 56.9835 14.0580 58.0770 ;
        RECT 13.9240 56.9835 13.9500 58.0770 ;
        RECT 13.8160 56.9835 13.8420 58.0770 ;
        RECT 13.7080 56.9835 13.7340 58.0770 ;
        RECT 13.6000 56.9835 13.6260 58.0770 ;
        RECT 13.4920 56.9835 13.5180 58.0770 ;
        RECT 13.3840 56.9835 13.4100 58.0770 ;
        RECT 13.2760 56.9835 13.3020 58.0770 ;
        RECT 13.1680 56.9835 13.1940 58.0770 ;
        RECT 13.0600 56.9835 13.0860 58.0770 ;
        RECT 12.9520 56.9835 12.9780 58.0770 ;
        RECT 12.8440 56.9835 12.8700 58.0770 ;
        RECT 12.7360 56.9835 12.7620 58.0770 ;
        RECT 12.6280 56.9835 12.6540 58.0770 ;
        RECT 12.5200 56.9835 12.5460 58.0770 ;
        RECT 12.4120 56.9835 12.4380 58.0770 ;
        RECT 12.3040 56.9835 12.3300 58.0770 ;
        RECT 12.1960 56.9835 12.2220 58.0770 ;
        RECT 12.0880 56.9835 12.1140 58.0770 ;
        RECT 11.9800 56.9835 12.0060 58.0770 ;
        RECT 11.8720 56.9835 11.8980 58.0770 ;
        RECT 11.7640 56.9835 11.7900 58.0770 ;
        RECT 11.6560 56.9835 11.6820 58.0770 ;
        RECT 11.5480 56.9835 11.5740 58.0770 ;
        RECT 11.4400 56.9835 11.4660 58.0770 ;
        RECT 11.3320 56.9835 11.3580 58.0770 ;
        RECT 11.2240 56.9835 11.2500 58.0770 ;
        RECT 11.1160 56.9835 11.1420 58.0770 ;
        RECT 11.0080 56.9835 11.0340 58.0770 ;
        RECT 10.9000 56.9835 10.9260 58.0770 ;
        RECT 10.7920 56.9835 10.8180 58.0770 ;
        RECT 10.6840 56.9835 10.7100 58.0770 ;
        RECT 10.5760 56.9835 10.6020 58.0770 ;
        RECT 10.4680 56.9835 10.4940 58.0770 ;
        RECT 10.3600 56.9835 10.3860 58.0770 ;
        RECT 10.2520 56.9835 10.2780 58.0770 ;
        RECT 10.1440 56.9835 10.1700 58.0770 ;
        RECT 10.0360 56.9835 10.0620 58.0770 ;
        RECT 9.9280 56.9835 9.9540 58.0770 ;
        RECT 9.8200 56.9835 9.8460 58.0770 ;
        RECT 9.7120 56.9835 9.7380 58.0770 ;
        RECT 9.6040 56.9835 9.6300 58.0770 ;
        RECT 9.4960 56.9835 9.5220 58.0770 ;
        RECT 9.3880 56.9835 9.4140 58.0770 ;
        RECT 9.2800 56.9835 9.3060 58.0770 ;
        RECT 9.1720 56.9835 9.1980 58.0770 ;
        RECT 9.0640 56.9835 9.0900 58.0770 ;
        RECT 8.9560 56.9835 8.9820 58.0770 ;
        RECT 8.8480 56.9835 8.8740 58.0770 ;
        RECT 8.7400 56.9835 8.7660 58.0770 ;
        RECT 8.6320 56.9835 8.6580 58.0770 ;
        RECT 8.5240 56.9835 8.5500 58.0770 ;
        RECT 8.4160 56.9835 8.4420 58.0770 ;
        RECT 8.3080 56.9835 8.3340 58.0770 ;
        RECT 8.2000 56.9835 8.2260 58.0770 ;
        RECT 8.0920 56.9835 8.1180 58.0770 ;
        RECT 7.9840 56.9835 8.0100 58.0770 ;
        RECT 7.8760 56.9835 7.9020 58.0770 ;
        RECT 7.7680 56.9835 7.7940 58.0770 ;
        RECT 7.6600 56.9835 7.6860 58.0770 ;
        RECT 7.5520 56.9835 7.5780 58.0770 ;
        RECT 7.4440 56.9835 7.4700 58.0770 ;
        RECT 7.3360 56.9835 7.3620 58.0770 ;
        RECT 7.2280 56.9835 7.2540 58.0770 ;
        RECT 7.1200 56.9835 7.1460 58.0770 ;
        RECT 7.0120 56.9835 7.0380 58.0770 ;
        RECT 6.9040 56.9835 6.9300 58.0770 ;
        RECT 6.7960 56.9835 6.8220 58.0770 ;
        RECT 6.6880 56.9835 6.7140 58.0770 ;
        RECT 6.5800 56.9835 6.6060 58.0770 ;
        RECT 6.4720 56.9835 6.4980 58.0770 ;
        RECT 6.3640 56.9835 6.3900 58.0770 ;
        RECT 6.2560 56.9835 6.2820 58.0770 ;
        RECT 6.1480 56.9835 6.1740 58.0770 ;
        RECT 6.0400 56.9835 6.0660 58.0770 ;
        RECT 5.9320 56.9835 5.9580 58.0770 ;
        RECT 5.8240 56.9835 5.8500 58.0770 ;
        RECT 5.7160 56.9835 5.7420 58.0770 ;
        RECT 5.6080 56.9835 5.6340 58.0770 ;
        RECT 5.5000 56.9835 5.5260 58.0770 ;
        RECT 5.3920 56.9835 5.4180 58.0770 ;
        RECT 5.2840 56.9835 5.3100 58.0770 ;
        RECT 5.1760 56.9835 5.2020 58.0770 ;
        RECT 5.0680 56.9835 5.0940 58.0770 ;
        RECT 4.9600 56.9835 4.9860 58.0770 ;
        RECT 4.8520 56.9835 4.8780 58.0770 ;
        RECT 4.7440 56.9835 4.7700 58.0770 ;
        RECT 4.6360 56.9835 4.6620 58.0770 ;
        RECT 4.5280 56.9835 4.5540 58.0770 ;
        RECT 4.4200 56.9835 4.4460 58.0770 ;
        RECT 4.3120 56.9835 4.3380 58.0770 ;
        RECT 4.2040 56.9835 4.2300 58.0770 ;
        RECT 4.0960 56.9835 4.1220 58.0770 ;
        RECT 3.9880 56.9835 4.0140 58.0770 ;
        RECT 3.8800 56.9835 3.9060 58.0770 ;
        RECT 3.7720 56.9835 3.7980 58.0770 ;
        RECT 3.6640 56.9835 3.6900 58.0770 ;
        RECT 3.5560 56.9835 3.5820 58.0770 ;
        RECT 3.4480 56.9835 3.4740 58.0770 ;
        RECT 3.3400 56.9835 3.3660 58.0770 ;
        RECT 3.2320 56.9835 3.2580 58.0770 ;
        RECT 3.1240 56.9835 3.1500 58.0770 ;
        RECT 3.0160 56.9835 3.0420 58.0770 ;
        RECT 2.9080 56.9835 2.9340 58.0770 ;
        RECT 2.8000 56.9835 2.8260 58.0770 ;
        RECT 2.6920 56.9835 2.7180 58.0770 ;
        RECT 2.5840 56.9835 2.6100 58.0770 ;
        RECT 2.4760 56.9835 2.5020 58.0770 ;
        RECT 2.3680 56.9835 2.3940 58.0770 ;
        RECT 2.2600 56.9835 2.2860 58.0770 ;
        RECT 2.1520 56.9835 2.1780 58.0770 ;
        RECT 2.0440 56.9835 2.0700 58.0770 ;
        RECT 1.9360 56.9835 1.9620 58.0770 ;
        RECT 1.8280 56.9835 1.8540 58.0770 ;
        RECT 1.7200 56.9835 1.7460 58.0770 ;
        RECT 1.6120 56.9835 1.6380 58.0770 ;
        RECT 1.5040 56.9835 1.5300 58.0770 ;
        RECT 1.3960 56.9835 1.4220 58.0770 ;
        RECT 1.2880 56.9835 1.3140 58.0770 ;
        RECT 1.1800 56.9835 1.2060 58.0770 ;
        RECT 1.0720 56.9835 1.0980 58.0770 ;
        RECT 0.9640 56.9835 0.9900 58.0770 ;
        RECT 0.8560 56.9835 0.8820 58.0770 ;
        RECT 0.7480 56.9835 0.7740 58.0770 ;
        RECT 0.6400 56.9835 0.6660 58.0770 ;
        RECT 0.5320 56.9835 0.5580 58.0770 ;
        RECT 0.4240 56.9835 0.4500 58.0770 ;
        RECT 0.3160 56.9835 0.3420 58.0770 ;
        RECT 0.2080 56.9835 0.2340 58.0770 ;
        RECT 0.0050 56.9835 0.0900 58.0770 ;
        RECT 15.5530 58.0635 15.6810 59.1570 ;
        RECT 15.5390 58.7290 15.6810 59.0515 ;
        RECT 15.3190 58.4560 15.4530 59.1570 ;
        RECT 15.2960 58.7910 15.4530 59.0490 ;
        RECT 15.3190 58.0635 15.4170 59.1570 ;
        RECT 15.3190 58.1845 15.4310 58.4240 ;
        RECT 15.3190 58.0635 15.4530 58.1525 ;
        RECT 15.0940 58.5140 15.2280 59.1570 ;
        RECT 15.0940 58.0635 15.1920 59.1570 ;
        RECT 14.6770 58.0635 14.7600 59.1570 ;
        RECT 14.6770 58.1520 14.7740 59.0875 ;
        RECT 30.2680 58.0635 30.3530 59.1570 ;
        RECT 30.1240 58.0635 30.1500 59.1570 ;
        RECT 30.0160 58.0635 30.0420 59.1570 ;
        RECT 29.9080 58.0635 29.9340 59.1570 ;
        RECT 29.8000 58.0635 29.8260 59.1570 ;
        RECT 29.6920 58.0635 29.7180 59.1570 ;
        RECT 29.5840 58.0635 29.6100 59.1570 ;
        RECT 29.4760 58.0635 29.5020 59.1570 ;
        RECT 29.3680 58.0635 29.3940 59.1570 ;
        RECT 29.2600 58.0635 29.2860 59.1570 ;
        RECT 29.1520 58.0635 29.1780 59.1570 ;
        RECT 29.0440 58.0635 29.0700 59.1570 ;
        RECT 28.9360 58.0635 28.9620 59.1570 ;
        RECT 28.8280 58.0635 28.8540 59.1570 ;
        RECT 28.7200 58.0635 28.7460 59.1570 ;
        RECT 28.6120 58.0635 28.6380 59.1570 ;
        RECT 28.5040 58.0635 28.5300 59.1570 ;
        RECT 28.3960 58.0635 28.4220 59.1570 ;
        RECT 28.2880 58.0635 28.3140 59.1570 ;
        RECT 28.1800 58.0635 28.2060 59.1570 ;
        RECT 28.0720 58.0635 28.0980 59.1570 ;
        RECT 27.9640 58.0635 27.9900 59.1570 ;
        RECT 27.8560 58.0635 27.8820 59.1570 ;
        RECT 27.7480 58.0635 27.7740 59.1570 ;
        RECT 27.6400 58.0635 27.6660 59.1570 ;
        RECT 27.5320 58.0635 27.5580 59.1570 ;
        RECT 27.4240 58.0635 27.4500 59.1570 ;
        RECT 27.3160 58.0635 27.3420 59.1570 ;
        RECT 27.2080 58.0635 27.2340 59.1570 ;
        RECT 27.1000 58.0635 27.1260 59.1570 ;
        RECT 26.9920 58.0635 27.0180 59.1570 ;
        RECT 26.8840 58.0635 26.9100 59.1570 ;
        RECT 26.7760 58.0635 26.8020 59.1570 ;
        RECT 26.6680 58.0635 26.6940 59.1570 ;
        RECT 26.5600 58.0635 26.5860 59.1570 ;
        RECT 26.4520 58.0635 26.4780 59.1570 ;
        RECT 26.3440 58.0635 26.3700 59.1570 ;
        RECT 26.2360 58.0635 26.2620 59.1570 ;
        RECT 26.1280 58.0635 26.1540 59.1570 ;
        RECT 26.0200 58.0635 26.0460 59.1570 ;
        RECT 25.9120 58.0635 25.9380 59.1570 ;
        RECT 25.8040 58.0635 25.8300 59.1570 ;
        RECT 25.6960 58.0635 25.7220 59.1570 ;
        RECT 25.5880 58.0635 25.6140 59.1570 ;
        RECT 25.4800 58.0635 25.5060 59.1570 ;
        RECT 25.3720 58.0635 25.3980 59.1570 ;
        RECT 25.2640 58.0635 25.2900 59.1570 ;
        RECT 25.1560 58.0635 25.1820 59.1570 ;
        RECT 25.0480 58.0635 25.0740 59.1570 ;
        RECT 24.9400 58.0635 24.9660 59.1570 ;
        RECT 24.8320 58.0635 24.8580 59.1570 ;
        RECT 24.7240 58.0635 24.7500 59.1570 ;
        RECT 24.6160 58.0635 24.6420 59.1570 ;
        RECT 24.5080 58.0635 24.5340 59.1570 ;
        RECT 24.4000 58.0635 24.4260 59.1570 ;
        RECT 24.2920 58.0635 24.3180 59.1570 ;
        RECT 24.1840 58.0635 24.2100 59.1570 ;
        RECT 24.0760 58.0635 24.1020 59.1570 ;
        RECT 23.9680 58.0635 23.9940 59.1570 ;
        RECT 23.8600 58.0635 23.8860 59.1570 ;
        RECT 23.7520 58.0635 23.7780 59.1570 ;
        RECT 23.6440 58.0635 23.6700 59.1570 ;
        RECT 23.5360 58.0635 23.5620 59.1570 ;
        RECT 23.4280 58.0635 23.4540 59.1570 ;
        RECT 23.3200 58.0635 23.3460 59.1570 ;
        RECT 23.2120 58.0635 23.2380 59.1570 ;
        RECT 23.1040 58.0635 23.1300 59.1570 ;
        RECT 22.9960 58.0635 23.0220 59.1570 ;
        RECT 22.8880 58.0635 22.9140 59.1570 ;
        RECT 22.7800 58.0635 22.8060 59.1570 ;
        RECT 22.6720 58.0635 22.6980 59.1570 ;
        RECT 22.5640 58.0635 22.5900 59.1570 ;
        RECT 22.4560 58.0635 22.4820 59.1570 ;
        RECT 22.3480 58.0635 22.3740 59.1570 ;
        RECT 22.2400 58.0635 22.2660 59.1570 ;
        RECT 22.1320 58.0635 22.1580 59.1570 ;
        RECT 22.0240 58.0635 22.0500 59.1570 ;
        RECT 21.9160 58.0635 21.9420 59.1570 ;
        RECT 21.8080 58.0635 21.8340 59.1570 ;
        RECT 21.7000 58.0635 21.7260 59.1570 ;
        RECT 21.5920 58.0635 21.6180 59.1570 ;
        RECT 21.4840 58.0635 21.5100 59.1570 ;
        RECT 21.3760 58.0635 21.4020 59.1570 ;
        RECT 21.2680 58.0635 21.2940 59.1570 ;
        RECT 21.1600 58.0635 21.1860 59.1570 ;
        RECT 21.0520 58.0635 21.0780 59.1570 ;
        RECT 20.9440 58.0635 20.9700 59.1570 ;
        RECT 20.8360 58.0635 20.8620 59.1570 ;
        RECT 20.7280 58.0635 20.7540 59.1570 ;
        RECT 20.6200 58.0635 20.6460 59.1570 ;
        RECT 20.5120 58.0635 20.5380 59.1570 ;
        RECT 20.4040 58.0635 20.4300 59.1570 ;
        RECT 20.2960 58.0635 20.3220 59.1570 ;
        RECT 20.1880 58.0635 20.2140 59.1570 ;
        RECT 20.0800 58.0635 20.1060 59.1570 ;
        RECT 19.9720 58.0635 19.9980 59.1570 ;
        RECT 19.8640 58.0635 19.8900 59.1570 ;
        RECT 19.7560 58.0635 19.7820 59.1570 ;
        RECT 19.6480 58.0635 19.6740 59.1570 ;
        RECT 19.5400 58.0635 19.5660 59.1570 ;
        RECT 19.4320 58.0635 19.4580 59.1570 ;
        RECT 19.3240 58.0635 19.3500 59.1570 ;
        RECT 19.2160 58.0635 19.2420 59.1570 ;
        RECT 19.1080 58.0635 19.1340 59.1570 ;
        RECT 19.0000 58.0635 19.0260 59.1570 ;
        RECT 18.8920 58.0635 18.9180 59.1570 ;
        RECT 18.7840 58.0635 18.8100 59.1570 ;
        RECT 18.6760 58.0635 18.7020 59.1570 ;
        RECT 18.5680 58.0635 18.5940 59.1570 ;
        RECT 18.4600 58.0635 18.4860 59.1570 ;
        RECT 18.3520 58.0635 18.3780 59.1570 ;
        RECT 18.2440 58.0635 18.2700 59.1570 ;
        RECT 18.1360 58.0635 18.1620 59.1570 ;
        RECT 18.0280 58.0635 18.0540 59.1570 ;
        RECT 17.9200 58.0635 17.9460 59.1570 ;
        RECT 17.8120 58.0635 17.8380 59.1570 ;
        RECT 17.7040 58.0635 17.7300 59.1570 ;
        RECT 17.5960 58.0635 17.6220 59.1570 ;
        RECT 17.4880 58.0635 17.5140 59.1570 ;
        RECT 17.3800 58.0635 17.4060 59.1570 ;
        RECT 17.2720 58.0635 17.2980 59.1570 ;
        RECT 17.1640 58.0635 17.1900 59.1570 ;
        RECT 17.0560 58.0635 17.0820 59.1570 ;
        RECT 16.9480 58.0635 16.9740 59.1570 ;
        RECT 16.8400 58.0635 16.8660 59.1570 ;
        RECT 16.7320 58.0635 16.7580 59.1570 ;
        RECT 16.6240 58.0635 16.6500 59.1570 ;
        RECT 16.5160 58.0635 16.5420 59.1570 ;
        RECT 16.4080 58.0635 16.4340 59.1570 ;
        RECT 16.3000 58.0635 16.3260 59.1570 ;
        RECT 16.0870 58.0635 16.1640 59.1570 ;
        RECT 14.1940 58.0635 14.2710 59.1570 ;
        RECT 14.0320 58.0635 14.0580 59.1570 ;
        RECT 13.9240 58.0635 13.9500 59.1570 ;
        RECT 13.8160 58.0635 13.8420 59.1570 ;
        RECT 13.7080 58.0635 13.7340 59.1570 ;
        RECT 13.6000 58.0635 13.6260 59.1570 ;
        RECT 13.4920 58.0635 13.5180 59.1570 ;
        RECT 13.3840 58.0635 13.4100 59.1570 ;
        RECT 13.2760 58.0635 13.3020 59.1570 ;
        RECT 13.1680 58.0635 13.1940 59.1570 ;
        RECT 13.0600 58.0635 13.0860 59.1570 ;
        RECT 12.9520 58.0635 12.9780 59.1570 ;
        RECT 12.8440 58.0635 12.8700 59.1570 ;
        RECT 12.7360 58.0635 12.7620 59.1570 ;
        RECT 12.6280 58.0635 12.6540 59.1570 ;
        RECT 12.5200 58.0635 12.5460 59.1570 ;
        RECT 12.4120 58.0635 12.4380 59.1570 ;
        RECT 12.3040 58.0635 12.3300 59.1570 ;
        RECT 12.1960 58.0635 12.2220 59.1570 ;
        RECT 12.0880 58.0635 12.1140 59.1570 ;
        RECT 11.9800 58.0635 12.0060 59.1570 ;
        RECT 11.8720 58.0635 11.8980 59.1570 ;
        RECT 11.7640 58.0635 11.7900 59.1570 ;
        RECT 11.6560 58.0635 11.6820 59.1570 ;
        RECT 11.5480 58.0635 11.5740 59.1570 ;
        RECT 11.4400 58.0635 11.4660 59.1570 ;
        RECT 11.3320 58.0635 11.3580 59.1570 ;
        RECT 11.2240 58.0635 11.2500 59.1570 ;
        RECT 11.1160 58.0635 11.1420 59.1570 ;
        RECT 11.0080 58.0635 11.0340 59.1570 ;
        RECT 10.9000 58.0635 10.9260 59.1570 ;
        RECT 10.7920 58.0635 10.8180 59.1570 ;
        RECT 10.6840 58.0635 10.7100 59.1570 ;
        RECT 10.5760 58.0635 10.6020 59.1570 ;
        RECT 10.4680 58.0635 10.4940 59.1570 ;
        RECT 10.3600 58.0635 10.3860 59.1570 ;
        RECT 10.2520 58.0635 10.2780 59.1570 ;
        RECT 10.1440 58.0635 10.1700 59.1570 ;
        RECT 10.0360 58.0635 10.0620 59.1570 ;
        RECT 9.9280 58.0635 9.9540 59.1570 ;
        RECT 9.8200 58.0635 9.8460 59.1570 ;
        RECT 9.7120 58.0635 9.7380 59.1570 ;
        RECT 9.6040 58.0635 9.6300 59.1570 ;
        RECT 9.4960 58.0635 9.5220 59.1570 ;
        RECT 9.3880 58.0635 9.4140 59.1570 ;
        RECT 9.2800 58.0635 9.3060 59.1570 ;
        RECT 9.1720 58.0635 9.1980 59.1570 ;
        RECT 9.0640 58.0635 9.0900 59.1570 ;
        RECT 8.9560 58.0635 8.9820 59.1570 ;
        RECT 8.8480 58.0635 8.8740 59.1570 ;
        RECT 8.7400 58.0635 8.7660 59.1570 ;
        RECT 8.6320 58.0635 8.6580 59.1570 ;
        RECT 8.5240 58.0635 8.5500 59.1570 ;
        RECT 8.4160 58.0635 8.4420 59.1570 ;
        RECT 8.3080 58.0635 8.3340 59.1570 ;
        RECT 8.2000 58.0635 8.2260 59.1570 ;
        RECT 8.0920 58.0635 8.1180 59.1570 ;
        RECT 7.9840 58.0635 8.0100 59.1570 ;
        RECT 7.8760 58.0635 7.9020 59.1570 ;
        RECT 7.7680 58.0635 7.7940 59.1570 ;
        RECT 7.6600 58.0635 7.6860 59.1570 ;
        RECT 7.5520 58.0635 7.5780 59.1570 ;
        RECT 7.4440 58.0635 7.4700 59.1570 ;
        RECT 7.3360 58.0635 7.3620 59.1570 ;
        RECT 7.2280 58.0635 7.2540 59.1570 ;
        RECT 7.1200 58.0635 7.1460 59.1570 ;
        RECT 7.0120 58.0635 7.0380 59.1570 ;
        RECT 6.9040 58.0635 6.9300 59.1570 ;
        RECT 6.7960 58.0635 6.8220 59.1570 ;
        RECT 6.6880 58.0635 6.7140 59.1570 ;
        RECT 6.5800 58.0635 6.6060 59.1570 ;
        RECT 6.4720 58.0635 6.4980 59.1570 ;
        RECT 6.3640 58.0635 6.3900 59.1570 ;
        RECT 6.2560 58.0635 6.2820 59.1570 ;
        RECT 6.1480 58.0635 6.1740 59.1570 ;
        RECT 6.0400 58.0635 6.0660 59.1570 ;
        RECT 5.9320 58.0635 5.9580 59.1570 ;
        RECT 5.8240 58.0635 5.8500 59.1570 ;
        RECT 5.7160 58.0635 5.7420 59.1570 ;
        RECT 5.6080 58.0635 5.6340 59.1570 ;
        RECT 5.5000 58.0635 5.5260 59.1570 ;
        RECT 5.3920 58.0635 5.4180 59.1570 ;
        RECT 5.2840 58.0635 5.3100 59.1570 ;
        RECT 5.1760 58.0635 5.2020 59.1570 ;
        RECT 5.0680 58.0635 5.0940 59.1570 ;
        RECT 4.9600 58.0635 4.9860 59.1570 ;
        RECT 4.8520 58.0635 4.8780 59.1570 ;
        RECT 4.7440 58.0635 4.7700 59.1570 ;
        RECT 4.6360 58.0635 4.6620 59.1570 ;
        RECT 4.5280 58.0635 4.5540 59.1570 ;
        RECT 4.4200 58.0635 4.4460 59.1570 ;
        RECT 4.3120 58.0635 4.3380 59.1570 ;
        RECT 4.2040 58.0635 4.2300 59.1570 ;
        RECT 4.0960 58.0635 4.1220 59.1570 ;
        RECT 3.9880 58.0635 4.0140 59.1570 ;
        RECT 3.8800 58.0635 3.9060 59.1570 ;
        RECT 3.7720 58.0635 3.7980 59.1570 ;
        RECT 3.6640 58.0635 3.6900 59.1570 ;
        RECT 3.5560 58.0635 3.5820 59.1570 ;
        RECT 3.4480 58.0635 3.4740 59.1570 ;
        RECT 3.3400 58.0635 3.3660 59.1570 ;
        RECT 3.2320 58.0635 3.2580 59.1570 ;
        RECT 3.1240 58.0635 3.1500 59.1570 ;
        RECT 3.0160 58.0635 3.0420 59.1570 ;
        RECT 2.9080 58.0635 2.9340 59.1570 ;
        RECT 2.8000 58.0635 2.8260 59.1570 ;
        RECT 2.6920 58.0635 2.7180 59.1570 ;
        RECT 2.5840 58.0635 2.6100 59.1570 ;
        RECT 2.4760 58.0635 2.5020 59.1570 ;
        RECT 2.3680 58.0635 2.3940 59.1570 ;
        RECT 2.2600 58.0635 2.2860 59.1570 ;
        RECT 2.1520 58.0635 2.1780 59.1570 ;
        RECT 2.0440 58.0635 2.0700 59.1570 ;
        RECT 1.9360 58.0635 1.9620 59.1570 ;
        RECT 1.8280 58.0635 1.8540 59.1570 ;
        RECT 1.7200 58.0635 1.7460 59.1570 ;
        RECT 1.6120 58.0635 1.6380 59.1570 ;
        RECT 1.5040 58.0635 1.5300 59.1570 ;
        RECT 1.3960 58.0635 1.4220 59.1570 ;
        RECT 1.2880 58.0635 1.3140 59.1570 ;
        RECT 1.1800 58.0635 1.2060 59.1570 ;
        RECT 1.0720 58.0635 1.0980 59.1570 ;
        RECT 0.9640 58.0635 0.9900 59.1570 ;
        RECT 0.8560 58.0635 0.8820 59.1570 ;
        RECT 0.7480 58.0635 0.7740 59.1570 ;
        RECT 0.6400 58.0635 0.6660 59.1570 ;
        RECT 0.5320 58.0635 0.5580 59.1570 ;
        RECT 0.4240 58.0635 0.4500 59.1570 ;
        RECT 0.3160 58.0635 0.3420 59.1570 ;
        RECT 0.2080 58.0635 0.2340 59.1570 ;
        RECT 0.0050 58.0635 0.0900 59.1570 ;
        RECT 15.5530 59.1435 15.6810 60.2370 ;
        RECT 15.5390 59.8090 15.6810 60.1315 ;
        RECT 15.3190 59.5360 15.4530 60.2370 ;
        RECT 15.2960 59.8710 15.4530 60.1290 ;
        RECT 15.3190 59.1435 15.4170 60.2370 ;
        RECT 15.3190 59.2645 15.4310 59.5040 ;
        RECT 15.3190 59.1435 15.4530 59.2325 ;
        RECT 15.0940 59.5940 15.2280 60.2370 ;
        RECT 15.0940 59.1435 15.1920 60.2370 ;
        RECT 14.6770 59.1435 14.7600 60.2370 ;
        RECT 14.6770 59.2320 14.7740 60.1675 ;
        RECT 30.2680 59.1435 30.3530 60.2370 ;
        RECT 30.1240 59.1435 30.1500 60.2370 ;
        RECT 30.0160 59.1435 30.0420 60.2370 ;
        RECT 29.9080 59.1435 29.9340 60.2370 ;
        RECT 29.8000 59.1435 29.8260 60.2370 ;
        RECT 29.6920 59.1435 29.7180 60.2370 ;
        RECT 29.5840 59.1435 29.6100 60.2370 ;
        RECT 29.4760 59.1435 29.5020 60.2370 ;
        RECT 29.3680 59.1435 29.3940 60.2370 ;
        RECT 29.2600 59.1435 29.2860 60.2370 ;
        RECT 29.1520 59.1435 29.1780 60.2370 ;
        RECT 29.0440 59.1435 29.0700 60.2370 ;
        RECT 28.9360 59.1435 28.9620 60.2370 ;
        RECT 28.8280 59.1435 28.8540 60.2370 ;
        RECT 28.7200 59.1435 28.7460 60.2370 ;
        RECT 28.6120 59.1435 28.6380 60.2370 ;
        RECT 28.5040 59.1435 28.5300 60.2370 ;
        RECT 28.3960 59.1435 28.4220 60.2370 ;
        RECT 28.2880 59.1435 28.3140 60.2370 ;
        RECT 28.1800 59.1435 28.2060 60.2370 ;
        RECT 28.0720 59.1435 28.0980 60.2370 ;
        RECT 27.9640 59.1435 27.9900 60.2370 ;
        RECT 27.8560 59.1435 27.8820 60.2370 ;
        RECT 27.7480 59.1435 27.7740 60.2370 ;
        RECT 27.6400 59.1435 27.6660 60.2370 ;
        RECT 27.5320 59.1435 27.5580 60.2370 ;
        RECT 27.4240 59.1435 27.4500 60.2370 ;
        RECT 27.3160 59.1435 27.3420 60.2370 ;
        RECT 27.2080 59.1435 27.2340 60.2370 ;
        RECT 27.1000 59.1435 27.1260 60.2370 ;
        RECT 26.9920 59.1435 27.0180 60.2370 ;
        RECT 26.8840 59.1435 26.9100 60.2370 ;
        RECT 26.7760 59.1435 26.8020 60.2370 ;
        RECT 26.6680 59.1435 26.6940 60.2370 ;
        RECT 26.5600 59.1435 26.5860 60.2370 ;
        RECT 26.4520 59.1435 26.4780 60.2370 ;
        RECT 26.3440 59.1435 26.3700 60.2370 ;
        RECT 26.2360 59.1435 26.2620 60.2370 ;
        RECT 26.1280 59.1435 26.1540 60.2370 ;
        RECT 26.0200 59.1435 26.0460 60.2370 ;
        RECT 25.9120 59.1435 25.9380 60.2370 ;
        RECT 25.8040 59.1435 25.8300 60.2370 ;
        RECT 25.6960 59.1435 25.7220 60.2370 ;
        RECT 25.5880 59.1435 25.6140 60.2370 ;
        RECT 25.4800 59.1435 25.5060 60.2370 ;
        RECT 25.3720 59.1435 25.3980 60.2370 ;
        RECT 25.2640 59.1435 25.2900 60.2370 ;
        RECT 25.1560 59.1435 25.1820 60.2370 ;
        RECT 25.0480 59.1435 25.0740 60.2370 ;
        RECT 24.9400 59.1435 24.9660 60.2370 ;
        RECT 24.8320 59.1435 24.8580 60.2370 ;
        RECT 24.7240 59.1435 24.7500 60.2370 ;
        RECT 24.6160 59.1435 24.6420 60.2370 ;
        RECT 24.5080 59.1435 24.5340 60.2370 ;
        RECT 24.4000 59.1435 24.4260 60.2370 ;
        RECT 24.2920 59.1435 24.3180 60.2370 ;
        RECT 24.1840 59.1435 24.2100 60.2370 ;
        RECT 24.0760 59.1435 24.1020 60.2370 ;
        RECT 23.9680 59.1435 23.9940 60.2370 ;
        RECT 23.8600 59.1435 23.8860 60.2370 ;
        RECT 23.7520 59.1435 23.7780 60.2370 ;
        RECT 23.6440 59.1435 23.6700 60.2370 ;
        RECT 23.5360 59.1435 23.5620 60.2370 ;
        RECT 23.4280 59.1435 23.4540 60.2370 ;
        RECT 23.3200 59.1435 23.3460 60.2370 ;
        RECT 23.2120 59.1435 23.2380 60.2370 ;
        RECT 23.1040 59.1435 23.1300 60.2370 ;
        RECT 22.9960 59.1435 23.0220 60.2370 ;
        RECT 22.8880 59.1435 22.9140 60.2370 ;
        RECT 22.7800 59.1435 22.8060 60.2370 ;
        RECT 22.6720 59.1435 22.6980 60.2370 ;
        RECT 22.5640 59.1435 22.5900 60.2370 ;
        RECT 22.4560 59.1435 22.4820 60.2370 ;
        RECT 22.3480 59.1435 22.3740 60.2370 ;
        RECT 22.2400 59.1435 22.2660 60.2370 ;
        RECT 22.1320 59.1435 22.1580 60.2370 ;
        RECT 22.0240 59.1435 22.0500 60.2370 ;
        RECT 21.9160 59.1435 21.9420 60.2370 ;
        RECT 21.8080 59.1435 21.8340 60.2370 ;
        RECT 21.7000 59.1435 21.7260 60.2370 ;
        RECT 21.5920 59.1435 21.6180 60.2370 ;
        RECT 21.4840 59.1435 21.5100 60.2370 ;
        RECT 21.3760 59.1435 21.4020 60.2370 ;
        RECT 21.2680 59.1435 21.2940 60.2370 ;
        RECT 21.1600 59.1435 21.1860 60.2370 ;
        RECT 21.0520 59.1435 21.0780 60.2370 ;
        RECT 20.9440 59.1435 20.9700 60.2370 ;
        RECT 20.8360 59.1435 20.8620 60.2370 ;
        RECT 20.7280 59.1435 20.7540 60.2370 ;
        RECT 20.6200 59.1435 20.6460 60.2370 ;
        RECT 20.5120 59.1435 20.5380 60.2370 ;
        RECT 20.4040 59.1435 20.4300 60.2370 ;
        RECT 20.2960 59.1435 20.3220 60.2370 ;
        RECT 20.1880 59.1435 20.2140 60.2370 ;
        RECT 20.0800 59.1435 20.1060 60.2370 ;
        RECT 19.9720 59.1435 19.9980 60.2370 ;
        RECT 19.8640 59.1435 19.8900 60.2370 ;
        RECT 19.7560 59.1435 19.7820 60.2370 ;
        RECT 19.6480 59.1435 19.6740 60.2370 ;
        RECT 19.5400 59.1435 19.5660 60.2370 ;
        RECT 19.4320 59.1435 19.4580 60.2370 ;
        RECT 19.3240 59.1435 19.3500 60.2370 ;
        RECT 19.2160 59.1435 19.2420 60.2370 ;
        RECT 19.1080 59.1435 19.1340 60.2370 ;
        RECT 19.0000 59.1435 19.0260 60.2370 ;
        RECT 18.8920 59.1435 18.9180 60.2370 ;
        RECT 18.7840 59.1435 18.8100 60.2370 ;
        RECT 18.6760 59.1435 18.7020 60.2370 ;
        RECT 18.5680 59.1435 18.5940 60.2370 ;
        RECT 18.4600 59.1435 18.4860 60.2370 ;
        RECT 18.3520 59.1435 18.3780 60.2370 ;
        RECT 18.2440 59.1435 18.2700 60.2370 ;
        RECT 18.1360 59.1435 18.1620 60.2370 ;
        RECT 18.0280 59.1435 18.0540 60.2370 ;
        RECT 17.9200 59.1435 17.9460 60.2370 ;
        RECT 17.8120 59.1435 17.8380 60.2370 ;
        RECT 17.7040 59.1435 17.7300 60.2370 ;
        RECT 17.5960 59.1435 17.6220 60.2370 ;
        RECT 17.4880 59.1435 17.5140 60.2370 ;
        RECT 17.3800 59.1435 17.4060 60.2370 ;
        RECT 17.2720 59.1435 17.2980 60.2370 ;
        RECT 17.1640 59.1435 17.1900 60.2370 ;
        RECT 17.0560 59.1435 17.0820 60.2370 ;
        RECT 16.9480 59.1435 16.9740 60.2370 ;
        RECT 16.8400 59.1435 16.8660 60.2370 ;
        RECT 16.7320 59.1435 16.7580 60.2370 ;
        RECT 16.6240 59.1435 16.6500 60.2370 ;
        RECT 16.5160 59.1435 16.5420 60.2370 ;
        RECT 16.4080 59.1435 16.4340 60.2370 ;
        RECT 16.3000 59.1435 16.3260 60.2370 ;
        RECT 16.0870 59.1435 16.1640 60.2370 ;
        RECT 14.1940 59.1435 14.2710 60.2370 ;
        RECT 14.0320 59.1435 14.0580 60.2370 ;
        RECT 13.9240 59.1435 13.9500 60.2370 ;
        RECT 13.8160 59.1435 13.8420 60.2370 ;
        RECT 13.7080 59.1435 13.7340 60.2370 ;
        RECT 13.6000 59.1435 13.6260 60.2370 ;
        RECT 13.4920 59.1435 13.5180 60.2370 ;
        RECT 13.3840 59.1435 13.4100 60.2370 ;
        RECT 13.2760 59.1435 13.3020 60.2370 ;
        RECT 13.1680 59.1435 13.1940 60.2370 ;
        RECT 13.0600 59.1435 13.0860 60.2370 ;
        RECT 12.9520 59.1435 12.9780 60.2370 ;
        RECT 12.8440 59.1435 12.8700 60.2370 ;
        RECT 12.7360 59.1435 12.7620 60.2370 ;
        RECT 12.6280 59.1435 12.6540 60.2370 ;
        RECT 12.5200 59.1435 12.5460 60.2370 ;
        RECT 12.4120 59.1435 12.4380 60.2370 ;
        RECT 12.3040 59.1435 12.3300 60.2370 ;
        RECT 12.1960 59.1435 12.2220 60.2370 ;
        RECT 12.0880 59.1435 12.1140 60.2370 ;
        RECT 11.9800 59.1435 12.0060 60.2370 ;
        RECT 11.8720 59.1435 11.8980 60.2370 ;
        RECT 11.7640 59.1435 11.7900 60.2370 ;
        RECT 11.6560 59.1435 11.6820 60.2370 ;
        RECT 11.5480 59.1435 11.5740 60.2370 ;
        RECT 11.4400 59.1435 11.4660 60.2370 ;
        RECT 11.3320 59.1435 11.3580 60.2370 ;
        RECT 11.2240 59.1435 11.2500 60.2370 ;
        RECT 11.1160 59.1435 11.1420 60.2370 ;
        RECT 11.0080 59.1435 11.0340 60.2370 ;
        RECT 10.9000 59.1435 10.9260 60.2370 ;
        RECT 10.7920 59.1435 10.8180 60.2370 ;
        RECT 10.6840 59.1435 10.7100 60.2370 ;
        RECT 10.5760 59.1435 10.6020 60.2370 ;
        RECT 10.4680 59.1435 10.4940 60.2370 ;
        RECT 10.3600 59.1435 10.3860 60.2370 ;
        RECT 10.2520 59.1435 10.2780 60.2370 ;
        RECT 10.1440 59.1435 10.1700 60.2370 ;
        RECT 10.0360 59.1435 10.0620 60.2370 ;
        RECT 9.9280 59.1435 9.9540 60.2370 ;
        RECT 9.8200 59.1435 9.8460 60.2370 ;
        RECT 9.7120 59.1435 9.7380 60.2370 ;
        RECT 9.6040 59.1435 9.6300 60.2370 ;
        RECT 9.4960 59.1435 9.5220 60.2370 ;
        RECT 9.3880 59.1435 9.4140 60.2370 ;
        RECT 9.2800 59.1435 9.3060 60.2370 ;
        RECT 9.1720 59.1435 9.1980 60.2370 ;
        RECT 9.0640 59.1435 9.0900 60.2370 ;
        RECT 8.9560 59.1435 8.9820 60.2370 ;
        RECT 8.8480 59.1435 8.8740 60.2370 ;
        RECT 8.7400 59.1435 8.7660 60.2370 ;
        RECT 8.6320 59.1435 8.6580 60.2370 ;
        RECT 8.5240 59.1435 8.5500 60.2370 ;
        RECT 8.4160 59.1435 8.4420 60.2370 ;
        RECT 8.3080 59.1435 8.3340 60.2370 ;
        RECT 8.2000 59.1435 8.2260 60.2370 ;
        RECT 8.0920 59.1435 8.1180 60.2370 ;
        RECT 7.9840 59.1435 8.0100 60.2370 ;
        RECT 7.8760 59.1435 7.9020 60.2370 ;
        RECT 7.7680 59.1435 7.7940 60.2370 ;
        RECT 7.6600 59.1435 7.6860 60.2370 ;
        RECT 7.5520 59.1435 7.5780 60.2370 ;
        RECT 7.4440 59.1435 7.4700 60.2370 ;
        RECT 7.3360 59.1435 7.3620 60.2370 ;
        RECT 7.2280 59.1435 7.2540 60.2370 ;
        RECT 7.1200 59.1435 7.1460 60.2370 ;
        RECT 7.0120 59.1435 7.0380 60.2370 ;
        RECT 6.9040 59.1435 6.9300 60.2370 ;
        RECT 6.7960 59.1435 6.8220 60.2370 ;
        RECT 6.6880 59.1435 6.7140 60.2370 ;
        RECT 6.5800 59.1435 6.6060 60.2370 ;
        RECT 6.4720 59.1435 6.4980 60.2370 ;
        RECT 6.3640 59.1435 6.3900 60.2370 ;
        RECT 6.2560 59.1435 6.2820 60.2370 ;
        RECT 6.1480 59.1435 6.1740 60.2370 ;
        RECT 6.0400 59.1435 6.0660 60.2370 ;
        RECT 5.9320 59.1435 5.9580 60.2370 ;
        RECT 5.8240 59.1435 5.8500 60.2370 ;
        RECT 5.7160 59.1435 5.7420 60.2370 ;
        RECT 5.6080 59.1435 5.6340 60.2370 ;
        RECT 5.5000 59.1435 5.5260 60.2370 ;
        RECT 5.3920 59.1435 5.4180 60.2370 ;
        RECT 5.2840 59.1435 5.3100 60.2370 ;
        RECT 5.1760 59.1435 5.2020 60.2370 ;
        RECT 5.0680 59.1435 5.0940 60.2370 ;
        RECT 4.9600 59.1435 4.9860 60.2370 ;
        RECT 4.8520 59.1435 4.8780 60.2370 ;
        RECT 4.7440 59.1435 4.7700 60.2370 ;
        RECT 4.6360 59.1435 4.6620 60.2370 ;
        RECT 4.5280 59.1435 4.5540 60.2370 ;
        RECT 4.4200 59.1435 4.4460 60.2370 ;
        RECT 4.3120 59.1435 4.3380 60.2370 ;
        RECT 4.2040 59.1435 4.2300 60.2370 ;
        RECT 4.0960 59.1435 4.1220 60.2370 ;
        RECT 3.9880 59.1435 4.0140 60.2370 ;
        RECT 3.8800 59.1435 3.9060 60.2370 ;
        RECT 3.7720 59.1435 3.7980 60.2370 ;
        RECT 3.6640 59.1435 3.6900 60.2370 ;
        RECT 3.5560 59.1435 3.5820 60.2370 ;
        RECT 3.4480 59.1435 3.4740 60.2370 ;
        RECT 3.3400 59.1435 3.3660 60.2370 ;
        RECT 3.2320 59.1435 3.2580 60.2370 ;
        RECT 3.1240 59.1435 3.1500 60.2370 ;
        RECT 3.0160 59.1435 3.0420 60.2370 ;
        RECT 2.9080 59.1435 2.9340 60.2370 ;
        RECT 2.8000 59.1435 2.8260 60.2370 ;
        RECT 2.6920 59.1435 2.7180 60.2370 ;
        RECT 2.5840 59.1435 2.6100 60.2370 ;
        RECT 2.4760 59.1435 2.5020 60.2370 ;
        RECT 2.3680 59.1435 2.3940 60.2370 ;
        RECT 2.2600 59.1435 2.2860 60.2370 ;
        RECT 2.1520 59.1435 2.1780 60.2370 ;
        RECT 2.0440 59.1435 2.0700 60.2370 ;
        RECT 1.9360 59.1435 1.9620 60.2370 ;
        RECT 1.8280 59.1435 1.8540 60.2370 ;
        RECT 1.7200 59.1435 1.7460 60.2370 ;
        RECT 1.6120 59.1435 1.6380 60.2370 ;
        RECT 1.5040 59.1435 1.5300 60.2370 ;
        RECT 1.3960 59.1435 1.4220 60.2370 ;
        RECT 1.2880 59.1435 1.3140 60.2370 ;
        RECT 1.1800 59.1435 1.2060 60.2370 ;
        RECT 1.0720 59.1435 1.0980 60.2370 ;
        RECT 0.9640 59.1435 0.9900 60.2370 ;
        RECT 0.8560 59.1435 0.8820 60.2370 ;
        RECT 0.7480 59.1435 0.7740 60.2370 ;
        RECT 0.6400 59.1435 0.6660 60.2370 ;
        RECT 0.5320 59.1435 0.5580 60.2370 ;
        RECT 0.4240 59.1435 0.4500 60.2370 ;
        RECT 0.3160 59.1435 0.3420 60.2370 ;
        RECT 0.2080 59.1435 0.2340 60.2370 ;
        RECT 0.0050 59.1435 0.0900 60.2370 ;
        RECT 15.5530 60.2235 15.6810 61.3170 ;
        RECT 15.5390 60.8890 15.6810 61.2115 ;
        RECT 15.3190 60.6160 15.4530 61.3170 ;
        RECT 15.2960 60.9510 15.4530 61.2090 ;
        RECT 15.3190 60.2235 15.4170 61.3170 ;
        RECT 15.3190 60.3445 15.4310 60.5840 ;
        RECT 15.3190 60.2235 15.4530 60.3125 ;
        RECT 15.0940 60.6740 15.2280 61.3170 ;
        RECT 15.0940 60.2235 15.1920 61.3170 ;
        RECT 14.6770 60.2235 14.7600 61.3170 ;
        RECT 14.6770 60.3120 14.7740 61.2475 ;
        RECT 30.2680 60.2235 30.3530 61.3170 ;
        RECT 30.1240 60.2235 30.1500 61.3170 ;
        RECT 30.0160 60.2235 30.0420 61.3170 ;
        RECT 29.9080 60.2235 29.9340 61.3170 ;
        RECT 29.8000 60.2235 29.8260 61.3170 ;
        RECT 29.6920 60.2235 29.7180 61.3170 ;
        RECT 29.5840 60.2235 29.6100 61.3170 ;
        RECT 29.4760 60.2235 29.5020 61.3170 ;
        RECT 29.3680 60.2235 29.3940 61.3170 ;
        RECT 29.2600 60.2235 29.2860 61.3170 ;
        RECT 29.1520 60.2235 29.1780 61.3170 ;
        RECT 29.0440 60.2235 29.0700 61.3170 ;
        RECT 28.9360 60.2235 28.9620 61.3170 ;
        RECT 28.8280 60.2235 28.8540 61.3170 ;
        RECT 28.7200 60.2235 28.7460 61.3170 ;
        RECT 28.6120 60.2235 28.6380 61.3170 ;
        RECT 28.5040 60.2235 28.5300 61.3170 ;
        RECT 28.3960 60.2235 28.4220 61.3170 ;
        RECT 28.2880 60.2235 28.3140 61.3170 ;
        RECT 28.1800 60.2235 28.2060 61.3170 ;
        RECT 28.0720 60.2235 28.0980 61.3170 ;
        RECT 27.9640 60.2235 27.9900 61.3170 ;
        RECT 27.8560 60.2235 27.8820 61.3170 ;
        RECT 27.7480 60.2235 27.7740 61.3170 ;
        RECT 27.6400 60.2235 27.6660 61.3170 ;
        RECT 27.5320 60.2235 27.5580 61.3170 ;
        RECT 27.4240 60.2235 27.4500 61.3170 ;
        RECT 27.3160 60.2235 27.3420 61.3170 ;
        RECT 27.2080 60.2235 27.2340 61.3170 ;
        RECT 27.1000 60.2235 27.1260 61.3170 ;
        RECT 26.9920 60.2235 27.0180 61.3170 ;
        RECT 26.8840 60.2235 26.9100 61.3170 ;
        RECT 26.7760 60.2235 26.8020 61.3170 ;
        RECT 26.6680 60.2235 26.6940 61.3170 ;
        RECT 26.5600 60.2235 26.5860 61.3170 ;
        RECT 26.4520 60.2235 26.4780 61.3170 ;
        RECT 26.3440 60.2235 26.3700 61.3170 ;
        RECT 26.2360 60.2235 26.2620 61.3170 ;
        RECT 26.1280 60.2235 26.1540 61.3170 ;
        RECT 26.0200 60.2235 26.0460 61.3170 ;
        RECT 25.9120 60.2235 25.9380 61.3170 ;
        RECT 25.8040 60.2235 25.8300 61.3170 ;
        RECT 25.6960 60.2235 25.7220 61.3170 ;
        RECT 25.5880 60.2235 25.6140 61.3170 ;
        RECT 25.4800 60.2235 25.5060 61.3170 ;
        RECT 25.3720 60.2235 25.3980 61.3170 ;
        RECT 25.2640 60.2235 25.2900 61.3170 ;
        RECT 25.1560 60.2235 25.1820 61.3170 ;
        RECT 25.0480 60.2235 25.0740 61.3170 ;
        RECT 24.9400 60.2235 24.9660 61.3170 ;
        RECT 24.8320 60.2235 24.8580 61.3170 ;
        RECT 24.7240 60.2235 24.7500 61.3170 ;
        RECT 24.6160 60.2235 24.6420 61.3170 ;
        RECT 24.5080 60.2235 24.5340 61.3170 ;
        RECT 24.4000 60.2235 24.4260 61.3170 ;
        RECT 24.2920 60.2235 24.3180 61.3170 ;
        RECT 24.1840 60.2235 24.2100 61.3170 ;
        RECT 24.0760 60.2235 24.1020 61.3170 ;
        RECT 23.9680 60.2235 23.9940 61.3170 ;
        RECT 23.8600 60.2235 23.8860 61.3170 ;
        RECT 23.7520 60.2235 23.7780 61.3170 ;
        RECT 23.6440 60.2235 23.6700 61.3170 ;
        RECT 23.5360 60.2235 23.5620 61.3170 ;
        RECT 23.4280 60.2235 23.4540 61.3170 ;
        RECT 23.3200 60.2235 23.3460 61.3170 ;
        RECT 23.2120 60.2235 23.2380 61.3170 ;
        RECT 23.1040 60.2235 23.1300 61.3170 ;
        RECT 22.9960 60.2235 23.0220 61.3170 ;
        RECT 22.8880 60.2235 22.9140 61.3170 ;
        RECT 22.7800 60.2235 22.8060 61.3170 ;
        RECT 22.6720 60.2235 22.6980 61.3170 ;
        RECT 22.5640 60.2235 22.5900 61.3170 ;
        RECT 22.4560 60.2235 22.4820 61.3170 ;
        RECT 22.3480 60.2235 22.3740 61.3170 ;
        RECT 22.2400 60.2235 22.2660 61.3170 ;
        RECT 22.1320 60.2235 22.1580 61.3170 ;
        RECT 22.0240 60.2235 22.0500 61.3170 ;
        RECT 21.9160 60.2235 21.9420 61.3170 ;
        RECT 21.8080 60.2235 21.8340 61.3170 ;
        RECT 21.7000 60.2235 21.7260 61.3170 ;
        RECT 21.5920 60.2235 21.6180 61.3170 ;
        RECT 21.4840 60.2235 21.5100 61.3170 ;
        RECT 21.3760 60.2235 21.4020 61.3170 ;
        RECT 21.2680 60.2235 21.2940 61.3170 ;
        RECT 21.1600 60.2235 21.1860 61.3170 ;
        RECT 21.0520 60.2235 21.0780 61.3170 ;
        RECT 20.9440 60.2235 20.9700 61.3170 ;
        RECT 20.8360 60.2235 20.8620 61.3170 ;
        RECT 20.7280 60.2235 20.7540 61.3170 ;
        RECT 20.6200 60.2235 20.6460 61.3170 ;
        RECT 20.5120 60.2235 20.5380 61.3170 ;
        RECT 20.4040 60.2235 20.4300 61.3170 ;
        RECT 20.2960 60.2235 20.3220 61.3170 ;
        RECT 20.1880 60.2235 20.2140 61.3170 ;
        RECT 20.0800 60.2235 20.1060 61.3170 ;
        RECT 19.9720 60.2235 19.9980 61.3170 ;
        RECT 19.8640 60.2235 19.8900 61.3170 ;
        RECT 19.7560 60.2235 19.7820 61.3170 ;
        RECT 19.6480 60.2235 19.6740 61.3170 ;
        RECT 19.5400 60.2235 19.5660 61.3170 ;
        RECT 19.4320 60.2235 19.4580 61.3170 ;
        RECT 19.3240 60.2235 19.3500 61.3170 ;
        RECT 19.2160 60.2235 19.2420 61.3170 ;
        RECT 19.1080 60.2235 19.1340 61.3170 ;
        RECT 19.0000 60.2235 19.0260 61.3170 ;
        RECT 18.8920 60.2235 18.9180 61.3170 ;
        RECT 18.7840 60.2235 18.8100 61.3170 ;
        RECT 18.6760 60.2235 18.7020 61.3170 ;
        RECT 18.5680 60.2235 18.5940 61.3170 ;
        RECT 18.4600 60.2235 18.4860 61.3170 ;
        RECT 18.3520 60.2235 18.3780 61.3170 ;
        RECT 18.2440 60.2235 18.2700 61.3170 ;
        RECT 18.1360 60.2235 18.1620 61.3170 ;
        RECT 18.0280 60.2235 18.0540 61.3170 ;
        RECT 17.9200 60.2235 17.9460 61.3170 ;
        RECT 17.8120 60.2235 17.8380 61.3170 ;
        RECT 17.7040 60.2235 17.7300 61.3170 ;
        RECT 17.5960 60.2235 17.6220 61.3170 ;
        RECT 17.4880 60.2235 17.5140 61.3170 ;
        RECT 17.3800 60.2235 17.4060 61.3170 ;
        RECT 17.2720 60.2235 17.2980 61.3170 ;
        RECT 17.1640 60.2235 17.1900 61.3170 ;
        RECT 17.0560 60.2235 17.0820 61.3170 ;
        RECT 16.9480 60.2235 16.9740 61.3170 ;
        RECT 16.8400 60.2235 16.8660 61.3170 ;
        RECT 16.7320 60.2235 16.7580 61.3170 ;
        RECT 16.6240 60.2235 16.6500 61.3170 ;
        RECT 16.5160 60.2235 16.5420 61.3170 ;
        RECT 16.4080 60.2235 16.4340 61.3170 ;
        RECT 16.3000 60.2235 16.3260 61.3170 ;
        RECT 16.0870 60.2235 16.1640 61.3170 ;
        RECT 14.1940 60.2235 14.2710 61.3170 ;
        RECT 14.0320 60.2235 14.0580 61.3170 ;
        RECT 13.9240 60.2235 13.9500 61.3170 ;
        RECT 13.8160 60.2235 13.8420 61.3170 ;
        RECT 13.7080 60.2235 13.7340 61.3170 ;
        RECT 13.6000 60.2235 13.6260 61.3170 ;
        RECT 13.4920 60.2235 13.5180 61.3170 ;
        RECT 13.3840 60.2235 13.4100 61.3170 ;
        RECT 13.2760 60.2235 13.3020 61.3170 ;
        RECT 13.1680 60.2235 13.1940 61.3170 ;
        RECT 13.0600 60.2235 13.0860 61.3170 ;
        RECT 12.9520 60.2235 12.9780 61.3170 ;
        RECT 12.8440 60.2235 12.8700 61.3170 ;
        RECT 12.7360 60.2235 12.7620 61.3170 ;
        RECT 12.6280 60.2235 12.6540 61.3170 ;
        RECT 12.5200 60.2235 12.5460 61.3170 ;
        RECT 12.4120 60.2235 12.4380 61.3170 ;
        RECT 12.3040 60.2235 12.3300 61.3170 ;
        RECT 12.1960 60.2235 12.2220 61.3170 ;
        RECT 12.0880 60.2235 12.1140 61.3170 ;
        RECT 11.9800 60.2235 12.0060 61.3170 ;
        RECT 11.8720 60.2235 11.8980 61.3170 ;
        RECT 11.7640 60.2235 11.7900 61.3170 ;
        RECT 11.6560 60.2235 11.6820 61.3170 ;
        RECT 11.5480 60.2235 11.5740 61.3170 ;
        RECT 11.4400 60.2235 11.4660 61.3170 ;
        RECT 11.3320 60.2235 11.3580 61.3170 ;
        RECT 11.2240 60.2235 11.2500 61.3170 ;
        RECT 11.1160 60.2235 11.1420 61.3170 ;
        RECT 11.0080 60.2235 11.0340 61.3170 ;
        RECT 10.9000 60.2235 10.9260 61.3170 ;
        RECT 10.7920 60.2235 10.8180 61.3170 ;
        RECT 10.6840 60.2235 10.7100 61.3170 ;
        RECT 10.5760 60.2235 10.6020 61.3170 ;
        RECT 10.4680 60.2235 10.4940 61.3170 ;
        RECT 10.3600 60.2235 10.3860 61.3170 ;
        RECT 10.2520 60.2235 10.2780 61.3170 ;
        RECT 10.1440 60.2235 10.1700 61.3170 ;
        RECT 10.0360 60.2235 10.0620 61.3170 ;
        RECT 9.9280 60.2235 9.9540 61.3170 ;
        RECT 9.8200 60.2235 9.8460 61.3170 ;
        RECT 9.7120 60.2235 9.7380 61.3170 ;
        RECT 9.6040 60.2235 9.6300 61.3170 ;
        RECT 9.4960 60.2235 9.5220 61.3170 ;
        RECT 9.3880 60.2235 9.4140 61.3170 ;
        RECT 9.2800 60.2235 9.3060 61.3170 ;
        RECT 9.1720 60.2235 9.1980 61.3170 ;
        RECT 9.0640 60.2235 9.0900 61.3170 ;
        RECT 8.9560 60.2235 8.9820 61.3170 ;
        RECT 8.8480 60.2235 8.8740 61.3170 ;
        RECT 8.7400 60.2235 8.7660 61.3170 ;
        RECT 8.6320 60.2235 8.6580 61.3170 ;
        RECT 8.5240 60.2235 8.5500 61.3170 ;
        RECT 8.4160 60.2235 8.4420 61.3170 ;
        RECT 8.3080 60.2235 8.3340 61.3170 ;
        RECT 8.2000 60.2235 8.2260 61.3170 ;
        RECT 8.0920 60.2235 8.1180 61.3170 ;
        RECT 7.9840 60.2235 8.0100 61.3170 ;
        RECT 7.8760 60.2235 7.9020 61.3170 ;
        RECT 7.7680 60.2235 7.7940 61.3170 ;
        RECT 7.6600 60.2235 7.6860 61.3170 ;
        RECT 7.5520 60.2235 7.5780 61.3170 ;
        RECT 7.4440 60.2235 7.4700 61.3170 ;
        RECT 7.3360 60.2235 7.3620 61.3170 ;
        RECT 7.2280 60.2235 7.2540 61.3170 ;
        RECT 7.1200 60.2235 7.1460 61.3170 ;
        RECT 7.0120 60.2235 7.0380 61.3170 ;
        RECT 6.9040 60.2235 6.9300 61.3170 ;
        RECT 6.7960 60.2235 6.8220 61.3170 ;
        RECT 6.6880 60.2235 6.7140 61.3170 ;
        RECT 6.5800 60.2235 6.6060 61.3170 ;
        RECT 6.4720 60.2235 6.4980 61.3170 ;
        RECT 6.3640 60.2235 6.3900 61.3170 ;
        RECT 6.2560 60.2235 6.2820 61.3170 ;
        RECT 6.1480 60.2235 6.1740 61.3170 ;
        RECT 6.0400 60.2235 6.0660 61.3170 ;
        RECT 5.9320 60.2235 5.9580 61.3170 ;
        RECT 5.8240 60.2235 5.8500 61.3170 ;
        RECT 5.7160 60.2235 5.7420 61.3170 ;
        RECT 5.6080 60.2235 5.6340 61.3170 ;
        RECT 5.5000 60.2235 5.5260 61.3170 ;
        RECT 5.3920 60.2235 5.4180 61.3170 ;
        RECT 5.2840 60.2235 5.3100 61.3170 ;
        RECT 5.1760 60.2235 5.2020 61.3170 ;
        RECT 5.0680 60.2235 5.0940 61.3170 ;
        RECT 4.9600 60.2235 4.9860 61.3170 ;
        RECT 4.8520 60.2235 4.8780 61.3170 ;
        RECT 4.7440 60.2235 4.7700 61.3170 ;
        RECT 4.6360 60.2235 4.6620 61.3170 ;
        RECT 4.5280 60.2235 4.5540 61.3170 ;
        RECT 4.4200 60.2235 4.4460 61.3170 ;
        RECT 4.3120 60.2235 4.3380 61.3170 ;
        RECT 4.2040 60.2235 4.2300 61.3170 ;
        RECT 4.0960 60.2235 4.1220 61.3170 ;
        RECT 3.9880 60.2235 4.0140 61.3170 ;
        RECT 3.8800 60.2235 3.9060 61.3170 ;
        RECT 3.7720 60.2235 3.7980 61.3170 ;
        RECT 3.6640 60.2235 3.6900 61.3170 ;
        RECT 3.5560 60.2235 3.5820 61.3170 ;
        RECT 3.4480 60.2235 3.4740 61.3170 ;
        RECT 3.3400 60.2235 3.3660 61.3170 ;
        RECT 3.2320 60.2235 3.2580 61.3170 ;
        RECT 3.1240 60.2235 3.1500 61.3170 ;
        RECT 3.0160 60.2235 3.0420 61.3170 ;
        RECT 2.9080 60.2235 2.9340 61.3170 ;
        RECT 2.8000 60.2235 2.8260 61.3170 ;
        RECT 2.6920 60.2235 2.7180 61.3170 ;
        RECT 2.5840 60.2235 2.6100 61.3170 ;
        RECT 2.4760 60.2235 2.5020 61.3170 ;
        RECT 2.3680 60.2235 2.3940 61.3170 ;
        RECT 2.2600 60.2235 2.2860 61.3170 ;
        RECT 2.1520 60.2235 2.1780 61.3170 ;
        RECT 2.0440 60.2235 2.0700 61.3170 ;
        RECT 1.9360 60.2235 1.9620 61.3170 ;
        RECT 1.8280 60.2235 1.8540 61.3170 ;
        RECT 1.7200 60.2235 1.7460 61.3170 ;
        RECT 1.6120 60.2235 1.6380 61.3170 ;
        RECT 1.5040 60.2235 1.5300 61.3170 ;
        RECT 1.3960 60.2235 1.4220 61.3170 ;
        RECT 1.2880 60.2235 1.3140 61.3170 ;
        RECT 1.1800 60.2235 1.2060 61.3170 ;
        RECT 1.0720 60.2235 1.0980 61.3170 ;
        RECT 0.9640 60.2235 0.9900 61.3170 ;
        RECT 0.8560 60.2235 0.8820 61.3170 ;
        RECT 0.7480 60.2235 0.7740 61.3170 ;
        RECT 0.6400 60.2235 0.6660 61.3170 ;
        RECT 0.5320 60.2235 0.5580 61.3170 ;
        RECT 0.4240 60.2235 0.4500 61.3170 ;
        RECT 0.3160 60.2235 0.3420 61.3170 ;
        RECT 0.2080 60.2235 0.2340 61.3170 ;
        RECT 0.0050 60.2235 0.0900 61.3170 ;
        RECT 15.5530 61.3035 15.6810 62.3970 ;
        RECT 15.5390 61.9690 15.6810 62.2915 ;
        RECT 15.3190 61.6960 15.4530 62.3970 ;
        RECT 15.2960 62.0310 15.4530 62.2890 ;
        RECT 15.3190 61.3035 15.4170 62.3970 ;
        RECT 15.3190 61.4245 15.4310 61.6640 ;
        RECT 15.3190 61.3035 15.4530 61.3925 ;
        RECT 15.0940 61.7540 15.2280 62.3970 ;
        RECT 15.0940 61.3035 15.1920 62.3970 ;
        RECT 14.6770 61.3035 14.7600 62.3970 ;
        RECT 14.6770 61.3920 14.7740 62.3275 ;
        RECT 30.2680 61.3035 30.3530 62.3970 ;
        RECT 30.1240 61.3035 30.1500 62.3970 ;
        RECT 30.0160 61.3035 30.0420 62.3970 ;
        RECT 29.9080 61.3035 29.9340 62.3970 ;
        RECT 29.8000 61.3035 29.8260 62.3970 ;
        RECT 29.6920 61.3035 29.7180 62.3970 ;
        RECT 29.5840 61.3035 29.6100 62.3970 ;
        RECT 29.4760 61.3035 29.5020 62.3970 ;
        RECT 29.3680 61.3035 29.3940 62.3970 ;
        RECT 29.2600 61.3035 29.2860 62.3970 ;
        RECT 29.1520 61.3035 29.1780 62.3970 ;
        RECT 29.0440 61.3035 29.0700 62.3970 ;
        RECT 28.9360 61.3035 28.9620 62.3970 ;
        RECT 28.8280 61.3035 28.8540 62.3970 ;
        RECT 28.7200 61.3035 28.7460 62.3970 ;
        RECT 28.6120 61.3035 28.6380 62.3970 ;
        RECT 28.5040 61.3035 28.5300 62.3970 ;
        RECT 28.3960 61.3035 28.4220 62.3970 ;
        RECT 28.2880 61.3035 28.3140 62.3970 ;
        RECT 28.1800 61.3035 28.2060 62.3970 ;
        RECT 28.0720 61.3035 28.0980 62.3970 ;
        RECT 27.9640 61.3035 27.9900 62.3970 ;
        RECT 27.8560 61.3035 27.8820 62.3970 ;
        RECT 27.7480 61.3035 27.7740 62.3970 ;
        RECT 27.6400 61.3035 27.6660 62.3970 ;
        RECT 27.5320 61.3035 27.5580 62.3970 ;
        RECT 27.4240 61.3035 27.4500 62.3970 ;
        RECT 27.3160 61.3035 27.3420 62.3970 ;
        RECT 27.2080 61.3035 27.2340 62.3970 ;
        RECT 27.1000 61.3035 27.1260 62.3970 ;
        RECT 26.9920 61.3035 27.0180 62.3970 ;
        RECT 26.8840 61.3035 26.9100 62.3970 ;
        RECT 26.7760 61.3035 26.8020 62.3970 ;
        RECT 26.6680 61.3035 26.6940 62.3970 ;
        RECT 26.5600 61.3035 26.5860 62.3970 ;
        RECT 26.4520 61.3035 26.4780 62.3970 ;
        RECT 26.3440 61.3035 26.3700 62.3970 ;
        RECT 26.2360 61.3035 26.2620 62.3970 ;
        RECT 26.1280 61.3035 26.1540 62.3970 ;
        RECT 26.0200 61.3035 26.0460 62.3970 ;
        RECT 25.9120 61.3035 25.9380 62.3970 ;
        RECT 25.8040 61.3035 25.8300 62.3970 ;
        RECT 25.6960 61.3035 25.7220 62.3970 ;
        RECT 25.5880 61.3035 25.6140 62.3970 ;
        RECT 25.4800 61.3035 25.5060 62.3970 ;
        RECT 25.3720 61.3035 25.3980 62.3970 ;
        RECT 25.2640 61.3035 25.2900 62.3970 ;
        RECT 25.1560 61.3035 25.1820 62.3970 ;
        RECT 25.0480 61.3035 25.0740 62.3970 ;
        RECT 24.9400 61.3035 24.9660 62.3970 ;
        RECT 24.8320 61.3035 24.8580 62.3970 ;
        RECT 24.7240 61.3035 24.7500 62.3970 ;
        RECT 24.6160 61.3035 24.6420 62.3970 ;
        RECT 24.5080 61.3035 24.5340 62.3970 ;
        RECT 24.4000 61.3035 24.4260 62.3970 ;
        RECT 24.2920 61.3035 24.3180 62.3970 ;
        RECT 24.1840 61.3035 24.2100 62.3970 ;
        RECT 24.0760 61.3035 24.1020 62.3970 ;
        RECT 23.9680 61.3035 23.9940 62.3970 ;
        RECT 23.8600 61.3035 23.8860 62.3970 ;
        RECT 23.7520 61.3035 23.7780 62.3970 ;
        RECT 23.6440 61.3035 23.6700 62.3970 ;
        RECT 23.5360 61.3035 23.5620 62.3970 ;
        RECT 23.4280 61.3035 23.4540 62.3970 ;
        RECT 23.3200 61.3035 23.3460 62.3970 ;
        RECT 23.2120 61.3035 23.2380 62.3970 ;
        RECT 23.1040 61.3035 23.1300 62.3970 ;
        RECT 22.9960 61.3035 23.0220 62.3970 ;
        RECT 22.8880 61.3035 22.9140 62.3970 ;
        RECT 22.7800 61.3035 22.8060 62.3970 ;
        RECT 22.6720 61.3035 22.6980 62.3970 ;
        RECT 22.5640 61.3035 22.5900 62.3970 ;
        RECT 22.4560 61.3035 22.4820 62.3970 ;
        RECT 22.3480 61.3035 22.3740 62.3970 ;
        RECT 22.2400 61.3035 22.2660 62.3970 ;
        RECT 22.1320 61.3035 22.1580 62.3970 ;
        RECT 22.0240 61.3035 22.0500 62.3970 ;
        RECT 21.9160 61.3035 21.9420 62.3970 ;
        RECT 21.8080 61.3035 21.8340 62.3970 ;
        RECT 21.7000 61.3035 21.7260 62.3970 ;
        RECT 21.5920 61.3035 21.6180 62.3970 ;
        RECT 21.4840 61.3035 21.5100 62.3970 ;
        RECT 21.3760 61.3035 21.4020 62.3970 ;
        RECT 21.2680 61.3035 21.2940 62.3970 ;
        RECT 21.1600 61.3035 21.1860 62.3970 ;
        RECT 21.0520 61.3035 21.0780 62.3970 ;
        RECT 20.9440 61.3035 20.9700 62.3970 ;
        RECT 20.8360 61.3035 20.8620 62.3970 ;
        RECT 20.7280 61.3035 20.7540 62.3970 ;
        RECT 20.6200 61.3035 20.6460 62.3970 ;
        RECT 20.5120 61.3035 20.5380 62.3970 ;
        RECT 20.4040 61.3035 20.4300 62.3970 ;
        RECT 20.2960 61.3035 20.3220 62.3970 ;
        RECT 20.1880 61.3035 20.2140 62.3970 ;
        RECT 20.0800 61.3035 20.1060 62.3970 ;
        RECT 19.9720 61.3035 19.9980 62.3970 ;
        RECT 19.8640 61.3035 19.8900 62.3970 ;
        RECT 19.7560 61.3035 19.7820 62.3970 ;
        RECT 19.6480 61.3035 19.6740 62.3970 ;
        RECT 19.5400 61.3035 19.5660 62.3970 ;
        RECT 19.4320 61.3035 19.4580 62.3970 ;
        RECT 19.3240 61.3035 19.3500 62.3970 ;
        RECT 19.2160 61.3035 19.2420 62.3970 ;
        RECT 19.1080 61.3035 19.1340 62.3970 ;
        RECT 19.0000 61.3035 19.0260 62.3970 ;
        RECT 18.8920 61.3035 18.9180 62.3970 ;
        RECT 18.7840 61.3035 18.8100 62.3970 ;
        RECT 18.6760 61.3035 18.7020 62.3970 ;
        RECT 18.5680 61.3035 18.5940 62.3970 ;
        RECT 18.4600 61.3035 18.4860 62.3970 ;
        RECT 18.3520 61.3035 18.3780 62.3970 ;
        RECT 18.2440 61.3035 18.2700 62.3970 ;
        RECT 18.1360 61.3035 18.1620 62.3970 ;
        RECT 18.0280 61.3035 18.0540 62.3970 ;
        RECT 17.9200 61.3035 17.9460 62.3970 ;
        RECT 17.8120 61.3035 17.8380 62.3970 ;
        RECT 17.7040 61.3035 17.7300 62.3970 ;
        RECT 17.5960 61.3035 17.6220 62.3970 ;
        RECT 17.4880 61.3035 17.5140 62.3970 ;
        RECT 17.3800 61.3035 17.4060 62.3970 ;
        RECT 17.2720 61.3035 17.2980 62.3970 ;
        RECT 17.1640 61.3035 17.1900 62.3970 ;
        RECT 17.0560 61.3035 17.0820 62.3970 ;
        RECT 16.9480 61.3035 16.9740 62.3970 ;
        RECT 16.8400 61.3035 16.8660 62.3970 ;
        RECT 16.7320 61.3035 16.7580 62.3970 ;
        RECT 16.6240 61.3035 16.6500 62.3970 ;
        RECT 16.5160 61.3035 16.5420 62.3970 ;
        RECT 16.4080 61.3035 16.4340 62.3970 ;
        RECT 16.3000 61.3035 16.3260 62.3970 ;
        RECT 16.0870 61.3035 16.1640 62.3970 ;
        RECT 14.1940 61.3035 14.2710 62.3970 ;
        RECT 14.0320 61.3035 14.0580 62.3970 ;
        RECT 13.9240 61.3035 13.9500 62.3970 ;
        RECT 13.8160 61.3035 13.8420 62.3970 ;
        RECT 13.7080 61.3035 13.7340 62.3970 ;
        RECT 13.6000 61.3035 13.6260 62.3970 ;
        RECT 13.4920 61.3035 13.5180 62.3970 ;
        RECT 13.3840 61.3035 13.4100 62.3970 ;
        RECT 13.2760 61.3035 13.3020 62.3970 ;
        RECT 13.1680 61.3035 13.1940 62.3970 ;
        RECT 13.0600 61.3035 13.0860 62.3970 ;
        RECT 12.9520 61.3035 12.9780 62.3970 ;
        RECT 12.8440 61.3035 12.8700 62.3970 ;
        RECT 12.7360 61.3035 12.7620 62.3970 ;
        RECT 12.6280 61.3035 12.6540 62.3970 ;
        RECT 12.5200 61.3035 12.5460 62.3970 ;
        RECT 12.4120 61.3035 12.4380 62.3970 ;
        RECT 12.3040 61.3035 12.3300 62.3970 ;
        RECT 12.1960 61.3035 12.2220 62.3970 ;
        RECT 12.0880 61.3035 12.1140 62.3970 ;
        RECT 11.9800 61.3035 12.0060 62.3970 ;
        RECT 11.8720 61.3035 11.8980 62.3970 ;
        RECT 11.7640 61.3035 11.7900 62.3970 ;
        RECT 11.6560 61.3035 11.6820 62.3970 ;
        RECT 11.5480 61.3035 11.5740 62.3970 ;
        RECT 11.4400 61.3035 11.4660 62.3970 ;
        RECT 11.3320 61.3035 11.3580 62.3970 ;
        RECT 11.2240 61.3035 11.2500 62.3970 ;
        RECT 11.1160 61.3035 11.1420 62.3970 ;
        RECT 11.0080 61.3035 11.0340 62.3970 ;
        RECT 10.9000 61.3035 10.9260 62.3970 ;
        RECT 10.7920 61.3035 10.8180 62.3970 ;
        RECT 10.6840 61.3035 10.7100 62.3970 ;
        RECT 10.5760 61.3035 10.6020 62.3970 ;
        RECT 10.4680 61.3035 10.4940 62.3970 ;
        RECT 10.3600 61.3035 10.3860 62.3970 ;
        RECT 10.2520 61.3035 10.2780 62.3970 ;
        RECT 10.1440 61.3035 10.1700 62.3970 ;
        RECT 10.0360 61.3035 10.0620 62.3970 ;
        RECT 9.9280 61.3035 9.9540 62.3970 ;
        RECT 9.8200 61.3035 9.8460 62.3970 ;
        RECT 9.7120 61.3035 9.7380 62.3970 ;
        RECT 9.6040 61.3035 9.6300 62.3970 ;
        RECT 9.4960 61.3035 9.5220 62.3970 ;
        RECT 9.3880 61.3035 9.4140 62.3970 ;
        RECT 9.2800 61.3035 9.3060 62.3970 ;
        RECT 9.1720 61.3035 9.1980 62.3970 ;
        RECT 9.0640 61.3035 9.0900 62.3970 ;
        RECT 8.9560 61.3035 8.9820 62.3970 ;
        RECT 8.8480 61.3035 8.8740 62.3970 ;
        RECT 8.7400 61.3035 8.7660 62.3970 ;
        RECT 8.6320 61.3035 8.6580 62.3970 ;
        RECT 8.5240 61.3035 8.5500 62.3970 ;
        RECT 8.4160 61.3035 8.4420 62.3970 ;
        RECT 8.3080 61.3035 8.3340 62.3970 ;
        RECT 8.2000 61.3035 8.2260 62.3970 ;
        RECT 8.0920 61.3035 8.1180 62.3970 ;
        RECT 7.9840 61.3035 8.0100 62.3970 ;
        RECT 7.8760 61.3035 7.9020 62.3970 ;
        RECT 7.7680 61.3035 7.7940 62.3970 ;
        RECT 7.6600 61.3035 7.6860 62.3970 ;
        RECT 7.5520 61.3035 7.5780 62.3970 ;
        RECT 7.4440 61.3035 7.4700 62.3970 ;
        RECT 7.3360 61.3035 7.3620 62.3970 ;
        RECT 7.2280 61.3035 7.2540 62.3970 ;
        RECT 7.1200 61.3035 7.1460 62.3970 ;
        RECT 7.0120 61.3035 7.0380 62.3970 ;
        RECT 6.9040 61.3035 6.9300 62.3970 ;
        RECT 6.7960 61.3035 6.8220 62.3970 ;
        RECT 6.6880 61.3035 6.7140 62.3970 ;
        RECT 6.5800 61.3035 6.6060 62.3970 ;
        RECT 6.4720 61.3035 6.4980 62.3970 ;
        RECT 6.3640 61.3035 6.3900 62.3970 ;
        RECT 6.2560 61.3035 6.2820 62.3970 ;
        RECT 6.1480 61.3035 6.1740 62.3970 ;
        RECT 6.0400 61.3035 6.0660 62.3970 ;
        RECT 5.9320 61.3035 5.9580 62.3970 ;
        RECT 5.8240 61.3035 5.8500 62.3970 ;
        RECT 5.7160 61.3035 5.7420 62.3970 ;
        RECT 5.6080 61.3035 5.6340 62.3970 ;
        RECT 5.5000 61.3035 5.5260 62.3970 ;
        RECT 5.3920 61.3035 5.4180 62.3970 ;
        RECT 5.2840 61.3035 5.3100 62.3970 ;
        RECT 5.1760 61.3035 5.2020 62.3970 ;
        RECT 5.0680 61.3035 5.0940 62.3970 ;
        RECT 4.9600 61.3035 4.9860 62.3970 ;
        RECT 4.8520 61.3035 4.8780 62.3970 ;
        RECT 4.7440 61.3035 4.7700 62.3970 ;
        RECT 4.6360 61.3035 4.6620 62.3970 ;
        RECT 4.5280 61.3035 4.5540 62.3970 ;
        RECT 4.4200 61.3035 4.4460 62.3970 ;
        RECT 4.3120 61.3035 4.3380 62.3970 ;
        RECT 4.2040 61.3035 4.2300 62.3970 ;
        RECT 4.0960 61.3035 4.1220 62.3970 ;
        RECT 3.9880 61.3035 4.0140 62.3970 ;
        RECT 3.8800 61.3035 3.9060 62.3970 ;
        RECT 3.7720 61.3035 3.7980 62.3970 ;
        RECT 3.6640 61.3035 3.6900 62.3970 ;
        RECT 3.5560 61.3035 3.5820 62.3970 ;
        RECT 3.4480 61.3035 3.4740 62.3970 ;
        RECT 3.3400 61.3035 3.3660 62.3970 ;
        RECT 3.2320 61.3035 3.2580 62.3970 ;
        RECT 3.1240 61.3035 3.1500 62.3970 ;
        RECT 3.0160 61.3035 3.0420 62.3970 ;
        RECT 2.9080 61.3035 2.9340 62.3970 ;
        RECT 2.8000 61.3035 2.8260 62.3970 ;
        RECT 2.6920 61.3035 2.7180 62.3970 ;
        RECT 2.5840 61.3035 2.6100 62.3970 ;
        RECT 2.4760 61.3035 2.5020 62.3970 ;
        RECT 2.3680 61.3035 2.3940 62.3970 ;
        RECT 2.2600 61.3035 2.2860 62.3970 ;
        RECT 2.1520 61.3035 2.1780 62.3970 ;
        RECT 2.0440 61.3035 2.0700 62.3970 ;
        RECT 1.9360 61.3035 1.9620 62.3970 ;
        RECT 1.8280 61.3035 1.8540 62.3970 ;
        RECT 1.7200 61.3035 1.7460 62.3970 ;
        RECT 1.6120 61.3035 1.6380 62.3970 ;
        RECT 1.5040 61.3035 1.5300 62.3970 ;
        RECT 1.3960 61.3035 1.4220 62.3970 ;
        RECT 1.2880 61.3035 1.3140 62.3970 ;
        RECT 1.1800 61.3035 1.2060 62.3970 ;
        RECT 1.0720 61.3035 1.0980 62.3970 ;
        RECT 0.9640 61.3035 0.9900 62.3970 ;
        RECT 0.8560 61.3035 0.8820 62.3970 ;
        RECT 0.7480 61.3035 0.7740 62.3970 ;
        RECT 0.6400 61.3035 0.6660 62.3970 ;
        RECT 0.5320 61.3035 0.5580 62.3970 ;
        RECT 0.4240 61.3035 0.4500 62.3970 ;
        RECT 0.3160 61.3035 0.3420 62.3970 ;
        RECT 0.2080 61.3035 0.2340 62.3970 ;
        RECT 0.0050 61.3035 0.0900 62.3970 ;
        RECT 15.5530 62.3835 15.6810 63.4770 ;
        RECT 15.5390 63.0490 15.6810 63.3715 ;
        RECT 15.3190 62.7760 15.4530 63.4770 ;
        RECT 15.2960 63.1110 15.4530 63.3690 ;
        RECT 15.3190 62.3835 15.4170 63.4770 ;
        RECT 15.3190 62.5045 15.4310 62.7440 ;
        RECT 15.3190 62.3835 15.4530 62.4725 ;
        RECT 15.0940 62.8340 15.2280 63.4770 ;
        RECT 15.0940 62.3835 15.1920 63.4770 ;
        RECT 14.6770 62.3835 14.7600 63.4770 ;
        RECT 14.6770 62.4720 14.7740 63.4075 ;
        RECT 30.2680 62.3835 30.3530 63.4770 ;
        RECT 30.1240 62.3835 30.1500 63.4770 ;
        RECT 30.0160 62.3835 30.0420 63.4770 ;
        RECT 29.9080 62.3835 29.9340 63.4770 ;
        RECT 29.8000 62.3835 29.8260 63.4770 ;
        RECT 29.6920 62.3835 29.7180 63.4770 ;
        RECT 29.5840 62.3835 29.6100 63.4770 ;
        RECT 29.4760 62.3835 29.5020 63.4770 ;
        RECT 29.3680 62.3835 29.3940 63.4770 ;
        RECT 29.2600 62.3835 29.2860 63.4770 ;
        RECT 29.1520 62.3835 29.1780 63.4770 ;
        RECT 29.0440 62.3835 29.0700 63.4770 ;
        RECT 28.9360 62.3835 28.9620 63.4770 ;
        RECT 28.8280 62.3835 28.8540 63.4770 ;
        RECT 28.7200 62.3835 28.7460 63.4770 ;
        RECT 28.6120 62.3835 28.6380 63.4770 ;
        RECT 28.5040 62.3835 28.5300 63.4770 ;
        RECT 28.3960 62.3835 28.4220 63.4770 ;
        RECT 28.2880 62.3835 28.3140 63.4770 ;
        RECT 28.1800 62.3835 28.2060 63.4770 ;
        RECT 28.0720 62.3835 28.0980 63.4770 ;
        RECT 27.9640 62.3835 27.9900 63.4770 ;
        RECT 27.8560 62.3835 27.8820 63.4770 ;
        RECT 27.7480 62.3835 27.7740 63.4770 ;
        RECT 27.6400 62.3835 27.6660 63.4770 ;
        RECT 27.5320 62.3835 27.5580 63.4770 ;
        RECT 27.4240 62.3835 27.4500 63.4770 ;
        RECT 27.3160 62.3835 27.3420 63.4770 ;
        RECT 27.2080 62.3835 27.2340 63.4770 ;
        RECT 27.1000 62.3835 27.1260 63.4770 ;
        RECT 26.9920 62.3835 27.0180 63.4770 ;
        RECT 26.8840 62.3835 26.9100 63.4770 ;
        RECT 26.7760 62.3835 26.8020 63.4770 ;
        RECT 26.6680 62.3835 26.6940 63.4770 ;
        RECT 26.5600 62.3835 26.5860 63.4770 ;
        RECT 26.4520 62.3835 26.4780 63.4770 ;
        RECT 26.3440 62.3835 26.3700 63.4770 ;
        RECT 26.2360 62.3835 26.2620 63.4770 ;
        RECT 26.1280 62.3835 26.1540 63.4770 ;
        RECT 26.0200 62.3835 26.0460 63.4770 ;
        RECT 25.9120 62.3835 25.9380 63.4770 ;
        RECT 25.8040 62.3835 25.8300 63.4770 ;
        RECT 25.6960 62.3835 25.7220 63.4770 ;
        RECT 25.5880 62.3835 25.6140 63.4770 ;
        RECT 25.4800 62.3835 25.5060 63.4770 ;
        RECT 25.3720 62.3835 25.3980 63.4770 ;
        RECT 25.2640 62.3835 25.2900 63.4770 ;
        RECT 25.1560 62.3835 25.1820 63.4770 ;
        RECT 25.0480 62.3835 25.0740 63.4770 ;
        RECT 24.9400 62.3835 24.9660 63.4770 ;
        RECT 24.8320 62.3835 24.8580 63.4770 ;
        RECT 24.7240 62.3835 24.7500 63.4770 ;
        RECT 24.6160 62.3835 24.6420 63.4770 ;
        RECT 24.5080 62.3835 24.5340 63.4770 ;
        RECT 24.4000 62.3835 24.4260 63.4770 ;
        RECT 24.2920 62.3835 24.3180 63.4770 ;
        RECT 24.1840 62.3835 24.2100 63.4770 ;
        RECT 24.0760 62.3835 24.1020 63.4770 ;
        RECT 23.9680 62.3835 23.9940 63.4770 ;
        RECT 23.8600 62.3835 23.8860 63.4770 ;
        RECT 23.7520 62.3835 23.7780 63.4770 ;
        RECT 23.6440 62.3835 23.6700 63.4770 ;
        RECT 23.5360 62.3835 23.5620 63.4770 ;
        RECT 23.4280 62.3835 23.4540 63.4770 ;
        RECT 23.3200 62.3835 23.3460 63.4770 ;
        RECT 23.2120 62.3835 23.2380 63.4770 ;
        RECT 23.1040 62.3835 23.1300 63.4770 ;
        RECT 22.9960 62.3835 23.0220 63.4770 ;
        RECT 22.8880 62.3835 22.9140 63.4770 ;
        RECT 22.7800 62.3835 22.8060 63.4770 ;
        RECT 22.6720 62.3835 22.6980 63.4770 ;
        RECT 22.5640 62.3835 22.5900 63.4770 ;
        RECT 22.4560 62.3835 22.4820 63.4770 ;
        RECT 22.3480 62.3835 22.3740 63.4770 ;
        RECT 22.2400 62.3835 22.2660 63.4770 ;
        RECT 22.1320 62.3835 22.1580 63.4770 ;
        RECT 22.0240 62.3835 22.0500 63.4770 ;
        RECT 21.9160 62.3835 21.9420 63.4770 ;
        RECT 21.8080 62.3835 21.8340 63.4770 ;
        RECT 21.7000 62.3835 21.7260 63.4770 ;
        RECT 21.5920 62.3835 21.6180 63.4770 ;
        RECT 21.4840 62.3835 21.5100 63.4770 ;
        RECT 21.3760 62.3835 21.4020 63.4770 ;
        RECT 21.2680 62.3835 21.2940 63.4770 ;
        RECT 21.1600 62.3835 21.1860 63.4770 ;
        RECT 21.0520 62.3835 21.0780 63.4770 ;
        RECT 20.9440 62.3835 20.9700 63.4770 ;
        RECT 20.8360 62.3835 20.8620 63.4770 ;
        RECT 20.7280 62.3835 20.7540 63.4770 ;
        RECT 20.6200 62.3835 20.6460 63.4770 ;
        RECT 20.5120 62.3835 20.5380 63.4770 ;
        RECT 20.4040 62.3835 20.4300 63.4770 ;
        RECT 20.2960 62.3835 20.3220 63.4770 ;
        RECT 20.1880 62.3835 20.2140 63.4770 ;
        RECT 20.0800 62.3835 20.1060 63.4770 ;
        RECT 19.9720 62.3835 19.9980 63.4770 ;
        RECT 19.8640 62.3835 19.8900 63.4770 ;
        RECT 19.7560 62.3835 19.7820 63.4770 ;
        RECT 19.6480 62.3835 19.6740 63.4770 ;
        RECT 19.5400 62.3835 19.5660 63.4770 ;
        RECT 19.4320 62.3835 19.4580 63.4770 ;
        RECT 19.3240 62.3835 19.3500 63.4770 ;
        RECT 19.2160 62.3835 19.2420 63.4770 ;
        RECT 19.1080 62.3835 19.1340 63.4770 ;
        RECT 19.0000 62.3835 19.0260 63.4770 ;
        RECT 18.8920 62.3835 18.9180 63.4770 ;
        RECT 18.7840 62.3835 18.8100 63.4770 ;
        RECT 18.6760 62.3835 18.7020 63.4770 ;
        RECT 18.5680 62.3835 18.5940 63.4770 ;
        RECT 18.4600 62.3835 18.4860 63.4770 ;
        RECT 18.3520 62.3835 18.3780 63.4770 ;
        RECT 18.2440 62.3835 18.2700 63.4770 ;
        RECT 18.1360 62.3835 18.1620 63.4770 ;
        RECT 18.0280 62.3835 18.0540 63.4770 ;
        RECT 17.9200 62.3835 17.9460 63.4770 ;
        RECT 17.8120 62.3835 17.8380 63.4770 ;
        RECT 17.7040 62.3835 17.7300 63.4770 ;
        RECT 17.5960 62.3835 17.6220 63.4770 ;
        RECT 17.4880 62.3835 17.5140 63.4770 ;
        RECT 17.3800 62.3835 17.4060 63.4770 ;
        RECT 17.2720 62.3835 17.2980 63.4770 ;
        RECT 17.1640 62.3835 17.1900 63.4770 ;
        RECT 17.0560 62.3835 17.0820 63.4770 ;
        RECT 16.9480 62.3835 16.9740 63.4770 ;
        RECT 16.8400 62.3835 16.8660 63.4770 ;
        RECT 16.7320 62.3835 16.7580 63.4770 ;
        RECT 16.6240 62.3835 16.6500 63.4770 ;
        RECT 16.5160 62.3835 16.5420 63.4770 ;
        RECT 16.4080 62.3835 16.4340 63.4770 ;
        RECT 16.3000 62.3835 16.3260 63.4770 ;
        RECT 16.0870 62.3835 16.1640 63.4770 ;
        RECT 14.1940 62.3835 14.2710 63.4770 ;
        RECT 14.0320 62.3835 14.0580 63.4770 ;
        RECT 13.9240 62.3835 13.9500 63.4770 ;
        RECT 13.8160 62.3835 13.8420 63.4770 ;
        RECT 13.7080 62.3835 13.7340 63.4770 ;
        RECT 13.6000 62.3835 13.6260 63.4770 ;
        RECT 13.4920 62.3835 13.5180 63.4770 ;
        RECT 13.3840 62.3835 13.4100 63.4770 ;
        RECT 13.2760 62.3835 13.3020 63.4770 ;
        RECT 13.1680 62.3835 13.1940 63.4770 ;
        RECT 13.0600 62.3835 13.0860 63.4770 ;
        RECT 12.9520 62.3835 12.9780 63.4770 ;
        RECT 12.8440 62.3835 12.8700 63.4770 ;
        RECT 12.7360 62.3835 12.7620 63.4770 ;
        RECT 12.6280 62.3835 12.6540 63.4770 ;
        RECT 12.5200 62.3835 12.5460 63.4770 ;
        RECT 12.4120 62.3835 12.4380 63.4770 ;
        RECT 12.3040 62.3835 12.3300 63.4770 ;
        RECT 12.1960 62.3835 12.2220 63.4770 ;
        RECT 12.0880 62.3835 12.1140 63.4770 ;
        RECT 11.9800 62.3835 12.0060 63.4770 ;
        RECT 11.8720 62.3835 11.8980 63.4770 ;
        RECT 11.7640 62.3835 11.7900 63.4770 ;
        RECT 11.6560 62.3835 11.6820 63.4770 ;
        RECT 11.5480 62.3835 11.5740 63.4770 ;
        RECT 11.4400 62.3835 11.4660 63.4770 ;
        RECT 11.3320 62.3835 11.3580 63.4770 ;
        RECT 11.2240 62.3835 11.2500 63.4770 ;
        RECT 11.1160 62.3835 11.1420 63.4770 ;
        RECT 11.0080 62.3835 11.0340 63.4770 ;
        RECT 10.9000 62.3835 10.9260 63.4770 ;
        RECT 10.7920 62.3835 10.8180 63.4770 ;
        RECT 10.6840 62.3835 10.7100 63.4770 ;
        RECT 10.5760 62.3835 10.6020 63.4770 ;
        RECT 10.4680 62.3835 10.4940 63.4770 ;
        RECT 10.3600 62.3835 10.3860 63.4770 ;
        RECT 10.2520 62.3835 10.2780 63.4770 ;
        RECT 10.1440 62.3835 10.1700 63.4770 ;
        RECT 10.0360 62.3835 10.0620 63.4770 ;
        RECT 9.9280 62.3835 9.9540 63.4770 ;
        RECT 9.8200 62.3835 9.8460 63.4770 ;
        RECT 9.7120 62.3835 9.7380 63.4770 ;
        RECT 9.6040 62.3835 9.6300 63.4770 ;
        RECT 9.4960 62.3835 9.5220 63.4770 ;
        RECT 9.3880 62.3835 9.4140 63.4770 ;
        RECT 9.2800 62.3835 9.3060 63.4770 ;
        RECT 9.1720 62.3835 9.1980 63.4770 ;
        RECT 9.0640 62.3835 9.0900 63.4770 ;
        RECT 8.9560 62.3835 8.9820 63.4770 ;
        RECT 8.8480 62.3835 8.8740 63.4770 ;
        RECT 8.7400 62.3835 8.7660 63.4770 ;
        RECT 8.6320 62.3835 8.6580 63.4770 ;
        RECT 8.5240 62.3835 8.5500 63.4770 ;
        RECT 8.4160 62.3835 8.4420 63.4770 ;
        RECT 8.3080 62.3835 8.3340 63.4770 ;
        RECT 8.2000 62.3835 8.2260 63.4770 ;
        RECT 8.0920 62.3835 8.1180 63.4770 ;
        RECT 7.9840 62.3835 8.0100 63.4770 ;
        RECT 7.8760 62.3835 7.9020 63.4770 ;
        RECT 7.7680 62.3835 7.7940 63.4770 ;
        RECT 7.6600 62.3835 7.6860 63.4770 ;
        RECT 7.5520 62.3835 7.5780 63.4770 ;
        RECT 7.4440 62.3835 7.4700 63.4770 ;
        RECT 7.3360 62.3835 7.3620 63.4770 ;
        RECT 7.2280 62.3835 7.2540 63.4770 ;
        RECT 7.1200 62.3835 7.1460 63.4770 ;
        RECT 7.0120 62.3835 7.0380 63.4770 ;
        RECT 6.9040 62.3835 6.9300 63.4770 ;
        RECT 6.7960 62.3835 6.8220 63.4770 ;
        RECT 6.6880 62.3835 6.7140 63.4770 ;
        RECT 6.5800 62.3835 6.6060 63.4770 ;
        RECT 6.4720 62.3835 6.4980 63.4770 ;
        RECT 6.3640 62.3835 6.3900 63.4770 ;
        RECT 6.2560 62.3835 6.2820 63.4770 ;
        RECT 6.1480 62.3835 6.1740 63.4770 ;
        RECT 6.0400 62.3835 6.0660 63.4770 ;
        RECT 5.9320 62.3835 5.9580 63.4770 ;
        RECT 5.8240 62.3835 5.8500 63.4770 ;
        RECT 5.7160 62.3835 5.7420 63.4770 ;
        RECT 5.6080 62.3835 5.6340 63.4770 ;
        RECT 5.5000 62.3835 5.5260 63.4770 ;
        RECT 5.3920 62.3835 5.4180 63.4770 ;
        RECT 5.2840 62.3835 5.3100 63.4770 ;
        RECT 5.1760 62.3835 5.2020 63.4770 ;
        RECT 5.0680 62.3835 5.0940 63.4770 ;
        RECT 4.9600 62.3835 4.9860 63.4770 ;
        RECT 4.8520 62.3835 4.8780 63.4770 ;
        RECT 4.7440 62.3835 4.7700 63.4770 ;
        RECT 4.6360 62.3835 4.6620 63.4770 ;
        RECT 4.5280 62.3835 4.5540 63.4770 ;
        RECT 4.4200 62.3835 4.4460 63.4770 ;
        RECT 4.3120 62.3835 4.3380 63.4770 ;
        RECT 4.2040 62.3835 4.2300 63.4770 ;
        RECT 4.0960 62.3835 4.1220 63.4770 ;
        RECT 3.9880 62.3835 4.0140 63.4770 ;
        RECT 3.8800 62.3835 3.9060 63.4770 ;
        RECT 3.7720 62.3835 3.7980 63.4770 ;
        RECT 3.6640 62.3835 3.6900 63.4770 ;
        RECT 3.5560 62.3835 3.5820 63.4770 ;
        RECT 3.4480 62.3835 3.4740 63.4770 ;
        RECT 3.3400 62.3835 3.3660 63.4770 ;
        RECT 3.2320 62.3835 3.2580 63.4770 ;
        RECT 3.1240 62.3835 3.1500 63.4770 ;
        RECT 3.0160 62.3835 3.0420 63.4770 ;
        RECT 2.9080 62.3835 2.9340 63.4770 ;
        RECT 2.8000 62.3835 2.8260 63.4770 ;
        RECT 2.6920 62.3835 2.7180 63.4770 ;
        RECT 2.5840 62.3835 2.6100 63.4770 ;
        RECT 2.4760 62.3835 2.5020 63.4770 ;
        RECT 2.3680 62.3835 2.3940 63.4770 ;
        RECT 2.2600 62.3835 2.2860 63.4770 ;
        RECT 2.1520 62.3835 2.1780 63.4770 ;
        RECT 2.0440 62.3835 2.0700 63.4770 ;
        RECT 1.9360 62.3835 1.9620 63.4770 ;
        RECT 1.8280 62.3835 1.8540 63.4770 ;
        RECT 1.7200 62.3835 1.7460 63.4770 ;
        RECT 1.6120 62.3835 1.6380 63.4770 ;
        RECT 1.5040 62.3835 1.5300 63.4770 ;
        RECT 1.3960 62.3835 1.4220 63.4770 ;
        RECT 1.2880 62.3835 1.3140 63.4770 ;
        RECT 1.1800 62.3835 1.2060 63.4770 ;
        RECT 1.0720 62.3835 1.0980 63.4770 ;
        RECT 0.9640 62.3835 0.9900 63.4770 ;
        RECT 0.8560 62.3835 0.8820 63.4770 ;
        RECT 0.7480 62.3835 0.7740 63.4770 ;
        RECT 0.6400 62.3835 0.6660 63.4770 ;
        RECT 0.5320 62.3835 0.5580 63.4770 ;
        RECT 0.4240 62.3835 0.4500 63.4770 ;
        RECT 0.3160 62.3835 0.3420 63.4770 ;
        RECT 0.2080 62.3835 0.2340 63.4770 ;
        RECT 0.0050 62.3835 0.0900 63.4770 ;
        RECT 15.5530 63.4635 15.6810 64.5570 ;
        RECT 15.5390 64.1290 15.6810 64.4515 ;
        RECT 15.3190 63.8560 15.4530 64.5570 ;
        RECT 15.2960 64.1910 15.4530 64.4490 ;
        RECT 15.3190 63.4635 15.4170 64.5570 ;
        RECT 15.3190 63.5845 15.4310 63.8240 ;
        RECT 15.3190 63.4635 15.4530 63.5525 ;
        RECT 15.0940 63.9140 15.2280 64.5570 ;
        RECT 15.0940 63.4635 15.1920 64.5570 ;
        RECT 14.6770 63.4635 14.7600 64.5570 ;
        RECT 14.6770 63.5520 14.7740 64.4875 ;
        RECT 30.2680 63.4635 30.3530 64.5570 ;
        RECT 30.1240 63.4635 30.1500 64.5570 ;
        RECT 30.0160 63.4635 30.0420 64.5570 ;
        RECT 29.9080 63.4635 29.9340 64.5570 ;
        RECT 29.8000 63.4635 29.8260 64.5570 ;
        RECT 29.6920 63.4635 29.7180 64.5570 ;
        RECT 29.5840 63.4635 29.6100 64.5570 ;
        RECT 29.4760 63.4635 29.5020 64.5570 ;
        RECT 29.3680 63.4635 29.3940 64.5570 ;
        RECT 29.2600 63.4635 29.2860 64.5570 ;
        RECT 29.1520 63.4635 29.1780 64.5570 ;
        RECT 29.0440 63.4635 29.0700 64.5570 ;
        RECT 28.9360 63.4635 28.9620 64.5570 ;
        RECT 28.8280 63.4635 28.8540 64.5570 ;
        RECT 28.7200 63.4635 28.7460 64.5570 ;
        RECT 28.6120 63.4635 28.6380 64.5570 ;
        RECT 28.5040 63.4635 28.5300 64.5570 ;
        RECT 28.3960 63.4635 28.4220 64.5570 ;
        RECT 28.2880 63.4635 28.3140 64.5570 ;
        RECT 28.1800 63.4635 28.2060 64.5570 ;
        RECT 28.0720 63.4635 28.0980 64.5570 ;
        RECT 27.9640 63.4635 27.9900 64.5570 ;
        RECT 27.8560 63.4635 27.8820 64.5570 ;
        RECT 27.7480 63.4635 27.7740 64.5570 ;
        RECT 27.6400 63.4635 27.6660 64.5570 ;
        RECT 27.5320 63.4635 27.5580 64.5570 ;
        RECT 27.4240 63.4635 27.4500 64.5570 ;
        RECT 27.3160 63.4635 27.3420 64.5570 ;
        RECT 27.2080 63.4635 27.2340 64.5570 ;
        RECT 27.1000 63.4635 27.1260 64.5570 ;
        RECT 26.9920 63.4635 27.0180 64.5570 ;
        RECT 26.8840 63.4635 26.9100 64.5570 ;
        RECT 26.7760 63.4635 26.8020 64.5570 ;
        RECT 26.6680 63.4635 26.6940 64.5570 ;
        RECT 26.5600 63.4635 26.5860 64.5570 ;
        RECT 26.4520 63.4635 26.4780 64.5570 ;
        RECT 26.3440 63.4635 26.3700 64.5570 ;
        RECT 26.2360 63.4635 26.2620 64.5570 ;
        RECT 26.1280 63.4635 26.1540 64.5570 ;
        RECT 26.0200 63.4635 26.0460 64.5570 ;
        RECT 25.9120 63.4635 25.9380 64.5570 ;
        RECT 25.8040 63.4635 25.8300 64.5570 ;
        RECT 25.6960 63.4635 25.7220 64.5570 ;
        RECT 25.5880 63.4635 25.6140 64.5570 ;
        RECT 25.4800 63.4635 25.5060 64.5570 ;
        RECT 25.3720 63.4635 25.3980 64.5570 ;
        RECT 25.2640 63.4635 25.2900 64.5570 ;
        RECT 25.1560 63.4635 25.1820 64.5570 ;
        RECT 25.0480 63.4635 25.0740 64.5570 ;
        RECT 24.9400 63.4635 24.9660 64.5570 ;
        RECT 24.8320 63.4635 24.8580 64.5570 ;
        RECT 24.7240 63.4635 24.7500 64.5570 ;
        RECT 24.6160 63.4635 24.6420 64.5570 ;
        RECT 24.5080 63.4635 24.5340 64.5570 ;
        RECT 24.4000 63.4635 24.4260 64.5570 ;
        RECT 24.2920 63.4635 24.3180 64.5570 ;
        RECT 24.1840 63.4635 24.2100 64.5570 ;
        RECT 24.0760 63.4635 24.1020 64.5570 ;
        RECT 23.9680 63.4635 23.9940 64.5570 ;
        RECT 23.8600 63.4635 23.8860 64.5570 ;
        RECT 23.7520 63.4635 23.7780 64.5570 ;
        RECT 23.6440 63.4635 23.6700 64.5570 ;
        RECT 23.5360 63.4635 23.5620 64.5570 ;
        RECT 23.4280 63.4635 23.4540 64.5570 ;
        RECT 23.3200 63.4635 23.3460 64.5570 ;
        RECT 23.2120 63.4635 23.2380 64.5570 ;
        RECT 23.1040 63.4635 23.1300 64.5570 ;
        RECT 22.9960 63.4635 23.0220 64.5570 ;
        RECT 22.8880 63.4635 22.9140 64.5570 ;
        RECT 22.7800 63.4635 22.8060 64.5570 ;
        RECT 22.6720 63.4635 22.6980 64.5570 ;
        RECT 22.5640 63.4635 22.5900 64.5570 ;
        RECT 22.4560 63.4635 22.4820 64.5570 ;
        RECT 22.3480 63.4635 22.3740 64.5570 ;
        RECT 22.2400 63.4635 22.2660 64.5570 ;
        RECT 22.1320 63.4635 22.1580 64.5570 ;
        RECT 22.0240 63.4635 22.0500 64.5570 ;
        RECT 21.9160 63.4635 21.9420 64.5570 ;
        RECT 21.8080 63.4635 21.8340 64.5570 ;
        RECT 21.7000 63.4635 21.7260 64.5570 ;
        RECT 21.5920 63.4635 21.6180 64.5570 ;
        RECT 21.4840 63.4635 21.5100 64.5570 ;
        RECT 21.3760 63.4635 21.4020 64.5570 ;
        RECT 21.2680 63.4635 21.2940 64.5570 ;
        RECT 21.1600 63.4635 21.1860 64.5570 ;
        RECT 21.0520 63.4635 21.0780 64.5570 ;
        RECT 20.9440 63.4635 20.9700 64.5570 ;
        RECT 20.8360 63.4635 20.8620 64.5570 ;
        RECT 20.7280 63.4635 20.7540 64.5570 ;
        RECT 20.6200 63.4635 20.6460 64.5570 ;
        RECT 20.5120 63.4635 20.5380 64.5570 ;
        RECT 20.4040 63.4635 20.4300 64.5570 ;
        RECT 20.2960 63.4635 20.3220 64.5570 ;
        RECT 20.1880 63.4635 20.2140 64.5570 ;
        RECT 20.0800 63.4635 20.1060 64.5570 ;
        RECT 19.9720 63.4635 19.9980 64.5570 ;
        RECT 19.8640 63.4635 19.8900 64.5570 ;
        RECT 19.7560 63.4635 19.7820 64.5570 ;
        RECT 19.6480 63.4635 19.6740 64.5570 ;
        RECT 19.5400 63.4635 19.5660 64.5570 ;
        RECT 19.4320 63.4635 19.4580 64.5570 ;
        RECT 19.3240 63.4635 19.3500 64.5570 ;
        RECT 19.2160 63.4635 19.2420 64.5570 ;
        RECT 19.1080 63.4635 19.1340 64.5570 ;
        RECT 19.0000 63.4635 19.0260 64.5570 ;
        RECT 18.8920 63.4635 18.9180 64.5570 ;
        RECT 18.7840 63.4635 18.8100 64.5570 ;
        RECT 18.6760 63.4635 18.7020 64.5570 ;
        RECT 18.5680 63.4635 18.5940 64.5570 ;
        RECT 18.4600 63.4635 18.4860 64.5570 ;
        RECT 18.3520 63.4635 18.3780 64.5570 ;
        RECT 18.2440 63.4635 18.2700 64.5570 ;
        RECT 18.1360 63.4635 18.1620 64.5570 ;
        RECT 18.0280 63.4635 18.0540 64.5570 ;
        RECT 17.9200 63.4635 17.9460 64.5570 ;
        RECT 17.8120 63.4635 17.8380 64.5570 ;
        RECT 17.7040 63.4635 17.7300 64.5570 ;
        RECT 17.5960 63.4635 17.6220 64.5570 ;
        RECT 17.4880 63.4635 17.5140 64.5570 ;
        RECT 17.3800 63.4635 17.4060 64.5570 ;
        RECT 17.2720 63.4635 17.2980 64.5570 ;
        RECT 17.1640 63.4635 17.1900 64.5570 ;
        RECT 17.0560 63.4635 17.0820 64.5570 ;
        RECT 16.9480 63.4635 16.9740 64.5570 ;
        RECT 16.8400 63.4635 16.8660 64.5570 ;
        RECT 16.7320 63.4635 16.7580 64.5570 ;
        RECT 16.6240 63.4635 16.6500 64.5570 ;
        RECT 16.5160 63.4635 16.5420 64.5570 ;
        RECT 16.4080 63.4635 16.4340 64.5570 ;
        RECT 16.3000 63.4635 16.3260 64.5570 ;
        RECT 16.0870 63.4635 16.1640 64.5570 ;
        RECT 14.1940 63.4635 14.2710 64.5570 ;
        RECT 14.0320 63.4635 14.0580 64.5570 ;
        RECT 13.9240 63.4635 13.9500 64.5570 ;
        RECT 13.8160 63.4635 13.8420 64.5570 ;
        RECT 13.7080 63.4635 13.7340 64.5570 ;
        RECT 13.6000 63.4635 13.6260 64.5570 ;
        RECT 13.4920 63.4635 13.5180 64.5570 ;
        RECT 13.3840 63.4635 13.4100 64.5570 ;
        RECT 13.2760 63.4635 13.3020 64.5570 ;
        RECT 13.1680 63.4635 13.1940 64.5570 ;
        RECT 13.0600 63.4635 13.0860 64.5570 ;
        RECT 12.9520 63.4635 12.9780 64.5570 ;
        RECT 12.8440 63.4635 12.8700 64.5570 ;
        RECT 12.7360 63.4635 12.7620 64.5570 ;
        RECT 12.6280 63.4635 12.6540 64.5570 ;
        RECT 12.5200 63.4635 12.5460 64.5570 ;
        RECT 12.4120 63.4635 12.4380 64.5570 ;
        RECT 12.3040 63.4635 12.3300 64.5570 ;
        RECT 12.1960 63.4635 12.2220 64.5570 ;
        RECT 12.0880 63.4635 12.1140 64.5570 ;
        RECT 11.9800 63.4635 12.0060 64.5570 ;
        RECT 11.8720 63.4635 11.8980 64.5570 ;
        RECT 11.7640 63.4635 11.7900 64.5570 ;
        RECT 11.6560 63.4635 11.6820 64.5570 ;
        RECT 11.5480 63.4635 11.5740 64.5570 ;
        RECT 11.4400 63.4635 11.4660 64.5570 ;
        RECT 11.3320 63.4635 11.3580 64.5570 ;
        RECT 11.2240 63.4635 11.2500 64.5570 ;
        RECT 11.1160 63.4635 11.1420 64.5570 ;
        RECT 11.0080 63.4635 11.0340 64.5570 ;
        RECT 10.9000 63.4635 10.9260 64.5570 ;
        RECT 10.7920 63.4635 10.8180 64.5570 ;
        RECT 10.6840 63.4635 10.7100 64.5570 ;
        RECT 10.5760 63.4635 10.6020 64.5570 ;
        RECT 10.4680 63.4635 10.4940 64.5570 ;
        RECT 10.3600 63.4635 10.3860 64.5570 ;
        RECT 10.2520 63.4635 10.2780 64.5570 ;
        RECT 10.1440 63.4635 10.1700 64.5570 ;
        RECT 10.0360 63.4635 10.0620 64.5570 ;
        RECT 9.9280 63.4635 9.9540 64.5570 ;
        RECT 9.8200 63.4635 9.8460 64.5570 ;
        RECT 9.7120 63.4635 9.7380 64.5570 ;
        RECT 9.6040 63.4635 9.6300 64.5570 ;
        RECT 9.4960 63.4635 9.5220 64.5570 ;
        RECT 9.3880 63.4635 9.4140 64.5570 ;
        RECT 9.2800 63.4635 9.3060 64.5570 ;
        RECT 9.1720 63.4635 9.1980 64.5570 ;
        RECT 9.0640 63.4635 9.0900 64.5570 ;
        RECT 8.9560 63.4635 8.9820 64.5570 ;
        RECT 8.8480 63.4635 8.8740 64.5570 ;
        RECT 8.7400 63.4635 8.7660 64.5570 ;
        RECT 8.6320 63.4635 8.6580 64.5570 ;
        RECT 8.5240 63.4635 8.5500 64.5570 ;
        RECT 8.4160 63.4635 8.4420 64.5570 ;
        RECT 8.3080 63.4635 8.3340 64.5570 ;
        RECT 8.2000 63.4635 8.2260 64.5570 ;
        RECT 8.0920 63.4635 8.1180 64.5570 ;
        RECT 7.9840 63.4635 8.0100 64.5570 ;
        RECT 7.8760 63.4635 7.9020 64.5570 ;
        RECT 7.7680 63.4635 7.7940 64.5570 ;
        RECT 7.6600 63.4635 7.6860 64.5570 ;
        RECT 7.5520 63.4635 7.5780 64.5570 ;
        RECT 7.4440 63.4635 7.4700 64.5570 ;
        RECT 7.3360 63.4635 7.3620 64.5570 ;
        RECT 7.2280 63.4635 7.2540 64.5570 ;
        RECT 7.1200 63.4635 7.1460 64.5570 ;
        RECT 7.0120 63.4635 7.0380 64.5570 ;
        RECT 6.9040 63.4635 6.9300 64.5570 ;
        RECT 6.7960 63.4635 6.8220 64.5570 ;
        RECT 6.6880 63.4635 6.7140 64.5570 ;
        RECT 6.5800 63.4635 6.6060 64.5570 ;
        RECT 6.4720 63.4635 6.4980 64.5570 ;
        RECT 6.3640 63.4635 6.3900 64.5570 ;
        RECT 6.2560 63.4635 6.2820 64.5570 ;
        RECT 6.1480 63.4635 6.1740 64.5570 ;
        RECT 6.0400 63.4635 6.0660 64.5570 ;
        RECT 5.9320 63.4635 5.9580 64.5570 ;
        RECT 5.8240 63.4635 5.8500 64.5570 ;
        RECT 5.7160 63.4635 5.7420 64.5570 ;
        RECT 5.6080 63.4635 5.6340 64.5570 ;
        RECT 5.5000 63.4635 5.5260 64.5570 ;
        RECT 5.3920 63.4635 5.4180 64.5570 ;
        RECT 5.2840 63.4635 5.3100 64.5570 ;
        RECT 5.1760 63.4635 5.2020 64.5570 ;
        RECT 5.0680 63.4635 5.0940 64.5570 ;
        RECT 4.9600 63.4635 4.9860 64.5570 ;
        RECT 4.8520 63.4635 4.8780 64.5570 ;
        RECT 4.7440 63.4635 4.7700 64.5570 ;
        RECT 4.6360 63.4635 4.6620 64.5570 ;
        RECT 4.5280 63.4635 4.5540 64.5570 ;
        RECT 4.4200 63.4635 4.4460 64.5570 ;
        RECT 4.3120 63.4635 4.3380 64.5570 ;
        RECT 4.2040 63.4635 4.2300 64.5570 ;
        RECT 4.0960 63.4635 4.1220 64.5570 ;
        RECT 3.9880 63.4635 4.0140 64.5570 ;
        RECT 3.8800 63.4635 3.9060 64.5570 ;
        RECT 3.7720 63.4635 3.7980 64.5570 ;
        RECT 3.6640 63.4635 3.6900 64.5570 ;
        RECT 3.5560 63.4635 3.5820 64.5570 ;
        RECT 3.4480 63.4635 3.4740 64.5570 ;
        RECT 3.3400 63.4635 3.3660 64.5570 ;
        RECT 3.2320 63.4635 3.2580 64.5570 ;
        RECT 3.1240 63.4635 3.1500 64.5570 ;
        RECT 3.0160 63.4635 3.0420 64.5570 ;
        RECT 2.9080 63.4635 2.9340 64.5570 ;
        RECT 2.8000 63.4635 2.8260 64.5570 ;
        RECT 2.6920 63.4635 2.7180 64.5570 ;
        RECT 2.5840 63.4635 2.6100 64.5570 ;
        RECT 2.4760 63.4635 2.5020 64.5570 ;
        RECT 2.3680 63.4635 2.3940 64.5570 ;
        RECT 2.2600 63.4635 2.2860 64.5570 ;
        RECT 2.1520 63.4635 2.1780 64.5570 ;
        RECT 2.0440 63.4635 2.0700 64.5570 ;
        RECT 1.9360 63.4635 1.9620 64.5570 ;
        RECT 1.8280 63.4635 1.8540 64.5570 ;
        RECT 1.7200 63.4635 1.7460 64.5570 ;
        RECT 1.6120 63.4635 1.6380 64.5570 ;
        RECT 1.5040 63.4635 1.5300 64.5570 ;
        RECT 1.3960 63.4635 1.4220 64.5570 ;
        RECT 1.2880 63.4635 1.3140 64.5570 ;
        RECT 1.1800 63.4635 1.2060 64.5570 ;
        RECT 1.0720 63.4635 1.0980 64.5570 ;
        RECT 0.9640 63.4635 0.9900 64.5570 ;
        RECT 0.8560 63.4635 0.8820 64.5570 ;
        RECT 0.7480 63.4635 0.7740 64.5570 ;
        RECT 0.6400 63.4635 0.6660 64.5570 ;
        RECT 0.5320 63.4635 0.5580 64.5570 ;
        RECT 0.4240 63.4635 0.4500 64.5570 ;
        RECT 0.3160 63.4635 0.3420 64.5570 ;
        RECT 0.2080 63.4635 0.2340 64.5570 ;
        RECT 0.0050 63.4635 0.0900 64.5570 ;
        RECT 15.5530 64.5435 15.6810 65.6370 ;
        RECT 15.5390 65.2090 15.6810 65.5315 ;
        RECT 15.3190 64.9360 15.4530 65.6370 ;
        RECT 15.2960 65.2710 15.4530 65.5290 ;
        RECT 15.3190 64.5435 15.4170 65.6370 ;
        RECT 15.3190 64.6645 15.4310 64.9040 ;
        RECT 15.3190 64.5435 15.4530 64.6325 ;
        RECT 15.0940 64.9940 15.2280 65.6370 ;
        RECT 15.0940 64.5435 15.1920 65.6370 ;
        RECT 14.6770 64.5435 14.7600 65.6370 ;
        RECT 14.6770 64.6320 14.7740 65.5675 ;
        RECT 30.2680 64.5435 30.3530 65.6370 ;
        RECT 30.1240 64.5435 30.1500 65.6370 ;
        RECT 30.0160 64.5435 30.0420 65.6370 ;
        RECT 29.9080 64.5435 29.9340 65.6370 ;
        RECT 29.8000 64.5435 29.8260 65.6370 ;
        RECT 29.6920 64.5435 29.7180 65.6370 ;
        RECT 29.5840 64.5435 29.6100 65.6370 ;
        RECT 29.4760 64.5435 29.5020 65.6370 ;
        RECT 29.3680 64.5435 29.3940 65.6370 ;
        RECT 29.2600 64.5435 29.2860 65.6370 ;
        RECT 29.1520 64.5435 29.1780 65.6370 ;
        RECT 29.0440 64.5435 29.0700 65.6370 ;
        RECT 28.9360 64.5435 28.9620 65.6370 ;
        RECT 28.8280 64.5435 28.8540 65.6370 ;
        RECT 28.7200 64.5435 28.7460 65.6370 ;
        RECT 28.6120 64.5435 28.6380 65.6370 ;
        RECT 28.5040 64.5435 28.5300 65.6370 ;
        RECT 28.3960 64.5435 28.4220 65.6370 ;
        RECT 28.2880 64.5435 28.3140 65.6370 ;
        RECT 28.1800 64.5435 28.2060 65.6370 ;
        RECT 28.0720 64.5435 28.0980 65.6370 ;
        RECT 27.9640 64.5435 27.9900 65.6370 ;
        RECT 27.8560 64.5435 27.8820 65.6370 ;
        RECT 27.7480 64.5435 27.7740 65.6370 ;
        RECT 27.6400 64.5435 27.6660 65.6370 ;
        RECT 27.5320 64.5435 27.5580 65.6370 ;
        RECT 27.4240 64.5435 27.4500 65.6370 ;
        RECT 27.3160 64.5435 27.3420 65.6370 ;
        RECT 27.2080 64.5435 27.2340 65.6370 ;
        RECT 27.1000 64.5435 27.1260 65.6370 ;
        RECT 26.9920 64.5435 27.0180 65.6370 ;
        RECT 26.8840 64.5435 26.9100 65.6370 ;
        RECT 26.7760 64.5435 26.8020 65.6370 ;
        RECT 26.6680 64.5435 26.6940 65.6370 ;
        RECT 26.5600 64.5435 26.5860 65.6370 ;
        RECT 26.4520 64.5435 26.4780 65.6370 ;
        RECT 26.3440 64.5435 26.3700 65.6370 ;
        RECT 26.2360 64.5435 26.2620 65.6370 ;
        RECT 26.1280 64.5435 26.1540 65.6370 ;
        RECT 26.0200 64.5435 26.0460 65.6370 ;
        RECT 25.9120 64.5435 25.9380 65.6370 ;
        RECT 25.8040 64.5435 25.8300 65.6370 ;
        RECT 25.6960 64.5435 25.7220 65.6370 ;
        RECT 25.5880 64.5435 25.6140 65.6370 ;
        RECT 25.4800 64.5435 25.5060 65.6370 ;
        RECT 25.3720 64.5435 25.3980 65.6370 ;
        RECT 25.2640 64.5435 25.2900 65.6370 ;
        RECT 25.1560 64.5435 25.1820 65.6370 ;
        RECT 25.0480 64.5435 25.0740 65.6370 ;
        RECT 24.9400 64.5435 24.9660 65.6370 ;
        RECT 24.8320 64.5435 24.8580 65.6370 ;
        RECT 24.7240 64.5435 24.7500 65.6370 ;
        RECT 24.6160 64.5435 24.6420 65.6370 ;
        RECT 24.5080 64.5435 24.5340 65.6370 ;
        RECT 24.4000 64.5435 24.4260 65.6370 ;
        RECT 24.2920 64.5435 24.3180 65.6370 ;
        RECT 24.1840 64.5435 24.2100 65.6370 ;
        RECT 24.0760 64.5435 24.1020 65.6370 ;
        RECT 23.9680 64.5435 23.9940 65.6370 ;
        RECT 23.8600 64.5435 23.8860 65.6370 ;
        RECT 23.7520 64.5435 23.7780 65.6370 ;
        RECT 23.6440 64.5435 23.6700 65.6370 ;
        RECT 23.5360 64.5435 23.5620 65.6370 ;
        RECT 23.4280 64.5435 23.4540 65.6370 ;
        RECT 23.3200 64.5435 23.3460 65.6370 ;
        RECT 23.2120 64.5435 23.2380 65.6370 ;
        RECT 23.1040 64.5435 23.1300 65.6370 ;
        RECT 22.9960 64.5435 23.0220 65.6370 ;
        RECT 22.8880 64.5435 22.9140 65.6370 ;
        RECT 22.7800 64.5435 22.8060 65.6370 ;
        RECT 22.6720 64.5435 22.6980 65.6370 ;
        RECT 22.5640 64.5435 22.5900 65.6370 ;
        RECT 22.4560 64.5435 22.4820 65.6370 ;
        RECT 22.3480 64.5435 22.3740 65.6370 ;
        RECT 22.2400 64.5435 22.2660 65.6370 ;
        RECT 22.1320 64.5435 22.1580 65.6370 ;
        RECT 22.0240 64.5435 22.0500 65.6370 ;
        RECT 21.9160 64.5435 21.9420 65.6370 ;
        RECT 21.8080 64.5435 21.8340 65.6370 ;
        RECT 21.7000 64.5435 21.7260 65.6370 ;
        RECT 21.5920 64.5435 21.6180 65.6370 ;
        RECT 21.4840 64.5435 21.5100 65.6370 ;
        RECT 21.3760 64.5435 21.4020 65.6370 ;
        RECT 21.2680 64.5435 21.2940 65.6370 ;
        RECT 21.1600 64.5435 21.1860 65.6370 ;
        RECT 21.0520 64.5435 21.0780 65.6370 ;
        RECT 20.9440 64.5435 20.9700 65.6370 ;
        RECT 20.8360 64.5435 20.8620 65.6370 ;
        RECT 20.7280 64.5435 20.7540 65.6370 ;
        RECT 20.6200 64.5435 20.6460 65.6370 ;
        RECT 20.5120 64.5435 20.5380 65.6370 ;
        RECT 20.4040 64.5435 20.4300 65.6370 ;
        RECT 20.2960 64.5435 20.3220 65.6370 ;
        RECT 20.1880 64.5435 20.2140 65.6370 ;
        RECT 20.0800 64.5435 20.1060 65.6370 ;
        RECT 19.9720 64.5435 19.9980 65.6370 ;
        RECT 19.8640 64.5435 19.8900 65.6370 ;
        RECT 19.7560 64.5435 19.7820 65.6370 ;
        RECT 19.6480 64.5435 19.6740 65.6370 ;
        RECT 19.5400 64.5435 19.5660 65.6370 ;
        RECT 19.4320 64.5435 19.4580 65.6370 ;
        RECT 19.3240 64.5435 19.3500 65.6370 ;
        RECT 19.2160 64.5435 19.2420 65.6370 ;
        RECT 19.1080 64.5435 19.1340 65.6370 ;
        RECT 19.0000 64.5435 19.0260 65.6370 ;
        RECT 18.8920 64.5435 18.9180 65.6370 ;
        RECT 18.7840 64.5435 18.8100 65.6370 ;
        RECT 18.6760 64.5435 18.7020 65.6370 ;
        RECT 18.5680 64.5435 18.5940 65.6370 ;
        RECT 18.4600 64.5435 18.4860 65.6370 ;
        RECT 18.3520 64.5435 18.3780 65.6370 ;
        RECT 18.2440 64.5435 18.2700 65.6370 ;
        RECT 18.1360 64.5435 18.1620 65.6370 ;
        RECT 18.0280 64.5435 18.0540 65.6370 ;
        RECT 17.9200 64.5435 17.9460 65.6370 ;
        RECT 17.8120 64.5435 17.8380 65.6370 ;
        RECT 17.7040 64.5435 17.7300 65.6370 ;
        RECT 17.5960 64.5435 17.6220 65.6370 ;
        RECT 17.4880 64.5435 17.5140 65.6370 ;
        RECT 17.3800 64.5435 17.4060 65.6370 ;
        RECT 17.2720 64.5435 17.2980 65.6370 ;
        RECT 17.1640 64.5435 17.1900 65.6370 ;
        RECT 17.0560 64.5435 17.0820 65.6370 ;
        RECT 16.9480 64.5435 16.9740 65.6370 ;
        RECT 16.8400 64.5435 16.8660 65.6370 ;
        RECT 16.7320 64.5435 16.7580 65.6370 ;
        RECT 16.6240 64.5435 16.6500 65.6370 ;
        RECT 16.5160 64.5435 16.5420 65.6370 ;
        RECT 16.4080 64.5435 16.4340 65.6370 ;
        RECT 16.3000 64.5435 16.3260 65.6370 ;
        RECT 16.0870 64.5435 16.1640 65.6370 ;
        RECT 14.1940 64.5435 14.2710 65.6370 ;
        RECT 14.0320 64.5435 14.0580 65.6370 ;
        RECT 13.9240 64.5435 13.9500 65.6370 ;
        RECT 13.8160 64.5435 13.8420 65.6370 ;
        RECT 13.7080 64.5435 13.7340 65.6370 ;
        RECT 13.6000 64.5435 13.6260 65.6370 ;
        RECT 13.4920 64.5435 13.5180 65.6370 ;
        RECT 13.3840 64.5435 13.4100 65.6370 ;
        RECT 13.2760 64.5435 13.3020 65.6370 ;
        RECT 13.1680 64.5435 13.1940 65.6370 ;
        RECT 13.0600 64.5435 13.0860 65.6370 ;
        RECT 12.9520 64.5435 12.9780 65.6370 ;
        RECT 12.8440 64.5435 12.8700 65.6370 ;
        RECT 12.7360 64.5435 12.7620 65.6370 ;
        RECT 12.6280 64.5435 12.6540 65.6370 ;
        RECT 12.5200 64.5435 12.5460 65.6370 ;
        RECT 12.4120 64.5435 12.4380 65.6370 ;
        RECT 12.3040 64.5435 12.3300 65.6370 ;
        RECT 12.1960 64.5435 12.2220 65.6370 ;
        RECT 12.0880 64.5435 12.1140 65.6370 ;
        RECT 11.9800 64.5435 12.0060 65.6370 ;
        RECT 11.8720 64.5435 11.8980 65.6370 ;
        RECT 11.7640 64.5435 11.7900 65.6370 ;
        RECT 11.6560 64.5435 11.6820 65.6370 ;
        RECT 11.5480 64.5435 11.5740 65.6370 ;
        RECT 11.4400 64.5435 11.4660 65.6370 ;
        RECT 11.3320 64.5435 11.3580 65.6370 ;
        RECT 11.2240 64.5435 11.2500 65.6370 ;
        RECT 11.1160 64.5435 11.1420 65.6370 ;
        RECT 11.0080 64.5435 11.0340 65.6370 ;
        RECT 10.9000 64.5435 10.9260 65.6370 ;
        RECT 10.7920 64.5435 10.8180 65.6370 ;
        RECT 10.6840 64.5435 10.7100 65.6370 ;
        RECT 10.5760 64.5435 10.6020 65.6370 ;
        RECT 10.4680 64.5435 10.4940 65.6370 ;
        RECT 10.3600 64.5435 10.3860 65.6370 ;
        RECT 10.2520 64.5435 10.2780 65.6370 ;
        RECT 10.1440 64.5435 10.1700 65.6370 ;
        RECT 10.0360 64.5435 10.0620 65.6370 ;
        RECT 9.9280 64.5435 9.9540 65.6370 ;
        RECT 9.8200 64.5435 9.8460 65.6370 ;
        RECT 9.7120 64.5435 9.7380 65.6370 ;
        RECT 9.6040 64.5435 9.6300 65.6370 ;
        RECT 9.4960 64.5435 9.5220 65.6370 ;
        RECT 9.3880 64.5435 9.4140 65.6370 ;
        RECT 9.2800 64.5435 9.3060 65.6370 ;
        RECT 9.1720 64.5435 9.1980 65.6370 ;
        RECT 9.0640 64.5435 9.0900 65.6370 ;
        RECT 8.9560 64.5435 8.9820 65.6370 ;
        RECT 8.8480 64.5435 8.8740 65.6370 ;
        RECT 8.7400 64.5435 8.7660 65.6370 ;
        RECT 8.6320 64.5435 8.6580 65.6370 ;
        RECT 8.5240 64.5435 8.5500 65.6370 ;
        RECT 8.4160 64.5435 8.4420 65.6370 ;
        RECT 8.3080 64.5435 8.3340 65.6370 ;
        RECT 8.2000 64.5435 8.2260 65.6370 ;
        RECT 8.0920 64.5435 8.1180 65.6370 ;
        RECT 7.9840 64.5435 8.0100 65.6370 ;
        RECT 7.8760 64.5435 7.9020 65.6370 ;
        RECT 7.7680 64.5435 7.7940 65.6370 ;
        RECT 7.6600 64.5435 7.6860 65.6370 ;
        RECT 7.5520 64.5435 7.5780 65.6370 ;
        RECT 7.4440 64.5435 7.4700 65.6370 ;
        RECT 7.3360 64.5435 7.3620 65.6370 ;
        RECT 7.2280 64.5435 7.2540 65.6370 ;
        RECT 7.1200 64.5435 7.1460 65.6370 ;
        RECT 7.0120 64.5435 7.0380 65.6370 ;
        RECT 6.9040 64.5435 6.9300 65.6370 ;
        RECT 6.7960 64.5435 6.8220 65.6370 ;
        RECT 6.6880 64.5435 6.7140 65.6370 ;
        RECT 6.5800 64.5435 6.6060 65.6370 ;
        RECT 6.4720 64.5435 6.4980 65.6370 ;
        RECT 6.3640 64.5435 6.3900 65.6370 ;
        RECT 6.2560 64.5435 6.2820 65.6370 ;
        RECT 6.1480 64.5435 6.1740 65.6370 ;
        RECT 6.0400 64.5435 6.0660 65.6370 ;
        RECT 5.9320 64.5435 5.9580 65.6370 ;
        RECT 5.8240 64.5435 5.8500 65.6370 ;
        RECT 5.7160 64.5435 5.7420 65.6370 ;
        RECT 5.6080 64.5435 5.6340 65.6370 ;
        RECT 5.5000 64.5435 5.5260 65.6370 ;
        RECT 5.3920 64.5435 5.4180 65.6370 ;
        RECT 5.2840 64.5435 5.3100 65.6370 ;
        RECT 5.1760 64.5435 5.2020 65.6370 ;
        RECT 5.0680 64.5435 5.0940 65.6370 ;
        RECT 4.9600 64.5435 4.9860 65.6370 ;
        RECT 4.8520 64.5435 4.8780 65.6370 ;
        RECT 4.7440 64.5435 4.7700 65.6370 ;
        RECT 4.6360 64.5435 4.6620 65.6370 ;
        RECT 4.5280 64.5435 4.5540 65.6370 ;
        RECT 4.4200 64.5435 4.4460 65.6370 ;
        RECT 4.3120 64.5435 4.3380 65.6370 ;
        RECT 4.2040 64.5435 4.2300 65.6370 ;
        RECT 4.0960 64.5435 4.1220 65.6370 ;
        RECT 3.9880 64.5435 4.0140 65.6370 ;
        RECT 3.8800 64.5435 3.9060 65.6370 ;
        RECT 3.7720 64.5435 3.7980 65.6370 ;
        RECT 3.6640 64.5435 3.6900 65.6370 ;
        RECT 3.5560 64.5435 3.5820 65.6370 ;
        RECT 3.4480 64.5435 3.4740 65.6370 ;
        RECT 3.3400 64.5435 3.3660 65.6370 ;
        RECT 3.2320 64.5435 3.2580 65.6370 ;
        RECT 3.1240 64.5435 3.1500 65.6370 ;
        RECT 3.0160 64.5435 3.0420 65.6370 ;
        RECT 2.9080 64.5435 2.9340 65.6370 ;
        RECT 2.8000 64.5435 2.8260 65.6370 ;
        RECT 2.6920 64.5435 2.7180 65.6370 ;
        RECT 2.5840 64.5435 2.6100 65.6370 ;
        RECT 2.4760 64.5435 2.5020 65.6370 ;
        RECT 2.3680 64.5435 2.3940 65.6370 ;
        RECT 2.2600 64.5435 2.2860 65.6370 ;
        RECT 2.1520 64.5435 2.1780 65.6370 ;
        RECT 2.0440 64.5435 2.0700 65.6370 ;
        RECT 1.9360 64.5435 1.9620 65.6370 ;
        RECT 1.8280 64.5435 1.8540 65.6370 ;
        RECT 1.7200 64.5435 1.7460 65.6370 ;
        RECT 1.6120 64.5435 1.6380 65.6370 ;
        RECT 1.5040 64.5435 1.5300 65.6370 ;
        RECT 1.3960 64.5435 1.4220 65.6370 ;
        RECT 1.2880 64.5435 1.3140 65.6370 ;
        RECT 1.1800 64.5435 1.2060 65.6370 ;
        RECT 1.0720 64.5435 1.0980 65.6370 ;
        RECT 0.9640 64.5435 0.9900 65.6370 ;
        RECT 0.8560 64.5435 0.8820 65.6370 ;
        RECT 0.7480 64.5435 0.7740 65.6370 ;
        RECT 0.6400 64.5435 0.6660 65.6370 ;
        RECT 0.5320 64.5435 0.5580 65.6370 ;
        RECT 0.4240 64.5435 0.4500 65.6370 ;
        RECT 0.3160 64.5435 0.3420 65.6370 ;
        RECT 0.2080 64.5435 0.2340 65.6370 ;
        RECT 0.0050 64.5435 0.0900 65.6370 ;
        RECT 15.5530 65.6235 15.6810 66.7170 ;
        RECT 15.5390 66.2890 15.6810 66.6115 ;
        RECT 15.3190 66.0160 15.4530 66.7170 ;
        RECT 15.2960 66.3510 15.4530 66.6090 ;
        RECT 15.3190 65.6235 15.4170 66.7170 ;
        RECT 15.3190 65.7445 15.4310 65.9840 ;
        RECT 15.3190 65.6235 15.4530 65.7125 ;
        RECT 15.0940 66.0740 15.2280 66.7170 ;
        RECT 15.0940 65.6235 15.1920 66.7170 ;
        RECT 14.6770 65.6235 14.7600 66.7170 ;
        RECT 14.6770 65.7120 14.7740 66.6475 ;
        RECT 30.2680 65.6235 30.3530 66.7170 ;
        RECT 30.1240 65.6235 30.1500 66.7170 ;
        RECT 30.0160 65.6235 30.0420 66.7170 ;
        RECT 29.9080 65.6235 29.9340 66.7170 ;
        RECT 29.8000 65.6235 29.8260 66.7170 ;
        RECT 29.6920 65.6235 29.7180 66.7170 ;
        RECT 29.5840 65.6235 29.6100 66.7170 ;
        RECT 29.4760 65.6235 29.5020 66.7170 ;
        RECT 29.3680 65.6235 29.3940 66.7170 ;
        RECT 29.2600 65.6235 29.2860 66.7170 ;
        RECT 29.1520 65.6235 29.1780 66.7170 ;
        RECT 29.0440 65.6235 29.0700 66.7170 ;
        RECT 28.9360 65.6235 28.9620 66.7170 ;
        RECT 28.8280 65.6235 28.8540 66.7170 ;
        RECT 28.7200 65.6235 28.7460 66.7170 ;
        RECT 28.6120 65.6235 28.6380 66.7170 ;
        RECT 28.5040 65.6235 28.5300 66.7170 ;
        RECT 28.3960 65.6235 28.4220 66.7170 ;
        RECT 28.2880 65.6235 28.3140 66.7170 ;
        RECT 28.1800 65.6235 28.2060 66.7170 ;
        RECT 28.0720 65.6235 28.0980 66.7170 ;
        RECT 27.9640 65.6235 27.9900 66.7170 ;
        RECT 27.8560 65.6235 27.8820 66.7170 ;
        RECT 27.7480 65.6235 27.7740 66.7170 ;
        RECT 27.6400 65.6235 27.6660 66.7170 ;
        RECT 27.5320 65.6235 27.5580 66.7170 ;
        RECT 27.4240 65.6235 27.4500 66.7170 ;
        RECT 27.3160 65.6235 27.3420 66.7170 ;
        RECT 27.2080 65.6235 27.2340 66.7170 ;
        RECT 27.1000 65.6235 27.1260 66.7170 ;
        RECT 26.9920 65.6235 27.0180 66.7170 ;
        RECT 26.8840 65.6235 26.9100 66.7170 ;
        RECT 26.7760 65.6235 26.8020 66.7170 ;
        RECT 26.6680 65.6235 26.6940 66.7170 ;
        RECT 26.5600 65.6235 26.5860 66.7170 ;
        RECT 26.4520 65.6235 26.4780 66.7170 ;
        RECT 26.3440 65.6235 26.3700 66.7170 ;
        RECT 26.2360 65.6235 26.2620 66.7170 ;
        RECT 26.1280 65.6235 26.1540 66.7170 ;
        RECT 26.0200 65.6235 26.0460 66.7170 ;
        RECT 25.9120 65.6235 25.9380 66.7170 ;
        RECT 25.8040 65.6235 25.8300 66.7170 ;
        RECT 25.6960 65.6235 25.7220 66.7170 ;
        RECT 25.5880 65.6235 25.6140 66.7170 ;
        RECT 25.4800 65.6235 25.5060 66.7170 ;
        RECT 25.3720 65.6235 25.3980 66.7170 ;
        RECT 25.2640 65.6235 25.2900 66.7170 ;
        RECT 25.1560 65.6235 25.1820 66.7170 ;
        RECT 25.0480 65.6235 25.0740 66.7170 ;
        RECT 24.9400 65.6235 24.9660 66.7170 ;
        RECT 24.8320 65.6235 24.8580 66.7170 ;
        RECT 24.7240 65.6235 24.7500 66.7170 ;
        RECT 24.6160 65.6235 24.6420 66.7170 ;
        RECT 24.5080 65.6235 24.5340 66.7170 ;
        RECT 24.4000 65.6235 24.4260 66.7170 ;
        RECT 24.2920 65.6235 24.3180 66.7170 ;
        RECT 24.1840 65.6235 24.2100 66.7170 ;
        RECT 24.0760 65.6235 24.1020 66.7170 ;
        RECT 23.9680 65.6235 23.9940 66.7170 ;
        RECT 23.8600 65.6235 23.8860 66.7170 ;
        RECT 23.7520 65.6235 23.7780 66.7170 ;
        RECT 23.6440 65.6235 23.6700 66.7170 ;
        RECT 23.5360 65.6235 23.5620 66.7170 ;
        RECT 23.4280 65.6235 23.4540 66.7170 ;
        RECT 23.3200 65.6235 23.3460 66.7170 ;
        RECT 23.2120 65.6235 23.2380 66.7170 ;
        RECT 23.1040 65.6235 23.1300 66.7170 ;
        RECT 22.9960 65.6235 23.0220 66.7170 ;
        RECT 22.8880 65.6235 22.9140 66.7170 ;
        RECT 22.7800 65.6235 22.8060 66.7170 ;
        RECT 22.6720 65.6235 22.6980 66.7170 ;
        RECT 22.5640 65.6235 22.5900 66.7170 ;
        RECT 22.4560 65.6235 22.4820 66.7170 ;
        RECT 22.3480 65.6235 22.3740 66.7170 ;
        RECT 22.2400 65.6235 22.2660 66.7170 ;
        RECT 22.1320 65.6235 22.1580 66.7170 ;
        RECT 22.0240 65.6235 22.0500 66.7170 ;
        RECT 21.9160 65.6235 21.9420 66.7170 ;
        RECT 21.8080 65.6235 21.8340 66.7170 ;
        RECT 21.7000 65.6235 21.7260 66.7170 ;
        RECT 21.5920 65.6235 21.6180 66.7170 ;
        RECT 21.4840 65.6235 21.5100 66.7170 ;
        RECT 21.3760 65.6235 21.4020 66.7170 ;
        RECT 21.2680 65.6235 21.2940 66.7170 ;
        RECT 21.1600 65.6235 21.1860 66.7170 ;
        RECT 21.0520 65.6235 21.0780 66.7170 ;
        RECT 20.9440 65.6235 20.9700 66.7170 ;
        RECT 20.8360 65.6235 20.8620 66.7170 ;
        RECT 20.7280 65.6235 20.7540 66.7170 ;
        RECT 20.6200 65.6235 20.6460 66.7170 ;
        RECT 20.5120 65.6235 20.5380 66.7170 ;
        RECT 20.4040 65.6235 20.4300 66.7170 ;
        RECT 20.2960 65.6235 20.3220 66.7170 ;
        RECT 20.1880 65.6235 20.2140 66.7170 ;
        RECT 20.0800 65.6235 20.1060 66.7170 ;
        RECT 19.9720 65.6235 19.9980 66.7170 ;
        RECT 19.8640 65.6235 19.8900 66.7170 ;
        RECT 19.7560 65.6235 19.7820 66.7170 ;
        RECT 19.6480 65.6235 19.6740 66.7170 ;
        RECT 19.5400 65.6235 19.5660 66.7170 ;
        RECT 19.4320 65.6235 19.4580 66.7170 ;
        RECT 19.3240 65.6235 19.3500 66.7170 ;
        RECT 19.2160 65.6235 19.2420 66.7170 ;
        RECT 19.1080 65.6235 19.1340 66.7170 ;
        RECT 19.0000 65.6235 19.0260 66.7170 ;
        RECT 18.8920 65.6235 18.9180 66.7170 ;
        RECT 18.7840 65.6235 18.8100 66.7170 ;
        RECT 18.6760 65.6235 18.7020 66.7170 ;
        RECT 18.5680 65.6235 18.5940 66.7170 ;
        RECT 18.4600 65.6235 18.4860 66.7170 ;
        RECT 18.3520 65.6235 18.3780 66.7170 ;
        RECT 18.2440 65.6235 18.2700 66.7170 ;
        RECT 18.1360 65.6235 18.1620 66.7170 ;
        RECT 18.0280 65.6235 18.0540 66.7170 ;
        RECT 17.9200 65.6235 17.9460 66.7170 ;
        RECT 17.8120 65.6235 17.8380 66.7170 ;
        RECT 17.7040 65.6235 17.7300 66.7170 ;
        RECT 17.5960 65.6235 17.6220 66.7170 ;
        RECT 17.4880 65.6235 17.5140 66.7170 ;
        RECT 17.3800 65.6235 17.4060 66.7170 ;
        RECT 17.2720 65.6235 17.2980 66.7170 ;
        RECT 17.1640 65.6235 17.1900 66.7170 ;
        RECT 17.0560 65.6235 17.0820 66.7170 ;
        RECT 16.9480 65.6235 16.9740 66.7170 ;
        RECT 16.8400 65.6235 16.8660 66.7170 ;
        RECT 16.7320 65.6235 16.7580 66.7170 ;
        RECT 16.6240 65.6235 16.6500 66.7170 ;
        RECT 16.5160 65.6235 16.5420 66.7170 ;
        RECT 16.4080 65.6235 16.4340 66.7170 ;
        RECT 16.3000 65.6235 16.3260 66.7170 ;
        RECT 16.0870 65.6235 16.1640 66.7170 ;
        RECT 14.1940 65.6235 14.2710 66.7170 ;
        RECT 14.0320 65.6235 14.0580 66.7170 ;
        RECT 13.9240 65.6235 13.9500 66.7170 ;
        RECT 13.8160 65.6235 13.8420 66.7170 ;
        RECT 13.7080 65.6235 13.7340 66.7170 ;
        RECT 13.6000 65.6235 13.6260 66.7170 ;
        RECT 13.4920 65.6235 13.5180 66.7170 ;
        RECT 13.3840 65.6235 13.4100 66.7170 ;
        RECT 13.2760 65.6235 13.3020 66.7170 ;
        RECT 13.1680 65.6235 13.1940 66.7170 ;
        RECT 13.0600 65.6235 13.0860 66.7170 ;
        RECT 12.9520 65.6235 12.9780 66.7170 ;
        RECT 12.8440 65.6235 12.8700 66.7170 ;
        RECT 12.7360 65.6235 12.7620 66.7170 ;
        RECT 12.6280 65.6235 12.6540 66.7170 ;
        RECT 12.5200 65.6235 12.5460 66.7170 ;
        RECT 12.4120 65.6235 12.4380 66.7170 ;
        RECT 12.3040 65.6235 12.3300 66.7170 ;
        RECT 12.1960 65.6235 12.2220 66.7170 ;
        RECT 12.0880 65.6235 12.1140 66.7170 ;
        RECT 11.9800 65.6235 12.0060 66.7170 ;
        RECT 11.8720 65.6235 11.8980 66.7170 ;
        RECT 11.7640 65.6235 11.7900 66.7170 ;
        RECT 11.6560 65.6235 11.6820 66.7170 ;
        RECT 11.5480 65.6235 11.5740 66.7170 ;
        RECT 11.4400 65.6235 11.4660 66.7170 ;
        RECT 11.3320 65.6235 11.3580 66.7170 ;
        RECT 11.2240 65.6235 11.2500 66.7170 ;
        RECT 11.1160 65.6235 11.1420 66.7170 ;
        RECT 11.0080 65.6235 11.0340 66.7170 ;
        RECT 10.9000 65.6235 10.9260 66.7170 ;
        RECT 10.7920 65.6235 10.8180 66.7170 ;
        RECT 10.6840 65.6235 10.7100 66.7170 ;
        RECT 10.5760 65.6235 10.6020 66.7170 ;
        RECT 10.4680 65.6235 10.4940 66.7170 ;
        RECT 10.3600 65.6235 10.3860 66.7170 ;
        RECT 10.2520 65.6235 10.2780 66.7170 ;
        RECT 10.1440 65.6235 10.1700 66.7170 ;
        RECT 10.0360 65.6235 10.0620 66.7170 ;
        RECT 9.9280 65.6235 9.9540 66.7170 ;
        RECT 9.8200 65.6235 9.8460 66.7170 ;
        RECT 9.7120 65.6235 9.7380 66.7170 ;
        RECT 9.6040 65.6235 9.6300 66.7170 ;
        RECT 9.4960 65.6235 9.5220 66.7170 ;
        RECT 9.3880 65.6235 9.4140 66.7170 ;
        RECT 9.2800 65.6235 9.3060 66.7170 ;
        RECT 9.1720 65.6235 9.1980 66.7170 ;
        RECT 9.0640 65.6235 9.0900 66.7170 ;
        RECT 8.9560 65.6235 8.9820 66.7170 ;
        RECT 8.8480 65.6235 8.8740 66.7170 ;
        RECT 8.7400 65.6235 8.7660 66.7170 ;
        RECT 8.6320 65.6235 8.6580 66.7170 ;
        RECT 8.5240 65.6235 8.5500 66.7170 ;
        RECT 8.4160 65.6235 8.4420 66.7170 ;
        RECT 8.3080 65.6235 8.3340 66.7170 ;
        RECT 8.2000 65.6235 8.2260 66.7170 ;
        RECT 8.0920 65.6235 8.1180 66.7170 ;
        RECT 7.9840 65.6235 8.0100 66.7170 ;
        RECT 7.8760 65.6235 7.9020 66.7170 ;
        RECT 7.7680 65.6235 7.7940 66.7170 ;
        RECT 7.6600 65.6235 7.6860 66.7170 ;
        RECT 7.5520 65.6235 7.5780 66.7170 ;
        RECT 7.4440 65.6235 7.4700 66.7170 ;
        RECT 7.3360 65.6235 7.3620 66.7170 ;
        RECT 7.2280 65.6235 7.2540 66.7170 ;
        RECT 7.1200 65.6235 7.1460 66.7170 ;
        RECT 7.0120 65.6235 7.0380 66.7170 ;
        RECT 6.9040 65.6235 6.9300 66.7170 ;
        RECT 6.7960 65.6235 6.8220 66.7170 ;
        RECT 6.6880 65.6235 6.7140 66.7170 ;
        RECT 6.5800 65.6235 6.6060 66.7170 ;
        RECT 6.4720 65.6235 6.4980 66.7170 ;
        RECT 6.3640 65.6235 6.3900 66.7170 ;
        RECT 6.2560 65.6235 6.2820 66.7170 ;
        RECT 6.1480 65.6235 6.1740 66.7170 ;
        RECT 6.0400 65.6235 6.0660 66.7170 ;
        RECT 5.9320 65.6235 5.9580 66.7170 ;
        RECT 5.8240 65.6235 5.8500 66.7170 ;
        RECT 5.7160 65.6235 5.7420 66.7170 ;
        RECT 5.6080 65.6235 5.6340 66.7170 ;
        RECT 5.5000 65.6235 5.5260 66.7170 ;
        RECT 5.3920 65.6235 5.4180 66.7170 ;
        RECT 5.2840 65.6235 5.3100 66.7170 ;
        RECT 5.1760 65.6235 5.2020 66.7170 ;
        RECT 5.0680 65.6235 5.0940 66.7170 ;
        RECT 4.9600 65.6235 4.9860 66.7170 ;
        RECT 4.8520 65.6235 4.8780 66.7170 ;
        RECT 4.7440 65.6235 4.7700 66.7170 ;
        RECT 4.6360 65.6235 4.6620 66.7170 ;
        RECT 4.5280 65.6235 4.5540 66.7170 ;
        RECT 4.4200 65.6235 4.4460 66.7170 ;
        RECT 4.3120 65.6235 4.3380 66.7170 ;
        RECT 4.2040 65.6235 4.2300 66.7170 ;
        RECT 4.0960 65.6235 4.1220 66.7170 ;
        RECT 3.9880 65.6235 4.0140 66.7170 ;
        RECT 3.8800 65.6235 3.9060 66.7170 ;
        RECT 3.7720 65.6235 3.7980 66.7170 ;
        RECT 3.6640 65.6235 3.6900 66.7170 ;
        RECT 3.5560 65.6235 3.5820 66.7170 ;
        RECT 3.4480 65.6235 3.4740 66.7170 ;
        RECT 3.3400 65.6235 3.3660 66.7170 ;
        RECT 3.2320 65.6235 3.2580 66.7170 ;
        RECT 3.1240 65.6235 3.1500 66.7170 ;
        RECT 3.0160 65.6235 3.0420 66.7170 ;
        RECT 2.9080 65.6235 2.9340 66.7170 ;
        RECT 2.8000 65.6235 2.8260 66.7170 ;
        RECT 2.6920 65.6235 2.7180 66.7170 ;
        RECT 2.5840 65.6235 2.6100 66.7170 ;
        RECT 2.4760 65.6235 2.5020 66.7170 ;
        RECT 2.3680 65.6235 2.3940 66.7170 ;
        RECT 2.2600 65.6235 2.2860 66.7170 ;
        RECT 2.1520 65.6235 2.1780 66.7170 ;
        RECT 2.0440 65.6235 2.0700 66.7170 ;
        RECT 1.9360 65.6235 1.9620 66.7170 ;
        RECT 1.8280 65.6235 1.8540 66.7170 ;
        RECT 1.7200 65.6235 1.7460 66.7170 ;
        RECT 1.6120 65.6235 1.6380 66.7170 ;
        RECT 1.5040 65.6235 1.5300 66.7170 ;
        RECT 1.3960 65.6235 1.4220 66.7170 ;
        RECT 1.2880 65.6235 1.3140 66.7170 ;
        RECT 1.1800 65.6235 1.2060 66.7170 ;
        RECT 1.0720 65.6235 1.0980 66.7170 ;
        RECT 0.9640 65.6235 0.9900 66.7170 ;
        RECT 0.8560 65.6235 0.8820 66.7170 ;
        RECT 0.7480 65.6235 0.7740 66.7170 ;
        RECT 0.6400 65.6235 0.6660 66.7170 ;
        RECT 0.5320 65.6235 0.5580 66.7170 ;
        RECT 0.4240 65.6235 0.4500 66.7170 ;
        RECT 0.3160 65.6235 0.3420 66.7170 ;
        RECT 0.2080 65.6235 0.2340 66.7170 ;
        RECT 0.0050 65.6235 0.0900 66.7170 ;
        RECT 15.5530 66.7035 15.6810 67.7970 ;
        RECT 15.5390 67.3690 15.6810 67.6915 ;
        RECT 15.3190 67.0960 15.4530 67.7970 ;
        RECT 15.2960 67.4310 15.4530 67.6890 ;
        RECT 15.3190 66.7035 15.4170 67.7970 ;
        RECT 15.3190 66.8245 15.4310 67.0640 ;
        RECT 15.3190 66.7035 15.4530 66.7925 ;
        RECT 15.0940 67.1540 15.2280 67.7970 ;
        RECT 15.0940 66.7035 15.1920 67.7970 ;
        RECT 14.6770 66.7035 14.7600 67.7970 ;
        RECT 14.6770 66.7920 14.7740 67.7275 ;
        RECT 30.2680 66.7035 30.3530 67.7970 ;
        RECT 30.1240 66.7035 30.1500 67.7970 ;
        RECT 30.0160 66.7035 30.0420 67.7970 ;
        RECT 29.9080 66.7035 29.9340 67.7970 ;
        RECT 29.8000 66.7035 29.8260 67.7970 ;
        RECT 29.6920 66.7035 29.7180 67.7970 ;
        RECT 29.5840 66.7035 29.6100 67.7970 ;
        RECT 29.4760 66.7035 29.5020 67.7970 ;
        RECT 29.3680 66.7035 29.3940 67.7970 ;
        RECT 29.2600 66.7035 29.2860 67.7970 ;
        RECT 29.1520 66.7035 29.1780 67.7970 ;
        RECT 29.0440 66.7035 29.0700 67.7970 ;
        RECT 28.9360 66.7035 28.9620 67.7970 ;
        RECT 28.8280 66.7035 28.8540 67.7970 ;
        RECT 28.7200 66.7035 28.7460 67.7970 ;
        RECT 28.6120 66.7035 28.6380 67.7970 ;
        RECT 28.5040 66.7035 28.5300 67.7970 ;
        RECT 28.3960 66.7035 28.4220 67.7970 ;
        RECT 28.2880 66.7035 28.3140 67.7970 ;
        RECT 28.1800 66.7035 28.2060 67.7970 ;
        RECT 28.0720 66.7035 28.0980 67.7970 ;
        RECT 27.9640 66.7035 27.9900 67.7970 ;
        RECT 27.8560 66.7035 27.8820 67.7970 ;
        RECT 27.7480 66.7035 27.7740 67.7970 ;
        RECT 27.6400 66.7035 27.6660 67.7970 ;
        RECT 27.5320 66.7035 27.5580 67.7970 ;
        RECT 27.4240 66.7035 27.4500 67.7970 ;
        RECT 27.3160 66.7035 27.3420 67.7970 ;
        RECT 27.2080 66.7035 27.2340 67.7970 ;
        RECT 27.1000 66.7035 27.1260 67.7970 ;
        RECT 26.9920 66.7035 27.0180 67.7970 ;
        RECT 26.8840 66.7035 26.9100 67.7970 ;
        RECT 26.7760 66.7035 26.8020 67.7970 ;
        RECT 26.6680 66.7035 26.6940 67.7970 ;
        RECT 26.5600 66.7035 26.5860 67.7970 ;
        RECT 26.4520 66.7035 26.4780 67.7970 ;
        RECT 26.3440 66.7035 26.3700 67.7970 ;
        RECT 26.2360 66.7035 26.2620 67.7970 ;
        RECT 26.1280 66.7035 26.1540 67.7970 ;
        RECT 26.0200 66.7035 26.0460 67.7970 ;
        RECT 25.9120 66.7035 25.9380 67.7970 ;
        RECT 25.8040 66.7035 25.8300 67.7970 ;
        RECT 25.6960 66.7035 25.7220 67.7970 ;
        RECT 25.5880 66.7035 25.6140 67.7970 ;
        RECT 25.4800 66.7035 25.5060 67.7970 ;
        RECT 25.3720 66.7035 25.3980 67.7970 ;
        RECT 25.2640 66.7035 25.2900 67.7970 ;
        RECT 25.1560 66.7035 25.1820 67.7970 ;
        RECT 25.0480 66.7035 25.0740 67.7970 ;
        RECT 24.9400 66.7035 24.9660 67.7970 ;
        RECT 24.8320 66.7035 24.8580 67.7970 ;
        RECT 24.7240 66.7035 24.7500 67.7970 ;
        RECT 24.6160 66.7035 24.6420 67.7970 ;
        RECT 24.5080 66.7035 24.5340 67.7970 ;
        RECT 24.4000 66.7035 24.4260 67.7970 ;
        RECT 24.2920 66.7035 24.3180 67.7970 ;
        RECT 24.1840 66.7035 24.2100 67.7970 ;
        RECT 24.0760 66.7035 24.1020 67.7970 ;
        RECT 23.9680 66.7035 23.9940 67.7970 ;
        RECT 23.8600 66.7035 23.8860 67.7970 ;
        RECT 23.7520 66.7035 23.7780 67.7970 ;
        RECT 23.6440 66.7035 23.6700 67.7970 ;
        RECT 23.5360 66.7035 23.5620 67.7970 ;
        RECT 23.4280 66.7035 23.4540 67.7970 ;
        RECT 23.3200 66.7035 23.3460 67.7970 ;
        RECT 23.2120 66.7035 23.2380 67.7970 ;
        RECT 23.1040 66.7035 23.1300 67.7970 ;
        RECT 22.9960 66.7035 23.0220 67.7970 ;
        RECT 22.8880 66.7035 22.9140 67.7970 ;
        RECT 22.7800 66.7035 22.8060 67.7970 ;
        RECT 22.6720 66.7035 22.6980 67.7970 ;
        RECT 22.5640 66.7035 22.5900 67.7970 ;
        RECT 22.4560 66.7035 22.4820 67.7970 ;
        RECT 22.3480 66.7035 22.3740 67.7970 ;
        RECT 22.2400 66.7035 22.2660 67.7970 ;
        RECT 22.1320 66.7035 22.1580 67.7970 ;
        RECT 22.0240 66.7035 22.0500 67.7970 ;
        RECT 21.9160 66.7035 21.9420 67.7970 ;
        RECT 21.8080 66.7035 21.8340 67.7970 ;
        RECT 21.7000 66.7035 21.7260 67.7970 ;
        RECT 21.5920 66.7035 21.6180 67.7970 ;
        RECT 21.4840 66.7035 21.5100 67.7970 ;
        RECT 21.3760 66.7035 21.4020 67.7970 ;
        RECT 21.2680 66.7035 21.2940 67.7970 ;
        RECT 21.1600 66.7035 21.1860 67.7970 ;
        RECT 21.0520 66.7035 21.0780 67.7970 ;
        RECT 20.9440 66.7035 20.9700 67.7970 ;
        RECT 20.8360 66.7035 20.8620 67.7970 ;
        RECT 20.7280 66.7035 20.7540 67.7970 ;
        RECT 20.6200 66.7035 20.6460 67.7970 ;
        RECT 20.5120 66.7035 20.5380 67.7970 ;
        RECT 20.4040 66.7035 20.4300 67.7970 ;
        RECT 20.2960 66.7035 20.3220 67.7970 ;
        RECT 20.1880 66.7035 20.2140 67.7970 ;
        RECT 20.0800 66.7035 20.1060 67.7970 ;
        RECT 19.9720 66.7035 19.9980 67.7970 ;
        RECT 19.8640 66.7035 19.8900 67.7970 ;
        RECT 19.7560 66.7035 19.7820 67.7970 ;
        RECT 19.6480 66.7035 19.6740 67.7970 ;
        RECT 19.5400 66.7035 19.5660 67.7970 ;
        RECT 19.4320 66.7035 19.4580 67.7970 ;
        RECT 19.3240 66.7035 19.3500 67.7970 ;
        RECT 19.2160 66.7035 19.2420 67.7970 ;
        RECT 19.1080 66.7035 19.1340 67.7970 ;
        RECT 19.0000 66.7035 19.0260 67.7970 ;
        RECT 18.8920 66.7035 18.9180 67.7970 ;
        RECT 18.7840 66.7035 18.8100 67.7970 ;
        RECT 18.6760 66.7035 18.7020 67.7970 ;
        RECT 18.5680 66.7035 18.5940 67.7970 ;
        RECT 18.4600 66.7035 18.4860 67.7970 ;
        RECT 18.3520 66.7035 18.3780 67.7970 ;
        RECT 18.2440 66.7035 18.2700 67.7970 ;
        RECT 18.1360 66.7035 18.1620 67.7970 ;
        RECT 18.0280 66.7035 18.0540 67.7970 ;
        RECT 17.9200 66.7035 17.9460 67.7970 ;
        RECT 17.8120 66.7035 17.8380 67.7970 ;
        RECT 17.7040 66.7035 17.7300 67.7970 ;
        RECT 17.5960 66.7035 17.6220 67.7970 ;
        RECT 17.4880 66.7035 17.5140 67.7970 ;
        RECT 17.3800 66.7035 17.4060 67.7970 ;
        RECT 17.2720 66.7035 17.2980 67.7970 ;
        RECT 17.1640 66.7035 17.1900 67.7970 ;
        RECT 17.0560 66.7035 17.0820 67.7970 ;
        RECT 16.9480 66.7035 16.9740 67.7970 ;
        RECT 16.8400 66.7035 16.8660 67.7970 ;
        RECT 16.7320 66.7035 16.7580 67.7970 ;
        RECT 16.6240 66.7035 16.6500 67.7970 ;
        RECT 16.5160 66.7035 16.5420 67.7970 ;
        RECT 16.4080 66.7035 16.4340 67.7970 ;
        RECT 16.3000 66.7035 16.3260 67.7970 ;
        RECT 16.0870 66.7035 16.1640 67.7970 ;
        RECT 14.1940 66.7035 14.2710 67.7970 ;
        RECT 14.0320 66.7035 14.0580 67.7970 ;
        RECT 13.9240 66.7035 13.9500 67.7970 ;
        RECT 13.8160 66.7035 13.8420 67.7970 ;
        RECT 13.7080 66.7035 13.7340 67.7970 ;
        RECT 13.6000 66.7035 13.6260 67.7970 ;
        RECT 13.4920 66.7035 13.5180 67.7970 ;
        RECT 13.3840 66.7035 13.4100 67.7970 ;
        RECT 13.2760 66.7035 13.3020 67.7970 ;
        RECT 13.1680 66.7035 13.1940 67.7970 ;
        RECT 13.0600 66.7035 13.0860 67.7970 ;
        RECT 12.9520 66.7035 12.9780 67.7970 ;
        RECT 12.8440 66.7035 12.8700 67.7970 ;
        RECT 12.7360 66.7035 12.7620 67.7970 ;
        RECT 12.6280 66.7035 12.6540 67.7970 ;
        RECT 12.5200 66.7035 12.5460 67.7970 ;
        RECT 12.4120 66.7035 12.4380 67.7970 ;
        RECT 12.3040 66.7035 12.3300 67.7970 ;
        RECT 12.1960 66.7035 12.2220 67.7970 ;
        RECT 12.0880 66.7035 12.1140 67.7970 ;
        RECT 11.9800 66.7035 12.0060 67.7970 ;
        RECT 11.8720 66.7035 11.8980 67.7970 ;
        RECT 11.7640 66.7035 11.7900 67.7970 ;
        RECT 11.6560 66.7035 11.6820 67.7970 ;
        RECT 11.5480 66.7035 11.5740 67.7970 ;
        RECT 11.4400 66.7035 11.4660 67.7970 ;
        RECT 11.3320 66.7035 11.3580 67.7970 ;
        RECT 11.2240 66.7035 11.2500 67.7970 ;
        RECT 11.1160 66.7035 11.1420 67.7970 ;
        RECT 11.0080 66.7035 11.0340 67.7970 ;
        RECT 10.9000 66.7035 10.9260 67.7970 ;
        RECT 10.7920 66.7035 10.8180 67.7970 ;
        RECT 10.6840 66.7035 10.7100 67.7970 ;
        RECT 10.5760 66.7035 10.6020 67.7970 ;
        RECT 10.4680 66.7035 10.4940 67.7970 ;
        RECT 10.3600 66.7035 10.3860 67.7970 ;
        RECT 10.2520 66.7035 10.2780 67.7970 ;
        RECT 10.1440 66.7035 10.1700 67.7970 ;
        RECT 10.0360 66.7035 10.0620 67.7970 ;
        RECT 9.9280 66.7035 9.9540 67.7970 ;
        RECT 9.8200 66.7035 9.8460 67.7970 ;
        RECT 9.7120 66.7035 9.7380 67.7970 ;
        RECT 9.6040 66.7035 9.6300 67.7970 ;
        RECT 9.4960 66.7035 9.5220 67.7970 ;
        RECT 9.3880 66.7035 9.4140 67.7970 ;
        RECT 9.2800 66.7035 9.3060 67.7970 ;
        RECT 9.1720 66.7035 9.1980 67.7970 ;
        RECT 9.0640 66.7035 9.0900 67.7970 ;
        RECT 8.9560 66.7035 8.9820 67.7970 ;
        RECT 8.8480 66.7035 8.8740 67.7970 ;
        RECT 8.7400 66.7035 8.7660 67.7970 ;
        RECT 8.6320 66.7035 8.6580 67.7970 ;
        RECT 8.5240 66.7035 8.5500 67.7970 ;
        RECT 8.4160 66.7035 8.4420 67.7970 ;
        RECT 8.3080 66.7035 8.3340 67.7970 ;
        RECT 8.2000 66.7035 8.2260 67.7970 ;
        RECT 8.0920 66.7035 8.1180 67.7970 ;
        RECT 7.9840 66.7035 8.0100 67.7970 ;
        RECT 7.8760 66.7035 7.9020 67.7970 ;
        RECT 7.7680 66.7035 7.7940 67.7970 ;
        RECT 7.6600 66.7035 7.6860 67.7970 ;
        RECT 7.5520 66.7035 7.5780 67.7970 ;
        RECT 7.4440 66.7035 7.4700 67.7970 ;
        RECT 7.3360 66.7035 7.3620 67.7970 ;
        RECT 7.2280 66.7035 7.2540 67.7970 ;
        RECT 7.1200 66.7035 7.1460 67.7970 ;
        RECT 7.0120 66.7035 7.0380 67.7970 ;
        RECT 6.9040 66.7035 6.9300 67.7970 ;
        RECT 6.7960 66.7035 6.8220 67.7970 ;
        RECT 6.6880 66.7035 6.7140 67.7970 ;
        RECT 6.5800 66.7035 6.6060 67.7970 ;
        RECT 6.4720 66.7035 6.4980 67.7970 ;
        RECT 6.3640 66.7035 6.3900 67.7970 ;
        RECT 6.2560 66.7035 6.2820 67.7970 ;
        RECT 6.1480 66.7035 6.1740 67.7970 ;
        RECT 6.0400 66.7035 6.0660 67.7970 ;
        RECT 5.9320 66.7035 5.9580 67.7970 ;
        RECT 5.8240 66.7035 5.8500 67.7970 ;
        RECT 5.7160 66.7035 5.7420 67.7970 ;
        RECT 5.6080 66.7035 5.6340 67.7970 ;
        RECT 5.5000 66.7035 5.5260 67.7970 ;
        RECT 5.3920 66.7035 5.4180 67.7970 ;
        RECT 5.2840 66.7035 5.3100 67.7970 ;
        RECT 5.1760 66.7035 5.2020 67.7970 ;
        RECT 5.0680 66.7035 5.0940 67.7970 ;
        RECT 4.9600 66.7035 4.9860 67.7970 ;
        RECT 4.8520 66.7035 4.8780 67.7970 ;
        RECT 4.7440 66.7035 4.7700 67.7970 ;
        RECT 4.6360 66.7035 4.6620 67.7970 ;
        RECT 4.5280 66.7035 4.5540 67.7970 ;
        RECT 4.4200 66.7035 4.4460 67.7970 ;
        RECT 4.3120 66.7035 4.3380 67.7970 ;
        RECT 4.2040 66.7035 4.2300 67.7970 ;
        RECT 4.0960 66.7035 4.1220 67.7970 ;
        RECT 3.9880 66.7035 4.0140 67.7970 ;
        RECT 3.8800 66.7035 3.9060 67.7970 ;
        RECT 3.7720 66.7035 3.7980 67.7970 ;
        RECT 3.6640 66.7035 3.6900 67.7970 ;
        RECT 3.5560 66.7035 3.5820 67.7970 ;
        RECT 3.4480 66.7035 3.4740 67.7970 ;
        RECT 3.3400 66.7035 3.3660 67.7970 ;
        RECT 3.2320 66.7035 3.2580 67.7970 ;
        RECT 3.1240 66.7035 3.1500 67.7970 ;
        RECT 3.0160 66.7035 3.0420 67.7970 ;
        RECT 2.9080 66.7035 2.9340 67.7970 ;
        RECT 2.8000 66.7035 2.8260 67.7970 ;
        RECT 2.6920 66.7035 2.7180 67.7970 ;
        RECT 2.5840 66.7035 2.6100 67.7970 ;
        RECT 2.4760 66.7035 2.5020 67.7970 ;
        RECT 2.3680 66.7035 2.3940 67.7970 ;
        RECT 2.2600 66.7035 2.2860 67.7970 ;
        RECT 2.1520 66.7035 2.1780 67.7970 ;
        RECT 2.0440 66.7035 2.0700 67.7970 ;
        RECT 1.9360 66.7035 1.9620 67.7970 ;
        RECT 1.8280 66.7035 1.8540 67.7970 ;
        RECT 1.7200 66.7035 1.7460 67.7970 ;
        RECT 1.6120 66.7035 1.6380 67.7970 ;
        RECT 1.5040 66.7035 1.5300 67.7970 ;
        RECT 1.3960 66.7035 1.4220 67.7970 ;
        RECT 1.2880 66.7035 1.3140 67.7970 ;
        RECT 1.1800 66.7035 1.2060 67.7970 ;
        RECT 1.0720 66.7035 1.0980 67.7970 ;
        RECT 0.9640 66.7035 0.9900 67.7970 ;
        RECT 0.8560 66.7035 0.8820 67.7970 ;
        RECT 0.7480 66.7035 0.7740 67.7970 ;
        RECT 0.6400 66.7035 0.6660 67.7970 ;
        RECT 0.5320 66.7035 0.5580 67.7970 ;
        RECT 0.4240 66.7035 0.4500 67.7970 ;
        RECT 0.3160 66.7035 0.3420 67.7970 ;
        RECT 0.2080 66.7035 0.2340 67.7970 ;
        RECT 0.0050 66.7035 0.0900 67.7970 ;
        RECT 15.5530 67.7835 15.6810 68.8770 ;
        RECT 15.5390 68.4490 15.6810 68.7715 ;
        RECT 15.3190 68.1760 15.4530 68.8770 ;
        RECT 15.2960 68.5110 15.4530 68.7690 ;
        RECT 15.3190 67.7835 15.4170 68.8770 ;
        RECT 15.3190 67.9045 15.4310 68.1440 ;
        RECT 15.3190 67.7835 15.4530 67.8725 ;
        RECT 15.0940 68.2340 15.2280 68.8770 ;
        RECT 15.0940 67.7835 15.1920 68.8770 ;
        RECT 14.6770 67.7835 14.7600 68.8770 ;
        RECT 14.6770 67.8720 14.7740 68.8075 ;
        RECT 30.2680 67.7835 30.3530 68.8770 ;
        RECT 30.1240 67.7835 30.1500 68.8770 ;
        RECT 30.0160 67.7835 30.0420 68.8770 ;
        RECT 29.9080 67.7835 29.9340 68.8770 ;
        RECT 29.8000 67.7835 29.8260 68.8770 ;
        RECT 29.6920 67.7835 29.7180 68.8770 ;
        RECT 29.5840 67.7835 29.6100 68.8770 ;
        RECT 29.4760 67.7835 29.5020 68.8770 ;
        RECT 29.3680 67.7835 29.3940 68.8770 ;
        RECT 29.2600 67.7835 29.2860 68.8770 ;
        RECT 29.1520 67.7835 29.1780 68.8770 ;
        RECT 29.0440 67.7835 29.0700 68.8770 ;
        RECT 28.9360 67.7835 28.9620 68.8770 ;
        RECT 28.8280 67.7835 28.8540 68.8770 ;
        RECT 28.7200 67.7835 28.7460 68.8770 ;
        RECT 28.6120 67.7835 28.6380 68.8770 ;
        RECT 28.5040 67.7835 28.5300 68.8770 ;
        RECT 28.3960 67.7835 28.4220 68.8770 ;
        RECT 28.2880 67.7835 28.3140 68.8770 ;
        RECT 28.1800 67.7835 28.2060 68.8770 ;
        RECT 28.0720 67.7835 28.0980 68.8770 ;
        RECT 27.9640 67.7835 27.9900 68.8770 ;
        RECT 27.8560 67.7835 27.8820 68.8770 ;
        RECT 27.7480 67.7835 27.7740 68.8770 ;
        RECT 27.6400 67.7835 27.6660 68.8770 ;
        RECT 27.5320 67.7835 27.5580 68.8770 ;
        RECT 27.4240 67.7835 27.4500 68.8770 ;
        RECT 27.3160 67.7835 27.3420 68.8770 ;
        RECT 27.2080 67.7835 27.2340 68.8770 ;
        RECT 27.1000 67.7835 27.1260 68.8770 ;
        RECT 26.9920 67.7835 27.0180 68.8770 ;
        RECT 26.8840 67.7835 26.9100 68.8770 ;
        RECT 26.7760 67.7835 26.8020 68.8770 ;
        RECT 26.6680 67.7835 26.6940 68.8770 ;
        RECT 26.5600 67.7835 26.5860 68.8770 ;
        RECT 26.4520 67.7835 26.4780 68.8770 ;
        RECT 26.3440 67.7835 26.3700 68.8770 ;
        RECT 26.2360 67.7835 26.2620 68.8770 ;
        RECT 26.1280 67.7835 26.1540 68.8770 ;
        RECT 26.0200 67.7835 26.0460 68.8770 ;
        RECT 25.9120 67.7835 25.9380 68.8770 ;
        RECT 25.8040 67.7835 25.8300 68.8770 ;
        RECT 25.6960 67.7835 25.7220 68.8770 ;
        RECT 25.5880 67.7835 25.6140 68.8770 ;
        RECT 25.4800 67.7835 25.5060 68.8770 ;
        RECT 25.3720 67.7835 25.3980 68.8770 ;
        RECT 25.2640 67.7835 25.2900 68.8770 ;
        RECT 25.1560 67.7835 25.1820 68.8770 ;
        RECT 25.0480 67.7835 25.0740 68.8770 ;
        RECT 24.9400 67.7835 24.9660 68.8770 ;
        RECT 24.8320 67.7835 24.8580 68.8770 ;
        RECT 24.7240 67.7835 24.7500 68.8770 ;
        RECT 24.6160 67.7835 24.6420 68.8770 ;
        RECT 24.5080 67.7835 24.5340 68.8770 ;
        RECT 24.4000 67.7835 24.4260 68.8770 ;
        RECT 24.2920 67.7835 24.3180 68.8770 ;
        RECT 24.1840 67.7835 24.2100 68.8770 ;
        RECT 24.0760 67.7835 24.1020 68.8770 ;
        RECT 23.9680 67.7835 23.9940 68.8770 ;
        RECT 23.8600 67.7835 23.8860 68.8770 ;
        RECT 23.7520 67.7835 23.7780 68.8770 ;
        RECT 23.6440 67.7835 23.6700 68.8770 ;
        RECT 23.5360 67.7835 23.5620 68.8770 ;
        RECT 23.4280 67.7835 23.4540 68.8770 ;
        RECT 23.3200 67.7835 23.3460 68.8770 ;
        RECT 23.2120 67.7835 23.2380 68.8770 ;
        RECT 23.1040 67.7835 23.1300 68.8770 ;
        RECT 22.9960 67.7835 23.0220 68.8770 ;
        RECT 22.8880 67.7835 22.9140 68.8770 ;
        RECT 22.7800 67.7835 22.8060 68.8770 ;
        RECT 22.6720 67.7835 22.6980 68.8770 ;
        RECT 22.5640 67.7835 22.5900 68.8770 ;
        RECT 22.4560 67.7835 22.4820 68.8770 ;
        RECT 22.3480 67.7835 22.3740 68.8770 ;
        RECT 22.2400 67.7835 22.2660 68.8770 ;
        RECT 22.1320 67.7835 22.1580 68.8770 ;
        RECT 22.0240 67.7835 22.0500 68.8770 ;
        RECT 21.9160 67.7835 21.9420 68.8770 ;
        RECT 21.8080 67.7835 21.8340 68.8770 ;
        RECT 21.7000 67.7835 21.7260 68.8770 ;
        RECT 21.5920 67.7835 21.6180 68.8770 ;
        RECT 21.4840 67.7835 21.5100 68.8770 ;
        RECT 21.3760 67.7835 21.4020 68.8770 ;
        RECT 21.2680 67.7835 21.2940 68.8770 ;
        RECT 21.1600 67.7835 21.1860 68.8770 ;
        RECT 21.0520 67.7835 21.0780 68.8770 ;
        RECT 20.9440 67.7835 20.9700 68.8770 ;
        RECT 20.8360 67.7835 20.8620 68.8770 ;
        RECT 20.7280 67.7835 20.7540 68.8770 ;
        RECT 20.6200 67.7835 20.6460 68.8770 ;
        RECT 20.5120 67.7835 20.5380 68.8770 ;
        RECT 20.4040 67.7835 20.4300 68.8770 ;
        RECT 20.2960 67.7835 20.3220 68.8770 ;
        RECT 20.1880 67.7835 20.2140 68.8770 ;
        RECT 20.0800 67.7835 20.1060 68.8770 ;
        RECT 19.9720 67.7835 19.9980 68.8770 ;
        RECT 19.8640 67.7835 19.8900 68.8770 ;
        RECT 19.7560 67.7835 19.7820 68.8770 ;
        RECT 19.6480 67.7835 19.6740 68.8770 ;
        RECT 19.5400 67.7835 19.5660 68.8770 ;
        RECT 19.4320 67.7835 19.4580 68.8770 ;
        RECT 19.3240 67.7835 19.3500 68.8770 ;
        RECT 19.2160 67.7835 19.2420 68.8770 ;
        RECT 19.1080 67.7835 19.1340 68.8770 ;
        RECT 19.0000 67.7835 19.0260 68.8770 ;
        RECT 18.8920 67.7835 18.9180 68.8770 ;
        RECT 18.7840 67.7835 18.8100 68.8770 ;
        RECT 18.6760 67.7835 18.7020 68.8770 ;
        RECT 18.5680 67.7835 18.5940 68.8770 ;
        RECT 18.4600 67.7835 18.4860 68.8770 ;
        RECT 18.3520 67.7835 18.3780 68.8770 ;
        RECT 18.2440 67.7835 18.2700 68.8770 ;
        RECT 18.1360 67.7835 18.1620 68.8770 ;
        RECT 18.0280 67.7835 18.0540 68.8770 ;
        RECT 17.9200 67.7835 17.9460 68.8770 ;
        RECT 17.8120 67.7835 17.8380 68.8770 ;
        RECT 17.7040 67.7835 17.7300 68.8770 ;
        RECT 17.5960 67.7835 17.6220 68.8770 ;
        RECT 17.4880 67.7835 17.5140 68.8770 ;
        RECT 17.3800 67.7835 17.4060 68.8770 ;
        RECT 17.2720 67.7835 17.2980 68.8770 ;
        RECT 17.1640 67.7835 17.1900 68.8770 ;
        RECT 17.0560 67.7835 17.0820 68.8770 ;
        RECT 16.9480 67.7835 16.9740 68.8770 ;
        RECT 16.8400 67.7835 16.8660 68.8770 ;
        RECT 16.7320 67.7835 16.7580 68.8770 ;
        RECT 16.6240 67.7835 16.6500 68.8770 ;
        RECT 16.5160 67.7835 16.5420 68.8770 ;
        RECT 16.4080 67.7835 16.4340 68.8770 ;
        RECT 16.3000 67.7835 16.3260 68.8770 ;
        RECT 16.0870 67.7835 16.1640 68.8770 ;
        RECT 14.1940 67.7835 14.2710 68.8770 ;
        RECT 14.0320 67.7835 14.0580 68.8770 ;
        RECT 13.9240 67.7835 13.9500 68.8770 ;
        RECT 13.8160 67.7835 13.8420 68.8770 ;
        RECT 13.7080 67.7835 13.7340 68.8770 ;
        RECT 13.6000 67.7835 13.6260 68.8770 ;
        RECT 13.4920 67.7835 13.5180 68.8770 ;
        RECT 13.3840 67.7835 13.4100 68.8770 ;
        RECT 13.2760 67.7835 13.3020 68.8770 ;
        RECT 13.1680 67.7835 13.1940 68.8770 ;
        RECT 13.0600 67.7835 13.0860 68.8770 ;
        RECT 12.9520 67.7835 12.9780 68.8770 ;
        RECT 12.8440 67.7835 12.8700 68.8770 ;
        RECT 12.7360 67.7835 12.7620 68.8770 ;
        RECT 12.6280 67.7835 12.6540 68.8770 ;
        RECT 12.5200 67.7835 12.5460 68.8770 ;
        RECT 12.4120 67.7835 12.4380 68.8770 ;
        RECT 12.3040 67.7835 12.3300 68.8770 ;
        RECT 12.1960 67.7835 12.2220 68.8770 ;
        RECT 12.0880 67.7835 12.1140 68.8770 ;
        RECT 11.9800 67.7835 12.0060 68.8770 ;
        RECT 11.8720 67.7835 11.8980 68.8770 ;
        RECT 11.7640 67.7835 11.7900 68.8770 ;
        RECT 11.6560 67.7835 11.6820 68.8770 ;
        RECT 11.5480 67.7835 11.5740 68.8770 ;
        RECT 11.4400 67.7835 11.4660 68.8770 ;
        RECT 11.3320 67.7835 11.3580 68.8770 ;
        RECT 11.2240 67.7835 11.2500 68.8770 ;
        RECT 11.1160 67.7835 11.1420 68.8770 ;
        RECT 11.0080 67.7835 11.0340 68.8770 ;
        RECT 10.9000 67.7835 10.9260 68.8770 ;
        RECT 10.7920 67.7835 10.8180 68.8770 ;
        RECT 10.6840 67.7835 10.7100 68.8770 ;
        RECT 10.5760 67.7835 10.6020 68.8770 ;
        RECT 10.4680 67.7835 10.4940 68.8770 ;
        RECT 10.3600 67.7835 10.3860 68.8770 ;
        RECT 10.2520 67.7835 10.2780 68.8770 ;
        RECT 10.1440 67.7835 10.1700 68.8770 ;
        RECT 10.0360 67.7835 10.0620 68.8770 ;
        RECT 9.9280 67.7835 9.9540 68.8770 ;
        RECT 9.8200 67.7835 9.8460 68.8770 ;
        RECT 9.7120 67.7835 9.7380 68.8770 ;
        RECT 9.6040 67.7835 9.6300 68.8770 ;
        RECT 9.4960 67.7835 9.5220 68.8770 ;
        RECT 9.3880 67.7835 9.4140 68.8770 ;
        RECT 9.2800 67.7835 9.3060 68.8770 ;
        RECT 9.1720 67.7835 9.1980 68.8770 ;
        RECT 9.0640 67.7835 9.0900 68.8770 ;
        RECT 8.9560 67.7835 8.9820 68.8770 ;
        RECT 8.8480 67.7835 8.8740 68.8770 ;
        RECT 8.7400 67.7835 8.7660 68.8770 ;
        RECT 8.6320 67.7835 8.6580 68.8770 ;
        RECT 8.5240 67.7835 8.5500 68.8770 ;
        RECT 8.4160 67.7835 8.4420 68.8770 ;
        RECT 8.3080 67.7835 8.3340 68.8770 ;
        RECT 8.2000 67.7835 8.2260 68.8770 ;
        RECT 8.0920 67.7835 8.1180 68.8770 ;
        RECT 7.9840 67.7835 8.0100 68.8770 ;
        RECT 7.8760 67.7835 7.9020 68.8770 ;
        RECT 7.7680 67.7835 7.7940 68.8770 ;
        RECT 7.6600 67.7835 7.6860 68.8770 ;
        RECT 7.5520 67.7835 7.5780 68.8770 ;
        RECT 7.4440 67.7835 7.4700 68.8770 ;
        RECT 7.3360 67.7835 7.3620 68.8770 ;
        RECT 7.2280 67.7835 7.2540 68.8770 ;
        RECT 7.1200 67.7835 7.1460 68.8770 ;
        RECT 7.0120 67.7835 7.0380 68.8770 ;
        RECT 6.9040 67.7835 6.9300 68.8770 ;
        RECT 6.7960 67.7835 6.8220 68.8770 ;
        RECT 6.6880 67.7835 6.7140 68.8770 ;
        RECT 6.5800 67.7835 6.6060 68.8770 ;
        RECT 6.4720 67.7835 6.4980 68.8770 ;
        RECT 6.3640 67.7835 6.3900 68.8770 ;
        RECT 6.2560 67.7835 6.2820 68.8770 ;
        RECT 6.1480 67.7835 6.1740 68.8770 ;
        RECT 6.0400 67.7835 6.0660 68.8770 ;
        RECT 5.9320 67.7835 5.9580 68.8770 ;
        RECT 5.8240 67.7835 5.8500 68.8770 ;
        RECT 5.7160 67.7835 5.7420 68.8770 ;
        RECT 5.6080 67.7835 5.6340 68.8770 ;
        RECT 5.5000 67.7835 5.5260 68.8770 ;
        RECT 5.3920 67.7835 5.4180 68.8770 ;
        RECT 5.2840 67.7835 5.3100 68.8770 ;
        RECT 5.1760 67.7835 5.2020 68.8770 ;
        RECT 5.0680 67.7835 5.0940 68.8770 ;
        RECT 4.9600 67.7835 4.9860 68.8770 ;
        RECT 4.8520 67.7835 4.8780 68.8770 ;
        RECT 4.7440 67.7835 4.7700 68.8770 ;
        RECT 4.6360 67.7835 4.6620 68.8770 ;
        RECT 4.5280 67.7835 4.5540 68.8770 ;
        RECT 4.4200 67.7835 4.4460 68.8770 ;
        RECT 4.3120 67.7835 4.3380 68.8770 ;
        RECT 4.2040 67.7835 4.2300 68.8770 ;
        RECT 4.0960 67.7835 4.1220 68.8770 ;
        RECT 3.9880 67.7835 4.0140 68.8770 ;
        RECT 3.8800 67.7835 3.9060 68.8770 ;
        RECT 3.7720 67.7835 3.7980 68.8770 ;
        RECT 3.6640 67.7835 3.6900 68.8770 ;
        RECT 3.5560 67.7835 3.5820 68.8770 ;
        RECT 3.4480 67.7835 3.4740 68.8770 ;
        RECT 3.3400 67.7835 3.3660 68.8770 ;
        RECT 3.2320 67.7835 3.2580 68.8770 ;
        RECT 3.1240 67.7835 3.1500 68.8770 ;
        RECT 3.0160 67.7835 3.0420 68.8770 ;
        RECT 2.9080 67.7835 2.9340 68.8770 ;
        RECT 2.8000 67.7835 2.8260 68.8770 ;
        RECT 2.6920 67.7835 2.7180 68.8770 ;
        RECT 2.5840 67.7835 2.6100 68.8770 ;
        RECT 2.4760 67.7835 2.5020 68.8770 ;
        RECT 2.3680 67.7835 2.3940 68.8770 ;
        RECT 2.2600 67.7835 2.2860 68.8770 ;
        RECT 2.1520 67.7835 2.1780 68.8770 ;
        RECT 2.0440 67.7835 2.0700 68.8770 ;
        RECT 1.9360 67.7835 1.9620 68.8770 ;
        RECT 1.8280 67.7835 1.8540 68.8770 ;
        RECT 1.7200 67.7835 1.7460 68.8770 ;
        RECT 1.6120 67.7835 1.6380 68.8770 ;
        RECT 1.5040 67.7835 1.5300 68.8770 ;
        RECT 1.3960 67.7835 1.4220 68.8770 ;
        RECT 1.2880 67.7835 1.3140 68.8770 ;
        RECT 1.1800 67.7835 1.2060 68.8770 ;
        RECT 1.0720 67.7835 1.0980 68.8770 ;
        RECT 0.9640 67.7835 0.9900 68.8770 ;
        RECT 0.8560 67.7835 0.8820 68.8770 ;
        RECT 0.7480 67.7835 0.7740 68.8770 ;
        RECT 0.6400 67.7835 0.6660 68.8770 ;
        RECT 0.5320 67.7835 0.5580 68.8770 ;
        RECT 0.4240 67.7835 0.4500 68.8770 ;
        RECT 0.3160 67.7835 0.3420 68.8770 ;
        RECT 0.2080 67.7835 0.2340 68.8770 ;
        RECT 0.0050 67.7835 0.0900 68.8770 ;
        RECT 15.5530 68.8635 15.6810 69.9570 ;
        RECT 15.5390 69.5290 15.6810 69.8515 ;
        RECT 15.3190 69.2560 15.4530 69.9570 ;
        RECT 15.2960 69.5910 15.4530 69.8490 ;
        RECT 15.3190 68.8635 15.4170 69.9570 ;
        RECT 15.3190 68.9845 15.4310 69.2240 ;
        RECT 15.3190 68.8635 15.4530 68.9525 ;
        RECT 15.0940 69.3140 15.2280 69.9570 ;
        RECT 15.0940 68.8635 15.1920 69.9570 ;
        RECT 14.6770 68.8635 14.7600 69.9570 ;
        RECT 14.6770 68.9520 14.7740 69.8875 ;
        RECT 30.2680 68.8635 30.3530 69.9570 ;
        RECT 30.1240 68.8635 30.1500 69.9570 ;
        RECT 30.0160 68.8635 30.0420 69.9570 ;
        RECT 29.9080 68.8635 29.9340 69.9570 ;
        RECT 29.8000 68.8635 29.8260 69.9570 ;
        RECT 29.6920 68.8635 29.7180 69.9570 ;
        RECT 29.5840 68.8635 29.6100 69.9570 ;
        RECT 29.4760 68.8635 29.5020 69.9570 ;
        RECT 29.3680 68.8635 29.3940 69.9570 ;
        RECT 29.2600 68.8635 29.2860 69.9570 ;
        RECT 29.1520 68.8635 29.1780 69.9570 ;
        RECT 29.0440 68.8635 29.0700 69.9570 ;
        RECT 28.9360 68.8635 28.9620 69.9570 ;
        RECT 28.8280 68.8635 28.8540 69.9570 ;
        RECT 28.7200 68.8635 28.7460 69.9570 ;
        RECT 28.6120 68.8635 28.6380 69.9570 ;
        RECT 28.5040 68.8635 28.5300 69.9570 ;
        RECT 28.3960 68.8635 28.4220 69.9570 ;
        RECT 28.2880 68.8635 28.3140 69.9570 ;
        RECT 28.1800 68.8635 28.2060 69.9570 ;
        RECT 28.0720 68.8635 28.0980 69.9570 ;
        RECT 27.9640 68.8635 27.9900 69.9570 ;
        RECT 27.8560 68.8635 27.8820 69.9570 ;
        RECT 27.7480 68.8635 27.7740 69.9570 ;
        RECT 27.6400 68.8635 27.6660 69.9570 ;
        RECT 27.5320 68.8635 27.5580 69.9570 ;
        RECT 27.4240 68.8635 27.4500 69.9570 ;
        RECT 27.3160 68.8635 27.3420 69.9570 ;
        RECT 27.2080 68.8635 27.2340 69.9570 ;
        RECT 27.1000 68.8635 27.1260 69.9570 ;
        RECT 26.9920 68.8635 27.0180 69.9570 ;
        RECT 26.8840 68.8635 26.9100 69.9570 ;
        RECT 26.7760 68.8635 26.8020 69.9570 ;
        RECT 26.6680 68.8635 26.6940 69.9570 ;
        RECT 26.5600 68.8635 26.5860 69.9570 ;
        RECT 26.4520 68.8635 26.4780 69.9570 ;
        RECT 26.3440 68.8635 26.3700 69.9570 ;
        RECT 26.2360 68.8635 26.2620 69.9570 ;
        RECT 26.1280 68.8635 26.1540 69.9570 ;
        RECT 26.0200 68.8635 26.0460 69.9570 ;
        RECT 25.9120 68.8635 25.9380 69.9570 ;
        RECT 25.8040 68.8635 25.8300 69.9570 ;
        RECT 25.6960 68.8635 25.7220 69.9570 ;
        RECT 25.5880 68.8635 25.6140 69.9570 ;
        RECT 25.4800 68.8635 25.5060 69.9570 ;
        RECT 25.3720 68.8635 25.3980 69.9570 ;
        RECT 25.2640 68.8635 25.2900 69.9570 ;
        RECT 25.1560 68.8635 25.1820 69.9570 ;
        RECT 25.0480 68.8635 25.0740 69.9570 ;
        RECT 24.9400 68.8635 24.9660 69.9570 ;
        RECT 24.8320 68.8635 24.8580 69.9570 ;
        RECT 24.7240 68.8635 24.7500 69.9570 ;
        RECT 24.6160 68.8635 24.6420 69.9570 ;
        RECT 24.5080 68.8635 24.5340 69.9570 ;
        RECT 24.4000 68.8635 24.4260 69.9570 ;
        RECT 24.2920 68.8635 24.3180 69.9570 ;
        RECT 24.1840 68.8635 24.2100 69.9570 ;
        RECT 24.0760 68.8635 24.1020 69.9570 ;
        RECT 23.9680 68.8635 23.9940 69.9570 ;
        RECT 23.8600 68.8635 23.8860 69.9570 ;
        RECT 23.7520 68.8635 23.7780 69.9570 ;
        RECT 23.6440 68.8635 23.6700 69.9570 ;
        RECT 23.5360 68.8635 23.5620 69.9570 ;
        RECT 23.4280 68.8635 23.4540 69.9570 ;
        RECT 23.3200 68.8635 23.3460 69.9570 ;
        RECT 23.2120 68.8635 23.2380 69.9570 ;
        RECT 23.1040 68.8635 23.1300 69.9570 ;
        RECT 22.9960 68.8635 23.0220 69.9570 ;
        RECT 22.8880 68.8635 22.9140 69.9570 ;
        RECT 22.7800 68.8635 22.8060 69.9570 ;
        RECT 22.6720 68.8635 22.6980 69.9570 ;
        RECT 22.5640 68.8635 22.5900 69.9570 ;
        RECT 22.4560 68.8635 22.4820 69.9570 ;
        RECT 22.3480 68.8635 22.3740 69.9570 ;
        RECT 22.2400 68.8635 22.2660 69.9570 ;
        RECT 22.1320 68.8635 22.1580 69.9570 ;
        RECT 22.0240 68.8635 22.0500 69.9570 ;
        RECT 21.9160 68.8635 21.9420 69.9570 ;
        RECT 21.8080 68.8635 21.8340 69.9570 ;
        RECT 21.7000 68.8635 21.7260 69.9570 ;
        RECT 21.5920 68.8635 21.6180 69.9570 ;
        RECT 21.4840 68.8635 21.5100 69.9570 ;
        RECT 21.3760 68.8635 21.4020 69.9570 ;
        RECT 21.2680 68.8635 21.2940 69.9570 ;
        RECT 21.1600 68.8635 21.1860 69.9570 ;
        RECT 21.0520 68.8635 21.0780 69.9570 ;
        RECT 20.9440 68.8635 20.9700 69.9570 ;
        RECT 20.8360 68.8635 20.8620 69.9570 ;
        RECT 20.7280 68.8635 20.7540 69.9570 ;
        RECT 20.6200 68.8635 20.6460 69.9570 ;
        RECT 20.5120 68.8635 20.5380 69.9570 ;
        RECT 20.4040 68.8635 20.4300 69.9570 ;
        RECT 20.2960 68.8635 20.3220 69.9570 ;
        RECT 20.1880 68.8635 20.2140 69.9570 ;
        RECT 20.0800 68.8635 20.1060 69.9570 ;
        RECT 19.9720 68.8635 19.9980 69.9570 ;
        RECT 19.8640 68.8635 19.8900 69.9570 ;
        RECT 19.7560 68.8635 19.7820 69.9570 ;
        RECT 19.6480 68.8635 19.6740 69.9570 ;
        RECT 19.5400 68.8635 19.5660 69.9570 ;
        RECT 19.4320 68.8635 19.4580 69.9570 ;
        RECT 19.3240 68.8635 19.3500 69.9570 ;
        RECT 19.2160 68.8635 19.2420 69.9570 ;
        RECT 19.1080 68.8635 19.1340 69.9570 ;
        RECT 19.0000 68.8635 19.0260 69.9570 ;
        RECT 18.8920 68.8635 18.9180 69.9570 ;
        RECT 18.7840 68.8635 18.8100 69.9570 ;
        RECT 18.6760 68.8635 18.7020 69.9570 ;
        RECT 18.5680 68.8635 18.5940 69.9570 ;
        RECT 18.4600 68.8635 18.4860 69.9570 ;
        RECT 18.3520 68.8635 18.3780 69.9570 ;
        RECT 18.2440 68.8635 18.2700 69.9570 ;
        RECT 18.1360 68.8635 18.1620 69.9570 ;
        RECT 18.0280 68.8635 18.0540 69.9570 ;
        RECT 17.9200 68.8635 17.9460 69.9570 ;
        RECT 17.8120 68.8635 17.8380 69.9570 ;
        RECT 17.7040 68.8635 17.7300 69.9570 ;
        RECT 17.5960 68.8635 17.6220 69.9570 ;
        RECT 17.4880 68.8635 17.5140 69.9570 ;
        RECT 17.3800 68.8635 17.4060 69.9570 ;
        RECT 17.2720 68.8635 17.2980 69.9570 ;
        RECT 17.1640 68.8635 17.1900 69.9570 ;
        RECT 17.0560 68.8635 17.0820 69.9570 ;
        RECT 16.9480 68.8635 16.9740 69.9570 ;
        RECT 16.8400 68.8635 16.8660 69.9570 ;
        RECT 16.7320 68.8635 16.7580 69.9570 ;
        RECT 16.6240 68.8635 16.6500 69.9570 ;
        RECT 16.5160 68.8635 16.5420 69.9570 ;
        RECT 16.4080 68.8635 16.4340 69.9570 ;
        RECT 16.3000 68.8635 16.3260 69.9570 ;
        RECT 16.0870 68.8635 16.1640 69.9570 ;
        RECT 14.1940 68.8635 14.2710 69.9570 ;
        RECT 14.0320 68.8635 14.0580 69.9570 ;
        RECT 13.9240 68.8635 13.9500 69.9570 ;
        RECT 13.8160 68.8635 13.8420 69.9570 ;
        RECT 13.7080 68.8635 13.7340 69.9570 ;
        RECT 13.6000 68.8635 13.6260 69.9570 ;
        RECT 13.4920 68.8635 13.5180 69.9570 ;
        RECT 13.3840 68.8635 13.4100 69.9570 ;
        RECT 13.2760 68.8635 13.3020 69.9570 ;
        RECT 13.1680 68.8635 13.1940 69.9570 ;
        RECT 13.0600 68.8635 13.0860 69.9570 ;
        RECT 12.9520 68.8635 12.9780 69.9570 ;
        RECT 12.8440 68.8635 12.8700 69.9570 ;
        RECT 12.7360 68.8635 12.7620 69.9570 ;
        RECT 12.6280 68.8635 12.6540 69.9570 ;
        RECT 12.5200 68.8635 12.5460 69.9570 ;
        RECT 12.4120 68.8635 12.4380 69.9570 ;
        RECT 12.3040 68.8635 12.3300 69.9570 ;
        RECT 12.1960 68.8635 12.2220 69.9570 ;
        RECT 12.0880 68.8635 12.1140 69.9570 ;
        RECT 11.9800 68.8635 12.0060 69.9570 ;
        RECT 11.8720 68.8635 11.8980 69.9570 ;
        RECT 11.7640 68.8635 11.7900 69.9570 ;
        RECT 11.6560 68.8635 11.6820 69.9570 ;
        RECT 11.5480 68.8635 11.5740 69.9570 ;
        RECT 11.4400 68.8635 11.4660 69.9570 ;
        RECT 11.3320 68.8635 11.3580 69.9570 ;
        RECT 11.2240 68.8635 11.2500 69.9570 ;
        RECT 11.1160 68.8635 11.1420 69.9570 ;
        RECT 11.0080 68.8635 11.0340 69.9570 ;
        RECT 10.9000 68.8635 10.9260 69.9570 ;
        RECT 10.7920 68.8635 10.8180 69.9570 ;
        RECT 10.6840 68.8635 10.7100 69.9570 ;
        RECT 10.5760 68.8635 10.6020 69.9570 ;
        RECT 10.4680 68.8635 10.4940 69.9570 ;
        RECT 10.3600 68.8635 10.3860 69.9570 ;
        RECT 10.2520 68.8635 10.2780 69.9570 ;
        RECT 10.1440 68.8635 10.1700 69.9570 ;
        RECT 10.0360 68.8635 10.0620 69.9570 ;
        RECT 9.9280 68.8635 9.9540 69.9570 ;
        RECT 9.8200 68.8635 9.8460 69.9570 ;
        RECT 9.7120 68.8635 9.7380 69.9570 ;
        RECT 9.6040 68.8635 9.6300 69.9570 ;
        RECT 9.4960 68.8635 9.5220 69.9570 ;
        RECT 9.3880 68.8635 9.4140 69.9570 ;
        RECT 9.2800 68.8635 9.3060 69.9570 ;
        RECT 9.1720 68.8635 9.1980 69.9570 ;
        RECT 9.0640 68.8635 9.0900 69.9570 ;
        RECT 8.9560 68.8635 8.9820 69.9570 ;
        RECT 8.8480 68.8635 8.8740 69.9570 ;
        RECT 8.7400 68.8635 8.7660 69.9570 ;
        RECT 8.6320 68.8635 8.6580 69.9570 ;
        RECT 8.5240 68.8635 8.5500 69.9570 ;
        RECT 8.4160 68.8635 8.4420 69.9570 ;
        RECT 8.3080 68.8635 8.3340 69.9570 ;
        RECT 8.2000 68.8635 8.2260 69.9570 ;
        RECT 8.0920 68.8635 8.1180 69.9570 ;
        RECT 7.9840 68.8635 8.0100 69.9570 ;
        RECT 7.8760 68.8635 7.9020 69.9570 ;
        RECT 7.7680 68.8635 7.7940 69.9570 ;
        RECT 7.6600 68.8635 7.6860 69.9570 ;
        RECT 7.5520 68.8635 7.5780 69.9570 ;
        RECT 7.4440 68.8635 7.4700 69.9570 ;
        RECT 7.3360 68.8635 7.3620 69.9570 ;
        RECT 7.2280 68.8635 7.2540 69.9570 ;
        RECT 7.1200 68.8635 7.1460 69.9570 ;
        RECT 7.0120 68.8635 7.0380 69.9570 ;
        RECT 6.9040 68.8635 6.9300 69.9570 ;
        RECT 6.7960 68.8635 6.8220 69.9570 ;
        RECT 6.6880 68.8635 6.7140 69.9570 ;
        RECT 6.5800 68.8635 6.6060 69.9570 ;
        RECT 6.4720 68.8635 6.4980 69.9570 ;
        RECT 6.3640 68.8635 6.3900 69.9570 ;
        RECT 6.2560 68.8635 6.2820 69.9570 ;
        RECT 6.1480 68.8635 6.1740 69.9570 ;
        RECT 6.0400 68.8635 6.0660 69.9570 ;
        RECT 5.9320 68.8635 5.9580 69.9570 ;
        RECT 5.8240 68.8635 5.8500 69.9570 ;
        RECT 5.7160 68.8635 5.7420 69.9570 ;
        RECT 5.6080 68.8635 5.6340 69.9570 ;
        RECT 5.5000 68.8635 5.5260 69.9570 ;
        RECT 5.3920 68.8635 5.4180 69.9570 ;
        RECT 5.2840 68.8635 5.3100 69.9570 ;
        RECT 5.1760 68.8635 5.2020 69.9570 ;
        RECT 5.0680 68.8635 5.0940 69.9570 ;
        RECT 4.9600 68.8635 4.9860 69.9570 ;
        RECT 4.8520 68.8635 4.8780 69.9570 ;
        RECT 4.7440 68.8635 4.7700 69.9570 ;
        RECT 4.6360 68.8635 4.6620 69.9570 ;
        RECT 4.5280 68.8635 4.5540 69.9570 ;
        RECT 4.4200 68.8635 4.4460 69.9570 ;
        RECT 4.3120 68.8635 4.3380 69.9570 ;
        RECT 4.2040 68.8635 4.2300 69.9570 ;
        RECT 4.0960 68.8635 4.1220 69.9570 ;
        RECT 3.9880 68.8635 4.0140 69.9570 ;
        RECT 3.8800 68.8635 3.9060 69.9570 ;
        RECT 3.7720 68.8635 3.7980 69.9570 ;
        RECT 3.6640 68.8635 3.6900 69.9570 ;
        RECT 3.5560 68.8635 3.5820 69.9570 ;
        RECT 3.4480 68.8635 3.4740 69.9570 ;
        RECT 3.3400 68.8635 3.3660 69.9570 ;
        RECT 3.2320 68.8635 3.2580 69.9570 ;
        RECT 3.1240 68.8635 3.1500 69.9570 ;
        RECT 3.0160 68.8635 3.0420 69.9570 ;
        RECT 2.9080 68.8635 2.9340 69.9570 ;
        RECT 2.8000 68.8635 2.8260 69.9570 ;
        RECT 2.6920 68.8635 2.7180 69.9570 ;
        RECT 2.5840 68.8635 2.6100 69.9570 ;
        RECT 2.4760 68.8635 2.5020 69.9570 ;
        RECT 2.3680 68.8635 2.3940 69.9570 ;
        RECT 2.2600 68.8635 2.2860 69.9570 ;
        RECT 2.1520 68.8635 2.1780 69.9570 ;
        RECT 2.0440 68.8635 2.0700 69.9570 ;
        RECT 1.9360 68.8635 1.9620 69.9570 ;
        RECT 1.8280 68.8635 1.8540 69.9570 ;
        RECT 1.7200 68.8635 1.7460 69.9570 ;
        RECT 1.6120 68.8635 1.6380 69.9570 ;
        RECT 1.5040 68.8635 1.5300 69.9570 ;
        RECT 1.3960 68.8635 1.4220 69.9570 ;
        RECT 1.2880 68.8635 1.3140 69.9570 ;
        RECT 1.1800 68.8635 1.2060 69.9570 ;
        RECT 1.0720 68.8635 1.0980 69.9570 ;
        RECT 0.9640 68.8635 0.9900 69.9570 ;
        RECT 0.8560 68.8635 0.8820 69.9570 ;
        RECT 0.7480 68.8635 0.7740 69.9570 ;
        RECT 0.6400 68.8635 0.6660 69.9570 ;
        RECT 0.5320 68.8635 0.5580 69.9570 ;
        RECT 0.4240 68.8635 0.4500 69.9570 ;
        RECT 0.3160 68.8635 0.3420 69.9570 ;
        RECT 0.2080 68.8635 0.2340 69.9570 ;
        RECT 0.0050 68.8635 0.0900 69.9570 ;
        RECT 15.5530 69.9435 15.6810 71.0370 ;
        RECT 15.5390 70.6090 15.6810 70.9315 ;
        RECT 15.3190 70.3360 15.4530 71.0370 ;
        RECT 15.2960 70.6710 15.4530 70.9290 ;
        RECT 15.3190 69.9435 15.4170 71.0370 ;
        RECT 15.3190 70.0645 15.4310 70.3040 ;
        RECT 15.3190 69.9435 15.4530 70.0325 ;
        RECT 15.0940 70.3940 15.2280 71.0370 ;
        RECT 15.0940 69.9435 15.1920 71.0370 ;
        RECT 14.6770 69.9435 14.7600 71.0370 ;
        RECT 14.6770 70.0320 14.7740 70.9675 ;
        RECT 30.2680 69.9435 30.3530 71.0370 ;
        RECT 30.1240 69.9435 30.1500 71.0370 ;
        RECT 30.0160 69.9435 30.0420 71.0370 ;
        RECT 29.9080 69.9435 29.9340 71.0370 ;
        RECT 29.8000 69.9435 29.8260 71.0370 ;
        RECT 29.6920 69.9435 29.7180 71.0370 ;
        RECT 29.5840 69.9435 29.6100 71.0370 ;
        RECT 29.4760 69.9435 29.5020 71.0370 ;
        RECT 29.3680 69.9435 29.3940 71.0370 ;
        RECT 29.2600 69.9435 29.2860 71.0370 ;
        RECT 29.1520 69.9435 29.1780 71.0370 ;
        RECT 29.0440 69.9435 29.0700 71.0370 ;
        RECT 28.9360 69.9435 28.9620 71.0370 ;
        RECT 28.8280 69.9435 28.8540 71.0370 ;
        RECT 28.7200 69.9435 28.7460 71.0370 ;
        RECT 28.6120 69.9435 28.6380 71.0370 ;
        RECT 28.5040 69.9435 28.5300 71.0370 ;
        RECT 28.3960 69.9435 28.4220 71.0370 ;
        RECT 28.2880 69.9435 28.3140 71.0370 ;
        RECT 28.1800 69.9435 28.2060 71.0370 ;
        RECT 28.0720 69.9435 28.0980 71.0370 ;
        RECT 27.9640 69.9435 27.9900 71.0370 ;
        RECT 27.8560 69.9435 27.8820 71.0370 ;
        RECT 27.7480 69.9435 27.7740 71.0370 ;
        RECT 27.6400 69.9435 27.6660 71.0370 ;
        RECT 27.5320 69.9435 27.5580 71.0370 ;
        RECT 27.4240 69.9435 27.4500 71.0370 ;
        RECT 27.3160 69.9435 27.3420 71.0370 ;
        RECT 27.2080 69.9435 27.2340 71.0370 ;
        RECT 27.1000 69.9435 27.1260 71.0370 ;
        RECT 26.9920 69.9435 27.0180 71.0370 ;
        RECT 26.8840 69.9435 26.9100 71.0370 ;
        RECT 26.7760 69.9435 26.8020 71.0370 ;
        RECT 26.6680 69.9435 26.6940 71.0370 ;
        RECT 26.5600 69.9435 26.5860 71.0370 ;
        RECT 26.4520 69.9435 26.4780 71.0370 ;
        RECT 26.3440 69.9435 26.3700 71.0370 ;
        RECT 26.2360 69.9435 26.2620 71.0370 ;
        RECT 26.1280 69.9435 26.1540 71.0370 ;
        RECT 26.0200 69.9435 26.0460 71.0370 ;
        RECT 25.9120 69.9435 25.9380 71.0370 ;
        RECT 25.8040 69.9435 25.8300 71.0370 ;
        RECT 25.6960 69.9435 25.7220 71.0370 ;
        RECT 25.5880 69.9435 25.6140 71.0370 ;
        RECT 25.4800 69.9435 25.5060 71.0370 ;
        RECT 25.3720 69.9435 25.3980 71.0370 ;
        RECT 25.2640 69.9435 25.2900 71.0370 ;
        RECT 25.1560 69.9435 25.1820 71.0370 ;
        RECT 25.0480 69.9435 25.0740 71.0370 ;
        RECT 24.9400 69.9435 24.9660 71.0370 ;
        RECT 24.8320 69.9435 24.8580 71.0370 ;
        RECT 24.7240 69.9435 24.7500 71.0370 ;
        RECT 24.6160 69.9435 24.6420 71.0370 ;
        RECT 24.5080 69.9435 24.5340 71.0370 ;
        RECT 24.4000 69.9435 24.4260 71.0370 ;
        RECT 24.2920 69.9435 24.3180 71.0370 ;
        RECT 24.1840 69.9435 24.2100 71.0370 ;
        RECT 24.0760 69.9435 24.1020 71.0370 ;
        RECT 23.9680 69.9435 23.9940 71.0370 ;
        RECT 23.8600 69.9435 23.8860 71.0370 ;
        RECT 23.7520 69.9435 23.7780 71.0370 ;
        RECT 23.6440 69.9435 23.6700 71.0370 ;
        RECT 23.5360 69.9435 23.5620 71.0370 ;
        RECT 23.4280 69.9435 23.4540 71.0370 ;
        RECT 23.3200 69.9435 23.3460 71.0370 ;
        RECT 23.2120 69.9435 23.2380 71.0370 ;
        RECT 23.1040 69.9435 23.1300 71.0370 ;
        RECT 22.9960 69.9435 23.0220 71.0370 ;
        RECT 22.8880 69.9435 22.9140 71.0370 ;
        RECT 22.7800 69.9435 22.8060 71.0370 ;
        RECT 22.6720 69.9435 22.6980 71.0370 ;
        RECT 22.5640 69.9435 22.5900 71.0370 ;
        RECT 22.4560 69.9435 22.4820 71.0370 ;
        RECT 22.3480 69.9435 22.3740 71.0370 ;
        RECT 22.2400 69.9435 22.2660 71.0370 ;
        RECT 22.1320 69.9435 22.1580 71.0370 ;
        RECT 22.0240 69.9435 22.0500 71.0370 ;
        RECT 21.9160 69.9435 21.9420 71.0370 ;
        RECT 21.8080 69.9435 21.8340 71.0370 ;
        RECT 21.7000 69.9435 21.7260 71.0370 ;
        RECT 21.5920 69.9435 21.6180 71.0370 ;
        RECT 21.4840 69.9435 21.5100 71.0370 ;
        RECT 21.3760 69.9435 21.4020 71.0370 ;
        RECT 21.2680 69.9435 21.2940 71.0370 ;
        RECT 21.1600 69.9435 21.1860 71.0370 ;
        RECT 21.0520 69.9435 21.0780 71.0370 ;
        RECT 20.9440 69.9435 20.9700 71.0370 ;
        RECT 20.8360 69.9435 20.8620 71.0370 ;
        RECT 20.7280 69.9435 20.7540 71.0370 ;
        RECT 20.6200 69.9435 20.6460 71.0370 ;
        RECT 20.5120 69.9435 20.5380 71.0370 ;
        RECT 20.4040 69.9435 20.4300 71.0370 ;
        RECT 20.2960 69.9435 20.3220 71.0370 ;
        RECT 20.1880 69.9435 20.2140 71.0370 ;
        RECT 20.0800 69.9435 20.1060 71.0370 ;
        RECT 19.9720 69.9435 19.9980 71.0370 ;
        RECT 19.8640 69.9435 19.8900 71.0370 ;
        RECT 19.7560 69.9435 19.7820 71.0370 ;
        RECT 19.6480 69.9435 19.6740 71.0370 ;
        RECT 19.5400 69.9435 19.5660 71.0370 ;
        RECT 19.4320 69.9435 19.4580 71.0370 ;
        RECT 19.3240 69.9435 19.3500 71.0370 ;
        RECT 19.2160 69.9435 19.2420 71.0370 ;
        RECT 19.1080 69.9435 19.1340 71.0370 ;
        RECT 19.0000 69.9435 19.0260 71.0370 ;
        RECT 18.8920 69.9435 18.9180 71.0370 ;
        RECT 18.7840 69.9435 18.8100 71.0370 ;
        RECT 18.6760 69.9435 18.7020 71.0370 ;
        RECT 18.5680 69.9435 18.5940 71.0370 ;
        RECT 18.4600 69.9435 18.4860 71.0370 ;
        RECT 18.3520 69.9435 18.3780 71.0370 ;
        RECT 18.2440 69.9435 18.2700 71.0370 ;
        RECT 18.1360 69.9435 18.1620 71.0370 ;
        RECT 18.0280 69.9435 18.0540 71.0370 ;
        RECT 17.9200 69.9435 17.9460 71.0370 ;
        RECT 17.8120 69.9435 17.8380 71.0370 ;
        RECT 17.7040 69.9435 17.7300 71.0370 ;
        RECT 17.5960 69.9435 17.6220 71.0370 ;
        RECT 17.4880 69.9435 17.5140 71.0370 ;
        RECT 17.3800 69.9435 17.4060 71.0370 ;
        RECT 17.2720 69.9435 17.2980 71.0370 ;
        RECT 17.1640 69.9435 17.1900 71.0370 ;
        RECT 17.0560 69.9435 17.0820 71.0370 ;
        RECT 16.9480 69.9435 16.9740 71.0370 ;
        RECT 16.8400 69.9435 16.8660 71.0370 ;
        RECT 16.7320 69.9435 16.7580 71.0370 ;
        RECT 16.6240 69.9435 16.6500 71.0370 ;
        RECT 16.5160 69.9435 16.5420 71.0370 ;
        RECT 16.4080 69.9435 16.4340 71.0370 ;
        RECT 16.3000 69.9435 16.3260 71.0370 ;
        RECT 16.0870 69.9435 16.1640 71.0370 ;
        RECT 14.1940 69.9435 14.2710 71.0370 ;
        RECT 14.0320 69.9435 14.0580 71.0370 ;
        RECT 13.9240 69.9435 13.9500 71.0370 ;
        RECT 13.8160 69.9435 13.8420 71.0370 ;
        RECT 13.7080 69.9435 13.7340 71.0370 ;
        RECT 13.6000 69.9435 13.6260 71.0370 ;
        RECT 13.4920 69.9435 13.5180 71.0370 ;
        RECT 13.3840 69.9435 13.4100 71.0370 ;
        RECT 13.2760 69.9435 13.3020 71.0370 ;
        RECT 13.1680 69.9435 13.1940 71.0370 ;
        RECT 13.0600 69.9435 13.0860 71.0370 ;
        RECT 12.9520 69.9435 12.9780 71.0370 ;
        RECT 12.8440 69.9435 12.8700 71.0370 ;
        RECT 12.7360 69.9435 12.7620 71.0370 ;
        RECT 12.6280 69.9435 12.6540 71.0370 ;
        RECT 12.5200 69.9435 12.5460 71.0370 ;
        RECT 12.4120 69.9435 12.4380 71.0370 ;
        RECT 12.3040 69.9435 12.3300 71.0370 ;
        RECT 12.1960 69.9435 12.2220 71.0370 ;
        RECT 12.0880 69.9435 12.1140 71.0370 ;
        RECT 11.9800 69.9435 12.0060 71.0370 ;
        RECT 11.8720 69.9435 11.8980 71.0370 ;
        RECT 11.7640 69.9435 11.7900 71.0370 ;
        RECT 11.6560 69.9435 11.6820 71.0370 ;
        RECT 11.5480 69.9435 11.5740 71.0370 ;
        RECT 11.4400 69.9435 11.4660 71.0370 ;
        RECT 11.3320 69.9435 11.3580 71.0370 ;
        RECT 11.2240 69.9435 11.2500 71.0370 ;
        RECT 11.1160 69.9435 11.1420 71.0370 ;
        RECT 11.0080 69.9435 11.0340 71.0370 ;
        RECT 10.9000 69.9435 10.9260 71.0370 ;
        RECT 10.7920 69.9435 10.8180 71.0370 ;
        RECT 10.6840 69.9435 10.7100 71.0370 ;
        RECT 10.5760 69.9435 10.6020 71.0370 ;
        RECT 10.4680 69.9435 10.4940 71.0370 ;
        RECT 10.3600 69.9435 10.3860 71.0370 ;
        RECT 10.2520 69.9435 10.2780 71.0370 ;
        RECT 10.1440 69.9435 10.1700 71.0370 ;
        RECT 10.0360 69.9435 10.0620 71.0370 ;
        RECT 9.9280 69.9435 9.9540 71.0370 ;
        RECT 9.8200 69.9435 9.8460 71.0370 ;
        RECT 9.7120 69.9435 9.7380 71.0370 ;
        RECT 9.6040 69.9435 9.6300 71.0370 ;
        RECT 9.4960 69.9435 9.5220 71.0370 ;
        RECT 9.3880 69.9435 9.4140 71.0370 ;
        RECT 9.2800 69.9435 9.3060 71.0370 ;
        RECT 9.1720 69.9435 9.1980 71.0370 ;
        RECT 9.0640 69.9435 9.0900 71.0370 ;
        RECT 8.9560 69.9435 8.9820 71.0370 ;
        RECT 8.8480 69.9435 8.8740 71.0370 ;
        RECT 8.7400 69.9435 8.7660 71.0370 ;
        RECT 8.6320 69.9435 8.6580 71.0370 ;
        RECT 8.5240 69.9435 8.5500 71.0370 ;
        RECT 8.4160 69.9435 8.4420 71.0370 ;
        RECT 8.3080 69.9435 8.3340 71.0370 ;
        RECT 8.2000 69.9435 8.2260 71.0370 ;
        RECT 8.0920 69.9435 8.1180 71.0370 ;
        RECT 7.9840 69.9435 8.0100 71.0370 ;
        RECT 7.8760 69.9435 7.9020 71.0370 ;
        RECT 7.7680 69.9435 7.7940 71.0370 ;
        RECT 7.6600 69.9435 7.6860 71.0370 ;
        RECT 7.5520 69.9435 7.5780 71.0370 ;
        RECT 7.4440 69.9435 7.4700 71.0370 ;
        RECT 7.3360 69.9435 7.3620 71.0370 ;
        RECT 7.2280 69.9435 7.2540 71.0370 ;
        RECT 7.1200 69.9435 7.1460 71.0370 ;
        RECT 7.0120 69.9435 7.0380 71.0370 ;
        RECT 6.9040 69.9435 6.9300 71.0370 ;
        RECT 6.7960 69.9435 6.8220 71.0370 ;
        RECT 6.6880 69.9435 6.7140 71.0370 ;
        RECT 6.5800 69.9435 6.6060 71.0370 ;
        RECT 6.4720 69.9435 6.4980 71.0370 ;
        RECT 6.3640 69.9435 6.3900 71.0370 ;
        RECT 6.2560 69.9435 6.2820 71.0370 ;
        RECT 6.1480 69.9435 6.1740 71.0370 ;
        RECT 6.0400 69.9435 6.0660 71.0370 ;
        RECT 5.9320 69.9435 5.9580 71.0370 ;
        RECT 5.8240 69.9435 5.8500 71.0370 ;
        RECT 5.7160 69.9435 5.7420 71.0370 ;
        RECT 5.6080 69.9435 5.6340 71.0370 ;
        RECT 5.5000 69.9435 5.5260 71.0370 ;
        RECT 5.3920 69.9435 5.4180 71.0370 ;
        RECT 5.2840 69.9435 5.3100 71.0370 ;
        RECT 5.1760 69.9435 5.2020 71.0370 ;
        RECT 5.0680 69.9435 5.0940 71.0370 ;
        RECT 4.9600 69.9435 4.9860 71.0370 ;
        RECT 4.8520 69.9435 4.8780 71.0370 ;
        RECT 4.7440 69.9435 4.7700 71.0370 ;
        RECT 4.6360 69.9435 4.6620 71.0370 ;
        RECT 4.5280 69.9435 4.5540 71.0370 ;
        RECT 4.4200 69.9435 4.4460 71.0370 ;
        RECT 4.3120 69.9435 4.3380 71.0370 ;
        RECT 4.2040 69.9435 4.2300 71.0370 ;
        RECT 4.0960 69.9435 4.1220 71.0370 ;
        RECT 3.9880 69.9435 4.0140 71.0370 ;
        RECT 3.8800 69.9435 3.9060 71.0370 ;
        RECT 3.7720 69.9435 3.7980 71.0370 ;
        RECT 3.6640 69.9435 3.6900 71.0370 ;
        RECT 3.5560 69.9435 3.5820 71.0370 ;
        RECT 3.4480 69.9435 3.4740 71.0370 ;
        RECT 3.3400 69.9435 3.3660 71.0370 ;
        RECT 3.2320 69.9435 3.2580 71.0370 ;
        RECT 3.1240 69.9435 3.1500 71.0370 ;
        RECT 3.0160 69.9435 3.0420 71.0370 ;
        RECT 2.9080 69.9435 2.9340 71.0370 ;
        RECT 2.8000 69.9435 2.8260 71.0370 ;
        RECT 2.6920 69.9435 2.7180 71.0370 ;
        RECT 2.5840 69.9435 2.6100 71.0370 ;
        RECT 2.4760 69.9435 2.5020 71.0370 ;
        RECT 2.3680 69.9435 2.3940 71.0370 ;
        RECT 2.2600 69.9435 2.2860 71.0370 ;
        RECT 2.1520 69.9435 2.1780 71.0370 ;
        RECT 2.0440 69.9435 2.0700 71.0370 ;
        RECT 1.9360 69.9435 1.9620 71.0370 ;
        RECT 1.8280 69.9435 1.8540 71.0370 ;
        RECT 1.7200 69.9435 1.7460 71.0370 ;
        RECT 1.6120 69.9435 1.6380 71.0370 ;
        RECT 1.5040 69.9435 1.5300 71.0370 ;
        RECT 1.3960 69.9435 1.4220 71.0370 ;
        RECT 1.2880 69.9435 1.3140 71.0370 ;
        RECT 1.1800 69.9435 1.2060 71.0370 ;
        RECT 1.0720 69.9435 1.0980 71.0370 ;
        RECT 0.9640 69.9435 0.9900 71.0370 ;
        RECT 0.8560 69.9435 0.8820 71.0370 ;
        RECT 0.7480 69.9435 0.7740 71.0370 ;
        RECT 0.6400 69.9435 0.6660 71.0370 ;
        RECT 0.5320 69.9435 0.5580 71.0370 ;
        RECT 0.4240 69.9435 0.4500 71.0370 ;
        RECT 0.3160 69.9435 0.3420 71.0370 ;
        RECT 0.2080 69.9435 0.2340 71.0370 ;
        RECT 0.0050 69.9435 0.0900 71.0370 ;
        RECT 15.5530 71.0235 15.6810 72.1170 ;
        RECT 15.5390 71.6890 15.6810 72.0115 ;
        RECT 15.3190 71.4160 15.4530 72.1170 ;
        RECT 15.2960 71.7510 15.4530 72.0090 ;
        RECT 15.3190 71.0235 15.4170 72.1170 ;
        RECT 15.3190 71.1445 15.4310 71.3840 ;
        RECT 15.3190 71.0235 15.4530 71.1125 ;
        RECT 15.0940 71.4740 15.2280 72.1170 ;
        RECT 15.0940 71.0235 15.1920 72.1170 ;
        RECT 14.6770 71.0235 14.7600 72.1170 ;
        RECT 14.6770 71.1120 14.7740 72.0475 ;
        RECT 30.2680 71.0235 30.3530 72.1170 ;
        RECT 30.1240 71.0235 30.1500 72.1170 ;
        RECT 30.0160 71.0235 30.0420 72.1170 ;
        RECT 29.9080 71.0235 29.9340 72.1170 ;
        RECT 29.8000 71.0235 29.8260 72.1170 ;
        RECT 29.6920 71.0235 29.7180 72.1170 ;
        RECT 29.5840 71.0235 29.6100 72.1170 ;
        RECT 29.4760 71.0235 29.5020 72.1170 ;
        RECT 29.3680 71.0235 29.3940 72.1170 ;
        RECT 29.2600 71.0235 29.2860 72.1170 ;
        RECT 29.1520 71.0235 29.1780 72.1170 ;
        RECT 29.0440 71.0235 29.0700 72.1170 ;
        RECT 28.9360 71.0235 28.9620 72.1170 ;
        RECT 28.8280 71.0235 28.8540 72.1170 ;
        RECT 28.7200 71.0235 28.7460 72.1170 ;
        RECT 28.6120 71.0235 28.6380 72.1170 ;
        RECT 28.5040 71.0235 28.5300 72.1170 ;
        RECT 28.3960 71.0235 28.4220 72.1170 ;
        RECT 28.2880 71.0235 28.3140 72.1170 ;
        RECT 28.1800 71.0235 28.2060 72.1170 ;
        RECT 28.0720 71.0235 28.0980 72.1170 ;
        RECT 27.9640 71.0235 27.9900 72.1170 ;
        RECT 27.8560 71.0235 27.8820 72.1170 ;
        RECT 27.7480 71.0235 27.7740 72.1170 ;
        RECT 27.6400 71.0235 27.6660 72.1170 ;
        RECT 27.5320 71.0235 27.5580 72.1170 ;
        RECT 27.4240 71.0235 27.4500 72.1170 ;
        RECT 27.3160 71.0235 27.3420 72.1170 ;
        RECT 27.2080 71.0235 27.2340 72.1170 ;
        RECT 27.1000 71.0235 27.1260 72.1170 ;
        RECT 26.9920 71.0235 27.0180 72.1170 ;
        RECT 26.8840 71.0235 26.9100 72.1170 ;
        RECT 26.7760 71.0235 26.8020 72.1170 ;
        RECT 26.6680 71.0235 26.6940 72.1170 ;
        RECT 26.5600 71.0235 26.5860 72.1170 ;
        RECT 26.4520 71.0235 26.4780 72.1170 ;
        RECT 26.3440 71.0235 26.3700 72.1170 ;
        RECT 26.2360 71.0235 26.2620 72.1170 ;
        RECT 26.1280 71.0235 26.1540 72.1170 ;
        RECT 26.0200 71.0235 26.0460 72.1170 ;
        RECT 25.9120 71.0235 25.9380 72.1170 ;
        RECT 25.8040 71.0235 25.8300 72.1170 ;
        RECT 25.6960 71.0235 25.7220 72.1170 ;
        RECT 25.5880 71.0235 25.6140 72.1170 ;
        RECT 25.4800 71.0235 25.5060 72.1170 ;
        RECT 25.3720 71.0235 25.3980 72.1170 ;
        RECT 25.2640 71.0235 25.2900 72.1170 ;
        RECT 25.1560 71.0235 25.1820 72.1170 ;
        RECT 25.0480 71.0235 25.0740 72.1170 ;
        RECT 24.9400 71.0235 24.9660 72.1170 ;
        RECT 24.8320 71.0235 24.8580 72.1170 ;
        RECT 24.7240 71.0235 24.7500 72.1170 ;
        RECT 24.6160 71.0235 24.6420 72.1170 ;
        RECT 24.5080 71.0235 24.5340 72.1170 ;
        RECT 24.4000 71.0235 24.4260 72.1170 ;
        RECT 24.2920 71.0235 24.3180 72.1170 ;
        RECT 24.1840 71.0235 24.2100 72.1170 ;
        RECT 24.0760 71.0235 24.1020 72.1170 ;
        RECT 23.9680 71.0235 23.9940 72.1170 ;
        RECT 23.8600 71.0235 23.8860 72.1170 ;
        RECT 23.7520 71.0235 23.7780 72.1170 ;
        RECT 23.6440 71.0235 23.6700 72.1170 ;
        RECT 23.5360 71.0235 23.5620 72.1170 ;
        RECT 23.4280 71.0235 23.4540 72.1170 ;
        RECT 23.3200 71.0235 23.3460 72.1170 ;
        RECT 23.2120 71.0235 23.2380 72.1170 ;
        RECT 23.1040 71.0235 23.1300 72.1170 ;
        RECT 22.9960 71.0235 23.0220 72.1170 ;
        RECT 22.8880 71.0235 22.9140 72.1170 ;
        RECT 22.7800 71.0235 22.8060 72.1170 ;
        RECT 22.6720 71.0235 22.6980 72.1170 ;
        RECT 22.5640 71.0235 22.5900 72.1170 ;
        RECT 22.4560 71.0235 22.4820 72.1170 ;
        RECT 22.3480 71.0235 22.3740 72.1170 ;
        RECT 22.2400 71.0235 22.2660 72.1170 ;
        RECT 22.1320 71.0235 22.1580 72.1170 ;
        RECT 22.0240 71.0235 22.0500 72.1170 ;
        RECT 21.9160 71.0235 21.9420 72.1170 ;
        RECT 21.8080 71.0235 21.8340 72.1170 ;
        RECT 21.7000 71.0235 21.7260 72.1170 ;
        RECT 21.5920 71.0235 21.6180 72.1170 ;
        RECT 21.4840 71.0235 21.5100 72.1170 ;
        RECT 21.3760 71.0235 21.4020 72.1170 ;
        RECT 21.2680 71.0235 21.2940 72.1170 ;
        RECT 21.1600 71.0235 21.1860 72.1170 ;
        RECT 21.0520 71.0235 21.0780 72.1170 ;
        RECT 20.9440 71.0235 20.9700 72.1170 ;
        RECT 20.8360 71.0235 20.8620 72.1170 ;
        RECT 20.7280 71.0235 20.7540 72.1170 ;
        RECT 20.6200 71.0235 20.6460 72.1170 ;
        RECT 20.5120 71.0235 20.5380 72.1170 ;
        RECT 20.4040 71.0235 20.4300 72.1170 ;
        RECT 20.2960 71.0235 20.3220 72.1170 ;
        RECT 20.1880 71.0235 20.2140 72.1170 ;
        RECT 20.0800 71.0235 20.1060 72.1170 ;
        RECT 19.9720 71.0235 19.9980 72.1170 ;
        RECT 19.8640 71.0235 19.8900 72.1170 ;
        RECT 19.7560 71.0235 19.7820 72.1170 ;
        RECT 19.6480 71.0235 19.6740 72.1170 ;
        RECT 19.5400 71.0235 19.5660 72.1170 ;
        RECT 19.4320 71.0235 19.4580 72.1170 ;
        RECT 19.3240 71.0235 19.3500 72.1170 ;
        RECT 19.2160 71.0235 19.2420 72.1170 ;
        RECT 19.1080 71.0235 19.1340 72.1170 ;
        RECT 19.0000 71.0235 19.0260 72.1170 ;
        RECT 18.8920 71.0235 18.9180 72.1170 ;
        RECT 18.7840 71.0235 18.8100 72.1170 ;
        RECT 18.6760 71.0235 18.7020 72.1170 ;
        RECT 18.5680 71.0235 18.5940 72.1170 ;
        RECT 18.4600 71.0235 18.4860 72.1170 ;
        RECT 18.3520 71.0235 18.3780 72.1170 ;
        RECT 18.2440 71.0235 18.2700 72.1170 ;
        RECT 18.1360 71.0235 18.1620 72.1170 ;
        RECT 18.0280 71.0235 18.0540 72.1170 ;
        RECT 17.9200 71.0235 17.9460 72.1170 ;
        RECT 17.8120 71.0235 17.8380 72.1170 ;
        RECT 17.7040 71.0235 17.7300 72.1170 ;
        RECT 17.5960 71.0235 17.6220 72.1170 ;
        RECT 17.4880 71.0235 17.5140 72.1170 ;
        RECT 17.3800 71.0235 17.4060 72.1170 ;
        RECT 17.2720 71.0235 17.2980 72.1170 ;
        RECT 17.1640 71.0235 17.1900 72.1170 ;
        RECT 17.0560 71.0235 17.0820 72.1170 ;
        RECT 16.9480 71.0235 16.9740 72.1170 ;
        RECT 16.8400 71.0235 16.8660 72.1170 ;
        RECT 16.7320 71.0235 16.7580 72.1170 ;
        RECT 16.6240 71.0235 16.6500 72.1170 ;
        RECT 16.5160 71.0235 16.5420 72.1170 ;
        RECT 16.4080 71.0235 16.4340 72.1170 ;
        RECT 16.3000 71.0235 16.3260 72.1170 ;
        RECT 16.0870 71.0235 16.1640 72.1170 ;
        RECT 14.1940 71.0235 14.2710 72.1170 ;
        RECT 14.0320 71.0235 14.0580 72.1170 ;
        RECT 13.9240 71.0235 13.9500 72.1170 ;
        RECT 13.8160 71.0235 13.8420 72.1170 ;
        RECT 13.7080 71.0235 13.7340 72.1170 ;
        RECT 13.6000 71.0235 13.6260 72.1170 ;
        RECT 13.4920 71.0235 13.5180 72.1170 ;
        RECT 13.3840 71.0235 13.4100 72.1170 ;
        RECT 13.2760 71.0235 13.3020 72.1170 ;
        RECT 13.1680 71.0235 13.1940 72.1170 ;
        RECT 13.0600 71.0235 13.0860 72.1170 ;
        RECT 12.9520 71.0235 12.9780 72.1170 ;
        RECT 12.8440 71.0235 12.8700 72.1170 ;
        RECT 12.7360 71.0235 12.7620 72.1170 ;
        RECT 12.6280 71.0235 12.6540 72.1170 ;
        RECT 12.5200 71.0235 12.5460 72.1170 ;
        RECT 12.4120 71.0235 12.4380 72.1170 ;
        RECT 12.3040 71.0235 12.3300 72.1170 ;
        RECT 12.1960 71.0235 12.2220 72.1170 ;
        RECT 12.0880 71.0235 12.1140 72.1170 ;
        RECT 11.9800 71.0235 12.0060 72.1170 ;
        RECT 11.8720 71.0235 11.8980 72.1170 ;
        RECT 11.7640 71.0235 11.7900 72.1170 ;
        RECT 11.6560 71.0235 11.6820 72.1170 ;
        RECT 11.5480 71.0235 11.5740 72.1170 ;
        RECT 11.4400 71.0235 11.4660 72.1170 ;
        RECT 11.3320 71.0235 11.3580 72.1170 ;
        RECT 11.2240 71.0235 11.2500 72.1170 ;
        RECT 11.1160 71.0235 11.1420 72.1170 ;
        RECT 11.0080 71.0235 11.0340 72.1170 ;
        RECT 10.9000 71.0235 10.9260 72.1170 ;
        RECT 10.7920 71.0235 10.8180 72.1170 ;
        RECT 10.6840 71.0235 10.7100 72.1170 ;
        RECT 10.5760 71.0235 10.6020 72.1170 ;
        RECT 10.4680 71.0235 10.4940 72.1170 ;
        RECT 10.3600 71.0235 10.3860 72.1170 ;
        RECT 10.2520 71.0235 10.2780 72.1170 ;
        RECT 10.1440 71.0235 10.1700 72.1170 ;
        RECT 10.0360 71.0235 10.0620 72.1170 ;
        RECT 9.9280 71.0235 9.9540 72.1170 ;
        RECT 9.8200 71.0235 9.8460 72.1170 ;
        RECT 9.7120 71.0235 9.7380 72.1170 ;
        RECT 9.6040 71.0235 9.6300 72.1170 ;
        RECT 9.4960 71.0235 9.5220 72.1170 ;
        RECT 9.3880 71.0235 9.4140 72.1170 ;
        RECT 9.2800 71.0235 9.3060 72.1170 ;
        RECT 9.1720 71.0235 9.1980 72.1170 ;
        RECT 9.0640 71.0235 9.0900 72.1170 ;
        RECT 8.9560 71.0235 8.9820 72.1170 ;
        RECT 8.8480 71.0235 8.8740 72.1170 ;
        RECT 8.7400 71.0235 8.7660 72.1170 ;
        RECT 8.6320 71.0235 8.6580 72.1170 ;
        RECT 8.5240 71.0235 8.5500 72.1170 ;
        RECT 8.4160 71.0235 8.4420 72.1170 ;
        RECT 8.3080 71.0235 8.3340 72.1170 ;
        RECT 8.2000 71.0235 8.2260 72.1170 ;
        RECT 8.0920 71.0235 8.1180 72.1170 ;
        RECT 7.9840 71.0235 8.0100 72.1170 ;
        RECT 7.8760 71.0235 7.9020 72.1170 ;
        RECT 7.7680 71.0235 7.7940 72.1170 ;
        RECT 7.6600 71.0235 7.6860 72.1170 ;
        RECT 7.5520 71.0235 7.5780 72.1170 ;
        RECT 7.4440 71.0235 7.4700 72.1170 ;
        RECT 7.3360 71.0235 7.3620 72.1170 ;
        RECT 7.2280 71.0235 7.2540 72.1170 ;
        RECT 7.1200 71.0235 7.1460 72.1170 ;
        RECT 7.0120 71.0235 7.0380 72.1170 ;
        RECT 6.9040 71.0235 6.9300 72.1170 ;
        RECT 6.7960 71.0235 6.8220 72.1170 ;
        RECT 6.6880 71.0235 6.7140 72.1170 ;
        RECT 6.5800 71.0235 6.6060 72.1170 ;
        RECT 6.4720 71.0235 6.4980 72.1170 ;
        RECT 6.3640 71.0235 6.3900 72.1170 ;
        RECT 6.2560 71.0235 6.2820 72.1170 ;
        RECT 6.1480 71.0235 6.1740 72.1170 ;
        RECT 6.0400 71.0235 6.0660 72.1170 ;
        RECT 5.9320 71.0235 5.9580 72.1170 ;
        RECT 5.8240 71.0235 5.8500 72.1170 ;
        RECT 5.7160 71.0235 5.7420 72.1170 ;
        RECT 5.6080 71.0235 5.6340 72.1170 ;
        RECT 5.5000 71.0235 5.5260 72.1170 ;
        RECT 5.3920 71.0235 5.4180 72.1170 ;
        RECT 5.2840 71.0235 5.3100 72.1170 ;
        RECT 5.1760 71.0235 5.2020 72.1170 ;
        RECT 5.0680 71.0235 5.0940 72.1170 ;
        RECT 4.9600 71.0235 4.9860 72.1170 ;
        RECT 4.8520 71.0235 4.8780 72.1170 ;
        RECT 4.7440 71.0235 4.7700 72.1170 ;
        RECT 4.6360 71.0235 4.6620 72.1170 ;
        RECT 4.5280 71.0235 4.5540 72.1170 ;
        RECT 4.4200 71.0235 4.4460 72.1170 ;
        RECT 4.3120 71.0235 4.3380 72.1170 ;
        RECT 4.2040 71.0235 4.2300 72.1170 ;
        RECT 4.0960 71.0235 4.1220 72.1170 ;
        RECT 3.9880 71.0235 4.0140 72.1170 ;
        RECT 3.8800 71.0235 3.9060 72.1170 ;
        RECT 3.7720 71.0235 3.7980 72.1170 ;
        RECT 3.6640 71.0235 3.6900 72.1170 ;
        RECT 3.5560 71.0235 3.5820 72.1170 ;
        RECT 3.4480 71.0235 3.4740 72.1170 ;
        RECT 3.3400 71.0235 3.3660 72.1170 ;
        RECT 3.2320 71.0235 3.2580 72.1170 ;
        RECT 3.1240 71.0235 3.1500 72.1170 ;
        RECT 3.0160 71.0235 3.0420 72.1170 ;
        RECT 2.9080 71.0235 2.9340 72.1170 ;
        RECT 2.8000 71.0235 2.8260 72.1170 ;
        RECT 2.6920 71.0235 2.7180 72.1170 ;
        RECT 2.5840 71.0235 2.6100 72.1170 ;
        RECT 2.4760 71.0235 2.5020 72.1170 ;
        RECT 2.3680 71.0235 2.3940 72.1170 ;
        RECT 2.2600 71.0235 2.2860 72.1170 ;
        RECT 2.1520 71.0235 2.1780 72.1170 ;
        RECT 2.0440 71.0235 2.0700 72.1170 ;
        RECT 1.9360 71.0235 1.9620 72.1170 ;
        RECT 1.8280 71.0235 1.8540 72.1170 ;
        RECT 1.7200 71.0235 1.7460 72.1170 ;
        RECT 1.6120 71.0235 1.6380 72.1170 ;
        RECT 1.5040 71.0235 1.5300 72.1170 ;
        RECT 1.3960 71.0235 1.4220 72.1170 ;
        RECT 1.2880 71.0235 1.3140 72.1170 ;
        RECT 1.1800 71.0235 1.2060 72.1170 ;
        RECT 1.0720 71.0235 1.0980 72.1170 ;
        RECT 0.9640 71.0235 0.9900 72.1170 ;
        RECT 0.8560 71.0235 0.8820 72.1170 ;
        RECT 0.7480 71.0235 0.7740 72.1170 ;
        RECT 0.6400 71.0235 0.6660 72.1170 ;
        RECT 0.5320 71.0235 0.5580 72.1170 ;
        RECT 0.4240 71.0235 0.4500 72.1170 ;
        RECT 0.3160 71.0235 0.3420 72.1170 ;
        RECT 0.2080 71.0235 0.2340 72.1170 ;
        RECT 0.0050 71.0235 0.0900 72.1170 ;
        RECT 15.5530 72.1035 15.6810 73.1970 ;
        RECT 15.5390 72.7690 15.6810 73.0915 ;
        RECT 15.3190 72.4960 15.4530 73.1970 ;
        RECT 15.2960 72.8310 15.4530 73.0890 ;
        RECT 15.3190 72.1035 15.4170 73.1970 ;
        RECT 15.3190 72.2245 15.4310 72.4640 ;
        RECT 15.3190 72.1035 15.4530 72.1925 ;
        RECT 15.0940 72.5540 15.2280 73.1970 ;
        RECT 15.0940 72.1035 15.1920 73.1970 ;
        RECT 14.6770 72.1035 14.7600 73.1970 ;
        RECT 14.6770 72.1920 14.7740 73.1275 ;
        RECT 30.2680 72.1035 30.3530 73.1970 ;
        RECT 30.1240 72.1035 30.1500 73.1970 ;
        RECT 30.0160 72.1035 30.0420 73.1970 ;
        RECT 29.9080 72.1035 29.9340 73.1970 ;
        RECT 29.8000 72.1035 29.8260 73.1970 ;
        RECT 29.6920 72.1035 29.7180 73.1970 ;
        RECT 29.5840 72.1035 29.6100 73.1970 ;
        RECT 29.4760 72.1035 29.5020 73.1970 ;
        RECT 29.3680 72.1035 29.3940 73.1970 ;
        RECT 29.2600 72.1035 29.2860 73.1970 ;
        RECT 29.1520 72.1035 29.1780 73.1970 ;
        RECT 29.0440 72.1035 29.0700 73.1970 ;
        RECT 28.9360 72.1035 28.9620 73.1970 ;
        RECT 28.8280 72.1035 28.8540 73.1970 ;
        RECT 28.7200 72.1035 28.7460 73.1970 ;
        RECT 28.6120 72.1035 28.6380 73.1970 ;
        RECT 28.5040 72.1035 28.5300 73.1970 ;
        RECT 28.3960 72.1035 28.4220 73.1970 ;
        RECT 28.2880 72.1035 28.3140 73.1970 ;
        RECT 28.1800 72.1035 28.2060 73.1970 ;
        RECT 28.0720 72.1035 28.0980 73.1970 ;
        RECT 27.9640 72.1035 27.9900 73.1970 ;
        RECT 27.8560 72.1035 27.8820 73.1970 ;
        RECT 27.7480 72.1035 27.7740 73.1970 ;
        RECT 27.6400 72.1035 27.6660 73.1970 ;
        RECT 27.5320 72.1035 27.5580 73.1970 ;
        RECT 27.4240 72.1035 27.4500 73.1970 ;
        RECT 27.3160 72.1035 27.3420 73.1970 ;
        RECT 27.2080 72.1035 27.2340 73.1970 ;
        RECT 27.1000 72.1035 27.1260 73.1970 ;
        RECT 26.9920 72.1035 27.0180 73.1970 ;
        RECT 26.8840 72.1035 26.9100 73.1970 ;
        RECT 26.7760 72.1035 26.8020 73.1970 ;
        RECT 26.6680 72.1035 26.6940 73.1970 ;
        RECT 26.5600 72.1035 26.5860 73.1970 ;
        RECT 26.4520 72.1035 26.4780 73.1970 ;
        RECT 26.3440 72.1035 26.3700 73.1970 ;
        RECT 26.2360 72.1035 26.2620 73.1970 ;
        RECT 26.1280 72.1035 26.1540 73.1970 ;
        RECT 26.0200 72.1035 26.0460 73.1970 ;
        RECT 25.9120 72.1035 25.9380 73.1970 ;
        RECT 25.8040 72.1035 25.8300 73.1970 ;
        RECT 25.6960 72.1035 25.7220 73.1970 ;
        RECT 25.5880 72.1035 25.6140 73.1970 ;
        RECT 25.4800 72.1035 25.5060 73.1970 ;
        RECT 25.3720 72.1035 25.3980 73.1970 ;
        RECT 25.2640 72.1035 25.2900 73.1970 ;
        RECT 25.1560 72.1035 25.1820 73.1970 ;
        RECT 25.0480 72.1035 25.0740 73.1970 ;
        RECT 24.9400 72.1035 24.9660 73.1970 ;
        RECT 24.8320 72.1035 24.8580 73.1970 ;
        RECT 24.7240 72.1035 24.7500 73.1970 ;
        RECT 24.6160 72.1035 24.6420 73.1970 ;
        RECT 24.5080 72.1035 24.5340 73.1970 ;
        RECT 24.4000 72.1035 24.4260 73.1970 ;
        RECT 24.2920 72.1035 24.3180 73.1970 ;
        RECT 24.1840 72.1035 24.2100 73.1970 ;
        RECT 24.0760 72.1035 24.1020 73.1970 ;
        RECT 23.9680 72.1035 23.9940 73.1970 ;
        RECT 23.8600 72.1035 23.8860 73.1970 ;
        RECT 23.7520 72.1035 23.7780 73.1970 ;
        RECT 23.6440 72.1035 23.6700 73.1970 ;
        RECT 23.5360 72.1035 23.5620 73.1970 ;
        RECT 23.4280 72.1035 23.4540 73.1970 ;
        RECT 23.3200 72.1035 23.3460 73.1970 ;
        RECT 23.2120 72.1035 23.2380 73.1970 ;
        RECT 23.1040 72.1035 23.1300 73.1970 ;
        RECT 22.9960 72.1035 23.0220 73.1970 ;
        RECT 22.8880 72.1035 22.9140 73.1970 ;
        RECT 22.7800 72.1035 22.8060 73.1970 ;
        RECT 22.6720 72.1035 22.6980 73.1970 ;
        RECT 22.5640 72.1035 22.5900 73.1970 ;
        RECT 22.4560 72.1035 22.4820 73.1970 ;
        RECT 22.3480 72.1035 22.3740 73.1970 ;
        RECT 22.2400 72.1035 22.2660 73.1970 ;
        RECT 22.1320 72.1035 22.1580 73.1970 ;
        RECT 22.0240 72.1035 22.0500 73.1970 ;
        RECT 21.9160 72.1035 21.9420 73.1970 ;
        RECT 21.8080 72.1035 21.8340 73.1970 ;
        RECT 21.7000 72.1035 21.7260 73.1970 ;
        RECT 21.5920 72.1035 21.6180 73.1970 ;
        RECT 21.4840 72.1035 21.5100 73.1970 ;
        RECT 21.3760 72.1035 21.4020 73.1970 ;
        RECT 21.2680 72.1035 21.2940 73.1970 ;
        RECT 21.1600 72.1035 21.1860 73.1970 ;
        RECT 21.0520 72.1035 21.0780 73.1970 ;
        RECT 20.9440 72.1035 20.9700 73.1970 ;
        RECT 20.8360 72.1035 20.8620 73.1970 ;
        RECT 20.7280 72.1035 20.7540 73.1970 ;
        RECT 20.6200 72.1035 20.6460 73.1970 ;
        RECT 20.5120 72.1035 20.5380 73.1970 ;
        RECT 20.4040 72.1035 20.4300 73.1970 ;
        RECT 20.2960 72.1035 20.3220 73.1970 ;
        RECT 20.1880 72.1035 20.2140 73.1970 ;
        RECT 20.0800 72.1035 20.1060 73.1970 ;
        RECT 19.9720 72.1035 19.9980 73.1970 ;
        RECT 19.8640 72.1035 19.8900 73.1970 ;
        RECT 19.7560 72.1035 19.7820 73.1970 ;
        RECT 19.6480 72.1035 19.6740 73.1970 ;
        RECT 19.5400 72.1035 19.5660 73.1970 ;
        RECT 19.4320 72.1035 19.4580 73.1970 ;
        RECT 19.3240 72.1035 19.3500 73.1970 ;
        RECT 19.2160 72.1035 19.2420 73.1970 ;
        RECT 19.1080 72.1035 19.1340 73.1970 ;
        RECT 19.0000 72.1035 19.0260 73.1970 ;
        RECT 18.8920 72.1035 18.9180 73.1970 ;
        RECT 18.7840 72.1035 18.8100 73.1970 ;
        RECT 18.6760 72.1035 18.7020 73.1970 ;
        RECT 18.5680 72.1035 18.5940 73.1970 ;
        RECT 18.4600 72.1035 18.4860 73.1970 ;
        RECT 18.3520 72.1035 18.3780 73.1970 ;
        RECT 18.2440 72.1035 18.2700 73.1970 ;
        RECT 18.1360 72.1035 18.1620 73.1970 ;
        RECT 18.0280 72.1035 18.0540 73.1970 ;
        RECT 17.9200 72.1035 17.9460 73.1970 ;
        RECT 17.8120 72.1035 17.8380 73.1970 ;
        RECT 17.7040 72.1035 17.7300 73.1970 ;
        RECT 17.5960 72.1035 17.6220 73.1970 ;
        RECT 17.4880 72.1035 17.5140 73.1970 ;
        RECT 17.3800 72.1035 17.4060 73.1970 ;
        RECT 17.2720 72.1035 17.2980 73.1970 ;
        RECT 17.1640 72.1035 17.1900 73.1970 ;
        RECT 17.0560 72.1035 17.0820 73.1970 ;
        RECT 16.9480 72.1035 16.9740 73.1970 ;
        RECT 16.8400 72.1035 16.8660 73.1970 ;
        RECT 16.7320 72.1035 16.7580 73.1970 ;
        RECT 16.6240 72.1035 16.6500 73.1970 ;
        RECT 16.5160 72.1035 16.5420 73.1970 ;
        RECT 16.4080 72.1035 16.4340 73.1970 ;
        RECT 16.3000 72.1035 16.3260 73.1970 ;
        RECT 16.0870 72.1035 16.1640 73.1970 ;
        RECT 14.1940 72.1035 14.2710 73.1970 ;
        RECT 14.0320 72.1035 14.0580 73.1970 ;
        RECT 13.9240 72.1035 13.9500 73.1970 ;
        RECT 13.8160 72.1035 13.8420 73.1970 ;
        RECT 13.7080 72.1035 13.7340 73.1970 ;
        RECT 13.6000 72.1035 13.6260 73.1970 ;
        RECT 13.4920 72.1035 13.5180 73.1970 ;
        RECT 13.3840 72.1035 13.4100 73.1970 ;
        RECT 13.2760 72.1035 13.3020 73.1970 ;
        RECT 13.1680 72.1035 13.1940 73.1970 ;
        RECT 13.0600 72.1035 13.0860 73.1970 ;
        RECT 12.9520 72.1035 12.9780 73.1970 ;
        RECT 12.8440 72.1035 12.8700 73.1970 ;
        RECT 12.7360 72.1035 12.7620 73.1970 ;
        RECT 12.6280 72.1035 12.6540 73.1970 ;
        RECT 12.5200 72.1035 12.5460 73.1970 ;
        RECT 12.4120 72.1035 12.4380 73.1970 ;
        RECT 12.3040 72.1035 12.3300 73.1970 ;
        RECT 12.1960 72.1035 12.2220 73.1970 ;
        RECT 12.0880 72.1035 12.1140 73.1970 ;
        RECT 11.9800 72.1035 12.0060 73.1970 ;
        RECT 11.8720 72.1035 11.8980 73.1970 ;
        RECT 11.7640 72.1035 11.7900 73.1970 ;
        RECT 11.6560 72.1035 11.6820 73.1970 ;
        RECT 11.5480 72.1035 11.5740 73.1970 ;
        RECT 11.4400 72.1035 11.4660 73.1970 ;
        RECT 11.3320 72.1035 11.3580 73.1970 ;
        RECT 11.2240 72.1035 11.2500 73.1970 ;
        RECT 11.1160 72.1035 11.1420 73.1970 ;
        RECT 11.0080 72.1035 11.0340 73.1970 ;
        RECT 10.9000 72.1035 10.9260 73.1970 ;
        RECT 10.7920 72.1035 10.8180 73.1970 ;
        RECT 10.6840 72.1035 10.7100 73.1970 ;
        RECT 10.5760 72.1035 10.6020 73.1970 ;
        RECT 10.4680 72.1035 10.4940 73.1970 ;
        RECT 10.3600 72.1035 10.3860 73.1970 ;
        RECT 10.2520 72.1035 10.2780 73.1970 ;
        RECT 10.1440 72.1035 10.1700 73.1970 ;
        RECT 10.0360 72.1035 10.0620 73.1970 ;
        RECT 9.9280 72.1035 9.9540 73.1970 ;
        RECT 9.8200 72.1035 9.8460 73.1970 ;
        RECT 9.7120 72.1035 9.7380 73.1970 ;
        RECT 9.6040 72.1035 9.6300 73.1970 ;
        RECT 9.4960 72.1035 9.5220 73.1970 ;
        RECT 9.3880 72.1035 9.4140 73.1970 ;
        RECT 9.2800 72.1035 9.3060 73.1970 ;
        RECT 9.1720 72.1035 9.1980 73.1970 ;
        RECT 9.0640 72.1035 9.0900 73.1970 ;
        RECT 8.9560 72.1035 8.9820 73.1970 ;
        RECT 8.8480 72.1035 8.8740 73.1970 ;
        RECT 8.7400 72.1035 8.7660 73.1970 ;
        RECT 8.6320 72.1035 8.6580 73.1970 ;
        RECT 8.5240 72.1035 8.5500 73.1970 ;
        RECT 8.4160 72.1035 8.4420 73.1970 ;
        RECT 8.3080 72.1035 8.3340 73.1970 ;
        RECT 8.2000 72.1035 8.2260 73.1970 ;
        RECT 8.0920 72.1035 8.1180 73.1970 ;
        RECT 7.9840 72.1035 8.0100 73.1970 ;
        RECT 7.8760 72.1035 7.9020 73.1970 ;
        RECT 7.7680 72.1035 7.7940 73.1970 ;
        RECT 7.6600 72.1035 7.6860 73.1970 ;
        RECT 7.5520 72.1035 7.5780 73.1970 ;
        RECT 7.4440 72.1035 7.4700 73.1970 ;
        RECT 7.3360 72.1035 7.3620 73.1970 ;
        RECT 7.2280 72.1035 7.2540 73.1970 ;
        RECT 7.1200 72.1035 7.1460 73.1970 ;
        RECT 7.0120 72.1035 7.0380 73.1970 ;
        RECT 6.9040 72.1035 6.9300 73.1970 ;
        RECT 6.7960 72.1035 6.8220 73.1970 ;
        RECT 6.6880 72.1035 6.7140 73.1970 ;
        RECT 6.5800 72.1035 6.6060 73.1970 ;
        RECT 6.4720 72.1035 6.4980 73.1970 ;
        RECT 6.3640 72.1035 6.3900 73.1970 ;
        RECT 6.2560 72.1035 6.2820 73.1970 ;
        RECT 6.1480 72.1035 6.1740 73.1970 ;
        RECT 6.0400 72.1035 6.0660 73.1970 ;
        RECT 5.9320 72.1035 5.9580 73.1970 ;
        RECT 5.8240 72.1035 5.8500 73.1970 ;
        RECT 5.7160 72.1035 5.7420 73.1970 ;
        RECT 5.6080 72.1035 5.6340 73.1970 ;
        RECT 5.5000 72.1035 5.5260 73.1970 ;
        RECT 5.3920 72.1035 5.4180 73.1970 ;
        RECT 5.2840 72.1035 5.3100 73.1970 ;
        RECT 5.1760 72.1035 5.2020 73.1970 ;
        RECT 5.0680 72.1035 5.0940 73.1970 ;
        RECT 4.9600 72.1035 4.9860 73.1970 ;
        RECT 4.8520 72.1035 4.8780 73.1970 ;
        RECT 4.7440 72.1035 4.7700 73.1970 ;
        RECT 4.6360 72.1035 4.6620 73.1970 ;
        RECT 4.5280 72.1035 4.5540 73.1970 ;
        RECT 4.4200 72.1035 4.4460 73.1970 ;
        RECT 4.3120 72.1035 4.3380 73.1970 ;
        RECT 4.2040 72.1035 4.2300 73.1970 ;
        RECT 4.0960 72.1035 4.1220 73.1970 ;
        RECT 3.9880 72.1035 4.0140 73.1970 ;
        RECT 3.8800 72.1035 3.9060 73.1970 ;
        RECT 3.7720 72.1035 3.7980 73.1970 ;
        RECT 3.6640 72.1035 3.6900 73.1970 ;
        RECT 3.5560 72.1035 3.5820 73.1970 ;
        RECT 3.4480 72.1035 3.4740 73.1970 ;
        RECT 3.3400 72.1035 3.3660 73.1970 ;
        RECT 3.2320 72.1035 3.2580 73.1970 ;
        RECT 3.1240 72.1035 3.1500 73.1970 ;
        RECT 3.0160 72.1035 3.0420 73.1970 ;
        RECT 2.9080 72.1035 2.9340 73.1970 ;
        RECT 2.8000 72.1035 2.8260 73.1970 ;
        RECT 2.6920 72.1035 2.7180 73.1970 ;
        RECT 2.5840 72.1035 2.6100 73.1970 ;
        RECT 2.4760 72.1035 2.5020 73.1970 ;
        RECT 2.3680 72.1035 2.3940 73.1970 ;
        RECT 2.2600 72.1035 2.2860 73.1970 ;
        RECT 2.1520 72.1035 2.1780 73.1970 ;
        RECT 2.0440 72.1035 2.0700 73.1970 ;
        RECT 1.9360 72.1035 1.9620 73.1970 ;
        RECT 1.8280 72.1035 1.8540 73.1970 ;
        RECT 1.7200 72.1035 1.7460 73.1970 ;
        RECT 1.6120 72.1035 1.6380 73.1970 ;
        RECT 1.5040 72.1035 1.5300 73.1970 ;
        RECT 1.3960 72.1035 1.4220 73.1970 ;
        RECT 1.2880 72.1035 1.3140 73.1970 ;
        RECT 1.1800 72.1035 1.2060 73.1970 ;
        RECT 1.0720 72.1035 1.0980 73.1970 ;
        RECT 0.9640 72.1035 0.9900 73.1970 ;
        RECT 0.8560 72.1035 0.8820 73.1970 ;
        RECT 0.7480 72.1035 0.7740 73.1970 ;
        RECT 0.6400 72.1035 0.6660 73.1970 ;
        RECT 0.5320 72.1035 0.5580 73.1970 ;
        RECT 0.4240 72.1035 0.4500 73.1970 ;
        RECT 0.3160 72.1035 0.3420 73.1970 ;
        RECT 0.2080 72.1035 0.2340 73.1970 ;
        RECT 0.0050 72.1035 0.0900 73.1970 ;
        RECT 15.5530 73.1835 15.6810 74.2770 ;
        RECT 15.5390 73.8490 15.6810 74.1715 ;
        RECT 15.3190 73.5760 15.4530 74.2770 ;
        RECT 15.2960 73.9110 15.4530 74.1690 ;
        RECT 15.3190 73.1835 15.4170 74.2770 ;
        RECT 15.3190 73.3045 15.4310 73.5440 ;
        RECT 15.3190 73.1835 15.4530 73.2725 ;
        RECT 15.0940 73.6340 15.2280 74.2770 ;
        RECT 15.0940 73.1835 15.1920 74.2770 ;
        RECT 14.6770 73.1835 14.7600 74.2770 ;
        RECT 14.6770 73.2720 14.7740 74.2075 ;
        RECT 30.2680 73.1835 30.3530 74.2770 ;
        RECT 30.1240 73.1835 30.1500 74.2770 ;
        RECT 30.0160 73.1835 30.0420 74.2770 ;
        RECT 29.9080 73.1835 29.9340 74.2770 ;
        RECT 29.8000 73.1835 29.8260 74.2770 ;
        RECT 29.6920 73.1835 29.7180 74.2770 ;
        RECT 29.5840 73.1835 29.6100 74.2770 ;
        RECT 29.4760 73.1835 29.5020 74.2770 ;
        RECT 29.3680 73.1835 29.3940 74.2770 ;
        RECT 29.2600 73.1835 29.2860 74.2770 ;
        RECT 29.1520 73.1835 29.1780 74.2770 ;
        RECT 29.0440 73.1835 29.0700 74.2770 ;
        RECT 28.9360 73.1835 28.9620 74.2770 ;
        RECT 28.8280 73.1835 28.8540 74.2770 ;
        RECT 28.7200 73.1835 28.7460 74.2770 ;
        RECT 28.6120 73.1835 28.6380 74.2770 ;
        RECT 28.5040 73.1835 28.5300 74.2770 ;
        RECT 28.3960 73.1835 28.4220 74.2770 ;
        RECT 28.2880 73.1835 28.3140 74.2770 ;
        RECT 28.1800 73.1835 28.2060 74.2770 ;
        RECT 28.0720 73.1835 28.0980 74.2770 ;
        RECT 27.9640 73.1835 27.9900 74.2770 ;
        RECT 27.8560 73.1835 27.8820 74.2770 ;
        RECT 27.7480 73.1835 27.7740 74.2770 ;
        RECT 27.6400 73.1835 27.6660 74.2770 ;
        RECT 27.5320 73.1835 27.5580 74.2770 ;
        RECT 27.4240 73.1835 27.4500 74.2770 ;
        RECT 27.3160 73.1835 27.3420 74.2770 ;
        RECT 27.2080 73.1835 27.2340 74.2770 ;
        RECT 27.1000 73.1835 27.1260 74.2770 ;
        RECT 26.9920 73.1835 27.0180 74.2770 ;
        RECT 26.8840 73.1835 26.9100 74.2770 ;
        RECT 26.7760 73.1835 26.8020 74.2770 ;
        RECT 26.6680 73.1835 26.6940 74.2770 ;
        RECT 26.5600 73.1835 26.5860 74.2770 ;
        RECT 26.4520 73.1835 26.4780 74.2770 ;
        RECT 26.3440 73.1835 26.3700 74.2770 ;
        RECT 26.2360 73.1835 26.2620 74.2770 ;
        RECT 26.1280 73.1835 26.1540 74.2770 ;
        RECT 26.0200 73.1835 26.0460 74.2770 ;
        RECT 25.9120 73.1835 25.9380 74.2770 ;
        RECT 25.8040 73.1835 25.8300 74.2770 ;
        RECT 25.6960 73.1835 25.7220 74.2770 ;
        RECT 25.5880 73.1835 25.6140 74.2770 ;
        RECT 25.4800 73.1835 25.5060 74.2770 ;
        RECT 25.3720 73.1835 25.3980 74.2770 ;
        RECT 25.2640 73.1835 25.2900 74.2770 ;
        RECT 25.1560 73.1835 25.1820 74.2770 ;
        RECT 25.0480 73.1835 25.0740 74.2770 ;
        RECT 24.9400 73.1835 24.9660 74.2770 ;
        RECT 24.8320 73.1835 24.8580 74.2770 ;
        RECT 24.7240 73.1835 24.7500 74.2770 ;
        RECT 24.6160 73.1835 24.6420 74.2770 ;
        RECT 24.5080 73.1835 24.5340 74.2770 ;
        RECT 24.4000 73.1835 24.4260 74.2770 ;
        RECT 24.2920 73.1835 24.3180 74.2770 ;
        RECT 24.1840 73.1835 24.2100 74.2770 ;
        RECT 24.0760 73.1835 24.1020 74.2770 ;
        RECT 23.9680 73.1835 23.9940 74.2770 ;
        RECT 23.8600 73.1835 23.8860 74.2770 ;
        RECT 23.7520 73.1835 23.7780 74.2770 ;
        RECT 23.6440 73.1835 23.6700 74.2770 ;
        RECT 23.5360 73.1835 23.5620 74.2770 ;
        RECT 23.4280 73.1835 23.4540 74.2770 ;
        RECT 23.3200 73.1835 23.3460 74.2770 ;
        RECT 23.2120 73.1835 23.2380 74.2770 ;
        RECT 23.1040 73.1835 23.1300 74.2770 ;
        RECT 22.9960 73.1835 23.0220 74.2770 ;
        RECT 22.8880 73.1835 22.9140 74.2770 ;
        RECT 22.7800 73.1835 22.8060 74.2770 ;
        RECT 22.6720 73.1835 22.6980 74.2770 ;
        RECT 22.5640 73.1835 22.5900 74.2770 ;
        RECT 22.4560 73.1835 22.4820 74.2770 ;
        RECT 22.3480 73.1835 22.3740 74.2770 ;
        RECT 22.2400 73.1835 22.2660 74.2770 ;
        RECT 22.1320 73.1835 22.1580 74.2770 ;
        RECT 22.0240 73.1835 22.0500 74.2770 ;
        RECT 21.9160 73.1835 21.9420 74.2770 ;
        RECT 21.8080 73.1835 21.8340 74.2770 ;
        RECT 21.7000 73.1835 21.7260 74.2770 ;
        RECT 21.5920 73.1835 21.6180 74.2770 ;
        RECT 21.4840 73.1835 21.5100 74.2770 ;
        RECT 21.3760 73.1835 21.4020 74.2770 ;
        RECT 21.2680 73.1835 21.2940 74.2770 ;
        RECT 21.1600 73.1835 21.1860 74.2770 ;
        RECT 21.0520 73.1835 21.0780 74.2770 ;
        RECT 20.9440 73.1835 20.9700 74.2770 ;
        RECT 20.8360 73.1835 20.8620 74.2770 ;
        RECT 20.7280 73.1835 20.7540 74.2770 ;
        RECT 20.6200 73.1835 20.6460 74.2770 ;
        RECT 20.5120 73.1835 20.5380 74.2770 ;
        RECT 20.4040 73.1835 20.4300 74.2770 ;
        RECT 20.2960 73.1835 20.3220 74.2770 ;
        RECT 20.1880 73.1835 20.2140 74.2770 ;
        RECT 20.0800 73.1835 20.1060 74.2770 ;
        RECT 19.9720 73.1835 19.9980 74.2770 ;
        RECT 19.8640 73.1835 19.8900 74.2770 ;
        RECT 19.7560 73.1835 19.7820 74.2770 ;
        RECT 19.6480 73.1835 19.6740 74.2770 ;
        RECT 19.5400 73.1835 19.5660 74.2770 ;
        RECT 19.4320 73.1835 19.4580 74.2770 ;
        RECT 19.3240 73.1835 19.3500 74.2770 ;
        RECT 19.2160 73.1835 19.2420 74.2770 ;
        RECT 19.1080 73.1835 19.1340 74.2770 ;
        RECT 19.0000 73.1835 19.0260 74.2770 ;
        RECT 18.8920 73.1835 18.9180 74.2770 ;
        RECT 18.7840 73.1835 18.8100 74.2770 ;
        RECT 18.6760 73.1835 18.7020 74.2770 ;
        RECT 18.5680 73.1835 18.5940 74.2770 ;
        RECT 18.4600 73.1835 18.4860 74.2770 ;
        RECT 18.3520 73.1835 18.3780 74.2770 ;
        RECT 18.2440 73.1835 18.2700 74.2770 ;
        RECT 18.1360 73.1835 18.1620 74.2770 ;
        RECT 18.0280 73.1835 18.0540 74.2770 ;
        RECT 17.9200 73.1835 17.9460 74.2770 ;
        RECT 17.8120 73.1835 17.8380 74.2770 ;
        RECT 17.7040 73.1835 17.7300 74.2770 ;
        RECT 17.5960 73.1835 17.6220 74.2770 ;
        RECT 17.4880 73.1835 17.5140 74.2770 ;
        RECT 17.3800 73.1835 17.4060 74.2770 ;
        RECT 17.2720 73.1835 17.2980 74.2770 ;
        RECT 17.1640 73.1835 17.1900 74.2770 ;
        RECT 17.0560 73.1835 17.0820 74.2770 ;
        RECT 16.9480 73.1835 16.9740 74.2770 ;
        RECT 16.8400 73.1835 16.8660 74.2770 ;
        RECT 16.7320 73.1835 16.7580 74.2770 ;
        RECT 16.6240 73.1835 16.6500 74.2770 ;
        RECT 16.5160 73.1835 16.5420 74.2770 ;
        RECT 16.4080 73.1835 16.4340 74.2770 ;
        RECT 16.3000 73.1835 16.3260 74.2770 ;
        RECT 16.0870 73.1835 16.1640 74.2770 ;
        RECT 14.1940 73.1835 14.2710 74.2770 ;
        RECT 14.0320 73.1835 14.0580 74.2770 ;
        RECT 13.9240 73.1835 13.9500 74.2770 ;
        RECT 13.8160 73.1835 13.8420 74.2770 ;
        RECT 13.7080 73.1835 13.7340 74.2770 ;
        RECT 13.6000 73.1835 13.6260 74.2770 ;
        RECT 13.4920 73.1835 13.5180 74.2770 ;
        RECT 13.3840 73.1835 13.4100 74.2770 ;
        RECT 13.2760 73.1835 13.3020 74.2770 ;
        RECT 13.1680 73.1835 13.1940 74.2770 ;
        RECT 13.0600 73.1835 13.0860 74.2770 ;
        RECT 12.9520 73.1835 12.9780 74.2770 ;
        RECT 12.8440 73.1835 12.8700 74.2770 ;
        RECT 12.7360 73.1835 12.7620 74.2770 ;
        RECT 12.6280 73.1835 12.6540 74.2770 ;
        RECT 12.5200 73.1835 12.5460 74.2770 ;
        RECT 12.4120 73.1835 12.4380 74.2770 ;
        RECT 12.3040 73.1835 12.3300 74.2770 ;
        RECT 12.1960 73.1835 12.2220 74.2770 ;
        RECT 12.0880 73.1835 12.1140 74.2770 ;
        RECT 11.9800 73.1835 12.0060 74.2770 ;
        RECT 11.8720 73.1835 11.8980 74.2770 ;
        RECT 11.7640 73.1835 11.7900 74.2770 ;
        RECT 11.6560 73.1835 11.6820 74.2770 ;
        RECT 11.5480 73.1835 11.5740 74.2770 ;
        RECT 11.4400 73.1835 11.4660 74.2770 ;
        RECT 11.3320 73.1835 11.3580 74.2770 ;
        RECT 11.2240 73.1835 11.2500 74.2770 ;
        RECT 11.1160 73.1835 11.1420 74.2770 ;
        RECT 11.0080 73.1835 11.0340 74.2770 ;
        RECT 10.9000 73.1835 10.9260 74.2770 ;
        RECT 10.7920 73.1835 10.8180 74.2770 ;
        RECT 10.6840 73.1835 10.7100 74.2770 ;
        RECT 10.5760 73.1835 10.6020 74.2770 ;
        RECT 10.4680 73.1835 10.4940 74.2770 ;
        RECT 10.3600 73.1835 10.3860 74.2770 ;
        RECT 10.2520 73.1835 10.2780 74.2770 ;
        RECT 10.1440 73.1835 10.1700 74.2770 ;
        RECT 10.0360 73.1835 10.0620 74.2770 ;
        RECT 9.9280 73.1835 9.9540 74.2770 ;
        RECT 9.8200 73.1835 9.8460 74.2770 ;
        RECT 9.7120 73.1835 9.7380 74.2770 ;
        RECT 9.6040 73.1835 9.6300 74.2770 ;
        RECT 9.4960 73.1835 9.5220 74.2770 ;
        RECT 9.3880 73.1835 9.4140 74.2770 ;
        RECT 9.2800 73.1835 9.3060 74.2770 ;
        RECT 9.1720 73.1835 9.1980 74.2770 ;
        RECT 9.0640 73.1835 9.0900 74.2770 ;
        RECT 8.9560 73.1835 8.9820 74.2770 ;
        RECT 8.8480 73.1835 8.8740 74.2770 ;
        RECT 8.7400 73.1835 8.7660 74.2770 ;
        RECT 8.6320 73.1835 8.6580 74.2770 ;
        RECT 8.5240 73.1835 8.5500 74.2770 ;
        RECT 8.4160 73.1835 8.4420 74.2770 ;
        RECT 8.3080 73.1835 8.3340 74.2770 ;
        RECT 8.2000 73.1835 8.2260 74.2770 ;
        RECT 8.0920 73.1835 8.1180 74.2770 ;
        RECT 7.9840 73.1835 8.0100 74.2770 ;
        RECT 7.8760 73.1835 7.9020 74.2770 ;
        RECT 7.7680 73.1835 7.7940 74.2770 ;
        RECT 7.6600 73.1835 7.6860 74.2770 ;
        RECT 7.5520 73.1835 7.5780 74.2770 ;
        RECT 7.4440 73.1835 7.4700 74.2770 ;
        RECT 7.3360 73.1835 7.3620 74.2770 ;
        RECT 7.2280 73.1835 7.2540 74.2770 ;
        RECT 7.1200 73.1835 7.1460 74.2770 ;
        RECT 7.0120 73.1835 7.0380 74.2770 ;
        RECT 6.9040 73.1835 6.9300 74.2770 ;
        RECT 6.7960 73.1835 6.8220 74.2770 ;
        RECT 6.6880 73.1835 6.7140 74.2770 ;
        RECT 6.5800 73.1835 6.6060 74.2770 ;
        RECT 6.4720 73.1835 6.4980 74.2770 ;
        RECT 6.3640 73.1835 6.3900 74.2770 ;
        RECT 6.2560 73.1835 6.2820 74.2770 ;
        RECT 6.1480 73.1835 6.1740 74.2770 ;
        RECT 6.0400 73.1835 6.0660 74.2770 ;
        RECT 5.9320 73.1835 5.9580 74.2770 ;
        RECT 5.8240 73.1835 5.8500 74.2770 ;
        RECT 5.7160 73.1835 5.7420 74.2770 ;
        RECT 5.6080 73.1835 5.6340 74.2770 ;
        RECT 5.5000 73.1835 5.5260 74.2770 ;
        RECT 5.3920 73.1835 5.4180 74.2770 ;
        RECT 5.2840 73.1835 5.3100 74.2770 ;
        RECT 5.1760 73.1835 5.2020 74.2770 ;
        RECT 5.0680 73.1835 5.0940 74.2770 ;
        RECT 4.9600 73.1835 4.9860 74.2770 ;
        RECT 4.8520 73.1835 4.8780 74.2770 ;
        RECT 4.7440 73.1835 4.7700 74.2770 ;
        RECT 4.6360 73.1835 4.6620 74.2770 ;
        RECT 4.5280 73.1835 4.5540 74.2770 ;
        RECT 4.4200 73.1835 4.4460 74.2770 ;
        RECT 4.3120 73.1835 4.3380 74.2770 ;
        RECT 4.2040 73.1835 4.2300 74.2770 ;
        RECT 4.0960 73.1835 4.1220 74.2770 ;
        RECT 3.9880 73.1835 4.0140 74.2770 ;
        RECT 3.8800 73.1835 3.9060 74.2770 ;
        RECT 3.7720 73.1835 3.7980 74.2770 ;
        RECT 3.6640 73.1835 3.6900 74.2770 ;
        RECT 3.5560 73.1835 3.5820 74.2770 ;
        RECT 3.4480 73.1835 3.4740 74.2770 ;
        RECT 3.3400 73.1835 3.3660 74.2770 ;
        RECT 3.2320 73.1835 3.2580 74.2770 ;
        RECT 3.1240 73.1835 3.1500 74.2770 ;
        RECT 3.0160 73.1835 3.0420 74.2770 ;
        RECT 2.9080 73.1835 2.9340 74.2770 ;
        RECT 2.8000 73.1835 2.8260 74.2770 ;
        RECT 2.6920 73.1835 2.7180 74.2770 ;
        RECT 2.5840 73.1835 2.6100 74.2770 ;
        RECT 2.4760 73.1835 2.5020 74.2770 ;
        RECT 2.3680 73.1835 2.3940 74.2770 ;
        RECT 2.2600 73.1835 2.2860 74.2770 ;
        RECT 2.1520 73.1835 2.1780 74.2770 ;
        RECT 2.0440 73.1835 2.0700 74.2770 ;
        RECT 1.9360 73.1835 1.9620 74.2770 ;
        RECT 1.8280 73.1835 1.8540 74.2770 ;
        RECT 1.7200 73.1835 1.7460 74.2770 ;
        RECT 1.6120 73.1835 1.6380 74.2770 ;
        RECT 1.5040 73.1835 1.5300 74.2770 ;
        RECT 1.3960 73.1835 1.4220 74.2770 ;
        RECT 1.2880 73.1835 1.3140 74.2770 ;
        RECT 1.1800 73.1835 1.2060 74.2770 ;
        RECT 1.0720 73.1835 1.0980 74.2770 ;
        RECT 0.9640 73.1835 0.9900 74.2770 ;
        RECT 0.8560 73.1835 0.8820 74.2770 ;
        RECT 0.7480 73.1835 0.7740 74.2770 ;
        RECT 0.6400 73.1835 0.6660 74.2770 ;
        RECT 0.5320 73.1835 0.5580 74.2770 ;
        RECT 0.4240 73.1835 0.4500 74.2770 ;
        RECT 0.3160 73.1835 0.3420 74.2770 ;
        RECT 0.2080 73.1835 0.2340 74.2770 ;
        RECT 0.0050 73.1835 0.0900 74.2770 ;
        RECT 15.5530 74.2635 15.6810 75.3570 ;
        RECT 15.5390 74.9290 15.6810 75.2515 ;
        RECT 15.3190 74.6560 15.4530 75.3570 ;
        RECT 15.2960 74.9910 15.4530 75.2490 ;
        RECT 15.3190 74.2635 15.4170 75.3570 ;
        RECT 15.3190 74.3845 15.4310 74.6240 ;
        RECT 15.3190 74.2635 15.4530 74.3525 ;
        RECT 15.0940 74.7140 15.2280 75.3570 ;
        RECT 15.0940 74.2635 15.1920 75.3570 ;
        RECT 14.6770 74.2635 14.7600 75.3570 ;
        RECT 14.6770 74.3520 14.7740 75.2875 ;
        RECT 30.2680 74.2635 30.3530 75.3570 ;
        RECT 30.1240 74.2635 30.1500 75.3570 ;
        RECT 30.0160 74.2635 30.0420 75.3570 ;
        RECT 29.9080 74.2635 29.9340 75.3570 ;
        RECT 29.8000 74.2635 29.8260 75.3570 ;
        RECT 29.6920 74.2635 29.7180 75.3570 ;
        RECT 29.5840 74.2635 29.6100 75.3570 ;
        RECT 29.4760 74.2635 29.5020 75.3570 ;
        RECT 29.3680 74.2635 29.3940 75.3570 ;
        RECT 29.2600 74.2635 29.2860 75.3570 ;
        RECT 29.1520 74.2635 29.1780 75.3570 ;
        RECT 29.0440 74.2635 29.0700 75.3570 ;
        RECT 28.9360 74.2635 28.9620 75.3570 ;
        RECT 28.8280 74.2635 28.8540 75.3570 ;
        RECT 28.7200 74.2635 28.7460 75.3570 ;
        RECT 28.6120 74.2635 28.6380 75.3570 ;
        RECT 28.5040 74.2635 28.5300 75.3570 ;
        RECT 28.3960 74.2635 28.4220 75.3570 ;
        RECT 28.2880 74.2635 28.3140 75.3570 ;
        RECT 28.1800 74.2635 28.2060 75.3570 ;
        RECT 28.0720 74.2635 28.0980 75.3570 ;
        RECT 27.9640 74.2635 27.9900 75.3570 ;
        RECT 27.8560 74.2635 27.8820 75.3570 ;
        RECT 27.7480 74.2635 27.7740 75.3570 ;
        RECT 27.6400 74.2635 27.6660 75.3570 ;
        RECT 27.5320 74.2635 27.5580 75.3570 ;
        RECT 27.4240 74.2635 27.4500 75.3570 ;
        RECT 27.3160 74.2635 27.3420 75.3570 ;
        RECT 27.2080 74.2635 27.2340 75.3570 ;
        RECT 27.1000 74.2635 27.1260 75.3570 ;
        RECT 26.9920 74.2635 27.0180 75.3570 ;
        RECT 26.8840 74.2635 26.9100 75.3570 ;
        RECT 26.7760 74.2635 26.8020 75.3570 ;
        RECT 26.6680 74.2635 26.6940 75.3570 ;
        RECT 26.5600 74.2635 26.5860 75.3570 ;
        RECT 26.4520 74.2635 26.4780 75.3570 ;
        RECT 26.3440 74.2635 26.3700 75.3570 ;
        RECT 26.2360 74.2635 26.2620 75.3570 ;
        RECT 26.1280 74.2635 26.1540 75.3570 ;
        RECT 26.0200 74.2635 26.0460 75.3570 ;
        RECT 25.9120 74.2635 25.9380 75.3570 ;
        RECT 25.8040 74.2635 25.8300 75.3570 ;
        RECT 25.6960 74.2635 25.7220 75.3570 ;
        RECT 25.5880 74.2635 25.6140 75.3570 ;
        RECT 25.4800 74.2635 25.5060 75.3570 ;
        RECT 25.3720 74.2635 25.3980 75.3570 ;
        RECT 25.2640 74.2635 25.2900 75.3570 ;
        RECT 25.1560 74.2635 25.1820 75.3570 ;
        RECT 25.0480 74.2635 25.0740 75.3570 ;
        RECT 24.9400 74.2635 24.9660 75.3570 ;
        RECT 24.8320 74.2635 24.8580 75.3570 ;
        RECT 24.7240 74.2635 24.7500 75.3570 ;
        RECT 24.6160 74.2635 24.6420 75.3570 ;
        RECT 24.5080 74.2635 24.5340 75.3570 ;
        RECT 24.4000 74.2635 24.4260 75.3570 ;
        RECT 24.2920 74.2635 24.3180 75.3570 ;
        RECT 24.1840 74.2635 24.2100 75.3570 ;
        RECT 24.0760 74.2635 24.1020 75.3570 ;
        RECT 23.9680 74.2635 23.9940 75.3570 ;
        RECT 23.8600 74.2635 23.8860 75.3570 ;
        RECT 23.7520 74.2635 23.7780 75.3570 ;
        RECT 23.6440 74.2635 23.6700 75.3570 ;
        RECT 23.5360 74.2635 23.5620 75.3570 ;
        RECT 23.4280 74.2635 23.4540 75.3570 ;
        RECT 23.3200 74.2635 23.3460 75.3570 ;
        RECT 23.2120 74.2635 23.2380 75.3570 ;
        RECT 23.1040 74.2635 23.1300 75.3570 ;
        RECT 22.9960 74.2635 23.0220 75.3570 ;
        RECT 22.8880 74.2635 22.9140 75.3570 ;
        RECT 22.7800 74.2635 22.8060 75.3570 ;
        RECT 22.6720 74.2635 22.6980 75.3570 ;
        RECT 22.5640 74.2635 22.5900 75.3570 ;
        RECT 22.4560 74.2635 22.4820 75.3570 ;
        RECT 22.3480 74.2635 22.3740 75.3570 ;
        RECT 22.2400 74.2635 22.2660 75.3570 ;
        RECT 22.1320 74.2635 22.1580 75.3570 ;
        RECT 22.0240 74.2635 22.0500 75.3570 ;
        RECT 21.9160 74.2635 21.9420 75.3570 ;
        RECT 21.8080 74.2635 21.8340 75.3570 ;
        RECT 21.7000 74.2635 21.7260 75.3570 ;
        RECT 21.5920 74.2635 21.6180 75.3570 ;
        RECT 21.4840 74.2635 21.5100 75.3570 ;
        RECT 21.3760 74.2635 21.4020 75.3570 ;
        RECT 21.2680 74.2635 21.2940 75.3570 ;
        RECT 21.1600 74.2635 21.1860 75.3570 ;
        RECT 21.0520 74.2635 21.0780 75.3570 ;
        RECT 20.9440 74.2635 20.9700 75.3570 ;
        RECT 20.8360 74.2635 20.8620 75.3570 ;
        RECT 20.7280 74.2635 20.7540 75.3570 ;
        RECT 20.6200 74.2635 20.6460 75.3570 ;
        RECT 20.5120 74.2635 20.5380 75.3570 ;
        RECT 20.4040 74.2635 20.4300 75.3570 ;
        RECT 20.2960 74.2635 20.3220 75.3570 ;
        RECT 20.1880 74.2635 20.2140 75.3570 ;
        RECT 20.0800 74.2635 20.1060 75.3570 ;
        RECT 19.9720 74.2635 19.9980 75.3570 ;
        RECT 19.8640 74.2635 19.8900 75.3570 ;
        RECT 19.7560 74.2635 19.7820 75.3570 ;
        RECT 19.6480 74.2635 19.6740 75.3570 ;
        RECT 19.5400 74.2635 19.5660 75.3570 ;
        RECT 19.4320 74.2635 19.4580 75.3570 ;
        RECT 19.3240 74.2635 19.3500 75.3570 ;
        RECT 19.2160 74.2635 19.2420 75.3570 ;
        RECT 19.1080 74.2635 19.1340 75.3570 ;
        RECT 19.0000 74.2635 19.0260 75.3570 ;
        RECT 18.8920 74.2635 18.9180 75.3570 ;
        RECT 18.7840 74.2635 18.8100 75.3570 ;
        RECT 18.6760 74.2635 18.7020 75.3570 ;
        RECT 18.5680 74.2635 18.5940 75.3570 ;
        RECT 18.4600 74.2635 18.4860 75.3570 ;
        RECT 18.3520 74.2635 18.3780 75.3570 ;
        RECT 18.2440 74.2635 18.2700 75.3570 ;
        RECT 18.1360 74.2635 18.1620 75.3570 ;
        RECT 18.0280 74.2635 18.0540 75.3570 ;
        RECT 17.9200 74.2635 17.9460 75.3570 ;
        RECT 17.8120 74.2635 17.8380 75.3570 ;
        RECT 17.7040 74.2635 17.7300 75.3570 ;
        RECT 17.5960 74.2635 17.6220 75.3570 ;
        RECT 17.4880 74.2635 17.5140 75.3570 ;
        RECT 17.3800 74.2635 17.4060 75.3570 ;
        RECT 17.2720 74.2635 17.2980 75.3570 ;
        RECT 17.1640 74.2635 17.1900 75.3570 ;
        RECT 17.0560 74.2635 17.0820 75.3570 ;
        RECT 16.9480 74.2635 16.9740 75.3570 ;
        RECT 16.8400 74.2635 16.8660 75.3570 ;
        RECT 16.7320 74.2635 16.7580 75.3570 ;
        RECT 16.6240 74.2635 16.6500 75.3570 ;
        RECT 16.5160 74.2635 16.5420 75.3570 ;
        RECT 16.4080 74.2635 16.4340 75.3570 ;
        RECT 16.3000 74.2635 16.3260 75.3570 ;
        RECT 16.0870 74.2635 16.1640 75.3570 ;
        RECT 14.1940 74.2635 14.2710 75.3570 ;
        RECT 14.0320 74.2635 14.0580 75.3570 ;
        RECT 13.9240 74.2635 13.9500 75.3570 ;
        RECT 13.8160 74.2635 13.8420 75.3570 ;
        RECT 13.7080 74.2635 13.7340 75.3570 ;
        RECT 13.6000 74.2635 13.6260 75.3570 ;
        RECT 13.4920 74.2635 13.5180 75.3570 ;
        RECT 13.3840 74.2635 13.4100 75.3570 ;
        RECT 13.2760 74.2635 13.3020 75.3570 ;
        RECT 13.1680 74.2635 13.1940 75.3570 ;
        RECT 13.0600 74.2635 13.0860 75.3570 ;
        RECT 12.9520 74.2635 12.9780 75.3570 ;
        RECT 12.8440 74.2635 12.8700 75.3570 ;
        RECT 12.7360 74.2635 12.7620 75.3570 ;
        RECT 12.6280 74.2635 12.6540 75.3570 ;
        RECT 12.5200 74.2635 12.5460 75.3570 ;
        RECT 12.4120 74.2635 12.4380 75.3570 ;
        RECT 12.3040 74.2635 12.3300 75.3570 ;
        RECT 12.1960 74.2635 12.2220 75.3570 ;
        RECT 12.0880 74.2635 12.1140 75.3570 ;
        RECT 11.9800 74.2635 12.0060 75.3570 ;
        RECT 11.8720 74.2635 11.8980 75.3570 ;
        RECT 11.7640 74.2635 11.7900 75.3570 ;
        RECT 11.6560 74.2635 11.6820 75.3570 ;
        RECT 11.5480 74.2635 11.5740 75.3570 ;
        RECT 11.4400 74.2635 11.4660 75.3570 ;
        RECT 11.3320 74.2635 11.3580 75.3570 ;
        RECT 11.2240 74.2635 11.2500 75.3570 ;
        RECT 11.1160 74.2635 11.1420 75.3570 ;
        RECT 11.0080 74.2635 11.0340 75.3570 ;
        RECT 10.9000 74.2635 10.9260 75.3570 ;
        RECT 10.7920 74.2635 10.8180 75.3570 ;
        RECT 10.6840 74.2635 10.7100 75.3570 ;
        RECT 10.5760 74.2635 10.6020 75.3570 ;
        RECT 10.4680 74.2635 10.4940 75.3570 ;
        RECT 10.3600 74.2635 10.3860 75.3570 ;
        RECT 10.2520 74.2635 10.2780 75.3570 ;
        RECT 10.1440 74.2635 10.1700 75.3570 ;
        RECT 10.0360 74.2635 10.0620 75.3570 ;
        RECT 9.9280 74.2635 9.9540 75.3570 ;
        RECT 9.8200 74.2635 9.8460 75.3570 ;
        RECT 9.7120 74.2635 9.7380 75.3570 ;
        RECT 9.6040 74.2635 9.6300 75.3570 ;
        RECT 9.4960 74.2635 9.5220 75.3570 ;
        RECT 9.3880 74.2635 9.4140 75.3570 ;
        RECT 9.2800 74.2635 9.3060 75.3570 ;
        RECT 9.1720 74.2635 9.1980 75.3570 ;
        RECT 9.0640 74.2635 9.0900 75.3570 ;
        RECT 8.9560 74.2635 8.9820 75.3570 ;
        RECT 8.8480 74.2635 8.8740 75.3570 ;
        RECT 8.7400 74.2635 8.7660 75.3570 ;
        RECT 8.6320 74.2635 8.6580 75.3570 ;
        RECT 8.5240 74.2635 8.5500 75.3570 ;
        RECT 8.4160 74.2635 8.4420 75.3570 ;
        RECT 8.3080 74.2635 8.3340 75.3570 ;
        RECT 8.2000 74.2635 8.2260 75.3570 ;
        RECT 8.0920 74.2635 8.1180 75.3570 ;
        RECT 7.9840 74.2635 8.0100 75.3570 ;
        RECT 7.8760 74.2635 7.9020 75.3570 ;
        RECT 7.7680 74.2635 7.7940 75.3570 ;
        RECT 7.6600 74.2635 7.6860 75.3570 ;
        RECT 7.5520 74.2635 7.5780 75.3570 ;
        RECT 7.4440 74.2635 7.4700 75.3570 ;
        RECT 7.3360 74.2635 7.3620 75.3570 ;
        RECT 7.2280 74.2635 7.2540 75.3570 ;
        RECT 7.1200 74.2635 7.1460 75.3570 ;
        RECT 7.0120 74.2635 7.0380 75.3570 ;
        RECT 6.9040 74.2635 6.9300 75.3570 ;
        RECT 6.7960 74.2635 6.8220 75.3570 ;
        RECT 6.6880 74.2635 6.7140 75.3570 ;
        RECT 6.5800 74.2635 6.6060 75.3570 ;
        RECT 6.4720 74.2635 6.4980 75.3570 ;
        RECT 6.3640 74.2635 6.3900 75.3570 ;
        RECT 6.2560 74.2635 6.2820 75.3570 ;
        RECT 6.1480 74.2635 6.1740 75.3570 ;
        RECT 6.0400 74.2635 6.0660 75.3570 ;
        RECT 5.9320 74.2635 5.9580 75.3570 ;
        RECT 5.8240 74.2635 5.8500 75.3570 ;
        RECT 5.7160 74.2635 5.7420 75.3570 ;
        RECT 5.6080 74.2635 5.6340 75.3570 ;
        RECT 5.5000 74.2635 5.5260 75.3570 ;
        RECT 5.3920 74.2635 5.4180 75.3570 ;
        RECT 5.2840 74.2635 5.3100 75.3570 ;
        RECT 5.1760 74.2635 5.2020 75.3570 ;
        RECT 5.0680 74.2635 5.0940 75.3570 ;
        RECT 4.9600 74.2635 4.9860 75.3570 ;
        RECT 4.8520 74.2635 4.8780 75.3570 ;
        RECT 4.7440 74.2635 4.7700 75.3570 ;
        RECT 4.6360 74.2635 4.6620 75.3570 ;
        RECT 4.5280 74.2635 4.5540 75.3570 ;
        RECT 4.4200 74.2635 4.4460 75.3570 ;
        RECT 4.3120 74.2635 4.3380 75.3570 ;
        RECT 4.2040 74.2635 4.2300 75.3570 ;
        RECT 4.0960 74.2635 4.1220 75.3570 ;
        RECT 3.9880 74.2635 4.0140 75.3570 ;
        RECT 3.8800 74.2635 3.9060 75.3570 ;
        RECT 3.7720 74.2635 3.7980 75.3570 ;
        RECT 3.6640 74.2635 3.6900 75.3570 ;
        RECT 3.5560 74.2635 3.5820 75.3570 ;
        RECT 3.4480 74.2635 3.4740 75.3570 ;
        RECT 3.3400 74.2635 3.3660 75.3570 ;
        RECT 3.2320 74.2635 3.2580 75.3570 ;
        RECT 3.1240 74.2635 3.1500 75.3570 ;
        RECT 3.0160 74.2635 3.0420 75.3570 ;
        RECT 2.9080 74.2635 2.9340 75.3570 ;
        RECT 2.8000 74.2635 2.8260 75.3570 ;
        RECT 2.6920 74.2635 2.7180 75.3570 ;
        RECT 2.5840 74.2635 2.6100 75.3570 ;
        RECT 2.4760 74.2635 2.5020 75.3570 ;
        RECT 2.3680 74.2635 2.3940 75.3570 ;
        RECT 2.2600 74.2635 2.2860 75.3570 ;
        RECT 2.1520 74.2635 2.1780 75.3570 ;
        RECT 2.0440 74.2635 2.0700 75.3570 ;
        RECT 1.9360 74.2635 1.9620 75.3570 ;
        RECT 1.8280 74.2635 1.8540 75.3570 ;
        RECT 1.7200 74.2635 1.7460 75.3570 ;
        RECT 1.6120 74.2635 1.6380 75.3570 ;
        RECT 1.5040 74.2635 1.5300 75.3570 ;
        RECT 1.3960 74.2635 1.4220 75.3570 ;
        RECT 1.2880 74.2635 1.3140 75.3570 ;
        RECT 1.1800 74.2635 1.2060 75.3570 ;
        RECT 1.0720 74.2635 1.0980 75.3570 ;
        RECT 0.9640 74.2635 0.9900 75.3570 ;
        RECT 0.8560 74.2635 0.8820 75.3570 ;
        RECT 0.7480 74.2635 0.7740 75.3570 ;
        RECT 0.6400 74.2635 0.6660 75.3570 ;
        RECT 0.5320 74.2635 0.5580 75.3570 ;
        RECT 0.4240 74.2635 0.4500 75.3570 ;
        RECT 0.3160 74.2635 0.3420 75.3570 ;
        RECT 0.2080 74.2635 0.2340 75.3570 ;
        RECT 0.0050 74.2635 0.0900 75.3570 ;
        RECT 15.5530 75.3435 15.6810 76.4370 ;
        RECT 15.5390 76.0090 15.6810 76.3315 ;
        RECT 15.3190 75.7360 15.4530 76.4370 ;
        RECT 15.2960 76.0710 15.4530 76.3290 ;
        RECT 15.3190 75.3435 15.4170 76.4370 ;
        RECT 15.3190 75.4645 15.4310 75.7040 ;
        RECT 15.3190 75.3435 15.4530 75.4325 ;
        RECT 15.0940 75.7940 15.2280 76.4370 ;
        RECT 15.0940 75.3435 15.1920 76.4370 ;
        RECT 14.6770 75.3435 14.7600 76.4370 ;
        RECT 14.6770 75.4320 14.7740 76.3675 ;
        RECT 30.2680 75.3435 30.3530 76.4370 ;
        RECT 30.1240 75.3435 30.1500 76.4370 ;
        RECT 30.0160 75.3435 30.0420 76.4370 ;
        RECT 29.9080 75.3435 29.9340 76.4370 ;
        RECT 29.8000 75.3435 29.8260 76.4370 ;
        RECT 29.6920 75.3435 29.7180 76.4370 ;
        RECT 29.5840 75.3435 29.6100 76.4370 ;
        RECT 29.4760 75.3435 29.5020 76.4370 ;
        RECT 29.3680 75.3435 29.3940 76.4370 ;
        RECT 29.2600 75.3435 29.2860 76.4370 ;
        RECT 29.1520 75.3435 29.1780 76.4370 ;
        RECT 29.0440 75.3435 29.0700 76.4370 ;
        RECT 28.9360 75.3435 28.9620 76.4370 ;
        RECT 28.8280 75.3435 28.8540 76.4370 ;
        RECT 28.7200 75.3435 28.7460 76.4370 ;
        RECT 28.6120 75.3435 28.6380 76.4370 ;
        RECT 28.5040 75.3435 28.5300 76.4370 ;
        RECT 28.3960 75.3435 28.4220 76.4370 ;
        RECT 28.2880 75.3435 28.3140 76.4370 ;
        RECT 28.1800 75.3435 28.2060 76.4370 ;
        RECT 28.0720 75.3435 28.0980 76.4370 ;
        RECT 27.9640 75.3435 27.9900 76.4370 ;
        RECT 27.8560 75.3435 27.8820 76.4370 ;
        RECT 27.7480 75.3435 27.7740 76.4370 ;
        RECT 27.6400 75.3435 27.6660 76.4370 ;
        RECT 27.5320 75.3435 27.5580 76.4370 ;
        RECT 27.4240 75.3435 27.4500 76.4370 ;
        RECT 27.3160 75.3435 27.3420 76.4370 ;
        RECT 27.2080 75.3435 27.2340 76.4370 ;
        RECT 27.1000 75.3435 27.1260 76.4370 ;
        RECT 26.9920 75.3435 27.0180 76.4370 ;
        RECT 26.8840 75.3435 26.9100 76.4370 ;
        RECT 26.7760 75.3435 26.8020 76.4370 ;
        RECT 26.6680 75.3435 26.6940 76.4370 ;
        RECT 26.5600 75.3435 26.5860 76.4370 ;
        RECT 26.4520 75.3435 26.4780 76.4370 ;
        RECT 26.3440 75.3435 26.3700 76.4370 ;
        RECT 26.2360 75.3435 26.2620 76.4370 ;
        RECT 26.1280 75.3435 26.1540 76.4370 ;
        RECT 26.0200 75.3435 26.0460 76.4370 ;
        RECT 25.9120 75.3435 25.9380 76.4370 ;
        RECT 25.8040 75.3435 25.8300 76.4370 ;
        RECT 25.6960 75.3435 25.7220 76.4370 ;
        RECT 25.5880 75.3435 25.6140 76.4370 ;
        RECT 25.4800 75.3435 25.5060 76.4370 ;
        RECT 25.3720 75.3435 25.3980 76.4370 ;
        RECT 25.2640 75.3435 25.2900 76.4370 ;
        RECT 25.1560 75.3435 25.1820 76.4370 ;
        RECT 25.0480 75.3435 25.0740 76.4370 ;
        RECT 24.9400 75.3435 24.9660 76.4370 ;
        RECT 24.8320 75.3435 24.8580 76.4370 ;
        RECT 24.7240 75.3435 24.7500 76.4370 ;
        RECT 24.6160 75.3435 24.6420 76.4370 ;
        RECT 24.5080 75.3435 24.5340 76.4370 ;
        RECT 24.4000 75.3435 24.4260 76.4370 ;
        RECT 24.2920 75.3435 24.3180 76.4370 ;
        RECT 24.1840 75.3435 24.2100 76.4370 ;
        RECT 24.0760 75.3435 24.1020 76.4370 ;
        RECT 23.9680 75.3435 23.9940 76.4370 ;
        RECT 23.8600 75.3435 23.8860 76.4370 ;
        RECT 23.7520 75.3435 23.7780 76.4370 ;
        RECT 23.6440 75.3435 23.6700 76.4370 ;
        RECT 23.5360 75.3435 23.5620 76.4370 ;
        RECT 23.4280 75.3435 23.4540 76.4370 ;
        RECT 23.3200 75.3435 23.3460 76.4370 ;
        RECT 23.2120 75.3435 23.2380 76.4370 ;
        RECT 23.1040 75.3435 23.1300 76.4370 ;
        RECT 22.9960 75.3435 23.0220 76.4370 ;
        RECT 22.8880 75.3435 22.9140 76.4370 ;
        RECT 22.7800 75.3435 22.8060 76.4370 ;
        RECT 22.6720 75.3435 22.6980 76.4370 ;
        RECT 22.5640 75.3435 22.5900 76.4370 ;
        RECT 22.4560 75.3435 22.4820 76.4370 ;
        RECT 22.3480 75.3435 22.3740 76.4370 ;
        RECT 22.2400 75.3435 22.2660 76.4370 ;
        RECT 22.1320 75.3435 22.1580 76.4370 ;
        RECT 22.0240 75.3435 22.0500 76.4370 ;
        RECT 21.9160 75.3435 21.9420 76.4370 ;
        RECT 21.8080 75.3435 21.8340 76.4370 ;
        RECT 21.7000 75.3435 21.7260 76.4370 ;
        RECT 21.5920 75.3435 21.6180 76.4370 ;
        RECT 21.4840 75.3435 21.5100 76.4370 ;
        RECT 21.3760 75.3435 21.4020 76.4370 ;
        RECT 21.2680 75.3435 21.2940 76.4370 ;
        RECT 21.1600 75.3435 21.1860 76.4370 ;
        RECT 21.0520 75.3435 21.0780 76.4370 ;
        RECT 20.9440 75.3435 20.9700 76.4370 ;
        RECT 20.8360 75.3435 20.8620 76.4370 ;
        RECT 20.7280 75.3435 20.7540 76.4370 ;
        RECT 20.6200 75.3435 20.6460 76.4370 ;
        RECT 20.5120 75.3435 20.5380 76.4370 ;
        RECT 20.4040 75.3435 20.4300 76.4370 ;
        RECT 20.2960 75.3435 20.3220 76.4370 ;
        RECT 20.1880 75.3435 20.2140 76.4370 ;
        RECT 20.0800 75.3435 20.1060 76.4370 ;
        RECT 19.9720 75.3435 19.9980 76.4370 ;
        RECT 19.8640 75.3435 19.8900 76.4370 ;
        RECT 19.7560 75.3435 19.7820 76.4370 ;
        RECT 19.6480 75.3435 19.6740 76.4370 ;
        RECT 19.5400 75.3435 19.5660 76.4370 ;
        RECT 19.4320 75.3435 19.4580 76.4370 ;
        RECT 19.3240 75.3435 19.3500 76.4370 ;
        RECT 19.2160 75.3435 19.2420 76.4370 ;
        RECT 19.1080 75.3435 19.1340 76.4370 ;
        RECT 19.0000 75.3435 19.0260 76.4370 ;
        RECT 18.8920 75.3435 18.9180 76.4370 ;
        RECT 18.7840 75.3435 18.8100 76.4370 ;
        RECT 18.6760 75.3435 18.7020 76.4370 ;
        RECT 18.5680 75.3435 18.5940 76.4370 ;
        RECT 18.4600 75.3435 18.4860 76.4370 ;
        RECT 18.3520 75.3435 18.3780 76.4370 ;
        RECT 18.2440 75.3435 18.2700 76.4370 ;
        RECT 18.1360 75.3435 18.1620 76.4370 ;
        RECT 18.0280 75.3435 18.0540 76.4370 ;
        RECT 17.9200 75.3435 17.9460 76.4370 ;
        RECT 17.8120 75.3435 17.8380 76.4370 ;
        RECT 17.7040 75.3435 17.7300 76.4370 ;
        RECT 17.5960 75.3435 17.6220 76.4370 ;
        RECT 17.4880 75.3435 17.5140 76.4370 ;
        RECT 17.3800 75.3435 17.4060 76.4370 ;
        RECT 17.2720 75.3435 17.2980 76.4370 ;
        RECT 17.1640 75.3435 17.1900 76.4370 ;
        RECT 17.0560 75.3435 17.0820 76.4370 ;
        RECT 16.9480 75.3435 16.9740 76.4370 ;
        RECT 16.8400 75.3435 16.8660 76.4370 ;
        RECT 16.7320 75.3435 16.7580 76.4370 ;
        RECT 16.6240 75.3435 16.6500 76.4370 ;
        RECT 16.5160 75.3435 16.5420 76.4370 ;
        RECT 16.4080 75.3435 16.4340 76.4370 ;
        RECT 16.3000 75.3435 16.3260 76.4370 ;
        RECT 16.0870 75.3435 16.1640 76.4370 ;
        RECT 14.1940 75.3435 14.2710 76.4370 ;
        RECT 14.0320 75.3435 14.0580 76.4370 ;
        RECT 13.9240 75.3435 13.9500 76.4370 ;
        RECT 13.8160 75.3435 13.8420 76.4370 ;
        RECT 13.7080 75.3435 13.7340 76.4370 ;
        RECT 13.6000 75.3435 13.6260 76.4370 ;
        RECT 13.4920 75.3435 13.5180 76.4370 ;
        RECT 13.3840 75.3435 13.4100 76.4370 ;
        RECT 13.2760 75.3435 13.3020 76.4370 ;
        RECT 13.1680 75.3435 13.1940 76.4370 ;
        RECT 13.0600 75.3435 13.0860 76.4370 ;
        RECT 12.9520 75.3435 12.9780 76.4370 ;
        RECT 12.8440 75.3435 12.8700 76.4370 ;
        RECT 12.7360 75.3435 12.7620 76.4370 ;
        RECT 12.6280 75.3435 12.6540 76.4370 ;
        RECT 12.5200 75.3435 12.5460 76.4370 ;
        RECT 12.4120 75.3435 12.4380 76.4370 ;
        RECT 12.3040 75.3435 12.3300 76.4370 ;
        RECT 12.1960 75.3435 12.2220 76.4370 ;
        RECT 12.0880 75.3435 12.1140 76.4370 ;
        RECT 11.9800 75.3435 12.0060 76.4370 ;
        RECT 11.8720 75.3435 11.8980 76.4370 ;
        RECT 11.7640 75.3435 11.7900 76.4370 ;
        RECT 11.6560 75.3435 11.6820 76.4370 ;
        RECT 11.5480 75.3435 11.5740 76.4370 ;
        RECT 11.4400 75.3435 11.4660 76.4370 ;
        RECT 11.3320 75.3435 11.3580 76.4370 ;
        RECT 11.2240 75.3435 11.2500 76.4370 ;
        RECT 11.1160 75.3435 11.1420 76.4370 ;
        RECT 11.0080 75.3435 11.0340 76.4370 ;
        RECT 10.9000 75.3435 10.9260 76.4370 ;
        RECT 10.7920 75.3435 10.8180 76.4370 ;
        RECT 10.6840 75.3435 10.7100 76.4370 ;
        RECT 10.5760 75.3435 10.6020 76.4370 ;
        RECT 10.4680 75.3435 10.4940 76.4370 ;
        RECT 10.3600 75.3435 10.3860 76.4370 ;
        RECT 10.2520 75.3435 10.2780 76.4370 ;
        RECT 10.1440 75.3435 10.1700 76.4370 ;
        RECT 10.0360 75.3435 10.0620 76.4370 ;
        RECT 9.9280 75.3435 9.9540 76.4370 ;
        RECT 9.8200 75.3435 9.8460 76.4370 ;
        RECT 9.7120 75.3435 9.7380 76.4370 ;
        RECT 9.6040 75.3435 9.6300 76.4370 ;
        RECT 9.4960 75.3435 9.5220 76.4370 ;
        RECT 9.3880 75.3435 9.4140 76.4370 ;
        RECT 9.2800 75.3435 9.3060 76.4370 ;
        RECT 9.1720 75.3435 9.1980 76.4370 ;
        RECT 9.0640 75.3435 9.0900 76.4370 ;
        RECT 8.9560 75.3435 8.9820 76.4370 ;
        RECT 8.8480 75.3435 8.8740 76.4370 ;
        RECT 8.7400 75.3435 8.7660 76.4370 ;
        RECT 8.6320 75.3435 8.6580 76.4370 ;
        RECT 8.5240 75.3435 8.5500 76.4370 ;
        RECT 8.4160 75.3435 8.4420 76.4370 ;
        RECT 8.3080 75.3435 8.3340 76.4370 ;
        RECT 8.2000 75.3435 8.2260 76.4370 ;
        RECT 8.0920 75.3435 8.1180 76.4370 ;
        RECT 7.9840 75.3435 8.0100 76.4370 ;
        RECT 7.8760 75.3435 7.9020 76.4370 ;
        RECT 7.7680 75.3435 7.7940 76.4370 ;
        RECT 7.6600 75.3435 7.6860 76.4370 ;
        RECT 7.5520 75.3435 7.5780 76.4370 ;
        RECT 7.4440 75.3435 7.4700 76.4370 ;
        RECT 7.3360 75.3435 7.3620 76.4370 ;
        RECT 7.2280 75.3435 7.2540 76.4370 ;
        RECT 7.1200 75.3435 7.1460 76.4370 ;
        RECT 7.0120 75.3435 7.0380 76.4370 ;
        RECT 6.9040 75.3435 6.9300 76.4370 ;
        RECT 6.7960 75.3435 6.8220 76.4370 ;
        RECT 6.6880 75.3435 6.7140 76.4370 ;
        RECT 6.5800 75.3435 6.6060 76.4370 ;
        RECT 6.4720 75.3435 6.4980 76.4370 ;
        RECT 6.3640 75.3435 6.3900 76.4370 ;
        RECT 6.2560 75.3435 6.2820 76.4370 ;
        RECT 6.1480 75.3435 6.1740 76.4370 ;
        RECT 6.0400 75.3435 6.0660 76.4370 ;
        RECT 5.9320 75.3435 5.9580 76.4370 ;
        RECT 5.8240 75.3435 5.8500 76.4370 ;
        RECT 5.7160 75.3435 5.7420 76.4370 ;
        RECT 5.6080 75.3435 5.6340 76.4370 ;
        RECT 5.5000 75.3435 5.5260 76.4370 ;
        RECT 5.3920 75.3435 5.4180 76.4370 ;
        RECT 5.2840 75.3435 5.3100 76.4370 ;
        RECT 5.1760 75.3435 5.2020 76.4370 ;
        RECT 5.0680 75.3435 5.0940 76.4370 ;
        RECT 4.9600 75.3435 4.9860 76.4370 ;
        RECT 4.8520 75.3435 4.8780 76.4370 ;
        RECT 4.7440 75.3435 4.7700 76.4370 ;
        RECT 4.6360 75.3435 4.6620 76.4370 ;
        RECT 4.5280 75.3435 4.5540 76.4370 ;
        RECT 4.4200 75.3435 4.4460 76.4370 ;
        RECT 4.3120 75.3435 4.3380 76.4370 ;
        RECT 4.2040 75.3435 4.2300 76.4370 ;
        RECT 4.0960 75.3435 4.1220 76.4370 ;
        RECT 3.9880 75.3435 4.0140 76.4370 ;
        RECT 3.8800 75.3435 3.9060 76.4370 ;
        RECT 3.7720 75.3435 3.7980 76.4370 ;
        RECT 3.6640 75.3435 3.6900 76.4370 ;
        RECT 3.5560 75.3435 3.5820 76.4370 ;
        RECT 3.4480 75.3435 3.4740 76.4370 ;
        RECT 3.3400 75.3435 3.3660 76.4370 ;
        RECT 3.2320 75.3435 3.2580 76.4370 ;
        RECT 3.1240 75.3435 3.1500 76.4370 ;
        RECT 3.0160 75.3435 3.0420 76.4370 ;
        RECT 2.9080 75.3435 2.9340 76.4370 ;
        RECT 2.8000 75.3435 2.8260 76.4370 ;
        RECT 2.6920 75.3435 2.7180 76.4370 ;
        RECT 2.5840 75.3435 2.6100 76.4370 ;
        RECT 2.4760 75.3435 2.5020 76.4370 ;
        RECT 2.3680 75.3435 2.3940 76.4370 ;
        RECT 2.2600 75.3435 2.2860 76.4370 ;
        RECT 2.1520 75.3435 2.1780 76.4370 ;
        RECT 2.0440 75.3435 2.0700 76.4370 ;
        RECT 1.9360 75.3435 1.9620 76.4370 ;
        RECT 1.8280 75.3435 1.8540 76.4370 ;
        RECT 1.7200 75.3435 1.7460 76.4370 ;
        RECT 1.6120 75.3435 1.6380 76.4370 ;
        RECT 1.5040 75.3435 1.5300 76.4370 ;
        RECT 1.3960 75.3435 1.4220 76.4370 ;
        RECT 1.2880 75.3435 1.3140 76.4370 ;
        RECT 1.1800 75.3435 1.2060 76.4370 ;
        RECT 1.0720 75.3435 1.0980 76.4370 ;
        RECT 0.9640 75.3435 0.9900 76.4370 ;
        RECT 0.8560 75.3435 0.8820 76.4370 ;
        RECT 0.7480 75.3435 0.7740 76.4370 ;
        RECT 0.6400 75.3435 0.6660 76.4370 ;
        RECT 0.5320 75.3435 0.5580 76.4370 ;
        RECT 0.4240 75.3435 0.4500 76.4370 ;
        RECT 0.3160 75.3435 0.3420 76.4370 ;
        RECT 0.2080 75.3435 0.2340 76.4370 ;
        RECT 0.0050 75.3435 0.0900 76.4370 ;
        RECT 15.5530 76.4235 15.6810 77.5170 ;
        RECT 15.5390 77.0890 15.6810 77.4115 ;
        RECT 15.3190 76.8160 15.4530 77.5170 ;
        RECT 15.2960 77.1510 15.4530 77.4090 ;
        RECT 15.3190 76.4235 15.4170 77.5170 ;
        RECT 15.3190 76.5445 15.4310 76.7840 ;
        RECT 15.3190 76.4235 15.4530 76.5125 ;
        RECT 15.0940 76.8740 15.2280 77.5170 ;
        RECT 15.0940 76.4235 15.1920 77.5170 ;
        RECT 14.6770 76.4235 14.7600 77.5170 ;
        RECT 14.6770 76.5120 14.7740 77.4475 ;
        RECT 30.2680 76.4235 30.3530 77.5170 ;
        RECT 30.1240 76.4235 30.1500 77.5170 ;
        RECT 30.0160 76.4235 30.0420 77.5170 ;
        RECT 29.9080 76.4235 29.9340 77.5170 ;
        RECT 29.8000 76.4235 29.8260 77.5170 ;
        RECT 29.6920 76.4235 29.7180 77.5170 ;
        RECT 29.5840 76.4235 29.6100 77.5170 ;
        RECT 29.4760 76.4235 29.5020 77.5170 ;
        RECT 29.3680 76.4235 29.3940 77.5170 ;
        RECT 29.2600 76.4235 29.2860 77.5170 ;
        RECT 29.1520 76.4235 29.1780 77.5170 ;
        RECT 29.0440 76.4235 29.0700 77.5170 ;
        RECT 28.9360 76.4235 28.9620 77.5170 ;
        RECT 28.8280 76.4235 28.8540 77.5170 ;
        RECT 28.7200 76.4235 28.7460 77.5170 ;
        RECT 28.6120 76.4235 28.6380 77.5170 ;
        RECT 28.5040 76.4235 28.5300 77.5170 ;
        RECT 28.3960 76.4235 28.4220 77.5170 ;
        RECT 28.2880 76.4235 28.3140 77.5170 ;
        RECT 28.1800 76.4235 28.2060 77.5170 ;
        RECT 28.0720 76.4235 28.0980 77.5170 ;
        RECT 27.9640 76.4235 27.9900 77.5170 ;
        RECT 27.8560 76.4235 27.8820 77.5170 ;
        RECT 27.7480 76.4235 27.7740 77.5170 ;
        RECT 27.6400 76.4235 27.6660 77.5170 ;
        RECT 27.5320 76.4235 27.5580 77.5170 ;
        RECT 27.4240 76.4235 27.4500 77.5170 ;
        RECT 27.3160 76.4235 27.3420 77.5170 ;
        RECT 27.2080 76.4235 27.2340 77.5170 ;
        RECT 27.1000 76.4235 27.1260 77.5170 ;
        RECT 26.9920 76.4235 27.0180 77.5170 ;
        RECT 26.8840 76.4235 26.9100 77.5170 ;
        RECT 26.7760 76.4235 26.8020 77.5170 ;
        RECT 26.6680 76.4235 26.6940 77.5170 ;
        RECT 26.5600 76.4235 26.5860 77.5170 ;
        RECT 26.4520 76.4235 26.4780 77.5170 ;
        RECT 26.3440 76.4235 26.3700 77.5170 ;
        RECT 26.2360 76.4235 26.2620 77.5170 ;
        RECT 26.1280 76.4235 26.1540 77.5170 ;
        RECT 26.0200 76.4235 26.0460 77.5170 ;
        RECT 25.9120 76.4235 25.9380 77.5170 ;
        RECT 25.8040 76.4235 25.8300 77.5170 ;
        RECT 25.6960 76.4235 25.7220 77.5170 ;
        RECT 25.5880 76.4235 25.6140 77.5170 ;
        RECT 25.4800 76.4235 25.5060 77.5170 ;
        RECT 25.3720 76.4235 25.3980 77.5170 ;
        RECT 25.2640 76.4235 25.2900 77.5170 ;
        RECT 25.1560 76.4235 25.1820 77.5170 ;
        RECT 25.0480 76.4235 25.0740 77.5170 ;
        RECT 24.9400 76.4235 24.9660 77.5170 ;
        RECT 24.8320 76.4235 24.8580 77.5170 ;
        RECT 24.7240 76.4235 24.7500 77.5170 ;
        RECT 24.6160 76.4235 24.6420 77.5170 ;
        RECT 24.5080 76.4235 24.5340 77.5170 ;
        RECT 24.4000 76.4235 24.4260 77.5170 ;
        RECT 24.2920 76.4235 24.3180 77.5170 ;
        RECT 24.1840 76.4235 24.2100 77.5170 ;
        RECT 24.0760 76.4235 24.1020 77.5170 ;
        RECT 23.9680 76.4235 23.9940 77.5170 ;
        RECT 23.8600 76.4235 23.8860 77.5170 ;
        RECT 23.7520 76.4235 23.7780 77.5170 ;
        RECT 23.6440 76.4235 23.6700 77.5170 ;
        RECT 23.5360 76.4235 23.5620 77.5170 ;
        RECT 23.4280 76.4235 23.4540 77.5170 ;
        RECT 23.3200 76.4235 23.3460 77.5170 ;
        RECT 23.2120 76.4235 23.2380 77.5170 ;
        RECT 23.1040 76.4235 23.1300 77.5170 ;
        RECT 22.9960 76.4235 23.0220 77.5170 ;
        RECT 22.8880 76.4235 22.9140 77.5170 ;
        RECT 22.7800 76.4235 22.8060 77.5170 ;
        RECT 22.6720 76.4235 22.6980 77.5170 ;
        RECT 22.5640 76.4235 22.5900 77.5170 ;
        RECT 22.4560 76.4235 22.4820 77.5170 ;
        RECT 22.3480 76.4235 22.3740 77.5170 ;
        RECT 22.2400 76.4235 22.2660 77.5170 ;
        RECT 22.1320 76.4235 22.1580 77.5170 ;
        RECT 22.0240 76.4235 22.0500 77.5170 ;
        RECT 21.9160 76.4235 21.9420 77.5170 ;
        RECT 21.8080 76.4235 21.8340 77.5170 ;
        RECT 21.7000 76.4235 21.7260 77.5170 ;
        RECT 21.5920 76.4235 21.6180 77.5170 ;
        RECT 21.4840 76.4235 21.5100 77.5170 ;
        RECT 21.3760 76.4235 21.4020 77.5170 ;
        RECT 21.2680 76.4235 21.2940 77.5170 ;
        RECT 21.1600 76.4235 21.1860 77.5170 ;
        RECT 21.0520 76.4235 21.0780 77.5170 ;
        RECT 20.9440 76.4235 20.9700 77.5170 ;
        RECT 20.8360 76.4235 20.8620 77.5170 ;
        RECT 20.7280 76.4235 20.7540 77.5170 ;
        RECT 20.6200 76.4235 20.6460 77.5170 ;
        RECT 20.5120 76.4235 20.5380 77.5170 ;
        RECT 20.4040 76.4235 20.4300 77.5170 ;
        RECT 20.2960 76.4235 20.3220 77.5170 ;
        RECT 20.1880 76.4235 20.2140 77.5170 ;
        RECT 20.0800 76.4235 20.1060 77.5170 ;
        RECT 19.9720 76.4235 19.9980 77.5170 ;
        RECT 19.8640 76.4235 19.8900 77.5170 ;
        RECT 19.7560 76.4235 19.7820 77.5170 ;
        RECT 19.6480 76.4235 19.6740 77.5170 ;
        RECT 19.5400 76.4235 19.5660 77.5170 ;
        RECT 19.4320 76.4235 19.4580 77.5170 ;
        RECT 19.3240 76.4235 19.3500 77.5170 ;
        RECT 19.2160 76.4235 19.2420 77.5170 ;
        RECT 19.1080 76.4235 19.1340 77.5170 ;
        RECT 19.0000 76.4235 19.0260 77.5170 ;
        RECT 18.8920 76.4235 18.9180 77.5170 ;
        RECT 18.7840 76.4235 18.8100 77.5170 ;
        RECT 18.6760 76.4235 18.7020 77.5170 ;
        RECT 18.5680 76.4235 18.5940 77.5170 ;
        RECT 18.4600 76.4235 18.4860 77.5170 ;
        RECT 18.3520 76.4235 18.3780 77.5170 ;
        RECT 18.2440 76.4235 18.2700 77.5170 ;
        RECT 18.1360 76.4235 18.1620 77.5170 ;
        RECT 18.0280 76.4235 18.0540 77.5170 ;
        RECT 17.9200 76.4235 17.9460 77.5170 ;
        RECT 17.8120 76.4235 17.8380 77.5170 ;
        RECT 17.7040 76.4235 17.7300 77.5170 ;
        RECT 17.5960 76.4235 17.6220 77.5170 ;
        RECT 17.4880 76.4235 17.5140 77.5170 ;
        RECT 17.3800 76.4235 17.4060 77.5170 ;
        RECT 17.2720 76.4235 17.2980 77.5170 ;
        RECT 17.1640 76.4235 17.1900 77.5170 ;
        RECT 17.0560 76.4235 17.0820 77.5170 ;
        RECT 16.9480 76.4235 16.9740 77.5170 ;
        RECT 16.8400 76.4235 16.8660 77.5170 ;
        RECT 16.7320 76.4235 16.7580 77.5170 ;
        RECT 16.6240 76.4235 16.6500 77.5170 ;
        RECT 16.5160 76.4235 16.5420 77.5170 ;
        RECT 16.4080 76.4235 16.4340 77.5170 ;
        RECT 16.3000 76.4235 16.3260 77.5170 ;
        RECT 16.0870 76.4235 16.1640 77.5170 ;
        RECT 14.1940 76.4235 14.2710 77.5170 ;
        RECT 14.0320 76.4235 14.0580 77.5170 ;
        RECT 13.9240 76.4235 13.9500 77.5170 ;
        RECT 13.8160 76.4235 13.8420 77.5170 ;
        RECT 13.7080 76.4235 13.7340 77.5170 ;
        RECT 13.6000 76.4235 13.6260 77.5170 ;
        RECT 13.4920 76.4235 13.5180 77.5170 ;
        RECT 13.3840 76.4235 13.4100 77.5170 ;
        RECT 13.2760 76.4235 13.3020 77.5170 ;
        RECT 13.1680 76.4235 13.1940 77.5170 ;
        RECT 13.0600 76.4235 13.0860 77.5170 ;
        RECT 12.9520 76.4235 12.9780 77.5170 ;
        RECT 12.8440 76.4235 12.8700 77.5170 ;
        RECT 12.7360 76.4235 12.7620 77.5170 ;
        RECT 12.6280 76.4235 12.6540 77.5170 ;
        RECT 12.5200 76.4235 12.5460 77.5170 ;
        RECT 12.4120 76.4235 12.4380 77.5170 ;
        RECT 12.3040 76.4235 12.3300 77.5170 ;
        RECT 12.1960 76.4235 12.2220 77.5170 ;
        RECT 12.0880 76.4235 12.1140 77.5170 ;
        RECT 11.9800 76.4235 12.0060 77.5170 ;
        RECT 11.8720 76.4235 11.8980 77.5170 ;
        RECT 11.7640 76.4235 11.7900 77.5170 ;
        RECT 11.6560 76.4235 11.6820 77.5170 ;
        RECT 11.5480 76.4235 11.5740 77.5170 ;
        RECT 11.4400 76.4235 11.4660 77.5170 ;
        RECT 11.3320 76.4235 11.3580 77.5170 ;
        RECT 11.2240 76.4235 11.2500 77.5170 ;
        RECT 11.1160 76.4235 11.1420 77.5170 ;
        RECT 11.0080 76.4235 11.0340 77.5170 ;
        RECT 10.9000 76.4235 10.9260 77.5170 ;
        RECT 10.7920 76.4235 10.8180 77.5170 ;
        RECT 10.6840 76.4235 10.7100 77.5170 ;
        RECT 10.5760 76.4235 10.6020 77.5170 ;
        RECT 10.4680 76.4235 10.4940 77.5170 ;
        RECT 10.3600 76.4235 10.3860 77.5170 ;
        RECT 10.2520 76.4235 10.2780 77.5170 ;
        RECT 10.1440 76.4235 10.1700 77.5170 ;
        RECT 10.0360 76.4235 10.0620 77.5170 ;
        RECT 9.9280 76.4235 9.9540 77.5170 ;
        RECT 9.8200 76.4235 9.8460 77.5170 ;
        RECT 9.7120 76.4235 9.7380 77.5170 ;
        RECT 9.6040 76.4235 9.6300 77.5170 ;
        RECT 9.4960 76.4235 9.5220 77.5170 ;
        RECT 9.3880 76.4235 9.4140 77.5170 ;
        RECT 9.2800 76.4235 9.3060 77.5170 ;
        RECT 9.1720 76.4235 9.1980 77.5170 ;
        RECT 9.0640 76.4235 9.0900 77.5170 ;
        RECT 8.9560 76.4235 8.9820 77.5170 ;
        RECT 8.8480 76.4235 8.8740 77.5170 ;
        RECT 8.7400 76.4235 8.7660 77.5170 ;
        RECT 8.6320 76.4235 8.6580 77.5170 ;
        RECT 8.5240 76.4235 8.5500 77.5170 ;
        RECT 8.4160 76.4235 8.4420 77.5170 ;
        RECT 8.3080 76.4235 8.3340 77.5170 ;
        RECT 8.2000 76.4235 8.2260 77.5170 ;
        RECT 8.0920 76.4235 8.1180 77.5170 ;
        RECT 7.9840 76.4235 8.0100 77.5170 ;
        RECT 7.8760 76.4235 7.9020 77.5170 ;
        RECT 7.7680 76.4235 7.7940 77.5170 ;
        RECT 7.6600 76.4235 7.6860 77.5170 ;
        RECT 7.5520 76.4235 7.5780 77.5170 ;
        RECT 7.4440 76.4235 7.4700 77.5170 ;
        RECT 7.3360 76.4235 7.3620 77.5170 ;
        RECT 7.2280 76.4235 7.2540 77.5170 ;
        RECT 7.1200 76.4235 7.1460 77.5170 ;
        RECT 7.0120 76.4235 7.0380 77.5170 ;
        RECT 6.9040 76.4235 6.9300 77.5170 ;
        RECT 6.7960 76.4235 6.8220 77.5170 ;
        RECT 6.6880 76.4235 6.7140 77.5170 ;
        RECT 6.5800 76.4235 6.6060 77.5170 ;
        RECT 6.4720 76.4235 6.4980 77.5170 ;
        RECT 6.3640 76.4235 6.3900 77.5170 ;
        RECT 6.2560 76.4235 6.2820 77.5170 ;
        RECT 6.1480 76.4235 6.1740 77.5170 ;
        RECT 6.0400 76.4235 6.0660 77.5170 ;
        RECT 5.9320 76.4235 5.9580 77.5170 ;
        RECT 5.8240 76.4235 5.8500 77.5170 ;
        RECT 5.7160 76.4235 5.7420 77.5170 ;
        RECT 5.6080 76.4235 5.6340 77.5170 ;
        RECT 5.5000 76.4235 5.5260 77.5170 ;
        RECT 5.3920 76.4235 5.4180 77.5170 ;
        RECT 5.2840 76.4235 5.3100 77.5170 ;
        RECT 5.1760 76.4235 5.2020 77.5170 ;
        RECT 5.0680 76.4235 5.0940 77.5170 ;
        RECT 4.9600 76.4235 4.9860 77.5170 ;
        RECT 4.8520 76.4235 4.8780 77.5170 ;
        RECT 4.7440 76.4235 4.7700 77.5170 ;
        RECT 4.6360 76.4235 4.6620 77.5170 ;
        RECT 4.5280 76.4235 4.5540 77.5170 ;
        RECT 4.4200 76.4235 4.4460 77.5170 ;
        RECT 4.3120 76.4235 4.3380 77.5170 ;
        RECT 4.2040 76.4235 4.2300 77.5170 ;
        RECT 4.0960 76.4235 4.1220 77.5170 ;
        RECT 3.9880 76.4235 4.0140 77.5170 ;
        RECT 3.8800 76.4235 3.9060 77.5170 ;
        RECT 3.7720 76.4235 3.7980 77.5170 ;
        RECT 3.6640 76.4235 3.6900 77.5170 ;
        RECT 3.5560 76.4235 3.5820 77.5170 ;
        RECT 3.4480 76.4235 3.4740 77.5170 ;
        RECT 3.3400 76.4235 3.3660 77.5170 ;
        RECT 3.2320 76.4235 3.2580 77.5170 ;
        RECT 3.1240 76.4235 3.1500 77.5170 ;
        RECT 3.0160 76.4235 3.0420 77.5170 ;
        RECT 2.9080 76.4235 2.9340 77.5170 ;
        RECT 2.8000 76.4235 2.8260 77.5170 ;
        RECT 2.6920 76.4235 2.7180 77.5170 ;
        RECT 2.5840 76.4235 2.6100 77.5170 ;
        RECT 2.4760 76.4235 2.5020 77.5170 ;
        RECT 2.3680 76.4235 2.3940 77.5170 ;
        RECT 2.2600 76.4235 2.2860 77.5170 ;
        RECT 2.1520 76.4235 2.1780 77.5170 ;
        RECT 2.0440 76.4235 2.0700 77.5170 ;
        RECT 1.9360 76.4235 1.9620 77.5170 ;
        RECT 1.8280 76.4235 1.8540 77.5170 ;
        RECT 1.7200 76.4235 1.7460 77.5170 ;
        RECT 1.6120 76.4235 1.6380 77.5170 ;
        RECT 1.5040 76.4235 1.5300 77.5170 ;
        RECT 1.3960 76.4235 1.4220 77.5170 ;
        RECT 1.2880 76.4235 1.3140 77.5170 ;
        RECT 1.1800 76.4235 1.2060 77.5170 ;
        RECT 1.0720 76.4235 1.0980 77.5170 ;
        RECT 0.9640 76.4235 0.9900 77.5170 ;
        RECT 0.8560 76.4235 0.8820 77.5170 ;
        RECT 0.7480 76.4235 0.7740 77.5170 ;
        RECT 0.6400 76.4235 0.6660 77.5170 ;
        RECT 0.5320 76.4235 0.5580 77.5170 ;
        RECT 0.4240 76.4235 0.4500 77.5170 ;
        RECT 0.3160 76.4235 0.3420 77.5170 ;
        RECT 0.2080 76.4235 0.2340 77.5170 ;
        RECT 0.0050 76.4235 0.0900 77.5170 ;
  LAYER V3 SPACING 0.018  ;
      RECT 0.0050 1.2200 30.3530 1.3500 ;
      RECT 30.2360 0.2565 30.3530 1.3500 ;
      RECT 16.2140 1.1240 30.2180 1.3500 ;
      RECT 14.8820 1.1240 16.1960 1.3500 ;
      RECT 14.1620 0.2565 14.7920 1.3500 ;
      RECT 0.1400 1.1240 14.1440 1.3500 ;
      RECT 0.0050 0.2565 0.1220 1.3500 ;
      RECT 30.2000 0.2565 30.3530 1.1720 ;
      RECT 16.2680 0.2565 30.1820 1.3500 ;
      RECT 15.5210 0.2565 16.2500 1.1720 ;
      RECT 15.2870 0.4520 15.4850 1.3500 ;
      RECT 14.1080 0.3560 15.2600 1.1720 ;
      RECT 0.1760 0.2565 14.0900 1.3500 ;
      RECT 0.0050 0.2565 0.1580 1.1720 ;
      RECT 15.4670 0.2565 30.3530 1.0760 ;
      RECT 0.0050 0.3560 15.4490 1.0760 ;
      RECT 15.2420 0.2565 30.3530 0.4280 ;
      RECT 0.0050 0.2565 15.2240 1.0760 ;
      RECT 0.0050 0.2565 30.3530 0.3320 ;
      RECT 0.0050 2.3000 30.3530 2.4300 ;
      RECT 30.2360 1.3365 30.3530 2.4300 ;
      RECT 16.2140 2.2040 30.2180 2.4300 ;
      RECT 14.8820 2.2040 16.1960 2.4300 ;
      RECT 14.1620 1.3365 14.7920 2.4300 ;
      RECT 0.1400 2.2040 14.1440 2.4300 ;
      RECT 0.0050 1.3365 0.1220 2.4300 ;
      RECT 30.2000 1.3365 30.3530 2.2520 ;
      RECT 16.2680 1.3365 30.1820 2.4300 ;
      RECT 15.5210 1.3365 16.2500 2.2520 ;
      RECT 15.2870 1.5320 15.4850 2.4300 ;
      RECT 14.1080 1.4360 15.2600 2.2520 ;
      RECT 0.1760 1.3365 14.0900 2.4300 ;
      RECT 0.0050 1.3365 0.1580 2.2520 ;
      RECT 15.4670 1.3365 30.3530 2.1560 ;
      RECT 0.0050 1.4360 15.4490 2.1560 ;
      RECT 15.2420 1.3365 30.3530 1.5080 ;
      RECT 0.0050 1.3365 15.2240 2.1560 ;
      RECT 0.0050 1.3365 30.3530 1.4120 ;
      RECT 0.0050 3.3800 30.3530 3.5100 ;
      RECT 30.2360 2.4165 30.3530 3.5100 ;
      RECT 16.2140 3.2840 30.2180 3.5100 ;
      RECT 14.8820 3.2840 16.1960 3.5100 ;
      RECT 14.1620 2.4165 14.7920 3.5100 ;
      RECT 0.1400 3.2840 14.1440 3.5100 ;
      RECT 0.0050 2.4165 0.1220 3.5100 ;
      RECT 30.2000 2.4165 30.3530 3.3320 ;
      RECT 16.2680 2.4165 30.1820 3.5100 ;
      RECT 15.5210 2.4165 16.2500 3.3320 ;
      RECT 15.2870 2.6120 15.4850 3.5100 ;
      RECT 14.1080 2.5160 15.2600 3.3320 ;
      RECT 0.1760 2.4165 14.0900 3.5100 ;
      RECT 0.0050 2.4165 0.1580 3.3320 ;
      RECT 15.4670 2.4165 30.3530 3.2360 ;
      RECT 0.0050 2.5160 15.4490 3.2360 ;
      RECT 15.2420 2.4165 30.3530 2.5880 ;
      RECT 0.0050 2.4165 15.2240 3.2360 ;
      RECT 0.0050 2.4165 30.3530 2.4920 ;
      RECT 0.0050 4.4600 30.3530 4.5900 ;
      RECT 30.2360 3.4965 30.3530 4.5900 ;
      RECT 16.2140 4.3640 30.2180 4.5900 ;
      RECT 14.8820 4.3640 16.1960 4.5900 ;
      RECT 14.1620 3.4965 14.7920 4.5900 ;
      RECT 0.1400 4.3640 14.1440 4.5900 ;
      RECT 0.0050 3.4965 0.1220 4.5900 ;
      RECT 30.2000 3.4965 30.3530 4.4120 ;
      RECT 16.2680 3.4965 30.1820 4.5900 ;
      RECT 15.5210 3.4965 16.2500 4.4120 ;
      RECT 15.2870 3.6920 15.4850 4.5900 ;
      RECT 14.1080 3.5960 15.2600 4.4120 ;
      RECT 0.1760 3.4965 14.0900 4.5900 ;
      RECT 0.0050 3.4965 0.1580 4.4120 ;
      RECT 15.4670 3.4965 30.3530 4.3160 ;
      RECT 0.0050 3.5960 15.4490 4.3160 ;
      RECT 15.2420 3.4965 30.3530 3.6680 ;
      RECT 0.0050 3.4965 15.2240 4.3160 ;
      RECT 0.0050 3.4965 30.3530 3.5720 ;
      RECT 0.0050 5.5400 30.3530 5.6700 ;
      RECT 30.2360 4.5765 30.3530 5.6700 ;
      RECT 16.2140 5.4440 30.2180 5.6700 ;
      RECT 14.8820 5.4440 16.1960 5.6700 ;
      RECT 14.1620 4.5765 14.7920 5.6700 ;
      RECT 0.1400 5.4440 14.1440 5.6700 ;
      RECT 0.0050 4.5765 0.1220 5.6700 ;
      RECT 30.2000 4.5765 30.3530 5.4920 ;
      RECT 16.2680 4.5765 30.1820 5.6700 ;
      RECT 15.5210 4.5765 16.2500 5.4920 ;
      RECT 15.2870 4.7720 15.4850 5.6700 ;
      RECT 14.1080 4.6760 15.2600 5.4920 ;
      RECT 0.1760 4.5765 14.0900 5.6700 ;
      RECT 0.0050 4.5765 0.1580 5.4920 ;
      RECT 15.4670 4.5765 30.3530 5.3960 ;
      RECT 0.0050 4.6760 15.4490 5.3960 ;
      RECT 15.2420 4.5765 30.3530 4.7480 ;
      RECT 0.0050 4.5765 15.2240 5.3960 ;
      RECT 0.0050 4.5765 30.3530 4.6520 ;
      RECT 0.0050 6.6200 30.3530 6.7500 ;
      RECT 30.2360 5.6565 30.3530 6.7500 ;
      RECT 16.2140 6.5240 30.2180 6.7500 ;
      RECT 14.8820 6.5240 16.1960 6.7500 ;
      RECT 14.1620 5.6565 14.7920 6.7500 ;
      RECT 0.1400 6.5240 14.1440 6.7500 ;
      RECT 0.0050 5.6565 0.1220 6.7500 ;
      RECT 30.2000 5.6565 30.3530 6.5720 ;
      RECT 16.2680 5.6565 30.1820 6.7500 ;
      RECT 15.5210 5.6565 16.2500 6.5720 ;
      RECT 15.2870 5.8520 15.4850 6.7500 ;
      RECT 14.1080 5.7560 15.2600 6.5720 ;
      RECT 0.1760 5.6565 14.0900 6.7500 ;
      RECT 0.0050 5.6565 0.1580 6.5720 ;
      RECT 15.4670 5.6565 30.3530 6.4760 ;
      RECT 0.0050 5.7560 15.4490 6.4760 ;
      RECT 15.2420 5.6565 30.3530 5.8280 ;
      RECT 0.0050 5.6565 15.2240 6.4760 ;
      RECT 0.0050 5.6565 30.3530 5.7320 ;
      RECT 0.0050 7.7000 30.3530 7.8300 ;
      RECT 30.2360 6.7365 30.3530 7.8300 ;
      RECT 16.2140 7.6040 30.2180 7.8300 ;
      RECT 14.8820 7.6040 16.1960 7.8300 ;
      RECT 14.1620 6.7365 14.7920 7.8300 ;
      RECT 0.1400 7.6040 14.1440 7.8300 ;
      RECT 0.0050 6.7365 0.1220 7.8300 ;
      RECT 30.2000 6.7365 30.3530 7.6520 ;
      RECT 16.2680 6.7365 30.1820 7.8300 ;
      RECT 15.5210 6.7365 16.2500 7.6520 ;
      RECT 15.2870 6.9320 15.4850 7.8300 ;
      RECT 14.1080 6.8360 15.2600 7.6520 ;
      RECT 0.1760 6.7365 14.0900 7.8300 ;
      RECT 0.0050 6.7365 0.1580 7.6520 ;
      RECT 15.4670 6.7365 30.3530 7.5560 ;
      RECT 0.0050 6.8360 15.4490 7.5560 ;
      RECT 15.2420 6.7365 30.3530 6.9080 ;
      RECT 0.0050 6.7365 15.2240 7.5560 ;
      RECT 0.0050 6.7365 30.3530 6.8120 ;
      RECT 0.0050 8.7800 30.3530 8.9100 ;
      RECT 30.2360 7.8165 30.3530 8.9100 ;
      RECT 16.2140 8.6840 30.2180 8.9100 ;
      RECT 14.8820 8.6840 16.1960 8.9100 ;
      RECT 14.1620 7.8165 14.7920 8.9100 ;
      RECT 0.1400 8.6840 14.1440 8.9100 ;
      RECT 0.0050 7.8165 0.1220 8.9100 ;
      RECT 30.2000 7.8165 30.3530 8.7320 ;
      RECT 16.2680 7.8165 30.1820 8.9100 ;
      RECT 15.5210 7.8165 16.2500 8.7320 ;
      RECT 15.2870 8.0120 15.4850 8.9100 ;
      RECT 14.1080 7.9160 15.2600 8.7320 ;
      RECT 0.1760 7.8165 14.0900 8.9100 ;
      RECT 0.0050 7.8165 0.1580 8.7320 ;
      RECT 15.4670 7.8165 30.3530 8.6360 ;
      RECT 0.0050 7.9160 15.4490 8.6360 ;
      RECT 15.2420 7.8165 30.3530 7.9880 ;
      RECT 0.0050 7.8165 15.2240 8.6360 ;
      RECT 0.0050 7.8165 30.3530 7.8920 ;
      RECT 0.0050 9.8600 30.3530 9.9900 ;
      RECT 30.2360 8.8965 30.3530 9.9900 ;
      RECT 16.2140 9.7640 30.2180 9.9900 ;
      RECT 14.8820 9.7640 16.1960 9.9900 ;
      RECT 14.1620 8.8965 14.7920 9.9900 ;
      RECT 0.1400 9.7640 14.1440 9.9900 ;
      RECT 0.0050 8.8965 0.1220 9.9900 ;
      RECT 30.2000 8.8965 30.3530 9.8120 ;
      RECT 16.2680 8.8965 30.1820 9.9900 ;
      RECT 15.5210 8.8965 16.2500 9.8120 ;
      RECT 15.2870 9.0920 15.4850 9.9900 ;
      RECT 14.1080 8.9960 15.2600 9.8120 ;
      RECT 0.1760 8.8965 14.0900 9.9900 ;
      RECT 0.0050 8.8965 0.1580 9.8120 ;
      RECT 15.4670 8.8965 30.3530 9.7160 ;
      RECT 0.0050 8.9960 15.4490 9.7160 ;
      RECT 15.2420 8.8965 30.3530 9.0680 ;
      RECT 0.0050 8.8965 15.2240 9.7160 ;
      RECT 0.0050 8.8965 30.3530 8.9720 ;
      RECT 0.0050 10.9400 30.3530 11.0700 ;
      RECT 30.2360 9.9765 30.3530 11.0700 ;
      RECT 16.2140 10.8440 30.2180 11.0700 ;
      RECT 14.8820 10.8440 16.1960 11.0700 ;
      RECT 14.1620 9.9765 14.7920 11.0700 ;
      RECT 0.1400 10.8440 14.1440 11.0700 ;
      RECT 0.0050 9.9765 0.1220 11.0700 ;
      RECT 30.2000 9.9765 30.3530 10.8920 ;
      RECT 16.2680 9.9765 30.1820 11.0700 ;
      RECT 15.5210 9.9765 16.2500 10.8920 ;
      RECT 15.2870 10.1720 15.4850 11.0700 ;
      RECT 14.1080 10.0760 15.2600 10.8920 ;
      RECT 0.1760 9.9765 14.0900 11.0700 ;
      RECT 0.0050 9.9765 0.1580 10.8920 ;
      RECT 15.4670 9.9765 30.3530 10.7960 ;
      RECT 0.0050 10.0760 15.4490 10.7960 ;
      RECT 15.2420 9.9765 30.3530 10.1480 ;
      RECT 0.0050 9.9765 15.2240 10.7960 ;
      RECT 0.0050 9.9765 30.3530 10.0520 ;
      RECT 0.0050 12.0200 30.3530 12.1500 ;
      RECT 30.2360 11.0565 30.3530 12.1500 ;
      RECT 16.2140 11.9240 30.2180 12.1500 ;
      RECT 14.8820 11.9240 16.1960 12.1500 ;
      RECT 14.1620 11.0565 14.7920 12.1500 ;
      RECT 0.1400 11.9240 14.1440 12.1500 ;
      RECT 0.0050 11.0565 0.1220 12.1500 ;
      RECT 30.2000 11.0565 30.3530 11.9720 ;
      RECT 16.2680 11.0565 30.1820 12.1500 ;
      RECT 15.5210 11.0565 16.2500 11.9720 ;
      RECT 15.2870 11.2520 15.4850 12.1500 ;
      RECT 14.1080 11.1560 15.2600 11.9720 ;
      RECT 0.1760 11.0565 14.0900 12.1500 ;
      RECT 0.0050 11.0565 0.1580 11.9720 ;
      RECT 15.4670 11.0565 30.3530 11.8760 ;
      RECT 0.0050 11.1560 15.4490 11.8760 ;
      RECT 15.2420 11.0565 30.3530 11.2280 ;
      RECT 0.0050 11.0565 15.2240 11.8760 ;
      RECT 0.0050 11.0565 30.3530 11.1320 ;
      RECT 0.0050 13.1000 30.3530 13.2300 ;
      RECT 30.2360 12.1365 30.3530 13.2300 ;
      RECT 16.2140 13.0040 30.2180 13.2300 ;
      RECT 14.8820 13.0040 16.1960 13.2300 ;
      RECT 14.1620 12.1365 14.7920 13.2300 ;
      RECT 0.1400 13.0040 14.1440 13.2300 ;
      RECT 0.0050 12.1365 0.1220 13.2300 ;
      RECT 30.2000 12.1365 30.3530 13.0520 ;
      RECT 16.2680 12.1365 30.1820 13.2300 ;
      RECT 15.5210 12.1365 16.2500 13.0520 ;
      RECT 15.2870 12.3320 15.4850 13.2300 ;
      RECT 14.1080 12.2360 15.2600 13.0520 ;
      RECT 0.1760 12.1365 14.0900 13.2300 ;
      RECT 0.0050 12.1365 0.1580 13.0520 ;
      RECT 15.4670 12.1365 30.3530 12.9560 ;
      RECT 0.0050 12.2360 15.4490 12.9560 ;
      RECT 15.2420 12.1365 30.3530 12.3080 ;
      RECT 0.0050 12.1365 15.2240 12.9560 ;
      RECT 0.0050 12.1365 30.3530 12.2120 ;
      RECT 0.0050 14.1800 30.3530 14.3100 ;
      RECT 30.2360 13.2165 30.3530 14.3100 ;
      RECT 16.2140 14.0840 30.2180 14.3100 ;
      RECT 14.8820 14.0840 16.1960 14.3100 ;
      RECT 14.1620 13.2165 14.7920 14.3100 ;
      RECT 0.1400 14.0840 14.1440 14.3100 ;
      RECT 0.0050 13.2165 0.1220 14.3100 ;
      RECT 30.2000 13.2165 30.3530 14.1320 ;
      RECT 16.2680 13.2165 30.1820 14.3100 ;
      RECT 15.5210 13.2165 16.2500 14.1320 ;
      RECT 15.2870 13.4120 15.4850 14.3100 ;
      RECT 14.1080 13.3160 15.2600 14.1320 ;
      RECT 0.1760 13.2165 14.0900 14.3100 ;
      RECT 0.0050 13.2165 0.1580 14.1320 ;
      RECT 15.4670 13.2165 30.3530 14.0360 ;
      RECT 0.0050 13.3160 15.4490 14.0360 ;
      RECT 15.2420 13.2165 30.3530 13.3880 ;
      RECT 0.0050 13.2165 15.2240 14.0360 ;
      RECT 0.0050 13.2165 30.3530 13.2920 ;
      RECT 0.0050 15.2600 30.3530 15.3900 ;
      RECT 30.2360 14.2965 30.3530 15.3900 ;
      RECT 16.2140 15.1640 30.2180 15.3900 ;
      RECT 14.8820 15.1640 16.1960 15.3900 ;
      RECT 14.1620 14.2965 14.7920 15.3900 ;
      RECT 0.1400 15.1640 14.1440 15.3900 ;
      RECT 0.0050 14.2965 0.1220 15.3900 ;
      RECT 30.2000 14.2965 30.3530 15.2120 ;
      RECT 16.2680 14.2965 30.1820 15.3900 ;
      RECT 15.5210 14.2965 16.2500 15.2120 ;
      RECT 15.2870 14.4920 15.4850 15.3900 ;
      RECT 14.1080 14.3960 15.2600 15.2120 ;
      RECT 0.1760 14.2965 14.0900 15.3900 ;
      RECT 0.0050 14.2965 0.1580 15.2120 ;
      RECT 15.4670 14.2965 30.3530 15.1160 ;
      RECT 0.0050 14.3960 15.4490 15.1160 ;
      RECT 15.2420 14.2965 30.3530 14.4680 ;
      RECT 0.0050 14.2965 15.2240 15.1160 ;
      RECT 0.0050 14.2965 30.3530 14.3720 ;
      RECT 0.0050 16.3400 30.3530 16.4700 ;
      RECT 30.2360 15.3765 30.3530 16.4700 ;
      RECT 16.2140 16.2440 30.2180 16.4700 ;
      RECT 14.8820 16.2440 16.1960 16.4700 ;
      RECT 14.1620 15.3765 14.7920 16.4700 ;
      RECT 0.1400 16.2440 14.1440 16.4700 ;
      RECT 0.0050 15.3765 0.1220 16.4700 ;
      RECT 30.2000 15.3765 30.3530 16.2920 ;
      RECT 16.2680 15.3765 30.1820 16.4700 ;
      RECT 15.5210 15.3765 16.2500 16.2920 ;
      RECT 15.2870 15.5720 15.4850 16.4700 ;
      RECT 14.1080 15.4760 15.2600 16.2920 ;
      RECT 0.1760 15.3765 14.0900 16.4700 ;
      RECT 0.0050 15.3765 0.1580 16.2920 ;
      RECT 15.4670 15.3765 30.3530 16.1960 ;
      RECT 0.0050 15.4760 15.4490 16.1960 ;
      RECT 15.2420 15.3765 30.3530 15.5480 ;
      RECT 0.0050 15.3765 15.2240 16.1960 ;
      RECT 0.0050 15.3765 30.3530 15.4520 ;
      RECT 0.0050 17.4200 30.3530 17.5500 ;
      RECT 30.2360 16.4565 30.3530 17.5500 ;
      RECT 16.2140 17.3240 30.2180 17.5500 ;
      RECT 14.8820 17.3240 16.1960 17.5500 ;
      RECT 14.1620 16.4565 14.7920 17.5500 ;
      RECT 0.1400 17.3240 14.1440 17.5500 ;
      RECT 0.0050 16.4565 0.1220 17.5500 ;
      RECT 30.2000 16.4565 30.3530 17.3720 ;
      RECT 16.2680 16.4565 30.1820 17.5500 ;
      RECT 15.5210 16.4565 16.2500 17.3720 ;
      RECT 15.2870 16.6520 15.4850 17.5500 ;
      RECT 14.1080 16.5560 15.2600 17.3720 ;
      RECT 0.1760 16.4565 14.0900 17.5500 ;
      RECT 0.0050 16.4565 0.1580 17.3720 ;
      RECT 15.4670 16.4565 30.3530 17.2760 ;
      RECT 0.0050 16.5560 15.4490 17.2760 ;
      RECT 15.2420 16.4565 30.3530 16.6280 ;
      RECT 0.0050 16.4565 15.2240 17.2760 ;
      RECT 0.0050 16.4565 30.3530 16.5320 ;
      RECT 0.0050 18.5000 30.3530 18.6300 ;
      RECT 30.2360 17.5365 30.3530 18.6300 ;
      RECT 16.2140 18.4040 30.2180 18.6300 ;
      RECT 14.8820 18.4040 16.1960 18.6300 ;
      RECT 14.1620 17.5365 14.7920 18.6300 ;
      RECT 0.1400 18.4040 14.1440 18.6300 ;
      RECT 0.0050 17.5365 0.1220 18.6300 ;
      RECT 30.2000 17.5365 30.3530 18.4520 ;
      RECT 16.2680 17.5365 30.1820 18.6300 ;
      RECT 15.5210 17.5365 16.2500 18.4520 ;
      RECT 15.2870 17.7320 15.4850 18.6300 ;
      RECT 14.1080 17.6360 15.2600 18.4520 ;
      RECT 0.1760 17.5365 14.0900 18.6300 ;
      RECT 0.0050 17.5365 0.1580 18.4520 ;
      RECT 15.4670 17.5365 30.3530 18.3560 ;
      RECT 0.0050 17.6360 15.4490 18.3560 ;
      RECT 15.2420 17.5365 30.3530 17.7080 ;
      RECT 0.0050 17.5365 15.2240 18.3560 ;
      RECT 0.0050 17.5365 30.3530 17.6120 ;
      RECT 0.0050 19.5800 30.3530 19.7100 ;
      RECT 30.2360 18.6165 30.3530 19.7100 ;
      RECT 16.2140 19.4840 30.2180 19.7100 ;
      RECT 14.8820 19.4840 16.1960 19.7100 ;
      RECT 14.1620 18.6165 14.7920 19.7100 ;
      RECT 0.1400 19.4840 14.1440 19.7100 ;
      RECT 0.0050 18.6165 0.1220 19.7100 ;
      RECT 30.2000 18.6165 30.3530 19.5320 ;
      RECT 16.2680 18.6165 30.1820 19.7100 ;
      RECT 15.5210 18.6165 16.2500 19.5320 ;
      RECT 15.2870 18.8120 15.4850 19.7100 ;
      RECT 14.1080 18.7160 15.2600 19.5320 ;
      RECT 0.1760 18.6165 14.0900 19.7100 ;
      RECT 0.0050 18.6165 0.1580 19.5320 ;
      RECT 15.4670 18.6165 30.3530 19.4360 ;
      RECT 0.0050 18.7160 15.4490 19.4360 ;
      RECT 15.2420 18.6165 30.3530 18.7880 ;
      RECT 0.0050 18.6165 15.2240 19.4360 ;
      RECT 0.0050 18.6165 30.3530 18.6920 ;
      RECT 0.0050 20.6600 30.3530 20.7900 ;
      RECT 30.2360 19.6965 30.3530 20.7900 ;
      RECT 16.2140 20.5640 30.2180 20.7900 ;
      RECT 14.8820 20.5640 16.1960 20.7900 ;
      RECT 14.1620 19.6965 14.7920 20.7900 ;
      RECT 0.1400 20.5640 14.1440 20.7900 ;
      RECT 0.0050 19.6965 0.1220 20.7900 ;
      RECT 30.2000 19.6965 30.3530 20.6120 ;
      RECT 16.2680 19.6965 30.1820 20.7900 ;
      RECT 15.5210 19.6965 16.2500 20.6120 ;
      RECT 15.2870 19.8920 15.4850 20.7900 ;
      RECT 14.1080 19.7960 15.2600 20.6120 ;
      RECT 0.1760 19.6965 14.0900 20.7900 ;
      RECT 0.0050 19.6965 0.1580 20.6120 ;
      RECT 15.4670 19.6965 30.3530 20.5160 ;
      RECT 0.0050 19.7960 15.4490 20.5160 ;
      RECT 15.2420 19.6965 30.3530 19.8680 ;
      RECT 0.0050 19.6965 15.2240 20.5160 ;
      RECT 0.0050 19.6965 30.3530 19.7720 ;
      RECT 0.0050 21.7400 30.3530 21.8700 ;
      RECT 30.2360 20.7765 30.3530 21.8700 ;
      RECT 16.2140 21.6440 30.2180 21.8700 ;
      RECT 14.8820 21.6440 16.1960 21.8700 ;
      RECT 14.1620 20.7765 14.7920 21.8700 ;
      RECT 0.1400 21.6440 14.1440 21.8700 ;
      RECT 0.0050 20.7765 0.1220 21.8700 ;
      RECT 30.2000 20.7765 30.3530 21.6920 ;
      RECT 16.2680 20.7765 30.1820 21.8700 ;
      RECT 15.5210 20.7765 16.2500 21.6920 ;
      RECT 15.2870 20.9720 15.4850 21.8700 ;
      RECT 14.1080 20.8760 15.2600 21.6920 ;
      RECT 0.1760 20.7765 14.0900 21.8700 ;
      RECT 0.0050 20.7765 0.1580 21.6920 ;
      RECT 15.4670 20.7765 30.3530 21.5960 ;
      RECT 0.0050 20.8760 15.4490 21.5960 ;
      RECT 15.2420 20.7765 30.3530 20.9480 ;
      RECT 0.0050 20.7765 15.2240 21.5960 ;
      RECT 0.0050 20.7765 30.3530 20.8520 ;
      RECT 0.0050 22.8200 30.3530 22.9500 ;
      RECT 30.2360 21.8565 30.3530 22.9500 ;
      RECT 16.2140 22.7240 30.2180 22.9500 ;
      RECT 14.8820 22.7240 16.1960 22.9500 ;
      RECT 14.1620 21.8565 14.7920 22.9500 ;
      RECT 0.1400 22.7240 14.1440 22.9500 ;
      RECT 0.0050 21.8565 0.1220 22.9500 ;
      RECT 30.2000 21.8565 30.3530 22.7720 ;
      RECT 16.2680 21.8565 30.1820 22.9500 ;
      RECT 15.5210 21.8565 16.2500 22.7720 ;
      RECT 15.2870 22.0520 15.4850 22.9500 ;
      RECT 14.1080 21.9560 15.2600 22.7720 ;
      RECT 0.1760 21.8565 14.0900 22.9500 ;
      RECT 0.0050 21.8565 0.1580 22.7720 ;
      RECT 15.4670 21.8565 30.3530 22.6760 ;
      RECT 0.0050 21.9560 15.4490 22.6760 ;
      RECT 15.2420 21.8565 30.3530 22.0280 ;
      RECT 0.0050 21.8565 15.2240 22.6760 ;
      RECT 0.0050 21.8565 30.3530 21.9320 ;
      RECT 0.0050 23.9000 30.3530 24.0300 ;
      RECT 30.2360 22.9365 30.3530 24.0300 ;
      RECT 16.2140 23.8040 30.2180 24.0300 ;
      RECT 14.8820 23.8040 16.1960 24.0300 ;
      RECT 14.1620 22.9365 14.7920 24.0300 ;
      RECT 0.1400 23.8040 14.1440 24.0300 ;
      RECT 0.0050 22.9365 0.1220 24.0300 ;
      RECT 30.2000 22.9365 30.3530 23.8520 ;
      RECT 16.2680 22.9365 30.1820 24.0300 ;
      RECT 15.5210 22.9365 16.2500 23.8520 ;
      RECT 15.2870 23.1320 15.4850 24.0300 ;
      RECT 14.1080 23.0360 15.2600 23.8520 ;
      RECT 0.1760 22.9365 14.0900 24.0300 ;
      RECT 0.0050 22.9365 0.1580 23.8520 ;
      RECT 15.4670 22.9365 30.3530 23.7560 ;
      RECT 0.0050 23.0360 15.4490 23.7560 ;
      RECT 15.2420 22.9365 30.3530 23.1080 ;
      RECT 0.0050 22.9365 15.2240 23.7560 ;
      RECT 0.0050 22.9365 30.3530 23.0120 ;
      RECT 0.0050 24.9800 30.3530 25.1100 ;
      RECT 30.2360 24.0165 30.3530 25.1100 ;
      RECT 16.2140 24.8840 30.2180 25.1100 ;
      RECT 14.8820 24.8840 16.1960 25.1100 ;
      RECT 14.1620 24.0165 14.7920 25.1100 ;
      RECT 0.1400 24.8840 14.1440 25.1100 ;
      RECT 0.0050 24.0165 0.1220 25.1100 ;
      RECT 30.2000 24.0165 30.3530 24.9320 ;
      RECT 16.2680 24.0165 30.1820 25.1100 ;
      RECT 15.5210 24.0165 16.2500 24.9320 ;
      RECT 15.2870 24.2120 15.4850 25.1100 ;
      RECT 14.1080 24.1160 15.2600 24.9320 ;
      RECT 0.1760 24.0165 14.0900 25.1100 ;
      RECT 0.0050 24.0165 0.1580 24.9320 ;
      RECT 15.4670 24.0165 30.3530 24.8360 ;
      RECT 0.0050 24.1160 15.4490 24.8360 ;
      RECT 15.2420 24.0165 30.3530 24.1880 ;
      RECT 0.0050 24.0165 15.2240 24.8360 ;
      RECT 0.0050 24.0165 30.3530 24.0920 ;
      RECT 0.0050 26.0600 30.3530 26.1900 ;
      RECT 30.2360 25.0965 30.3530 26.1900 ;
      RECT 16.2140 25.9640 30.2180 26.1900 ;
      RECT 14.8820 25.9640 16.1960 26.1900 ;
      RECT 14.1620 25.0965 14.7920 26.1900 ;
      RECT 0.1400 25.9640 14.1440 26.1900 ;
      RECT 0.0050 25.0965 0.1220 26.1900 ;
      RECT 30.2000 25.0965 30.3530 26.0120 ;
      RECT 16.2680 25.0965 30.1820 26.1900 ;
      RECT 15.5210 25.0965 16.2500 26.0120 ;
      RECT 15.2870 25.2920 15.4850 26.1900 ;
      RECT 14.1080 25.1960 15.2600 26.0120 ;
      RECT 0.1760 25.0965 14.0900 26.1900 ;
      RECT 0.0050 25.0965 0.1580 26.0120 ;
      RECT 15.4670 25.0965 30.3530 25.9160 ;
      RECT 0.0050 25.1960 15.4490 25.9160 ;
      RECT 15.2420 25.0965 30.3530 25.2680 ;
      RECT 0.0050 25.0965 15.2240 25.9160 ;
      RECT 0.0050 25.0965 30.3530 25.1720 ;
      RECT 0.0050 27.1400 30.3530 27.2700 ;
      RECT 30.2360 26.1765 30.3530 27.2700 ;
      RECT 16.2140 27.0440 30.2180 27.2700 ;
      RECT 14.8820 27.0440 16.1960 27.2700 ;
      RECT 14.1620 26.1765 14.7920 27.2700 ;
      RECT 0.1400 27.0440 14.1440 27.2700 ;
      RECT 0.0050 26.1765 0.1220 27.2700 ;
      RECT 30.2000 26.1765 30.3530 27.0920 ;
      RECT 16.2680 26.1765 30.1820 27.2700 ;
      RECT 15.5210 26.1765 16.2500 27.0920 ;
      RECT 15.2870 26.3720 15.4850 27.2700 ;
      RECT 14.1080 26.2760 15.2600 27.0920 ;
      RECT 0.1760 26.1765 14.0900 27.2700 ;
      RECT 0.0050 26.1765 0.1580 27.0920 ;
      RECT 15.4670 26.1765 30.3530 26.9960 ;
      RECT 0.0050 26.2760 15.4490 26.9960 ;
      RECT 15.2420 26.1765 30.3530 26.3480 ;
      RECT 0.0050 26.1765 15.2240 26.9960 ;
      RECT 0.0050 26.1765 30.3530 26.2520 ;
      RECT 0.0050 28.2200 30.3530 28.3500 ;
      RECT 30.2360 27.2565 30.3530 28.3500 ;
      RECT 16.2140 28.1240 30.2180 28.3500 ;
      RECT 14.8820 28.1240 16.1960 28.3500 ;
      RECT 14.1620 27.2565 14.7920 28.3500 ;
      RECT 0.1400 28.1240 14.1440 28.3500 ;
      RECT 0.0050 27.2565 0.1220 28.3500 ;
      RECT 30.2000 27.2565 30.3530 28.1720 ;
      RECT 16.2680 27.2565 30.1820 28.3500 ;
      RECT 15.5210 27.2565 16.2500 28.1720 ;
      RECT 15.2870 27.4520 15.4850 28.3500 ;
      RECT 14.1080 27.3560 15.2600 28.1720 ;
      RECT 0.1760 27.2565 14.0900 28.3500 ;
      RECT 0.0050 27.2565 0.1580 28.1720 ;
      RECT 15.4670 27.2565 30.3530 28.0760 ;
      RECT 0.0050 27.3560 15.4490 28.0760 ;
      RECT 15.2420 27.2565 30.3530 27.4280 ;
      RECT 0.0050 27.2565 15.2240 28.0760 ;
      RECT 0.0050 27.2565 30.3530 27.3320 ;
      RECT 0.0050 29.3000 30.3530 29.4300 ;
      RECT 30.2360 28.3365 30.3530 29.4300 ;
      RECT 16.2140 29.2040 30.2180 29.4300 ;
      RECT 14.8820 29.2040 16.1960 29.4300 ;
      RECT 14.1620 28.3365 14.7920 29.4300 ;
      RECT 0.1400 29.2040 14.1440 29.4300 ;
      RECT 0.0050 28.3365 0.1220 29.4300 ;
      RECT 30.2000 28.3365 30.3530 29.2520 ;
      RECT 16.2680 28.3365 30.1820 29.4300 ;
      RECT 15.5210 28.3365 16.2500 29.2520 ;
      RECT 15.2870 28.5320 15.4850 29.4300 ;
      RECT 14.1080 28.4360 15.2600 29.2520 ;
      RECT 0.1760 28.3365 14.0900 29.4300 ;
      RECT 0.0050 28.3365 0.1580 29.2520 ;
      RECT 15.4670 28.3365 30.3530 29.1560 ;
      RECT 0.0050 28.4360 15.4490 29.1560 ;
      RECT 15.2420 28.3365 30.3530 28.5080 ;
      RECT 0.0050 28.3365 15.2240 29.1560 ;
      RECT 0.0050 28.3365 30.3530 28.4120 ;
      RECT 0.0050 30.3800 30.3530 30.5100 ;
      RECT 30.2360 29.4165 30.3530 30.5100 ;
      RECT 16.2140 30.2840 30.2180 30.5100 ;
      RECT 14.8820 30.2840 16.1960 30.5100 ;
      RECT 14.1620 29.4165 14.7920 30.5100 ;
      RECT 0.1400 30.2840 14.1440 30.5100 ;
      RECT 0.0050 29.4165 0.1220 30.5100 ;
      RECT 30.2000 29.4165 30.3530 30.3320 ;
      RECT 16.2680 29.4165 30.1820 30.5100 ;
      RECT 15.5210 29.4165 16.2500 30.3320 ;
      RECT 15.2870 29.6120 15.4850 30.5100 ;
      RECT 14.1080 29.5160 15.2600 30.3320 ;
      RECT 0.1760 29.4165 14.0900 30.5100 ;
      RECT 0.0050 29.4165 0.1580 30.3320 ;
      RECT 15.4670 29.4165 30.3530 30.2360 ;
      RECT 0.0050 29.5160 15.4490 30.2360 ;
      RECT 15.2420 29.4165 30.3530 29.5880 ;
      RECT 0.0050 29.4165 15.2240 30.2360 ;
      RECT 0.0050 29.4165 30.3530 29.4920 ;
      RECT 0.0050 31.4600 30.3530 31.5900 ;
      RECT 30.2360 30.4965 30.3530 31.5900 ;
      RECT 16.2140 31.3640 30.2180 31.5900 ;
      RECT 14.8820 31.3640 16.1960 31.5900 ;
      RECT 14.1620 30.4965 14.7920 31.5900 ;
      RECT 0.1400 31.3640 14.1440 31.5900 ;
      RECT 0.0050 30.4965 0.1220 31.5900 ;
      RECT 30.2000 30.4965 30.3530 31.4120 ;
      RECT 16.2680 30.4965 30.1820 31.5900 ;
      RECT 15.5210 30.4965 16.2500 31.4120 ;
      RECT 15.2870 30.6920 15.4850 31.5900 ;
      RECT 14.1080 30.5960 15.2600 31.4120 ;
      RECT 0.1760 30.4965 14.0900 31.5900 ;
      RECT 0.0050 30.4965 0.1580 31.4120 ;
      RECT 15.4670 30.4965 30.3530 31.3160 ;
      RECT 0.0050 30.5960 15.4490 31.3160 ;
      RECT 15.2420 30.4965 30.3530 30.6680 ;
      RECT 0.0050 30.4965 15.2240 31.3160 ;
      RECT 0.0050 30.4965 30.3530 30.5720 ;
      RECT 0.0050 32.5400 30.3530 32.6700 ;
      RECT 30.2360 31.5765 30.3530 32.6700 ;
      RECT 16.2140 32.4440 30.2180 32.6700 ;
      RECT 14.8820 32.4440 16.1960 32.6700 ;
      RECT 14.1620 31.5765 14.7920 32.6700 ;
      RECT 0.1400 32.4440 14.1440 32.6700 ;
      RECT 0.0050 31.5765 0.1220 32.6700 ;
      RECT 30.2000 31.5765 30.3530 32.4920 ;
      RECT 16.2680 31.5765 30.1820 32.6700 ;
      RECT 15.5210 31.5765 16.2500 32.4920 ;
      RECT 15.2870 31.7720 15.4850 32.6700 ;
      RECT 14.1080 31.6760 15.2600 32.4920 ;
      RECT 0.1760 31.5765 14.0900 32.6700 ;
      RECT 0.0050 31.5765 0.1580 32.4920 ;
      RECT 15.4670 31.5765 30.3530 32.3960 ;
      RECT 0.0050 31.6760 15.4490 32.3960 ;
      RECT 15.2420 31.5765 30.3530 31.7480 ;
      RECT 0.0050 31.5765 15.2240 32.3960 ;
      RECT 0.0050 31.5765 30.3530 31.6520 ;
      RECT 0.0050 33.6200 30.3530 33.7500 ;
      RECT 30.2360 32.6565 30.3530 33.7500 ;
      RECT 16.2140 33.5240 30.2180 33.7500 ;
      RECT 14.8820 33.5240 16.1960 33.7500 ;
      RECT 14.1620 32.6565 14.7920 33.7500 ;
      RECT 0.1400 33.5240 14.1440 33.7500 ;
      RECT 0.0050 32.6565 0.1220 33.7500 ;
      RECT 30.2000 32.6565 30.3530 33.5720 ;
      RECT 16.2680 32.6565 30.1820 33.7500 ;
      RECT 15.5210 32.6565 16.2500 33.5720 ;
      RECT 15.2870 32.8520 15.4850 33.7500 ;
      RECT 14.1080 32.7560 15.2600 33.5720 ;
      RECT 0.1760 32.6565 14.0900 33.7500 ;
      RECT 0.0050 32.6565 0.1580 33.5720 ;
      RECT 15.4670 32.6565 30.3530 33.4760 ;
      RECT 0.0050 32.7560 15.4490 33.4760 ;
      RECT 15.2420 32.6565 30.3530 32.8280 ;
      RECT 0.0050 32.6565 15.2240 33.4760 ;
      RECT 0.0050 32.6565 30.3530 32.7320 ;
      RECT 0.0050 34.7000 30.3530 34.8300 ;
      RECT 30.2360 33.7365 30.3530 34.8300 ;
      RECT 16.2140 34.6040 30.2180 34.8300 ;
      RECT 14.8820 34.6040 16.1960 34.8300 ;
      RECT 14.1620 33.7365 14.7920 34.8300 ;
      RECT 0.1400 34.6040 14.1440 34.8300 ;
      RECT 0.0050 33.7365 0.1220 34.8300 ;
      RECT 30.2000 33.7365 30.3530 34.6520 ;
      RECT 16.2680 33.7365 30.1820 34.8300 ;
      RECT 15.5210 33.7365 16.2500 34.6520 ;
      RECT 15.2870 33.9320 15.4850 34.8300 ;
      RECT 14.1080 33.8360 15.2600 34.6520 ;
      RECT 0.1760 33.7365 14.0900 34.8300 ;
      RECT 0.0050 33.7365 0.1580 34.6520 ;
      RECT 15.4670 33.7365 30.3530 34.5560 ;
      RECT 0.0050 33.8360 15.4490 34.5560 ;
      RECT 15.2420 33.7365 30.3530 33.9080 ;
      RECT 0.0050 33.7365 15.2240 34.5560 ;
      RECT 0.0050 33.7365 30.3530 33.8120 ;
      RECT 0.0000 42.1735 30.3480 43.5070 ;
      RECT 17.7210 34.8535 30.3480 43.5070 ;
      RECT 15.5210 36.3175 30.3480 43.5070 ;
      RECT 16.4250 36.1255 30.3480 43.5070 ;
      RECT 15.4690 34.8535 15.5030 43.5070 ;
      RECT 15.4170 34.8535 15.4510 43.5070 ;
      RECT 15.3650 34.8535 15.3990 43.5070 ;
      RECT 15.3130 34.8535 15.3470 43.5070 ;
      RECT 0.0000 36.4135 15.2950 43.5070 ;
      RECT 0.0000 39.0055 30.3480 41.9575 ;
      RECT 14.1570 35.8375 15.8310 38.7895 ;
      RECT 0.0000 36.1255 14.1390 43.5070 ;
      RECT 0.0000 36.2215 16.4070 36.3895 ;
      RECT 16.2090 36.1255 30.3480 36.2935 ;
      RECT 0.0000 36.1255 16.1910 36.3895 ;
      RECT 17.5050 34.8535 17.7030 43.5070 ;
      RECT 13.7250 35.9335 17.4870 36.1975 ;
      RECT 12.8610 35.5495 13.7070 43.5070 ;
      RECT 0.0000 34.8535 12.8430 43.5070 ;
      RECT 17.2890 34.8535 30.3480 36.1015 ;
      RECT 17.0730 35.5495 30.3480 36.1015 ;
      RECT 15.8490 35.8375 17.0550 36.1975 ;
      RECT 0.0000 35.8375 15.8310 36.1015 ;
      RECT 16.8570 34.8535 17.2710 35.9095 ;
      RECT 16.2630 35.5495 30.3480 35.9095 ;
      RECT 15.5210 35.5495 16.2450 35.9095 ;
      RECT 14.1030 35.5495 15.2950 36.3895 ;
      RECT 0.0000 35.5495 14.0850 36.1015 ;
      RECT 15.5610 35.5015 16.8390 35.6215 ;
      RECT 14.3730 35.5015 15.5430 35.6215 ;
      RECT 13.5090 35.5015 14.3550 35.6215 ;
      RECT 13.0770 35.5015 13.4910 43.5070 ;
      RECT 0.0000 34.8535 13.0590 36.1015 ;
      RECT 16.6410 34.8535 30.3480 35.5255 ;
      RECT 15.1650 34.8535 16.6230 35.5255 ;
      RECT 14.1930 34.8535 15.1470 35.5255 ;
      RECT 13.2930 34.8535 14.1750 35.5255 ;
      RECT 0.0000 34.8535 13.2750 35.5255 ;
      RECT 0.0000 34.8535 30.3480 35.4775 ;
        RECT 0.0050 43.9070 30.3530 44.0370 ;
        RECT 30.2360 42.9435 30.3530 44.0370 ;
        RECT 16.2140 43.8110 30.2180 44.0370 ;
        RECT 14.8820 43.8110 16.1960 44.0370 ;
        RECT 14.1620 42.9435 14.7920 44.0370 ;
        RECT 0.1400 43.8110 14.1440 44.0370 ;
        RECT 0.0050 42.9435 0.1220 44.0370 ;
        RECT 30.2000 42.9435 30.3530 43.8590 ;
        RECT 16.2680 42.9435 30.1820 44.0370 ;
        RECT 15.5210 42.9435 16.2500 43.8590 ;
        RECT 15.2870 43.1390 15.4850 44.0370 ;
        RECT 14.1080 43.0430 15.2600 43.8590 ;
        RECT 0.1760 42.9435 14.0900 44.0370 ;
        RECT 0.0050 42.9435 0.1580 43.8590 ;
        RECT 15.4670 42.9435 30.3530 43.7630 ;
        RECT 0.0050 43.0430 15.4490 43.7630 ;
        RECT 15.2420 42.9435 30.3530 43.1150 ;
        RECT 0.0050 42.9435 15.2240 43.7630 ;
        RECT 0.0050 42.9435 30.3530 43.0190 ;
        RECT 0.0050 44.9870 30.3530 45.1170 ;
        RECT 30.2360 44.0235 30.3530 45.1170 ;
        RECT 16.2140 44.8910 30.2180 45.1170 ;
        RECT 14.8820 44.8910 16.1960 45.1170 ;
        RECT 14.1620 44.0235 14.7920 45.1170 ;
        RECT 0.1400 44.8910 14.1440 45.1170 ;
        RECT 0.0050 44.0235 0.1220 45.1170 ;
        RECT 30.2000 44.0235 30.3530 44.9390 ;
        RECT 16.2680 44.0235 30.1820 45.1170 ;
        RECT 15.5210 44.0235 16.2500 44.9390 ;
        RECT 15.2870 44.2190 15.4850 45.1170 ;
        RECT 14.1080 44.1230 15.2600 44.9390 ;
        RECT 0.1760 44.0235 14.0900 45.1170 ;
        RECT 0.0050 44.0235 0.1580 44.9390 ;
        RECT 15.4670 44.0235 30.3530 44.8430 ;
        RECT 0.0050 44.1230 15.4490 44.8430 ;
        RECT 15.2420 44.0235 30.3530 44.1950 ;
        RECT 0.0050 44.0235 15.2240 44.8430 ;
        RECT 0.0050 44.0235 30.3530 44.0990 ;
        RECT 0.0050 46.0670 30.3530 46.1970 ;
        RECT 30.2360 45.1035 30.3530 46.1970 ;
        RECT 16.2140 45.9710 30.2180 46.1970 ;
        RECT 14.8820 45.9710 16.1960 46.1970 ;
        RECT 14.1620 45.1035 14.7920 46.1970 ;
        RECT 0.1400 45.9710 14.1440 46.1970 ;
        RECT 0.0050 45.1035 0.1220 46.1970 ;
        RECT 30.2000 45.1035 30.3530 46.0190 ;
        RECT 16.2680 45.1035 30.1820 46.1970 ;
        RECT 15.5210 45.1035 16.2500 46.0190 ;
        RECT 15.2870 45.2990 15.4850 46.1970 ;
        RECT 14.1080 45.2030 15.2600 46.0190 ;
        RECT 0.1760 45.1035 14.0900 46.1970 ;
        RECT 0.0050 45.1035 0.1580 46.0190 ;
        RECT 15.4670 45.1035 30.3530 45.9230 ;
        RECT 0.0050 45.2030 15.4490 45.9230 ;
        RECT 15.2420 45.1035 30.3530 45.2750 ;
        RECT 0.0050 45.1035 15.2240 45.9230 ;
        RECT 0.0050 45.1035 30.3530 45.1790 ;
        RECT 0.0050 47.1470 30.3530 47.2770 ;
        RECT 30.2360 46.1835 30.3530 47.2770 ;
        RECT 16.2140 47.0510 30.2180 47.2770 ;
        RECT 14.8820 47.0510 16.1960 47.2770 ;
        RECT 14.1620 46.1835 14.7920 47.2770 ;
        RECT 0.1400 47.0510 14.1440 47.2770 ;
        RECT 0.0050 46.1835 0.1220 47.2770 ;
        RECT 30.2000 46.1835 30.3530 47.0990 ;
        RECT 16.2680 46.1835 30.1820 47.2770 ;
        RECT 15.5210 46.1835 16.2500 47.0990 ;
        RECT 15.2870 46.3790 15.4850 47.2770 ;
        RECT 14.1080 46.2830 15.2600 47.0990 ;
        RECT 0.1760 46.1835 14.0900 47.2770 ;
        RECT 0.0050 46.1835 0.1580 47.0990 ;
        RECT 15.4670 46.1835 30.3530 47.0030 ;
        RECT 0.0050 46.2830 15.4490 47.0030 ;
        RECT 15.2420 46.1835 30.3530 46.3550 ;
        RECT 0.0050 46.1835 15.2240 47.0030 ;
        RECT 0.0050 46.1835 30.3530 46.2590 ;
        RECT 0.0050 48.2270 30.3530 48.3570 ;
        RECT 30.2360 47.2635 30.3530 48.3570 ;
        RECT 16.2140 48.1310 30.2180 48.3570 ;
        RECT 14.8820 48.1310 16.1960 48.3570 ;
        RECT 14.1620 47.2635 14.7920 48.3570 ;
        RECT 0.1400 48.1310 14.1440 48.3570 ;
        RECT 0.0050 47.2635 0.1220 48.3570 ;
        RECT 30.2000 47.2635 30.3530 48.1790 ;
        RECT 16.2680 47.2635 30.1820 48.3570 ;
        RECT 15.5210 47.2635 16.2500 48.1790 ;
        RECT 15.2870 47.4590 15.4850 48.3570 ;
        RECT 14.1080 47.3630 15.2600 48.1790 ;
        RECT 0.1760 47.2635 14.0900 48.3570 ;
        RECT 0.0050 47.2635 0.1580 48.1790 ;
        RECT 15.4670 47.2635 30.3530 48.0830 ;
        RECT 0.0050 47.3630 15.4490 48.0830 ;
        RECT 15.2420 47.2635 30.3530 47.4350 ;
        RECT 0.0050 47.2635 15.2240 48.0830 ;
        RECT 0.0050 47.2635 30.3530 47.3390 ;
        RECT 0.0050 49.3070 30.3530 49.4370 ;
        RECT 30.2360 48.3435 30.3530 49.4370 ;
        RECT 16.2140 49.2110 30.2180 49.4370 ;
        RECT 14.8820 49.2110 16.1960 49.4370 ;
        RECT 14.1620 48.3435 14.7920 49.4370 ;
        RECT 0.1400 49.2110 14.1440 49.4370 ;
        RECT 0.0050 48.3435 0.1220 49.4370 ;
        RECT 30.2000 48.3435 30.3530 49.2590 ;
        RECT 16.2680 48.3435 30.1820 49.4370 ;
        RECT 15.5210 48.3435 16.2500 49.2590 ;
        RECT 15.2870 48.5390 15.4850 49.4370 ;
        RECT 14.1080 48.4430 15.2600 49.2590 ;
        RECT 0.1760 48.3435 14.0900 49.4370 ;
        RECT 0.0050 48.3435 0.1580 49.2590 ;
        RECT 15.4670 48.3435 30.3530 49.1630 ;
        RECT 0.0050 48.4430 15.4490 49.1630 ;
        RECT 15.2420 48.3435 30.3530 48.5150 ;
        RECT 0.0050 48.3435 15.2240 49.1630 ;
        RECT 0.0050 48.3435 30.3530 48.4190 ;
        RECT 0.0050 50.3870 30.3530 50.5170 ;
        RECT 30.2360 49.4235 30.3530 50.5170 ;
        RECT 16.2140 50.2910 30.2180 50.5170 ;
        RECT 14.8820 50.2910 16.1960 50.5170 ;
        RECT 14.1620 49.4235 14.7920 50.5170 ;
        RECT 0.1400 50.2910 14.1440 50.5170 ;
        RECT 0.0050 49.4235 0.1220 50.5170 ;
        RECT 30.2000 49.4235 30.3530 50.3390 ;
        RECT 16.2680 49.4235 30.1820 50.5170 ;
        RECT 15.5210 49.4235 16.2500 50.3390 ;
        RECT 15.2870 49.6190 15.4850 50.5170 ;
        RECT 14.1080 49.5230 15.2600 50.3390 ;
        RECT 0.1760 49.4235 14.0900 50.5170 ;
        RECT 0.0050 49.4235 0.1580 50.3390 ;
        RECT 15.4670 49.4235 30.3530 50.2430 ;
        RECT 0.0050 49.5230 15.4490 50.2430 ;
        RECT 15.2420 49.4235 30.3530 49.5950 ;
        RECT 0.0050 49.4235 15.2240 50.2430 ;
        RECT 0.0050 49.4235 30.3530 49.4990 ;
        RECT 0.0050 51.4670 30.3530 51.5970 ;
        RECT 30.2360 50.5035 30.3530 51.5970 ;
        RECT 16.2140 51.3710 30.2180 51.5970 ;
        RECT 14.8820 51.3710 16.1960 51.5970 ;
        RECT 14.1620 50.5035 14.7920 51.5970 ;
        RECT 0.1400 51.3710 14.1440 51.5970 ;
        RECT 0.0050 50.5035 0.1220 51.5970 ;
        RECT 30.2000 50.5035 30.3530 51.4190 ;
        RECT 16.2680 50.5035 30.1820 51.5970 ;
        RECT 15.5210 50.5035 16.2500 51.4190 ;
        RECT 15.2870 50.6990 15.4850 51.5970 ;
        RECT 14.1080 50.6030 15.2600 51.4190 ;
        RECT 0.1760 50.5035 14.0900 51.5970 ;
        RECT 0.0050 50.5035 0.1580 51.4190 ;
        RECT 15.4670 50.5035 30.3530 51.3230 ;
        RECT 0.0050 50.6030 15.4490 51.3230 ;
        RECT 15.2420 50.5035 30.3530 50.6750 ;
        RECT 0.0050 50.5035 15.2240 51.3230 ;
        RECT 0.0050 50.5035 30.3530 50.5790 ;
        RECT 0.0050 52.5470 30.3530 52.6770 ;
        RECT 30.2360 51.5835 30.3530 52.6770 ;
        RECT 16.2140 52.4510 30.2180 52.6770 ;
        RECT 14.8820 52.4510 16.1960 52.6770 ;
        RECT 14.1620 51.5835 14.7920 52.6770 ;
        RECT 0.1400 52.4510 14.1440 52.6770 ;
        RECT 0.0050 51.5835 0.1220 52.6770 ;
        RECT 30.2000 51.5835 30.3530 52.4990 ;
        RECT 16.2680 51.5835 30.1820 52.6770 ;
        RECT 15.5210 51.5835 16.2500 52.4990 ;
        RECT 15.2870 51.7790 15.4850 52.6770 ;
        RECT 14.1080 51.6830 15.2600 52.4990 ;
        RECT 0.1760 51.5835 14.0900 52.6770 ;
        RECT 0.0050 51.5835 0.1580 52.4990 ;
        RECT 15.4670 51.5835 30.3530 52.4030 ;
        RECT 0.0050 51.6830 15.4490 52.4030 ;
        RECT 15.2420 51.5835 30.3530 51.7550 ;
        RECT 0.0050 51.5835 15.2240 52.4030 ;
        RECT 0.0050 51.5835 30.3530 51.6590 ;
        RECT 0.0050 53.6270 30.3530 53.7570 ;
        RECT 30.2360 52.6635 30.3530 53.7570 ;
        RECT 16.2140 53.5310 30.2180 53.7570 ;
        RECT 14.8820 53.5310 16.1960 53.7570 ;
        RECT 14.1620 52.6635 14.7920 53.7570 ;
        RECT 0.1400 53.5310 14.1440 53.7570 ;
        RECT 0.0050 52.6635 0.1220 53.7570 ;
        RECT 30.2000 52.6635 30.3530 53.5790 ;
        RECT 16.2680 52.6635 30.1820 53.7570 ;
        RECT 15.5210 52.6635 16.2500 53.5790 ;
        RECT 15.2870 52.8590 15.4850 53.7570 ;
        RECT 14.1080 52.7630 15.2600 53.5790 ;
        RECT 0.1760 52.6635 14.0900 53.7570 ;
        RECT 0.0050 52.6635 0.1580 53.5790 ;
        RECT 15.4670 52.6635 30.3530 53.4830 ;
        RECT 0.0050 52.7630 15.4490 53.4830 ;
        RECT 15.2420 52.6635 30.3530 52.8350 ;
        RECT 0.0050 52.6635 15.2240 53.4830 ;
        RECT 0.0050 52.6635 30.3530 52.7390 ;
        RECT 0.0050 54.7070 30.3530 54.8370 ;
        RECT 30.2360 53.7435 30.3530 54.8370 ;
        RECT 16.2140 54.6110 30.2180 54.8370 ;
        RECT 14.8820 54.6110 16.1960 54.8370 ;
        RECT 14.1620 53.7435 14.7920 54.8370 ;
        RECT 0.1400 54.6110 14.1440 54.8370 ;
        RECT 0.0050 53.7435 0.1220 54.8370 ;
        RECT 30.2000 53.7435 30.3530 54.6590 ;
        RECT 16.2680 53.7435 30.1820 54.8370 ;
        RECT 15.5210 53.7435 16.2500 54.6590 ;
        RECT 15.2870 53.9390 15.4850 54.8370 ;
        RECT 14.1080 53.8430 15.2600 54.6590 ;
        RECT 0.1760 53.7435 14.0900 54.8370 ;
        RECT 0.0050 53.7435 0.1580 54.6590 ;
        RECT 15.4670 53.7435 30.3530 54.5630 ;
        RECT 0.0050 53.8430 15.4490 54.5630 ;
        RECT 15.2420 53.7435 30.3530 53.9150 ;
        RECT 0.0050 53.7435 15.2240 54.5630 ;
        RECT 0.0050 53.7435 30.3530 53.8190 ;
        RECT 0.0050 55.7870 30.3530 55.9170 ;
        RECT 30.2360 54.8235 30.3530 55.9170 ;
        RECT 16.2140 55.6910 30.2180 55.9170 ;
        RECT 14.8820 55.6910 16.1960 55.9170 ;
        RECT 14.1620 54.8235 14.7920 55.9170 ;
        RECT 0.1400 55.6910 14.1440 55.9170 ;
        RECT 0.0050 54.8235 0.1220 55.9170 ;
        RECT 30.2000 54.8235 30.3530 55.7390 ;
        RECT 16.2680 54.8235 30.1820 55.9170 ;
        RECT 15.5210 54.8235 16.2500 55.7390 ;
        RECT 15.2870 55.0190 15.4850 55.9170 ;
        RECT 14.1080 54.9230 15.2600 55.7390 ;
        RECT 0.1760 54.8235 14.0900 55.9170 ;
        RECT 0.0050 54.8235 0.1580 55.7390 ;
        RECT 15.4670 54.8235 30.3530 55.6430 ;
        RECT 0.0050 54.9230 15.4490 55.6430 ;
        RECT 15.2420 54.8235 30.3530 54.9950 ;
        RECT 0.0050 54.8235 15.2240 55.6430 ;
        RECT 0.0050 54.8235 30.3530 54.8990 ;
        RECT 0.0050 56.8670 30.3530 56.9970 ;
        RECT 30.2360 55.9035 30.3530 56.9970 ;
        RECT 16.2140 56.7710 30.2180 56.9970 ;
        RECT 14.8820 56.7710 16.1960 56.9970 ;
        RECT 14.1620 55.9035 14.7920 56.9970 ;
        RECT 0.1400 56.7710 14.1440 56.9970 ;
        RECT 0.0050 55.9035 0.1220 56.9970 ;
        RECT 30.2000 55.9035 30.3530 56.8190 ;
        RECT 16.2680 55.9035 30.1820 56.9970 ;
        RECT 15.5210 55.9035 16.2500 56.8190 ;
        RECT 15.2870 56.0990 15.4850 56.9970 ;
        RECT 14.1080 56.0030 15.2600 56.8190 ;
        RECT 0.1760 55.9035 14.0900 56.9970 ;
        RECT 0.0050 55.9035 0.1580 56.8190 ;
        RECT 15.4670 55.9035 30.3530 56.7230 ;
        RECT 0.0050 56.0030 15.4490 56.7230 ;
        RECT 15.2420 55.9035 30.3530 56.0750 ;
        RECT 0.0050 55.9035 15.2240 56.7230 ;
        RECT 0.0050 55.9035 30.3530 55.9790 ;
        RECT 0.0050 57.9470 30.3530 58.0770 ;
        RECT 30.2360 56.9835 30.3530 58.0770 ;
        RECT 16.2140 57.8510 30.2180 58.0770 ;
        RECT 14.8820 57.8510 16.1960 58.0770 ;
        RECT 14.1620 56.9835 14.7920 58.0770 ;
        RECT 0.1400 57.8510 14.1440 58.0770 ;
        RECT 0.0050 56.9835 0.1220 58.0770 ;
        RECT 30.2000 56.9835 30.3530 57.8990 ;
        RECT 16.2680 56.9835 30.1820 58.0770 ;
        RECT 15.5210 56.9835 16.2500 57.8990 ;
        RECT 15.2870 57.1790 15.4850 58.0770 ;
        RECT 14.1080 57.0830 15.2600 57.8990 ;
        RECT 0.1760 56.9835 14.0900 58.0770 ;
        RECT 0.0050 56.9835 0.1580 57.8990 ;
        RECT 15.4670 56.9835 30.3530 57.8030 ;
        RECT 0.0050 57.0830 15.4490 57.8030 ;
        RECT 15.2420 56.9835 30.3530 57.1550 ;
        RECT 0.0050 56.9835 15.2240 57.8030 ;
        RECT 0.0050 56.9835 30.3530 57.0590 ;
        RECT 0.0050 59.0270 30.3530 59.1570 ;
        RECT 30.2360 58.0635 30.3530 59.1570 ;
        RECT 16.2140 58.9310 30.2180 59.1570 ;
        RECT 14.8820 58.9310 16.1960 59.1570 ;
        RECT 14.1620 58.0635 14.7920 59.1570 ;
        RECT 0.1400 58.9310 14.1440 59.1570 ;
        RECT 0.0050 58.0635 0.1220 59.1570 ;
        RECT 30.2000 58.0635 30.3530 58.9790 ;
        RECT 16.2680 58.0635 30.1820 59.1570 ;
        RECT 15.5210 58.0635 16.2500 58.9790 ;
        RECT 15.2870 58.2590 15.4850 59.1570 ;
        RECT 14.1080 58.1630 15.2600 58.9790 ;
        RECT 0.1760 58.0635 14.0900 59.1570 ;
        RECT 0.0050 58.0635 0.1580 58.9790 ;
        RECT 15.4670 58.0635 30.3530 58.8830 ;
        RECT 0.0050 58.1630 15.4490 58.8830 ;
        RECT 15.2420 58.0635 30.3530 58.2350 ;
        RECT 0.0050 58.0635 15.2240 58.8830 ;
        RECT 0.0050 58.0635 30.3530 58.1390 ;
        RECT 0.0050 60.1070 30.3530 60.2370 ;
        RECT 30.2360 59.1435 30.3530 60.2370 ;
        RECT 16.2140 60.0110 30.2180 60.2370 ;
        RECT 14.8820 60.0110 16.1960 60.2370 ;
        RECT 14.1620 59.1435 14.7920 60.2370 ;
        RECT 0.1400 60.0110 14.1440 60.2370 ;
        RECT 0.0050 59.1435 0.1220 60.2370 ;
        RECT 30.2000 59.1435 30.3530 60.0590 ;
        RECT 16.2680 59.1435 30.1820 60.2370 ;
        RECT 15.5210 59.1435 16.2500 60.0590 ;
        RECT 15.2870 59.3390 15.4850 60.2370 ;
        RECT 14.1080 59.2430 15.2600 60.0590 ;
        RECT 0.1760 59.1435 14.0900 60.2370 ;
        RECT 0.0050 59.1435 0.1580 60.0590 ;
        RECT 15.4670 59.1435 30.3530 59.9630 ;
        RECT 0.0050 59.2430 15.4490 59.9630 ;
        RECT 15.2420 59.1435 30.3530 59.3150 ;
        RECT 0.0050 59.1435 15.2240 59.9630 ;
        RECT 0.0050 59.1435 30.3530 59.2190 ;
        RECT 0.0050 61.1870 30.3530 61.3170 ;
        RECT 30.2360 60.2235 30.3530 61.3170 ;
        RECT 16.2140 61.0910 30.2180 61.3170 ;
        RECT 14.8820 61.0910 16.1960 61.3170 ;
        RECT 14.1620 60.2235 14.7920 61.3170 ;
        RECT 0.1400 61.0910 14.1440 61.3170 ;
        RECT 0.0050 60.2235 0.1220 61.3170 ;
        RECT 30.2000 60.2235 30.3530 61.1390 ;
        RECT 16.2680 60.2235 30.1820 61.3170 ;
        RECT 15.5210 60.2235 16.2500 61.1390 ;
        RECT 15.2870 60.4190 15.4850 61.3170 ;
        RECT 14.1080 60.3230 15.2600 61.1390 ;
        RECT 0.1760 60.2235 14.0900 61.3170 ;
        RECT 0.0050 60.2235 0.1580 61.1390 ;
        RECT 15.4670 60.2235 30.3530 61.0430 ;
        RECT 0.0050 60.3230 15.4490 61.0430 ;
        RECT 15.2420 60.2235 30.3530 60.3950 ;
        RECT 0.0050 60.2235 15.2240 61.0430 ;
        RECT 0.0050 60.2235 30.3530 60.2990 ;
        RECT 0.0050 62.2670 30.3530 62.3970 ;
        RECT 30.2360 61.3035 30.3530 62.3970 ;
        RECT 16.2140 62.1710 30.2180 62.3970 ;
        RECT 14.8820 62.1710 16.1960 62.3970 ;
        RECT 14.1620 61.3035 14.7920 62.3970 ;
        RECT 0.1400 62.1710 14.1440 62.3970 ;
        RECT 0.0050 61.3035 0.1220 62.3970 ;
        RECT 30.2000 61.3035 30.3530 62.2190 ;
        RECT 16.2680 61.3035 30.1820 62.3970 ;
        RECT 15.5210 61.3035 16.2500 62.2190 ;
        RECT 15.2870 61.4990 15.4850 62.3970 ;
        RECT 14.1080 61.4030 15.2600 62.2190 ;
        RECT 0.1760 61.3035 14.0900 62.3970 ;
        RECT 0.0050 61.3035 0.1580 62.2190 ;
        RECT 15.4670 61.3035 30.3530 62.1230 ;
        RECT 0.0050 61.4030 15.4490 62.1230 ;
        RECT 15.2420 61.3035 30.3530 61.4750 ;
        RECT 0.0050 61.3035 15.2240 62.1230 ;
        RECT 0.0050 61.3035 30.3530 61.3790 ;
        RECT 0.0050 63.3470 30.3530 63.4770 ;
        RECT 30.2360 62.3835 30.3530 63.4770 ;
        RECT 16.2140 63.2510 30.2180 63.4770 ;
        RECT 14.8820 63.2510 16.1960 63.4770 ;
        RECT 14.1620 62.3835 14.7920 63.4770 ;
        RECT 0.1400 63.2510 14.1440 63.4770 ;
        RECT 0.0050 62.3835 0.1220 63.4770 ;
        RECT 30.2000 62.3835 30.3530 63.2990 ;
        RECT 16.2680 62.3835 30.1820 63.4770 ;
        RECT 15.5210 62.3835 16.2500 63.2990 ;
        RECT 15.2870 62.5790 15.4850 63.4770 ;
        RECT 14.1080 62.4830 15.2600 63.2990 ;
        RECT 0.1760 62.3835 14.0900 63.4770 ;
        RECT 0.0050 62.3835 0.1580 63.2990 ;
        RECT 15.4670 62.3835 30.3530 63.2030 ;
        RECT 0.0050 62.4830 15.4490 63.2030 ;
        RECT 15.2420 62.3835 30.3530 62.5550 ;
        RECT 0.0050 62.3835 15.2240 63.2030 ;
        RECT 0.0050 62.3835 30.3530 62.4590 ;
        RECT 0.0050 64.4270 30.3530 64.5570 ;
        RECT 30.2360 63.4635 30.3530 64.5570 ;
        RECT 16.2140 64.3310 30.2180 64.5570 ;
        RECT 14.8820 64.3310 16.1960 64.5570 ;
        RECT 14.1620 63.4635 14.7920 64.5570 ;
        RECT 0.1400 64.3310 14.1440 64.5570 ;
        RECT 0.0050 63.4635 0.1220 64.5570 ;
        RECT 30.2000 63.4635 30.3530 64.3790 ;
        RECT 16.2680 63.4635 30.1820 64.5570 ;
        RECT 15.5210 63.4635 16.2500 64.3790 ;
        RECT 15.2870 63.6590 15.4850 64.5570 ;
        RECT 14.1080 63.5630 15.2600 64.3790 ;
        RECT 0.1760 63.4635 14.0900 64.5570 ;
        RECT 0.0050 63.4635 0.1580 64.3790 ;
        RECT 15.4670 63.4635 30.3530 64.2830 ;
        RECT 0.0050 63.5630 15.4490 64.2830 ;
        RECT 15.2420 63.4635 30.3530 63.6350 ;
        RECT 0.0050 63.4635 15.2240 64.2830 ;
        RECT 0.0050 63.4635 30.3530 63.5390 ;
        RECT 0.0050 65.5070 30.3530 65.6370 ;
        RECT 30.2360 64.5435 30.3530 65.6370 ;
        RECT 16.2140 65.4110 30.2180 65.6370 ;
        RECT 14.8820 65.4110 16.1960 65.6370 ;
        RECT 14.1620 64.5435 14.7920 65.6370 ;
        RECT 0.1400 65.4110 14.1440 65.6370 ;
        RECT 0.0050 64.5435 0.1220 65.6370 ;
        RECT 30.2000 64.5435 30.3530 65.4590 ;
        RECT 16.2680 64.5435 30.1820 65.6370 ;
        RECT 15.5210 64.5435 16.2500 65.4590 ;
        RECT 15.2870 64.7390 15.4850 65.6370 ;
        RECT 14.1080 64.6430 15.2600 65.4590 ;
        RECT 0.1760 64.5435 14.0900 65.6370 ;
        RECT 0.0050 64.5435 0.1580 65.4590 ;
        RECT 15.4670 64.5435 30.3530 65.3630 ;
        RECT 0.0050 64.6430 15.4490 65.3630 ;
        RECT 15.2420 64.5435 30.3530 64.7150 ;
        RECT 0.0050 64.5435 15.2240 65.3630 ;
        RECT 0.0050 64.5435 30.3530 64.6190 ;
        RECT 0.0050 66.5870 30.3530 66.7170 ;
        RECT 30.2360 65.6235 30.3530 66.7170 ;
        RECT 16.2140 66.4910 30.2180 66.7170 ;
        RECT 14.8820 66.4910 16.1960 66.7170 ;
        RECT 14.1620 65.6235 14.7920 66.7170 ;
        RECT 0.1400 66.4910 14.1440 66.7170 ;
        RECT 0.0050 65.6235 0.1220 66.7170 ;
        RECT 30.2000 65.6235 30.3530 66.5390 ;
        RECT 16.2680 65.6235 30.1820 66.7170 ;
        RECT 15.5210 65.6235 16.2500 66.5390 ;
        RECT 15.2870 65.8190 15.4850 66.7170 ;
        RECT 14.1080 65.7230 15.2600 66.5390 ;
        RECT 0.1760 65.6235 14.0900 66.7170 ;
        RECT 0.0050 65.6235 0.1580 66.5390 ;
        RECT 15.4670 65.6235 30.3530 66.4430 ;
        RECT 0.0050 65.7230 15.4490 66.4430 ;
        RECT 15.2420 65.6235 30.3530 65.7950 ;
        RECT 0.0050 65.6235 15.2240 66.4430 ;
        RECT 0.0050 65.6235 30.3530 65.6990 ;
        RECT 0.0050 67.6670 30.3530 67.7970 ;
        RECT 30.2360 66.7035 30.3530 67.7970 ;
        RECT 16.2140 67.5710 30.2180 67.7970 ;
        RECT 14.8820 67.5710 16.1960 67.7970 ;
        RECT 14.1620 66.7035 14.7920 67.7970 ;
        RECT 0.1400 67.5710 14.1440 67.7970 ;
        RECT 0.0050 66.7035 0.1220 67.7970 ;
        RECT 30.2000 66.7035 30.3530 67.6190 ;
        RECT 16.2680 66.7035 30.1820 67.7970 ;
        RECT 15.5210 66.7035 16.2500 67.6190 ;
        RECT 15.2870 66.8990 15.4850 67.7970 ;
        RECT 14.1080 66.8030 15.2600 67.6190 ;
        RECT 0.1760 66.7035 14.0900 67.7970 ;
        RECT 0.0050 66.7035 0.1580 67.6190 ;
        RECT 15.4670 66.7035 30.3530 67.5230 ;
        RECT 0.0050 66.8030 15.4490 67.5230 ;
        RECT 15.2420 66.7035 30.3530 66.8750 ;
        RECT 0.0050 66.7035 15.2240 67.5230 ;
        RECT 0.0050 66.7035 30.3530 66.7790 ;
        RECT 0.0050 68.7470 30.3530 68.8770 ;
        RECT 30.2360 67.7835 30.3530 68.8770 ;
        RECT 16.2140 68.6510 30.2180 68.8770 ;
        RECT 14.8820 68.6510 16.1960 68.8770 ;
        RECT 14.1620 67.7835 14.7920 68.8770 ;
        RECT 0.1400 68.6510 14.1440 68.8770 ;
        RECT 0.0050 67.7835 0.1220 68.8770 ;
        RECT 30.2000 67.7835 30.3530 68.6990 ;
        RECT 16.2680 67.7835 30.1820 68.8770 ;
        RECT 15.5210 67.7835 16.2500 68.6990 ;
        RECT 15.2870 67.9790 15.4850 68.8770 ;
        RECT 14.1080 67.8830 15.2600 68.6990 ;
        RECT 0.1760 67.7835 14.0900 68.8770 ;
        RECT 0.0050 67.7835 0.1580 68.6990 ;
        RECT 15.4670 67.7835 30.3530 68.6030 ;
        RECT 0.0050 67.8830 15.4490 68.6030 ;
        RECT 15.2420 67.7835 30.3530 67.9550 ;
        RECT 0.0050 67.7835 15.2240 68.6030 ;
        RECT 0.0050 67.7835 30.3530 67.8590 ;
        RECT 0.0050 69.8270 30.3530 69.9570 ;
        RECT 30.2360 68.8635 30.3530 69.9570 ;
        RECT 16.2140 69.7310 30.2180 69.9570 ;
        RECT 14.8820 69.7310 16.1960 69.9570 ;
        RECT 14.1620 68.8635 14.7920 69.9570 ;
        RECT 0.1400 69.7310 14.1440 69.9570 ;
        RECT 0.0050 68.8635 0.1220 69.9570 ;
        RECT 30.2000 68.8635 30.3530 69.7790 ;
        RECT 16.2680 68.8635 30.1820 69.9570 ;
        RECT 15.5210 68.8635 16.2500 69.7790 ;
        RECT 15.2870 69.0590 15.4850 69.9570 ;
        RECT 14.1080 68.9630 15.2600 69.7790 ;
        RECT 0.1760 68.8635 14.0900 69.9570 ;
        RECT 0.0050 68.8635 0.1580 69.7790 ;
        RECT 15.4670 68.8635 30.3530 69.6830 ;
        RECT 0.0050 68.9630 15.4490 69.6830 ;
        RECT 15.2420 68.8635 30.3530 69.0350 ;
        RECT 0.0050 68.8635 15.2240 69.6830 ;
        RECT 0.0050 68.8635 30.3530 68.9390 ;
        RECT 0.0050 70.9070 30.3530 71.0370 ;
        RECT 30.2360 69.9435 30.3530 71.0370 ;
        RECT 16.2140 70.8110 30.2180 71.0370 ;
        RECT 14.8820 70.8110 16.1960 71.0370 ;
        RECT 14.1620 69.9435 14.7920 71.0370 ;
        RECT 0.1400 70.8110 14.1440 71.0370 ;
        RECT 0.0050 69.9435 0.1220 71.0370 ;
        RECT 30.2000 69.9435 30.3530 70.8590 ;
        RECT 16.2680 69.9435 30.1820 71.0370 ;
        RECT 15.5210 69.9435 16.2500 70.8590 ;
        RECT 15.2870 70.1390 15.4850 71.0370 ;
        RECT 14.1080 70.0430 15.2600 70.8590 ;
        RECT 0.1760 69.9435 14.0900 71.0370 ;
        RECT 0.0050 69.9435 0.1580 70.8590 ;
        RECT 15.4670 69.9435 30.3530 70.7630 ;
        RECT 0.0050 70.0430 15.4490 70.7630 ;
        RECT 15.2420 69.9435 30.3530 70.1150 ;
        RECT 0.0050 69.9435 15.2240 70.7630 ;
        RECT 0.0050 69.9435 30.3530 70.0190 ;
        RECT 0.0050 71.9870 30.3530 72.1170 ;
        RECT 30.2360 71.0235 30.3530 72.1170 ;
        RECT 16.2140 71.8910 30.2180 72.1170 ;
        RECT 14.8820 71.8910 16.1960 72.1170 ;
        RECT 14.1620 71.0235 14.7920 72.1170 ;
        RECT 0.1400 71.8910 14.1440 72.1170 ;
        RECT 0.0050 71.0235 0.1220 72.1170 ;
        RECT 30.2000 71.0235 30.3530 71.9390 ;
        RECT 16.2680 71.0235 30.1820 72.1170 ;
        RECT 15.5210 71.0235 16.2500 71.9390 ;
        RECT 15.2870 71.2190 15.4850 72.1170 ;
        RECT 14.1080 71.1230 15.2600 71.9390 ;
        RECT 0.1760 71.0235 14.0900 72.1170 ;
        RECT 0.0050 71.0235 0.1580 71.9390 ;
        RECT 15.4670 71.0235 30.3530 71.8430 ;
        RECT 0.0050 71.1230 15.4490 71.8430 ;
        RECT 15.2420 71.0235 30.3530 71.1950 ;
        RECT 0.0050 71.0235 15.2240 71.8430 ;
        RECT 0.0050 71.0235 30.3530 71.0990 ;
        RECT 0.0050 73.0670 30.3530 73.1970 ;
        RECT 30.2360 72.1035 30.3530 73.1970 ;
        RECT 16.2140 72.9710 30.2180 73.1970 ;
        RECT 14.8820 72.9710 16.1960 73.1970 ;
        RECT 14.1620 72.1035 14.7920 73.1970 ;
        RECT 0.1400 72.9710 14.1440 73.1970 ;
        RECT 0.0050 72.1035 0.1220 73.1970 ;
        RECT 30.2000 72.1035 30.3530 73.0190 ;
        RECT 16.2680 72.1035 30.1820 73.1970 ;
        RECT 15.5210 72.1035 16.2500 73.0190 ;
        RECT 15.2870 72.2990 15.4850 73.1970 ;
        RECT 14.1080 72.2030 15.2600 73.0190 ;
        RECT 0.1760 72.1035 14.0900 73.1970 ;
        RECT 0.0050 72.1035 0.1580 73.0190 ;
        RECT 15.4670 72.1035 30.3530 72.9230 ;
        RECT 0.0050 72.2030 15.4490 72.9230 ;
        RECT 15.2420 72.1035 30.3530 72.2750 ;
        RECT 0.0050 72.1035 15.2240 72.9230 ;
        RECT 0.0050 72.1035 30.3530 72.1790 ;
        RECT 0.0050 74.1470 30.3530 74.2770 ;
        RECT 30.2360 73.1835 30.3530 74.2770 ;
        RECT 16.2140 74.0510 30.2180 74.2770 ;
        RECT 14.8820 74.0510 16.1960 74.2770 ;
        RECT 14.1620 73.1835 14.7920 74.2770 ;
        RECT 0.1400 74.0510 14.1440 74.2770 ;
        RECT 0.0050 73.1835 0.1220 74.2770 ;
        RECT 30.2000 73.1835 30.3530 74.0990 ;
        RECT 16.2680 73.1835 30.1820 74.2770 ;
        RECT 15.5210 73.1835 16.2500 74.0990 ;
        RECT 15.2870 73.3790 15.4850 74.2770 ;
        RECT 14.1080 73.2830 15.2600 74.0990 ;
        RECT 0.1760 73.1835 14.0900 74.2770 ;
        RECT 0.0050 73.1835 0.1580 74.0990 ;
        RECT 15.4670 73.1835 30.3530 74.0030 ;
        RECT 0.0050 73.2830 15.4490 74.0030 ;
        RECT 15.2420 73.1835 30.3530 73.3550 ;
        RECT 0.0050 73.1835 15.2240 74.0030 ;
        RECT 0.0050 73.1835 30.3530 73.2590 ;
        RECT 0.0050 75.2270 30.3530 75.3570 ;
        RECT 30.2360 74.2635 30.3530 75.3570 ;
        RECT 16.2140 75.1310 30.2180 75.3570 ;
        RECT 14.8820 75.1310 16.1960 75.3570 ;
        RECT 14.1620 74.2635 14.7920 75.3570 ;
        RECT 0.1400 75.1310 14.1440 75.3570 ;
        RECT 0.0050 74.2635 0.1220 75.3570 ;
        RECT 30.2000 74.2635 30.3530 75.1790 ;
        RECT 16.2680 74.2635 30.1820 75.3570 ;
        RECT 15.5210 74.2635 16.2500 75.1790 ;
        RECT 15.2870 74.4590 15.4850 75.3570 ;
        RECT 14.1080 74.3630 15.2600 75.1790 ;
        RECT 0.1760 74.2635 14.0900 75.3570 ;
        RECT 0.0050 74.2635 0.1580 75.1790 ;
        RECT 15.4670 74.2635 30.3530 75.0830 ;
        RECT 0.0050 74.3630 15.4490 75.0830 ;
        RECT 15.2420 74.2635 30.3530 74.4350 ;
        RECT 0.0050 74.2635 15.2240 75.0830 ;
        RECT 0.0050 74.2635 30.3530 74.3390 ;
        RECT 0.0050 76.3070 30.3530 76.4370 ;
        RECT 30.2360 75.3435 30.3530 76.4370 ;
        RECT 16.2140 76.2110 30.2180 76.4370 ;
        RECT 14.8820 76.2110 16.1960 76.4370 ;
        RECT 14.1620 75.3435 14.7920 76.4370 ;
        RECT 0.1400 76.2110 14.1440 76.4370 ;
        RECT 0.0050 75.3435 0.1220 76.4370 ;
        RECT 30.2000 75.3435 30.3530 76.2590 ;
        RECT 16.2680 75.3435 30.1820 76.4370 ;
        RECT 15.5210 75.3435 16.2500 76.2590 ;
        RECT 15.2870 75.5390 15.4850 76.4370 ;
        RECT 14.1080 75.4430 15.2600 76.2590 ;
        RECT 0.1760 75.3435 14.0900 76.4370 ;
        RECT 0.0050 75.3435 0.1580 76.2590 ;
        RECT 15.4670 75.3435 30.3530 76.1630 ;
        RECT 0.0050 75.4430 15.4490 76.1630 ;
        RECT 15.2420 75.3435 30.3530 75.5150 ;
        RECT 0.0050 75.3435 15.2240 76.1630 ;
        RECT 0.0050 75.3435 30.3530 75.4190 ;
        RECT 0.0050 77.3870 30.3530 77.5170 ;
        RECT 30.2360 76.4235 30.3530 77.5170 ;
        RECT 16.2140 77.2910 30.2180 77.5170 ;
        RECT 14.8820 77.2910 16.1960 77.5170 ;
        RECT 14.1620 76.4235 14.7920 77.5170 ;
        RECT 0.1400 77.2910 14.1440 77.5170 ;
        RECT 0.0050 76.4235 0.1220 77.5170 ;
        RECT 30.2000 76.4235 30.3530 77.3390 ;
        RECT 16.2680 76.4235 30.1820 77.5170 ;
        RECT 15.5210 76.4235 16.2500 77.3390 ;
        RECT 15.2870 76.6190 15.4850 77.5170 ;
        RECT 14.1080 76.5230 15.2600 77.3390 ;
        RECT 0.1760 76.4235 14.0900 77.5170 ;
        RECT 0.0050 76.4235 0.1580 77.3390 ;
        RECT 15.4670 76.4235 30.3530 77.2430 ;
        RECT 0.0050 76.5230 15.4490 77.2430 ;
        RECT 15.2420 76.4235 30.3530 76.5950 ;
        RECT 0.0050 76.4235 15.2240 77.2430 ;
        RECT 0.0050 76.4235 30.3530 76.4990 ;
  LAYER M4  ;
      RECT 1.6000 36.5665 28.8355 36.5905 ;
      RECT 1.6000 36.8545 28.8355 36.8785 ;
      RECT 1.6000 37.2385 28.8355 37.2625 ;
      RECT 1.6000 37.3345 28.8355 37.3585 ;
      RECT 1.6000 37.6705 28.8355 37.6945 ;
      RECT 1.6000 38.0545 28.8355 38.0785 ;
      RECT 1.6000 38.1505 28.8355 38.1745 ;
      RECT 10.4760 35.1895 19.8720 35.4055 ;
      RECT 17.8670 35.5255 17.9510 35.5495 ;
      RECT 17.6785 35.9575 17.8085 35.9815 ;
      RECT 17.6870 36.9025 17.8040 36.9265 ;
      RECT 17.6865 36.6150 17.8035 36.6390 ;
      RECT 17.0375 35.9575 17.6085 35.9815 ;
      RECT 17.0975 36.7225 17.2055 36.7465 ;
      RECT 15.7750 37.1095 16.8680 37.1335 ;
      RECT 16.4630 36.6775 16.5470 36.7015 ;
      RECT 15.6790 37.8775 16.5470 37.9015 ;
      RECT 16.4630 37.9735 16.5470 37.9975 ;
      RECT 16.2850 36.1975 16.3690 36.2215 ;
      RECT 16.2470 37.5415 16.3310 37.5655 ;
      RECT 16.2470 38.2615 16.3310 38.2855 ;
      RECT 15.9780 34.9095 16.2410 34.9335 ;
      RECT 16.1090 38.6935 16.2210 38.7175 ;
      RECT 16.0690 36.1015 16.1530 36.1255 ;
      RECT 15.8550 34.8135 16.1180 34.8375 ;
      RECT 15.8550 43.4185 16.1180 43.4425 ;
      RECT 15.8710 37.5895 16.1150 37.6135 ;
      RECT 16.0310 37.7335 16.1150 37.7575 ;
      RECT 14.5750 37.9735 16.1150 37.9975 ;
      RECT 16.0310 38.2615 16.1150 38.2855 ;
      RECT 15.7970 43.3225 16.0600 43.3465 ;
      RECT 15.7960 34.7175 16.0590 34.7415 ;
      RECT 14.3100 38.3575 16.0380 38.5735 ;
      RECT 14.3100 41.5255 16.0380 41.7415 ;
      RECT 15.7580 34.6215 16.0210 34.6455 ;
      RECT 15.7580 43.1305 16.0210 43.1545 ;
      RECT 15.9230 38.6935 16.0070 38.7175 ;
      RECT 15.1510 39.0775 16.0070 39.1015 ;
      RECT 15.5350 41.3335 16.0070 41.3575 ;
      RECT 15.9230 41.4295 16.0070 41.4535 ;
      RECT 15.7100 34.5255 15.9730 34.5495 ;
      RECT 15.7100 43.0345 15.9730 43.0585 ;
      RECT 15.4870 40.4215 15.9320 40.4455 ;
      RECT 15.6660 34.4295 15.9290 34.4535 ;
      RECT 15.6660 43.3705 15.9290 43.3945 ;
      RECT 15.6170 34.7655 15.8800 34.7895 ;
      RECT 15.6170 43.2745 15.8800 43.2985 ;
      RECT 15.7480 37.7335 15.8690 37.7575 ;
      RECT 15.7270 39.8455 15.8600 39.8695 ;
      RECT 15.5700 34.6695 15.8330 34.6935 ;
      RECT 15.5700 43.1785 15.8330 43.2025 ;
      RECT 15.5350 34.3815 15.7980 34.4055 ;
      RECT 15.5350 43.0825 15.7980 43.1065 ;
      RECT 14.7190 41.4295 15.7880 41.4535 ;
      RECT 15.7040 42.5815 15.7880 42.6055 ;
      RECT 15.4790 34.2375 15.7420 34.2615 ;
      RECT 15.4790 42.9865 15.7420 43.0105 ;
      RECT 15.6310 38.6935 15.7160 38.7175 ;
      RECT 14.5270 39.2695 15.6440 39.2935 ;
      RECT 15.1720 37.1095 15.6290 37.1335 ;
      RECT 14.9990 34.9575 15.2660 34.9815 ;
      RECT 14.9990 42.8425 15.2660 42.8665 ;
      RECT 15.1360 38.6455 15.2450 38.6695 ;
      RECT 14.9760 34.8615 15.2180 34.8855 ;
      RECT 14.9760 43.4665 15.2180 43.4905 ;
      RECT 14.9200 34.3815 15.1620 34.4055 ;
      RECT 14.9490 43.5625 15.1620 43.5865 ;
      RECT 15.0650 38.2615 15.1490 38.2855 ;
      RECT 14.8660 34.4775 15.1140 34.5015 ;
      RECT 14.8660 43.4185 15.1140 43.4425 ;
      RECT 14.6320 40.8535 15.0530 40.8775 ;
      RECT 14.6000 34.8135 14.8670 34.8375 ;
      RECT 14.6000 43.5625 14.8670 43.5865 ;
      RECT 14.7400 39.4135 14.8610 39.4375 ;
      RECT 14.7320 42.5815 14.8160 42.6055 ;
      RECT 14.5660 34.7175 14.8130 34.7415 ;
      RECT 14.4990 43.1305 14.8130 43.1545 ;
      RECT 14.5400 34.6215 14.7700 34.6455 ;
      RECT 14.5280 43.4665 14.7700 43.4905 ;
      RECT 14.4870 34.5255 14.7170 34.5495 ;
      RECT 14.6330 40.9975 14.7170 41.0215 ;
      RECT 14.4370 43.0345 14.7170 43.0585 ;
      RECT 14.4420 34.4295 14.6720 34.4535 ;
      RECT 14.4420 43.3705 14.6720 43.3945 ;
      RECT 13.4800 38.2615 14.6690 38.2855 ;
      RECT 14.4040 34.6695 14.6340 34.6935 ;
      RECT 14.4040 43.2745 14.6340 43.2985 ;
      RECT 14.3860 34.5735 14.5790 34.5975 ;
      RECT 14.3860 43.1785 14.5790 43.2025 ;
      RECT 14.3370 34.4775 14.5300 34.5015 ;
      RECT 14.3370 43.0825 14.5300 43.1065 ;
      RECT 14.3410 39.1735 14.5250 39.1975 ;
      RECT 14.2850 34.3815 14.4780 34.4055 ;
      RECT 14.2850 42.9865 14.4780 43.0105 ;
      RECT 13.8010 36.4855 14.4770 36.5095 ;
      RECT 14.3410 39.2695 14.4250 39.2935 ;
      RECT 14.0720 34.9095 14.3350 34.9335 ;
      RECT 14.1950 37.1095 14.2790 37.1335 ;
      RECT 14.1260 38.6935 14.2380 38.7175 ;
      RECT 13.7630 36.6775 13.8470 36.7015 ;
  LAYER V4  ;
      RECT 17.9160 35.5255 17.9400 35.5495 ;
      RECT 17.9160 36.5665 17.9400 36.5905 ;
      RECT 17.7480 36.6150 17.7720 36.6390 ;
      RECT 17.7480 36.9025 17.7720 36.9265 ;
      RECT 17.7475 35.9575 17.7715 35.9815 ;
      RECT 17.1135 35.9575 17.1375 35.9815 ;
      RECT 17.1135 36.7225 17.1375 36.7465 ;
      RECT 16.5120 36.6775 16.5360 36.7015 ;
      RECT 16.5120 36.8545 16.5360 36.8785 ;
      RECT 16.5120 37.8775 16.5360 37.9015 ;
      RECT 16.5120 37.9735 16.5360 37.9975 ;
      RECT 16.2960 36.1975 16.3200 36.2215 ;
      RECT 16.2960 37.2385 16.3200 37.2625 ;
      RECT 16.2960 37.5415 16.3200 37.5655 ;
      RECT 16.2960 37.6705 16.3200 37.6945 ;
      RECT 16.2960 38.0545 16.3200 38.0785 ;
      RECT 16.2960 38.2615 16.3200 38.2855 ;
      RECT 16.1270 34.9095 16.1510 34.9335 ;
      RECT 16.1280 35.1895 16.1510 35.4055 ;
      RECT 16.1270 38.6935 16.1510 38.7175 ;
      RECT 16.0800 36.1015 16.1040 36.1255 ;
      RECT 16.0800 37.3345 16.1040 37.3585 ;
      RECT 16.0800 37.5895 16.1040 37.6135 ;
      RECT 16.0800 37.7335 16.1040 37.7575 ;
      RECT 16.0800 37.9735 16.1040 37.9975 ;
      RECT 16.0800 38.2615 16.1040 38.2855 ;
      RECT 15.9720 38.6935 15.9960 38.7175 ;
      RECT 15.9720 39.0775 15.9960 39.1015 ;
      RECT 15.9720 41.3335 15.9960 41.3575 ;
      RECT 15.9720 41.4295 15.9960 41.4535 ;
      RECT 15.8820 34.8135 15.9060 34.8375 ;
      RECT 15.8820 37.5895 15.9060 37.6135 ;
      RECT 15.8820 43.4185 15.9060 43.4425 ;
      RECT 15.8340 34.7175 15.8580 34.7415 ;
      RECT 15.8340 37.7335 15.8580 37.7575 ;
      RECT 15.8340 43.3225 15.8580 43.3465 ;
      RECT 15.7860 34.6215 15.8100 34.6455 ;
      RECT 15.7860 37.1095 15.8100 37.1335 ;
      RECT 15.7860 43.1305 15.8100 43.1545 ;
      RECT 15.7380 34.5255 15.7620 34.5495 ;
      RECT 15.7380 39.8455 15.7620 39.8695 ;
      RECT 15.7380 42.5815 15.7620 42.6055 ;
      RECT 15.7380 43.0345 15.7620 43.0585 ;
      RECT 15.6900 34.4295 15.7140 34.4535 ;
      RECT 15.6900 37.8775 15.7140 37.9015 ;
      RECT 15.6900 43.3705 15.7140 43.3945 ;
      RECT 15.6420 34.7655 15.6660 34.7895 ;
      RECT 15.6420 38.6935 15.6660 38.7175 ;
      RECT 15.6420 43.2745 15.6660 43.2985 ;
      RECT 15.5940 34.6695 15.6180 34.6935 ;
      RECT 15.5940 37.1095 15.6180 37.1335 ;
      RECT 15.5940 43.1785 15.6180 43.2025 ;
      RECT 15.5460 34.3815 15.5700 34.4055 ;
      RECT 15.5460 41.3335 15.5700 41.3575 ;
      RECT 15.5460 43.0825 15.5700 43.1065 ;
      RECT 15.4980 34.2375 15.5220 34.2615 ;
      RECT 15.4980 40.4215 15.5220 40.4455 ;
      RECT 15.4980 42.9865 15.5220 43.0105 ;
      RECT 15.2100 34.9575 15.2340 34.9815 ;
      RECT 15.2100 38.6455 15.2340 38.6695 ;
      RECT 15.2100 42.8425 15.2340 42.8665 ;
      RECT 15.1620 34.8615 15.1860 34.8855 ;
      RECT 15.1620 39.0775 15.1860 39.1015 ;
      RECT 15.1620 43.4665 15.1860 43.4905 ;
      RECT 15.1140 34.3815 15.1380 34.4055 ;
      RECT 15.1140 38.2615 15.1380 38.2855 ;
      RECT 15.1140 43.5625 15.1380 43.5865 ;
      RECT 15.0180 34.4775 15.0420 34.5015 ;
      RECT 15.0180 40.8535 15.0420 40.8775 ;
      RECT 15.0180 43.4185 15.0420 43.4425 ;
      RECT 14.8260 34.8135 14.8500 34.8375 ;
      RECT 14.8260 39.4135 14.8500 39.4375 ;
      RECT 14.8260 43.5625 14.8500 43.5865 ;
      RECT 14.7780 34.7175 14.8020 34.7415 ;
      RECT 14.7780 42.5815 14.8020 42.6055 ;
      RECT 14.7780 43.1305 14.8020 43.1545 ;
      RECT 14.7300 34.6215 14.7540 34.6455 ;
      RECT 14.7300 41.4295 14.7540 41.4535 ;
      RECT 14.7300 43.4665 14.7540 43.4905 ;
      RECT 14.6820 34.5255 14.7060 34.5495 ;
      RECT 14.6820 40.9975 14.7060 41.0215 ;
      RECT 14.6820 43.0345 14.7060 43.0585 ;
      RECT 14.6340 34.4295 14.6580 34.4535 ;
      RECT 14.6340 38.2615 14.6580 38.2855 ;
      RECT 14.6340 43.3705 14.6580 43.3945 ;
      RECT 14.5860 34.6695 14.6100 34.6935 ;
      RECT 14.5860 37.9735 14.6100 37.9975 ;
      RECT 14.5860 43.2745 14.6100 43.2985 ;
      RECT 14.5380 34.5735 14.5620 34.5975 ;
      RECT 14.5380 39.2695 14.5620 39.2935 ;
      RECT 14.5380 43.1785 14.5620 43.2025 ;
      RECT 14.4900 34.4775 14.5140 34.5015 ;
      RECT 14.4900 39.1735 14.5140 39.1975 ;
      RECT 14.4900 43.0825 14.5140 43.1065 ;
      RECT 14.4420 34.3815 14.4660 34.4055 ;
      RECT 14.4420 36.4855 14.4660 36.5095 ;
      RECT 14.4420 42.9865 14.4660 43.0105 ;
      RECT 14.3520 39.1735 14.3760 39.1975 ;
      RECT 14.3520 39.2695 14.3760 39.2935 ;
      RECT 14.2440 37.1095 14.2680 37.1335 ;
      RECT 14.2440 38.1505 14.2680 38.1745 ;
      RECT 14.1840 34.9095 14.2080 34.9335 ;
      RECT 14.1850 35.1895 14.2080 35.4055 ;
      RECT 14.1840 38.6935 14.2080 38.7175 ;
      RECT 13.8120 36.4855 13.8360 36.5095 ;
      RECT 13.8120 36.6775 13.8360 36.7015 ;
  LAYER M5  ;
      RECT 17.9160 35.5145 17.9400 36.6015 ;
      RECT 17.7475 35.9120 17.7715 36.9725 ;
      RECT 17.1135 35.9160 17.1375 36.7870 ;
      RECT 16.5120 36.6665 16.5360 36.8895 ;
      RECT 16.5120 37.8665 16.5360 38.0085 ;
      RECT 16.2960 36.1865 16.3200 37.2735 ;
      RECT 16.2960 37.5305 16.3200 37.7055 ;
      RECT 16.2960 38.0435 16.3200 38.2965 ;
      RECT 16.1270 34.8915 16.1510 38.7355 ;
      RECT 16.0800 36.0905 16.1040 37.3695 ;
      RECT 16.0800 37.5785 16.1040 37.7685 ;
      RECT 16.0800 37.9625 16.1040 38.2965 ;
      RECT 15.9720 38.6825 15.9960 39.1125 ;
      RECT 15.9720 41.3225 15.9960 41.4645 ;
      RECT 15.8820 34.1610 15.9060 43.6625 ;
      RECT 15.8340 34.1610 15.8580 43.6615 ;
      RECT 15.7860 34.1610 15.8100 43.6615 ;
      RECT 15.7380 34.1610 15.7620 43.6325 ;
      RECT 15.6900 34.1610 15.7140 43.6295 ;
      RECT 15.6420 34.1610 15.6660 43.6315 ;
      RECT 15.5940 34.1610 15.6180 43.6245 ;
      RECT 15.5460 34.1610 15.5700 43.6405 ;
      RECT 15.4980 34.1610 15.5220 43.6395 ;
      RECT 15.2100 34.3665 15.2340 43.6955 ;
      RECT 15.1620 34.3675 15.1860 43.6965 ;
      RECT 15.1140 34.3665 15.1380 43.6955 ;
      RECT 15.0180 34.3825 15.0420 43.6965 ;
      RECT 14.8260 34.3815 14.8500 43.6495 ;
      RECT 14.7780 34.3815 14.8020 43.6495 ;
      RECT 14.7300 34.3815 14.7540 43.6495 ;
      RECT 14.6820 34.3815 14.7060 43.6495 ;
      RECT 14.6340 34.3815 14.6580 43.6495 ;
      RECT 14.5860 34.3525 14.6100 43.6495 ;
      RECT 14.5380 34.3085 14.5620 43.3635 ;
      RECT 14.4900 34.2715 14.5140 43.3175 ;
      RECT 14.4420 34.2175 14.4660 43.2635 ;
      RECT 14.3520 39.1625 14.3760 39.3045 ;
      RECT 14.2440 37.0985 14.2680 38.1855 ;
      RECT 14.1840 34.8915 14.2080 38.7355 ;
      RECT 13.8120 36.4745 13.8360 36.7125 ;
  LAYER M2  ;
    RECT 0.108 0.036 30.2400 77.7240 ;
  LAYER M1  ;
    RECT 0.108 0.036 30.2400 77.7240 ;
  END
END srambank_256x4x64_6t122 
