VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_64x4x80_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_64x4x80_6t122 0 0 ; 
  SIZE 38.448 BY 380.16 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.688 38.036 4.88 ; 
        RECT 0.404 9.008 38.036 9.2 ; 
        RECT 0.404 13.328 38.036 13.52 ; 
        RECT 0.404 17.648 38.036 17.84 ; 
        RECT 0.404 21.968 38.036 22.16 ; 
        RECT 0.404 26.288 38.036 26.48 ; 
        RECT 0.404 30.608 38.036 30.8 ; 
        RECT 0.404 34.928 38.036 35.12 ; 
        RECT 0.404 39.248 38.036 39.44 ; 
        RECT 0.404 43.568 38.036 43.76 ; 
        RECT 0.404 47.888 38.036 48.08 ; 
        RECT 0.404 52.208 38.036 52.4 ; 
        RECT 0.404 56.528 38.036 56.72 ; 
        RECT 0.404 60.848 38.036 61.04 ; 
        RECT 0.404 65.168 38.036 65.36 ; 
        RECT 0.404 69.488 38.036 69.68 ; 
        RECT 0.404 73.808 38.036 74 ; 
        RECT 0.404 78.128 38.036 78.32 ; 
        RECT 0.404 82.448 38.036 82.64 ; 
        RECT 0.404 86.768 38.036 86.96 ; 
        RECT 0.404 91.088 38.036 91.28 ; 
        RECT 0.404 95.408 38.036 95.6 ; 
        RECT 0.404 99.728 38.036 99.92 ; 
        RECT 0.404 104.048 38.036 104.24 ; 
        RECT 0.404 108.368 38.036 108.56 ; 
        RECT 0.404 112.688 38.036 112.88 ; 
        RECT 0.404 117.008 38.036 117.2 ; 
        RECT 0.404 121.328 38.036 121.52 ; 
        RECT 0.404 125.648 38.036 125.84 ; 
        RECT 0.404 129.968 38.036 130.16 ; 
        RECT 0.404 134.288 38.036 134.48 ; 
        RECT 0.404 138.608 38.036 138.8 ; 
        RECT 0.404 142.928 38.036 143.12 ; 
        RECT 0.404 147.248 38.036 147.44 ; 
        RECT 0.404 151.568 38.036 151.76 ; 
        RECT 0.404 155.888 38.036 156.08 ; 
        RECT 0.404 160.208 38.036 160.4 ; 
        RECT 0.404 164.528 38.036 164.72 ; 
        RECT 0.404 168.848 38.036 169.04 ; 
        RECT 0.404 173.168 38.036 173.36 ; 
        RECT 0.432 175.116 38.016 175.98 ; 
        RECT 22.44 173.996 23.492 174.092 ; 
        RECT 22.964 189.132 23.412 189.228 ; 
        RECT 15.768 187.788 22.68 188.652 ; 
        RECT 15.768 200.46 22.68 201.324 ; 
        RECT 0.404 209.996 38.036 210.188 ; 
        RECT 0.404 214.316 38.036 214.508 ; 
        RECT 0.404 218.636 38.036 218.828 ; 
        RECT 0.404 222.956 38.036 223.148 ; 
        RECT 0.404 227.276 38.036 227.468 ; 
        RECT 0.404 231.596 38.036 231.788 ; 
        RECT 0.404 235.916 38.036 236.108 ; 
        RECT 0.404 240.236 38.036 240.428 ; 
        RECT 0.404 244.556 38.036 244.748 ; 
        RECT 0.404 248.876 38.036 249.068 ; 
        RECT 0.404 253.196 38.036 253.388 ; 
        RECT 0.404 257.516 38.036 257.708 ; 
        RECT 0.404 261.836 38.036 262.028 ; 
        RECT 0.404 266.156 38.036 266.348 ; 
        RECT 0.404 270.476 38.036 270.668 ; 
        RECT 0.404 274.796 38.036 274.988 ; 
        RECT 0.404 279.116 38.036 279.308 ; 
        RECT 0.404 283.436 38.036 283.628 ; 
        RECT 0.404 287.756 38.036 287.948 ; 
        RECT 0.404 292.076 38.036 292.268 ; 
        RECT 0.404 296.396 38.036 296.588 ; 
        RECT 0.404 300.716 38.036 300.908 ; 
        RECT 0.404 305.036 38.036 305.228 ; 
        RECT 0.404 309.356 38.036 309.548 ; 
        RECT 0.404 313.676 38.036 313.868 ; 
        RECT 0.404 317.996 38.036 318.188 ; 
        RECT 0.404 322.316 38.036 322.508 ; 
        RECT 0.404 326.636 38.036 326.828 ; 
        RECT 0.404 330.956 38.036 331.148 ; 
        RECT 0.404 335.276 38.036 335.468 ; 
        RECT 0.404 339.596 38.036 339.788 ; 
        RECT 0.404 343.916 38.036 344.108 ; 
        RECT 0.404 348.236 38.036 348.428 ; 
        RECT 0.404 352.556 38.036 352.748 ; 
        RECT 0.404 356.876 38.036 357.068 ; 
        RECT 0.404 361.196 38.036 361.388 ; 
        RECT 0.404 365.516 38.036 365.708 ; 
        RECT 0.404 369.836 38.036 370.028 ; 
        RECT 0.404 374.156 38.036 374.348 ; 
        RECT 0.404 378.476 38.036 378.668 ; 
      LAYER M3 ; 
        RECT 37.908 0.866 37.98 5.506 ; 
        RECT 23.292 0.868 23.364 5.504 ; 
        RECT 17.676 1.012 18.036 5.468 ; 
        RECT 15.084 0.868 15.156 5.504 ; 
        RECT 0.468 0.866 0.54 5.506 ; 
        RECT 37.908 5.186 37.98 9.826 ; 
        RECT 23.292 5.188 23.364 9.824 ; 
        RECT 17.676 5.332 18.036 9.788 ; 
        RECT 15.084 5.188 15.156 9.824 ; 
        RECT 0.468 5.186 0.54 9.826 ; 
        RECT 37.908 9.506 37.98 14.146 ; 
        RECT 23.292 9.508 23.364 14.144 ; 
        RECT 17.676 9.652 18.036 14.108 ; 
        RECT 15.084 9.508 15.156 14.144 ; 
        RECT 0.468 9.506 0.54 14.146 ; 
        RECT 37.908 13.826 37.98 18.466 ; 
        RECT 23.292 13.828 23.364 18.464 ; 
        RECT 17.676 13.972 18.036 18.428 ; 
        RECT 15.084 13.828 15.156 18.464 ; 
        RECT 0.468 13.826 0.54 18.466 ; 
        RECT 37.908 18.146 37.98 22.786 ; 
        RECT 23.292 18.148 23.364 22.784 ; 
        RECT 17.676 18.292 18.036 22.748 ; 
        RECT 15.084 18.148 15.156 22.784 ; 
        RECT 0.468 18.146 0.54 22.786 ; 
        RECT 37.908 22.466 37.98 27.106 ; 
        RECT 23.292 22.468 23.364 27.104 ; 
        RECT 17.676 22.612 18.036 27.068 ; 
        RECT 15.084 22.468 15.156 27.104 ; 
        RECT 0.468 22.466 0.54 27.106 ; 
        RECT 37.908 26.786 37.98 31.426 ; 
        RECT 23.292 26.788 23.364 31.424 ; 
        RECT 17.676 26.932 18.036 31.388 ; 
        RECT 15.084 26.788 15.156 31.424 ; 
        RECT 0.468 26.786 0.54 31.426 ; 
        RECT 37.908 31.106 37.98 35.746 ; 
        RECT 23.292 31.108 23.364 35.744 ; 
        RECT 17.676 31.252 18.036 35.708 ; 
        RECT 15.084 31.108 15.156 35.744 ; 
        RECT 0.468 31.106 0.54 35.746 ; 
        RECT 37.908 35.426 37.98 40.066 ; 
        RECT 23.292 35.428 23.364 40.064 ; 
        RECT 17.676 35.572 18.036 40.028 ; 
        RECT 15.084 35.428 15.156 40.064 ; 
        RECT 0.468 35.426 0.54 40.066 ; 
        RECT 37.908 39.746 37.98 44.386 ; 
        RECT 23.292 39.748 23.364 44.384 ; 
        RECT 17.676 39.892 18.036 44.348 ; 
        RECT 15.084 39.748 15.156 44.384 ; 
        RECT 0.468 39.746 0.54 44.386 ; 
        RECT 37.908 44.066 37.98 48.706 ; 
        RECT 23.292 44.068 23.364 48.704 ; 
        RECT 17.676 44.212 18.036 48.668 ; 
        RECT 15.084 44.068 15.156 48.704 ; 
        RECT 0.468 44.066 0.54 48.706 ; 
        RECT 37.908 48.386 37.98 53.026 ; 
        RECT 23.292 48.388 23.364 53.024 ; 
        RECT 17.676 48.532 18.036 52.988 ; 
        RECT 15.084 48.388 15.156 53.024 ; 
        RECT 0.468 48.386 0.54 53.026 ; 
        RECT 37.908 52.706 37.98 57.346 ; 
        RECT 23.292 52.708 23.364 57.344 ; 
        RECT 17.676 52.852 18.036 57.308 ; 
        RECT 15.084 52.708 15.156 57.344 ; 
        RECT 0.468 52.706 0.54 57.346 ; 
        RECT 37.908 57.026 37.98 61.666 ; 
        RECT 23.292 57.028 23.364 61.664 ; 
        RECT 17.676 57.172 18.036 61.628 ; 
        RECT 15.084 57.028 15.156 61.664 ; 
        RECT 0.468 57.026 0.54 61.666 ; 
        RECT 37.908 61.346 37.98 65.986 ; 
        RECT 23.292 61.348 23.364 65.984 ; 
        RECT 17.676 61.492 18.036 65.948 ; 
        RECT 15.084 61.348 15.156 65.984 ; 
        RECT 0.468 61.346 0.54 65.986 ; 
        RECT 37.908 65.666 37.98 70.306 ; 
        RECT 23.292 65.668 23.364 70.304 ; 
        RECT 17.676 65.812 18.036 70.268 ; 
        RECT 15.084 65.668 15.156 70.304 ; 
        RECT 0.468 65.666 0.54 70.306 ; 
        RECT 37.908 69.986 37.98 74.626 ; 
        RECT 23.292 69.988 23.364 74.624 ; 
        RECT 17.676 70.132 18.036 74.588 ; 
        RECT 15.084 69.988 15.156 74.624 ; 
        RECT 0.468 69.986 0.54 74.626 ; 
        RECT 37.908 74.306 37.98 78.946 ; 
        RECT 23.292 74.308 23.364 78.944 ; 
        RECT 17.676 74.452 18.036 78.908 ; 
        RECT 15.084 74.308 15.156 78.944 ; 
        RECT 0.468 74.306 0.54 78.946 ; 
        RECT 37.908 78.626 37.98 83.266 ; 
        RECT 23.292 78.628 23.364 83.264 ; 
        RECT 17.676 78.772 18.036 83.228 ; 
        RECT 15.084 78.628 15.156 83.264 ; 
        RECT 0.468 78.626 0.54 83.266 ; 
        RECT 37.908 82.946 37.98 87.586 ; 
        RECT 23.292 82.948 23.364 87.584 ; 
        RECT 17.676 83.092 18.036 87.548 ; 
        RECT 15.084 82.948 15.156 87.584 ; 
        RECT 0.468 82.946 0.54 87.586 ; 
        RECT 37.908 87.266 37.98 91.906 ; 
        RECT 23.292 87.268 23.364 91.904 ; 
        RECT 17.676 87.412 18.036 91.868 ; 
        RECT 15.084 87.268 15.156 91.904 ; 
        RECT 0.468 87.266 0.54 91.906 ; 
        RECT 37.908 91.586 37.98 96.226 ; 
        RECT 23.292 91.588 23.364 96.224 ; 
        RECT 17.676 91.732 18.036 96.188 ; 
        RECT 15.084 91.588 15.156 96.224 ; 
        RECT 0.468 91.586 0.54 96.226 ; 
        RECT 37.908 95.906 37.98 100.546 ; 
        RECT 23.292 95.908 23.364 100.544 ; 
        RECT 17.676 96.052 18.036 100.508 ; 
        RECT 15.084 95.908 15.156 100.544 ; 
        RECT 0.468 95.906 0.54 100.546 ; 
        RECT 37.908 100.226 37.98 104.866 ; 
        RECT 23.292 100.228 23.364 104.864 ; 
        RECT 17.676 100.372 18.036 104.828 ; 
        RECT 15.084 100.228 15.156 104.864 ; 
        RECT 0.468 100.226 0.54 104.866 ; 
        RECT 37.908 104.546 37.98 109.186 ; 
        RECT 23.292 104.548 23.364 109.184 ; 
        RECT 17.676 104.692 18.036 109.148 ; 
        RECT 15.084 104.548 15.156 109.184 ; 
        RECT 0.468 104.546 0.54 109.186 ; 
        RECT 37.908 108.866 37.98 113.506 ; 
        RECT 23.292 108.868 23.364 113.504 ; 
        RECT 17.676 109.012 18.036 113.468 ; 
        RECT 15.084 108.868 15.156 113.504 ; 
        RECT 0.468 108.866 0.54 113.506 ; 
        RECT 37.908 113.186 37.98 117.826 ; 
        RECT 23.292 113.188 23.364 117.824 ; 
        RECT 17.676 113.332 18.036 117.788 ; 
        RECT 15.084 113.188 15.156 117.824 ; 
        RECT 0.468 113.186 0.54 117.826 ; 
        RECT 37.908 117.506 37.98 122.146 ; 
        RECT 23.292 117.508 23.364 122.144 ; 
        RECT 17.676 117.652 18.036 122.108 ; 
        RECT 15.084 117.508 15.156 122.144 ; 
        RECT 0.468 117.506 0.54 122.146 ; 
        RECT 37.908 121.826 37.98 126.466 ; 
        RECT 23.292 121.828 23.364 126.464 ; 
        RECT 17.676 121.972 18.036 126.428 ; 
        RECT 15.084 121.828 15.156 126.464 ; 
        RECT 0.468 121.826 0.54 126.466 ; 
        RECT 37.908 126.146 37.98 130.786 ; 
        RECT 23.292 126.148 23.364 130.784 ; 
        RECT 17.676 126.292 18.036 130.748 ; 
        RECT 15.084 126.148 15.156 130.784 ; 
        RECT 0.468 126.146 0.54 130.786 ; 
        RECT 37.908 130.466 37.98 135.106 ; 
        RECT 23.292 130.468 23.364 135.104 ; 
        RECT 17.676 130.612 18.036 135.068 ; 
        RECT 15.084 130.468 15.156 135.104 ; 
        RECT 0.468 130.466 0.54 135.106 ; 
        RECT 37.908 134.786 37.98 139.426 ; 
        RECT 23.292 134.788 23.364 139.424 ; 
        RECT 17.676 134.932 18.036 139.388 ; 
        RECT 15.084 134.788 15.156 139.424 ; 
        RECT 0.468 134.786 0.54 139.426 ; 
        RECT 37.908 139.106 37.98 143.746 ; 
        RECT 23.292 139.108 23.364 143.744 ; 
        RECT 17.676 139.252 18.036 143.708 ; 
        RECT 15.084 139.108 15.156 143.744 ; 
        RECT 0.468 139.106 0.54 143.746 ; 
        RECT 37.908 143.426 37.98 148.066 ; 
        RECT 23.292 143.428 23.364 148.064 ; 
        RECT 17.676 143.572 18.036 148.028 ; 
        RECT 15.084 143.428 15.156 148.064 ; 
        RECT 0.468 143.426 0.54 148.066 ; 
        RECT 37.908 147.746 37.98 152.386 ; 
        RECT 23.292 147.748 23.364 152.384 ; 
        RECT 17.676 147.892 18.036 152.348 ; 
        RECT 15.084 147.748 15.156 152.384 ; 
        RECT 0.468 147.746 0.54 152.386 ; 
        RECT 37.908 152.066 37.98 156.706 ; 
        RECT 23.292 152.068 23.364 156.704 ; 
        RECT 17.676 152.212 18.036 156.668 ; 
        RECT 15.084 152.068 15.156 156.704 ; 
        RECT 0.468 152.066 0.54 156.706 ; 
        RECT 37.908 156.386 37.98 161.026 ; 
        RECT 23.292 156.388 23.364 161.024 ; 
        RECT 17.676 156.532 18.036 160.988 ; 
        RECT 15.084 156.388 15.156 161.024 ; 
        RECT 0.468 156.386 0.54 161.026 ; 
        RECT 37.908 160.706 37.98 165.346 ; 
        RECT 23.292 160.708 23.364 165.344 ; 
        RECT 17.676 160.852 18.036 165.308 ; 
        RECT 15.084 160.708 15.156 165.344 ; 
        RECT 0.468 160.706 0.54 165.346 ; 
        RECT 37.908 165.026 37.98 169.666 ; 
        RECT 23.292 165.028 23.364 169.664 ; 
        RECT 17.676 165.172 18.036 169.628 ; 
        RECT 15.084 165.028 15.156 169.664 ; 
        RECT 0.468 165.026 0.54 169.666 ; 
        RECT 37.908 169.346 37.98 173.986 ; 
        RECT 23.292 169.348 23.364 173.984 ; 
        RECT 17.676 169.492 18.036 173.948 ; 
        RECT 15.084 169.348 15.156 173.984 ; 
        RECT 0.468 169.346 0.54 173.986 ; 
        RECT 37.908 173.666 37.98 206.494 ; 
        RECT 23.292 173.984 23.364 174.35 ; 
        RECT 23.292 188.944 23.364 206.384 ; 
        RECT 17.82 174.96 18.756 205.292 ; 
        RECT 17.676 204.948 18.036 207.088 ; 
        RECT 17.676 173.84 18.036 175.98 ; 
        RECT 0.468 173.666 0.54 206.494 ; 
        RECT 37.908 206.174 37.98 210.814 ; 
        RECT 23.292 206.176 23.364 210.812 ; 
        RECT 17.676 206.32 18.036 210.776 ; 
        RECT 15.084 206.176 15.156 210.812 ; 
        RECT 0.468 206.174 0.54 210.814 ; 
        RECT 37.908 210.494 37.98 215.134 ; 
        RECT 23.292 210.496 23.364 215.132 ; 
        RECT 17.676 210.64 18.036 215.096 ; 
        RECT 15.084 210.496 15.156 215.132 ; 
        RECT 0.468 210.494 0.54 215.134 ; 
        RECT 37.908 214.814 37.98 219.454 ; 
        RECT 23.292 214.816 23.364 219.452 ; 
        RECT 17.676 214.96 18.036 219.416 ; 
        RECT 15.084 214.816 15.156 219.452 ; 
        RECT 0.468 214.814 0.54 219.454 ; 
        RECT 37.908 219.134 37.98 223.774 ; 
        RECT 23.292 219.136 23.364 223.772 ; 
        RECT 17.676 219.28 18.036 223.736 ; 
        RECT 15.084 219.136 15.156 223.772 ; 
        RECT 0.468 219.134 0.54 223.774 ; 
        RECT 37.908 223.454 37.98 228.094 ; 
        RECT 23.292 223.456 23.364 228.092 ; 
        RECT 17.676 223.6 18.036 228.056 ; 
        RECT 15.084 223.456 15.156 228.092 ; 
        RECT 0.468 223.454 0.54 228.094 ; 
        RECT 37.908 227.774 37.98 232.414 ; 
        RECT 23.292 227.776 23.364 232.412 ; 
        RECT 17.676 227.92 18.036 232.376 ; 
        RECT 15.084 227.776 15.156 232.412 ; 
        RECT 0.468 227.774 0.54 232.414 ; 
        RECT 37.908 232.094 37.98 236.734 ; 
        RECT 23.292 232.096 23.364 236.732 ; 
        RECT 17.676 232.24 18.036 236.696 ; 
        RECT 15.084 232.096 15.156 236.732 ; 
        RECT 0.468 232.094 0.54 236.734 ; 
        RECT 37.908 236.414 37.98 241.054 ; 
        RECT 23.292 236.416 23.364 241.052 ; 
        RECT 17.676 236.56 18.036 241.016 ; 
        RECT 15.084 236.416 15.156 241.052 ; 
        RECT 0.468 236.414 0.54 241.054 ; 
        RECT 37.908 240.734 37.98 245.374 ; 
        RECT 23.292 240.736 23.364 245.372 ; 
        RECT 17.676 240.88 18.036 245.336 ; 
        RECT 15.084 240.736 15.156 245.372 ; 
        RECT 0.468 240.734 0.54 245.374 ; 
        RECT 37.908 245.054 37.98 249.694 ; 
        RECT 23.292 245.056 23.364 249.692 ; 
        RECT 17.676 245.2 18.036 249.656 ; 
        RECT 15.084 245.056 15.156 249.692 ; 
        RECT 0.468 245.054 0.54 249.694 ; 
        RECT 37.908 249.374 37.98 254.014 ; 
        RECT 23.292 249.376 23.364 254.012 ; 
        RECT 17.676 249.52 18.036 253.976 ; 
        RECT 15.084 249.376 15.156 254.012 ; 
        RECT 0.468 249.374 0.54 254.014 ; 
        RECT 37.908 253.694 37.98 258.334 ; 
        RECT 23.292 253.696 23.364 258.332 ; 
        RECT 17.676 253.84 18.036 258.296 ; 
        RECT 15.084 253.696 15.156 258.332 ; 
        RECT 0.468 253.694 0.54 258.334 ; 
        RECT 37.908 258.014 37.98 262.654 ; 
        RECT 23.292 258.016 23.364 262.652 ; 
        RECT 17.676 258.16 18.036 262.616 ; 
        RECT 15.084 258.016 15.156 262.652 ; 
        RECT 0.468 258.014 0.54 262.654 ; 
        RECT 37.908 262.334 37.98 266.974 ; 
        RECT 23.292 262.336 23.364 266.972 ; 
        RECT 17.676 262.48 18.036 266.936 ; 
        RECT 15.084 262.336 15.156 266.972 ; 
        RECT 0.468 262.334 0.54 266.974 ; 
        RECT 37.908 266.654 37.98 271.294 ; 
        RECT 23.292 266.656 23.364 271.292 ; 
        RECT 17.676 266.8 18.036 271.256 ; 
        RECT 15.084 266.656 15.156 271.292 ; 
        RECT 0.468 266.654 0.54 271.294 ; 
        RECT 37.908 270.974 37.98 275.614 ; 
        RECT 23.292 270.976 23.364 275.612 ; 
        RECT 17.676 271.12 18.036 275.576 ; 
        RECT 15.084 270.976 15.156 275.612 ; 
        RECT 0.468 270.974 0.54 275.614 ; 
        RECT 37.908 275.294 37.98 279.934 ; 
        RECT 23.292 275.296 23.364 279.932 ; 
        RECT 17.676 275.44 18.036 279.896 ; 
        RECT 15.084 275.296 15.156 279.932 ; 
        RECT 0.468 275.294 0.54 279.934 ; 
        RECT 37.908 279.614 37.98 284.254 ; 
        RECT 23.292 279.616 23.364 284.252 ; 
        RECT 17.676 279.76 18.036 284.216 ; 
        RECT 15.084 279.616 15.156 284.252 ; 
        RECT 0.468 279.614 0.54 284.254 ; 
        RECT 37.908 283.934 37.98 288.574 ; 
        RECT 23.292 283.936 23.364 288.572 ; 
        RECT 17.676 284.08 18.036 288.536 ; 
        RECT 15.084 283.936 15.156 288.572 ; 
        RECT 0.468 283.934 0.54 288.574 ; 
        RECT 37.908 288.254 37.98 292.894 ; 
        RECT 23.292 288.256 23.364 292.892 ; 
        RECT 17.676 288.4 18.036 292.856 ; 
        RECT 15.084 288.256 15.156 292.892 ; 
        RECT 0.468 288.254 0.54 292.894 ; 
        RECT 37.908 292.574 37.98 297.214 ; 
        RECT 23.292 292.576 23.364 297.212 ; 
        RECT 17.676 292.72 18.036 297.176 ; 
        RECT 15.084 292.576 15.156 297.212 ; 
        RECT 0.468 292.574 0.54 297.214 ; 
        RECT 37.908 296.894 37.98 301.534 ; 
        RECT 23.292 296.896 23.364 301.532 ; 
        RECT 17.676 297.04 18.036 301.496 ; 
        RECT 15.084 296.896 15.156 301.532 ; 
        RECT 0.468 296.894 0.54 301.534 ; 
        RECT 37.908 301.214 37.98 305.854 ; 
        RECT 23.292 301.216 23.364 305.852 ; 
        RECT 17.676 301.36 18.036 305.816 ; 
        RECT 15.084 301.216 15.156 305.852 ; 
        RECT 0.468 301.214 0.54 305.854 ; 
        RECT 37.908 305.534 37.98 310.174 ; 
        RECT 23.292 305.536 23.364 310.172 ; 
        RECT 17.676 305.68 18.036 310.136 ; 
        RECT 15.084 305.536 15.156 310.172 ; 
        RECT 0.468 305.534 0.54 310.174 ; 
        RECT 37.908 309.854 37.98 314.494 ; 
        RECT 23.292 309.856 23.364 314.492 ; 
        RECT 17.676 310 18.036 314.456 ; 
        RECT 15.084 309.856 15.156 314.492 ; 
        RECT 0.468 309.854 0.54 314.494 ; 
        RECT 37.908 314.174 37.98 318.814 ; 
        RECT 23.292 314.176 23.364 318.812 ; 
        RECT 17.676 314.32 18.036 318.776 ; 
        RECT 15.084 314.176 15.156 318.812 ; 
        RECT 0.468 314.174 0.54 318.814 ; 
        RECT 37.908 318.494 37.98 323.134 ; 
        RECT 23.292 318.496 23.364 323.132 ; 
        RECT 17.676 318.64 18.036 323.096 ; 
        RECT 15.084 318.496 15.156 323.132 ; 
        RECT 0.468 318.494 0.54 323.134 ; 
        RECT 37.908 322.814 37.98 327.454 ; 
        RECT 23.292 322.816 23.364 327.452 ; 
        RECT 17.676 322.96 18.036 327.416 ; 
        RECT 15.084 322.816 15.156 327.452 ; 
        RECT 0.468 322.814 0.54 327.454 ; 
        RECT 37.908 327.134 37.98 331.774 ; 
        RECT 23.292 327.136 23.364 331.772 ; 
        RECT 17.676 327.28 18.036 331.736 ; 
        RECT 15.084 327.136 15.156 331.772 ; 
        RECT 0.468 327.134 0.54 331.774 ; 
        RECT 37.908 331.454 37.98 336.094 ; 
        RECT 23.292 331.456 23.364 336.092 ; 
        RECT 17.676 331.6 18.036 336.056 ; 
        RECT 15.084 331.456 15.156 336.092 ; 
        RECT 0.468 331.454 0.54 336.094 ; 
        RECT 37.908 335.774 37.98 340.414 ; 
        RECT 23.292 335.776 23.364 340.412 ; 
        RECT 17.676 335.92 18.036 340.376 ; 
        RECT 15.084 335.776 15.156 340.412 ; 
        RECT 0.468 335.774 0.54 340.414 ; 
        RECT 37.908 340.094 37.98 344.734 ; 
        RECT 23.292 340.096 23.364 344.732 ; 
        RECT 17.676 340.24 18.036 344.696 ; 
        RECT 15.084 340.096 15.156 344.732 ; 
        RECT 0.468 340.094 0.54 344.734 ; 
        RECT 37.908 344.414 37.98 349.054 ; 
        RECT 23.292 344.416 23.364 349.052 ; 
        RECT 17.676 344.56 18.036 349.016 ; 
        RECT 15.084 344.416 15.156 349.052 ; 
        RECT 0.468 344.414 0.54 349.054 ; 
        RECT 37.908 348.734 37.98 353.374 ; 
        RECT 23.292 348.736 23.364 353.372 ; 
        RECT 17.676 348.88 18.036 353.336 ; 
        RECT 15.084 348.736 15.156 353.372 ; 
        RECT 0.468 348.734 0.54 353.374 ; 
        RECT 37.908 353.054 37.98 357.694 ; 
        RECT 23.292 353.056 23.364 357.692 ; 
        RECT 17.676 353.2 18.036 357.656 ; 
        RECT 15.084 353.056 15.156 357.692 ; 
        RECT 0.468 353.054 0.54 357.694 ; 
        RECT 37.908 357.374 37.98 362.014 ; 
        RECT 23.292 357.376 23.364 362.012 ; 
        RECT 17.676 357.52 18.036 361.976 ; 
        RECT 15.084 357.376 15.156 362.012 ; 
        RECT 0.468 357.374 0.54 362.014 ; 
        RECT 37.908 361.694 37.98 366.334 ; 
        RECT 23.292 361.696 23.364 366.332 ; 
        RECT 17.676 361.84 18.036 366.296 ; 
        RECT 15.084 361.696 15.156 366.332 ; 
        RECT 0.468 361.694 0.54 366.334 ; 
        RECT 37.908 366.014 37.98 370.654 ; 
        RECT 23.292 366.016 23.364 370.652 ; 
        RECT 17.676 366.16 18.036 370.616 ; 
        RECT 15.084 366.016 15.156 370.652 ; 
        RECT 0.468 366.014 0.54 370.654 ; 
        RECT 37.908 370.334 37.98 374.974 ; 
        RECT 23.292 370.336 23.364 374.972 ; 
        RECT 17.676 370.48 18.036 374.936 ; 
        RECT 15.084 370.336 15.156 374.972 ; 
        RECT 0.468 370.334 0.54 374.974 ; 
        RECT 37.908 374.654 37.98 379.294 ; 
        RECT 23.292 374.656 23.364 379.292 ; 
        RECT 17.676 374.8 18.036 379.256 ; 
        RECT 15.084 374.656 15.156 379.292 ; 
        RECT 0.468 374.654 0.54 379.294 ; 
      LAYER V3 ; 
        RECT 0.468 4.688 0.54 4.88 ; 
        RECT 15.084 4.688 15.156 4.88 ; 
        RECT 17.676 4.688 18.036 4.88 ; 
        RECT 23.292 4.688 23.364 4.88 ; 
        RECT 37.908 4.688 37.98 4.88 ; 
        RECT 0.468 9.008 0.54 9.2 ; 
        RECT 15.084 9.008 15.156 9.2 ; 
        RECT 17.676 9.008 18.036 9.2 ; 
        RECT 23.292 9.008 23.364 9.2 ; 
        RECT 37.908 9.008 37.98 9.2 ; 
        RECT 0.468 13.328 0.54 13.52 ; 
        RECT 15.084 13.328 15.156 13.52 ; 
        RECT 17.676 13.328 18.036 13.52 ; 
        RECT 23.292 13.328 23.364 13.52 ; 
        RECT 37.908 13.328 37.98 13.52 ; 
        RECT 0.468 17.648 0.54 17.84 ; 
        RECT 15.084 17.648 15.156 17.84 ; 
        RECT 17.676 17.648 18.036 17.84 ; 
        RECT 23.292 17.648 23.364 17.84 ; 
        RECT 37.908 17.648 37.98 17.84 ; 
        RECT 0.468 21.968 0.54 22.16 ; 
        RECT 15.084 21.968 15.156 22.16 ; 
        RECT 17.676 21.968 18.036 22.16 ; 
        RECT 23.292 21.968 23.364 22.16 ; 
        RECT 37.908 21.968 37.98 22.16 ; 
        RECT 0.468 26.288 0.54 26.48 ; 
        RECT 15.084 26.288 15.156 26.48 ; 
        RECT 17.676 26.288 18.036 26.48 ; 
        RECT 23.292 26.288 23.364 26.48 ; 
        RECT 37.908 26.288 37.98 26.48 ; 
        RECT 0.468 30.608 0.54 30.8 ; 
        RECT 15.084 30.608 15.156 30.8 ; 
        RECT 17.676 30.608 18.036 30.8 ; 
        RECT 23.292 30.608 23.364 30.8 ; 
        RECT 37.908 30.608 37.98 30.8 ; 
        RECT 0.468 34.928 0.54 35.12 ; 
        RECT 15.084 34.928 15.156 35.12 ; 
        RECT 17.676 34.928 18.036 35.12 ; 
        RECT 23.292 34.928 23.364 35.12 ; 
        RECT 37.908 34.928 37.98 35.12 ; 
        RECT 0.468 39.248 0.54 39.44 ; 
        RECT 15.084 39.248 15.156 39.44 ; 
        RECT 17.676 39.248 18.036 39.44 ; 
        RECT 23.292 39.248 23.364 39.44 ; 
        RECT 37.908 39.248 37.98 39.44 ; 
        RECT 0.468 43.568 0.54 43.76 ; 
        RECT 15.084 43.568 15.156 43.76 ; 
        RECT 17.676 43.568 18.036 43.76 ; 
        RECT 23.292 43.568 23.364 43.76 ; 
        RECT 37.908 43.568 37.98 43.76 ; 
        RECT 0.468 47.888 0.54 48.08 ; 
        RECT 15.084 47.888 15.156 48.08 ; 
        RECT 17.676 47.888 18.036 48.08 ; 
        RECT 23.292 47.888 23.364 48.08 ; 
        RECT 37.908 47.888 37.98 48.08 ; 
        RECT 0.468 52.208 0.54 52.4 ; 
        RECT 15.084 52.208 15.156 52.4 ; 
        RECT 17.676 52.208 18.036 52.4 ; 
        RECT 23.292 52.208 23.364 52.4 ; 
        RECT 37.908 52.208 37.98 52.4 ; 
        RECT 0.468 56.528 0.54 56.72 ; 
        RECT 15.084 56.528 15.156 56.72 ; 
        RECT 17.676 56.528 18.036 56.72 ; 
        RECT 23.292 56.528 23.364 56.72 ; 
        RECT 37.908 56.528 37.98 56.72 ; 
        RECT 0.468 60.848 0.54 61.04 ; 
        RECT 15.084 60.848 15.156 61.04 ; 
        RECT 17.676 60.848 18.036 61.04 ; 
        RECT 23.292 60.848 23.364 61.04 ; 
        RECT 37.908 60.848 37.98 61.04 ; 
        RECT 0.468 65.168 0.54 65.36 ; 
        RECT 15.084 65.168 15.156 65.36 ; 
        RECT 17.676 65.168 18.036 65.36 ; 
        RECT 23.292 65.168 23.364 65.36 ; 
        RECT 37.908 65.168 37.98 65.36 ; 
        RECT 0.468 69.488 0.54 69.68 ; 
        RECT 15.084 69.488 15.156 69.68 ; 
        RECT 17.676 69.488 18.036 69.68 ; 
        RECT 23.292 69.488 23.364 69.68 ; 
        RECT 37.908 69.488 37.98 69.68 ; 
        RECT 0.468 73.808 0.54 74 ; 
        RECT 15.084 73.808 15.156 74 ; 
        RECT 17.676 73.808 18.036 74 ; 
        RECT 23.292 73.808 23.364 74 ; 
        RECT 37.908 73.808 37.98 74 ; 
        RECT 0.468 78.128 0.54 78.32 ; 
        RECT 15.084 78.128 15.156 78.32 ; 
        RECT 17.676 78.128 18.036 78.32 ; 
        RECT 23.292 78.128 23.364 78.32 ; 
        RECT 37.908 78.128 37.98 78.32 ; 
        RECT 0.468 82.448 0.54 82.64 ; 
        RECT 15.084 82.448 15.156 82.64 ; 
        RECT 17.676 82.448 18.036 82.64 ; 
        RECT 23.292 82.448 23.364 82.64 ; 
        RECT 37.908 82.448 37.98 82.64 ; 
        RECT 0.468 86.768 0.54 86.96 ; 
        RECT 15.084 86.768 15.156 86.96 ; 
        RECT 17.676 86.768 18.036 86.96 ; 
        RECT 23.292 86.768 23.364 86.96 ; 
        RECT 37.908 86.768 37.98 86.96 ; 
        RECT 0.468 91.088 0.54 91.28 ; 
        RECT 15.084 91.088 15.156 91.28 ; 
        RECT 17.676 91.088 18.036 91.28 ; 
        RECT 23.292 91.088 23.364 91.28 ; 
        RECT 37.908 91.088 37.98 91.28 ; 
        RECT 0.468 95.408 0.54 95.6 ; 
        RECT 15.084 95.408 15.156 95.6 ; 
        RECT 17.676 95.408 18.036 95.6 ; 
        RECT 23.292 95.408 23.364 95.6 ; 
        RECT 37.908 95.408 37.98 95.6 ; 
        RECT 0.468 99.728 0.54 99.92 ; 
        RECT 15.084 99.728 15.156 99.92 ; 
        RECT 17.676 99.728 18.036 99.92 ; 
        RECT 23.292 99.728 23.364 99.92 ; 
        RECT 37.908 99.728 37.98 99.92 ; 
        RECT 0.468 104.048 0.54 104.24 ; 
        RECT 15.084 104.048 15.156 104.24 ; 
        RECT 17.676 104.048 18.036 104.24 ; 
        RECT 23.292 104.048 23.364 104.24 ; 
        RECT 37.908 104.048 37.98 104.24 ; 
        RECT 0.468 108.368 0.54 108.56 ; 
        RECT 15.084 108.368 15.156 108.56 ; 
        RECT 17.676 108.368 18.036 108.56 ; 
        RECT 23.292 108.368 23.364 108.56 ; 
        RECT 37.908 108.368 37.98 108.56 ; 
        RECT 0.468 112.688 0.54 112.88 ; 
        RECT 15.084 112.688 15.156 112.88 ; 
        RECT 17.676 112.688 18.036 112.88 ; 
        RECT 23.292 112.688 23.364 112.88 ; 
        RECT 37.908 112.688 37.98 112.88 ; 
        RECT 0.468 117.008 0.54 117.2 ; 
        RECT 15.084 117.008 15.156 117.2 ; 
        RECT 17.676 117.008 18.036 117.2 ; 
        RECT 23.292 117.008 23.364 117.2 ; 
        RECT 37.908 117.008 37.98 117.2 ; 
        RECT 0.468 121.328 0.54 121.52 ; 
        RECT 15.084 121.328 15.156 121.52 ; 
        RECT 17.676 121.328 18.036 121.52 ; 
        RECT 23.292 121.328 23.364 121.52 ; 
        RECT 37.908 121.328 37.98 121.52 ; 
        RECT 0.468 125.648 0.54 125.84 ; 
        RECT 15.084 125.648 15.156 125.84 ; 
        RECT 17.676 125.648 18.036 125.84 ; 
        RECT 23.292 125.648 23.364 125.84 ; 
        RECT 37.908 125.648 37.98 125.84 ; 
        RECT 0.468 129.968 0.54 130.16 ; 
        RECT 15.084 129.968 15.156 130.16 ; 
        RECT 17.676 129.968 18.036 130.16 ; 
        RECT 23.292 129.968 23.364 130.16 ; 
        RECT 37.908 129.968 37.98 130.16 ; 
        RECT 0.468 134.288 0.54 134.48 ; 
        RECT 15.084 134.288 15.156 134.48 ; 
        RECT 17.676 134.288 18.036 134.48 ; 
        RECT 23.292 134.288 23.364 134.48 ; 
        RECT 37.908 134.288 37.98 134.48 ; 
        RECT 0.468 138.608 0.54 138.8 ; 
        RECT 15.084 138.608 15.156 138.8 ; 
        RECT 17.676 138.608 18.036 138.8 ; 
        RECT 23.292 138.608 23.364 138.8 ; 
        RECT 37.908 138.608 37.98 138.8 ; 
        RECT 0.468 142.928 0.54 143.12 ; 
        RECT 15.084 142.928 15.156 143.12 ; 
        RECT 17.676 142.928 18.036 143.12 ; 
        RECT 23.292 142.928 23.364 143.12 ; 
        RECT 37.908 142.928 37.98 143.12 ; 
        RECT 0.468 147.248 0.54 147.44 ; 
        RECT 15.084 147.248 15.156 147.44 ; 
        RECT 17.676 147.248 18.036 147.44 ; 
        RECT 23.292 147.248 23.364 147.44 ; 
        RECT 37.908 147.248 37.98 147.44 ; 
        RECT 0.468 151.568 0.54 151.76 ; 
        RECT 15.084 151.568 15.156 151.76 ; 
        RECT 17.676 151.568 18.036 151.76 ; 
        RECT 23.292 151.568 23.364 151.76 ; 
        RECT 37.908 151.568 37.98 151.76 ; 
        RECT 0.468 155.888 0.54 156.08 ; 
        RECT 15.084 155.888 15.156 156.08 ; 
        RECT 17.676 155.888 18.036 156.08 ; 
        RECT 23.292 155.888 23.364 156.08 ; 
        RECT 37.908 155.888 37.98 156.08 ; 
        RECT 0.468 160.208 0.54 160.4 ; 
        RECT 15.084 160.208 15.156 160.4 ; 
        RECT 17.676 160.208 18.036 160.4 ; 
        RECT 23.292 160.208 23.364 160.4 ; 
        RECT 37.908 160.208 37.98 160.4 ; 
        RECT 0.468 164.528 0.54 164.72 ; 
        RECT 15.084 164.528 15.156 164.72 ; 
        RECT 17.676 164.528 18.036 164.72 ; 
        RECT 23.292 164.528 23.364 164.72 ; 
        RECT 37.908 164.528 37.98 164.72 ; 
        RECT 0.468 168.848 0.54 169.04 ; 
        RECT 15.084 168.848 15.156 169.04 ; 
        RECT 17.676 168.848 18.036 169.04 ; 
        RECT 23.292 168.848 23.364 169.04 ; 
        RECT 37.908 168.848 37.98 169.04 ; 
        RECT 0.468 173.168 0.54 173.36 ; 
        RECT 15.084 173.168 15.156 173.36 ; 
        RECT 17.676 173.168 18.036 173.36 ; 
        RECT 23.292 173.168 23.364 173.36 ; 
        RECT 37.908 173.168 37.98 173.36 ; 
        RECT 0.468 175.116 0.54 175.98 ; 
        RECT 17.836 200.46 17.908 201.324 ; 
        RECT 17.836 187.788 17.908 188.652 ; 
        RECT 17.836 175.116 17.908 175.98 ; 
        RECT 18.044 200.46 18.116 201.324 ; 
        RECT 18.044 187.788 18.116 188.652 ; 
        RECT 18.044 175.116 18.116 175.98 ; 
        RECT 18.252 200.46 18.324 201.324 ; 
        RECT 18.252 187.788 18.324 188.652 ; 
        RECT 18.252 175.116 18.324 175.98 ; 
        RECT 18.46 200.46 18.532 201.324 ; 
        RECT 18.46 187.788 18.532 188.652 ; 
        RECT 18.46 175.116 18.532 175.98 ; 
        RECT 18.668 200.46 18.74 201.324 ; 
        RECT 18.668 187.788 18.74 188.652 ; 
        RECT 18.668 175.116 18.74 175.98 ; 
        RECT 23.292 189.132 23.364 189.228 ; 
        RECT 23.292 173.996 23.364 174.092 ; 
        RECT 0.468 209.996 0.54 210.188 ; 
        RECT 15.084 209.996 15.156 210.188 ; 
        RECT 17.676 209.996 18.036 210.188 ; 
        RECT 23.292 209.996 23.364 210.188 ; 
        RECT 37.908 209.996 37.98 210.188 ; 
        RECT 0.468 214.316 0.54 214.508 ; 
        RECT 15.084 214.316 15.156 214.508 ; 
        RECT 17.676 214.316 18.036 214.508 ; 
        RECT 23.292 214.316 23.364 214.508 ; 
        RECT 37.908 214.316 37.98 214.508 ; 
        RECT 0.468 218.636 0.54 218.828 ; 
        RECT 15.084 218.636 15.156 218.828 ; 
        RECT 17.676 218.636 18.036 218.828 ; 
        RECT 23.292 218.636 23.364 218.828 ; 
        RECT 37.908 218.636 37.98 218.828 ; 
        RECT 0.468 222.956 0.54 223.148 ; 
        RECT 15.084 222.956 15.156 223.148 ; 
        RECT 17.676 222.956 18.036 223.148 ; 
        RECT 23.292 222.956 23.364 223.148 ; 
        RECT 37.908 222.956 37.98 223.148 ; 
        RECT 0.468 227.276 0.54 227.468 ; 
        RECT 15.084 227.276 15.156 227.468 ; 
        RECT 17.676 227.276 18.036 227.468 ; 
        RECT 23.292 227.276 23.364 227.468 ; 
        RECT 37.908 227.276 37.98 227.468 ; 
        RECT 0.468 231.596 0.54 231.788 ; 
        RECT 15.084 231.596 15.156 231.788 ; 
        RECT 17.676 231.596 18.036 231.788 ; 
        RECT 23.292 231.596 23.364 231.788 ; 
        RECT 37.908 231.596 37.98 231.788 ; 
        RECT 0.468 235.916 0.54 236.108 ; 
        RECT 15.084 235.916 15.156 236.108 ; 
        RECT 17.676 235.916 18.036 236.108 ; 
        RECT 23.292 235.916 23.364 236.108 ; 
        RECT 37.908 235.916 37.98 236.108 ; 
        RECT 0.468 240.236 0.54 240.428 ; 
        RECT 15.084 240.236 15.156 240.428 ; 
        RECT 17.676 240.236 18.036 240.428 ; 
        RECT 23.292 240.236 23.364 240.428 ; 
        RECT 37.908 240.236 37.98 240.428 ; 
        RECT 0.468 244.556 0.54 244.748 ; 
        RECT 15.084 244.556 15.156 244.748 ; 
        RECT 17.676 244.556 18.036 244.748 ; 
        RECT 23.292 244.556 23.364 244.748 ; 
        RECT 37.908 244.556 37.98 244.748 ; 
        RECT 0.468 248.876 0.54 249.068 ; 
        RECT 15.084 248.876 15.156 249.068 ; 
        RECT 17.676 248.876 18.036 249.068 ; 
        RECT 23.292 248.876 23.364 249.068 ; 
        RECT 37.908 248.876 37.98 249.068 ; 
        RECT 0.468 253.196 0.54 253.388 ; 
        RECT 15.084 253.196 15.156 253.388 ; 
        RECT 17.676 253.196 18.036 253.388 ; 
        RECT 23.292 253.196 23.364 253.388 ; 
        RECT 37.908 253.196 37.98 253.388 ; 
        RECT 0.468 257.516 0.54 257.708 ; 
        RECT 15.084 257.516 15.156 257.708 ; 
        RECT 17.676 257.516 18.036 257.708 ; 
        RECT 23.292 257.516 23.364 257.708 ; 
        RECT 37.908 257.516 37.98 257.708 ; 
        RECT 0.468 261.836 0.54 262.028 ; 
        RECT 15.084 261.836 15.156 262.028 ; 
        RECT 17.676 261.836 18.036 262.028 ; 
        RECT 23.292 261.836 23.364 262.028 ; 
        RECT 37.908 261.836 37.98 262.028 ; 
        RECT 0.468 266.156 0.54 266.348 ; 
        RECT 15.084 266.156 15.156 266.348 ; 
        RECT 17.676 266.156 18.036 266.348 ; 
        RECT 23.292 266.156 23.364 266.348 ; 
        RECT 37.908 266.156 37.98 266.348 ; 
        RECT 0.468 270.476 0.54 270.668 ; 
        RECT 15.084 270.476 15.156 270.668 ; 
        RECT 17.676 270.476 18.036 270.668 ; 
        RECT 23.292 270.476 23.364 270.668 ; 
        RECT 37.908 270.476 37.98 270.668 ; 
        RECT 0.468 274.796 0.54 274.988 ; 
        RECT 15.084 274.796 15.156 274.988 ; 
        RECT 17.676 274.796 18.036 274.988 ; 
        RECT 23.292 274.796 23.364 274.988 ; 
        RECT 37.908 274.796 37.98 274.988 ; 
        RECT 0.468 279.116 0.54 279.308 ; 
        RECT 15.084 279.116 15.156 279.308 ; 
        RECT 17.676 279.116 18.036 279.308 ; 
        RECT 23.292 279.116 23.364 279.308 ; 
        RECT 37.908 279.116 37.98 279.308 ; 
        RECT 0.468 283.436 0.54 283.628 ; 
        RECT 15.084 283.436 15.156 283.628 ; 
        RECT 17.676 283.436 18.036 283.628 ; 
        RECT 23.292 283.436 23.364 283.628 ; 
        RECT 37.908 283.436 37.98 283.628 ; 
        RECT 0.468 287.756 0.54 287.948 ; 
        RECT 15.084 287.756 15.156 287.948 ; 
        RECT 17.676 287.756 18.036 287.948 ; 
        RECT 23.292 287.756 23.364 287.948 ; 
        RECT 37.908 287.756 37.98 287.948 ; 
        RECT 0.468 292.076 0.54 292.268 ; 
        RECT 15.084 292.076 15.156 292.268 ; 
        RECT 17.676 292.076 18.036 292.268 ; 
        RECT 23.292 292.076 23.364 292.268 ; 
        RECT 37.908 292.076 37.98 292.268 ; 
        RECT 0.468 296.396 0.54 296.588 ; 
        RECT 15.084 296.396 15.156 296.588 ; 
        RECT 17.676 296.396 18.036 296.588 ; 
        RECT 23.292 296.396 23.364 296.588 ; 
        RECT 37.908 296.396 37.98 296.588 ; 
        RECT 0.468 300.716 0.54 300.908 ; 
        RECT 15.084 300.716 15.156 300.908 ; 
        RECT 17.676 300.716 18.036 300.908 ; 
        RECT 23.292 300.716 23.364 300.908 ; 
        RECT 37.908 300.716 37.98 300.908 ; 
        RECT 0.468 305.036 0.54 305.228 ; 
        RECT 15.084 305.036 15.156 305.228 ; 
        RECT 17.676 305.036 18.036 305.228 ; 
        RECT 23.292 305.036 23.364 305.228 ; 
        RECT 37.908 305.036 37.98 305.228 ; 
        RECT 0.468 309.356 0.54 309.548 ; 
        RECT 15.084 309.356 15.156 309.548 ; 
        RECT 17.676 309.356 18.036 309.548 ; 
        RECT 23.292 309.356 23.364 309.548 ; 
        RECT 37.908 309.356 37.98 309.548 ; 
        RECT 0.468 313.676 0.54 313.868 ; 
        RECT 15.084 313.676 15.156 313.868 ; 
        RECT 17.676 313.676 18.036 313.868 ; 
        RECT 23.292 313.676 23.364 313.868 ; 
        RECT 37.908 313.676 37.98 313.868 ; 
        RECT 0.468 317.996 0.54 318.188 ; 
        RECT 15.084 317.996 15.156 318.188 ; 
        RECT 17.676 317.996 18.036 318.188 ; 
        RECT 23.292 317.996 23.364 318.188 ; 
        RECT 37.908 317.996 37.98 318.188 ; 
        RECT 0.468 322.316 0.54 322.508 ; 
        RECT 15.084 322.316 15.156 322.508 ; 
        RECT 17.676 322.316 18.036 322.508 ; 
        RECT 23.292 322.316 23.364 322.508 ; 
        RECT 37.908 322.316 37.98 322.508 ; 
        RECT 0.468 326.636 0.54 326.828 ; 
        RECT 15.084 326.636 15.156 326.828 ; 
        RECT 17.676 326.636 18.036 326.828 ; 
        RECT 23.292 326.636 23.364 326.828 ; 
        RECT 37.908 326.636 37.98 326.828 ; 
        RECT 0.468 330.956 0.54 331.148 ; 
        RECT 15.084 330.956 15.156 331.148 ; 
        RECT 17.676 330.956 18.036 331.148 ; 
        RECT 23.292 330.956 23.364 331.148 ; 
        RECT 37.908 330.956 37.98 331.148 ; 
        RECT 0.468 335.276 0.54 335.468 ; 
        RECT 15.084 335.276 15.156 335.468 ; 
        RECT 17.676 335.276 18.036 335.468 ; 
        RECT 23.292 335.276 23.364 335.468 ; 
        RECT 37.908 335.276 37.98 335.468 ; 
        RECT 0.468 339.596 0.54 339.788 ; 
        RECT 15.084 339.596 15.156 339.788 ; 
        RECT 17.676 339.596 18.036 339.788 ; 
        RECT 23.292 339.596 23.364 339.788 ; 
        RECT 37.908 339.596 37.98 339.788 ; 
        RECT 0.468 343.916 0.54 344.108 ; 
        RECT 15.084 343.916 15.156 344.108 ; 
        RECT 17.676 343.916 18.036 344.108 ; 
        RECT 23.292 343.916 23.364 344.108 ; 
        RECT 37.908 343.916 37.98 344.108 ; 
        RECT 0.468 348.236 0.54 348.428 ; 
        RECT 15.084 348.236 15.156 348.428 ; 
        RECT 17.676 348.236 18.036 348.428 ; 
        RECT 23.292 348.236 23.364 348.428 ; 
        RECT 37.908 348.236 37.98 348.428 ; 
        RECT 0.468 352.556 0.54 352.748 ; 
        RECT 15.084 352.556 15.156 352.748 ; 
        RECT 17.676 352.556 18.036 352.748 ; 
        RECT 23.292 352.556 23.364 352.748 ; 
        RECT 37.908 352.556 37.98 352.748 ; 
        RECT 0.468 356.876 0.54 357.068 ; 
        RECT 15.084 356.876 15.156 357.068 ; 
        RECT 17.676 356.876 18.036 357.068 ; 
        RECT 23.292 356.876 23.364 357.068 ; 
        RECT 37.908 356.876 37.98 357.068 ; 
        RECT 0.468 361.196 0.54 361.388 ; 
        RECT 15.084 361.196 15.156 361.388 ; 
        RECT 17.676 361.196 18.036 361.388 ; 
        RECT 23.292 361.196 23.364 361.388 ; 
        RECT 37.908 361.196 37.98 361.388 ; 
        RECT 0.468 365.516 0.54 365.708 ; 
        RECT 15.084 365.516 15.156 365.708 ; 
        RECT 17.676 365.516 18.036 365.708 ; 
        RECT 23.292 365.516 23.364 365.708 ; 
        RECT 37.908 365.516 37.98 365.708 ; 
        RECT 0.468 369.836 0.54 370.028 ; 
        RECT 15.084 369.836 15.156 370.028 ; 
        RECT 17.676 369.836 18.036 370.028 ; 
        RECT 23.292 369.836 23.364 370.028 ; 
        RECT 37.908 369.836 37.98 370.028 ; 
        RECT 0.468 374.156 0.54 374.348 ; 
        RECT 15.084 374.156 15.156 374.348 ; 
        RECT 17.676 374.156 18.036 374.348 ; 
        RECT 23.292 374.156 23.364 374.348 ; 
        RECT 37.908 374.156 37.98 374.348 ; 
        RECT 0.468 378.476 0.54 378.668 ; 
        RECT 15.084 378.476 15.156 378.668 ; 
        RECT 17.676 378.476 18.036 378.668 ; 
        RECT 23.292 378.476 23.364 378.668 ; 
        RECT 37.908 378.476 37.98 378.668 ; 
      LAYER M5 ; 
        RECT 23.036 173.924 23.132 189.3 ; 
      LAYER V4 ; 
        RECT 23.036 189.132 23.132 189.228 ; 
        RECT 23.036 173.996 23.132 174.092 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.304 38.016 4.496 ; 
        RECT 0.404 8.624 38.016 8.816 ; 
        RECT 0.404 12.944 38.016 13.136 ; 
        RECT 0.404 17.264 38.016 17.456 ; 
        RECT 0.404 21.584 38.016 21.776 ; 
        RECT 0.404 25.904 38.016 26.096 ; 
        RECT 0.404 30.224 38.016 30.416 ; 
        RECT 0.404 34.544 38.016 34.736 ; 
        RECT 0.404 38.864 38.016 39.056 ; 
        RECT 0.404 43.184 38.016 43.376 ; 
        RECT 0.404 47.504 38.016 47.696 ; 
        RECT 0.404 51.824 38.016 52.016 ; 
        RECT 0.404 56.144 38.016 56.336 ; 
        RECT 0.404 60.464 38.016 60.656 ; 
        RECT 0.404 64.784 38.016 64.976 ; 
        RECT 0.404 69.104 38.016 69.296 ; 
        RECT 0.404 73.424 38.016 73.616 ; 
        RECT 0.404 77.744 38.016 77.936 ; 
        RECT 0.404 82.064 38.016 82.256 ; 
        RECT 0.404 86.384 38.016 86.576 ; 
        RECT 0.404 90.704 38.016 90.896 ; 
        RECT 0.404 95.024 38.016 95.216 ; 
        RECT 0.404 99.344 38.016 99.536 ; 
        RECT 0.404 103.664 38.016 103.856 ; 
        RECT 0.404 107.984 38.016 108.176 ; 
        RECT 0.404 112.304 38.016 112.496 ; 
        RECT 0.404 116.624 38.016 116.816 ; 
        RECT 0.404 120.944 38.016 121.136 ; 
        RECT 0.404 125.264 38.016 125.456 ; 
        RECT 0.404 129.584 38.016 129.776 ; 
        RECT 0.404 133.904 38.016 134.096 ; 
        RECT 0.404 138.224 38.016 138.416 ; 
        RECT 0.404 142.544 38.016 142.736 ; 
        RECT 0.404 146.864 38.016 147.056 ; 
        RECT 0.404 151.184 38.016 151.376 ; 
        RECT 0.404 155.504 38.016 155.696 ; 
        RECT 0.404 159.824 38.016 160.016 ; 
        RECT 0.404 164.144 38.016 164.336 ; 
        RECT 0.404 168.464 38.016 168.656 ; 
        RECT 0.404 172.784 38.016 172.976 ; 
        RECT 0.432 176.844 38.016 177.708 ; 
        RECT 15.768 189.516 22.68 190.38 ; 
        RECT 15.768 202.188 22.68 203.052 ; 
        RECT 0.404 209.612 38.016 209.804 ; 
        RECT 0.404 213.932 38.016 214.124 ; 
        RECT 0.404 218.252 38.016 218.444 ; 
        RECT 0.404 222.572 38.016 222.764 ; 
        RECT 0.404 226.892 38.016 227.084 ; 
        RECT 0.404 231.212 38.016 231.404 ; 
        RECT 0.404 235.532 38.016 235.724 ; 
        RECT 0.404 239.852 38.016 240.044 ; 
        RECT 0.404 244.172 38.016 244.364 ; 
        RECT 0.404 248.492 38.016 248.684 ; 
        RECT 0.404 252.812 38.016 253.004 ; 
        RECT 0.404 257.132 38.016 257.324 ; 
        RECT 0.404 261.452 38.016 261.644 ; 
        RECT 0.404 265.772 38.016 265.964 ; 
        RECT 0.404 270.092 38.016 270.284 ; 
        RECT 0.404 274.412 38.016 274.604 ; 
        RECT 0.404 278.732 38.016 278.924 ; 
        RECT 0.404 283.052 38.016 283.244 ; 
        RECT 0.404 287.372 38.016 287.564 ; 
        RECT 0.404 291.692 38.016 291.884 ; 
        RECT 0.404 296.012 38.016 296.204 ; 
        RECT 0.404 300.332 38.016 300.524 ; 
        RECT 0.404 304.652 38.016 304.844 ; 
        RECT 0.404 308.972 38.016 309.164 ; 
        RECT 0.404 313.292 38.016 313.484 ; 
        RECT 0.404 317.612 38.016 317.804 ; 
        RECT 0.404 321.932 38.016 322.124 ; 
        RECT 0.404 326.252 38.016 326.444 ; 
        RECT 0.404 330.572 38.016 330.764 ; 
        RECT 0.404 334.892 38.016 335.084 ; 
        RECT 0.404 339.212 38.016 339.404 ; 
        RECT 0.404 343.532 38.016 343.724 ; 
        RECT 0.404 347.852 38.016 348.044 ; 
        RECT 0.404 352.172 38.016 352.364 ; 
        RECT 0.404 356.492 38.016 356.684 ; 
        RECT 0.404 360.812 38.016 361.004 ; 
        RECT 0.404 365.132 38.016 365.324 ; 
        RECT 0.404 369.452 38.016 369.644 ; 
        RECT 0.404 373.772 38.016 373.964 ; 
        RECT 0.404 378.092 38.016 378.284 ; 
      LAYER M3 ; 
        RECT 37.764 0.866 37.836 5.506 ; 
        RECT 23.508 0.866 23.58 5.506 ; 
        RECT 20.448 1.012 20.592 5.468 ; 
        RECT 19.836 1.012 19.944 5.468 ; 
        RECT 14.868 0.866 14.94 5.506 ; 
        RECT 0.612 0.866 0.684 5.506 ; 
        RECT 37.764 5.186 37.836 9.826 ; 
        RECT 23.508 5.186 23.58 9.826 ; 
        RECT 20.448 5.332 20.592 9.788 ; 
        RECT 19.836 5.332 19.944 9.788 ; 
        RECT 14.868 5.186 14.94 9.826 ; 
        RECT 0.612 5.186 0.684 9.826 ; 
        RECT 37.764 9.506 37.836 14.146 ; 
        RECT 23.508 9.506 23.58 14.146 ; 
        RECT 20.448 9.652 20.592 14.108 ; 
        RECT 19.836 9.652 19.944 14.108 ; 
        RECT 14.868 9.506 14.94 14.146 ; 
        RECT 0.612 9.506 0.684 14.146 ; 
        RECT 37.764 13.826 37.836 18.466 ; 
        RECT 23.508 13.826 23.58 18.466 ; 
        RECT 20.448 13.972 20.592 18.428 ; 
        RECT 19.836 13.972 19.944 18.428 ; 
        RECT 14.868 13.826 14.94 18.466 ; 
        RECT 0.612 13.826 0.684 18.466 ; 
        RECT 37.764 18.146 37.836 22.786 ; 
        RECT 23.508 18.146 23.58 22.786 ; 
        RECT 20.448 18.292 20.592 22.748 ; 
        RECT 19.836 18.292 19.944 22.748 ; 
        RECT 14.868 18.146 14.94 22.786 ; 
        RECT 0.612 18.146 0.684 22.786 ; 
        RECT 37.764 22.466 37.836 27.106 ; 
        RECT 23.508 22.466 23.58 27.106 ; 
        RECT 20.448 22.612 20.592 27.068 ; 
        RECT 19.836 22.612 19.944 27.068 ; 
        RECT 14.868 22.466 14.94 27.106 ; 
        RECT 0.612 22.466 0.684 27.106 ; 
        RECT 37.764 26.786 37.836 31.426 ; 
        RECT 23.508 26.786 23.58 31.426 ; 
        RECT 20.448 26.932 20.592 31.388 ; 
        RECT 19.836 26.932 19.944 31.388 ; 
        RECT 14.868 26.786 14.94 31.426 ; 
        RECT 0.612 26.786 0.684 31.426 ; 
        RECT 37.764 31.106 37.836 35.746 ; 
        RECT 23.508 31.106 23.58 35.746 ; 
        RECT 20.448 31.252 20.592 35.708 ; 
        RECT 19.836 31.252 19.944 35.708 ; 
        RECT 14.868 31.106 14.94 35.746 ; 
        RECT 0.612 31.106 0.684 35.746 ; 
        RECT 37.764 35.426 37.836 40.066 ; 
        RECT 23.508 35.426 23.58 40.066 ; 
        RECT 20.448 35.572 20.592 40.028 ; 
        RECT 19.836 35.572 19.944 40.028 ; 
        RECT 14.868 35.426 14.94 40.066 ; 
        RECT 0.612 35.426 0.684 40.066 ; 
        RECT 37.764 39.746 37.836 44.386 ; 
        RECT 23.508 39.746 23.58 44.386 ; 
        RECT 20.448 39.892 20.592 44.348 ; 
        RECT 19.836 39.892 19.944 44.348 ; 
        RECT 14.868 39.746 14.94 44.386 ; 
        RECT 0.612 39.746 0.684 44.386 ; 
        RECT 37.764 44.066 37.836 48.706 ; 
        RECT 23.508 44.066 23.58 48.706 ; 
        RECT 20.448 44.212 20.592 48.668 ; 
        RECT 19.836 44.212 19.944 48.668 ; 
        RECT 14.868 44.066 14.94 48.706 ; 
        RECT 0.612 44.066 0.684 48.706 ; 
        RECT 37.764 48.386 37.836 53.026 ; 
        RECT 23.508 48.386 23.58 53.026 ; 
        RECT 20.448 48.532 20.592 52.988 ; 
        RECT 19.836 48.532 19.944 52.988 ; 
        RECT 14.868 48.386 14.94 53.026 ; 
        RECT 0.612 48.386 0.684 53.026 ; 
        RECT 37.764 52.706 37.836 57.346 ; 
        RECT 23.508 52.706 23.58 57.346 ; 
        RECT 20.448 52.852 20.592 57.308 ; 
        RECT 19.836 52.852 19.944 57.308 ; 
        RECT 14.868 52.706 14.94 57.346 ; 
        RECT 0.612 52.706 0.684 57.346 ; 
        RECT 37.764 57.026 37.836 61.666 ; 
        RECT 23.508 57.026 23.58 61.666 ; 
        RECT 20.448 57.172 20.592 61.628 ; 
        RECT 19.836 57.172 19.944 61.628 ; 
        RECT 14.868 57.026 14.94 61.666 ; 
        RECT 0.612 57.026 0.684 61.666 ; 
        RECT 37.764 61.346 37.836 65.986 ; 
        RECT 23.508 61.346 23.58 65.986 ; 
        RECT 20.448 61.492 20.592 65.948 ; 
        RECT 19.836 61.492 19.944 65.948 ; 
        RECT 14.868 61.346 14.94 65.986 ; 
        RECT 0.612 61.346 0.684 65.986 ; 
        RECT 37.764 65.666 37.836 70.306 ; 
        RECT 23.508 65.666 23.58 70.306 ; 
        RECT 20.448 65.812 20.592 70.268 ; 
        RECT 19.836 65.812 19.944 70.268 ; 
        RECT 14.868 65.666 14.94 70.306 ; 
        RECT 0.612 65.666 0.684 70.306 ; 
        RECT 37.764 69.986 37.836 74.626 ; 
        RECT 23.508 69.986 23.58 74.626 ; 
        RECT 20.448 70.132 20.592 74.588 ; 
        RECT 19.836 70.132 19.944 74.588 ; 
        RECT 14.868 69.986 14.94 74.626 ; 
        RECT 0.612 69.986 0.684 74.626 ; 
        RECT 37.764 74.306 37.836 78.946 ; 
        RECT 23.508 74.306 23.58 78.946 ; 
        RECT 20.448 74.452 20.592 78.908 ; 
        RECT 19.836 74.452 19.944 78.908 ; 
        RECT 14.868 74.306 14.94 78.946 ; 
        RECT 0.612 74.306 0.684 78.946 ; 
        RECT 37.764 78.626 37.836 83.266 ; 
        RECT 23.508 78.626 23.58 83.266 ; 
        RECT 20.448 78.772 20.592 83.228 ; 
        RECT 19.836 78.772 19.944 83.228 ; 
        RECT 14.868 78.626 14.94 83.266 ; 
        RECT 0.612 78.626 0.684 83.266 ; 
        RECT 37.764 82.946 37.836 87.586 ; 
        RECT 23.508 82.946 23.58 87.586 ; 
        RECT 20.448 83.092 20.592 87.548 ; 
        RECT 19.836 83.092 19.944 87.548 ; 
        RECT 14.868 82.946 14.94 87.586 ; 
        RECT 0.612 82.946 0.684 87.586 ; 
        RECT 37.764 87.266 37.836 91.906 ; 
        RECT 23.508 87.266 23.58 91.906 ; 
        RECT 20.448 87.412 20.592 91.868 ; 
        RECT 19.836 87.412 19.944 91.868 ; 
        RECT 14.868 87.266 14.94 91.906 ; 
        RECT 0.612 87.266 0.684 91.906 ; 
        RECT 37.764 91.586 37.836 96.226 ; 
        RECT 23.508 91.586 23.58 96.226 ; 
        RECT 20.448 91.732 20.592 96.188 ; 
        RECT 19.836 91.732 19.944 96.188 ; 
        RECT 14.868 91.586 14.94 96.226 ; 
        RECT 0.612 91.586 0.684 96.226 ; 
        RECT 37.764 95.906 37.836 100.546 ; 
        RECT 23.508 95.906 23.58 100.546 ; 
        RECT 20.448 96.052 20.592 100.508 ; 
        RECT 19.836 96.052 19.944 100.508 ; 
        RECT 14.868 95.906 14.94 100.546 ; 
        RECT 0.612 95.906 0.684 100.546 ; 
        RECT 37.764 100.226 37.836 104.866 ; 
        RECT 23.508 100.226 23.58 104.866 ; 
        RECT 20.448 100.372 20.592 104.828 ; 
        RECT 19.836 100.372 19.944 104.828 ; 
        RECT 14.868 100.226 14.94 104.866 ; 
        RECT 0.612 100.226 0.684 104.866 ; 
        RECT 37.764 104.546 37.836 109.186 ; 
        RECT 23.508 104.546 23.58 109.186 ; 
        RECT 20.448 104.692 20.592 109.148 ; 
        RECT 19.836 104.692 19.944 109.148 ; 
        RECT 14.868 104.546 14.94 109.186 ; 
        RECT 0.612 104.546 0.684 109.186 ; 
        RECT 37.764 108.866 37.836 113.506 ; 
        RECT 23.508 108.866 23.58 113.506 ; 
        RECT 20.448 109.012 20.592 113.468 ; 
        RECT 19.836 109.012 19.944 113.468 ; 
        RECT 14.868 108.866 14.94 113.506 ; 
        RECT 0.612 108.866 0.684 113.506 ; 
        RECT 37.764 113.186 37.836 117.826 ; 
        RECT 23.508 113.186 23.58 117.826 ; 
        RECT 20.448 113.332 20.592 117.788 ; 
        RECT 19.836 113.332 19.944 117.788 ; 
        RECT 14.868 113.186 14.94 117.826 ; 
        RECT 0.612 113.186 0.684 117.826 ; 
        RECT 37.764 117.506 37.836 122.146 ; 
        RECT 23.508 117.506 23.58 122.146 ; 
        RECT 20.448 117.652 20.592 122.108 ; 
        RECT 19.836 117.652 19.944 122.108 ; 
        RECT 14.868 117.506 14.94 122.146 ; 
        RECT 0.612 117.506 0.684 122.146 ; 
        RECT 37.764 121.826 37.836 126.466 ; 
        RECT 23.508 121.826 23.58 126.466 ; 
        RECT 20.448 121.972 20.592 126.428 ; 
        RECT 19.836 121.972 19.944 126.428 ; 
        RECT 14.868 121.826 14.94 126.466 ; 
        RECT 0.612 121.826 0.684 126.466 ; 
        RECT 37.764 126.146 37.836 130.786 ; 
        RECT 23.508 126.146 23.58 130.786 ; 
        RECT 20.448 126.292 20.592 130.748 ; 
        RECT 19.836 126.292 19.944 130.748 ; 
        RECT 14.868 126.146 14.94 130.786 ; 
        RECT 0.612 126.146 0.684 130.786 ; 
        RECT 37.764 130.466 37.836 135.106 ; 
        RECT 23.508 130.466 23.58 135.106 ; 
        RECT 20.448 130.612 20.592 135.068 ; 
        RECT 19.836 130.612 19.944 135.068 ; 
        RECT 14.868 130.466 14.94 135.106 ; 
        RECT 0.612 130.466 0.684 135.106 ; 
        RECT 37.764 134.786 37.836 139.426 ; 
        RECT 23.508 134.786 23.58 139.426 ; 
        RECT 20.448 134.932 20.592 139.388 ; 
        RECT 19.836 134.932 19.944 139.388 ; 
        RECT 14.868 134.786 14.94 139.426 ; 
        RECT 0.612 134.786 0.684 139.426 ; 
        RECT 37.764 139.106 37.836 143.746 ; 
        RECT 23.508 139.106 23.58 143.746 ; 
        RECT 20.448 139.252 20.592 143.708 ; 
        RECT 19.836 139.252 19.944 143.708 ; 
        RECT 14.868 139.106 14.94 143.746 ; 
        RECT 0.612 139.106 0.684 143.746 ; 
        RECT 37.764 143.426 37.836 148.066 ; 
        RECT 23.508 143.426 23.58 148.066 ; 
        RECT 20.448 143.572 20.592 148.028 ; 
        RECT 19.836 143.572 19.944 148.028 ; 
        RECT 14.868 143.426 14.94 148.066 ; 
        RECT 0.612 143.426 0.684 148.066 ; 
        RECT 37.764 147.746 37.836 152.386 ; 
        RECT 23.508 147.746 23.58 152.386 ; 
        RECT 20.448 147.892 20.592 152.348 ; 
        RECT 19.836 147.892 19.944 152.348 ; 
        RECT 14.868 147.746 14.94 152.386 ; 
        RECT 0.612 147.746 0.684 152.386 ; 
        RECT 37.764 152.066 37.836 156.706 ; 
        RECT 23.508 152.066 23.58 156.706 ; 
        RECT 20.448 152.212 20.592 156.668 ; 
        RECT 19.836 152.212 19.944 156.668 ; 
        RECT 14.868 152.066 14.94 156.706 ; 
        RECT 0.612 152.066 0.684 156.706 ; 
        RECT 37.764 156.386 37.836 161.026 ; 
        RECT 23.508 156.386 23.58 161.026 ; 
        RECT 20.448 156.532 20.592 160.988 ; 
        RECT 19.836 156.532 19.944 160.988 ; 
        RECT 14.868 156.386 14.94 161.026 ; 
        RECT 0.612 156.386 0.684 161.026 ; 
        RECT 37.764 160.706 37.836 165.346 ; 
        RECT 23.508 160.706 23.58 165.346 ; 
        RECT 20.448 160.852 20.592 165.308 ; 
        RECT 19.836 160.852 19.944 165.308 ; 
        RECT 14.868 160.706 14.94 165.346 ; 
        RECT 0.612 160.706 0.684 165.346 ; 
        RECT 37.764 165.026 37.836 169.666 ; 
        RECT 23.508 165.026 23.58 169.666 ; 
        RECT 20.448 165.172 20.592 169.628 ; 
        RECT 19.836 165.172 19.944 169.628 ; 
        RECT 14.868 165.026 14.94 169.666 ; 
        RECT 0.612 165.026 0.684 169.666 ; 
        RECT 37.764 169.346 37.836 173.986 ; 
        RECT 23.508 169.346 23.58 173.986 ; 
        RECT 20.448 169.492 20.592 173.948 ; 
        RECT 19.836 169.492 19.944 173.948 ; 
        RECT 14.868 169.346 14.94 173.986 ; 
        RECT 0.612 169.346 0.684 173.986 ; 
        RECT 37.764 173.666 37.836 206.494 ; 
        RECT 23.508 173.666 23.58 206.494 ; 
        RECT 19.692 174.56 20.628 205.292 ; 
        RECT 20.448 173.84 20.592 206.388 ; 
        RECT 19.836 173.84 19.944 206.376 ; 
        RECT 14.868 173.666 14.94 206.494 ; 
        RECT 0.612 173.666 0.684 206.494 ; 
        RECT 37.764 206.174 37.836 210.814 ; 
        RECT 23.508 206.174 23.58 210.814 ; 
        RECT 20.448 206.32 20.592 210.776 ; 
        RECT 19.836 206.32 19.944 210.776 ; 
        RECT 14.868 206.174 14.94 210.814 ; 
        RECT 0.612 206.174 0.684 210.814 ; 
        RECT 37.764 210.494 37.836 215.134 ; 
        RECT 23.508 210.494 23.58 215.134 ; 
        RECT 20.448 210.64 20.592 215.096 ; 
        RECT 19.836 210.64 19.944 215.096 ; 
        RECT 14.868 210.494 14.94 215.134 ; 
        RECT 0.612 210.494 0.684 215.134 ; 
        RECT 37.764 214.814 37.836 219.454 ; 
        RECT 23.508 214.814 23.58 219.454 ; 
        RECT 20.448 214.96 20.592 219.416 ; 
        RECT 19.836 214.96 19.944 219.416 ; 
        RECT 14.868 214.814 14.94 219.454 ; 
        RECT 0.612 214.814 0.684 219.454 ; 
        RECT 37.764 219.134 37.836 223.774 ; 
        RECT 23.508 219.134 23.58 223.774 ; 
        RECT 20.448 219.28 20.592 223.736 ; 
        RECT 19.836 219.28 19.944 223.736 ; 
        RECT 14.868 219.134 14.94 223.774 ; 
        RECT 0.612 219.134 0.684 223.774 ; 
        RECT 37.764 223.454 37.836 228.094 ; 
        RECT 23.508 223.454 23.58 228.094 ; 
        RECT 20.448 223.6 20.592 228.056 ; 
        RECT 19.836 223.6 19.944 228.056 ; 
        RECT 14.868 223.454 14.94 228.094 ; 
        RECT 0.612 223.454 0.684 228.094 ; 
        RECT 37.764 227.774 37.836 232.414 ; 
        RECT 23.508 227.774 23.58 232.414 ; 
        RECT 20.448 227.92 20.592 232.376 ; 
        RECT 19.836 227.92 19.944 232.376 ; 
        RECT 14.868 227.774 14.94 232.414 ; 
        RECT 0.612 227.774 0.684 232.414 ; 
        RECT 37.764 232.094 37.836 236.734 ; 
        RECT 23.508 232.094 23.58 236.734 ; 
        RECT 20.448 232.24 20.592 236.696 ; 
        RECT 19.836 232.24 19.944 236.696 ; 
        RECT 14.868 232.094 14.94 236.734 ; 
        RECT 0.612 232.094 0.684 236.734 ; 
        RECT 37.764 236.414 37.836 241.054 ; 
        RECT 23.508 236.414 23.58 241.054 ; 
        RECT 20.448 236.56 20.592 241.016 ; 
        RECT 19.836 236.56 19.944 241.016 ; 
        RECT 14.868 236.414 14.94 241.054 ; 
        RECT 0.612 236.414 0.684 241.054 ; 
        RECT 37.764 240.734 37.836 245.374 ; 
        RECT 23.508 240.734 23.58 245.374 ; 
        RECT 20.448 240.88 20.592 245.336 ; 
        RECT 19.836 240.88 19.944 245.336 ; 
        RECT 14.868 240.734 14.94 245.374 ; 
        RECT 0.612 240.734 0.684 245.374 ; 
        RECT 37.764 245.054 37.836 249.694 ; 
        RECT 23.508 245.054 23.58 249.694 ; 
        RECT 20.448 245.2 20.592 249.656 ; 
        RECT 19.836 245.2 19.944 249.656 ; 
        RECT 14.868 245.054 14.94 249.694 ; 
        RECT 0.612 245.054 0.684 249.694 ; 
        RECT 37.764 249.374 37.836 254.014 ; 
        RECT 23.508 249.374 23.58 254.014 ; 
        RECT 20.448 249.52 20.592 253.976 ; 
        RECT 19.836 249.52 19.944 253.976 ; 
        RECT 14.868 249.374 14.94 254.014 ; 
        RECT 0.612 249.374 0.684 254.014 ; 
        RECT 37.764 253.694 37.836 258.334 ; 
        RECT 23.508 253.694 23.58 258.334 ; 
        RECT 20.448 253.84 20.592 258.296 ; 
        RECT 19.836 253.84 19.944 258.296 ; 
        RECT 14.868 253.694 14.94 258.334 ; 
        RECT 0.612 253.694 0.684 258.334 ; 
        RECT 37.764 258.014 37.836 262.654 ; 
        RECT 23.508 258.014 23.58 262.654 ; 
        RECT 20.448 258.16 20.592 262.616 ; 
        RECT 19.836 258.16 19.944 262.616 ; 
        RECT 14.868 258.014 14.94 262.654 ; 
        RECT 0.612 258.014 0.684 262.654 ; 
        RECT 37.764 262.334 37.836 266.974 ; 
        RECT 23.508 262.334 23.58 266.974 ; 
        RECT 20.448 262.48 20.592 266.936 ; 
        RECT 19.836 262.48 19.944 266.936 ; 
        RECT 14.868 262.334 14.94 266.974 ; 
        RECT 0.612 262.334 0.684 266.974 ; 
        RECT 37.764 266.654 37.836 271.294 ; 
        RECT 23.508 266.654 23.58 271.294 ; 
        RECT 20.448 266.8 20.592 271.256 ; 
        RECT 19.836 266.8 19.944 271.256 ; 
        RECT 14.868 266.654 14.94 271.294 ; 
        RECT 0.612 266.654 0.684 271.294 ; 
        RECT 37.764 270.974 37.836 275.614 ; 
        RECT 23.508 270.974 23.58 275.614 ; 
        RECT 20.448 271.12 20.592 275.576 ; 
        RECT 19.836 271.12 19.944 275.576 ; 
        RECT 14.868 270.974 14.94 275.614 ; 
        RECT 0.612 270.974 0.684 275.614 ; 
        RECT 37.764 275.294 37.836 279.934 ; 
        RECT 23.508 275.294 23.58 279.934 ; 
        RECT 20.448 275.44 20.592 279.896 ; 
        RECT 19.836 275.44 19.944 279.896 ; 
        RECT 14.868 275.294 14.94 279.934 ; 
        RECT 0.612 275.294 0.684 279.934 ; 
        RECT 37.764 279.614 37.836 284.254 ; 
        RECT 23.508 279.614 23.58 284.254 ; 
        RECT 20.448 279.76 20.592 284.216 ; 
        RECT 19.836 279.76 19.944 284.216 ; 
        RECT 14.868 279.614 14.94 284.254 ; 
        RECT 0.612 279.614 0.684 284.254 ; 
        RECT 37.764 283.934 37.836 288.574 ; 
        RECT 23.508 283.934 23.58 288.574 ; 
        RECT 20.448 284.08 20.592 288.536 ; 
        RECT 19.836 284.08 19.944 288.536 ; 
        RECT 14.868 283.934 14.94 288.574 ; 
        RECT 0.612 283.934 0.684 288.574 ; 
        RECT 37.764 288.254 37.836 292.894 ; 
        RECT 23.508 288.254 23.58 292.894 ; 
        RECT 20.448 288.4 20.592 292.856 ; 
        RECT 19.836 288.4 19.944 292.856 ; 
        RECT 14.868 288.254 14.94 292.894 ; 
        RECT 0.612 288.254 0.684 292.894 ; 
        RECT 37.764 292.574 37.836 297.214 ; 
        RECT 23.508 292.574 23.58 297.214 ; 
        RECT 20.448 292.72 20.592 297.176 ; 
        RECT 19.836 292.72 19.944 297.176 ; 
        RECT 14.868 292.574 14.94 297.214 ; 
        RECT 0.612 292.574 0.684 297.214 ; 
        RECT 37.764 296.894 37.836 301.534 ; 
        RECT 23.508 296.894 23.58 301.534 ; 
        RECT 20.448 297.04 20.592 301.496 ; 
        RECT 19.836 297.04 19.944 301.496 ; 
        RECT 14.868 296.894 14.94 301.534 ; 
        RECT 0.612 296.894 0.684 301.534 ; 
        RECT 37.764 301.214 37.836 305.854 ; 
        RECT 23.508 301.214 23.58 305.854 ; 
        RECT 20.448 301.36 20.592 305.816 ; 
        RECT 19.836 301.36 19.944 305.816 ; 
        RECT 14.868 301.214 14.94 305.854 ; 
        RECT 0.612 301.214 0.684 305.854 ; 
        RECT 37.764 305.534 37.836 310.174 ; 
        RECT 23.508 305.534 23.58 310.174 ; 
        RECT 20.448 305.68 20.592 310.136 ; 
        RECT 19.836 305.68 19.944 310.136 ; 
        RECT 14.868 305.534 14.94 310.174 ; 
        RECT 0.612 305.534 0.684 310.174 ; 
        RECT 37.764 309.854 37.836 314.494 ; 
        RECT 23.508 309.854 23.58 314.494 ; 
        RECT 20.448 310 20.592 314.456 ; 
        RECT 19.836 310 19.944 314.456 ; 
        RECT 14.868 309.854 14.94 314.494 ; 
        RECT 0.612 309.854 0.684 314.494 ; 
        RECT 37.764 314.174 37.836 318.814 ; 
        RECT 23.508 314.174 23.58 318.814 ; 
        RECT 20.448 314.32 20.592 318.776 ; 
        RECT 19.836 314.32 19.944 318.776 ; 
        RECT 14.868 314.174 14.94 318.814 ; 
        RECT 0.612 314.174 0.684 318.814 ; 
        RECT 37.764 318.494 37.836 323.134 ; 
        RECT 23.508 318.494 23.58 323.134 ; 
        RECT 20.448 318.64 20.592 323.096 ; 
        RECT 19.836 318.64 19.944 323.096 ; 
        RECT 14.868 318.494 14.94 323.134 ; 
        RECT 0.612 318.494 0.684 323.134 ; 
        RECT 37.764 322.814 37.836 327.454 ; 
        RECT 23.508 322.814 23.58 327.454 ; 
        RECT 20.448 322.96 20.592 327.416 ; 
        RECT 19.836 322.96 19.944 327.416 ; 
        RECT 14.868 322.814 14.94 327.454 ; 
        RECT 0.612 322.814 0.684 327.454 ; 
        RECT 37.764 327.134 37.836 331.774 ; 
        RECT 23.508 327.134 23.58 331.774 ; 
        RECT 20.448 327.28 20.592 331.736 ; 
        RECT 19.836 327.28 19.944 331.736 ; 
        RECT 14.868 327.134 14.94 331.774 ; 
        RECT 0.612 327.134 0.684 331.774 ; 
        RECT 37.764 331.454 37.836 336.094 ; 
        RECT 23.508 331.454 23.58 336.094 ; 
        RECT 20.448 331.6 20.592 336.056 ; 
        RECT 19.836 331.6 19.944 336.056 ; 
        RECT 14.868 331.454 14.94 336.094 ; 
        RECT 0.612 331.454 0.684 336.094 ; 
        RECT 37.764 335.774 37.836 340.414 ; 
        RECT 23.508 335.774 23.58 340.414 ; 
        RECT 20.448 335.92 20.592 340.376 ; 
        RECT 19.836 335.92 19.944 340.376 ; 
        RECT 14.868 335.774 14.94 340.414 ; 
        RECT 0.612 335.774 0.684 340.414 ; 
        RECT 37.764 340.094 37.836 344.734 ; 
        RECT 23.508 340.094 23.58 344.734 ; 
        RECT 20.448 340.24 20.592 344.696 ; 
        RECT 19.836 340.24 19.944 344.696 ; 
        RECT 14.868 340.094 14.94 344.734 ; 
        RECT 0.612 340.094 0.684 344.734 ; 
        RECT 37.764 344.414 37.836 349.054 ; 
        RECT 23.508 344.414 23.58 349.054 ; 
        RECT 20.448 344.56 20.592 349.016 ; 
        RECT 19.836 344.56 19.944 349.016 ; 
        RECT 14.868 344.414 14.94 349.054 ; 
        RECT 0.612 344.414 0.684 349.054 ; 
        RECT 37.764 348.734 37.836 353.374 ; 
        RECT 23.508 348.734 23.58 353.374 ; 
        RECT 20.448 348.88 20.592 353.336 ; 
        RECT 19.836 348.88 19.944 353.336 ; 
        RECT 14.868 348.734 14.94 353.374 ; 
        RECT 0.612 348.734 0.684 353.374 ; 
        RECT 37.764 353.054 37.836 357.694 ; 
        RECT 23.508 353.054 23.58 357.694 ; 
        RECT 20.448 353.2 20.592 357.656 ; 
        RECT 19.836 353.2 19.944 357.656 ; 
        RECT 14.868 353.054 14.94 357.694 ; 
        RECT 0.612 353.054 0.684 357.694 ; 
        RECT 37.764 357.374 37.836 362.014 ; 
        RECT 23.508 357.374 23.58 362.014 ; 
        RECT 20.448 357.52 20.592 361.976 ; 
        RECT 19.836 357.52 19.944 361.976 ; 
        RECT 14.868 357.374 14.94 362.014 ; 
        RECT 0.612 357.374 0.684 362.014 ; 
        RECT 37.764 361.694 37.836 366.334 ; 
        RECT 23.508 361.694 23.58 366.334 ; 
        RECT 20.448 361.84 20.592 366.296 ; 
        RECT 19.836 361.84 19.944 366.296 ; 
        RECT 14.868 361.694 14.94 366.334 ; 
        RECT 0.612 361.694 0.684 366.334 ; 
        RECT 37.764 366.014 37.836 370.654 ; 
        RECT 23.508 366.014 23.58 370.654 ; 
        RECT 20.448 366.16 20.592 370.616 ; 
        RECT 19.836 366.16 19.944 370.616 ; 
        RECT 14.868 366.014 14.94 370.654 ; 
        RECT 0.612 366.014 0.684 370.654 ; 
        RECT 37.764 370.334 37.836 374.974 ; 
        RECT 23.508 370.334 23.58 374.974 ; 
        RECT 20.448 370.48 20.592 374.936 ; 
        RECT 19.836 370.48 19.944 374.936 ; 
        RECT 14.868 370.334 14.94 374.974 ; 
        RECT 0.612 370.334 0.684 374.974 ; 
        RECT 37.764 374.654 37.836 379.294 ; 
        RECT 23.508 374.654 23.58 379.294 ; 
        RECT 20.448 374.8 20.592 379.256 ; 
        RECT 19.836 374.8 19.944 379.256 ; 
        RECT 14.868 374.654 14.94 379.294 ; 
        RECT 0.612 374.654 0.684 379.294 ; 
      LAYER V3 ; 
        RECT 0.612 4.304 0.684 4.496 ; 
        RECT 14.868 4.304 14.94 4.496 ; 
        RECT 19.836 4.304 19.944 4.496 ; 
        RECT 20.448 4.304 20.592 4.496 ; 
        RECT 23.508 4.304 23.58 4.496 ; 
        RECT 37.764 4.304 37.836 4.496 ; 
        RECT 0.612 8.624 0.684 8.816 ; 
        RECT 14.868 8.624 14.94 8.816 ; 
        RECT 19.836 8.624 19.944 8.816 ; 
        RECT 20.448 8.624 20.592 8.816 ; 
        RECT 23.508 8.624 23.58 8.816 ; 
        RECT 37.764 8.624 37.836 8.816 ; 
        RECT 0.612 12.944 0.684 13.136 ; 
        RECT 14.868 12.944 14.94 13.136 ; 
        RECT 19.836 12.944 19.944 13.136 ; 
        RECT 20.448 12.944 20.592 13.136 ; 
        RECT 23.508 12.944 23.58 13.136 ; 
        RECT 37.764 12.944 37.836 13.136 ; 
        RECT 0.612 17.264 0.684 17.456 ; 
        RECT 14.868 17.264 14.94 17.456 ; 
        RECT 19.836 17.264 19.944 17.456 ; 
        RECT 20.448 17.264 20.592 17.456 ; 
        RECT 23.508 17.264 23.58 17.456 ; 
        RECT 37.764 17.264 37.836 17.456 ; 
        RECT 0.612 21.584 0.684 21.776 ; 
        RECT 14.868 21.584 14.94 21.776 ; 
        RECT 19.836 21.584 19.944 21.776 ; 
        RECT 20.448 21.584 20.592 21.776 ; 
        RECT 23.508 21.584 23.58 21.776 ; 
        RECT 37.764 21.584 37.836 21.776 ; 
        RECT 0.612 25.904 0.684 26.096 ; 
        RECT 14.868 25.904 14.94 26.096 ; 
        RECT 19.836 25.904 19.944 26.096 ; 
        RECT 20.448 25.904 20.592 26.096 ; 
        RECT 23.508 25.904 23.58 26.096 ; 
        RECT 37.764 25.904 37.836 26.096 ; 
        RECT 0.612 30.224 0.684 30.416 ; 
        RECT 14.868 30.224 14.94 30.416 ; 
        RECT 19.836 30.224 19.944 30.416 ; 
        RECT 20.448 30.224 20.592 30.416 ; 
        RECT 23.508 30.224 23.58 30.416 ; 
        RECT 37.764 30.224 37.836 30.416 ; 
        RECT 0.612 34.544 0.684 34.736 ; 
        RECT 14.868 34.544 14.94 34.736 ; 
        RECT 19.836 34.544 19.944 34.736 ; 
        RECT 20.448 34.544 20.592 34.736 ; 
        RECT 23.508 34.544 23.58 34.736 ; 
        RECT 37.764 34.544 37.836 34.736 ; 
        RECT 0.612 38.864 0.684 39.056 ; 
        RECT 14.868 38.864 14.94 39.056 ; 
        RECT 19.836 38.864 19.944 39.056 ; 
        RECT 20.448 38.864 20.592 39.056 ; 
        RECT 23.508 38.864 23.58 39.056 ; 
        RECT 37.764 38.864 37.836 39.056 ; 
        RECT 0.612 43.184 0.684 43.376 ; 
        RECT 14.868 43.184 14.94 43.376 ; 
        RECT 19.836 43.184 19.944 43.376 ; 
        RECT 20.448 43.184 20.592 43.376 ; 
        RECT 23.508 43.184 23.58 43.376 ; 
        RECT 37.764 43.184 37.836 43.376 ; 
        RECT 0.612 47.504 0.684 47.696 ; 
        RECT 14.868 47.504 14.94 47.696 ; 
        RECT 19.836 47.504 19.944 47.696 ; 
        RECT 20.448 47.504 20.592 47.696 ; 
        RECT 23.508 47.504 23.58 47.696 ; 
        RECT 37.764 47.504 37.836 47.696 ; 
        RECT 0.612 51.824 0.684 52.016 ; 
        RECT 14.868 51.824 14.94 52.016 ; 
        RECT 19.836 51.824 19.944 52.016 ; 
        RECT 20.448 51.824 20.592 52.016 ; 
        RECT 23.508 51.824 23.58 52.016 ; 
        RECT 37.764 51.824 37.836 52.016 ; 
        RECT 0.612 56.144 0.684 56.336 ; 
        RECT 14.868 56.144 14.94 56.336 ; 
        RECT 19.836 56.144 19.944 56.336 ; 
        RECT 20.448 56.144 20.592 56.336 ; 
        RECT 23.508 56.144 23.58 56.336 ; 
        RECT 37.764 56.144 37.836 56.336 ; 
        RECT 0.612 60.464 0.684 60.656 ; 
        RECT 14.868 60.464 14.94 60.656 ; 
        RECT 19.836 60.464 19.944 60.656 ; 
        RECT 20.448 60.464 20.592 60.656 ; 
        RECT 23.508 60.464 23.58 60.656 ; 
        RECT 37.764 60.464 37.836 60.656 ; 
        RECT 0.612 64.784 0.684 64.976 ; 
        RECT 14.868 64.784 14.94 64.976 ; 
        RECT 19.836 64.784 19.944 64.976 ; 
        RECT 20.448 64.784 20.592 64.976 ; 
        RECT 23.508 64.784 23.58 64.976 ; 
        RECT 37.764 64.784 37.836 64.976 ; 
        RECT 0.612 69.104 0.684 69.296 ; 
        RECT 14.868 69.104 14.94 69.296 ; 
        RECT 19.836 69.104 19.944 69.296 ; 
        RECT 20.448 69.104 20.592 69.296 ; 
        RECT 23.508 69.104 23.58 69.296 ; 
        RECT 37.764 69.104 37.836 69.296 ; 
        RECT 0.612 73.424 0.684 73.616 ; 
        RECT 14.868 73.424 14.94 73.616 ; 
        RECT 19.836 73.424 19.944 73.616 ; 
        RECT 20.448 73.424 20.592 73.616 ; 
        RECT 23.508 73.424 23.58 73.616 ; 
        RECT 37.764 73.424 37.836 73.616 ; 
        RECT 0.612 77.744 0.684 77.936 ; 
        RECT 14.868 77.744 14.94 77.936 ; 
        RECT 19.836 77.744 19.944 77.936 ; 
        RECT 20.448 77.744 20.592 77.936 ; 
        RECT 23.508 77.744 23.58 77.936 ; 
        RECT 37.764 77.744 37.836 77.936 ; 
        RECT 0.612 82.064 0.684 82.256 ; 
        RECT 14.868 82.064 14.94 82.256 ; 
        RECT 19.836 82.064 19.944 82.256 ; 
        RECT 20.448 82.064 20.592 82.256 ; 
        RECT 23.508 82.064 23.58 82.256 ; 
        RECT 37.764 82.064 37.836 82.256 ; 
        RECT 0.612 86.384 0.684 86.576 ; 
        RECT 14.868 86.384 14.94 86.576 ; 
        RECT 19.836 86.384 19.944 86.576 ; 
        RECT 20.448 86.384 20.592 86.576 ; 
        RECT 23.508 86.384 23.58 86.576 ; 
        RECT 37.764 86.384 37.836 86.576 ; 
        RECT 0.612 90.704 0.684 90.896 ; 
        RECT 14.868 90.704 14.94 90.896 ; 
        RECT 19.836 90.704 19.944 90.896 ; 
        RECT 20.448 90.704 20.592 90.896 ; 
        RECT 23.508 90.704 23.58 90.896 ; 
        RECT 37.764 90.704 37.836 90.896 ; 
        RECT 0.612 95.024 0.684 95.216 ; 
        RECT 14.868 95.024 14.94 95.216 ; 
        RECT 19.836 95.024 19.944 95.216 ; 
        RECT 20.448 95.024 20.592 95.216 ; 
        RECT 23.508 95.024 23.58 95.216 ; 
        RECT 37.764 95.024 37.836 95.216 ; 
        RECT 0.612 99.344 0.684 99.536 ; 
        RECT 14.868 99.344 14.94 99.536 ; 
        RECT 19.836 99.344 19.944 99.536 ; 
        RECT 20.448 99.344 20.592 99.536 ; 
        RECT 23.508 99.344 23.58 99.536 ; 
        RECT 37.764 99.344 37.836 99.536 ; 
        RECT 0.612 103.664 0.684 103.856 ; 
        RECT 14.868 103.664 14.94 103.856 ; 
        RECT 19.836 103.664 19.944 103.856 ; 
        RECT 20.448 103.664 20.592 103.856 ; 
        RECT 23.508 103.664 23.58 103.856 ; 
        RECT 37.764 103.664 37.836 103.856 ; 
        RECT 0.612 107.984 0.684 108.176 ; 
        RECT 14.868 107.984 14.94 108.176 ; 
        RECT 19.836 107.984 19.944 108.176 ; 
        RECT 20.448 107.984 20.592 108.176 ; 
        RECT 23.508 107.984 23.58 108.176 ; 
        RECT 37.764 107.984 37.836 108.176 ; 
        RECT 0.612 112.304 0.684 112.496 ; 
        RECT 14.868 112.304 14.94 112.496 ; 
        RECT 19.836 112.304 19.944 112.496 ; 
        RECT 20.448 112.304 20.592 112.496 ; 
        RECT 23.508 112.304 23.58 112.496 ; 
        RECT 37.764 112.304 37.836 112.496 ; 
        RECT 0.612 116.624 0.684 116.816 ; 
        RECT 14.868 116.624 14.94 116.816 ; 
        RECT 19.836 116.624 19.944 116.816 ; 
        RECT 20.448 116.624 20.592 116.816 ; 
        RECT 23.508 116.624 23.58 116.816 ; 
        RECT 37.764 116.624 37.836 116.816 ; 
        RECT 0.612 120.944 0.684 121.136 ; 
        RECT 14.868 120.944 14.94 121.136 ; 
        RECT 19.836 120.944 19.944 121.136 ; 
        RECT 20.448 120.944 20.592 121.136 ; 
        RECT 23.508 120.944 23.58 121.136 ; 
        RECT 37.764 120.944 37.836 121.136 ; 
        RECT 0.612 125.264 0.684 125.456 ; 
        RECT 14.868 125.264 14.94 125.456 ; 
        RECT 19.836 125.264 19.944 125.456 ; 
        RECT 20.448 125.264 20.592 125.456 ; 
        RECT 23.508 125.264 23.58 125.456 ; 
        RECT 37.764 125.264 37.836 125.456 ; 
        RECT 0.612 129.584 0.684 129.776 ; 
        RECT 14.868 129.584 14.94 129.776 ; 
        RECT 19.836 129.584 19.944 129.776 ; 
        RECT 20.448 129.584 20.592 129.776 ; 
        RECT 23.508 129.584 23.58 129.776 ; 
        RECT 37.764 129.584 37.836 129.776 ; 
        RECT 0.612 133.904 0.684 134.096 ; 
        RECT 14.868 133.904 14.94 134.096 ; 
        RECT 19.836 133.904 19.944 134.096 ; 
        RECT 20.448 133.904 20.592 134.096 ; 
        RECT 23.508 133.904 23.58 134.096 ; 
        RECT 37.764 133.904 37.836 134.096 ; 
        RECT 0.612 138.224 0.684 138.416 ; 
        RECT 14.868 138.224 14.94 138.416 ; 
        RECT 19.836 138.224 19.944 138.416 ; 
        RECT 20.448 138.224 20.592 138.416 ; 
        RECT 23.508 138.224 23.58 138.416 ; 
        RECT 37.764 138.224 37.836 138.416 ; 
        RECT 0.612 142.544 0.684 142.736 ; 
        RECT 14.868 142.544 14.94 142.736 ; 
        RECT 19.836 142.544 19.944 142.736 ; 
        RECT 20.448 142.544 20.592 142.736 ; 
        RECT 23.508 142.544 23.58 142.736 ; 
        RECT 37.764 142.544 37.836 142.736 ; 
        RECT 0.612 146.864 0.684 147.056 ; 
        RECT 14.868 146.864 14.94 147.056 ; 
        RECT 19.836 146.864 19.944 147.056 ; 
        RECT 20.448 146.864 20.592 147.056 ; 
        RECT 23.508 146.864 23.58 147.056 ; 
        RECT 37.764 146.864 37.836 147.056 ; 
        RECT 0.612 151.184 0.684 151.376 ; 
        RECT 14.868 151.184 14.94 151.376 ; 
        RECT 19.836 151.184 19.944 151.376 ; 
        RECT 20.448 151.184 20.592 151.376 ; 
        RECT 23.508 151.184 23.58 151.376 ; 
        RECT 37.764 151.184 37.836 151.376 ; 
        RECT 0.612 155.504 0.684 155.696 ; 
        RECT 14.868 155.504 14.94 155.696 ; 
        RECT 19.836 155.504 19.944 155.696 ; 
        RECT 20.448 155.504 20.592 155.696 ; 
        RECT 23.508 155.504 23.58 155.696 ; 
        RECT 37.764 155.504 37.836 155.696 ; 
        RECT 0.612 159.824 0.684 160.016 ; 
        RECT 14.868 159.824 14.94 160.016 ; 
        RECT 19.836 159.824 19.944 160.016 ; 
        RECT 20.448 159.824 20.592 160.016 ; 
        RECT 23.508 159.824 23.58 160.016 ; 
        RECT 37.764 159.824 37.836 160.016 ; 
        RECT 0.612 164.144 0.684 164.336 ; 
        RECT 14.868 164.144 14.94 164.336 ; 
        RECT 19.836 164.144 19.944 164.336 ; 
        RECT 20.448 164.144 20.592 164.336 ; 
        RECT 23.508 164.144 23.58 164.336 ; 
        RECT 37.764 164.144 37.836 164.336 ; 
        RECT 0.612 168.464 0.684 168.656 ; 
        RECT 14.868 168.464 14.94 168.656 ; 
        RECT 19.836 168.464 19.944 168.656 ; 
        RECT 20.448 168.464 20.592 168.656 ; 
        RECT 23.508 168.464 23.58 168.656 ; 
        RECT 37.764 168.464 37.836 168.656 ; 
        RECT 0.612 172.784 0.684 172.976 ; 
        RECT 14.868 172.784 14.94 172.976 ; 
        RECT 19.836 172.784 19.944 172.976 ; 
        RECT 20.448 172.784 20.592 172.976 ; 
        RECT 23.508 172.784 23.58 172.976 ; 
        RECT 37.764 172.784 37.836 172.976 ; 
        RECT 0.612 176.844 0.684 177.708 ; 
        RECT 19.708 202.188 19.78 203.052 ; 
        RECT 19.708 189.516 19.78 190.38 ; 
        RECT 19.708 176.844 19.78 177.708 ; 
        RECT 19.916 202.188 19.988 203.052 ; 
        RECT 19.916 189.516 19.988 190.38 ; 
        RECT 19.916 176.844 19.988 177.708 ; 
        RECT 20.124 202.188 20.196 203.052 ; 
        RECT 20.124 189.516 20.196 190.38 ; 
        RECT 20.124 176.844 20.196 177.708 ; 
        RECT 20.332 202.188 20.404 203.052 ; 
        RECT 20.332 189.516 20.404 190.38 ; 
        RECT 20.332 176.844 20.404 177.708 ; 
        RECT 20.54 202.188 20.612 203.052 ; 
        RECT 20.54 189.516 20.612 190.38 ; 
        RECT 20.54 176.844 20.612 177.708 ; 
        RECT 0.612 209.612 0.684 209.804 ; 
        RECT 14.868 209.612 14.94 209.804 ; 
        RECT 19.836 209.612 19.944 209.804 ; 
        RECT 20.448 209.612 20.592 209.804 ; 
        RECT 23.508 209.612 23.58 209.804 ; 
        RECT 37.764 209.612 37.836 209.804 ; 
        RECT 0.612 213.932 0.684 214.124 ; 
        RECT 14.868 213.932 14.94 214.124 ; 
        RECT 19.836 213.932 19.944 214.124 ; 
        RECT 20.448 213.932 20.592 214.124 ; 
        RECT 23.508 213.932 23.58 214.124 ; 
        RECT 37.764 213.932 37.836 214.124 ; 
        RECT 0.612 218.252 0.684 218.444 ; 
        RECT 14.868 218.252 14.94 218.444 ; 
        RECT 19.836 218.252 19.944 218.444 ; 
        RECT 20.448 218.252 20.592 218.444 ; 
        RECT 23.508 218.252 23.58 218.444 ; 
        RECT 37.764 218.252 37.836 218.444 ; 
        RECT 0.612 222.572 0.684 222.764 ; 
        RECT 14.868 222.572 14.94 222.764 ; 
        RECT 19.836 222.572 19.944 222.764 ; 
        RECT 20.448 222.572 20.592 222.764 ; 
        RECT 23.508 222.572 23.58 222.764 ; 
        RECT 37.764 222.572 37.836 222.764 ; 
        RECT 0.612 226.892 0.684 227.084 ; 
        RECT 14.868 226.892 14.94 227.084 ; 
        RECT 19.836 226.892 19.944 227.084 ; 
        RECT 20.448 226.892 20.592 227.084 ; 
        RECT 23.508 226.892 23.58 227.084 ; 
        RECT 37.764 226.892 37.836 227.084 ; 
        RECT 0.612 231.212 0.684 231.404 ; 
        RECT 14.868 231.212 14.94 231.404 ; 
        RECT 19.836 231.212 19.944 231.404 ; 
        RECT 20.448 231.212 20.592 231.404 ; 
        RECT 23.508 231.212 23.58 231.404 ; 
        RECT 37.764 231.212 37.836 231.404 ; 
        RECT 0.612 235.532 0.684 235.724 ; 
        RECT 14.868 235.532 14.94 235.724 ; 
        RECT 19.836 235.532 19.944 235.724 ; 
        RECT 20.448 235.532 20.592 235.724 ; 
        RECT 23.508 235.532 23.58 235.724 ; 
        RECT 37.764 235.532 37.836 235.724 ; 
        RECT 0.612 239.852 0.684 240.044 ; 
        RECT 14.868 239.852 14.94 240.044 ; 
        RECT 19.836 239.852 19.944 240.044 ; 
        RECT 20.448 239.852 20.592 240.044 ; 
        RECT 23.508 239.852 23.58 240.044 ; 
        RECT 37.764 239.852 37.836 240.044 ; 
        RECT 0.612 244.172 0.684 244.364 ; 
        RECT 14.868 244.172 14.94 244.364 ; 
        RECT 19.836 244.172 19.944 244.364 ; 
        RECT 20.448 244.172 20.592 244.364 ; 
        RECT 23.508 244.172 23.58 244.364 ; 
        RECT 37.764 244.172 37.836 244.364 ; 
        RECT 0.612 248.492 0.684 248.684 ; 
        RECT 14.868 248.492 14.94 248.684 ; 
        RECT 19.836 248.492 19.944 248.684 ; 
        RECT 20.448 248.492 20.592 248.684 ; 
        RECT 23.508 248.492 23.58 248.684 ; 
        RECT 37.764 248.492 37.836 248.684 ; 
        RECT 0.612 252.812 0.684 253.004 ; 
        RECT 14.868 252.812 14.94 253.004 ; 
        RECT 19.836 252.812 19.944 253.004 ; 
        RECT 20.448 252.812 20.592 253.004 ; 
        RECT 23.508 252.812 23.58 253.004 ; 
        RECT 37.764 252.812 37.836 253.004 ; 
        RECT 0.612 257.132 0.684 257.324 ; 
        RECT 14.868 257.132 14.94 257.324 ; 
        RECT 19.836 257.132 19.944 257.324 ; 
        RECT 20.448 257.132 20.592 257.324 ; 
        RECT 23.508 257.132 23.58 257.324 ; 
        RECT 37.764 257.132 37.836 257.324 ; 
        RECT 0.612 261.452 0.684 261.644 ; 
        RECT 14.868 261.452 14.94 261.644 ; 
        RECT 19.836 261.452 19.944 261.644 ; 
        RECT 20.448 261.452 20.592 261.644 ; 
        RECT 23.508 261.452 23.58 261.644 ; 
        RECT 37.764 261.452 37.836 261.644 ; 
        RECT 0.612 265.772 0.684 265.964 ; 
        RECT 14.868 265.772 14.94 265.964 ; 
        RECT 19.836 265.772 19.944 265.964 ; 
        RECT 20.448 265.772 20.592 265.964 ; 
        RECT 23.508 265.772 23.58 265.964 ; 
        RECT 37.764 265.772 37.836 265.964 ; 
        RECT 0.612 270.092 0.684 270.284 ; 
        RECT 14.868 270.092 14.94 270.284 ; 
        RECT 19.836 270.092 19.944 270.284 ; 
        RECT 20.448 270.092 20.592 270.284 ; 
        RECT 23.508 270.092 23.58 270.284 ; 
        RECT 37.764 270.092 37.836 270.284 ; 
        RECT 0.612 274.412 0.684 274.604 ; 
        RECT 14.868 274.412 14.94 274.604 ; 
        RECT 19.836 274.412 19.944 274.604 ; 
        RECT 20.448 274.412 20.592 274.604 ; 
        RECT 23.508 274.412 23.58 274.604 ; 
        RECT 37.764 274.412 37.836 274.604 ; 
        RECT 0.612 278.732 0.684 278.924 ; 
        RECT 14.868 278.732 14.94 278.924 ; 
        RECT 19.836 278.732 19.944 278.924 ; 
        RECT 20.448 278.732 20.592 278.924 ; 
        RECT 23.508 278.732 23.58 278.924 ; 
        RECT 37.764 278.732 37.836 278.924 ; 
        RECT 0.612 283.052 0.684 283.244 ; 
        RECT 14.868 283.052 14.94 283.244 ; 
        RECT 19.836 283.052 19.944 283.244 ; 
        RECT 20.448 283.052 20.592 283.244 ; 
        RECT 23.508 283.052 23.58 283.244 ; 
        RECT 37.764 283.052 37.836 283.244 ; 
        RECT 0.612 287.372 0.684 287.564 ; 
        RECT 14.868 287.372 14.94 287.564 ; 
        RECT 19.836 287.372 19.944 287.564 ; 
        RECT 20.448 287.372 20.592 287.564 ; 
        RECT 23.508 287.372 23.58 287.564 ; 
        RECT 37.764 287.372 37.836 287.564 ; 
        RECT 0.612 291.692 0.684 291.884 ; 
        RECT 14.868 291.692 14.94 291.884 ; 
        RECT 19.836 291.692 19.944 291.884 ; 
        RECT 20.448 291.692 20.592 291.884 ; 
        RECT 23.508 291.692 23.58 291.884 ; 
        RECT 37.764 291.692 37.836 291.884 ; 
        RECT 0.612 296.012 0.684 296.204 ; 
        RECT 14.868 296.012 14.94 296.204 ; 
        RECT 19.836 296.012 19.944 296.204 ; 
        RECT 20.448 296.012 20.592 296.204 ; 
        RECT 23.508 296.012 23.58 296.204 ; 
        RECT 37.764 296.012 37.836 296.204 ; 
        RECT 0.612 300.332 0.684 300.524 ; 
        RECT 14.868 300.332 14.94 300.524 ; 
        RECT 19.836 300.332 19.944 300.524 ; 
        RECT 20.448 300.332 20.592 300.524 ; 
        RECT 23.508 300.332 23.58 300.524 ; 
        RECT 37.764 300.332 37.836 300.524 ; 
        RECT 0.612 304.652 0.684 304.844 ; 
        RECT 14.868 304.652 14.94 304.844 ; 
        RECT 19.836 304.652 19.944 304.844 ; 
        RECT 20.448 304.652 20.592 304.844 ; 
        RECT 23.508 304.652 23.58 304.844 ; 
        RECT 37.764 304.652 37.836 304.844 ; 
        RECT 0.612 308.972 0.684 309.164 ; 
        RECT 14.868 308.972 14.94 309.164 ; 
        RECT 19.836 308.972 19.944 309.164 ; 
        RECT 20.448 308.972 20.592 309.164 ; 
        RECT 23.508 308.972 23.58 309.164 ; 
        RECT 37.764 308.972 37.836 309.164 ; 
        RECT 0.612 313.292 0.684 313.484 ; 
        RECT 14.868 313.292 14.94 313.484 ; 
        RECT 19.836 313.292 19.944 313.484 ; 
        RECT 20.448 313.292 20.592 313.484 ; 
        RECT 23.508 313.292 23.58 313.484 ; 
        RECT 37.764 313.292 37.836 313.484 ; 
        RECT 0.612 317.612 0.684 317.804 ; 
        RECT 14.868 317.612 14.94 317.804 ; 
        RECT 19.836 317.612 19.944 317.804 ; 
        RECT 20.448 317.612 20.592 317.804 ; 
        RECT 23.508 317.612 23.58 317.804 ; 
        RECT 37.764 317.612 37.836 317.804 ; 
        RECT 0.612 321.932 0.684 322.124 ; 
        RECT 14.868 321.932 14.94 322.124 ; 
        RECT 19.836 321.932 19.944 322.124 ; 
        RECT 20.448 321.932 20.592 322.124 ; 
        RECT 23.508 321.932 23.58 322.124 ; 
        RECT 37.764 321.932 37.836 322.124 ; 
        RECT 0.612 326.252 0.684 326.444 ; 
        RECT 14.868 326.252 14.94 326.444 ; 
        RECT 19.836 326.252 19.944 326.444 ; 
        RECT 20.448 326.252 20.592 326.444 ; 
        RECT 23.508 326.252 23.58 326.444 ; 
        RECT 37.764 326.252 37.836 326.444 ; 
        RECT 0.612 330.572 0.684 330.764 ; 
        RECT 14.868 330.572 14.94 330.764 ; 
        RECT 19.836 330.572 19.944 330.764 ; 
        RECT 20.448 330.572 20.592 330.764 ; 
        RECT 23.508 330.572 23.58 330.764 ; 
        RECT 37.764 330.572 37.836 330.764 ; 
        RECT 0.612 334.892 0.684 335.084 ; 
        RECT 14.868 334.892 14.94 335.084 ; 
        RECT 19.836 334.892 19.944 335.084 ; 
        RECT 20.448 334.892 20.592 335.084 ; 
        RECT 23.508 334.892 23.58 335.084 ; 
        RECT 37.764 334.892 37.836 335.084 ; 
        RECT 0.612 339.212 0.684 339.404 ; 
        RECT 14.868 339.212 14.94 339.404 ; 
        RECT 19.836 339.212 19.944 339.404 ; 
        RECT 20.448 339.212 20.592 339.404 ; 
        RECT 23.508 339.212 23.58 339.404 ; 
        RECT 37.764 339.212 37.836 339.404 ; 
        RECT 0.612 343.532 0.684 343.724 ; 
        RECT 14.868 343.532 14.94 343.724 ; 
        RECT 19.836 343.532 19.944 343.724 ; 
        RECT 20.448 343.532 20.592 343.724 ; 
        RECT 23.508 343.532 23.58 343.724 ; 
        RECT 37.764 343.532 37.836 343.724 ; 
        RECT 0.612 347.852 0.684 348.044 ; 
        RECT 14.868 347.852 14.94 348.044 ; 
        RECT 19.836 347.852 19.944 348.044 ; 
        RECT 20.448 347.852 20.592 348.044 ; 
        RECT 23.508 347.852 23.58 348.044 ; 
        RECT 37.764 347.852 37.836 348.044 ; 
        RECT 0.612 352.172 0.684 352.364 ; 
        RECT 14.868 352.172 14.94 352.364 ; 
        RECT 19.836 352.172 19.944 352.364 ; 
        RECT 20.448 352.172 20.592 352.364 ; 
        RECT 23.508 352.172 23.58 352.364 ; 
        RECT 37.764 352.172 37.836 352.364 ; 
        RECT 0.612 356.492 0.684 356.684 ; 
        RECT 14.868 356.492 14.94 356.684 ; 
        RECT 19.836 356.492 19.944 356.684 ; 
        RECT 20.448 356.492 20.592 356.684 ; 
        RECT 23.508 356.492 23.58 356.684 ; 
        RECT 37.764 356.492 37.836 356.684 ; 
        RECT 0.612 360.812 0.684 361.004 ; 
        RECT 14.868 360.812 14.94 361.004 ; 
        RECT 19.836 360.812 19.944 361.004 ; 
        RECT 20.448 360.812 20.592 361.004 ; 
        RECT 23.508 360.812 23.58 361.004 ; 
        RECT 37.764 360.812 37.836 361.004 ; 
        RECT 0.612 365.132 0.684 365.324 ; 
        RECT 14.868 365.132 14.94 365.324 ; 
        RECT 19.836 365.132 19.944 365.324 ; 
        RECT 20.448 365.132 20.592 365.324 ; 
        RECT 23.508 365.132 23.58 365.324 ; 
        RECT 37.764 365.132 37.836 365.324 ; 
        RECT 0.612 369.452 0.684 369.644 ; 
        RECT 14.868 369.452 14.94 369.644 ; 
        RECT 19.836 369.452 19.944 369.644 ; 
        RECT 20.448 369.452 20.592 369.644 ; 
        RECT 23.508 369.452 23.58 369.644 ; 
        RECT 37.764 369.452 37.836 369.644 ; 
        RECT 0.612 373.772 0.684 373.964 ; 
        RECT 14.868 373.772 14.94 373.964 ; 
        RECT 19.836 373.772 19.944 373.964 ; 
        RECT 20.448 373.772 20.592 373.964 ; 
        RECT 23.508 373.772 23.58 373.964 ; 
        RECT 37.764 373.772 37.836 373.964 ; 
        RECT 0.612 378.092 0.684 378.284 ; 
        RECT 14.868 378.092 14.94 378.284 ; 
        RECT 19.836 378.092 19.944 378.284 ; 
        RECT 20.448 378.092 20.592 378.284 ; 
        RECT 23.508 378.092 23.58 378.284 ; 
        RECT 37.764 378.092 37.836 378.284 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.34 178.732 29.412 178.88 ; 
      LAYER M4 ; 
        RECT 29.132 178.764 29.468 178.86 ; 
      LAYER M5 ; 
        RECT 29.328 174.96 29.424 187.92 ; 
      LAYER V3 ; 
        RECT 29.34 178.764 29.412 178.86 ; 
      LAYER V4 ; 
        RECT 29.328 178.764 29.424 178.86 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.476 178.744 28.548 178.892 ; 
      LAYER M4 ; 
        RECT 28.268 178.764 28.604 178.86 ; 
      LAYER M5 ; 
        RECT 28.464 174.96 28.56 187.92 ; 
      LAYER V3 ; 
        RECT 28.476 178.764 28.548 178.86 ; 
      LAYER V4 ; 
        RECT 28.464 178.764 28.56 178.86 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.612 176.428 27.684 176.576 ; 
      LAYER M4 ; 
        RECT 27.404 176.46 27.74 176.556 ; 
      LAYER M5 ; 
        RECT 27.6 174.96 27.696 187.92 ; 
      LAYER V3 ; 
        RECT 27.612 176.46 27.684 176.556 ; 
      LAYER V4 ; 
        RECT 27.6 176.46 27.696 176.556 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.748 177.388 26.82 178.112 ; 
      LAYER M4 ; 
        RECT 26.54 177.996 26.876 178.092 ; 
      LAYER M5 ; 
        RECT 26.736 174.96 26.832 187.92 ; 
      LAYER V3 ; 
        RECT 26.748 177.996 26.82 178.092 ; 
      LAYER V4 ; 
        RECT 26.736 177.996 26.832 178.092 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.884 176.44 25.956 176.708 ; 
      LAYER M4 ; 
        RECT 25.676 176.46 26.012 176.556 ; 
      LAYER M5 ; 
        RECT 25.872 174.96 25.968 187.92 ; 
      LAYER V3 ; 
        RECT 25.884 176.46 25.956 176.556 ; 
      LAYER V4 ; 
        RECT 25.872 176.46 25.968 176.556 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.02 175.372 25.092 176.384 ; 
      LAYER M4 ; 
        RECT 24.812 176.268 25.148 176.364 ; 
      LAYER M5 ; 
        RECT 25.008 174.96 25.104 187.92 ; 
      LAYER V3 ; 
        RECT 25.02 176.268 25.092 176.364 ; 
      LAYER V4 ; 
        RECT 25.008 176.268 25.104 176.364 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.156 179.512 24.228 179.66 ; 
      LAYER M4 ; 
        RECT 23.948 179.532 24.284 179.628 ; 
      LAYER M5 ; 
        RECT 24.144 174.96 24.24 187.92 ; 
      LAYER V3 ; 
        RECT 24.156 179.532 24.228 179.628 ; 
      LAYER V4 ; 
        RECT 24.144 179.532 24.24 179.628 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 20.7 176.44 20.772 176.708 ; 
      LAYER M4 ; 
        RECT 19.564 176.46 20.816 176.556 ; 
      LAYER M5 ; 
        RECT 19.608 174.96 19.704 187.92 ; 
      LAYER V3 ; 
        RECT 20.7 176.46 20.772 176.556 ; 
      LAYER V4 ; 
        RECT 19.608 176.46 19.704 176.556 ; 
    END 
  END ADDRESS[7] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 19.116 175.372 19.188 176.384 ; 
      LAYER M4 ; 
        RECT 18.268 176.268 19.232 176.364 ; 
      LAYER M5 ; 
        RECT 18.312 174.96 18.408 187.92 ; 
      LAYER V3 ; 
        RECT 19.116 176.268 19.188 176.364 ; 
      LAYER V4 ; 
        RECT 18.312 176.268 18.408 176.364 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.948 176.44 16.02 176.708 ; 
      LAYER M4 ; 
        RECT 15.74 176.46 16.076 176.556 ; 
      LAYER M5 ; 
        RECT 15.936 174.96 16.032 187.92 ; 
      LAYER V3 ; 
        RECT 15.948 176.46 16.02 176.556 ; 
      LAYER V4 ; 
        RECT 15.936 176.46 16.032 176.556 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.084 179.896 15.156 180.092 ; 
      LAYER M4 ; 
        RECT 14.876 179.916 15.212 180.012 ; 
      LAYER M5 ; 
        RECT 15.072 174.96 15.168 187.92 ; 
      LAYER V3 ; 
        RECT 15.084 179.916 15.156 180.012 ; 
      LAYER V4 ; 
        RECT 15.072 179.916 15.168 180.012 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.228 175.372 15.3 176.384 ; 
      LAYER M4 ; 
        RECT 14.164 176.268 15.344 176.364 ; 
      LAYER M5 ; 
        RECT 14.208 174.96 14.304 187.92 ; 
      LAYER V3 ; 
        RECT 15.228 176.268 15.3 176.364 ; 
      LAYER V4 ; 
        RECT 14.208 176.268 14.304 176.364 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 13.356 178.732 13.428 178.88 ; 
      LAYER M4 ; 
        RECT 13.148 178.764 13.484 178.86 ; 
      LAYER M5 ; 
        RECT 13.344 174.96 13.44 187.92 ; 
      LAYER V3 ; 
        RECT 13.356 178.764 13.428 178.86 ; 
      LAYER V4 ; 
        RECT 13.344 178.764 13.44 178.86 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 12.492 176.44 12.564 177.356 ; 
      LAYER M4 ; 
        RECT 12.284 176.46 12.62 176.556 ; 
      LAYER M5 ; 
        RECT 12.48 174.96 12.576 187.92 ; 
      LAYER V3 ; 
        RECT 12.492 176.46 12.564 176.556 ; 
      LAYER V4 ; 
        RECT 12.48 176.46 12.576 176.556 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 11.628 175.372 11.7 176.384 ; 
      LAYER M4 ; 
        RECT 11.42 176.268 11.756 176.364 ; 
      LAYER M5 ; 
        RECT 11.616 174.96 11.712 187.92 ; 
      LAYER V3 ; 
        RECT 11.628 176.268 11.7 176.364 ; 
      LAYER V4 ; 
        RECT 11.616 176.268 11.712 176.364 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 10.764 176.428 10.836 176.576 ; 
      LAYER M4 ; 
        RECT 10.556 176.46 10.892 176.556 ; 
      LAYER M5 ; 
        RECT 10.752 174.96 10.848 187.92 ; 
      LAYER V3 ; 
        RECT 10.764 176.46 10.836 176.556 ; 
      LAYER V4 ; 
        RECT 10.752 176.46 10.848 176.556 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 9.9 178.732 9.972 178.88 ; 
      LAYER M4 ; 
        RECT 9.692 178.764 10.028 178.86 ; 
      LAYER M5 ; 
        RECT 9.888 174.96 9.984 187.92 ; 
      LAYER V3 ; 
        RECT 9.9 178.764 9.972 178.86 ; 
      LAYER V4 ; 
        RECT 9.888 178.764 9.984 178.86 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.712 20.544 1.808 ; 
      LAYER M3 ; 
        RECT 20.304 1.51 20.376 2.468 ; 
      LAYER V3 ; 
        RECT 20.304 1.712 20.376 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.328 20.816 1.424 ; 
      LAYER M3 ; 
        RECT 19.404 1.08 19.476 2.7 ; 
      LAYER V3 ; 
        RECT 19.404 1.328 19.476 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 6.032 20.544 6.128 ; 
      LAYER M3 ; 
        RECT 20.304 5.83 20.376 6.788 ; 
      LAYER V3 ; 
        RECT 20.304 6.032 20.376 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 5.648 20.816 5.744 ; 
      LAYER M3 ; 
        RECT 19.404 5.4 19.476 7.02 ; 
      LAYER V3 ; 
        RECT 19.404 5.648 19.476 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 10.352 20.544 10.448 ; 
      LAYER M3 ; 
        RECT 20.304 10.15 20.376 11.108 ; 
      LAYER V3 ; 
        RECT 20.304 10.352 20.376 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 9.968 20.816 10.064 ; 
      LAYER M3 ; 
        RECT 19.404 9.72 19.476 11.34 ; 
      LAYER V3 ; 
        RECT 19.404 9.968 19.476 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.672 20.544 14.768 ; 
      LAYER M3 ; 
        RECT 20.304 14.47 20.376 15.428 ; 
      LAYER V3 ; 
        RECT 20.304 14.672 20.376 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.288 20.816 14.384 ; 
      LAYER M3 ; 
        RECT 19.404 14.04 19.476 15.66 ; 
      LAYER V3 ; 
        RECT 19.404 14.288 19.476 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.992 20.544 19.088 ; 
      LAYER M3 ; 
        RECT 20.304 18.79 20.376 19.748 ; 
      LAYER V3 ; 
        RECT 20.304 18.992 20.376 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.608 20.816 18.704 ; 
      LAYER M3 ; 
        RECT 19.404 18.36 19.476 19.98 ; 
      LAYER V3 ; 
        RECT 19.404 18.608 19.476 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 23.312 20.544 23.408 ; 
      LAYER M3 ; 
        RECT 20.304 23.11 20.376 24.068 ; 
      LAYER V3 ; 
        RECT 20.304 23.312 20.376 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 22.928 20.816 23.024 ; 
      LAYER M3 ; 
        RECT 19.404 22.68 19.476 24.3 ; 
      LAYER V3 ; 
        RECT 19.404 22.928 19.476 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.632 20.544 27.728 ; 
      LAYER M3 ; 
        RECT 20.304 27.43 20.376 28.388 ; 
      LAYER V3 ; 
        RECT 20.304 27.632 20.376 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.248 20.816 27.344 ; 
      LAYER M3 ; 
        RECT 19.404 27 19.476 28.62 ; 
      LAYER V3 ; 
        RECT 19.404 27.248 19.476 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.952 20.544 32.048 ; 
      LAYER M3 ; 
        RECT 20.304 31.75 20.376 32.708 ; 
      LAYER V3 ; 
        RECT 20.304 31.952 20.376 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.568 20.816 31.664 ; 
      LAYER M3 ; 
        RECT 19.404 31.32 19.476 32.94 ; 
      LAYER V3 ; 
        RECT 19.404 31.568 19.476 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 36.272 20.544 36.368 ; 
      LAYER M3 ; 
        RECT 20.304 36.07 20.376 37.028 ; 
      LAYER V3 ; 
        RECT 20.304 36.272 20.376 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 35.888 20.816 35.984 ; 
      LAYER M3 ; 
        RECT 19.404 35.64 19.476 37.26 ; 
      LAYER V3 ; 
        RECT 19.404 35.888 19.476 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 40.592 20.544 40.688 ; 
      LAYER M3 ; 
        RECT 20.304 40.39 20.376 41.348 ; 
      LAYER V3 ; 
        RECT 20.304 40.592 20.376 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 40.208 20.816 40.304 ; 
      LAYER M3 ; 
        RECT 19.404 39.96 19.476 41.58 ; 
      LAYER V3 ; 
        RECT 19.404 40.208 19.476 40.304 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 44.912 20.544 45.008 ; 
      LAYER M3 ; 
        RECT 20.304 44.71 20.376 45.668 ; 
      LAYER V3 ; 
        RECT 20.304 44.912 20.376 45.008 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 44.528 20.816 44.624 ; 
      LAYER M3 ; 
        RECT 19.404 44.28 19.476 45.9 ; 
      LAYER V3 ; 
        RECT 19.404 44.528 19.476 44.624 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 49.232 20.544 49.328 ; 
      LAYER M3 ; 
        RECT 20.304 49.03 20.376 49.988 ; 
      LAYER V3 ; 
        RECT 20.304 49.232 20.376 49.328 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 48.848 20.816 48.944 ; 
      LAYER M3 ; 
        RECT 19.404 48.6 19.476 50.22 ; 
      LAYER V3 ; 
        RECT 19.404 48.848 19.476 48.944 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 53.552 20.544 53.648 ; 
      LAYER M3 ; 
        RECT 20.304 53.35 20.376 54.308 ; 
      LAYER V3 ; 
        RECT 20.304 53.552 20.376 53.648 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 53.168 20.816 53.264 ; 
      LAYER M3 ; 
        RECT 19.404 52.92 19.476 54.54 ; 
      LAYER V3 ; 
        RECT 19.404 53.168 19.476 53.264 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 57.872 20.544 57.968 ; 
      LAYER M3 ; 
        RECT 20.304 57.67 20.376 58.628 ; 
      LAYER V3 ; 
        RECT 20.304 57.872 20.376 57.968 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 57.488 20.816 57.584 ; 
      LAYER M3 ; 
        RECT 19.404 57.24 19.476 58.86 ; 
      LAYER V3 ; 
        RECT 19.404 57.488 19.476 57.584 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 62.192 20.544 62.288 ; 
      LAYER M3 ; 
        RECT 20.304 61.99 20.376 62.948 ; 
      LAYER V3 ; 
        RECT 20.304 62.192 20.376 62.288 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 61.808 20.816 61.904 ; 
      LAYER M3 ; 
        RECT 19.404 61.56 19.476 63.18 ; 
      LAYER V3 ; 
        RECT 19.404 61.808 19.476 61.904 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 66.512 20.544 66.608 ; 
      LAYER M3 ; 
        RECT 20.304 66.31 20.376 67.268 ; 
      LAYER V3 ; 
        RECT 20.304 66.512 20.376 66.608 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 66.128 20.816 66.224 ; 
      LAYER M3 ; 
        RECT 19.404 65.88 19.476 67.5 ; 
      LAYER V3 ; 
        RECT 19.404 66.128 19.476 66.224 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 70.832 20.544 70.928 ; 
      LAYER M3 ; 
        RECT 20.304 70.63 20.376 71.588 ; 
      LAYER V3 ; 
        RECT 20.304 70.832 20.376 70.928 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 70.448 20.816 70.544 ; 
      LAYER M3 ; 
        RECT 19.404 70.2 19.476 71.82 ; 
      LAYER V3 ; 
        RECT 19.404 70.448 19.476 70.544 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 75.152 20.544 75.248 ; 
      LAYER M3 ; 
        RECT 20.304 74.95 20.376 75.908 ; 
      LAYER V3 ; 
        RECT 20.304 75.152 20.376 75.248 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 74.768 20.816 74.864 ; 
      LAYER M3 ; 
        RECT 19.404 74.52 19.476 76.14 ; 
      LAYER V3 ; 
        RECT 19.404 74.768 19.476 74.864 ; 
    END 
  END wd[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 79.472 20.544 79.568 ; 
      LAYER M3 ; 
        RECT 20.304 79.27 20.376 80.228 ; 
      LAYER V3 ; 
        RECT 20.304 79.472 20.376 79.568 ; 
    END 
  END dataout[18] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 79.088 20.816 79.184 ; 
      LAYER M3 ; 
        RECT 19.404 78.84 19.476 80.46 ; 
      LAYER V3 ; 
        RECT 19.404 79.088 19.476 79.184 ; 
    END 
  END wd[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 83.792 20.544 83.888 ; 
      LAYER M3 ; 
        RECT 20.304 83.59 20.376 84.548 ; 
      LAYER V3 ; 
        RECT 20.304 83.792 20.376 83.888 ; 
    END 
  END dataout[19] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 83.408 20.816 83.504 ; 
      LAYER M3 ; 
        RECT 19.404 83.16 19.476 84.78 ; 
      LAYER V3 ; 
        RECT 19.404 83.408 19.476 83.504 ; 
    END 
  END wd[19] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 88.112 20.544 88.208 ; 
      LAYER M3 ; 
        RECT 20.304 87.91 20.376 88.868 ; 
      LAYER V3 ; 
        RECT 20.304 88.112 20.376 88.208 ; 
    END 
  END dataout[20] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 87.728 20.816 87.824 ; 
      LAYER M3 ; 
        RECT 19.404 87.48 19.476 89.1 ; 
      LAYER V3 ; 
        RECT 19.404 87.728 19.476 87.824 ; 
    END 
  END wd[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 92.432 20.544 92.528 ; 
      LAYER M3 ; 
        RECT 20.304 92.23 20.376 93.188 ; 
      LAYER V3 ; 
        RECT 20.304 92.432 20.376 92.528 ; 
    END 
  END dataout[21] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 92.048 20.816 92.144 ; 
      LAYER M3 ; 
        RECT 19.404 91.8 19.476 93.42 ; 
      LAYER V3 ; 
        RECT 19.404 92.048 19.476 92.144 ; 
    END 
  END wd[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 96.752 20.544 96.848 ; 
      LAYER M3 ; 
        RECT 20.304 96.55 20.376 97.508 ; 
      LAYER V3 ; 
        RECT 20.304 96.752 20.376 96.848 ; 
    END 
  END dataout[22] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 96.368 20.816 96.464 ; 
      LAYER M3 ; 
        RECT 19.404 96.12 19.476 97.74 ; 
      LAYER V3 ; 
        RECT 19.404 96.368 19.476 96.464 ; 
    END 
  END wd[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 101.072 20.544 101.168 ; 
      LAYER M3 ; 
        RECT 20.304 100.87 20.376 101.828 ; 
      LAYER V3 ; 
        RECT 20.304 101.072 20.376 101.168 ; 
    END 
  END dataout[23] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 100.688 20.816 100.784 ; 
      LAYER M3 ; 
        RECT 19.404 100.44 19.476 102.06 ; 
      LAYER V3 ; 
        RECT 19.404 100.688 19.476 100.784 ; 
    END 
  END wd[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 105.392 20.544 105.488 ; 
      LAYER M3 ; 
        RECT 20.304 105.19 20.376 106.148 ; 
      LAYER V3 ; 
        RECT 20.304 105.392 20.376 105.488 ; 
    END 
  END dataout[24] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 105.008 20.816 105.104 ; 
      LAYER M3 ; 
        RECT 19.404 104.76 19.476 106.38 ; 
      LAYER V3 ; 
        RECT 19.404 105.008 19.476 105.104 ; 
    END 
  END wd[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 109.712 20.544 109.808 ; 
      LAYER M3 ; 
        RECT 20.304 109.51 20.376 110.468 ; 
      LAYER V3 ; 
        RECT 20.304 109.712 20.376 109.808 ; 
    END 
  END dataout[25] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 109.328 20.816 109.424 ; 
      LAYER M3 ; 
        RECT 19.404 109.08 19.476 110.7 ; 
      LAYER V3 ; 
        RECT 19.404 109.328 19.476 109.424 ; 
    END 
  END wd[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 114.032 20.544 114.128 ; 
      LAYER M3 ; 
        RECT 20.304 113.83 20.376 114.788 ; 
      LAYER V3 ; 
        RECT 20.304 114.032 20.376 114.128 ; 
    END 
  END dataout[26] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 113.648 20.816 113.744 ; 
      LAYER M3 ; 
        RECT 19.404 113.4 19.476 115.02 ; 
      LAYER V3 ; 
        RECT 19.404 113.648 19.476 113.744 ; 
    END 
  END wd[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 118.352 20.544 118.448 ; 
      LAYER M3 ; 
        RECT 20.304 118.15 20.376 119.108 ; 
      LAYER V3 ; 
        RECT 20.304 118.352 20.376 118.448 ; 
    END 
  END dataout[27] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 117.968 20.816 118.064 ; 
      LAYER M3 ; 
        RECT 19.404 117.72 19.476 119.34 ; 
      LAYER V3 ; 
        RECT 19.404 117.968 19.476 118.064 ; 
    END 
  END wd[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 122.672 20.544 122.768 ; 
      LAYER M3 ; 
        RECT 20.304 122.47 20.376 123.428 ; 
      LAYER V3 ; 
        RECT 20.304 122.672 20.376 122.768 ; 
    END 
  END dataout[28] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 122.288 20.816 122.384 ; 
      LAYER M3 ; 
        RECT 19.404 122.04 19.476 123.66 ; 
      LAYER V3 ; 
        RECT 19.404 122.288 19.476 122.384 ; 
    END 
  END wd[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 126.992 20.544 127.088 ; 
      LAYER M3 ; 
        RECT 20.304 126.79 20.376 127.748 ; 
      LAYER V3 ; 
        RECT 20.304 126.992 20.376 127.088 ; 
    END 
  END dataout[29] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 126.608 20.816 126.704 ; 
      LAYER M3 ; 
        RECT 19.404 126.36 19.476 127.98 ; 
      LAYER V3 ; 
        RECT 19.404 126.608 19.476 126.704 ; 
    END 
  END wd[29] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 131.312 20.544 131.408 ; 
      LAYER M3 ; 
        RECT 20.304 131.11 20.376 132.068 ; 
      LAYER V3 ; 
        RECT 20.304 131.312 20.376 131.408 ; 
    END 
  END dataout[30] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 130.928 20.816 131.024 ; 
      LAYER M3 ; 
        RECT 19.404 130.68 19.476 132.3 ; 
      LAYER V3 ; 
        RECT 19.404 130.928 19.476 131.024 ; 
    END 
  END wd[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 135.632 20.544 135.728 ; 
      LAYER M3 ; 
        RECT 20.304 135.43 20.376 136.388 ; 
      LAYER V3 ; 
        RECT 20.304 135.632 20.376 135.728 ; 
    END 
  END dataout[31] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 135.248 20.816 135.344 ; 
      LAYER M3 ; 
        RECT 19.404 135 19.476 136.62 ; 
      LAYER V3 ; 
        RECT 19.404 135.248 19.476 135.344 ; 
    END 
  END wd[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 139.952 20.544 140.048 ; 
      LAYER M3 ; 
        RECT 20.304 139.75 20.376 140.708 ; 
      LAYER V3 ; 
        RECT 20.304 139.952 20.376 140.048 ; 
    END 
  END dataout[32] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 139.568 20.816 139.664 ; 
      LAYER M3 ; 
        RECT 19.404 139.32 19.476 140.94 ; 
      LAYER V3 ; 
        RECT 19.404 139.568 19.476 139.664 ; 
    END 
  END wd[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 144.272 20.544 144.368 ; 
      LAYER M3 ; 
        RECT 20.304 144.07 20.376 145.028 ; 
      LAYER V3 ; 
        RECT 20.304 144.272 20.376 144.368 ; 
    END 
  END dataout[33] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 143.888 20.816 143.984 ; 
      LAYER M3 ; 
        RECT 19.404 143.64 19.476 145.26 ; 
      LAYER V3 ; 
        RECT 19.404 143.888 19.476 143.984 ; 
    END 
  END wd[33] 
  PIN dataout[34] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 148.592 20.544 148.688 ; 
      LAYER M3 ; 
        RECT 20.304 148.39 20.376 149.348 ; 
      LAYER V3 ; 
        RECT 20.304 148.592 20.376 148.688 ; 
    END 
  END dataout[34] 
  PIN wd[34] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 148.208 20.816 148.304 ; 
      LAYER M3 ; 
        RECT 19.404 147.96 19.476 149.58 ; 
      LAYER V3 ; 
        RECT 19.404 148.208 19.476 148.304 ; 
    END 
  END wd[34] 
  PIN dataout[35] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 152.912 20.544 153.008 ; 
      LAYER M3 ; 
        RECT 20.304 152.71 20.376 153.668 ; 
      LAYER V3 ; 
        RECT 20.304 152.912 20.376 153.008 ; 
    END 
  END dataout[35] 
  PIN wd[35] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 152.528 20.816 152.624 ; 
      LAYER M3 ; 
        RECT 19.404 152.28 19.476 153.9 ; 
      LAYER V3 ; 
        RECT 19.404 152.528 19.476 152.624 ; 
    END 
  END wd[35] 
  PIN dataout[36] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 157.232 20.544 157.328 ; 
      LAYER M3 ; 
        RECT 20.304 157.03 20.376 157.988 ; 
      LAYER V3 ; 
        RECT 20.304 157.232 20.376 157.328 ; 
    END 
  END dataout[36] 
  PIN wd[36] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 156.848 20.816 156.944 ; 
      LAYER M3 ; 
        RECT 19.404 156.6 19.476 158.22 ; 
      LAYER V3 ; 
        RECT 19.404 156.848 19.476 156.944 ; 
    END 
  END wd[36] 
  PIN dataout[37] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 161.552 20.544 161.648 ; 
      LAYER M3 ; 
        RECT 20.304 161.35 20.376 162.308 ; 
      LAYER V3 ; 
        RECT 20.304 161.552 20.376 161.648 ; 
    END 
  END dataout[37] 
  PIN wd[37] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 161.168 20.816 161.264 ; 
      LAYER M3 ; 
        RECT 19.404 160.92 19.476 162.54 ; 
      LAYER V3 ; 
        RECT 19.404 161.168 19.476 161.264 ; 
    END 
  END wd[37] 
  PIN dataout[38] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 165.872 20.544 165.968 ; 
      LAYER M3 ; 
        RECT 20.304 165.67 20.376 166.628 ; 
      LAYER V3 ; 
        RECT 20.304 165.872 20.376 165.968 ; 
    END 
  END dataout[38] 
  PIN wd[38] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 165.488 20.816 165.584 ; 
      LAYER M3 ; 
        RECT 19.404 165.24 19.476 166.86 ; 
      LAYER V3 ; 
        RECT 19.404 165.488 19.476 165.584 ; 
    END 
  END wd[38] 
  PIN dataout[39] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 170.192 20.544 170.288 ; 
      LAYER M3 ; 
        RECT 20.304 169.99 20.376 170.948 ; 
      LAYER V3 ; 
        RECT 20.304 170.192 20.376 170.288 ; 
    END 
  END dataout[39] 
  PIN wd[39] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 169.808 20.816 169.904 ; 
      LAYER M3 ; 
        RECT 19.404 169.56 19.476 171.18 ; 
      LAYER V3 ; 
        RECT 19.404 169.808 19.476 169.904 ; 
    END 
  END wd[39] 
  PIN dataout[40] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 207.02 20.544 207.116 ; 
      LAYER M3 ; 
        RECT 20.304 206.818 20.376 207.776 ; 
      LAYER V3 ; 
        RECT 20.304 207.02 20.376 207.116 ; 
    END 
  END dataout[40] 
  PIN wd[40] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 206.636 20.816 206.732 ; 
      LAYER M3 ; 
        RECT 19.404 206.388 19.476 208.008 ; 
      LAYER V3 ; 
        RECT 19.404 206.636 19.476 206.732 ; 
    END 
  END wd[40] 
  PIN dataout[41] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 211.34 20.544 211.436 ; 
      LAYER M3 ; 
        RECT 20.304 211.138 20.376 212.096 ; 
      LAYER V3 ; 
        RECT 20.304 211.34 20.376 211.436 ; 
    END 
  END dataout[41] 
  PIN wd[41] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 210.956 20.816 211.052 ; 
      LAYER M3 ; 
        RECT 19.404 210.708 19.476 212.328 ; 
      LAYER V3 ; 
        RECT 19.404 210.956 19.476 211.052 ; 
    END 
  END wd[41] 
  PIN dataout[42] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 215.66 20.544 215.756 ; 
      LAYER M3 ; 
        RECT 20.304 215.458 20.376 216.416 ; 
      LAYER V3 ; 
        RECT 20.304 215.66 20.376 215.756 ; 
    END 
  END dataout[42] 
  PIN wd[42] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 215.276 20.816 215.372 ; 
      LAYER M3 ; 
        RECT 19.404 215.028 19.476 216.648 ; 
      LAYER V3 ; 
        RECT 19.404 215.276 19.476 215.372 ; 
    END 
  END wd[42] 
  PIN dataout[43] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 219.98 20.544 220.076 ; 
      LAYER M3 ; 
        RECT 20.304 219.778 20.376 220.736 ; 
      LAYER V3 ; 
        RECT 20.304 219.98 20.376 220.076 ; 
    END 
  END dataout[43] 
  PIN wd[43] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 219.596 20.816 219.692 ; 
      LAYER M3 ; 
        RECT 19.404 219.348 19.476 220.968 ; 
      LAYER V3 ; 
        RECT 19.404 219.596 19.476 219.692 ; 
    END 
  END wd[43] 
  PIN dataout[44] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 224.3 20.544 224.396 ; 
      LAYER M3 ; 
        RECT 20.304 224.098 20.376 225.056 ; 
      LAYER V3 ; 
        RECT 20.304 224.3 20.376 224.396 ; 
    END 
  END dataout[44] 
  PIN wd[44] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 223.916 20.816 224.012 ; 
      LAYER M3 ; 
        RECT 19.404 223.668 19.476 225.288 ; 
      LAYER V3 ; 
        RECT 19.404 223.916 19.476 224.012 ; 
    END 
  END wd[44] 
  PIN dataout[45] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 228.62 20.544 228.716 ; 
      LAYER M3 ; 
        RECT 20.304 228.418 20.376 229.376 ; 
      LAYER V3 ; 
        RECT 20.304 228.62 20.376 228.716 ; 
    END 
  END dataout[45] 
  PIN wd[45] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 228.236 20.816 228.332 ; 
      LAYER M3 ; 
        RECT 19.404 227.988 19.476 229.608 ; 
      LAYER V3 ; 
        RECT 19.404 228.236 19.476 228.332 ; 
    END 
  END wd[45] 
  PIN dataout[46] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 232.94 20.544 233.036 ; 
      LAYER M3 ; 
        RECT 20.304 232.738 20.376 233.696 ; 
      LAYER V3 ; 
        RECT 20.304 232.94 20.376 233.036 ; 
    END 
  END dataout[46] 
  PIN wd[46] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 232.556 20.816 232.652 ; 
      LAYER M3 ; 
        RECT 19.404 232.308 19.476 233.928 ; 
      LAYER V3 ; 
        RECT 19.404 232.556 19.476 232.652 ; 
    END 
  END wd[46] 
  PIN dataout[47] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 237.26 20.544 237.356 ; 
      LAYER M3 ; 
        RECT 20.304 237.058 20.376 238.016 ; 
      LAYER V3 ; 
        RECT 20.304 237.26 20.376 237.356 ; 
    END 
  END dataout[47] 
  PIN wd[47] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 236.876 20.816 236.972 ; 
      LAYER M3 ; 
        RECT 19.404 236.628 19.476 238.248 ; 
      LAYER V3 ; 
        RECT 19.404 236.876 19.476 236.972 ; 
    END 
  END wd[47] 
  PIN dataout[48] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 241.58 20.544 241.676 ; 
      LAYER M3 ; 
        RECT 20.304 241.378 20.376 242.336 ; 
      LAYER V3 ; 
        RECT 20.304 241.58 20.376 241.676 ; 
    END 
  END dataout[48] 
  PIN wd[48] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 241.196 20.816 241.292 ; 
      LAYER M3 ; 
        RECT 19.404 240.948 19.476 242.568 ; 
      LAYER V3 ; 
        RECT 19.404 241.196 19.476 241.292 ; 
    END 
  END wd[48] 
  PIN dataout[49] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 245.9 20.544 245.996 ; 
      LAYER M3 ; 
        RECT 20.304 245.698 20.376 246.656 ; 
      LAYER V3 ; 
        RECT 20.304 245.9 20.376 245.996 ; 
    END 
  END dataout[49] 
  PIN wd[49] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 245.516 20.816 245.612 ; 
      LAYER M3 ; 
        RECT 19.404 245.268 19.476 246.888 ; 
      LAYER V3 ; 
        RECT 19.404 245.516 19.476 245.612 ; 
    END 
  END wd[49] 
  PIN dataout[50] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 250.22 20.544 250.316 ; 
      LAYER M3 ; 
        RECT 20.304 250.018 20.376 250.976 ; 
      LAYER V3 ; 
        RECT 20.304 250.22 20.376 250.316 ; 
    END 
  END dataout[50] 
  PIN wd[50] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 249.836 20.816 249.932 ; 
      LAYER M3 ; 
        RECT 19.404 249.588 19.476 251.208 ; 
      LAYER V3 ; 
        RECT 19.404 249.836 19.476 249.932 ; 
    END 
  END wd[50] 
  PIN dataout[51] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 254.54 20.544 254.636 ; 
      LAYER M3 ; 
        RECT 20.304 254.338 20.376 255.296 ; 
      LAYER V3 ; 
        RECT 20.304 254.54 20.376 254.636 ; 
    END 
  END dataout[51] 
  PIN wd[51] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 254.156 20.816 254.252 ; 
      LAYER M3 ; 
        RECT 19.404 253.908 19.476 255.528 ; 
      LAYER V3 ; 
        RECT 19.404 254.156 19.476 254.252 ; 
    END 
  END wd[51] 
  PIN dataout[52] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 258.86 20.544 258.956 ; 
      LAYER M3 ; 
        RECT 20.304 258.658 20.376 259.616 ; 
      LAYER V3 ; 
        RECT 20.304 258.86 20.376 258.956 ; 
    END 
  END dataout[52] 
  PIN wd[52] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 258.476 20.816 258.572 ; 
      LAYER M3 ; 
        RECT 19.404 258.228 19.476 259.848 ; 
      LAYER V3 ; 
        RECT 19.404 258.476 19.476 258.572 ; 
    END 
  END wd[52] 
  PIN dataout[53] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 263.18 20.544 263.276 ; 
      LAYER M3 ; 
        RECT 20.304 262.978 20.376 263.936 ; 
      LAYER V3 ; 
        RECT 20.304 263.18 20.376 263.276 ; 
    END 
  END dataout[53] 
  PIN wd[53] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 262.796 20.816 262.892 ; 
      LAYER M3 ; 
        RECT 19.404 262.548 19.476 264.168 ; 
      LAYER V3 ; 
        RECT 19.404 262.796 19.476 262.892 ; 
    END 
  END wd[53] 
  PIN dataout[54] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 267.5 20.544 267.596 ; 
      LAYER M3 ; 
        RECT 20.304 267.298 20.376 268.256 ; 
      LAYER V3 ; 
        RECT 20.304 267.5 20.376 267.596 ; 
    END 
  END dataout[54] 
  PIN wd[54] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 267.116 20.816 267.212 ; 
      LAYER M3 ; 
        RECT 19.404 266.868 19.476 268.488 ; 
      LAYER V3 ; 
        RECT 19.404 267.116 19.476 267.212 ; 
    END 
  END wd[54] 
  PIN dataout[55] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 271.82 20.544 271.916 ; 
      LAYER M3 ; 
        RECT 20.304 271.618 20.376 272.576 ; 
      LAYER V3 ; 
        RECT 20.304 271.82 20.376 271.916 ; 
    END 
  END dataout[55] 
  PIN wd[55] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 271.436 20.816 271.532 ; 
      LAYER M3 ; 
        RECT 19.404 271.188 19.476 272.808 ; 
      LAYER V3 ; 
        RECT 19.404 271.436 19.476 271.532 ; 
    END 
  END wd[55] 
  PIN dataout[56] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 276.14 20.544 276.236 ; 
      LAYER M3 ; 
        RECT 20.304 275.938 20.376 276.896 ; 
      LAYER V3 ; 
        RECT 20.304 276.14 20.376 276.236 ; 
    END 
  END dataout[56] 
  PIN wd[56] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 275.756 20.816 275.852 ; 
      LAYER M3 ; 
        RECT 19.404 275.508 19.476 277.128 ; 
      LAYER V3 ; 
        RECT 19.404 275.756 19.476 275.852 ; 
    END 
  END wd[56] 
  PIN dataout[57] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 280.46 20.544 280.556 ; 
      LAYER M3 ; 
        RECT 20.304 280.258 20.376 281.216 ; 
      LAYER V3 ; 
        RECT 20.304 280.46 20.376 280.556 ; 
    END 
  END dataout[57] 
  PIN wd[57] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 280.076 20.816 280.172 ; 
      LAYER M3 ; 
        RECT 19.404 279.828 19.476 281.448 ; 
      LAYER V3 ; 
        RECT 19.404 280.076 19.476 280.172 ; 
    END 
  END wd[57] 
  PIN dataout[58] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 284.78 20.544 284.876 ; 
      LAYER M3 ; 
        RECT 20.304 284.578 20.376 285.536 ; 
      LAYER V3 ; 
        RECT 20.304 284.78 20.376 284.876 ; 
    END 
  END dataout[58] 
  PIN wd[58] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 284.396 20.816 284.492 ; 
      LAYER M3 ; 
        RECT 19.404 284.148 19.476 285.768 ; 
      LAYER V3 ; 
        RECT 19.404 284.396 19.476 284.492 ; 
    END 
  END wd[58] 
  PIN dataout[59] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 289.1 20.544 289.196 ; 
      LAYER M3 ; 
        RECT 20.304 288.898 20.376 289.856 ; 
      LAYER V3 ; 
        RECT 20.304 289.1 20.376 289.196 ; 
    END 
  END dataout[59] 
  PIN wd[59] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 288.716 20.816 288.812 ; 
      LAYER M3 ; 
        RECT 19.404 288.468 19.476 290.088 ; 
      LAYER V3 ; 
        RECT 19.404 288.716 19.476 288.812 ; 
    END 
  END wd[59] 
  PIN dataout[60] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 293.42 20.544 293.516 ; 
      LAYER M3 ; 
        RECT 20.304 293.218 20.376 294.176 ; 
      LAYER V3 ; 
        RECT 20.304 293.42 20.376 293.516 ; 
    END 
  END dataout[60] 
  PIN wd[60] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 293.036 20.816 293.132 ; 
      LAYER M3 ; 
        RECT 19.404 292.788 19.476 294.408 ; 
      LAYER V3 ; 
        RECT 19.404 293.036 19.476 293.132 ; 
    END 
  END wd[60] 
  PIN dataout[61] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 297.74 20.544 297.836 ; 
      LAYER M3 ; 
        RECT 20.304 297.538 20.376 298.496 ; 
      LAYER V3 ; 
        RECT 20.304 297.74 20.376 297.836 ; 
    END 
  END dataout[61] 
  PIN wd[61] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 297.356 20.816 297.452 ; 
      LAYER M3 ; 
        RECT 19.404 297.108 19.476 298.728 ; 
      LAYER V3 ; 
        RECT 19.404 297.356 19.476 297.452 ; 
    END 
  END wd[61] 
  PIN dataout[62] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 302.06 20.544 302.156 ; 
      LAYER M3 ; 
        RECT 20.304 301.858 20.376 302.816 ; 
      LAYER V3 ; 
        RECT 20.304 302.06 20.376 302.156 ; 
    END 
  END dataout[62] 
  PIN wd[62] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 301.676 20.816 301.772 ; 
      LAYER M3 ; 
        RECT 19.404 301.428 19.476 303.048 ; 
      LAYER V3 ; 
        RECT 19.404 301.676 19.476 301.772 ; 
    END 
  END wd[62] 
  PIN dataout[63] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 306.38 20.544 306.476 ; 
      LAYER M3 ; 
        RECT 20.304 306.178 20.376 307.136 ; 
      LAYER V3 ; 
        RECT 20.304 306.38 20.376 306.476 ; 
    END 
  END dataout[63] 
  PIN wd[63] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 305.996 20.816 306.092 ; 
      LAYER M3 ; 
        RECT 19.404 305.748 19.476 307.368 ; 
      LAYER V3 ; 
        RECT 19.404 305.996 19.476 306.092 ; 
    END 
  END wd[63] 
  PIN dataout[64] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 310.7 20.544 310.796 ; 
      LAYER M3 ; 
        RECT 20.304 310.498 20.376 311.456 ; 
      LAYER V3 ; 
        RECT 20.304 310.7 20.376 310.796 ; 
    END 
  END dataout[64] 
  PIN wd[64] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 310.316 20.816 310.412 ; 
      LAYER M3 ; 
        RECT 19.404 310.068 19.476 311.688 ; 
      LAYER V3 ; 
        RECT 19.404 310.316 19.476 310.412 ; 
    END 
  END wd[64] 
  PIN dataout[65] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 315.02 20.544 315.116 ; 
      LAYER M3 ; 
        RECT 20.304 314.818 20.376 315.776 ; 
      LAYER V3 ; 
        RECT 20.304 315.02 20.376 315.116 ; 
    END 
  END dataout[65] 
  PIN wd[65] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 314.636 20.816 314.732 ; 
      LAYER M3 ; 
        RECT 19.404 314.388 19.476 316.008 ; 
      LAYER V3 ; 
        RECT 19.404 314.636 19.476 314.732 ; 
    END 
  END wd[65] 
  PIN dataout[66] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 319.34 20.544 319.436 ; 
      LAYER M3 ; 
        RECT 20.304 319.138 20.376 320.096 ; 
      LAYER V3 ; 
        RECT 20.304 319.34 20.376 319.436 ; 
    END 
  END dataout[66] 
  PIN wd[66] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 318.956 20.816 319.052 ; 
      LAYER M3 ; 
        RECT 19.404 318.708 19.476 320.328 ; 
      LAYER V3 ; 
        RECT 19.404 318.956 19.476 319.052 ; 
    END 
  END wd[66] 
  PIN dataout[67] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 323.66 20.544 323.756 ; 
      LAYER M3 ; 
        RECT 20.304 323.458 20.376 324.416 ; 
      LAYER V3 ; 
        RECT 20.304 323.66 20.376 323.756 ; 
    END 
  END dataout[67] 
  PIN wd[67] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 323.276 20.816 323.372 ; 
      LAYER M3 ; 
        RECT 19.404 323.028 19.476 324.648 ; 
      LAYER V3 ; 
        RECT 19.404 323.276 19.476 323.372 ; 
    END 
  END wd[67] 
  PIN dataout[68] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 327.98 20.544 328.076 ; 
      LAYER M3 ; 
        RECT 20.304 327.778 20.376 328.736 ; 
      LAYER V3 ; 
        RECT 20.304 327.98 20.376 328.076 ; 
    END 
  END dataout[68] 
  PIN wd[68] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 327.596 20.816 327.692 ; 
      LAYER M3 ; 
        RECT 19.404 327.348 19.476 328.968 ; 
      LAYER V3 ; 
        RECT 19.404 327.596 19.476 327.692 ; 
    END 
  END wd[68] 
  PIN dataout[69] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 332.3 20.544 332.396 ; 
      LAYER M3 ; 
        RECT 20.304 332.098 20.376 333.056 ; 
      LAYER V3 ; 
        RECT 20.304 332.3 20.376 332.396 ; 
    END 
  END dataout[69] 
  PIN wd[69] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 331.916 20.816 332.012 ; 
      LAYER M3 ; 
        RECT 19.404 331.668 19.476 333.288 ; 
      LAYER V3 ; 
        RECT 19.404 331.916 19.476 332.012 ; 
    END 
  END wd[69] 
  PIN dataout[70] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 336.62 20.544 336.716 ; 
      LAYER M3 ; 
        RECT 20.304 336.418 20.376 337.376 ; 
      LAYER V3 ; 
        RECT 20.304 336.62 20.376 336.716 ; 
    END 
  END dataout[70] 
  PIN wd[70] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 336.236 20.816 336.332 ; 
      LAYER M3 ; 
        RECT 19.404 335.988 19.476 337.608 ; 
      LAYER V3 ; 
        RECT 19.404 336.236 19.476 336.332 ; 
    END 
  END wd[70] 
  PIN dataout[71] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 340.94 20.544 341.036 ; 
      LAYER M3 ; 
        RECT 20.304 340.738 20.376 341.696 ; 
      LAYER V3 ; 
        RECT 20.304 340.94 20.376 341.036 ; 
    END 
  END dataout[71] 
  PIN wd[71] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 340.556 20.816 340.652 ; 
      LAYER M3 ; 
        RECT 19.404 340.308 19.476 341.928 ; 
      LAYER V3 ; 
        RECT 19.404 340.556 19.476 340.652 ; 
    END 
  END wd[71] 
  PIN dataout[72] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 345.26 20.544 345.356 ; 
      LAYER M3 ; 
        RECT 20.304 345.058 20.376 346.016 ; 
      LAYER V3 ; 
        RECT 20.304 345.26 20.376 345.356 ; 
    END 
  END dataout[72] 
  PIN wd[72] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 344.876 20.816 344.972 ; 
      LAYER M3 ; 
        RECT 19.404 344.628 19.476 346.248 ; 
      LAYER V3 ; 
        RECT 19.404 344.876 19.476 344.972 ; 
    END 
  END wd[72] 
  PIN dataout[73] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 349.58 20.544 349.676 ; 
      LAYER M3 ; 
        RECT 20.304 349.378 20.376 350.336 ; 
      LAYER V3 ; 
        RECT 20.304 349.58 20.376 349.676 ; 
    END 
  END dataout[73] 
  PIN wd[73] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 349.196 20.816 349.292 ; 
      LAYER M3 ; 
        RECT 19.404 348.948 19.476 350.568 ; 
      LAYER V3 ; 
        RECT 19.404 349.196 19.476 349.292 ; 
    END 
  END wd[73] 
  PIN dataout[74] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 353.9 20.544 353.996 ; 
      LAYER M3 ; 
        RECT 20.304 353.698 20.376 354.656 ; 
      LAYER V3 ; 
        RECT 20.304 353.9 20.376 353.996 ; 
    END 
  END dataout[74] 
  PIN wd[74] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 353.516 20.816 353.612 ; 
      LAYER M3 ; 
        RECT 19.404 353.268 19.476 354.888 ; 
      LAYER V3 ; 
        RECT 19.404 353.516 19.476 353.612 ; 
    END 
  END wd[74] 
  PIN dataout[75] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 358.22 20.544 358.316 ; 
      LAYER M3 ; 
        RECT 20.304 358.018 20.376 358.976 ; 
      LAYER V3 ; 
        RECT 20.304 358.22 20.376 358.316 ; 
    END 
  END dataout[75] 
  PIN wd[75] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 357.836 20.816 357.932 ; 
      LAYER M3 ; 
        RECT 19.404 357.588 19.476 359.208 ; 
      LAYER V3 ; 
        RECT 19.404 357.836 19.476 357.932 ; 
    END 
  END wd[75] 
  PIN dataout[76] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 362.54 20.544 362.636 ; 
      LAYER M3 ; 
        RECT 20.304 362.338 20.376 363.296 ; 
      LAYER V3 ; 
        RECT 20.304 362.54 20.376 362.636 ; 
    END 
  END dataout[76] 
  PIN wd[76] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 362.156 20.816 362.252 ; 
      LAYER M3 ; 
        RECT 19.404 361.908 19.476 363.528 ; 
      LAYER V3 ; 
        RECT 19.404 362.156 19.476 362.252 ; 
    END 
  END wd[76] 
  PIN dataout[77] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 366.86 20.544 366.956 ; 
      LAYER M3 ; 
        RECT 20.304 366.658 20.376 367.616 ; 
      LAYER V3 ; 
        RECT 20.304 366.86 20.376 366.956 ; 
    END 
  END dataout[77] 
  PIN wd[77] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 366.476 20.816 366.572 ; 
      LAYER M3 ; 
        RECT 19.404 366.228 19.476 367.848 ; 
      LAYER V3 ; 
        RECT 19.404 366.476 19.476 366.572 ; 
    END 
  END wd[77] 
  PIN dataout[78] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 371.18 20.544 371.276 ; 
      LAYER M3 ; 
        RECT 20.304 370.978 20.376 371.936 ; 
      LAYER V3 ; 
        RECT 20.304 371.18 20.376 371.276 ; 
    END 
  END dataout[78] 
  PIN wd[78] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 370.796 20.816 370.892 ; 
      LAYER M3 ; 
        RECT 19.404 370.548 19.476 372.168 ; 
      LAYER V3 ; 
        RECT 19.404 370.796 19.476 370.892 ; 
    END 
  END wd[78] 
  PIN dataout[79] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 375.5 20.544 375.596 ; 
      LAYER M3 ; 
        RECT 20.304 375.298 20.376 376.256 ; 
      LAYER V3 ; 
        RECT 20.304 375.5 20.376 375.596 ; 
    END 
  END dataout[79] 
  PIN wd[79] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 375.116 20.816 375.212 ; 
      LAYER M3 ; 
        RECT 19.404 374.868 19.476 376.488 ; 
      LAYER V3 ; 
        RECT 19.404 375.116 19.476 375.212 ; 
    END 
  END wd[79] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.706 38.448 109.08 ; 
      RECT 0 109.026 38.448 113.4 ; 
      RECT 0 113.346 38.448 117.72 ; 
      RECT 0 117.666 38.448 122.04 ; 
      RECT 0 121.986 38.448 126.36 ; 
      RECT 0 126.306 38.448 130.68 ; 
      RECT 0 130.626 38.448 135 ; 
      RECT 0 134.946 38.448 139.32 ; 
      RECT 0 139.266 38.448 143.64 ; 
      RECT 0 143.586 38.448 147.96 ; 
      RECT 0 147.906 38.448 152.28 ; 
      RECT 0 152.226 38.448 156.6 ; 
      RECT 0 156.546 38.448 160.92 ; 
      RECT 0 160.866 38.448 165.24 ; 
      RECT 0 165.186 38.448 169.56 ; 
      RECT 0 169.506 38.448 173.88 ; 
      RECT 0 173.772 38.448 208.386 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
        RECT 0 240.894 38.448 245.268 ; 
        RECT 0 245.214 38.448 249.588 ; 
        RECT 0 249.534 38.448 253.908 ; 
        RECT 0 253.854 38.448 258.228 ; 
        RECT 0 258.174 38.448 262.548 ; 
        RECT 0 262.494 38.448 266.868 ; 
        RECT 0 266.814 38.448 271.188 ; 
        RECT 0 271.134 38.448 275.508 ; 
        RECT 0 275.454 38.448 279.828 ; 
        RECT 0 279.774 38.448 284.148 ; 
        RECT 0 284.094 38.448 288.468 ; 
        RECT 0 288.414 38.448 292.788 ; 
        RECT 0 292.734 38.448 297.108 ; 
        RECT 0 297.054 38.448 301.428 ; 
        RECT 0 301.374 38.448 305.748 ; 
        RECT 0 305.694 38.448 310.068 ; 
        RECT 0 310.014 38.448 314.388 ; 
        RECT 0 314.334 38.448 318.708 ; 
        RECT 0 318.654 38.448 323.028 ; 
        RECT 0 322.974 38.448 327.348 ; 
        RECT 0 327.294 38.448 331.668 ; 
        RECT 0 331.614 38.448 335.988 ; 
        RECT 0 335.934 38.448 340.308 ; 
        RECT 0 340.254 38.448 344.628 ; 
        RECT 0 344.574 38.448 348.948 ; 
        RECT 0 348.894 38.448 353.268 ; 
        RECT 0 353.214 38.448 357.588 ; 
        RECT 0 357.534 38.448 361.908 ; 
        RECT 0 361.854 38.448 366.228 ; 
        RECT 0 366.174 38.448 370.548 ; 
        RECT 0 370.494 38.448 374.868 ; 
        RECT 0 374.814 38.448 379.188 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.706 38.448 109.08 ; 
      RECT 0 109.026 38.448 113.4 ; 
      RECT 0 113.346 38.448 117.72 ; 
      RECT 0 117.666 38.448 122.04 ; 
      RECT 0 121.986 38.448 126.36 ; 
      RECT 0 126.306 38.448 130.68 ; 
      RECT 0 130.626 38.448 135 ; 
      RECT 0 134.946 38.448 139.32 ; 
      RECT 0 139.266 38.448 143.64 ; 
      RECT 0 143.586 38.448 147.96 ; 
      RECT 0 147.906 38.448 152.28 ; 
      RECT 0 152.226 38.448 156.6 ; 
      RECT 0 156.546 38.448 160.92 ; 
      RECT 0 160.866 38.448 165.24 ; 
      RECT 0 165.186 38.448 169.56 ; 
      RECT 0 169.506 38.448 173.88 ; 
      RECT 0 173.772 38.448 208.386 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
        RECT 0 240.894 38.448 245.268 ; 
        RECT 0 245.214 38.448 249.588 ; 
        RECT 0 249.534 38.448 253.908 ; 
        RECT 0 253.854 38.448 258.228 ; 
        RECT 0 258.174 38.448 262.548 ; 
        RECT 0 262.494 38.448 266.868 ; 
        RECT 0 266.814 38.448 271.188 ; 
        RECT 0 271.134 38.448 275.508 ; 
        RECT 0 275.454 38.448 279.828 ; 
        RECT 0 279.774 38.448 284.148 ; 
        RECT 0 284.094 38.448 288.468 ; 
        RECT 0 288.414 38.448 292.788 ; 
        RECT 0 292.734 38.448 297.108 ; 
        RECT 0 297.054 38.448 301.428 ; 
        RECT 0 301.374 38.448 305.748 ; 
        RECT 0 305.694 38.448 310.068 ; 
        RECT 0 310.014 38.448 314.388 ; 
        RECT 0 314.334 38.448 318.708 ; 
        RECT 0 318.654 38.448 323.028 ; 
        RECT 0 322.974 38.448 327.348 ; 
        RECT 0 327.294 38.448 331.668 ; 
        RECT 0 331.614 38.448 335.988 ; 
        RECT 0 335.934 38.448 340.308 ; 
        RECT 0 340.254 38.448 344.628 ; 
        RECT 0 344.574 38.448 348.948 ; 
        RECT 0 348.894 38.448 353.268 ; 
        RECT 0 353.214 38.448 357.588 ; 
        RECT 0 357.534 38.448 361.908 ; 
        RECT 0 361.854 38.448 366.228 ; 
        RECT 0 366.174 38.448 370.548 ; 
        RECT 0 370.494 38.448 374.868 ; 
        RECT 0 374.814 38.448 379.188 ; 
  LAYER V1 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.706 38.448 109.08 ; 
      RECT 0 109.026 38.448 113.4 ; 
      RECT 0 113.346 38.448 117.72 ; 
      RECT 0 117.666 38.448 122.04 ; 
      RECT 0 121.986 38.448 126.36 ; 
      RECT 0 126.306 38.448 130.68 ; 
      RECT 0 130.626 38.448 135 ; 
      RECT 0 134.946 38.448 139.32 ; 
      RECT 0 139.266 38.448 143.64 ; 
      RECT 0 143.586 38.448 147.96 ; 
      RECT 0 147.906 38.448 152.28 ; 
      RECT 0 152.226 38.448 156.6 ; 
      RECT 0 156.546 38.448 160.92 ; 
      RECT 0 160.866 38.448 165.24 ; 
      RECT 0 165.186 38.448 169.56 ; 
      RECT 0 169.506 38.448 173.88 ; 
      RECT 0 173.772 38.448 208.386 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
        RECT 0 240.894 38.448 245.268 ; 
        RECT 0 245.214 38.448 249.588 ; 
        RECT 0 249.534 38.448 253.908 ; 
        RECT 0 253.854 38.448 258.228 ; 
        RECT 0 258.174 38.448 262.548 ; 
        RECT 0 262.494 38.448 266.868 ; 
        RECT 0 266.814 38.448 271.188 ; 
        RECT 0 271.134 38.448 275.508 ; 
        RECT 0 275.454 38.448 279.828 ; 
        RECT 0 279.774 38.448 284.148 ; 
        RECT 0 284.094 38.448 288.468 ; 
        RECT 0 288.414 38.448 292.788 ; 
        RECT 0 292.734 38.448 297.108 ; 
        RECT 0 297.054 38.448 301.428 ; 
        RECT 0 301.374 38.448 305.748 ; 
        RECT 0 305.694 38.448 310.068 ; 
        RECT 0 310.014 38.448 314.388 ; 
        RECT 0 314.334 38.448 318.708 ; 
        RECT 0 318.654 38.448 323.028 ; 
        RECT 0 322.974 38.448 327.348 ; 
        RECT 0 327.294 38.448 331.668 ; 
        RECT 0 331.614 38.448 335.988 ; 
        RECT 0 335.934 38.448 340.308 ; 
        RECT 0 340.254 38.448 344.628 ; 
        RECT 0 344.574 38.448 348.948 ; 
        RECT 0 348.894 38.448 353.268 ; 
        RECT 0 353.214 38.448 357.588 ; 
        RECT 0 357.534 38.448 361.908 ; 
        RECT 0 361.854 38.448 366.228 ; 
        RECT 0 366.174 38.448 370.548 ; 
        RECT 0 370.494 38.448 374.868 ; 
        RECT 0 374.814 38.448 379.188 ; 
  LAYER V2 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.466 38.448 78.84 ; 
      RECT 0 78.786 38.448 83.16 ; 
      RECT 0 83.106 38.448 87.48 ; 
      RECT 0 87.426 38.448 91.8 ; 
      RECT 0 91.746 38.448 96.12 ; 
      RECT 0 96.066 38.448 100.44 ; 
      RECT 0 100.386 38.448 104.76 ; 
      RECT 0 104.706 38.448 109.08 ; 
      RECT 0 109.026 38.448 113.4 ; 
      RECT 0 113.346 38.448 117.72 ; 
      RECT 0 117.666 38.448 122.04 ; 
      RECT 0 121.986 38.448 126.36 ; 
      RECT 0 126.306 38.448 130.68 ; 
      RECT 0 130.626 38.448 135 ; 
      RECT 0 134.946 38.448 139.32 ; 
      RECT 0 139.266 38.448 143.64 ; 
      RECT 0 143.586 38.448 147.96 ; 
      RECT 0 147.906 38.448 152.28 ; 
      RECT 0 152.226 38.448 156.6 ; 
      RECT 0 156.546 38.448 160.92 ; 
      RECT 0 160.866 38.448 165.24 ; 
      RECT 0 165.186 38.448 169.56 ; 
      RECT 0 169.506 38.448 173.88 ; 
      RECT 0 173.772 38.448 208.386 ; 
        RECT 0 206.334 38.448 210.708 ; 
        RECT 0 210.654 38.448 215.028 ; 
        RECT 0 214.974 38.448 219.348 ; 
        RECT 0 219.294 38.448 223.668 ; 
        RECT 0 223.614 38.448 227.988 ; 
        RECT 0 227.934 38.448 232.308 ; 
        RECT 0 232.254 38.448 236.628 ; 
        RECT 0 236.574 38.448 240.948 ; 
        RECT 0 240.894 38.448 245.268 ; 
        RECT 0 245.214 38.448 249.588 ; 
        RECT 0 249.534 38.448 253.908 ; 
        RECT 0 253.854 38.448 258.228 ; 
        RECT 0 258.174 38.448 262.548 ; 
        RECT 0 262.494 38.448 266.868 ; 
        RECT 0 266.814 38.448 271.188 ; 
        RECT 0 271.134 38.448 275.508 ; 
        RECT 0 275.454 38.448 279.828 ; 
        RECT 0 279.774 38.448 284.148 ; 
        RECT 0 284.094 38.448 288.468 ; 
        RECT 0 288.414 38.448 292.788 ; 
        RECT 0 292.734 38.448 297.108 ; 
        RECT 0 297.054 38.448 301.428 ; 
        RECT 0 301.374 38.448 305.748 ; 
        RECT 0 305.694 38.448 310.068 ; 
        RECT 0 310.014 38.448 314.388 ; 
        RECT 0 314.334 38.448 318.708 ; 
        RECT 0 318.654 38.448 323.028 ; 
        RECT 0 322.974 38.448 327.348 ; 
        RECT 0 327.294 38.448 331.668 ; 
        RECT 0 331.614 38.448 335.988 ; 
        RECT 0 335.934 38.448 340.308 ; 
        RECT 0 340.254 38.448 344.628 ; 
        RECT 0 344.574 38.448 348.948 ; 
        RECT 0 348.894 38.448 353.268 ; 
        RECT 0 353.214 38.448 357.588 ; 
        RECT 0 357.534 38.448 361.908 ; 
        RECT 0 361.854 38.448 366.228 ; 
        RECT 0 366.174 38.448 370.548 ; 
        RECT 0 370.494 38.448 374.868 ; 
        RECT 0 374.814 38.448 379.188 ; 
  LAYER M3 ; 
      RECT 20.952 1.38 21.024 5.122 ; 
      RECT 20.808 1.38 20.88 5.122 ; 
      RECT 20.664 3.688 20.736 4.978 ; 
      RECT 20.196 4.476 20.268 4.914 ; 
      RECT 20.16 1.51 20.232 2.468 ; 
      RECT 20.016 3.834 20.088 4.448 ; 
      RECT 19.692 3.936 19.764 4.968 ; 
      RECT 17.532 1.38 17.604 5.122 ; 
      RECT 17.388 1.38 17.46 5.122 ; 
      RECT 17.244 2.104 17.316 4.376 ; 
      RECT 20.952 5.7 21.024 9.442 ; 
      RECT 20.808 5.7 20.88 9.442 ; 
      RECT 20.664 8.008 20.736 9.298 ; 
      RECT 20.196 8.796 20.268 9.234 ; 
      RECT 20.16 5.83 20.232 6.788 ; 
      RECT 20.016 8.154 20.088 8.768 ; 
      RECT 19.692 8.256 19.764 9.288 ; 
      RECT 17.532 5.7 17.604 9.442 ; 
      RECT 17.388 5.7 17.46 9.442 ; 
      RECT 17.244 6.424 17.316 8.696 ; 
      RECT 20.952 10.02 21.024 13.762 ; 
      RECT 20.808 10.02 20.88 13.762 ; 
      RECT 20.664 12.328 20.736 13.618 ; 
      RECT 20.196 13.116 20.268 13.554 ; 
      RECT 20.16 10.15 20.232 11.108 ; 
      RECT 20.016 12.474 20.088 13.088 ; 
      RECT 19.692 12.576 19.764 13.608 ; 
      RECT 17.532 10.02 17.604 13.762 ; 
      RECT 17.388 10.02 17.46 13.762 ; 
      RECT 17.244 10.744 17.316 13.016 ; 
      RECT 20.952 14.34 21.024 18.082 ; 
      RECT 20.808 14.34 20.88 18.082 ; 
      RECT 20.664 16.648 20.736 17.938 ; 
      RECT 20.196 17.436 20.268 17.874 ; 
      RECT 20.16 14.47 20.232 15.428 ; 
      RECT 20.016 16.794 20.088 17.408 ; 
      RECT 19.692 16.896 19.764 17.928 ; 
      RECT 17.532 14.34 17.604 18.082 ; 
      RECT 17.388 14.34 17.46 18.082 ; 
      RECT 17.244 15.064 17.316 17.336 ; 
      RECT 20.952 18.66 21.024 22.402 ; 
      RECT 20.808 18.66 20.88 22.402 ; 
      RECT 20.664 20.968 20.736 22.258 ; 
      RECT 20.196 21.756 20.268 22.194 ; 
      RECT 20.16 18.79 20.232 19.748 ; 
      RECT 20.016 21.114 20.088 21.728 ; 
      RECT 19.692 21.216 19.764 22.248 ; 
      RECT 17.532 18.66 17.604 22.402 ; 
      RECT 17.388 18.66 17.46 22.402 ; 
      RECT 17.244 19.384 17.316 21.656 ; 
      RECT 20.952 22.98 21.024 26.722 ; 
      RECT 20.808 22.98 20.88 26.722 ; 
      RECT 20.664 25.288 20.736 26.578 ; 
      RECT 20.196 26.076 20.268 26.514 ; 
      RECT 20.16 23.11 20.232 24.068 ; 
      RECT 20.016 25.434 20.088 26.048 ; 
      RECT 19.692 25.536 19.764 26.568 ; 
      RECT 17.532 22.98 17.604 26.722 ; 
      RECT 17.388 22.98 17.46 26.722 ; 
      RECT 17.244 23.704 17.316 25.976 ; 
      RECT 20.952 27.3 21.024 31.042 ; 
      RECT 20.808 27.3 20.88 31.042 ; 
      RECT 20.664 29.608 20.736 30.898 ; 
      RECT 20.196 30.396 20.268 30.834 ; 
      RECT 20.16 27.43 20.232 28.388 ; 
      RECT 20.016 29.754 20.088 30.368 ; 
      RECT 19.692 29.856 19.764 30.888 ; 
      RECT 17.532 27.3 17.604 31.042 ; 
      RECT 17.388 27.3 17.46 31.042 ; 
      RECT 17.244 28.024 17.316 30.296 ; 
      RECT 20.952 31.62 21.024 35.362 ; 
      RECT 20.808 31.62 20.88 35.362 ; 
      RECT 20.664 33.928 20.736 35.218 ; 
      RECT 20.196 34.716 20.268 35.154 ; 
      RECT 20.16 31.75 20.232 32.708 ; 
      RECT 20.016 34.074 20.088 34.688 ; 
      RECT 19.692 34.176 19.764 35.208 ; 
      RECT 17.532 31.62 17.604 35.362 ; 
      RECT 17.388 31.62 17.46 35.362 ; 
      RECT 17.244 32.344 17.316 34.616 ; 
      RECT 20.952 35.94 21.024 39.682 ; 
      RECT 20.808 35.94 20.88 39.682 ; 
      RECT 20.664 38.248 20.736 39.538 ; 
      RECT 20.196 39.036 20.268 39.474 ; 
      RECT 20.16 36.07 20.232 37.028 ; 
      RECT 20.016 38.394 20.088 39.008 ; 
      RECT 19.692 38.496 19.764 39.528 ; 
      RECT 17.532 35.94 17.604 39.682 ; 
      RECT 17.388 35.94 17.46 39.682 ; 
      RECT 17.244 36.664 17.316 38.936 ; 
      RECT 20.952 40.26 21.024 44.002 ; 
      RECT 20.808 40.26 20.88 44.002 ; 
      RECT 20.664 42.568 20.736 43.858 ; 
      RECT 20.196 43.356 20.268 43.794 ; 
      RECT 20.16 40.39 20.232 41.348 ; 
      RECT 20.016 42.714 20.088 43.328 ; 
      RECT 19.692 42.816 19.764 43.848 ; 
      RECT 17.532 40.26 17.604 44.002 ; 
      RECT 17.388 40.26 17.46 44.002 ; 
      RECT 17.244 40.984 17.316 43.256 ; 
      RECT 20.952 44.58 21.024 48.322 ; 
      RECT 20.808 44.58 20.88 48.322 ; 
      RECT 20.664 46.888 20.736 48.178 ; 
      RECT 20.196 47.676 20.268 48.114 ; 
      RECT 20.16 44.71 20.232 45.668 ; 
      RECT 20.016 47.034 20.088 47.648 ; 
      RECT 19.692 47.136 19.764 48.168 ; 
      RECT 17.532 44.58 17.604 48.322 ; 
      RECT 17.388 44.58 17.46 48.322 ; 
      RECT 17.244 45.304 17.316 47.576 ; 
      RECT 20.952 48.9 21.024 52.642 ; 
      RECT 20.808 48.9 20.88 52.642 ; 
      RECT 20.664 51.208 20.736 52.498 ; 
      RECT 20.196 51.996 20.268 52.434 ; 
      RECT 20.16 49.03 20.232 49.988 ; 
      RECT 20.016 51.354 20.088 51.968 ; 
      RECT 19.692 51.456 19.764 52.488 ; 
      RECT 17.532 48.9 17.604 52.642 ; 
      RECT 17.388 48.9 17.46 52.642 ; 
      RECT 17.244 49.624 17.316 51.896 ; 
      RECT 20.952 53.22 21.024 56.962 ; 
      RECT 20.808 53.22 20.88 56.962 ; 
      RECT 20.664 55.528 20.736 56.818 ; 
      RECT 20.196 56.316 20.268 56.754 ; 
      RECT 20.16 53.35 20.232 54.308 ; 
      RECT 20.016 55.674 20.088 56.288 ; 
      RECT 19.692 55.776 19.764 56.808 ; 
      RECT 17.532 53.22 17.604 56.962 ; 
      RECT 17.388 53.22 17.46 56.962 ; 
      RECT 17.244 53.944 17.316 56.216 ; 
      RECT 20.952 57.54 21.024 61.282 ; 
      RECT 20.808 57.54 20.88 61.282 ; 
      RECT 20.664 59.848 20.736 61.138 ; 
      RECT 20.196 60.636 20.268 61.074 ; 
      RECT 20.16 57.67 20.232 58.628 ; 
      RECT 20.016 59.994 20.088 60.608 ; 
      RECT 19.692 60.096 19.764 61.128 ; 
      RECT 17.532 57.54 17.604 61.282 ; 
      RECT 17.388 57.54 17.46 61.282 ; 
      RECT 17.244 58.264 17.316 60.536 ; 
      RECT 20.952 61.86 21.024 65.602 ; 
      RECT 20.808 61.86 20.88 65.602 ; 
      RECT 20.664 64.168 20.736 65.458 ; 
      RECT 20.196 64.956 20.268 65.394 ; 
      RECT 20.16 61.99 20.232 62.948 ; 
      RECT 20.016 64.314 20.088 64.928 ; 
      RECT 19.692 64.416 19.764 65.448 ; 
      RECT 17.532 61.86 17.604 65.602 ; 
      RECT 17.388 61.86 17.46 65.602 ; 
      RECT 17.244 62.584 17.316 64.856 ; 
      RECT 20.952 66.18 21.024 69.922 ; 
      RECT 20.808 66.18 20.88 69.922 ; 
      RECT 20.664 68.488 20.736 69.778 ; 
      RECT 20.196 69.276 20.268 69.714 ; 
      RECT 20.16 66.31 20.232 67.268 ; 
      RECT 20.016 68.634 20.088 69.248 ; 
      RECT 19.692 68.736 19.764 69.768 ; 
      RECT 17.532 66.18 17.604 69.922 ; 
      RECT 17.388 66.18 17.46 69.922 ; 
      RECT 17.244 66.904 17.316 69.176 ; 
      RECT 20.952 70.5 21.024 74.242 ; 
      RECT 20.808 70.5 20.88 74.242 ; 
      RECT 20.664 72.808 20.736 74.098 ; 
      RECT 20.196 73.596 20.268 74.034 ; 
      RECT 20.16 70.63 20.232 71.588 ; 
      RECT 20.016 72.954 20.088 73.568 ; 
      RECT 19.692 73.056 19.764 74.088 ; 
      RECT 17.532 70.5 17.604 74.242 ; 
      RECT 17.388 70.5 17.46 74.242 ; 
      RECT 17.244 71.224 17.316 73.496 ; 
      RECT 20.952 74.82 21.024 78.562 ; 
      RECT 20.808 74.82 20.88 78.562 ; 
      RECT 20.664 77.128 20.736 78.418 ; 
      RECT 20.196 77.916 20.268 78.354 ; 
      RECT 20.16 74.95 20.232 75.908 ; 
      RECT 20.016 77.274 20.088 77.888 ; 
      RECT 19.692 77.376 19.764 78.408 ; 
      RECT 17.532 74.82 17.604 78.562 ; 
      RECT 17.388 74.82 17.46 78.562 ; 
      RECT 17.244 75.544 17.316 77.816 ; 
      RECT 20.952 79.14 21.024 82.882 ; 
      RECT 20.808 79.14 20.88 82.882 ; 
      RECT 20.664 81.448 20.736 82.738 ; 
      RECT 20.196 82.236 20.268 82.674 ; 
      RECT 20.16 79.27 20.232 80.228 ; 
      RECT 20.016 81.594 20.088 82.208 ; 
      RECT 19.692 81.696 19.764 82.728 ; 
      RECT 17.532 79.14 17.604 82.882 ; 
      RECT 17.388 79.14 17.46 82.882 ; 
      RECT 17.244 79.864 17.316 82.136 ; 
      RECT 20.952 83.46 21.024 87.202 ; 
      RECT 20.808 83.46 20.88 87.202 ; 
      RECT 20.664 85.768 20.736 87.058 ; 
      RECT 20.196 86.556 20.268 86.994 ; 
      RECT 20.16 83.59 20.232 84.548 ; 
      RECT 20.016 85.914 20.088 86.528 ; 
      RECT 19.692 86.016 19.764 87.048 ; 
      RECT 17.532 83.46 17.604 87.202 ; 
      RECT 17.388 83.46 17.46 87.202 ; 
      RECT 17.244 84.184 17.316 86.456 ; 
      RECT 20.952 87.78 21.024 91.522 ; 
      RECT 20.808 87.78 20.88 91.522 ; 
      RECT 20.664 90.088 20.736 91.378 ; 
      RECT 20.196 90.876 20.268 91.314 ; 
      RECT 20.16 87.91 20.232 88.868 ; 
      RECT 20.016 90.234 20.088 90.848 ; 
      RECT 19.692 90.336 19.764 91.368 ; 
      RECT 17.532 87.78 17.604 91.522 ; 
      RECT 17.388 87.78 17.46 91.522 ; 
      RECT 17.244 88.504 17.316 90.776 ; 
      RECT 20.952 92.1 21.024 95.842 ; 
      RECT 20.808 92.1 20.88 95.842 ; 
      RECT 20.664 94.408 20.736 95.698 ; 
      RECT 20.196 95.196 20.268 95.634 ; 
      RECT 20.16 92.23 20.232 93.188 ; 
      RECT 20.016 94.554 20.088 95.168 ; 
      RECT 19.692 94.656 19.764 95.688 ; 
      RECT 17.532 92.1 17.604 95.842 ; 
      RECT 17.388 92.1 17.46 95.842 ; 
      RECT 17.244 92.824 17.316 95.096 ; 
      RECT 20.952 96.42 21.024 100.162 ; 
      RECT 20.808 96.42 20.88 100.162 ; 
      RECT 20.664 98.728 20.736 100.018 ; 
      RECT 20.196 99.516 20.268 99.954 ; 
      RECT 20.16 96.55 20.232 97.508 ; 
      RECT 20.016 98.874 20.088 99.488 ; 
      RECT 19.692 98.976 19.764 100.008 ; 
      RECT 17.532 96.42 17.604 100.162 ; 
      RECT 17.388 96.42 17.46 100.162 ; 
      RECT 17.244 97.144 17.316 99.416 ; 
      RECT 20.952 100.74 21.024 104.482 ; 
      RECT 20.808 100.74 20.88 104.482 ; 
      RECT 20.664 103.048 20.736 104.338 ; 
      RECT 20.196 103.836 20.268 104.274 ; 
      RECT 20.16 100.87 20.232 101.828 ; 
      RECT 20.016 103.194 20.088 103.808 ; 
      RECT 19.692 103.296 19.764 104.328 ; 
      RECT 17.532 100.74 17.604 104.482 ; 
      RECT 17.388 100.74 17.46 104.482 ; 
      RECT 17.244 101.464 17.316 103.736 ; 
      RECT 20.952 105.06 21.024 108.802 ; 
      RECT 20.808 105.06 20.88 108.802 ; 
      RECT 20.664 107.368 20.736 108.658 ; 
      RECT 20.196 108.156 20.268 108.594 ; 
      RECT 20.16 105.19 20.232 106.148 ; 
      RECT 20.016 107.514 20.088 108.128 ; 
      RECT 19.692 107.616 19.764 108.648 ; 
      RECT 17.532 105.06 17.604 108.802 ; 
      RECT 17.388 105.06 17.46 108.802 ; 
      RECT 17.244 105.784 17.316 108.056 ; 
      RECT 20.952 109.38 21.024 113.122 ; 
      RECT 20.808 109.38 20.88 113.122 ; 
      RECT 20.664 111.688 20.736 112.978 ; 
      RECT 20.196 112.476 20.268 112.914 ; 
      RECT 20.16 109.51 20.232 110.468 ; 
      RECT 20.016 111.834 20.088 112.448 ; 
      RECT 19.692 111.936 19.764 112.968 ; 
      RECT 17.532 109.38 17.604 113.122 ; 
      RECT 17.388 109.38 17.46 113.122 ; 
      RECT 17.244 110.104 17.316 112.376 ; 
      RECT 20.952 113.7 21.024 117.442 ; 
      RECT 20.808 113.7 20.88 117.442 ; 
      RECT 20.664 116.008 20.736 117.298 ; 
      RECT 20.196 116.796 20.268 117.234 ; 
      RECT 20.16 113.83 20.232 114.788 ; 
      RECT 20.016 116.154 20.088 116.768 ; 
      RECT 19.692 116.256 19.764 117.288 ; 
      RECT 17.532 113.7 17.604 117.442 ; 
      RECT 17.388 113.7 17.46 117.442 ; 
      RECT 17.244 114.424 17.316 116.696 ; 
      RECT 20.952 118.02 21.024 121.762 ; 
      RECT 20.808 118.02 20.88 121.762 ; 
      RECT 20.664 120.328 20.736 121.618 ; 
      RECT 20.196 121.116 20.268 121.554 ; 
      RECT 20.16 118.15 20.232 119.108 ; 
      RECT 20.016 120.474 20.088 121.088 ; 
      RECT 19.692 120.576 19.764 121.608 ; 
      RECT 17.532 118.02 17.604 121.762 ; 
      RECT 17.388 118.02 17.46 121.762 ; 
      RECT 17.244 118.744 17.316 121.016 ; 
      RECT 20.952 122.34 21.024 126.082 ; 
      RECT 20.808 122.34 20.88 126.082 ; 
      RECT 20.664 124.648 20.736 125.938 ; 
      RECT 20.196 125.436 20.268 125.874 ; 
      RECT 20.16 122.47 20.232 123.428 ; 
      RECT 20.016 124.794 20.088 125.408 ; 
      RECT 19.692 124.896 19.764 125.928 ; 
      RECT 17.532 122.34 17.604 126.082 ; 
      RECT 17.388 122.34 17.46 126.082 ; 
      RECT 17.244 123.064 17.316 125.336 ; 
      RECT 20.952 126.66 21.024 130.402 ; 
      RECT 20.808 126.66 20.88 130.402 ; 
      RECT 20.664 128.968 20.736 130.258 ; 
      RECT 20.196 129.756 20.268 130.194 ; 
      RECT 20.16 126.79 20.232 127.748 ; 
      RECT 20.016 129.114 20.088 129.728 ; 
      RECT 19.692 129.216 19.764 130.248 ; 
      RECT 17.532 126.66 17.604 130.402 ; 
      RECT 17.388 126.66 17.46 130.402 ; 
      RECT 17.244 127.384 17.316 129.656 ; 
      RECT 20.952 130.98 21.024 134.722 ; 
      RECT 20.808 130.98 20.88 134.722 ; 
      RECT 20.664 133.288 20.736 134.578 ; 
      RECT 20.196 134.076 20.268 134.514 ; 
      RECT 20.16 131.11 20.232 132.068 ; 
      RECT 20.016 133.434 20.088 134.048 ; 
      RECT 19.692 133.536 19.764 134.568 ; 
      RECT 17.532 130.98 17.604 134.722 ; 
      RECT 17.388 130.98 17.46 134.722 ; 
      RECT 17.244 131.704 17.316 133.976 ; 
      RECT 20.952 135.3 21.024 139.042 ; 
      RECT 20.808 135.3 20.88 139.042 ; 
      RECT 20.664 137.608 20.736 138.898 ; 
      RECT 20.196 138.396 20.268 138.834 ; 
      RECT 20.16 135.43 20.232 136.388 ; 
      RECT 20.016 137.754 20.088 138.368 ; 
      RECT 19.692 137.856 19.764 138.888 ; 
      RECT 17.532 135.3 17.604 139.042 ; 
      RECT 17.388 135.3 17.46 139.042 ; 
      RECT 17.244 136.024 17.316 138.296 ; 
      RECT 20.952 139.62 21.024 143.362 ; 
      RECT 20.808 139.62 20.88 143.362 ; 
      RECT 20.664 141.928 20.736 143.218 ; 
      RECT 20.196 142.716 20.268 143.154 ; 
      RECT 20.16 139.75 20.232 140.708 ; 
      RECT 20.016 142.074 20.088 142.688 ; 
      RECT 19.692 142.176 19.764 143.208 ; 
      RECT 17.532 139.62 17.604 143.362 ; 
      RECT 17.388 139.62 17.46 143.362 ; 
      RECT 17.244 140.344 17.316 142.616 ; 
      RECT 20.952 143.94 21.024 147.682 ; 
      RECT 20.808 143.94 20.88 147.682 ; 
      RECT 20.664 146.248 20.736 147.538 ; 
      RECT 20.196 147.036 20.268 147.474 ; 
      RECT 20.16 144.07 20.232 145.028 ; 
      RECT 20.016 146.394 20.088 147.008 ; 
      RECT 19.692 146.496 19.764 147.528 ; 
      RECT 17.532 143.94 17.604 147.682 ; 
      RECT 17.388 143.94 17.46 147.682 ; 
      RECT 17.244 144.664 17.316 146.936 ; 
      RECT 20.952 148.26 21.024 152.002 ; 
      RECT 20.808 148.26 20.88 152.002 ; 
      RECT 20.664 150.568 20.736 151.858 ; 
      RECT 20.196 151.356 20.268 151.794 ; 
      RECT 20.16 148.39 20.232 149.348 ; 
      RECT 20.016 150.714 20.088 151.328 ; 
      RECT 19.692 150.816 19.764 151.848 ; 
      RECT 17.532 148.26 17.604 152.002 ; 
      RECT 17.388 148.26 17.46 152.002 ; 
      RECT 17.244 148.984 17.316 151.256 ; 
      RECT 20.952 152.58 21.024 156.322 ; 
      RECT 20.808 152.58 20.88 156.322 ; 
      RECT 20.664 154.888 20.736 156.178 ; 
      RECT 20.196 155.676 20.268 156.114 ; 
      RECT 20.16 152.71 20.232 153.668 ; 
      RECT 20.016 155.034 20.088 155.648 ; 
      RECT 19.692 155.136 19.764 156.168 ; 
      RECT 17.532 152.58 17.604 156.322 ; 
      RECT 17.388 152.58 17.46 156.322 ; 
      RECT 17.244 153.304 17.316 155.576 ; 
      RECT 20.952 156.9 21.024 160.642 ; 
      RECT 20.808 156.9 20.88 160.642 ; 
      RECT 20.664 159.208 20.736 160.498 ; 
      RECT 20.196 159.996 20.268 160.434 ; 
      RECT 20.16 157.03 20.232 157.988 ; 
      RECT 20.016 159.354 20.088 159.968 ; 
      RECT 19.692 159.456 19.764 160.488 ; 
      RECT 17.532 156.9 17.604 160.642 ; 
      RECT 17.388 156.9 17.46 160.642 ; 
      RECT 17.244 157.624 17.316 159.896 ; 
      RECT 20.952 161.22 21.024 164.962 ; 
      RECT 20.808 161.22 20.88 164.962 ; 
      RECT 20.664 163.528 20.736 164.818 ; 
      RECT 20.196 164.316 20.268 164.754 ; 
      RECT 20.16 161.35 20.232 162.308 ; 
      RECT 20.016 163.674 20.088 164.288 ; 
      RECT 19.692 163.776 19.764 164.808 ; 
      RECT 17.532 161.22 17.604 164.962 ; 
      RECT 17.388 161.22 17.46 164.962 ; 
      RECT 17.244 161.944 17.316 164.216 ; 
      RECT 20.952 165.54 21.024 169.282 ; 
      RECT 20.808 165.54 20.88 169.282 ; 
      RECT 20.664 167.848 20.736 169.138 ; 
      RECT 20.196 168.636 20.268 169.074 ; 
      RECT 20.16 165.67 20.232 166.628 ; 
      RECT 20.016 167.994 20.088 168.608 ; 
      RECT 19.692 168.096 19.764 169.128 ; 
      RECT 17.532 165.54 17.604 169.282 ; 
      RECT 17.388 165.54 17.46 169.282 ; 
      RECT 17.244 166.264 17.316 168.536 ; 
      RECT 20.952 169.86 21.024 173.602 ; 
      RECT 20.808 169.86 20.88 173.602 ; 
      RECT 20.664 172.168 20.736 173.458 ; 
      RECT 20.196 172.956 20.268 173.394 ; 
      RECT 20.16 169.99 20.232 170.948 ; 
      RECT 20.016 172.314 20.088 172.928 ; 
      RECT 19.692 172.416 19.764 173.448 ; 
      RECT 17.532 169.86 17.604 173.602 ; 
      RECT 17.388 169.86 17.46 173.602 ; 
      RECT 17.244 170.584 17.316 172.856 ; 
      RECT 37.62 188.944 37.692 206.366 ; 
      RECT 37.476 183.684 37.548 183.96 ; 
      RECT 37.476 190.916 37.548 192.774 ; 
      RECT 37.332 173.666 37.404 206.494 ; 
      RECT 37.188 188.744 37.26 191.834 ; 
      RECT 37.188 192.0388 37.26 194.004 ; 
      RECT 37.188 194.204 37.26 195.69 ; 
      RECT 37.188 195.942 37.26 199.188 ; 
      RECT 37.044 189.086 37.116 191.654 ; 
      RECT 37.044 194.364 37.116 196.492 ; 
      RECT 36.9 173.666 36.972 175.066 ; 
      RECT 36.468 173.666 36.54 175.066 ; 
      RECT 36.036 173.666 36.108 175.066 ; 
      RECT 35.604 173.666 35.676 175.066 ; 
      RECT 35.172 173.666 35.244 175.066 ; 
      RECT 34.74 173.666 34.812 175.066 ; 
      RECT 34.308 173.666 34.38 175.066 ; 
      RECT 33.876 173.666 33.948 175.066 ; 
      RECT 33.444 173.666 33.516 175.066 ; 
      RECT 33.012 173.666 33.084 175.066 ; 
      RECT 32.58 173.666 32.652 175.066 ; 
      RECT 32.148 173.666 32.22 175.066 ; 
      RECT 31.716 173.666 31.788 175.066 ; 
      RECT 31.284 173.666 31.356 175.066 ; 
      RECT 30.852 173.666 30.924 175.066 ; 
      RECT 30.42 173.666 30.492 175.066 ; 
      RECT 29.988 173.666 30.06 175.066 ; 
      RECT 29.556 173.666 29.628 175.066 ; 
      RECT 29.124 173.666 29.196 175.066 ; 
      RECT 28.692 173.666 28.764 175.066 ; 
      RECT 28.26 173.666 28.332 175.066 ; 
      RECT 27.828 173.666 27.9 175.066 ; 
      RECT 27.396 173.666 27.468 175.066 ; 
      RECT 26.964 173.666 27.036 175.066 ; 
      RECT 26.532 173.666 26.604 175.066 ; 
      RECT 26.1 173.666 26.172 175.066 ; 
      RECT 25.668 173.666 25.74 175.066 ; 
      RECT 25.236 173.666 25.308 175.066 ; 
      RECT 24.804 173.666 24.876 175.066 ; 
      RECT 24.372 173.666 24.444 175.066 ; 
      RECT 24.228 188.82 24.3 191.6388 ; 
      RECT 24.228 194.608 24.3 199.332 ; 
      RECT 24.156 176.308 24.228 179.012 ; 
      RECT 24.156 181.996 24.228 183.188 ; 
      RECT 24.084 189.074 24.156 191.834 ; 
      RECT 24.084 192.038 24.156 196.004 ; 
      RECT 24.084 196.124 24.156 199.26 ; 
      RECT 23.94 173.666 24.012 206.494 ; 
      RECT 23.796 190.164 23.868 190.496 ; 
      RECT 23.724 176.74 23.796 179.264 ; 
      RECT 23.724 180.916 23.796 181.676 ; 
      RECT 23.724 184.444 23.796 184.64 ; 
      RECT 23.652 188.944 23.724 206.384 ; 
      RECT 23.292 175.228 23.364 178.436 ; 
      RECT 23.292 180.628 23.364 182.9 ; 
      RECT 23.148 180.916 23.22 182.396 ; 
      RECT 23.004 178.324 23.076 178.868 ; 
      RECT 23.004 182.284 23.076 183.188 ; 
      RECT 23.004 187.252 23.076 187.508 ; 
      RECT 22.86 178.732 22.932 178.88 ; 
      RECT 22.86 185.236 22.932 185.408 ; 
      RECT 22.86 187.372 22.932 187.52 ; 
      RECT 22.716 179.98 22.788 181.964 ; 
      RECT 22.716 182.14 22.788 182.9 ; 
      RECT 22.716 185.98 22.788 187.22 ; 
      RECT 22.572 195.1 22.644 198.02 ; 
      RECT 22.572 199.42 22.644 202.34 ; 
      RECT 21.276 178.468 21.348 179.66 ; 
      RECT 21.276 183.22 21.348 183.476 ; 
      RECT 21.276 184.3 21.348 186.14 ; 
      RECT 21.276 189.1 21.348 189.248 ; 
      RECT 21.276 197.26 21.348 198.452 ; 
      RECT 21.132 178.756 21.204 180.776 ; 
      RECT 21.132 181.852 21.204 185.06 ; 
      RECT 21.132 189.232 21.204 190.316 ; 
      RECT 21.132 190.636 21.204 191.54 ; 
      RECT 20.988 178.468 21.06 181.172 ; 
      RECT 20.988 181.564 21.06 182.9 ; 
      RECT 20.988 183.724 21.06 184.268 ; 
      RECT 20.988 186.46 21.06 189.668 ; 
      RECT 20.988 191.404 21.06 191.552 ; 
      RECT 20.988 200.068 21.06 201.404 ; 
      RECT 20.844 179.404 20.916 179.948 ; 
      RECT 20.844 186.964 20.916 190.892 ; 
      RECT 20.844 192.652 20.916 193.844 ; 
      RECT 20.844 199.42 20.916 200.468 ; 
      RECT 20.7 175.66 20.772 176.276 ; 
      RECT 20.7 178.9 20.772 186.044 ; 
      RECT 20.7 190.204 20.772 199.532 ; 
      RECT 20.7 200.356 20.772 204.788 ; 
      RECT 19.548 176.74 19.62 177.788 ; 
      RECT 19.548 178.324 19.62 178.58 ; 
      RECT 19.548 178.9 19.62 179.804 ; 
      RECT 19.548 179.98 19.62 180.74 ; 
      RECT 19.548 181.06 19.62 191.54 ; 
      RECT 19.548 191.716 19.62 196.94 ; 
      RECT 19.548 201.292 19.62 202.34 ; 
      RECT 19.404 180.736 19.476 181.82 ; 
      RECT 19.404 182.14 19.476 185.492 ; 
      RECT 19.404 186.172 19.476 189.524 ; 
      RECT 19.404 189.7 19.476 194.78 ; 
      RECT 19.404 195.604 19.476 196.292 ; 
      RECT 19.404 199.132 19.476 203.42 ; 
      RECT 19.26 181.06 19.332 182.144 ; 
      RECT 19.26 182.764 19.332 182.912 ; 
      RECT 19.26 185.884 19.332 189.812 ; 
      RECT 19.26 190.78 19.332 192.62 ; 
      RECT 19.26 194.02 19.332 196.976 ; 
      RECT 19.116 177.532 19.188 181.82 ; 
      RECT 19.116 188.188 19.188 189.056 ; 
      RECT 19.116 193.732 19.188 194.924 ; 
      RECT 18.972 180.124 19.044 181.964 ; 
      RECT 18.972 186.46 19.044 187.22 ; 
      RECT 18.972 187.384 19.044 187.532 ; 
      RECT 18.972 188.476 19.044 189.812 ; 
      RECT 18.972 190.348 19.044 195.716 ; 
      RECT 18.972 196.144 19.044 200.612 ; 
      RECT 18.828 177.82 18.9 178.58 ; 
      RECT 18.828 179.404 18.9 179.948 ; 
      RECT 18.828 181.06 18.9 193.7 ; 
      RECT 18.828 194.02 18.9 195.86 ; 
      RECT 18.828 198.34 18.9 200.18 ; 
      RECT 18.828 203.596 18.9 204.5 ; 
      RECT 18.684 173.772 18.756 174.388 ; 
      RECT 18.684 205.816 18.756 206.432 ; 
      RECT 18.54 173.772 18.612 173.972 ; 
      RECT 18.252 173.772 18.324 174.058 ; 
      RECT 18.252 206.094 18.324 206.494 ; 
      RECT 17.676 179.836 17.748 180.596 ; 
      RECT 17.676 182.788 17.748 184.268 ; 
      RECT 17.676 190.636 17.748 191.54 ; 
      RECT 17.676 192.796 17.748 197.372 ; 
      RECT 17.676 200.5 17.748 202.34 ; 
      RECT 17.676 204.652 17.748 204.8 ; 
      RECT 17.532 175.66 17.604 177.644 ; 
      RECT 17.532 191.98 17.604 192.128 ; 
      RECT 17.532 196.288 17.604 199.532 ; 
      RECT 17.388 177.532 17.46 178.58 ; 
      RECT 17.388 179.692 17.46 181.028 ; 
      RECT 17.388 181.852 17.46 182.252 ; 
      RECT 17.388 185.38 17.46 196.436 ; 
      RECT 17.388 196.972 17.46 197.876 ; 
      RECT 17.244 176.164 17.316 180.74 ; 
      RECT 17.244 195.1 17.316 195.86 ; 
      RECT 17.244 198.316 17.316 198.464 ; 
      RECT 17.244 199.42 17.316 202.628 ; 
      RECT 17.1 179.98 17.172 183.98 ; 
      RECT 17.1 197.74 17.172 197.888 ; 
      RECT 16.956 176.74 17.028 176.852 ; 
      RECT 15.66 178.324 15.732 179.948 ; 
      RECT 15.372 178.468 15.444 180.884 ; 
      RECT 15.228 177.82 15.3 178.076 ; 
      RECT 15.084 173.984 15.156 174.188 ; 
      RECT 15.084 186.46 15.156 187.22 ; 
      RECT 15.084 188.944 15.156 206.384 ; 
      RECT 14.724 188.944 14.796 206.384 ; 
      RECT 14.652 175.66 14.724 176.42 ; 
      RECT 14.652 178.756 14.724 187.796 ; 
      RECT 14.58 190.164 14.652 190.496 ; 
      RECT 14.436 173.666 14.508 206.494 ; 
      RECT 14.292 189.074 14.364 191.834 ; 
      RECT 14.292 192.038 14.364 196.004 ; 
      RECT 14.292 196.124 14.364 199.26 ; 
      RECT 14.22 175.66 14.292 177.644 ; 
      RECT 14.22 180.772 14.292 183.044 ; 
      RECT 14.22 184.3 14.292 187.22 ; 
      RECT 14.148 188.82 14.22 191.6388 ; 
      RECT 14.148 194.608 14.22 199.332 ; 
      RECT 14.004 173.666 14.076 175.066 ; 
      RECT 13.572 173.666 13.644 175.066 ; 
      RECT 13.14 173.666 13.212 175.066 ; 
      RECT 12.708 173.666 12.78 175.066 ; 
      RECT 12.276 173.666 12.348 175.066 ; 
      RECT 11.844 173.666 11.916 175.066 ; 
      RECT 11.412 173.666 11.484 175.066 ; 
      RECT 10.98 173.666 11.052 175.066 ; 
      RECT 10.548 173.666 10.62 175.066 ; 
      RECT 10.116 173.666 10.188 175.066 ; 
      RECT 9.684 173.666 9.756 175.066 ; 
      RECT 9.252 173.666 9.324 175.066 ; 
      RECT 8.82 173.666 8.892 175.066 ; 
      RECT 8.388 173.666 8.46 175.066 ; 
      RECT 7.956 173.666 8.028 175.066 ; 
      RECT 7.524 173.666 7.596 175.066 ; 
      RECT 7.092 173.666 7.164 175.066 ; 
      RECT 6.66 173.666 6.732 175.066 ; 
      RECT 6.228 173.666 6.3 175.066 ; 
      RECT 5.796 173.666 5.868 175.066 ; 
      RECT 5.364 173.666 5.436 175.066 ; 
      RECT 4.932 173.666 5.004 175.066 ; 
      RECT 4.5 173.666 4.572 175.066 ; 
      RECT 4.068 173.666 4.14 175.066 ; 
      RECT 3.636 173.666 3.708 175.066 ; 
      RECT 3.204 173.666 3.276 175.066 ; 
      RECT 2.772 173.666 2.844 175.066 ; 
      RECT 2.34 173.666 2.412 175.066 ; 
      RECT 1.908 173.666 1.98 175.066 ; 
      RECT 1.476 173.666 1.548 175.066 ; 
      RECT 1.332 189.086 1.404 191.654 ; 
      RECT 1.332 194.364 1.404 196.492 ; 
      RECT 1.26 177.82 1.332 178.724 ; 
      RECT 1.188 188.744 1.26 191.834 ; 
      RECT 1.188 192.0388 1.26 194.004 ; 
      RECT 1.188 194.204 1.26 195.69 ; 
      RECT 1.188 195.942 1.26 199.188 ; 
      RECT 1.044 173.666 1.116 206.494 ; 
      RECT 0.9 183.684 0.972 183.96 ; 
      RECT 0.9 190.916 0.972 192.774 ; 
      RECT 0.756 188.944 0.828 206.366 ; 
        RECT 20.952 206.688 21.024 210.43 ; 
        RECT 20.808 206.688 20.88 210.43 ; 
        RECT 20.664 208.996 20.736 210.286 ; 
        RECT 20.196 209.784 20.268 210.222 ; 
        RECT 20.16 206.818 20.232 207.776 ; 
        RECT 20.016 209.142 20.088 209.756 ; 
        RECT 19.692 209.244 19.764 210.276 ; 
        RECT 17.532 206.688 17.604 210.43 ; 
        RECT 17.388 206.688 17.46 210.43 ; 
        RECT 17.244 207.412 17.316 209.684 ; 
        RECT 20.952 211.008 21.024 214.75 ; 
        RECT 20.808 211.008 20.88 214.75 ; 
        RECT 20.664 213.316 20.736 214.606 ; 
        RECT 20.196 214.104 20.268 214.542 ; 
        RECT 20.16 211.138 20.232 212.096 ; 
        RECT 20.016 213.462 20.088 214.076 ; 
        RECT 19.692 213.564 19.764 214.596 ; 
        RECT 17.532 211.008 17.604 214.75 ; 
        RECT 17.388 211.008 17.46 214.75 ; 
        RECT 17.244 211.732 17.316 214.004 ; 
        RECT 20.952 215.328 21.024 219.07 ; 
        RECT 20.808 215.328 20.88 219.07 ; 
        RECT 20.664 217.636 20.736 218.926 ; 
        RECT 20.196 218.424 20.268 218.862 ; 
        RECT 20.16 215.458 20.232 216.416 ; 
        RECT 20.016 217.782 20.088 218.396 ; 
        RECT 19.692 217.884 19.764 218.916 ; 
        RECT 17.532 215.328 17.604 219.07 ; 
        RECT 17.388 215.328 17.46 219.07 ; 
        RECT 17.244 216.052 17.316 218.324 ; 
        RECT 20.952 219.648 21.024 223.39 ; 
        RECT 20.808 219.648 20.88 223.39 ; 
        RECT 20.664 221.956 20.736 223.246 ; 
        RECT 20.196 222.744 20.268 223.182 ; 
        RECT 20.16 219.778 20.232 220.736 ; 
        RECT 20.016 222.102 20.088 222.716 ; 
        RECT 19.692 222.204 19.764 223.236 ; 
        RECT 17.532 219.648 17.604 223.39 ; 
        RECT 17.388 219.648 17.46 223.39 ; 
        RECT 17.244 220.372 17.316 222.644 ; 
        RECT 20.952 223.968 21.024 227.71 ; 
        RECT 20.808 223.968 20.88 227.71 ; 
        RECT 20.664 226.276 20.736 227.566 ; 
        RECT 20.196 227.064 20.268 227.502 ; 
        RECT 20.16 224.098 20.232 225.056 ; 
        RECT 20.016 226.422 20.088 227.036 ; 
        RECT 19.692 226.524 19.764 227.556 ; 
        RECT 17.532 223.968 17.604 227.71 ; 
        RECT 17.388 223.968 17.46 227.71 ; 
        RECT 17.244 224.692 17.316 226.964 ; 
        RECT 20.952 228.288 21.024 232.03 ; 
        RECT 20.808 228.288 20.88 232.03 ; 
        RECT 20.664 230.596 20.736 231.886 ; 
        RECT 20.196 231.384 20.268 231.822 ; 
        RECT 20.16 228.418 20.232 229.376 ; 
        RECT 20.016 230.742 20.088 231.356 ; 
        RECT 19.692 230.844 19.764 231.876 ; 
        RECT 17.532 228.288 17.604 232.03 ; 
        RECT 17.388 228.288 17.46 232.03 ; 
        RECT 17.244 229.012 17.316 231.284 ; 
        RECT 20.952 232.608 21.024 236.35 ; 
        RECT 20.808 232.608 20.88 236.35 ; 
        RECT 20.664 234.916 20.736 236.206 ; 
        RECT 20.196 235.704 20.268 236.142 ; 
        RECT 20.16 232.738 20.232 233.696 ; 
        RECT 20.016 235.062 20.088 235.676 ; 
        RECT 19.692 235.164 19.764 236.196 ; 
        RECT 17.532 232.608 17.604 236.35 ; 
        RECT 17.388 232.608 17.46 236.35 ; 
        RECT 17.244 233.332 17.316 235.604 ; 
        RECT 20.952 236.928 21.024 240.67 ; 
        RECT 20.808 236.928 20.88 240.67 ; 
        RECT 20.664 239.236 20.736 240.526 ; 
        RECT 20.196 240.024 20.268 240.462 ; 
        RECT 20.16 237.058 20.232 238.016 ; 
        RECT 20.016 239.382 20.088 239.996 ; 
        RECT 19.692 239.484 19.764 240.516 ; 
        RECT 17.532 236.928 17.604 240.67 ; 
        RECT 17.388 236.928 17.46 240.67 ; 
        RECT 17.244 237.652 17.316 239.924 ; 
        RECT 20.952 241.248 21.024 244.99 ; 
        RECT 20.808 241.248 20.88 244.99 ; 
        RECT 20.664 243.556 20.736 244.846 ; 
        RECT 20.196 244.344 20.268 244.782 ; 
        RECT 20.16 241.378 20.232 242.336 ; 
        RECT 20.016 243.702 20.088 244.316 ; 
        RECT 19.692 243.804 19.764 244.836 ; 
        RECT 17.532 241.248 17.604 244.99 ; 
        RECT 17.388 241.248 17.46 244.99 ; 
        RECT 17.244 241.972 17.316 244.244 ; 
        RECT 20.952 245.568 21.024 249.31 ; 
        RECT 20.808 245.568 20.88 249.31 ; 
        RECT 20.664 247.876 20.736 249.166 ; 
        RECT 20.196 248.664 20.268 249.102 ; 
        RECT 20.16 245.698 20.232 246.656 ; 
        RECT 20.016 248.022 20.088 248.636 ; 
        RECT 19.692 248.124 19.764 249.156 ; 
        RECT 17.532 245.568 17.604 249.31 ; 
        RECT 17.388 245.568 17.46 249.31 ; 
        RECT 17.244 246.292 17.316 248.564 ; 
        RECT 20.952 249.888 21.024 253.63 ; 
        RECT 20.808 249.888 20.88 253.63 ; 
        RECT 20.664 252.196 20.736 253.486 ; 
        RECT 20.196 252.984 20.268 253.422 ; 
        RECT 20.16 250.018 20.232 250.976 ; 
        RECT 20.016 252.342 20.088 252.956 ; 
        RECT 19.692 252.444 19.764 253.476 ; 
        RECT 17.532 249.888 17.604 253.63 ; 
        RECT 17.388 249.888 17.46 253.63 ; 
        RECT 17.244 250.612 17.316 252.884 ; 
        RECT 20.952 254.208 21.024 257.95 ; 
        RECT 20.808 254.208 20.88 257.95 ; 
        RECT 20.664 256.516 20.736 257.806 ; 
        RECT 20.196 257.304 20.268 257.742 ; 
        RECT 20.16 254.338 20.232 255.296 ; 
        RECT 20.016 256.662 20.088 257.276 ; 
        RECT 19.692 256.764 19.764 257.796 ; 
        RECT 17.532 254.208 17.604 257.95 ; 
        RECT 17.388 254.208 17.46 257.95 ; 
        RECT 17.244 254.932 17.316 257.204 ; 
        RECT 20.952 258.528 21.024 262.27 ; 
        RECT 20.808 258.528 20.88 262.27 ; 
        RECT 20.664 260.836 20.736 262.126 ; 
        RECT 20.196 261.624 20.268 262.062 ; 
        RECT 20.16 258.658 20.232 259.616 ; 
        RECT 20.016 260.982 20.088 261.596 ; 
        RECT 19.692 261.084 19.764 262.116 ; 
        RECT 17.532 258.528 17.604 262.27 ; 
        RECT 17.388 258.528 17.46 262.27 ; 
        RECT 17.244 259.252 17.316 261.524 ; 
        RECT 20.952 262.848 21.024 266.59 ; 
        RECT 20.808 262.848 20.88 266.59 ; 
        RECT 20.664 265.156 20.736 266.446 ; 
        RECT 20.196 265.944 20.268 266.382 ; 
        RECT 20.16 262.978 20.232 263.936 ; 
        RECT 20.016 265.302 20.088 265.916 ; 
        RECT 19.692 265.404 19.764 266.436 ; 
        RECT 17.532 262.848 17.604 266.59 ; 
        RECT 17.388 262.848 17.46 266.59 ; 
        RECT 17.244 263.572 17.316 265.844 ; 
        RECT 20.952 267.168 21.024 270.91 ; 
        RECT 20.808 267.168 20.88 270.91 ; 
        RECT 20.664 269.476 20.736 270.766 ; 
        RECT 20.196 270.264 20.268 270.702 ; 
        RECT 20.16 267.298 20.232 268.256 ; 
        RECT 20.016 269.622 20.088 270.236 ; 
        RECT 19.692 269.724 19.764 270.756 ; 
        RECT 17.532 267.168 17.604 270.91 ; 
        RECT 17.388 267.168 17.46 270.91 ; 
        RECT 17.244 267.892 17.316 270.164 ; 
        RECT 20.952 271.488 21.024 275.23 ; 
        RECT 20.808 271.488 20.88 275.23 ; 
        RECT 20.664 273.796 20.736 275.086 ; 
        RECT 20.196 274.584 20.268 275.022 ; 
        RECT 20.16 271.618 20.232 272.576 ; 
        RECT 20.016 273.942 20.088 274.556 ; 
        RECT 19.692 274.044 19.764 275.076 ; 
        RECT 17.532 271.488 17.604 275.23 ; 
        RECT 17.388 271.488 17.46 275.23 ; 
        RECT 17.244 272.212 17.316 274.484 ; 
        RECT 20.952 275.808 21.024 279.55 ; 
        RECT 20.808 275.808 20.88 279.55 ; 
        RECT 20.664 278.116 20.736 279.406 ; 
        RECT 20.196 278.904 20.268 279.342 ; 
        RECT 20.16 275.938 20.232 276.896 ; 
        RECT 20.016 278.262 20.088 278.876 ; 
        RECT 19.692 278.364 19.764 279.396 ; 
        RECT 17.532 275.808 17.604 279.55 ; 
        RECT 17.388 275.808 17.46 279.55 ; 
        RECT 17.244 276.532 17.316 278.804 ; 
        RECT 20.952 280.128 21.024 283.87 ; 
        RECT 20.808 280.128 20.88 283.87 ; 
        RECT 20.664 282.436 20.736 283.726 ; 
        RECT 20.196 283.224 20.268 283.662 ; 
        RECT 20.16 280.258 20.232 281.216 ; 
        RECT 20.016 282.582 20.088 283.196 ; 
        RECT 19.692 282.684 19.764 283.716 ; 
        RECT 17.532 280.128 17.604 283.87 ; 
        RECT 17.388 280.128 17.46 283.87 ; 
        RECT 17.244 280.852 17.316 283.124 ; 
        RECT 20.952 284.448 21.024 288.19 ; 
        RECT 20.808 284.448 20.88 288.19 ; 
        RECT 20.664 286.756 20.736 288.046 ; 
        RECT 20.196 287.544 20.268 287.982 ; 
        RECT 20.16 284.578 20.232 285.536 ; 
        RECT 20.016 286.902 20.088 287.516 ; 
        RECT 19.692 287.004 19.764 288.036 ; 
        RECT 17.532 284.448 17.604 288.19 ; 
        RECT 17.388 284.448 17.46 288.19 ; 
        RECT 17.244 285.172 17.316 287.444 ; 
        RECT 20.952 288.768 21.024 292.51 ; 
        RECT 20.808 288.768 20.88 292.51 ; 
        RECT 20.664 291.076 20.736 292.366 ; 
        RECT 20.196 291.864 20.268 292.302 ; 
        RECT 20.16 288.898 20.232 289.856 ; 
        RECT 20.016 291.222 20.088 291.836 ; 
        RECT 19.692 291.324 19.764 292.356 ; 
        RECT 17.532 288.768 17.604 292.51 ; 
        RECT 17.388 288.768 17.46 292.51 ; 
        RECT 17.244 289.492 17.316 291.764 ; 
        RECT 20.952 293.088 21.024 296.83 ; 
        RECT 20.808 293.088 20.88 296.83 ; 
        RECT 20.664 295.396 20.736 296.686 ; 
        RECT 20.196 296.184 20.268 296.622 ; 
        RECT 20.16 293.218 20.232 294.176 ; 
        RECT 20.016 295.542 20.088 296.156 ; 
        RECT 19.692 295.644 19.764 296.676 ; 
        RECT 17.532 293.088 17.604 296.83 ; 
        RECT 17.388 293.088 17.46 296.83 ; 
        RECT 17.244 293.812 17.316 296.084 ; 
        RECT 20.952 297.408 21.024 301.15 ; 
        RECT 20.808 297.408 20.88 301.15 ; 
        RECT 20.664 299.716 20.736 301.006 ; 
        RECT 20.196 300.504 20.268 300.942 ; 
        RECT 20.16 297.538 20.232 298.496 ; 
        RECT 20.016 299.862 20.088 300.476 ; 
        RECT 19.692 299.964 19.764 300.996 ; 
        RECT 17.532 297.408 17.604 301.15 ; 
        RECT 17.388 297.408 17.46 301.15 ; 
        RECT 17.244 298.132 17.316 300.404 ; 
        RECT 20.952 301.728 21.024 305.47 ; 
        RECT 20.808 301.728 20.88 305.47 ; 
        RECT 20.664 304.036 20.736 305.326 ; 
        RECT 20.196 304.824 20.268 305.262 ; 
        RECT 20.16 301.858 20.232 302.816 ; 
        RECT 20.016 304.182 20.088 304.796 ; 
        RECT 19.692 304.284 19.764 305.316 ; 
        RECT 17.532 301.728 17.604 305.47 ; 
        RECT 17.388 301.728 17.46 305.47 ; 
        RECT 17.244 302.452 17.316 304.724 ; 
        RECT 20.952 306.048 21.024 309.79 ; 
        RECT 20.808 306.048 20.88 309.79 ; 
        RECT 20.664 308.356 20.736 309.646 ; 
        RECT 20.196 309.144 20.268 309.582 ; 
        RECT 20.16 306.178 20.232 307.136 ; 
        RECT 20.016 308.502 20.088 309.116 ; 
        RECT 19.692 308.604 19.764 309.636 ; 
        RECT 17.532 306.048 17.604 309.79 ; 
        RECT 17.388 306.048 17.46 309.79 ; 
        RECT 17.244 306.772 17.316 309.044 ; 
        RECT 20.952 310.368 21.024 314.11 ; 
        RECT 20.808 310.368 20.88 314.11 ; 
        RECT 20.664 312.676 20.736 313.966 ; 
        RECT 20.196 313.464 20.268 313.902 ; 
        RECT 20.16 310.498 20.232 311.456 ; 
        RECT 20.016 312.822 20.088 313.436 ; 
        RECT 19.692 312.924 19.764 313.956 ; 
        RECT 17.532 310.368 17.604 314.11 ; 
        RECT 17.388 310.368 17.46 314.11 ; 
        RECT 17.244 311.092 17.316 313.364 ; 
        RECT 20.952 314.688 21.024 318.43 ; 
        RECT 20.808 314.688 20.88 318.43 ; 
        RECT 20.664 316.996 20.736 318.286 ; 
        RECT 20.196 317.784 20.268 318.222 ; 
        RECT 20.16 314.818 20.232 315.776 ; 
        RECT 20.016 317.142 20.088 317.756 ; 
        RECT 19.692 317.244 19.764 318.276 ; 
        RECT 17.532 314.688 17.604 318.43 ; 
        RECT 17.388 314.688 17.46 318.43 ; 
        RECT 17.244 315.412 17.316 317.684 ; 
        RECT 20.952 319.008 21.024 322.75 ; 
        RECT 20.808 319.008 20.88 322.75 ; 
        RECT 20.664 321.316 20.736 322.606 ; 
        RECT 20.196 322.104 20.268 322.542 ; 
        RECT 20.16 319.138 20.232 320.096 ; 
        RECT 20.016 321.462 20.088 322.076 ; 
        RECT 19.692 321.564 19.764 322.596 ; 
        RECT 17.532 319.008 17.604 322.75 ; 
        RECT 17.388 319.008 17.46 322.75 ; 
        RECT 17.244 319.732 17.316 322.004 ; 
        RECT 20.952 323.328 21.024 327.07 ; 
        RECT 20.808 323.328 20.88 327.07 ; 
        RECT 20.664 325.636 20.736 326.926 ; 
        RECT 20.196 326.424 20.268 326.862 ; 
        RECT 20.16 323.458 20.232 324.416 ; 
        RECT 20.016 325.782 20.088 326.396 ; 
        RECT 19.692 325.884 19.764 326.916 ; 
        RECT 17.532 323.328 17.604 327.07 ; 
        RECT 17.388 323.328 17.46 327.07 ; 
        RECT 17.244 324.052 17.316 326.324 ; 
        RECT 20.952 327.648 21.024 331.39 ; 
        RECT 20.808 327.648 20.88 331.39 ; 
        RECT 20.664 329.956 20.736 331.246 ; 
        RECT 20.196 330.744 20.268 331.182 ; 
        RECT 20.16 327.778 20.232 328.736 ; 
        RECT 20.016 330.102 20.088 330.716 ; 
        RECT 19.692 330.204 19.764 331.236 ; 
        RECT 17.532 327.648 17.604 331.39 ; 
        RECT 17.388 327.648 17.46 331.39 ; 
        RECT 17.244 328.372 17.316 330.644 ; 
        RECT 20.952 331.968 21.024 335.71 ; 
        RECT 20.808 331.968 20.88 335.71 ; 
        RECT 20.664 334.276 20.736 335.566 ; 
        RECT 20.196 335.064 20.268 335.502 ; 
        RECT 20.16 332.098 20.232 333.056 ; 
        RECT 20.016 334.422 20.088 335.036 ; 
        RECT 19.692 334.524 19.764 335.556 ; 
        RECT 17.532 331.968 17.604 335.71 ; 
        RECT 17.388 331.968 17.46 335.71 ; 
        RECT 17.244 332.692 17.316 334.964 ; 
        RECT 20.952 336.288 21.024 340.03 ; 
        RECT 20.808 336.288 20.88 340.03 ; 
        RECT 20.664 338.596 20.736 339.886 ; 
        RECT 20.196 339.384 20.268 339.822 ; 
        RECT 20.16 336.418 20.232 337.376 ; 
        RECT 20.016 338.742 20.088 339.356 ; 
        RECT 19.692 338.844 19.764 339.876 ; 
        RECT 17.532 336.288 17.604 340.03 ; 
        RECT 17.388 336.288 17.46 340.03 ; 
        RECT 17.244 337.012 17.316 339.284 ; 
        RECT 20.952 340.608 21.024 344.35 ; 
        RECT 20.808 340.608 20.88 344.35 ; 
        RECT 20.664 342.916 20.736 344.206 ; 
        RECT 20.196 343.704 20.268 344.142 ; 
        RECT 20.16 340.738 20.232 341.696 ; 
        RECT 20.016 343.062 20.088 343.676 ; 
        RECT 19.692 343.164 19.764 344.196 ; 
        RECT 17.532 340.608 17.604 344.35 ; 
        RECT 17.388 340.608 17.46 344.35 ; 
        RECT 17.244 341.332 17.316 343.604 ; 
        RECT 20.952 344.928 21.024 348.67 ; 
        RECT 20.808 344.928 20.88 348.67 ; 
        RECT 20.664 347.236 20.736 348.526 ; 
        RECT 20.196 348.024 20.268 348.462 ; 
        RECT 20.16 345.058 20.232 346.016 ; 
        RECT 20.016 347.382 20.088 347.996 ; 
        RECT 19.692 347.484 19.764 348.516 ; 
        RECT 17.532 344.928 17.604 348.67 ; 
        RECT 17.388 344.928 17.46 348.67 ; 
        RECT 17.244 345.652 17.316 347.924 ; 
        RECT 20.952 349.248 21.024 352.99 ; 
        RECT 20.808 349.248 20.88 352.99 ; 
        RECT 20.664 351.556 20.736 352.846 ; 
        RECT 20.196 352.344 20.268 352.782 ; 
        RECT 20.16 349.378 20.232 350.336 ; 
        RECT 20.016 351.702 20.088 352.316 ; 
        RECT 19.692 351.804 19.764 352.836 ; 
        RECT 17.532 349.248 17.604 352.99 ; 
        RECT 17.388 349.248 17.46 352.99 ; 
        RECT 17.244 349.972 17.316 352.244 ; 
        RECT 20.952 353.568 21.024 357.31 ; 
        RECT 20.808 353.568 20.88 357.31 ; 
        RECT 20.664 355.876 20.736 357.166 ; 
        RECT 20.196 356.664 20.268 357.102 ; 
        RECT 20.16 353.698 20.232 354.656 ; 
        RECT 20.016 356.022 20.088 356.636 ; 
        RECT 19.692 356.124 19.764 357.156 ; 
        RECT 17.532 353.568 17.604 357.31 ; 
        RECT 17.388 353.568 17.46 357.31 ; 
        RECT 17.244 354.292 17.316 356.564 ; 
        RECT 20.952 357.888 21.024 361.63 ; 
        RECT 20.808 357.888 20.88 361.63 ; 
        RECT 20.664 360.196 20.736 361.486 ; 
        RECT 20.196 360.984 20.268 361.422 ; 
        RECT 20.16 358.018 20.232 358.976 ; 
        RECT 20.016 360.342 20.088 360.956 ; 
        RECT 19.692 360.444 19.764 361.476 ; 
        RECT 17.532 357.888 17.604 361.63 ; 
        RECT 17.388 357.888 17.46 361.63 ; 
        RECT 17.244 358.612 17.316 360.884 ; 
        RECT 20.952 362.208 21.024 365.95 ; 
        RECT 20.808 362.208 20.88 365.95 ; 
        RECT 20.664 364.516 20.736 365.806 ; 
        RECT 20.196 365.304 20.268 365.742 ; 
        RECT 20.16 362.338 20.232 363.296 ; 
        RECT 20.016 364.662 20.088 365.276 ; 
        RECT 19.692 364.764 19.764 365.796 ; 
        RECT 17.532 362.208 17.604 365.95 ; 
        RECT 17.388 362.208 17.46 365.95 ; 
        RECT 17.244 362.932 17.316 365.204 ; 
        RECT 20.952 366.528 21.024 370.27 ; 
        RECT 20.808 366.528 20.88 370.27 ; 
        RECT 20.664 368.836 20.736 370.126 ; 
        RECT 20.196 369.624 20.268 370.062 ; 
        RECT 20.16 366.658 20.232 367.616 ; 
        RECT 20.016 368.982 20.088 369.596 ; 
        RECT 19.692 369.084 19.764 370.116 ; 
        RECT 17.532 366.528 17.604 370.27 ; 
        RECT 17.388 366.528 17.46 370.27 ; 
        RECT 17.244 367.252 17.316 369.524 ; 
        RECT 20.952 370.848 21.024 374.59 ; 
        RECT 20.808 370.848 20.88 374.59 ; 
        RECT 20.664 373.156 20.736 374.446 ; 
        RECT 20.196 373.944 20.268 374.382 ; 
        RECT 20.16 370.978 20.232 371.936 ; 
        RECT 20.016 373.302 20.088 373.916 ; 
        RECT 19.692 373.404 19.764 374.436 ; 
        RECT 17.532 370.848 17.604 374.59 ; 
        RECT 17.388 370.848 17.46 374.59 ; 
        RECT 17.244 371.572 17.316 373.844 ; 
        RECT 20.952 375.168 21.024 378.91 ; 
        RECT 20.808 375.168 20.88 378.91 ; 
        RECT 20.664 377.476 20.736 378.766 ; 
        RECT 20.196 378.264 20.268 378.702 ; 
        RECT 20.16 375.298 20.232 376.256 ; 
        RECT 20.016 377.622 20.088 378.236 ; 
        RECT 19.692 377.724 19.764 378.756 ; 
        RECT 17.532 375.168 17.604 378.91 ; 
        RECT 17.388 375.168 17.46 378.91 ; 
        RECT 17.244 375.892 17.316 378.164 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 20.72 1.026 21.232 5.4 ; 
      RECT 20.664 3.688 21.232 4.978 ; 
      RECT 20.072 2.596 20.32 5.4 ; 
      RECT 20.016 3.834 20.32 4.448 ; 
      RECT 20.072 1.026 20.176 5.4 ; 
      RECT 20.072 1.51 20.232 2.468 ; 
      RECT 20.072 1.026 20.32 1.382 ; 
      RECT 18.884 2.828 19.708 5.4 ; 
      RECT 19.604 1.026 19.708 5.4 ; 
      RECT 18.884 3.936 19.764 4.968 ; 
      RECT 18.884 1.026 19.276 5.4 ; 
      RECT 17.216 1.026 17.548 5.4 ; 
      RECT 17.216 1.38 17.604 5.122 ; 
      RECT 38.108 1.026 38.448 5.4 ; 
      RECT 37.532 1.026 37.636 5.4 ; 
      RECT 37.1 1.026 37.204 5.4 ; 
      RECT 36.668 1.026 36.772 5.4 ; 
      RECT 36.236 1.026 36.34 5.4 ; 
      RECT 35.804 1.026 35.908 5.4 ; 
      RECT 35.372 1.026 35.476 5.4 ; 
      RECT 34.94 1.026 35.044 5.4 ; 
      RECT 34.508 1.026 34.612 5.4 ; 
      RECT 34.076 1.026 34.18 5.4 ; 
      RECT 33.644 1.026 33.748 5.4 ; 
      RECT 33.212 1.026 33.316 5.4 ; 
      RECT 32.78 1.026 32.884 5.4 ; 
      RECT 32.348 1.026 32.452 5.4 ; 
      RECT 31.916 1.026 32.02 5.4 ; 
      RECT 31.484 1.026 31.588 5.4 ; 
      RECT 31.052 1.026 31.156 5.4 ; 
      RECT 30.62 1.026 30.724 5.4 ; 
      RECT 30.188 1.026 30.292 5.4 ; 
      RECT 29.756 1.026 29.86 5.4 ; 
      RECT 29.324 1.026 29.428 5.4 ; 
      RECT 28.892 1.026 28.996 5.4 ; 
      RECT 28.46 1.026 28.564 5.4 ; 
      RECT 28.028 1.026 28.132 5.4 ; 
      RECT 27.596 1.026 27.7 5.4 ; 
      RECT 27.164 1.026 27.268 5.4 ; 
      RECT 26.732 1.026 26.836 5.4 ; 
      RECT 26.3 1.026 26.404 5.4 ; 
      RECT 25.868 1.026 25.972 5.4 ; 
      RECT 25.436 1.026 25.54 5.4 ; 
      RECT 25.004 1.026 25.108 5.4 ; 
      RECT 24.572 1.026 24.676 5.4 ; 
      RECT 24.14 1.026 24.244 5.4 ; 
      RECT 23.708 1.026 23.812 5.4 ; 
      RECT 22.856 1.026 23.164 5.4 ; 
      RECT 15.284 1.026 15.592 5.4 ; 
      RECT 14.636 1.026 14.74 5.4 ; 
      RECT 14.204 1.026 14.308 5.4 ; 
      RECT 13.772 1.026 13.876 5.4 ; 
      RECT 13.34 1.026 13.444 5.4 ; 
      RECT 12.908 1.026 13.012 5.4 ; 
      RECT 12.476 1.026 12.58 5.4 ; 
      RECT 12.044 1.026 12.148 5.4 ; 
      RECT 11.612 1.026 11.716 5.4 ; 
      RECT 11.18 1.026 11.284 5.4 ; 
      RECT 10.748 1.026 10.852 5.4 ; 
      RECT 10.316 1.026 10.42 5.4 ; 
      RECT 9.884 1.026 9.988 5.4 ; 
      RECT 9.452 1.026 9.556 5.4 ; 
      RECT 9.02 1.026 9.124 5.4 ; 
      RECT 8.588 1.026 8.692 5.4 ; 
      RECT 8.156 1.026 8.26 5.4 ; 
      RECT 7.724 1.026 7.828 5.4 ; 
      RECT 7.292 1.026 7.396 5.4 ; 
      RECT 6.86 1.026 6.964 5.4 ; 
      RECT 6.428 1.026 6.532 5.4 ; 
      RECT 5.996 1.026 6.1 5.4 ; 
      RECT 5.564 1.026 5.668 5.4 ; 
      RECT 5.132 1.026 5.236 5.4 ; 
      RECT 4.7 1.026 4.804 5.4 ; 
      RECT 4.268 1.026 4.372 5.4 ; 
      RECT 3.836 1.026 3.94 5.4 ; 
      RECT 3.404 1.026 3.508 5.4 ; 
      RECT 2.972 1.026 3.076 5.4 ; 
      RECT 2.54 1.026 2.644 5.4 ; 
      RECT 2.108 1.026 2.212 5.4 ; 
      RECT 1.676 1.026 1.78 5.4 ; 
      RECT 1.244 1.026 1.348 5.4 ; 
      RECT 0.812 1.026 0.916 5.4 ; 
      RECT 0 1.026 0.34 5.4 ; 
      RECT 20.72 5.346 21.232 9.72 ; 
      RECT 20.664 8.008 21.232 9.298 ; 
      RECT 20.072 6.916 20.32 9.72 ; 
      RECT 20.016 8.154 20.32 8.768 ; 
      RECT 20.072 5.346 20.176 9.72 ; 
      RECT 20.072 5.83 20.232 6.788 ; 
      RECT 20.072 5.346 20.32 5.702 ; 
      RECT 18.884 7.148 19.708 9.72 ; 
      RECT 19.604 5.346 19.708 9.72 ; 
      RECT 18.884 8.256 19.764 9.288 ; 
      RECT 18.884 5.346 19.276 9.72 ; 
      RECT 17.216 5.346 17.548 9.72 ; 
      RECT 17.216 5.7 17.604 9.442 ; 
      RECT 38.108 5.346 38.448 9.72 ; 
      RECT 37.532 5.346 37.636 9.72 ; 
      RECT 37.1 5.346 37.204 9.72 ; 
      RECT 36.668 5.346 36.772 9.72 ; 
      RECT 36.236 5.346 36.34 9.72 ; 
      RECT 35.804 5.346 35.908 9.72 ; 
      RECT 35.372 5.346 35.476 9.72 ; 
      RECT 34.94 5.346 35.044 9.72 ; 
      RECT 34.508 5.346 34.612 9.72 ; 
      RECT 34.076 5.346 34.18 9.72 ; 
      RECT 33.644 5.346 33.748 9.72 ; 
      RECT 33.212 5.346 33.316 9.72 ; 
      RECT 32.78 5.346 32.884 9.72 ; 
      RECT 32.348 5.346 32.452 9.72 ; 
      RECT 31.916 5.346 32.02 9.72 ; 
      RECT 31.484 5.346 31.588 9.72 ; 
      RECT 31.052 5.346 31.156 9.72 ; 
      RECT 30.62 5.346 30.724 9.72 ; 
      RECT 30.188 5.346 30.292 9.72 ; 
      RECT 29.756 5.346 29.86 9.72 ; 
      RECT 29.324 5.346 29.428 9.72 ; 
      RECT 28.892 5.346 28.996 9.72 ; 
      RECT 28.46 5.346 28.564 9.72 ; 
      RECT 28.028 5.346 28.132 9.72 ; 
      RECT 27.596 5.346 27.7 9.72 ; 
      RECT 27.164 5.346 27.268 9.72 ; 
      RECT 26.732 5.346 26.836 9.72 ; 
      RECT 26.3 5.346 26.404 9.72 ; 
      RECT 25.868 5.346 25.972 9.72 ; 
      RECT 25.436 5.346 25.54 9.72 ; 
      RECT 25.004 5.346 25.108 9.72 ; 
      RECT 24.572 5.346 24.676 9.72 ; 
      RECT 24.14 5.346 24.244 9.72 ; 
      RECT 23.708 5.346 23.812 9.72 ; 
      RECT 22.856 5.346 23.164 9.72 ; 
      RECT 15.284 5.346 15.592 9.72 ; 
      RECT 14.636 5.346 14.74 9.72 ; 
      RECT 14.204 5.346 14.308 9.72 ; 
      RECT 13.772 5.346 13.876 9.72 ; 
      RECT 13.34 5.346 13.444 9.72 ; 
      RECT 12.908 5.346 13.012 9.72 ; 
      RECT 12.476 5.346 12.58 9.72 ; 
      RECT 12.044 5.346 12.148 9.72 ; 
      RECT 11.612 5.346 11.716 9.72 ; 
      RECT 11.18 5.346 11.284 9.72 ; 
      RECT 10.748 5.346 10.852 9.72 ; 
      RECT 10.316 5.346 10.42 9.72 ; 
      RECT 9.884 5.346 9.988 9.72 ; 
      RECT 9.452 5.346 9.556 9.72 ; 
      RECT 9.02 5.346 9.124 9.72 ; 
      RECT 8.588 5.346 8.692 9.72 ; 
      RECT 8.156 5.346 8.26 9.72 ; 
      RECT 7.724 5.346 7.828 9.72 ; 
      RECT 7.292 5.346 7.396 9.72 ; 
      RECT 6.86 5.346 6.964 9.72 ; 
      RECT 6.428 5.346 6.532 9.72 ; 
      RECT 5.996 5.346 6.1 9.72 ; 
      RECT 5.564 5.346 5.668 9.72 ; 
      RECT 5.132 5.346 5.236 9.72 ; 
      RECT 4.7 5.346 4.804 9.72 ; 
      RECT 4.268 5.346 4.372 9.72 ; 
      RECT 3.836 5.346 3.94 9.72 ; 
      RECT 3.404 5.346 3.508 9.72 ; 
      RECT 2.972 5.346 3.076 9.72 ; 
      RECT 2.54 5.346 2.644 9.72 ; 
      RECT 2.108 5.346 2.212 9.72 ; 
      RECT 1.676 5.346 1.78 9.72 ; 
      RECT 1.244 5.346 1.348 9.72 ; 
      RECT 0.812 5.346 0.916 9.72 ; 
      RECT 0 5.346 0.34 9.72 ; 
      RECT 20.72 9.666 21.232 14.04 ; 
      RECT 20.664 12.328 21.232 13.618 ; 
      RECT 20.072 11.236 20.32 14.04 ; 
      RECT 20.016 12.474 20.32 13.088 ; 
      RECT 20.072 9.666 20.176 14.04 ; 
      RECT 20.072 10.15 20.232 11.108 ; 
      RECT 20.072 9.666 20.32 10.022 ; 
      RECT 18.884 11.468 19.708 14.04 ; 
      RECT 19.604 9.666 19.708 14.04 ; 
      RECT 18.884 12.576 19.764 13.608 ; 
      RECT 18.884 9.666 19.276 14.04 ; 
      RECT 17.216 9.666 17.548 14.04 ; 
      RECT 17.216 10.02 17.604 13.762 ; 
      RECT 38.108 9.666 38.448 14.04 ; 
      RECT 37.532 9.666 37.636 14.04 ; 
      RECT 37.1 9.666 37.204 14.04 ; 
      RECT 36.668 9.666 36.772 14.04 ; 
      RECT 36.236 9.666 36.34 14.04 ; 
      RECT 35.804 9.666 35.908 14.04 ; 
      RECT 35.372 9.666 35.476 14.04 ; 
      RECT 34.94 9.666 35.044 14.04 ; 
      RECT 34.508 9.666 34.612 14.04 ; 
      RECT 34.076 9.666 34.18 14.04 ; 
      RECT 33.644 9.666 33.748 14.04 ; 
      RECT 33.212 9.666 33.316 14.04 ; 
      RECT 32.78 9.666 32.884 14.04 ; 
      RECT 32.348 9.666 32.452 14.04 ; 
      RECT 31.916 9.666 32.02 14.04 ; 
      RECT 31.484 9.666 31.588 14.04 ; 
      RECT 31.052 9.666 31.156 14.04 ; 
      RECT 30.62 9.666 30.724 14.04 ; 
      RECT 30.188 9.666 30.292 14.04 ; 
      RECT 29.756 9.666 29.86 14.04 ; 
      RECT 29.324 9.666 29.428 14.04 ; 
      RECT 28.892 9.666 28.996 14.04 ; 
      RECT 28.46 9.666 28.564 14.04 ; 
      RECT 28.028 9.666 28.132 14.04 ; 
      RECT 27.596 9.666 27.7 14.04 ; 
      RECT 27.164 9.666 27.268 14.04 ; 
      RECT 26.732 9.666 26.836 14.04 ; 
      RECT 26.3 9.666 26.404 14.04 ; 
      RECT 25.868 9.666 25.972 14.04 ; 
      RECT 25.436 9.666 25.54 14.04 ; 
      RECT 25.004 9.666 25.108 14.04 ; 
      RECT 24.572 9.666 24.676 14.04 ; 
      RECT 24.14 9.666 24.244 14.04 ; 
      RECT 23.708 9.666 23.812 14.04 ; 
      RECT 22.856 9.666 23.164 14.04 ; 
      RECT 15.284 9.666 15.592 14.04 ; 
      RECT 14.636 9.666 14.74 14.04 ; 
      RECT 14.204 9.666 14.308 14.04 ; 
      RECT 13.772 9.666 13.876 14.04 ; 
      RECT 13.34 9.666 13.444 14.04 ; 
      RECT 12.908 9.666 13.012 14.04 ; 
      RECT 12.476 9.666 12.58 14.04 ; 
      RECT 12.044 9.666 12.148 14.04 ; 
      RECT 11.612 9.666 11.716 14.04 ; 
      RECT 11.18 9.666 11.284 14.04 ; 
      RECT 10.748 9.666 10.852 14.04 ; 
      RECT 10.316 9.666 10.42 14.04 ; 
      RECT 9.884 9.666 9.988 14.04 ; 
      RECT 9.452 9.666 9.556 14.04 ; 
      RECT 9.02 9.666 9.124 14.04 ; 
      RECT 8.588 9.666 8.692 14.04 ; 
      RECT 8.156 9.666 8.26 14.04 ; 
      RECT 7.724 9.666 7.828 14.04 ; 
      RECT 7.292 9.666 7.396 14.04 ; 
      RECT 6.86 9.666 6.964 14.04 ; 
      RECT 6.428 9.666 6.532 14.04 ; 
      RECT 5.996 9.666 6.1 14.04 ; 
      RECT 5.564 9.666 5.668 14.04 ; 
      RECT 5.132 9.666 5.236 14.04 ; 
      RECT 4.7 9.666 4.804 14.04 ; 
      RECT 4.268 9.666 4.372 14.04 ; 
      RECT 3.836 9.666 3.94 14.04 ; 
      RECT 3.404 9.666 3.508 14.04 ; 
      RECT 2.972 9.666 3.076 14.04 ; 
      RECT 2.54 9.666 2.644 14.04 ; 
      RECT 2.108 9.666 2.212 14.04 ; 
      RECT 1.676 9.666 1.78 14.04 ; 
      RECT 1.244 9.666 1.348 14.04 ; 
      RECT 0.812 9.666 0.916 14.04 ; 
      RECT 0 9.666 0.34 14.04 ; 
      RECT 20.72 13.986 21.232 18.36 ; 
      RECT 20.664 16.648 21.232 17.938 ; 
      RECT 20.072 15.556 20.32 18.36 ; 
      RECT 20.016 16.794 20.32 17.408 ; 
      RECT 20.072 13.986 20.176 18.36 ; 
      RECT 20.072 14.47 20.232 15.428 ; 
      RECT 20.072 13.986 20.32 14.342 ; 
      RECT 18.884 15.788 19.708 18.36 ; 
      RECT 19.604 13.986 19.708 18.36 ; 
      RECT 18.884 16.896 19.764 17.928 ; 
      RECT 18.884 13.986 19.276 18.36 ; 
      RECT 17.216 13.986 17.548 18.36 ; 
      RECT 17.216 14.34 17.604 18.082 ; 
      RECT 38.108 13.986 38.448 18.36 ; 
      RECT 37.532 13.986 37.636 18.36 ; 
      RECT 37.1 13.986 37.204 18.36 ; 
      RECT 36.668 13.986 36.772 18.36 ; 
      RECT 36.236 13.986 36.34 18.36 ; 
      RECT 35.804 13.986 35.908 18.36 ; 
      RECT 35.372 13.986 35.476 18.36 ; 
      RECT 34.94 13.986 35.044 18.36 ; 
      RECT 34.508 13.986 34.612 18.36 ; 
      RECT 34.076 13.986 34.18 18.36 ; 
      RECT 33.644 13.986 33.748 18.36 ; 
      RECT 33.212 13.986 33.316 18.36 ; 
      RECT 32.78 13.986 32.884 18.36 ; 
      RECT 32.348 13.986 32.452 18.36 ; 
      RECT 31.916 13.986 32.02 18.36 ; 
      RECT 31.484 13.986 31.588 18.36 ; 
      RECT 31.052 13.986 31.156 18.36 ; 
      RECT 30.62 13.986 30.724 18.36 ; 
      RECT 30.188 13.986 30.292 18.36 ; 
      RECT 29.756 13.986 29.86 18.36 ; 
      RECT 29.324 13.986 29.428 18.36 ; 
      RECT 28.892 13.986 28.996 18.36 ; 
      RECT 28.46 13.986 28.564 18.36 ; 
      RECT 28.028 13.986 28.132 18.36 ; 
      RECT 27.596 13.986 27.7 18.36 ; 
      RECT 27.164 13.986 27.268 18.36 ; 
      RECT 26.732 13.986 26.836 18.36 ; 
      RECT 26.3 13.986 26.404 18.36 ; 
      RECT 25.868 13.986 25.972 18.36 ; 
      RECT 25.436 13.986 25.54 18.36 ; 
      RECT 25.004 13.986 25.108 18.36 ; 
      RECT 24.572 13.986 24.676 18.36 ; 
      RECT 24.14 13.986 24.244 18.36 ; 
      RECT 23.708 13.986 23.812 18.36 ; 
      RECT 22.856 13.986 23.164 18.36 ; 
      RECT 15.284 13.986 15.592 18.36 ; 
      RECT 14.636 13.986 14.74 18.36 ; 
      RECT 14.204 13.986 14.308 18.36 ; 
      RECT 13.772 13.986 13.876 18.36 ; 
      RECT 13.34 13.986 13.444 18.36 ; 
      RECT 12.908 13.986 13.012 18.36 ; 
      RECT 12.476 13.986 12.58 18.36 ; 
      RECT 12.044 13.986 12.148 18.36 ; 
      RECT 11.612 13.986 11.716 18.36 ; 
      RECT 11.18 13.986 11.284 18.36 ; 
      RECT 10.748 13.986 10.852 18.36 ; 
      RECT 10.316 13.986 10.42 18.36 ; 
      RECT 9.884 13.986 9.988 18.36 ; 
      RECT 9.452 13.986 9.556 18.36 ; 
      RECT 9.02 13.986 9.124 18.36 ; 
      RECT 8.588 13.986 8.692 18.36 ; 
      RECT 8.156 13.986 8.26 18.36 ; 
      RECT 7.724 13.986 7.828 18.36 ; 
      RECT 7.292 13.986 7.396 18.36 ; 
      RECT 6.86 13.986 6.964 18.36 ; 
      RECT 6.428 13.986 6.532 18.36 ; 
      RECT 5.996 13.986 6.1 18.36 ; 
      RECT 5.564 13.986 5.668 18.36 ; 
      RECT 5.132 13.986 5.236 18.36 ; 
      RECT 4.7 13.986 4.804 18.36 ; 
      RECT 4.268 13.986 4.372 18.36 ; 
      RECT 3.836 13.986 3.94 18.36 ; 
      RECT 3.404 13.986 3.508 18.36 ; 
      RECT 2.972 13.986 3.076 18.36 ; 
      RECT 2.54 13.986 2.644 18.36 ; 
      RECT 2.108 13.986 2.212 18.36 ; 
      RECT 1.676 13.986 1.78 18.36 ; 
      RECT 1.244 13.986 1.348 18.36 ; 
      RECT 0.812 13.986 0.916 18.36 ; 
      RECT 0 13.986 0.34 18.36 ; 
      RECT 20.72 18.306 21.232 22.68 ; 
      RECT 20.664 20.968 21.232 22.258 ; 
      RECT 20.072 19.876 20.32 22.68 ; 
      RECT 20.016 21.114 20.32 21.728 ; 
      RECT 20.072 18.306 20.176 22.68 ; 
      RECT 20.072 18.79 20.232 19.748 ; 
      RECT 20.072 18.306 20.32 18.662 ; 
      RECT 18.884 20.108 19.708 22.68 ; 
      RECT 19.604 18.306 19.708 22.68 ; 
      RECT 18.884 21.216 19.764 22.248 ; 
      RECT 18.884 18.306 19.276 22.68 ; 
      RECT 17.216 18.306 17.548 22.68 ; 
      RECT 17.216 18.66 17.604 22.402 ; 
      RECT 38.108 18.306 38.448 22.68 ; 
      RECT 37.532 18.306 37.636 22.68 ; 
      RECT 37.1 18.306 37.204 22.68 ; 
      RECT 36.668 18.306 36.772 22.68 ; 
      RECT 36.236 18.306 36.34 22.68 ; 
      RECT 35.804 18.306 35.908 22.68 ; 
      RECT 35.372 18.306 35.476 22.68 ; 
      RECT 34.94 18.306 35.044 22.68 ; 
      RECT 34.508 18.306 34.612 22.68 ; 
      RECT 34.076 18.306 34.18 22.68 ; 
      RECT 33.644 18.306 33.748 22.68 ; 
      RECT 33.212 18.306 33.316 22.68 ; 
      RECT 32.78 18.306 32.884 22.68 ; 
      RECT 32.348 18.306 32.452 22.68 ; 
      RECT 31.916 18.306 32.02 22.68 ; 
      RECT 31.484 18.306 31.588 22.68 ; 
      RECT 31.052 18.306 31.156 22.68 ; 
      RECT 30.62 18.306 30.724 22.68 ; 
      RECT 30.188 18.306 30.292 22.68 ; 
      RECT 29.756 18.306 29.86 22.68 ; 
      RECT 29.324 18.306 29.428 22.68 ; 
      RECT 28.892 18.306 28.996 22.68 ; 
      RECT 28.46 18.306 28.564 22.68 ; 
      RECT 28.028 18.306 28.132 22.68 ; 
      RECT 27.596 18.306 27.7 22.68 ; 
      RECT 27.164 18.306 27.268 22.68 ; 
      RECT 26.732 18.306 26.836 22.68 ; 
      RECT 26.3 18.306 26.404 22.68 ; 
      RECT 25.868 18.306 25.972 22.68 ; 
      RECT 25.436 18.306 25.54 22.68 ; 
      RECT 25.004 18.306 25.108 22.68 ; 
      RECT 24.572 18.306 24.676 22.68 ; 
      RECT 24.14 18.306 24.244 22.68 ; 
      RECT 23.708 18.306 23.812 22.68 ; 
      RECT 22.856 18.306 23.164 22.68 ; 
      RECT 15.284 18.306 15.592 22.68 ; 
      RECT 14.636 18.306 14.74 22.68 ; 
      RECT 14.204 18.306 14.308 22.68 ; 
      RECT 13.772 18.306 13.876 22.68 ; 
      RECT 13.34 18.306 13.444 22.68 ; 
      RECT 12.908 18.306 13.012 22.68 ; 
      RECT 12.476 18.306 12.58 22.68 ; 
      RECT 12.044 18.306 12.148 22.68 ; 
      RECT 11.612 18.306 11.716 22.68 ; 
      RECT 11.18 18.306 11.284 22.68 ; 
      RECT 10.748 18.306 10.852 22.68 ; 
      RECT 10.316 18.306 10.42 22.68 ; 
      RECT 9.884 18.306 9.988 22.68 ; 
      RECT 9.452 18.306 9.556 22.68 ; 
      RECT 9.02 18.306 9.124 22.68 ; 
      RECT 8.588 18.306 8.692 22.68 ; 
      RECT 8.156 18.306 8.26 22.68 ; 
      RECT 7.724 18.306 7.828 22.68 ; 
      RECT 7.292 18.306 7.396 22.68 ; 
      RECT 6.86 18.306 6.964 22.68 ; 
      RECT 6.428 18.306 6.532 22.68 ; 
      RECT 5.996 18.306 6.1 22.68 ; 
      RECT 5.564 18.306 5.668 22.68 ; 
      RECT 5.132 18.306 5.236 22.68 ; 
      RECT 4.7 18.306 4.804 22.68 ; 
      RECT 4.268 18.306 4.372 22.68 ; 
      RECT 3.836 18.306 3.94 22.68 ; 
      RECT 3.404 18.306 3.508 22.68 ; 
      RECT 2.972 18.306 3.076 22.68 ; 
      RECT 2.54 18.306 2.644 22.68 ; 
      RECT 2.108 18.306 2.212 22.68 ; 
      RECT 1.676 18.306 1.78 22.68 ; 
      RECT 1.244 18.306 1.348 22.68 ; 
      RECT 0.812 18.306 0.916 22.68 ; 
      RECT 0 18.306 0.34 22.68 ; 
      RECT 20.72 22.626 21.232 27 ; 
      RECT 20.664 25.288 21.232 26.578 ; 
      RECT 20.072 24.196 20.32 27 ; 
      RECT 20.016 25.434 20.32 26.048 ; 
      RECT 20.072 22.626 20.176 27 ; 
      RECT 20.072 23.11 20.232 24.068 ; 
      RECT 20.072 22.626 20.32 22.982 ; 
      RECT 18.884 24.428 19.708 27 ; 
      RECT 19.604 22.626 19.708 27 ; 
      RECT 18.884 25.536 19.764 26.568 ; 
      RECT 18.884 22.626 19.276 27 ; 
      RECT 17.216 22.626 17.548 27 ; 
      RECT 17.216 22.98 17.604 26.722 ; 
      RECT 38.108 22.626 38.448 27 ; 
      RECT 37.532 22.626 37.636 27 ; 
      RECT 37.1 22.626 37.204 27 ; 
      RECT 36.668 22.626 36.772 27 ; 
      RECT 36.236 22.626 36.34 27 ; 
      RECT 35.804 22.626 35.908 27 ; 
      RECT 35.372 22.626 35.476 27 ; 
      RECT 34.94 22.626 35.044 27 ; 
      RECT 34.508 22.626 34.612 27 ; 
      RECT 34.076 22.626 34.18 27 ; 
      RECT 33.644 22.626 33.748 27 ; 
      RECT 33.212 22.626 33.316 27 ; 
      RECT 32.78 22.626 32.884 27 ; 
      RECT 32.348 22.626 32.452 27 ; 
      RECT 31.916 22.626 32.02 27 ; 
      RECT 31.484 22.626 31.588 27 ; 
      RECT 31.052 22.626 31.156 27 ; 
      RECT 30.62 22.626 30.724 27 ; 
      RECT 30.188 22.626 30.292 27 ; 
      RECT 29.756 22.626 29.86 27 ; 
      RECT 29.324 22.626 29.428 27 ; 
      RECT 28.892 22.626 28.996 27 ; 
      RECT 28.46 22.626 28.564 27 ; 
      RECT 28.028 22.626 28.132 27 ; 
      RECT 27.596 22.626 27.7 27 ; 
      RECT 27.164 22.626 27.268 27 ; 
      RECT 26.732 22.626 26.836 27 ; 
      RECT 26.3 22.626 26.404 27 ; 
      RECT 25.868 22.626 25.972 27 ; 
      RECT 25.436 22.626 25.54 27 ; 
      RECT 25.004 22.626 25.108 27 ; 
      RECT 24.572 22.626 24.676 27 ; 
      RECT 24.14 22.626 24.244 27 ; 
      RECT 23.708 22.626 23.812 27 ; 
      RECT 22.856 22.626 23.164 27 ; 
      RECT 15.284 22.626 15.592 27 ; 
      RECT 14.636 22.626 14.74 27 ; 
      RECT 14.204 22.626 14.308 27 ; 
      RECT 13.772 22.626 13.876 27 ; 
      RECT 13.34 22.626 13.444 27 ; 
      RECT 12.908 22.626 13.012 27 ; 
      RECT 12.476 22.626 12.58 27 ; 
      RECT 12.044 22.626 12.148 27 ; 
      RECT 11.612 22.626 11.716 27 ; 
      RECT 11.18 22.626 11.284 27 ; 
      RECT 10.748 22.626 10.852 27 ; 
      RECT 10.316 22.626 10.42 27 ; 
      RECT 9.884 22.626 9.988 27 ; 
      RECT 9.452 22.626 9.556 27 ; 
      RECT 9.02 22.626 9.124 27 ; 
      RECT 8.588 22.626 8.692 27 ; 
      RECT 8.156 22.626 8.26 27 ; 
      RECT 7.724 22.626 7.828 27 ; 
      RECT 7.292 22.626 7.396 27 ; 
      RECT 6.86 22.626 6.964 27 ; 
      RECT 6.428 22.626 6.532 27 ; 
      RECT 5.996 22.626 6.1 27 ; 
      RECT 5.564 22.626 5.668 27 ; 
      RECT 5.132 22.626 5.236 27 ; 
      RECT 4.7 22.626 4.804 27 ; 
      RECT 4.268 22.626 4.372 27 ; 
      RECT 3.836 22.626 3.94 27 ; 
      RECT 3.404 22.626 3.508 27 ; 
      RECT 2.972 22.626 3.076 27 ; 
      RECT 2.54 22.626 2.644 27 ; 
      RECT 2.108 22.626 2.212 27 ; 
      RECT 1.676 22.626 1.78 27 ; 
      RECT 1.244 22.626 1.348 27 ; 
      RECT 0.812 22.626 0.916 27 ; 
      RECT 0 22.626 0.34 27 ; 
      RECT 20.72 26.946 21.232 31.32 ; 
      RECT 20.664 29.608 21.232 30.898 ; 
      RECT 20.072 28.516 20.32 31.32 ; 
      RECT 20.016 29.754 20.32 30.368 ; 
      RECT 20.072 26.946 20.176 31.32 ; 
      RECT 20.072 27.43 20.232 28.388 ; 
      RECT 20.072 26.946 20.32 27.302 ; 
      RECT 18.884 28.748 19.708 31.32 ; 
      RECT 19.604 26.946 19.708 31.32 ; 
      RECT 18.884 29.856 19.764 30.888 ; 
      RECT 18.884 26.946 19.276 31.32 ; 
      RECT 17.216 26.946 17.548 31.32 ; 
      RECT 17.216 27.3 17.604 31.042 ; 
      RECT 38.108 26.946 38.448 31.32 ; 
      RECT 37.532 26.946 37.636 31.32 ; 
      RECT 37.1 26.946 37.204 31.32 ; 
      RECT 36.668 26.946 36.772 31.32 ; 
      RECT 36.236 26.946 36.34 31.32 ; 
      RECT 35.804 26.946 35.908 31.32 ; 
      RECT 35.372 26.946 35.476 31.32 ; 
      RECT 34.94 26.946 35.044 31.32 ; 
      RECT 34.508 26.946 34.612 31.32 ; 
      RECT 34.076 26.946 34.18 31.32 ; 
      RECT 33.644 26.946 33.748 31.32 ; 
      RECT 33.212 26.946 33.316 31.32 ; 
      RECT 32.78 26.946 32.884 31.32 ; 
      RECT 32.348 26.946 32.452 31.32 ; 
      RECT 31.916 26.946 32.02 31.32 ; 
      RECT 31.484 26.946 31.588 31.32 ; 
      RECT 31.052 26.946 31.156 31.32 ; 
      RECT 30.62 26.946 30.724 31.32 ; 
      RECT 30.188 26.946 30.292 31.32 ; 
      RECT 29.756 26.946 29.86 31.32 ; 
      RECT 29.324 26.946 29.428 31.32 ; 
      RECT 28.892 26.946 28.996 31.32 ; 
      RECT 28.46 26.946 28.564 31.32 ; 
      RECT 28.028 26.946 28.132 31.32 ; 
      RECT 27.596 26.946 27.7 31.32 ; 
      RECT 27.164 26.946 27.268 31.32 ; 
      RECT 26.732 26.946 26.836 31.32 ; 
      RECT 26.3 26.946 26.404 31.32 ; 
      RECT 25.868 26.946 25.972 31.32 ; 
      RECT 25.436 26.946 25.54 31.32 ; 
      RECT 25.004 26.946 25.108 31.32 ; 
      RECT 24.572 26.946 24.676 31.32 ; 
      RECT 24.14 26.946 24.244 31.32 ; 
      RECT 23.708 26.946 23.812 31.32 ; 
      RECT 22.856 26.946 23.164 31.32 ; 
      RECT 15.284 26.946 15.592 31.32 ; 
      RECT 14.636 26.946 14.74 31.32 ; 
      RECT 14.204 26.946 14.308 31.32 ; 
      RECT 13.772 26.946 13.876 31.32 ; 
      RECT 13.34 26.946 13.444 31.32 ; 
      RECT 12.908 26.946 13.012 31.32 ; 
      RECT 12.476 26.946 12.58 31.32 ; 
      RECT 12.044 26.946 12.148 31.32 ; 
      RECT 11.612 26.946 11.716 31.32 ; 
      RECT 11.18 26.946 11.284 31.32 ; 
      RECT 10.748 26.946 10.852 31.32 ; 
      RECT 10.316 26.946 10.42 31.32 ; 
      RECT 9.884 26.946 9.988 31.32 ; 
      RECT 9.452 26.946 9.556 31.32 ; 
      RECT 9.02 26.946 9.124 31.32 ; 
      RECT 8.588 26.946 8.692 31.32 ; 
      RECT 8.156 26.946 8.26 31.32 ; 
      RECT 7.724 26.946 7.828 31.32 ; 
      RECT 7.292 26.946 7.396 31.32 ; 
      RECT 6.86 26.946 6.964 31.32 ; 
      RECT 6.428 26.946 6.532 31.32 ; 
      RECT 5.996 26.946 6.1 31.32 ; 
      RECT 5.564 26.946 5.668 31.32 ; 
      RECT 5.132 26.946 5.236 31.32 ; 
      RECT 4.7 26.946 4.804 31.32 ; 
      RECT 4.268 26.946 4.372 31.32 ; 
      RECT 3.836 26.946 3.94 31.32 ; 
      RECT 3.404 26.946 3.508 31.32 ; 
      RECT 2.972 26.946 3.076 31.32 ; 
      RECT 2.54 26.946 2.644 31.32 ; 
      RECT 2.108 26.946 2.212 31.32 ; 
      RECT 1.676 26.946 1.78 31.32 ; 
      RECT 1.244 26.946 1.348 31.32 ; 
      RECT 0.812 26.946 0.916 31.32 ; 
      RECT 0 26.946 0.34 31.32 ; 
      RECT 20.72 31.266 21.232 35.64 ; 
      RECT 20.664 33.928 21.232 35.218 ; 
      RECT 20.072 32.836 20.32 35.64 ; 
      RECT 20.016 34.074 20.32 34.688 ; 
      RECT 20.072 31.266 20.176 35.64 ; 
      RECT 20.072 31.75 20.232 32.708 ; 
      RECT 20.072 31.266 20.32 31.622 ; 
      RECT 18.884 33.068 19.708 35.64 ; 
      RECT 19.604 31.266 19.708 35.64 ; 
      RECT 18.884 34.176 19.764 35.208 ; 
      RECT 18.884 31.266 19.276 35.64 ; 
      RECT 17.216 31.266 17.548 35.64 ; 
      RECT 17.216 31.62 17.604 35.362 ; 
      RECT 38.108 31.266 38.448 35.64 ; 
      RECT 37.532 31.266 37.636 35.64 ; 
      RECT 37.1 31.266 37.204 35.64 ; 
      RECT 36.668 31.266 36.772 35.64 ; 
      RECT 36.236 31.266 36.34 35.64 ; 
      RECT 35.804 31.266 35.908 35.64 ; 
      RECT 35.372 31.266 35.476 35.64 ; 
      RECT 34.94 31.266 35.044 35.64 ; 
      RECT 34.508 31.266 34.612 35.64 ; 
      RECT 34.076 31.266 34.18 35.64 ; 
      RECT 33.644 31.266 33.748 35.64 ; 
      RECT 33.212 31.266 33.316 35.64 ; 
      RECT 32.78 31.266 32.884 35.64 ; 
      RECT 32.348 31.266 32.452 35.64 ; 
      RECT 31.916 31.266 32.02 35.64 ; 
      RECT 31.484 31.266 31.588 35.64 ; 
      RECT 31.052 31.266 31.156 35.64 ; 
      RECT 30.62 31.266 30.724 35.64 ; 
      RECT 30.188 31.266 30.292 35.64 ; 
      RECT 29.756 31.266 29.86 35.64 ; 
      RECT 29.324 31.266 29.428 35.64 ; 
      RECT 28.892 31.266 28.996 35.64 ; 
      RECT 28.46 31.266 28.564 35.64 ; 
      RECT 28.028 31.266 28.132 35.64 ; 
      RECT 27.596 31.266 27.7 35.64 ; 
      RECT 27.164 31.266 27.268 35.64 ; 
      RECT 26.732 31.266 26.836 35.64 ; 
      RECT 26.3 31.266 26.404 35.64 ; 
      RECT 25.868 31.266 25.972 35.64 ; 
      RECT 25.436 31.266 25.54 35.64 ; 
      RECT 25.004 31.266 25.108 35.64 ; 
      RECT 24.572 31.266 24.676 35.64 ; 
      RECT 24.14 31.266 24.244 35.64 ; 
      RECT 23.708 31.266 23.812 35.64 ; 
      RECT 22.856 31.266 23.164 35.64 ; 
      RECT 15.284 31.266 15.592 35.64 ; 
      RECT 14.636 31.266 14.74 35.64 ; 
      RECT 14.204 31.266 14.308 35.64 ; 
      RECT 13.772 31.266 13.876 35.64 ; 
      RECT 13.34 31.266 13.444 35.64 ; 
      RECT 12.908 31.266 13.012 35.64 ; 
      RECT 12.476 31.266 12.58 35.64 ; 
      RECT 12.044 31.266 12.148 35.64 ; 
      RECT 11.612 31.266 11.716 35.64 ; 
      RECT 11.18 31.266 11.284 35.64 ; 
      RECT 10.748 31.266 10.852 35.64 ; 
      RECT 10.316 31.266 10.42 35.64 ; 
      RECT 9.884 31.266 9.988 35.64 ; 
      RECT 9.452 31.266 9.556 35.64 ; 
      RECT 9.02 31.266 9.124 35.64 ; 
      RECT 8.588 31.266 8.692 35.64 ; 
      RECT 8.156 31.266 8.26 35.64 ; 
      RECT 7.724 31.266 7.828 35.64 ; 
      RECT 7.292 31.266 7.396 35.64 ; 
      RECT 6.86 31.266 6.964 35.64 ; 
      RECT 6.428 31.266 6.532 35.64 ; 
      RECT 5.996 31.266 6.1 35.64 ; 
      RECT 5.564 31.266 5.668 35.64 ; 
      RECT 5.132 31.266 5.236 35.64 ; 
      RECT 4.7 31.266 4.804 35.64 ; 
      RECT 4.268 31.266 4.372 35.64 ; 
      RECT 3.836 31.266 3.94 35.64 ; 
      RECT 3.404 31.266 3.508 35.64 ; 
      RECT 2.972 31.266 3.076 35.64 ; 
      RECT 2.54 31.266 2.644 35.64 ; 
      RECT 2.108 31.266 2.212 35.64 ; 
      RECT 1.676 31.266 1.78 35.64 ; 
      RECT 1.244 31.266 1.348 35.64 ; 
      RECT 0.812 31.266 0.916 35.64 ; 
      RECT 0 31.266 0.34 35.64 ; 
      RECT 20.72 35.586 21.232 39.96 ; 
      RECT 20.664 38.248 21.232 39.538 ; 
      RECT 20.072 37.156 20.32 39.96 ; 
      RECT 20.016 38.394 20.32 39.008 ; 
      RECT 20.072 35.586 20.176 39.96 ; 
      RECT 20.072 36.07 20.232 37.028 ; 
      RECT 20.072 35.586 20.32 35.942 ; 
      RECT 18.884 37.388 19.708 39.96 ; 
      RECT 19.604 35.586 19.708 39.96 ; 
      RECT 18.884 38.496 19.764 39.528 ; 
      RECT 18.884 35.586 19.276 39.96 ; 
      RECT 17.216 35.586 17.548 39.96 ; 
      RECT 17.216 35.94 17.604 39.682 ; 
      RECT 38.108 35.586 38.448 39.96 ; 
      RECT 37.532 35.586 37.636 39.96 ; 
      RECT 37.1 35.586 37.204 39.96 ; 
      RECT 36.668 35.586 36.772 39.96 ; 
      RECT 36.236 35.586 36.34 39.96 ; 
      RECT 35.804 35.586 35.908 39.96 ; 
      RECT 35.372 35.586 35.476 39.96 ; 
      RECT 34.94 35.586 35.044 39.96 ; 
      RECT 34.508 35.586 34.612 39.96 ; 
      RECT 34.076 35.586 34.18 39.96 ; 
      RECT 33.644 35.586 33.748 39.96 ; 
      RECT 33.212 35.586 33.316 39.96 ; 
      RECT 32.78 35.586 32.884 39.96 ; 
      RECT 32.348 35.586 32.452 39.96 ; 
      RECT 31.916 35.586 32.02 39.96 ; 
      RECT 31.484 35.586 31.588 39.96 ; 
      RECT 31.052 35.586 31.156 39.96 ; 
      RECT 30.62 35.586 30.724 39.96 ; 
      RECT 30.188 35.586 30.292 39.96 ; 
      RECT 29.756 35.586 29.86 39.96 ; 
      RECT 29.324 35.586 29.428 39.96 ; 
      RECT 28.892 35.586 28.996 39.96 ; 
      RECT 28.46 35.586 28.564 39.96 ; 
      RECT 28.028 35.586 28.132 39.96 ; 
      RECT 27.596 35.586 27.7 39.96 ; 
      RECT 27.164 35.586 27.268 39.96 ; 
      RECT 26.732 35.586 26.836 39.96 ; 
      RECT 26.3 35.586 26.404 39.96 ; 
      RECT 25.868 35.586 25.972 39.96 ; 
      RECT 25.436 35.586 25.54 39.96 ; 
      RECT 25.004 35.586 25.108 39.96 ; 
      RECT 24.572 35.586 24.676 39.96 ; 
      RECT 24.14 35.586 24.244 39.96 ; 
      RECT 23.708 35.586 23.812 39.96 ; 
      RECT 22.856 35.586 23.164 39.96 ; 
      RECT 15.284 35.586 15.592 39.96 ; 
      RECT 14.636 35.586 14.74 39.96 ; 
      RECT 14.204 35.586 14.308 39.96 ; 
      RECT 13.772 35.586 13.876 39.96 ; 
      RECT 13.34 35.586 13.444 39.96 ; 
      RECT 12.908 35.586 13.012 39.96 ; 
      RECT 12.476 35.586 12.58 39.96 ; 
      RECT 12.044 35.586 12.148 39.96 ; 
      RECT 11.612 35.586 11.716 39.96 ; 
      RECT 11.18 35.586 11.284 39.96 ; 
      RECT 10.748 35.586 10.852 39.96 ; 
      RECT 10.316 35.586 10.42 39.96 ; 
      RECT 9.884 35.586 9.988 39.96 ; 
      RECT 9.452 35.586 9.556 39.96 ; 
      RECT 9.02 35.586 9.124 39.96 ; 
      RECT 8.588 35.586 8.692 39.96 ; 
      RECT 8.156 35.586 8.26 39.96 ; 
      RECT 7.724 35.586 7.828 39.96 ; 
      RECT 7.292 35.586 7.396 39.96 ; 
      RECT 6.86 35.586 6.964 39.96 ; 
      RECT 6.428 35.586 6.532 39.96 ; 
      RECT 5.996 35.586 6.1 39.96 ; 
      RECT 5.564 35.586 5.668 39.96 ; 
      RECT 5.132 35.586 5.236 39.96 ; 
      RECT 4.7 35.586 4.804 39.96 ; 
      RECT 4.268 35.586 4.372 39.96 ; 
      RECT 3.836 35.586 3.94 39.96 ; 
      RECT 3.404 35.586 3.508 39.96 ; 
      RECT 2.972 35.586 3.076 39.96 ; 
      RECT 2.54 35.586 2.644 39.96 ; 
      RECT 2.108 35.586 2.212 39.96 ; 
      RECT 1.676 35.586 1.78 39.96 ; 
      RECT 1.244 35.586 1.348 39.96 ; 
      RECT 0.812 35.586 0.916 39.96 ; 
      RECT 0 35.586 0.34 39.96 ; 
      RECT 20.72 39.906 21.232 44.28 ; 
      RECT 20.664 42.568 21.232 43.858 ; 
      RECT 20.072 41.476 20.32 44.28 ; 
      RECT 20.016 42.714 20.32 43.328 ; 
      RECT 20.072 39.906 20.176 44.28 ; 
      RECT 20.072 40.39 20.232 41.348 ; 
      RECT 20.072 39.906 20.32 40.262 ; 
      RECT 18.884 41.708 19.708 44.28 ; 
      RECT 19.604 39.906 19.708 44.28 ; 
      RECT 18.884 42.816 19.764 43.848 ; 
      RECT 18.884 39.906 19.276 44.28 ; 
      RECT 17.216 39.906 17.548 44.28 ; 
      RECT 17.216 40.26 17.604 44.002 ; 
      RECT 38.108 39.906 38.448 44.28 ; 
      RECT 37.532 39.906 37.636 44.28 ; 
      RECT 37.1 39.906 37.204 44.28 ; 
      RECT 36.668 39.906 36.772 44.28 ; 
      RECT 36.236 39.906 36.34 44.28 ; 
      RECT 35.804 39.906 35.908 44.28 ; 
      RECT 35.372 39.906 35.476 44.28 ; 
      RECT 34.94 39.906 35.044 44.28 ; 
      RECT 34.508 39.906 34.612 44.28 ; 
      RECT 34.076 39.906 34.18 44.28 ; 
      RECT 33.644 39.906 33.748 44.28 ; 
      RECT 33.212 39.906 33.316 44.28 ; 
      RECT 32.78 39.906 32.884 44.28 ; 
      RECT 32.348 39.906 32.452 44.28 ; 
      RECT 31.916 39.906 32.02 44.28 ; 
      RECT 31.484 39.906 31.588 44.28 ; 
      RECT 31.052 39.906 31.156 44.28 ; 
      RECT 30.62 39.906 30.724 44.28 ; 
      RECT 30.188 39.906 30.292 44.28 ; 
      RECT 29.756 39.906 29.86 44.28 ; 
      RECT 29.324 39.906 29.428 44.28 ; 
      RECT 28.892 39.906 28.996 44.28 ; 
      RECT 28.46 39.906 28.564 44.28 ; 
      RECT 28.028 39.906 28.132 44.28 ; 
      RECT 27.596 39.906 27.7 44.28 ; 
      RECT 27.164 39.906 27.268 44.28 ; 
      RECT 26.732 39.906 26.836 44.28 ; 
      RECT 26.3 39.906 26.404 44.28 ; 
      RECT 25.868 39.906 25.972 44.28 ; 
      RECT 25.436 39.906 25.54 44.28 ; 
      RECT 25.004 39.906 25.108 44.28 ; 
      RECT 24.572 39.906 24.676 44.28 ; 
      RECT 24.14 39.906 24.244 44.28 ; 
      RECT 23.708 39.906 23.812 44.28 ; 
      RECT 22.856 39.906 23.164 44.28 ; 
      RECT 15.284 39.906 15.592 44.28 ; 
      RECT 14.636 39.906 14.74 44.28 ; 
      RECT 14.204 39.906 14.308 44.28 ; 
      RECT 13.772 39.906 13.876 44.28 ; 
      RECT 13.34 39.906 13.444 44.28 ; 
      RECT 12.908 39.906 13.012 44.28 ; 
      RECT 12.476 39.906 12.58 44.28 ; 
      RECT 12.044 39.906 12.148 44.28 ; 
      RECT 11.612 39.906 11.716 44.28 ; 
      RECT 11.18 39.906 11.284 44.28 ; 
      RECT 10.748 39.906 10.852 44.28 ; 
      RECT 10.316 39.906 10.42 44.28 ; 
      RECT 9.884 39.906 9.988 44.28 ; 
      RECT 9.452 39.906 9.556 44.28 ; 
      RECT 9.02 39.906 9.124 44.28 ; 
      RECT 8.588 39.906 8.692 44.28 ; 
      RECT 8.156 39.906 8.26 44.28 ; 
      RECT 7.724 39.906 7.828 44.28 ; 
      RECT 7.292 39.906 7.396 44.28 ; 
      RECT 6.86 39.906 6.964 44.28 ; 
      RECT 6.428 39.906 6.532 44.28 ; 
      RECT 5.996 39.906 6.1 44.28 ; 
      RECT 5.564 39.906 5.668 44.28 ; 
      RECT 5.132 39.906 5.236 44.28 ; 
      RECT 4.7 39.906 4.804 44.28 ; 
      RECT 4.268 39.906 4.372 44.28 ; 
      RECT 3.836 39.906 3.94 44.28 ; 
      RECT 3.404 39.906 3.508 44.28 ; 
      RECT 2.972 39.906 3.076 44.28 ; 
      RECT 2.54 39.906 2.644 44.28 ; 
      RECT 2.108 39.906 2.212 44.28 ; 
      RECT 1.676 39.906 1.78 44.28 ; 
      RECT 1.244 39.906 1.348 44.28 ; 
      RECT 0.812 39.906 0.916 44.28 ; 
      RECT 0 39.906 0.34 44.28 ; 
      RECT 20.72 44.226 21.232 48.6 ; 
      RECT 20.664 46.888 21.232 48.178 ; 
      RECT 20.072 45.796 20.32 48.6 ; 
      RECT 20.016 47.034 20.32 47.648 ; 
      RECT 20.072 44.226 20.176 48.6 ; 
      RECT 20.072 44.71 20.232 45.668 ; 
      RECT 20.072 44.226 20.32 44.582 ; 
      RECT 18.884 46.028 19.708 48.6 ; 
      RECT 19.604 44.226 19.708 48.6 ; 
      RECT 18.884 47.136 19.764 48.168 ; 
      RECT 18.884 44.226 19.276 48.6 ; 
      RECT 17.216 44.226 17.548 48.6 ; 
      RECT 17.216 44.58 17.604 48.322 ; 
      RECT 38.108 44.226 38.448 48.6 ; 
      RECT 37.532 44.226 37.636 48.6 ; 
      RECT 37.1 44.226 37.204 48.6 ; 
      RECT 36.668 44.226 36.772 48.6 ; 
      RECT 36.236 44.226 36.34 48.6 ; 
      RECT 35.804 44.226 35.908 48.6 ; 
      RECT 35.372 44.226 35.476 48.6 ; 
      RECT 34.94 44.226 35.044 48.6 ; 
      RECT 34.508 44.226 34.612 48.6 ; 
      RECT 34.076 44.226 34.18 48.6 ; 
      RECT 33.644 44.226 33.748 48.6 ; 
      RECT 33.212 44.226 33.316 48.6 ; 
      RECT 32.78 44.226 32.884 48.6 ; 
      RECT 32.348 44.226 32.452 48.6 ; 
      RECT 31.916 44.226 32.02 48.6 ; 
      RECT 31.484 44.226 31.588 48.6 ; 
      RECT 31.052 44.226 31.156 48.6 ; 
      RECT 30.62 44.226 30.724 48.6 ; 
      RECT 30.188 44.226 30.292 48.6 ; 
      RECT 29.756 44.226 29.86 48.6 ; 
      RECT 29.324 44.226 29.428 48.6 ; 
      RECT 28.892 44.226 28.996 48.6 ; 
      RECT 28.46 44.226 28.564 48.6 ; 
      RECT 28.028 44.226 28.132 48.6 ; 
      RECT 27.596 44.226 27.7 48.6 ; 
      RECT 27.164 44.226 27.268 48.6 ; 
      RECT 26.732 44.226 26.836 48.6 ; 
      RECT 26.3 44.226 26.404 48.6 ; 
      RECT 25.868 44.226 25.972 48.6 ; 
      RECT 25.436 44.226 25.54 48.6 ; 
      RECT 25.004 44.226 25.108 48.6 ; 
      RECT 24.572 44.226 24.676 48.6 ; 
      RECT 24.14 44.226 24.244 48.6 ; 
      RECT 23.708 44.226 23.812 48.6 ; 
      RECT 22.856 44.226 23.164 48.6 ; 
      RECT 15.284 44.226 15.592 48.6 ; 
      RECT 14.636 44.226 14.74 48.6 ; 
      RECT 14.204 44.226 14.308 48.6 ; 
      RECT 13.772 44.226 13.876 48.6 ; 
      RECT 13.34 44.226 13.444 48.6 ; 
      RECT 12.908 44.226 13.012 48.6 ; 
      RECT 12.476 44.226 12.58 48.6 ; 
      RECT 12.044 44.226 12.148 48.6 ; 
      RECT 11.612 44.226 11.716 48.6 ; 
      RECT 11.18 44.226 11.284 48.6 ; 
      RECT 10.748 44.226 10.852 48.6 ; 
      RECT 10.316 44.226 10.42 48.6 ; 
      RECT 9.884 44.226 9.988 48.6 ; 
      RECT 9.452 44.226 9.556 48.6 ; 
      RECT 9.02 44.226 9.124 48.6 ; 
      RECT 8.588 44.226 8.692 48.6 ; 
      RECT 8.156 44.226 8.26 48.6 ; 
      RECT 7.724 44.226 7.828 48.6 ; 
      RECT 7.292 44.226 7.396 48.6 ; 
      RECT 6.86 44.226 6.964 48.6 ; 
      RECT 6.428 44.226 6.532 48.6 ; 
      RECT 5.996 44.226 6.1 48.6 ; 
      RECT 5.564 44.226 5.668 48.6 ; 
      RECT 5.132 44.226 5.236 48.6 ; 
      RECT 4.7 44.226 4.804 48.6 ; 
      RECT 4.268 44.226 4.372 48.6 ; 
      RECT 3.836 44.226 3.94 48.6 ; 
      RECT 3.404 44.226 3.508 48.6 ; 
      RECT 2.972 44.226 3.076 48.6 ; 
      RECT 2.54 44.226 2.644 48.6 ; 
      RECT 2.108 44.226 2.212 48.6 ; 
      RECT 1.676 44.226 1.78 48.6 ; 
      RECT 1.244 44.226 1.348 48.6 ; 
      RECT 0.812 44.226 0.916 48.6 ; 
      RECT 0 44.226 0.34 48.6 ; 
      RECT 20.72 48.546 21.232 52.92 ; 
      RECT 20.664 51.208 21.232 52.498 ; 
      RECT 20.072 50.116 20.32 52.92 ; 
      RECT 20.016 51.354 20.32 51.968 ; 
      RECT 20.072 48.546 20.176 52.92 ; 
      RECT 20.072 49.03 20.232 49.988 ; 
      RECT 20.072 48.546 20.32 48.902 ; 
      RECT 18.884 50.348 19.708 52.92 ; 
      RECT 19.604 48.546 19.708 52.92 ; 
      RECT 18.884 51.456 19.764 52.488 ; 
      RECT 18.884 48.546 19.276 52.92 ; 
      RECT 17.216 48.546 17.548 52.92 ; 
      RECT 17.216 48.9 17.604 52.642 ; 
      RECT 38.108 48.546 38.448 52.92 ; 
      RECT 37.532 48.546 37.636 52.92 ; 
      RECT 37.1 48.546 37.204 52.92 ; 
      RECT 36.668 48.546 36.772 52.92 ; 
      RECT 36.236 48.546 36.34 52.92 ; 
      RECT 35.804 48.546 35.908 52.92 ; 
      RECT 35.372 48.546 35.476 52.92 ; 
      RECT 34.94 48.546 35.044 52.92 ; 
      RECT 34.508 48.546 34.612 52.92 ; 
      RECT 34.076 48.546 34.18 52.92 ; 
      RECT 33.644 48.546 33.748 52.92 ; 
      RECT 33.212 48.546 33.316 52.92 ; 
      RECT 32.78 48.546 32.884 52.92 ; 
      RECT 32.348 48.546 32.452 52.92 ; 
      RECT 31.916 48.546 32.02 52.92 ; 
      RECT 31.484 48.546 31.588 52.92 ; 
      RECT 31.052 48.546 31.156 52.92 ; 
      RECT 30.62 48.546 30.724 52.92 ; 
      RECT 30.188 48.546 30.292 52.92 ; 
      RECT 29.756 48.546 29.86 52.92 ; 
      RECT 29.324 48.546 29.428 52.92 ; 
      RECT 28.892 48.546 28.996 52.92 ; 
      RECT 28.46 48.546 28.564 52.92 ; 
      RECT 28.028 48.546 28.132 52.92 ; 
      RECT 27.596 48.546 27.7 52.92 ; 
      RECT 27.164 48.546 27.268 52.92 ; 
      RECT 26.732 48.546 26.836 52.92 ; 
      RECT 26.3 48.546 26.404 52.92 ; 
      RECT 25.868 48.546 25.972 52.92 ; 
      RECT 25.436 48.546 25.54 52.92 ; 
      RECT 25.004 48.546 25.108 52.92 ; 
      RECT 24.572 48.546 24.676 52.92 ; 
      RECT 24.14 48.546 24.244 52.92 ; 
      RECT 23.708 48.546 23.812 52.92 ; 
      RECT 22.856 48.546 23.164 52.92 ; 
      RECT 15.284 48.546 15.592 52.92 ; 
      RECT 14.636 48.546 14.74 52.92 ; 
      RECT 14.204 48.546 14.308 52.92 ; 
      RECT 13.772 48.546 13.876 52.92 ; 
      RECT 13.34 48.546 13.444 52.92 ; 
      RECT 12.908 48.546 13.012 52.92 ; 
      RECT 12.476 48.546 12.58 52.92 ; 
      RECT 12.044 48.546 12.148 52.92 ; 
      RECT 11.612 48.546 11.716 52.92 ; 
      RECT 11.18 48.546 11.284 52.92 ; 
      RECT 10.748 48.546 10.852 52.92 ; 
      RECT 10.316 48.546 10.42 52.92 ; 
      RECT 9.884 48.546 9.988 52.92 ; 
      RECT 9.452 48.546 9.556 52.92 ; 
      RECT 9.02 48.546 9.124 52.92 ; 
      RECT 8.588 48.546 8.692 52.92 ; 
      RECT 8.156 48.546 8.26 52.92 ; 
      RECT 7.724 48.546 7.828 52.92 ; 
      RECT 7.292 48.546 7.396 52.92 ; 
      RECT 6.86 48.546 6.964 52.92 ; 
      RECT 6.428 48.546 6.532 52.92 ; 
      RECT 5.996 48.546 6.1 52.92 ; 
      RECT 5.564 48.546 5.668 52.92 ; 
      RECT 5.132 48.546 5.236 52.92 ; 
      RECT 4.7 48.546 4.804 52.92 ; 
      RECT 4.268 48.546 4.372 52.92 ; 
      RECT 3.836 48.546 3.94 52.92 ; 
      RECT 3.404 48.546 3.508 52.92 ; 
      RECT 2.972 48.546 3.076 52.92 ; 
      RECT 2.54 48.546 2.644 52.92 ; 
      RECT 2.108 48.546 2.212 52.92 ; 
      RECT 1.676 48.546 1.78 52.92 ; 
      RECT 1.244 48.546 1.348 52.92 ; 
      RECT 0.812 48.546 0.916 52.92 ; 
      RECT 0 48.546 0.34 52.92 ; 
      RECT 20.72 52.866 21.232 57.24 ; 
      RECT 20.664 55.528 21.232 56.818 ; 
      RECT 20.072 54.436 20.32 57.24 ; 
      RECT 20.016 55.674 20.32 56.288 ; 
      RECT 20.072 52.866 20.176 57.24 ; 
      RECT 20.072 53.35 20.232 54.308 ; 
      RECT 20.072 52.866 20.32 53.222 ; 
      RECT 18.884 54.668 19.708 57.24 ; 
      RECT 19.604 52.866 19.708 57.24 ; 
      RECT 18.884 55.776 19.764 56.808 ; 
      RECT 18.884 52.866 19.276 57.24 ; 
      RECT 17.216 52.866 17.548 57.24 ; 
      RECT 17.216 53.22 17.604 56.962 ; 
      RECT 38.108 52.866 38.448 57.24 ; 
      RECT 37.532 52.866 37.636 57.24 ; 
      RECT 37.1 52.866 37.204 57.24 ; 
      RECT 36.668 52.866 36.772 57.24 ; 
      RECT 36.236 52.866 36.34 57.24 ; 
      RECT 35.804 52.866 35.908 57.24 ; 
      RECT 35.372 52.866 35.476 57.24 ; 
      RECT 34.94 52.866 35.044 57.24 ; 
      RECT 34.508 52.866 34.612 57.24 ; 
      RECT 34.076 52.866 34.18 57.24 ; 
      RECT 33.644 52.866 33.748 57.24 ; 
      RECT 33.212 52.866 33.316 57.24 ; 
      RECT 32.78 52.866 32.884 57.24 ; 
      RECT 32.348 52.866 32.452 57.24 ; 
      RECT 31.916 52.866 32.02 57.24 ; 
      RECT 31.484 52.866 31.588 57.24 ; 
      RECT 31.052 52.866 31.156 57.24 ; 
      RECT 30.62 52.866 30.724 57.24 ; 
      RECT 30.188 52.866 30.292 57.24 ; 
      RECT 29.756 52.866 29.86 57.24 ; 
      RECT 29.324 52.866 29.428 57.24 ; 
      RECT 28.892 52.866 28.996 57.24 ; 
      RECT 28.46 52.866 28.564 57.24 ; 
      RECT 28.028 52.866 28.132 57.24 ; 
      RECT 27.596 52.866 27.7 57.24 ; 
      RECT 27.164 52.866 27.268 57.24 ; 
      RECT 26.732 52.866 26.836 57.24 ; 
      RECT 26.3 52.866 26.404 57.24 ; 
      RECT 25.868 52.866 25.972 57.24 ; 
      RECT 25.436 52.866 25.54 57.24 ; 
      RECT 25.004 52.866 25.108 57.24 ; 
      RECT 24.572 52.866 24.676 57.24 ; 
      RECT 24.14 52.866 24.244 57.24 ; 
      RECT 23.708 52.866 23.812 57.24 ; 
      RECT 22.856 52.866 23.164 57.24 ; 
      RECT 15.284 52.866 15.592 57.24 ; 
      RECT 14.636 52.866 14.74 57.24 ; 
      RECT 14.204 52.866 14.308 57.24 ; 
      RECT 13.772 52.866 13.876 57.24 ; 
      RECT 13.34 52.866 13.444 57.24 ; 
      RECT 12.908 52.866 13.012 57.24 ; 
      RECT 12.476 52.866 12.58 57.24 ; 
      RECT 12.044 52.866 12.148 57.24 ; 
      RECT 11.612 52.866 11.716 57.24 ; 
      RECT 11.18 52.866 11.284 57.24 ; 
      RECT 10.748 52.866 10.852 57.24 ; 
      RECT 10.316 52.866 10.42 57.24 ; 
      RECT 9.884 52.866 9.988 57.24 ; 
      RECT 9.452 52.866 9.556 57.24 ; 
      RECT 9.02 52.866 9.124 57.24 ; 
      RECT 8.588 52.866 8.692 57.24 ; 
      RECT 8.156 52.866 8.26 57.24 ; 
      RECT 7.724 52.866 7.828 57.24 ; 
      RECT 7.292 52.866 7.396 57.24 ; 
      RECT 6.86 52.866 6.964 57.24 ; 
      RECT 6.428 52.866 6.532 57.24 ; 
      RECT 5.996 52.866 6.1 57.24 ; 
      RECT 5.564 52.866 5.668 57.24 ; 
      RECT 5.132 52.866 5.236 57.24 ; 
      RECT 4.7 52.866 4.804 57.24 ; 
      RECT 4.268 52.866 4.372 57.24 ; 
      RECT 3.836 52.866 3.94 57.24 ; 
      RECT 3.404 52.866 3.508 57.24 ; 
      RECT 2.972 52.866 3.076 57.24 ; 
      RECT 2.54 52.866 2.644 57.24 ; 
      RECT 2.108 52.866 2.212 57.24 ; 
      RECT 1.676 52.866 1.78 57.24 ; 
      RECT 1.244 52.866 1.348 57.24 ; 
      RECT 0.812 52.866 0.916 57.24 ; 
      RECT 0 52.866 0.34 57.24 ; 
      RECT 20.72 57.186 21.232 61.56 ; 
      RECT 20.664 59.848 21.232 61.138 ; 
      RECT 20.072 58.756 20.32 61.56 ; 
      RECT 20.016 59.994 20.32 60.608 ; 
      RECT 20.072 57.186 20.176 61.56 ; 
      RECT 20.072 57.67 20.232 58.628 ; 
      RECT 20.072 57.186 20.32 57.542 ; 
      RECT 18.884 58.988 19.708 61.56 ; 
      RECT 19.604 57.186 19.708 61.56 ; 
      RECT 18.884 60.096 19.764 61.128 ; 
      RECT 18.884 57.186 19.276 61.56 ; 
      RECT 17.216 57.186 17.548 61.56 ; 
      RECT 17.216 57.54 17.604 61.282 ; 
      RECT 38.108 57.186 38.448 61.56 ; 
      RECT 37.532 57.186 37.636 61.56 ; 
      RECT 37.1 57.186 37.204 61.56 ; 
      RECT 36.668 57.186 36.772 61.56 ; 
      RECT 36.236 57.186 36.34 61.56 ; 
      RECT 35.804 57.186 35.908 61.56 ; 
      RECT 35.372 57.186 35.476 61.56 ; 
      RECT 34.94 57.186 35.044 61.56 ; 
      RECT 34.508 57.186 34.612 61.56 ; 
      RECT 34.076 57.186 34.18 61.56 ; 
      RECT 33.644 57.186 33.748 61.56 ; 
      RECT 33.212 57.186 33.316 61.56 ; 
      RECT 32.78 57.186 32.884 61.56 ; 
      RECT 32.348 57.186 32.452 61.56 ; 
      RECT 31.916 57.186 32.02 61.56 ; 
      RECT 31.484 57.186 31.588 61.56 ; 
      RECT 31.052 57.186 31.156 61.56 ; 
      RECT 30.62 57.186 30.724 61.56 ; 
      RECT 30.188 57.186 30.292 61.56 ; 
      RECT 29.756 57.186 29.86 61.56 ; 
      RECT 29.324 57.186 29.428 61.56 ; 
      RECT 28.892 57.186 28.996 61.56 ; 
      RECT 28.46 57.186 28.564 61.56 ; 
      RECT 28.028 57.186 28.132 61.56 ; 
      RECT 27.596 57.186 27.7 61.56 ; 
      RECT 27.164 57.186 27.268 61.56 ; 
      RECT 26.732 57.186 26.836 61.56 ; 
      RECT 26.3 57.186 26.404 61.56 ; 
      RECT 25.868 57.186 25.972 61.56 ; 
      RECT 25.436 57.186 25.54 61.56 ; 
      RECT 25.004 57.186 25.108 61.56 ; 
      RECT 24.572 57.186 24.676 61.56 ; 
      RECT 24.14 57.186 24.244 61.56 ; 
      RECT 23.708 57.186 23.812 61.56 ; 
      RECT 22.856 57.186 23.164 61.56 ; 
      RECT 15.284 57.186 15.592 61.56 ; 
      RECT 14.636 57.186 14.74 61.56 ; 
      RECT 14.204 57.186 14.308 61.56 ; 
      RECT 13.772 57.186 13.876 61.56 ; 
      RECT 13.34 57.186 13.444 61.56 ; 
      RECT 12.908 57.186 13.012 61.56 ; 
      RECT 12.476 57.186 12.58 61.56 ; 
      RECT 12.044 57.186 12.148 61.56 ; 
      RECT 11.612 57.186 11.716 61.56 ; 
      RECT 11.18 57.186 11.284 61.56 ; 
      RECT 10.748 57.186 10.852 61.56 ; 
      RECT 10.316 57.186 10.42 61.56 ; 
      RECT 9.884 57.186 9.988 61.56 ; 
      RECT 9.452 57.186 9.556 61.56 ; 
      RECT 9.02 57.186 9.124 61.56 ; 
      RECT 8.588 57.186 8.692 61.56 ; 
      RECT 8.156 57.186 8.26 61.56 ; 
      RECT 7.724 57.186 7.828 61.56 ; 
      RECT 7.292 57.186 7.396 61.56 ; 
      RECT 6.86 57.186 6.964 61.56 ; 
      RECT 6.428 57.186 6.532 61.56 ; 
      RECT 5.996 57.186 6.1 61.56 ; 
      RECT 5.564 57.186 5.668 61.56 ; 
      RECT 5.132 57.186 5.236 61.56 ; 
      RECT 4.7 57.186 4.804 61.56 ; 
      RECT 4.268 57.186 4.372 61.56 ; 
      RECT 3.836 57.186 3.94 61.56 ; 
      RECT 3.404 57.186 3.508 61.56 ; 
      RECT 2.972 57.186 3.076 61.56 ; 
      RECT 2.54 57.186 2.644 61.56 ; 
      RECT 2.108 57.186 2.212 61.56 ; 
      RECT 1.676 57.186 1.78 61.56 ; 
      RECT 1.244 57.186 1.348 61.56 ; 
      RECT 0.812 57.186 0.916 61.56 ; 
      RECT 0 57.186 0.34 61.56 ; 
      RECT 20.72 61.506 21.232 65.88 ; 
      RECT 20.664 64.168 21.232 65.458 ; 
      RECT 20.072 63.076 20.32 65.88 ; 
      RECT 20.016 64.314 20.32 64.928 ; 
      RECT 20.072 61.506 20.176 65.88 ; 
      RECT 20.072 61.99 20.232 62.948 ; 
      RECT 20.072 61.506 20.32 61.862 ; 
      RECT 18.884 63.308 19.708 65.88 ; 
      RECT 19.604 61.506 19.708 65.88 ; 
      RECT 18.884 64.416 19.764 65.448 ; 
      RECT 18.884 61.506 19.276 65.88 ; 
      RECT 17.216 61.506 17.548 65.88 ; 
      RECT 17.216 61.86 17.604 65.602 ; 
      RECT 38.108 61.506 38.448 65.88 ; 
      RECT 37.532 61.506 37.636 65.88 ; 
      RECT 37.1 61.506 37.204 65.88 ; 
      RECT 36.668 61.506 36.772 65.88 ; 
      RECT 36.236 61.506 36.34 65.88 ; 
      RECT 35.804 61.506 35.908 65.88 ; 
      RECT 35.372 61.506 35.476 65.88 ; 
      RECT 34.94 61.506 35.044 65.88 ; 
      RECT 34.508 61.506 34.612 65.88 ; 
      RECT 34.076 61.506 34.18 65.88 ; 
      RECT 33.644 61.506 33.748 65.88 ; 
      RECT 33.212 61.506 33.316 65.88 ; 
      RECT 32.78 61.506 32.884 65.88 ; 
      RECT 32.348 61.506 32.452 65.88 ; 
      RECT 31.916 61.506 32.02 65.88 ; 
      RECT 31.484 61.506 31.588 65.88 ; 
      RECT 31.052 61.506 31.156 65.88 ; 
      RECT 30.62 61.506 30.724 65.88 ; 
      RECT 30.188 61.506 30.292 65.88 ; 
      RECT 29.756 61.506 29.86 65.88 ; 
      RECT 29.324 61.506 29.428 65.88 ; 
      RECT 28.892 61.506 28.996 65.88 ; 
      RECT 28.46 61.506 28.564 65.88 ; 
      RECT 28.028 61.506 28.132 65.88 ; 
      RECT 27.596 61.506 27.7 65.88 ; 
      RECT 27.164 61.506 27.268 65.88 ; 
      RECT 26.732 61.506 26.836 65.88 ; 
      RECT 26.3 61.506 26.404 65.88 ; 
      RECT 25.868 61.506 25.972 65.88 ; 
      RECT 25.436 61.506 25.54 65.88 ; 
      RECT 25.004 61.506 25.108 65.88 ; 
      RECT 24.572 61.506 24.676 65.88 ; 
      RECT 24.14 61.506 24.244 65.88 ; 
      RECT 23.708 61.506 23.812 65.88 ; 
      RECT 22.856 61.506 23.164 65.88 ; 
      RECT 15.284 61.506 15.592 65.88 ; 
      RECT 14.636 61.506 14.74 65.88 ; 
      RECT 14.204 61.506 14.308 65.88 ; 
      RECT 13.772 61.506 13.876 65.88 ; 
      RECT 13.34 61.506 13.444 65.88 ; 
      RECT 12.908 61.506 13.012 65.88 ; 
      RECT 12.476 61.506 12.58 65.88 ; 
      RECT 12.044 61.506 12.148 65.88 ; 
      RECT 11.612 61.506 11.716 65.88 ; 
      RECT 11.18 61.506 11.284 65.88 ; 
      RECT 10.748 61.506 10.852 65.88 ; 
      RECT 10.316 61.506 10.42 65.88 ; 
      RECT 9.884 61.506 9.988 65.88 ; 
      RECT 9.452 61.506 9.556 65.88 ; 
      RECT 9.02 61.506 9.124 65.88 ; 
      RECT 8.588 61.506 8.692 65.88 ; 
      RECT 8.156 61.506 8.26 65.88 ; 
      RECT 7.724 61.506 7.828 65.88 ; 
      RECT 7.292 61.506 7.396 65.88 ; 
      RECT 6.86 61.506 6.964 65.88 ; 
      RECT 6.428 61.506 6.532 65.88 ; 
      RECT 5.996 61.506 6.1 65.88 ; 
      RECT 5.564 61.506 5.668 65.88 ; 
      RECT 5.132 61.506 5.236 65.88 ; 
      RECT 4.7 61.506 4.804 65.88 ; 
      RECT 4.268 61.506 4.372 65.88 ; 
      RECT 3.836 61.506 3.94 65.88 ; 
      RECT 3.404 61.506 3.508 65.88 ; 
      RECT 2.972 61.506 3.076 65.88 ; 
      RECT 2.54 61.506 2.644 65.88 ; 
      RECT 2.108 61.506 2.212 65.88 ; 
      RECT 1.676 61.506 1.78 65.88 ; 
      RECT 1.244 61.506 1.348 65.88 ; 
      RECT 0.812 61.506 0.916 65.88 ; 
      RECT 0 61.506 0.34 65.88 ; 
      RECT 20.72 65.826 21.232 70.2 ; 
      RECT 20.664 68.488 21.232 69.778 ; 
      RECT 20.072 67.396 20.32 70.2 ; 
      RECT 20.016 68.634 20.32 69.248 ; 
      RECT 20.072 65.826 20.176 70.2 ; 
      RECT 20.072 66.31 20.232 67.268 ; 
      RECT 20.072 65.826 20.32 66.182 ; 
      RECT 18.884 67.628 19.708 70.2 ; 
      RECT 19.604 65.826 19.708 70.2 ; 
      RECT 18.884 68.736 19.764 69.768 ; 
      RECT 18.884 65.826 19.276 70.2 ; 
      RECT 17.216 65.826 17.548 70.2 ; 
      RECT 17.216 66.18 17.604 69.922 ; 
      RECT 38.108 65.826 38.448 70.2 ; 
      RECT 37.532 65.826 37.636 70.2 ; 
      RECT 37.1 65.826 37.204 70.2 ; 
      RECT 36.668 65.826 36.772 70.2 ; 
      RECT 36.236 65.826 36.34 70.2 ; 
      RECT 35.804 65.826 35.908 70.2 ; 
      RECT 35.372 65.826 35.476 70.2 ; 
      RECT 34.94 65.826 35.044 70.2 ; 
      RECT 34.508 65.826 34.612 70.2 ; 
      RECT 34.076 65.826 34.18 70.2 ; 
      RECT 33.644 65.826 33.748 70.2 ; 
      RECT 33.212 65.826 33.316 70.2 ; 
      RECT 32.78 65.826 32.884 70.2 ; 
      RECT 32.348 65.826 32.452 70.2 ; 
      RECT 31.916 65.826 32.02 70.2 ; 
      RECT 31.484 65.826 31.588 70.2 ; 
      RECT 31.052 65.826 31.156 70.2 ; 
      RECT 30.62 65.826 30.724 70.2 ; 
      RECT 30.188 65.826 30.292 70.2 ; 
      RECT 29.756 65.826 29.86 70.2 ; 
      RECT 29.324 65.826 29.428 70.2 ; 
      RECT 28.892 65.826 28.996 70.2 ; 
      RECT 28.46 65.826 28.564 70.2 ; 
      RECT 28.028 65.826 28.132 70.2 ; 
      RECT 27.596 65.826 27.7 70.2 ; 
      RECT 27.164 65.826 27.268 70.2 ; 
      RECT 26.732 65.826 26.836 70.2 ; 
      RECT 26.3 65.826 26.404 70.2 ; 
      RECT 25.868 65.826 25.972 70.2 ; 
      RECT 25.436 65.826 25.54 70.2 ; 
      RECT 25.004 65.826 25.108 70.2 ; 
      RECT 24.572 65.826 24.676 70.2 ; 
      RECT 24.14 65.826 24.244 70.2 ; 
      RECT 23.708 65.826 23.812 70.2 ; 
      RECT 22.856 65.826 23.164 70.2 ; 
      RECT 15.284 65.826 15.592 70.2 ; 
      RECT 14.636 65.826 14.74 70.2 ; 
      RECT 14.204 65.826 14.308 70.2 ; 
      RECT 13.772 65.826 13.876 70.2 ; 
      RECT 13.34 65.826 13.444 70.2 ; 
      RECT 12.908 65.826 13.012 70.2 ; 
      RECT 12.476 65.826 12.58 70.2 ; 
      RECT 12.044 65.826 12.148 70.2 ; 
      RECT 11.612 65.826 11.716 70.2 ; 
      RECT 11.18 65.826 11.284 70.2 ; 
      RECT 10.748 65.826 10.852 70.2 ; 
      RECT 10.316 65.826 10.42 70.2 ; 
      RECT 9.884 65.826 9.988 70.2 ; 
      RECT 9.452 65.826 9.556 70.2 ; 
      RECT 9.02 65.826 9.124 70.2 ; 
      RECT 8.588 65.826 8.692 70.2 ; 
      RECT 8.156 65.826 8.26 70.2 ; 
      RECT 7.724 65.826 7.828 70.2 ; 
      RECT 7.292 65.826 7.396 70.2 ; 
      RECT 6.86 65.826 6.964 70.2 ; 
      RECT 6.428 65.826 6.532 70.2 ; 
      RECT 5.996 65.826 6.1 70.2 ; 
      RECT 5.564 65.826 5.668 70.2 ; 
      RECT 5.132 65.826 5.236 70.2 ; 
      RECT 4.7 65.826 4.804 70.2 ; 
      RECT 4.268 65.826 4.372 70.2 ; 
      RECT 3.836 65.826 3.94 70.2 ; 
      RECT 3.404 65.826 3.508 70.2 ; 
      RECT 2.972 65.826 3.076 70.2 ; 
      RECT 2.54 65.826 2.644 70.2 ; 
      RECT 2.108 65.826 2.212 70.2 ; 
      RECT 1.676 65.826 1.78 70.2 ; 
      RECT 1.244 65.826 1.348 70.2 ; 
      RECT 0.812 65.826 0.916 70.2 ; 
      RECT 0 65.826 0.34 70.2 ; 
      RECT 20.72 70.146 21.232 74.52 ; 
      RECT 20.664 72.808 21.232 74.098 ; 
      RECT 20.072 71.716 20.32 74.52 ; 
      RECT 20.016 72.954 20.32 73.568 ; 
      RECT 20.072 70.146 20.176 74.52 ; 
      RECT 20.072 70.63 20.232 71.588 ; 
      RECT 20.072 70.146 20.32 70.502 ; 
      RECT 18.884 71.948 19.708 74.52 ; 
      RECT 19.604 70.146 19.708 74.52 ; 
      RECT 18.884 73.056 19.764 74.088 ; 
      RECT 18.884 70.146 19.276 74.52 ; 
      RECT 17.216 70.146 17.548 74.52 ; 
      RECT 17.216 70.5 17.604 74.242 ; 
      RECT 38.108 70.146 38.448 74.52 ; 
      RECT 37.532 70.146 37.636 74.52 ; 
      RECT 37.1 70.146 37.204 74.52 ; 
      RECT 36.668 70.146 36.772 74.52 ; 
      RECT 36.236 70.146 36.34 74.52 ; 
      RECT 35.804 70.146 35.908 74.52 ; 
      RECT 35.372 70.146 35.476 74.52 ; 
      RECT 34.94 70.146 35.044 74.52 ; 
      RECT 34.508 70.146 34.612 74.52 ; 
      RECT 34.076 70.146 34.18 74.52 ; 
      RECT 33.644 70.146 33.748 74.52 ; 
      RECT 33.212 70.146 33.316 74.52 ; 
      RECT 32.78 70.146 32.884 74.52 ; 
      RECT 32.348 70.146 32.452 74.52 ; 
      RECT 31.916 70.146 32.02 74.52 ; 
      RECT 31.484 70.146 31.588 74.52 ; 
      RECT 31.052 70.146 31.156 74.52 ; 
      RECT 30.62 70.146 30.724 74.52 ; 
      RECT 30.188 70.146 30.292 74.52 ; 
      RECT 29.756 70.146 29.86 74.52 ; 
      RECT 29.324 70.146 29.428 74.52 ; 
      RECT 28.892 70.146 28.996 74.52 ; 
      RECT 28.46 70.146 28.564 74.52 ; 
      RECT 28.028 70.146 28.132 74.52 ; 
      RECT 27.596 70.146 27.7 74.52 ; 
      RECT 27.164 70.146 27.268 74.52 ; 
      RECT 26.732 70.146 26.836 74.52 ; 
      RECT 26.3 70.146 26.404 74.52 ; 
      RECT 25.868 70.146 25.972 74.52 ; 
      RECT 25.436 70.146 25.54 74.52 ; 
      RECT 25.004 70.146 25.108 74.52 ; 
      RECT 24.572 70.146 24.676 74.52 ; 
      RECT 24.14 70.146 24.244 74.52 ; 
      RECT 23.708 70.146 23.812 74.52 ; 
      RECT 22.856 70.146 23.164 74.52 ; 
      RECT 15.284 70.146 15.592 74.52 ; 
      RECT 14.636 70.146 14.74 74.52 ; 
      RECT 14.204 70.146 14.308 74.52 ; 
      RECT 13.772 70.146 13.876 74.52 ; 
      RECT 13.34 70.146 13.444 74.52 ; 
      RECT 12.908 70.146 13.012 74.52 ; 
      RECT 12.476 70.146 12.58 74.52 ; 
      RECT 12.044 70.146 12.148 74.52 ; 
      RECT 11.612 70.146 11.716 74.52 ; 
      RECT 11.18 70.146 11.284 74.52 ; 
      RECT 10.748 70.146 10.852 74.52 ; 
      RECT 10.316 70.146 10.42 74.52 ; 
      RECT 9.884 70.146 9.988 74.52 ; 
      RECT 9.452 70.146 9.556 74.52 ; 
      RECT 9.02 70.146 9.124 74.52 ; 
      RECT 8.588 70.146 8.692 74.52 ; 
      RECT 8.156 70.146 8.26 74.52 ; 
      RECT 7.724 70.146 7.828 74.52 ; 
      RECT 7.292 70.146 7.396 74.52 ; 
      RECT 6.86 70.146 6.964 74.52 ; 
      RECT 6.428 70.146 6.532 74.52 ; 
      RECT 5.996 70.146 6.1 74.52 ; 
      RECT 5.564 70.146 5.668 74.52 ; 
      RECT 5.132 70.146 5.236 74.52 ; 
      RECT 4.7 70.146 4.804 74.52 ; 
      RECT 4.268 70.146 4.372 74.52 ; 
      RECT 3.836 70.146 3.94 74.52 ; 
      RECT 3.404 70.146 3.508 74.52 ; 
      RECT 2.972 70.146 3.076 74.52 ; 
      RECT 2.54 70.146 2.644 74.52 ; 
      RECT 2.108 70.146 2.212 74.52 ; 
      RECT 1.676 70.146 1.78 74.52 ; 
      RECT 1.244 70.146 1.348 74.52 ; 
      RECT 0.812 70.146 0.916 74.52 ; 
      RECT 0 70.146 0.34 74.52 ; 
      RECT 20.72 74.466 21.232 78.84 ; 
      RECT 20.664 77.128 21.232 78.418 ; 
      RECT 20.072 76.036 20.32 78.84 ; 
      RECT 20.016 77.274 20.32 77.888 ; 
      RECT 20.072 74.466 20.176 78.84 ; 
      RECT 20.072 74.95 20.232 75.908 ; 
      RECT 20.072 74.466 20.32 74.822 ; 
      RECT 18.884 76.268 19.708 78.84 ; 
      RECT 19.604 74.466 19.708 78.84 ; 
      RECT 18.884 77.376 19.764 78.408 ; 
      RECT 18.884 74.466 19.276 78.84 ; 
      RECT 17.216 74.466 17.548 78.84 ; 
      RECT 17.216 74.82 17.604 78.562 ; 
      RECT 38.108 74.466 38.448 78.84 ; 
      RECT 37.532 74.466 37.636 78.84 ; 
      RECT 37.1 74.466 37.204 78.84 ; 
      RECT 36.668 74.466 36.772 78.84 ; 
      RECT 36.236 74.466 36.34 78.84 ; 
      RECT 35.804 74.466 35.908 78.84 ; 
      RECT 35.372 74.466 35.476 78.84 ; 
      RECT 34.94 74.466 35.044 78.84 ; 
      RECT 34.508 74.466 34.612 78.84 ; 
      RECT 34.076 74.466 34.18 78.84 ; 
      RECT 33.644 74.466 33.748 78.84 ; 
      RECT 33.212 74.466 33.316 78.84 ; 
      RECT 32.78 74.466 32.884 78.84 ; 
      RECT 32.348 74.466 32.452 78.84 ; 
      RECT 31.916 74.466 32.02 78.84 ; 
      RECT 31.484 74.466 31.588 78.84 ; 
      RECT 31.052 74.466 31.156 78.84 ; 
      RECT 30.62 74.466 30.724 78.84 ; 
      RECT 30.188 74.466 30.292 78.84 ; 
      RECT 29.756 74.466 29.86 78.84 ; 
      RECT 29.324 74.466 29.428 78.84 ; 
      RECT 28.892 74.466 28.996 78.84 ; 
      RECT 28.46 74.466 28.564 78.84 ; 
      RECT 28.028 74.466 28.132 78.84 ; 
      RECT 27.596 74.466 27.7 78.84 ; 
      RECT 27.164 74.466 27.268 78.84 ; 
      RECT 26.732 74.466 26.836 78.84 ; 
      RECT 26.3 74.466 26.404 78.84 ; 
      RECT 25.868 74.466 25.972 78.84 ; 
      RECT 25.436 74.466 25.54 78.84 ; 
      RECT 25.004 74.466 25.108 78.84 ; 
      RECT 24.572 74.466 24.676 78.84 ; 
      RECT 24.14 74.466 24.244 78.84 ; 
      RECT 23.708 74.466 23.812 78.84 ; 
      RECT 22.856 74.466 23.164 78.84 ; 
      RECT 15.284 74.466 15.592 78.84 ; 
      RECT 14.636 74.466 14.74 78.84 ; 
      RECT 14.204 74.466 14.308 78.84 ; 
      RECT 13.772 74.466 13.876 78.84 ; 
      RECT 13.34 74.466 13.444 78.84 ; 
      RECT 12.908 74.466 13.012 78.84 ; 
      RECT 12.476 74.466 12.58 78.84 ; 
      RECT 12.044 74.466 12.148 78.84 ; 
      RECT 11.612 74.466 11.716 78.84 ; 
      RECT 11.18 74.466 11.284 78.84 ; 
      RECT 10.748 74.466 10.852 78.84 ; 
      RECT 10.316 74.466 10.42 78.84 ; 
      RECT 9.884 74.466 9.988 78.84 ; 
      RECT 9.452 74.466 9.556 78.84 ; 
      RECT 9.02 74.466 9.124 78.84 ; 
      RECT 8.588 74.466 8.692 78.84 ; 
      RECT 8.156 74.466 8.26 78.84 ; 
      RECT 7.724 74.466 7.828 78.84 ; 
      RECT 7.292 74.466 7.396 78.84 ; 
      RECT 6.86 74.466 6.964 78.84 ; 
      RECT 6.428 74.466 6.532 78.84 ; 
      RECT 5.996 74.466 6.1 78.84 ; 
      RECT 5.564 74.466 5.668 78.84 ; 
      RECT 5.132 74.466 5.236 78.84 ; 
      RECT 4.7 74.466 4.804 78.84 ; 
      RECT 4.268 74.466 4.372 78.84 ; 
      RECT 3.836 74.466 3.94 78.84 ; 
      RECT 3.404 74.466 3.508 78.84 ; 
      RECT 2.972 74.466 3.076 78.84 ; 
      RECT 2.54 74.466 2.644 78.84 ; 
      RECT 2.108 74.466 2.212 78.84 ; 
      RECT 1.676 74.466 1.78 78.84 ; 
      RECT 1.244 74.466 1.348 78.84 ; 
      RECT 0.812 74.466 0.916 78.84 ; 
      RECT 0 74.466 0.34 78.84 ; 
      RECT 20.72 78.786 21.232 83.16 ; 
      RECT 20.664 81.448 21.232 82.738 ; 
      RECT 20.072 80.356 20.32 83.16 ; 
      RECT 20.016 81.594 20.32 82.208 ; 
      RECT 20.072 78.786 20.176 83.16 ; 
      RECT 20.072 79.27 20.232 80.228 ; 
      RECT 20.072 78.786 20.32 79.142 ; 
      RECT 18.884 80.588 19.708 83.16 ; 
      RECT 19.604 78.786 19.708 83.16 ; 
      RECT 18.884 81.696 19.764 82.728 ; 
      RECT 18.884 78.786 19.276 83.16 ; 
      RECT 17.216 78.786 17.548 83.16 ; 
      RECT 17.216 79.14 17.604 82.882 ; 
      RECT 38.108 78.786 38.448 83.16 ; 
      RECT 37.532 78.786 37.636 83.16 ; 
      RECT 37.1 78.786 37.204 83.16 ; 
      RECT 36.668 78.786 36.772 83.16 ; 
      RECT 36.236 78.786 36.34 83.16 ; 
      RECT 35.804 78.786 35.908 83.16 ; 
      RECT 35.372 78.786 35.476 83.16 ; 
      RECT 34.94 78.786 35.044 83.16 ; 
      RECT 34.508 78.786 34.612 83.16 ; 
      RECT 34.076 78.786 34.18 83.16 ; 
      RECT 33.644 78.786 33.748 83.16 ; 
      RECT 33.212 78.786 33.316 83.16 ; 
      RECT 32.78 78.786 32.884 83.16 ; 
      RECT 32.348 78.786 32.452 83.16 ; 
      RECT 31.916 78.786 32.02 83.16 ; 
      RECT 31.484 78.786 31.588 83.16 ; 
      RECT 31.052 78.786 31.156 83.16 ; 
      RECT 30.62 78.786 30.724 83.16 ; 
      RECT 30.188 78.786 30.292 83.16 ; 
      RECT 29.756 78.786 29.86 83.16 ; 
      RECT 29.324 78.786 29.428 83.16 ; 
      RECT 28.892 78.786 28.996 83.16 ; 
      RECT 28.46 78.786 28.564 83.16 ; 
      RECT 28.028 78.786 28.132 83.16 ; 
      RECT 27.596 78.786 27.7 83.16 ; 
      RECT 27.164 78.786 27.268 83.16 ; 
      RECT 26.732 78.786 26.836 83.16 ; 
      RECT 26.3 78.786 26.404 83.16 ; 
      RECT 25.868 78.786 25.972 83.16 ; 
      RECT 25.436 78.786 25.54 83.16 ; 
      RECT 25.004 78.786 25.108 83.16 ; 
      RECT 24.572 78.786 24.676 83.16 ; 
      RECT 24.14 78.786 24.244 83.16 ; 
      RECT 23.708 78.786 23.812 83.16 ; 
      RECT 22.856 78.786 23.164 83.16 ; 
      RECT 15.284 78.786 15.592 83.16 ; 
      RECT 14.636 78.786 14.74 83.16 ; 
      RECT 14.204 78.786 14.308 83.16 ; 
      RECT 13.772 78.786 13.876 83.16 ; 
      RECT 13.34 78.786 13.444 83.16 ; 
      RECT 12.908 78.786 13.012 83.16 ; 
      RECT 12.476 78.786 12.58 83.16 ; 
      RECT 12.044 78.786 12.148 83.16 ; 
      RECT 11.612 78.786 11.716 83.16 ; 
      RECT 11.18 78.786 11.284 83.16 ; 
      RECT 10.748 78.786 10.852 83.16 ; 
      RECT 10.316 78.786 10.42 83.16 ; 
      RECT 9.884 78.786 9.988 83.16 ; 
      RECT 9.452 78.786 9.556 83.16 ; 
      RECT 9.02 78.786 9.124 83.16 ; 
      RECT 8.588 78.786 8.692 83.16 ; 
      RECT 8.156 78.786 8.26 83.16 ; 
      RECT 7.724 78.786 7.828 83.16 ; 
      RECT 7.292 78.786 7.396 83.16 ; 
      RECT 6.86 78.786 6.964 83.16 ; 
      RECT 6.428 78.786 6.532 83.16 ; 
      RECT 5.996 78.786 6.1 83.16 ; 
      RECT 5.564 78.786 5.668 83.16 ; 
      RECT 5.132 78.786 5.236 83.16 ; 
      RECT 4.7 78.786 4.804 83.16 ; 
      RECT 4.268 78.786 4.372 83.16 ; 
      RECT 3.836 78.786 3.94 83.16 ; 
      RECT 3.404 78.786 3.508 83.16 ; 
      RECT 2.972 78.786 3.076 83.16 ; 
      RECT 2.54 78.786 2.644 83.16 ; 
      RECT 2.108 78.786 2.212 83.16 ; 
      RECT 1.676 78.786 1.78 83.16 ; 
      RECT 1.244 78.786 1.348 83.16 ; 
      RECT 0.812 78.786 0.916 83.16 ; 
      RECT 0 78.786 0.34 83.16 ; 
      RECT 20.72 83.106 21.232 87.48 ; 
      RECT 20.664 85.768 21.232 87.058 ; 
      RECT 20.072 84.676 20.32 87.48 ; 
      RECT 20.016 85.914 20.32 86.528 ; 
      RECT 20.072 83.106 20.176 87.48 ; 
      RECT 20.072 83.59 20.232 84.548 ; 
      RECT 20.072 83.106 20.32 83.462 ; 
      RECT 18.884 84.908 19.708 87.48 ; 
      RECT 19.604 83.106 19.708 87.48 ; 
      RECT 18.884 86.016 19.764 87.048 ; 
      RECT 18.884 83.106 19.276 87.48 ; 
      RECT 17.216 83.106 17.548 87.48 ; 
      RECT 17.216 83.46 17.604 87.202 ; 
      RECT 38.108 83.106 38.448 87.48 ; 
      RECT 37.532 83.106 37.636 87.48 ; 
      RECT 37.1 83.106 37.204 87.48 ; 
      RECT 36.668 83.106 36.772 87.48 ; 
      RECT 36.236 83.106 36.34 87.48 ; 
      RECT 35.804 83.106 35.908 87.48 ; 
      RECT 35.372 83.106 35.476 87.48 ; 
      RECT 34.94 83.106 35.044 87.48 ; 
      RECT 34.508 83.106 34.612 87.48 ; 
      RECT 34.076 83.106 34.18 87.48 ; 
      RECT 33.644 83.106 33.748 87.48 ; 
      RECT 33.212 83.106 33.316 87.48 ; 
      RECT 32.78 83.106 32.884 87.48 ; 
      RECT 32.348 83.106 32.452 87.48 ; 
      RECT 31.916 83.106 32.02 87.48 ; 
      RECT 31.484 83.106 31.588 87.48 ; 
      RECT 31.052 83.106 31.156 87.48 ; 
      RECT 30.62 83.106 30.724 87.48 ; 
      RECT 30.188 83.106 30.292 87.48 ; 
      RECT 29.756 83.106 29.86 87.48 ; 
      RECT 29.324 83.106 29.428 87.48 ; 
      RECT 28.892 83.106 28.996 87.48 ; 
      RECT 28.46 83.106 28.564 87.48 ; 
      RECT 28.028 83.106 28.132 87.48 ; 
      RECT 27.596 83.106 27.7 87.48 ; 
      RECT 27.164 83.106 27.268 87.48 ; 
      RECT 26.732 83.106 26.836 87.48 ; 
      RECT 26.3 83.106 26.404 87.48 ; 
      RECT 25.868 83.106 25.972 87.48 ; 
      RECT 25.436 83.106 25.54 87.48 ; 
      RECT 25.004 83.106 25.108 87.48 ; 
      RECT 24.572 83.106 24.676 87.48 ; 
      RECT 24.14 83.106 24.244 87.48 ; 
      RECT 23.708 83.106 23.812 87.48 ; 
      RECT 22.856 83.106 23.164 87.48 ; 
      RECT 15.284 83.106 15.592 87.48 ; 
      RECT 14.636 83.106 14.74 87.48 ; 
      RECT 14.204 83.106 14.308 87.48 ; 
      RECT 13.772 83.106 13.876 87.48 ; 
      RECT 13.34 83.106 13.444 87.48 ; 
      RECT 12.908 83.106 13.012 87.48 ; 
      RECT 12.476 83.106 12.58 87.48 ; 
      RECT 12.044 83.106 12.148 87.48 ; 
      RECT 11.612 83.106 11.716 87.48 ; 
      RECT 11.18 83.106 11.284 87.48 ; 
      RECT 10.748 83.106 10.852 87.48 ; 
      RECT 10.316 83.106 10.42 87.48 ; 
      RECT 9.884 83.106 9.988 87.48 ; 
      RECT 9.452 83.106 9.556 87.48 ; 
      RECT 9.02 83.106 9.124 87.48 ; 
      RECT 8.588 83.106 8.692 87.48 ; 
      RECT 8.156 83.106 8.26 87.48 ; 
      RECT 7.724 83.106 7.828 87.48 ; 
      RECT 7.292 83.106 7.396 87.48 ; 
      RECT 6.86 83.106 6.964 87.48 ; 
      RECT 6.428 83.106 6.532 87.48 ; 
      RECT 5.996 83.106 6.1 87.48 ; 
      RECT 5.564 83.106 5.668 87.48 ; 
      RECT 5.132 83.106 5.236 87.48 ; 
      RECT 4.7 83.106 4.804 87.48 ; 
      RECT 4.268 83.106 4.372 87.48 ; 
      RECT 3.836 83.106 3.94 87.48 ; 
      RECT 3.404 83.106 3.508 87.48 ; 
      RECT 2.972 83.106 3.076 87.48 ; 
      RECT 2.54 83.106 2.644 87.48 ; 
      RECT 2.108 83.106 2.212 87.48 ; 
      RECT 1.676 83.106 1.78 87.48 ; 
      RECT 1.244 83.106 1.348 87.48 ; 
      RECT 0.812 83.106 0.916 87.48 ; 
      RECT 0 83.106 0.34 87.48 ; 
      RECT 20.72 87.426 21.232 91.8 ; 
      RECT 20.664 90.088 21.232 91.378 ; 
      RECT 20.072 88.996 20.32 91.8 ; 
      RECT 20.016 90.234 20.32 90.848 ; 
      RECT 20.072 87.426 20.176 91.8 ; 
      RECT 20.072 87.91 20.232 88.868 ; 
      RECT 20.072 87.426 20.32 87.782 ; 
      RECT 18.884 89.228 19.708 91.8 ; 
      RECT 19.604 87.426 19.708 91.8 ; 
      RECT 18.884 90.336 19.764 91.368 ; 
      RECT 18.884 87.426 19.276 91.8 ; 
      RECT 17.216 87.426 17.548 91.8 ; 
      RECT 17.216 87.78 17.604 91.522 ; 
      RECT 38.108 87.426 38.448 91.8 ; 
      RECT 37.532 87.426 37.636 91.8 ; 
      RECT 37.1 87.426 37.204 91.8 ; 
      RECT 36.668 87.426 36.772 91.8 ; 
      RECT 36.236 87.426 36.34 91.8 ; 
      RECT 35.804 87.426 35.908 91.8 ; 
      RECT 35.372 87.426 35.476 91.8 ; 
      RECT 34.94 87.426 35.044 91.8 ; 
      RECT 34.508 87.426 34.612 91.8 ; 
      RECT 34.076 87.426 34.18 91.8 ; 
      RECT 33.644 87.426 33.748 91.8 ; 
      RECT 33.212 87.426 33.316 91.8 ; 
      RECT 32.78 87.426 32.884 91.8 ; 
      RECT 32.348 87.426 32.452 91.8 ; 
      RECT 31.916 87.426 32.02 91.8 ; 
      RECT 31.484 87.426 31.588 91.8 ; 
      RECT 31.052 87.426 31.156 91.8 ; 
      RECT 30.62 87.426 30.724 91.8 ; 
      RECT 30.188 87.426 30.292 91.8 ; 
      RECT 29.756 87.426 29.86 91.8 ; 
      RECT 29.324 87.426 29.428 91.8 ; 
      RECT 28.892 87.426 28.996 91.8 ; 
      RECT 28.46 87.426 28.564 91.8 ; 
      RECT 28.028 87.426 28.132 91.8 ; 
      RECT 27.596 87.426 27.7 91.8 ; 
      RECT 27.164 87.426 27.268 91.8 ; 
      RECT 26.732 87.426 26.836 91.8 ; 
      RECT 26.3 87.426 26.404 91.8 ; 
      RECT 25.868 87.426 25.972 91.8 ; 
      RECT 25.436 87.426 25.54 91.8 ; 
      RECT 25.004 87.426 25.108 91.8 ; 
      RECT 24.572 87.426 24.676 91.8 ; 
      RECT 24.14 87.426 24.244 91.8 ; 
      RECT 23.708 87.426 23.812 91.8 ; 
      RECT 22.856 87.426 23.164 91.8 ; 
      RECT 15.284 87.426 15.592 91.8 ; 
      RECT 14.636 87.426 14.74 91.8 ; 
      RECT 14.204 87.426 14.308 91.8 ; 
      RECT 13.772 87.426 13.876 91.8 ; 
      RECT 13.34 87.426 13.444 91.8 ; 
      RECT 12.908 87.426 13.012 91.8 ; 
      RECT 12.476 87.426 12.58 91.8 ; 
      RECT 12.044 87.426 12.148 91.8 ; 
      RECT 11.612 87.426 11.716 91.8 ; 
      RECT 11.18 87.426 11.284 91.8 ; 
      RECT 10.748 87.426 10.852 91.8 ; 
      RECT 10.316 87.426 10.42 91.8 ; 
      RECT 9.884 87.426 9.988 91.8 ; 
      RECT 9.452 87.426 9.556 91.8 ; 
      RECT 9.02 87.426 9.124 91.8 ; 
      RECT 8.588 87.426 8.692 91.8 ; 
      RECT 8.156 87.426 8.26 91.8 ; 
      RECT 7.724 87.426 7.828 91.8 ; 
      RECT 7.292 87.426 7.396 91.8 ; 
      RECT 6.86 87.426 6.964 91.8 ; 
      RECT 6.428 87.426 6.532 91.8 ; 
      RECT 5.996 87.426 6.1 91.8 ; 
      RECT 5.564 87.426 5.668 91.8 ; 
      RECT 5.132 87.426 5.236 91.8 ; 
      RECT 4.7 87.426 4.804 91.8 ; 
      RECT 4.268 87.426 4.372 91.8 ; 
      RECT 3.836 87.426 3.94 91.8 ; 
      RECT 3.404 87.426 3.508 91.8 ; 
      RECT 2.972 87.426 3.076 91.8 ; 
      RECT 2.54 87.426 2.644 91.8 ; 
      RECT 2.108 87.426 2.212 91.8 ; 
      RECT 1.676 87.426 1.78 91.8 ; 
      RECT 1.244 87.426 1.348 91.8 ; 
      RECT 0.812 87.426 0.916 91.8 ; 
      RECT 0 87.426 0.34 91.8 ; 
      RECT 20.72 91.746 21.232 96.12 ; 
      RECT 20.664 94.408 21.232 95.698 ; 
      RECT 20.072 93.316 20.32 96.12 ; 
      RECT 20.016 94.554 20.32 95.168 ; 
      RECT 20.072 91.746 20.176 96.12 ; 
      RECT 20.072 92.23 20.232 93.188 ; 
      RECT 20.072 91.746 20.32 92.102 ; 
      RECT 18.884 93.548 19.708 96.12 ; 
      RECT 19.604 91.746 19.708 96.12 ; 
      RECT 18.884 94.656 19.764 95.688 ; 
      RECT 18.884 91.746 19.276 96.12 ; 
      RECT 17.216 91.746 17.548 96.12 ; 
      RECT 17.216 92.1 17.604 95.842 ; 
      RECT 38.108 91.746 38.448 96.12 ; 
      RECT 37.532 91.746 37.636 96.12 ; 
      RECT 37.1 91.746 37.204 96.12 ; 
      RECT 36.668 91.746 36.772 96.12 ; 
      RECT 36.236 91.746 36.34 96.12 ; 
      RECT 35.804 91.746 35.908 96.12 ; 
      RECT 35.372 91.746 35.476 96.12 ; 
      RECT 34.94 91.746 35.044 96.12 ; 
      RECT 34.508 91.746 34.612 96.12 ; 
      RECT 34.076 91.746 34.18 96.12 ; 
      RECT 33.644 91.746 33.748 96.12 ; 
      RECT 33.212 91.746 33.316 96.12 ; 
      RECT 32.78 91.746 32.884 96.12 ; 
      RECT 32.348 91.746 32.452 96.12 ; 
      RECT 31.916 91.746 32.02 96.12 ; 
      RECT 31.484 91.746 31.588 96.12 ; 
      RECT 31.052 91.746 31.156 96.12 ; 
      RECT 30.62 91.746 30.724 96.12 ; 
      RECT 30.188 91.746 30.292 96.12 ; 
      RECT 29.756 91.746 29.86 96.12 ; 
      RECT 29.324 91.746 29.428 96.12 ; 
      RECT 28.892 91.746 28.996 96.12 ; 
      RECT 28.46 91.746 28.564 96.12 ; 
      RECT 28.028 91.746 28.132 96.12 ; 
      RECT 27.596 91.746 27.7 96.12 ; 
      RECT 27.164 91.746 27.268 96.12 ; 
      RECT 26.732 91.746 26.836 96.12 ; 
      RECT 26.3 91.746 26.404 96.12 ; 
      RECT 25.868 91.746 25.972 96.12 ; 
      RECT 25.436 91.746 25.54 96.12 ; 
      RECT 25.004 91.746 25.108 96.12 ; 
      RECT 24.572 91.746 24.676 96.12 ; 
      RECT 24.14 91.746 24.244 96.12 ; 
      RECT 23.708 91.746 23.812 96.12 ; 
      RECT 22.856 91.746 23.164 96.12 ; 
      RECT 15.284 91.746 15.592 96.12 ; 
      RECT 14.636 91.746 14.74 96.12 ; 
      RECT 14.204 91.746 14.308 96.12 ; 
      RECT 13.772 91.746 13.876 96.12 ; 
      RECT 13.34 91.746 13.444 96.12 ; 
      RECT 12.908 91.746 13.012 96.12 ; 
      RECT 12.476 91.746 12.58 96.12 ; 
      RECT 12.044 91.746 12.148 96.12 ; 
      RECT 11.612 91.746 11.716 96.12 ; 
      RECT 11.18 91.746 11.284 96.12 ; 
      RECT 10.748 91.746 10.852 96.12 ; 
      RECT 10.316 91.746 10.42 96.12 ; 
      RECT 9.884 91.746 9.988 96.12 ; 
      RECT 9.452 91.746 9.556 96.12 ; 
      RECT 9.02 91.746 9.124 96.12 ; 
      RECT 8.588 91.746 8.692 96.12 ; 
      RECT 8.156 91.746 8.26 96.12 ; 
      RECT 7.724 91.746 7.828 96.12 ; 
      RECT 7.292 91.746 7.396 96.12 ; 
      RECT 6.86 91.746 6.964 96.12 ; 
      RECT 6.428 91.746 6.532 96.12 ; 
      RECT 5.996 91.746 6.1 96.12 ; 
      RECT 5.564 91.746 5.668 96.12 ; 
      RECT 5.132 91.746 5.236 96.12 ; 
      RECT 4.7 91.746 4.804 96.12 ; 
      RECT 4.268 91.746 4.372 96.12 ; 
      RECT 3.836 91.746 3.94 96.12 ; 
      RECT 3.404 91.746 3.508 96.12 ; 
      RECT 2.972 91.746 3.076 96.12 ; 
      RECT 2.54 91.746 2.644 96.12 ; 
      RECT 2.108 91.746 2.212 96.12 ; 
      RECT 1.676 91.746 1.78 96.12 ; 
      RECT 1.244 91.746 1.348 96.12 ; 
      RECT 0.812 91.746 0.916 96.12 ; 
      RECT 0 91.746 0.34 96.12 ; 
      RECT 20.72 96.066 21.232 100.44 ; 
      RECT 20.664 98.728 21.232 100.018 ; 
      RECT 20.072 97.636 20.32 100.44 ; 
      RECT 20.016 98.874 20.32 99.488 ; 
      RECT 20.072 96.066 20.176 100.44 ; 
      RECT 20.072 96.55 20.232 97.508 ; 
      RECT 20.072 96.066 20.32 96.422 ; 
      RECT 18.884 97.868 19.708 100.44 ; 
      RECT 19.604 96.066 19.708 100.44 ; 
      RECT 18.884 98.976 19.764 100.008 ; 
      RECT 18.884 96.066 19.276 100.44 ; 
      RECT 17.216 96.066 17.548 100.44 ; 
      RECT 17.216 96.42 17.604 100.162 ; 
      RECT 38.108 96.066 38.448 100.44 ; 
      RECT 37.532 96.066 37.636 100.44 ; 
      RECT 37.1 96.066 37.204 100.44 ; 
      RECT 36.668 96.066 36.772 100.44 ; 
      RECT 36.236 96.066 36.34 100.44 ; 
      RECT 35.804 96.066 35.908 100.44 ; 
      RECT 35.372 96.066 35.476 100.44 ; 
      RECT 34.94 96.066 35.044 100.44 ; 
      RECT 34.508 96.066 34.612 100.44 ; 
      RECT 34.076 96.066 34.18 100.44 ; 
      RECT 33.644 96.066 33.748 100.44 ; 
      RECT 33.212 96.066 33.316 100.44 ; 
      RECT 32.78 96.066 32.884 100.44 ; 
      RECT 32.348 96.066 32.452 100.44 ; 
      RECT 31.916 96.066 32.02 100.44 ; 
      RECT 31.484 96.066 31.588 100.44 ; 
      RECT 31.052 96.066 31.156 100.44 ; 
      RECT 30.62 96.066 30.724 100.44 ; 
      RECT 30.188 96.066 30.292 100.44 ; 
      RECT 29.756 96.066 29.86 100.44 ; 
      RECT 29.324 96.066 29.428 100.44 ; 
      RECT 28.892 96.066 28.996 100.44 ; 
      RECT 28.46 96.066 28.564 100.44 ; 
      RECT 28.028 96.066 28.132 100.44 ; 
      RECT 27.596 96.066 27.7 100.44 ; 
      RECT 27.164 96.066 27.268 100.44 ; 
      RECT 26.732 96.066 26.836 100.44 ; 
      RECT 26.3 96.066 26.404 100.44 ; 
      RECT 25.868 96.066 25.972 100.44 ; 
      RECT 25.436 96.066 25.54 100.44 ; 
      RECT 25.004 96.066 25.108 100.44 ; 
      RECT 24.572 96.066 24.676 100.44 ; 
      RECT 24.14 96.066 24.244 100.44 ; 
      RECT 23.708 96.066 23.812 100.44 ; 
      RECT 22.856 96.066 23.164 100.44 ; 
      RECT 15.284 96.066 15.592 100.44 ; 
      RECT 14.636 96.066 14.74 100.44 ; 
      RECT 14.204 96.066 14.308 100.44 ; 
      RECT 13.772 96.066 13.876 100.44 ; 
      RECT 13.34 96.066 13.444 100.44 ; 
      RECT 12.908 96.066 13.012 100.44 ; 
      RECT 12.476 96.066 12.58 100.44 ; 
      RECT 12.044 96.066 12.148 100.44 ; 
      RECT 11.612 96.066 11.716 100.44 ; 
      RECT 11.18 96.066 11.284 100.44 ; 
      RECT 10.748 96.066 10.852 100.44 ; 
      RECT 10.316 96.066 10.42 100.44 ; 
      RECT 9.884 96.066 9.988 100.44 ; 
      RECT 9.452 96.066 9.556 100.44 ; 
      RECT 9.02 96.066 9.124 100.44 ; 
      RECT 8.588 96.066 8.692 100.44 ; 
      RECT 8.156 96.066 8.26 100.44 ; 
      RECT 7.724 96.066 7.828 100.44 ; 
      RECT 7.292 96.066 7.396 100.44 ; 
      RECT 6.86 96.066 6.964 100.44 ; 
      RECT 6.428 96.066 6.532 100.44 ; 
      RECT 5.996 96.066 6.1 100.44 ; 
      RECT 5.564 96.066 5.668 100.44 ; 
      RECT 5.132 96.066 5.236 100.44 ; 
      RECT 4.7 96.066 4.804 100.44 ; 
      RECT 4.268 96.066 4.372 100.44 ; 
      RECT 3.836 96.066 3.94 100.44 ; 
      RECT 3.404 96.066 3.508 100.44 ; 
      RECT 2.972 96.066 3.076 100.44 ; 
      RECT 2.54 96.066 2.644 100.44 ; 
      RECT 2.108 96.066 2.212 100.44 ; 
      RECT 1.676 96.066 1.78 100.44 ; 
      RECT 1.244 96.066 1.348 100.44 ; 
      RECT 0.812 96.066 0.916 100.44 ; 
      RECT 0 96.066 0.34 100.44 ; 
      RECT 20.72 100.386 21.232 104.76 ; 
      RECT 20.664 103.048 21.232 104.338 ; 
      RECT 20.072 101.956 20.32 104.76 ; 
      RECT 20.016 103.194 20.32 103.808 ; 
      RECT 20.072 100.386 20.176 104.76 ; 
      RECT 20.072 100.87 20.232 101.828 ; 
      RECT 20.072 100.386 20.32 100.742 ; 
      RECT 18.884 102.188 19.708 104.76 ; 
      RECT 19.604 100.386 19.708 104.76 ; 
      RECT 18.884 103.296 19.764 104.328 ; 
      RECT 18.884 100.386 19.276 104.76 ; 
      RECT 17.216 100.386 17.548 104.76 ; 
      RECT 17.216 100.74 17.604 104.482 ; 
      RECT 38.108 100.386 38.448 104.76 ; 
      RECT 37.532 100.386 37.636 104.76 ; 
      RECT 37.1 100.386 37.204 104.76 ; 
      RECT 36.668 100.386 36.772 104.76 ; 
      RECT 36.236 100.386 36.34 104.76 ; 
      RECT 35.804 100.386 35.908 104.76 ; 
      RECT 35.372 100.386 35.476 104.76 ; 
      RECT 34.94 100.386 35.044 104.76 ; 
      RECT 34.508 100.386 34.612 104.76 ; 
      RECT 34.076 100.386 34.18 104.76 ; 
      RECT 33.644 100.386 33.748 104.76 ; 
      RECT 33.212 100.386 33.316 104.76 ; 
      RECT 32.78 100.386 32.884 104.76 ; 
      RECT 32.348 100.386 32.452 104.76 ; 
      RECT 31.916 100.386 32.02 104.76 ; 
      RECT 31.484 100.386 31.588 104.76 ; 
      RECT 31.052 100.386 31.156 104.76 ; 
      RECT 30.62 100.386 30.724 104.76 ; 
      RECT 30.188 100.386 30.292 104.76 ; 
      RECT 29.756 100.386 29.86 104.76 ; 
      RECT 29.324 100.386 29.428 104.76 ; 
      RECT 28.892 100.386 28.996 104.76 ; 
      RECT 28.46 100.386 28.564 104.76 ; 
      RECT 28.028 100.386 28.132 104.76 ; 
      RECT 27.596 100.386 27.7 104.76 ; 
      RECT 27.164 100.386 27.268 104.76 ; 
      RECT 26.732 100.386 26.836 104.76 ; 
      RECT 26.3 100.386 26.404 104.76 ; 
      RECT 25.868 100.386 25.972 104.76 ; 
      RECT 25.436 100.386 25.54 104.76 ; 
      RECT 25.004 100.386 25.108 104.76 ; 
      RECT 24.572 100.386 24.676 104.76 ; 
      RECT 24.14 100.386 24.244 104.76 ; 
      RECT 23.708 100.386 23.812 104.76 ; 
      RECT 22.856 100.386 23.164 104.76 ; 
      RECT 15.284 100.386 15.592 104.76 ; 
      RECT 14.636 100.386 14.74 104.76 ; 
      RECT 14.204 100.386 14.308 104.76 ; 
      RECT 13.772 100.386 13.876 104.76 ; 
      RECT 13.34 100.386 13.444 104.76 ; 
      RECT 12.908 100.386 13.012 104.76 ; 
      RECT 12.476 100.386 12.58 104.76 ; 
      RECT 12.044 100.386 12.148 104.76 ; 
      RECT 11.612 100.386 11.716 104.76 ; 
      RECT 11.18 100.386 11.284 104.76 ; 
      RECT 10.748 100.386 10.852 104.76 ; 
      RECT 10.316 100.386 10.42 104.76 ; 
      RECT 9.884 100.386 9.988 104.76 ; 
      RECT 9.452 100.386 9.556 104.76 ; 
      RECT 9.02 100.386 9.124 104.76 ; 
      RECT 8.588 100.386 8.692 104.76 ; 
      RECT 8.156 100.386 8.26 104.76 ; 
      RECT 7.724 100.386 7.828 104.76 ; 
      RECT 7.292 100.386 7.396 104.76 ; 
      RECT 6.86 100.386 6.964 104.76 ; 
      RECT 6.428 100.386 6.532 104.76 ; 
      RECT 5.996 100.386 6.1 104.76 ; 
      RECT 5.564 100.386 5.668 104.76 ; 
      RECT 5.132 100.386 5.236 104.76 ; 
      RECT 4.7 100.386 4.804 104.76 ; 
      RECT 4.268 100.386 4.372 104.76 ; 
      RECT 3.836 100.386 3.94 104.76 ; 
      RECT 3.404 100.386 3.508 104.76 ; 
      RECT 2.972 100.386 3.076 104.76 ; 
      RECT 2.54 100.386 2.644 104.76 ; 
      RECT 2.108 100.386 2.212 104.76 ; 
      RECT 1.676 100.386 1.78 104.76 ; 
      RECT 1.244 100.386 1.348 104.76 ; 
      RECT 0.812 100.386 0.916 104.76 ; 
      RECT 0 100.386 0.34 104.76 ; 
      RECT 20.72 104.706 21.232 109.08 ; 
      RECT 20.664 107.368 21.232 108.658 ; 
      RECT 20.072 106.276 20.32 109.08 ; 
      RECT 20.016 107.514 20.32 108.128 ; 
      RECT 20.072 104.706 20.176 109.08 ; 
      RECT 20.072 105.19 20.232 106.148 ; 
      RECT 20.072 104.706 20.32 105.062 ; 
      RECT 18.884 106.508 19.708 109.08 ; 
      RECT 19.604 104.706 19.708 109.08 ; 
      RECT 18.884 107.616 19.764 108.648 ; 
      RECT 18.884 104.706 19.276 109.08 ; 
      RECT 17.216 104.706 17.548 109.08 ; 
      RECT 17.216 105.06 17.604 108.802 ; 
      RECT 38.108 104.706 38.448 109.08 ; 
      RECT 37.532 104.706 37.636 109.08 ; 
      RECT 37.1 104.706 37.204 109.08 ; 
      RECT 36.668 104.706 36.772 109.08 ; 
      RECT 36.236 104.706 36.34 109.08 ; 
      RECT 35.804 104.706 35.908 109.08 ; 
      RECT 35.372 104.706 35.476 109.08 ; 
      RECT 34.94 104.706 35.044 109.08 ; 
      RECT 34.508 104.706 34.612 109.08 ; 
      RECT 34.076 104.706 34.18 109.08 ; 
      RECT 33.644 104.706 33.748 109.08 ; 
      RECT 33.212 104.706 33.316 109.08 ; 
      RECT 32.78 104.706 32.884 109.08 ; 
      RECT 32.348 104.706 32.452 109.08 ; 
      RECT 31.916 104.706 32.02 109.08 ; 
      RECT 31.484 104.706 31.588 109.08 ; 
      RECT 31.052 104.706 31.156 109.08 ; 
      RECT 30.62 104.706 30.724 109.08 ; 
      RECT 30.188 104.706 30.292 109.08 ; 
      RECT 29.756 104.706 29.86 109.08 ; 
      RECT 29.324 104.706 29.428 109.08 ; 
      RECT 28.892 104.706 28.996 109.08 ; 
      RECT 28.46 104.706 28.564 109.08 ; 
      RECT 28.028 104.706 28.132 109.08 ; 
      RECT 27.596 104.706 27.7 109.08 ; 
      RECT 27.164 104.706 27.268 109.08 ; 
      RECT 26.732 104.706 26.836 109.08 ; 
      RECT 26.3 104.706 26.404 109.08 ; 
      RECT 25.868 104.706 25.972 109.08 ; 
      RECT 25.436 104.706 25.54 109.08 ; 
      RECT 25.004 104.706 25.108 109.08 ; 
      RECT 24.572 104.706 24.676 109.08 ; 
      RECT 24.14 104.706 24.244 109.08 ; 
      RECT 23.708 104.706 23.812 109.08 ; 
      RECT 22.856 104.706 23.164 109.08 ; 
      RECT 15.284 104.706 15.592 109.08 ; 
      RECT 14.636 104.706 14.74 109.08 ; 
      RECT 14.204 104.706 14.308 109.08 ; 
      RECT 13.772 104.706 13.876 109.08 ; 
      RECT 13.34 104.706 13.444 109.08 ; 
      RECT 12.908 104.706 13.012 109.08 ; 
      RECT 12.476 104.706 12.58 109.08 ; 
      RECT 12.044 104.706 12.148 109.08 ; 
      RECT 11.612 104.706 11.716 109.08 ; 
      RECT 11.18 104.706 11.284 109.08 ; 
      RECT 10.748 104.706 10.852 109.08 ; 
      RECT 10.316 104.706 10.42 109.08 ; 
      RECT 9.884 104.706 9.988 109.08 ; 
      RECT 9.452 104.706 9.556 109.08 ; 
      RECT 9.02 104.706 9.124 109.08 ; 
      RECT 8.588 104.706 8.692 109.08 ; 
      RECT 8.156 104.706 8.26 109.08 ; 
      RECT 7.724 104.706 7.828 109.08 ; 
      RECT 7.292 104.706 7.396 109.08 ; 
      RECT 6.86 104.706 6.964 109.08 ; 
      RECT 6.428 104.706 6.532 109.08 ; 
      RECT 5.996 104.706 6.1 109.08 ; 
      RECT 5.564 104.706 5.668 109.08 ; 
      RECT 5.132 104.706 5.236 109.08 ; 
      RECT 4.7 104.706 4.804 109.08 ; 
      RECT 4.268 104.706 4.372 109.08 ; 
      RECT 3.836 104.706 3.94 109.08 ; 
      RECT 3.404 104.706 3.508 109.08 ; 
      RECT 2.972 104.706 3.076 109.08 ; 
      RECT 2.54 104.706 2.644 109.08 ; 
      RECT 2.108 104.706 2.212 109.08 ; 
      RECT 1.676 104.706 1.78 109.08 ; 
      RECT 1.244 104.706 1.348 109.08 ; 
      RECT 0.812 104.706 0.916 109.08 ; 
      RECT 0 104.706 0.34 109.08 ; 
      RECT 20.72 109.026 21.232 113.4 ; 
      RECT 20.664 111.688 21.232 112.978 ; 
      RECT 20.072 110.596 20.32 113.4 ; 
      RECT 20.016 111.834 20.32 112.448 ; 
      RECT 20.072 109.026 20.176 113.4 ; 
      RECT 20.072 109.51 20.232 110.468 ; 
      RECT 20.072 109.026 20.32 109.382 ; 
      RECT 18.884 110.828 19.708 113.4 ; 
      RECT 19.604 109.026 19.708 113.4 ; 
      RECT 18.884 111.936 19.764 112.968 ; 
      RECT 18.884 109.026 19.276 113.4 ; 
      RECT 17.216 109.026 17.548 113.4 ; 
      RECT 17.216 109.38 17.604 113.122 ; 
      RECT 38.108 109.026 38.448 113.4 ; 
      RECT 37.532 109.026 37.636 113.4 ; 
      RECT 37.1 109.026 37.204 113.4 ; 
      RECT 36.668 109.026 36.772 113.4 ; 
      RECT 36.236 109.026 36.34 113.4 ; 
      RECT 35.804 109.026 35.908 113.4 ; 
      RECT 35.372 109.026 35.476 113.4 ; 
      RECT 34.94 109.026 35.044 113.4 ; 
      RECT 34.508 109.026 34.612 113.4 ; 
      RECT 34.076 109.026 34.18 113.4 ; 
      RECT 33.644 109.026 33.748 113.4 ; 
      RECT 33.212 109.026 33.316 113.4 ; 
      RECT 32.78 109.026 32.884 113.4 ; 
      RECT 32.348 109.026 32.452 113.4 ; 
      RECT 31.916 109.026 32.02 113.4 ; 
      RECT 31.484 109.026 31.588 113.4 ; 
      RECT 31.052 109.026 31.156 113.4 ; 
      RECT 30.62 109.026 30.724 113.4 ; 
      RECT 30.188 109.026 30.292 113.4 ; 
      RECT 29.756 109.026 29.86 113.4 ; 
      RECT 29.324 109.026 29.428 113.4 ; 
      RECT 28.892 109.026 28.996 113.4 ; 
      RECT 28.46 109.026 28.564 113.4 ; 
      RECT 28.028 109.026 28.132 113.4 ; 
      RECT 27.596 109.026 27.7 113.4 ; 
      RECT 27.164 109.026 27.268 113.4 ; 
      RECT 26.732 109.026 26.836 113.4 ; 
      RECT 26.3 109.026 26.404 113.4 ; 
      RECT 25.868 109.026 25.972 113.4 ; 
      RECT 25.436 109.026 25.54 113.4 ; 
      RECT 25.004 109.026 25.108 113.4 ; 
      RECT 24.572 109.026 24.676 113.4 ; 
      RECT 24.14 109.026 24.244 113.4 ; 
      RECT 23.708 109.026 23.812 113.4 ; 
      RECT 22.856 109.026 23.164 113.4 ; 
      RECT 15.284 109.026 15.592 113.4 ; 
      RECT 14.636 109.026 14.74 113.4 ; 
      RECT 14.204 109.026 14.308 113.4 ; 
      RECT 13.772 109.026 13.876 113.4 ; 
      RECT 13.34 109.026 13.444 113.4 ; 
      RECT 12.908 109.026 13.012 113.4 ; 
      RECT 12.476 109.026 12.58 113.4 ; 
      RECT 12.044 109.026 12.148 113.4 ; 
      RECT 11.612 109.026 11.716 113.4 ; 
      RECT 11.18 109.026 11.284 113.4 ; 
      RECT 10.748 109.026 10.852 113.4 ; 
      RECT 10.316 109.026 10.42 113.4 ; 
      RECT 9.884 109.026 9.988 113.4 ; 
      RECT 9.452 109.026 9.556 113.4 ; 
      RECT 9.02 109.026 9.124 113.4 ; 
      RECT 8.588 109.026 8.692 113.4 ; 
      RECT 8.156 109.026 8.26 113.4 ; 
      RECT 7.724 109.026 7.828 113.4 ; 
      RECT 7.292 109.026 7.396 113.4 ; 
      RECT 6.86 109.026 6.964 113.4 ; 
      RECT 6.428 109.026 6.532 113.4 ; 
      RECT 5.996 109.026 6.1 113.4 ; 
      RECT 5.564 109.026 5.668 113.4 ; 
      RECT 5.132 109.026 5.236 113.4 ; 
      RECT 4.7 109.026 4.804 113.4 ; 
      RECT 4.268 109.026 4.372 113.4 ; 
      RECT 3.836 109.026 3.94 113.4 ; 
      RECT 3.404 109.026 3.508 113.4 ; 
      RECT 2.972 109.026 3.076 113.4 ; 
      RECT 2.54 109.026 2.644 113.4 ; 
      RECT 2.108 109.026 2.212 113.4 ; 
      RECT 1.676 109.026 1.78 113.4 ; 
      RECT 1.244 109.026 1.348 113.4 ; 
      RECT 0.812 109.026 0.916 113.4 ; 
      RECT 0 109.026 0.34 113.4 ; 
      RECT 20.72 113.346 21.232 117.72 ; 
      RECT 20.664 116.008 21.232 117.298 ; 
      RECT 20.072 114.916 20.32 117.72 ; 
      RECT 20.016 116.154 20.32 116.768 ; 
      RECT 20.072 113.346 20.176 117.72 ; 
      RECT 20.072 113.83 20.232 114.788 ; 
      RECT 20.072 113.346 20.32 113.702 ; 
      RECT 18.884 115.148 19.708 117.72 ; 
      RECT 19.604 113.346 19.708 117.72 ; 
      RECT 18.884 116.256 19.764 117.288 ; 
      RECT 18.884 113.346 19.276 117.72 ; 
      RECT 17.216 113.346 17.548 117.72 ; 
      RECT 17.216 113.7 17.604 117.442 ; 
      RECT 38.108 113.346 38.448 117.72 ; 
      RECT 37.532 113.346 37.636 117.72 ; 
      RECT 37.1 113.346 37.204 117.72 ; 
      RECT 36.668 113.346 36.772 117.72 ; 
      RECT 36.236 113.346 36.34 117.72 ; 
      RECT 35.804 113.346 35.908 117.72 ; 
      RECT 35.372 113.346 35.476 117.72 ; 
      RECT 34.94 113.346 35.044 117.72 ; 
      RECT 34.508 113.346 34.612 117.72 ; 
      RECT 34.076 113.346 34.18 117.72 ; 
      RECT 33.644 113.346 33.748 117.72 ; 
      RECT 33.212 113.346 33.316 117.72 ; 
      RECT 32.78 113.346 32.884 117.72 ; 
      RECT 32.348 113.346 32.452 117.72 ; 
      RECT 31.916 113.346 32.02 117.72 ; 
      RECT 31.484 113.346 31.588 117.72 ; 
      RECT 31.052 113.346 31.156 117.72 ; 
      RECT 30.62 113.346 30.724 117.72 ; 
      RECT 30.188 113.346 30.292 117.72 ; 
      RECT 29.756 113.346 29.86 117.72 ; 
      RECT 29.324 113.346 29.428 117.72 ; 
      RECT 28.892 113.346 28.996 117.72 ; 
      RECT 28.46 113.346 28.564 117.72 ; 
      RECT 28.028 113.346 28.132 117.72 ; 
      RECT 27.596 113.346 27.7 117.72 ; 
      RECT 27.164 113.346 27.268 117.72 ; 
      RECT 26.732 113.346 26.836 117.72 ; 
      RECT 26.3 113.346 26.404 117.72 ; 
      RECT 25.868 113.346 25.972 117.72 ; 
      RECT 25.436 113.346 25.54 117.72 ; 
      RECT 25.004 113.346 25.108 117.72 ; 
      RECT 24.572 113.346 24.676 117.72 ; 
      RECT 24.14 113.346 24.244 117.72 ; 
      RECT 23.708 113.346 23.812 117.72 ; 
      RECT 22.856 113.346 23.164 117.72 ; 
      RECT 15.284 113.346 15.592 117.72 ; 
      RECT 14.636 113.346 14.74 117.72 ; 
      RECT 14.204 113.346 14.308 117.72 ; 
      RECT 13.772 113.346 13.876 117.72 ; 
      RECT 13.34 113.346 13.444 117.72 ; 
      RECT 12.908 113.346 13.012 117.72 ; 
      RECT 12.476 113.346 12.58 117.72 ; 
      RECT 12.044 113.346 12.148 117.72 ; 
      RECT 11.612 113.346 11.716 117.72 ; 
      RECT 11.18 113.346 11.284 117.72 ; 
      RECT 10.748 113.346 10.852 117.72 ; 
      RECT 10.316 113.346 10.42 117.72 ; 
      RECT 9.884 113.346 9.988 117.72 ; 
      RECT 9.452 113.346 9.556 117.72 ; 
      RECT 9.02 113.346 9.124 117.72 ; 
      RECT 8.588 113.346 8.692 117.72 ; 
      RECT 8.156 113.346 8.26 117.72 ; 
      RECT 7.724 113.346 7.828 117.72 ; 
      RECT 7.292 113.346 7.396 117.72 ; 
      RECT 6.86 113.346 6.964 117.72 ; 
      RECT 6.428 113.346 6.532 117.72 ; 
      RECT 5.996 113.346 6.1 117.72 ; 
      RECT 5.564 113.346 5.668 117.72 ; 
      RECT 5.132 113.346 5.236 117.72 ; 
      RECT 4.7 113.346 4.804 117.72 ; 
      RECT 4.268 113.346 4.372 117.72 ; 
      RECT 3.836 113.346 3.94 117.72 ; 
      RECT 3.404 113.346 3.508 117.72 ; 
      RECT 2.972 113.346 3.076 117.72 ; 
      RECT 2.54 113.346 2.644 117.72 ; 
      RECT 2.108 113.346 2.212 117.72 ; 
      RECT 1.676 113.346 1.78 117.72 ; 
      RECT 1.244 113.346 1.348 117.72 ; 
      RECT 0.812 113.346 0.916 117.72 ; 
      RECT 0 113.346 0.34 117.72 ; 
      RECT 20.72 117.666 21.232 122.04 ; 
      RECT 20.664 120.328 21.232 121.618 ; 
      RECT 20.072 119.236 20.32 122.04 ; 
      RECT 20.016 120.474 20.32 121.088 ; 
      RECT 20.072 117.666 20.176 122.04 ; 
      RECT 20.072 118.15 20.232 119.108 ; 
      RECT 20.072 117.666 20.32 118.022 ; 
      RECT 18.884 119.468 19.708 122.04 ; 
      RECT 19.604 117.666 19.708 122.04 ; 
      RECT 18.884 120.576 19.764 121.608 ; 
      RECT 18.884 117.666 19.276 122.04 ; 
      RECT 17.216 117.666 17.548 122.04 ; 
      RECT 17.216 118.02 17.604 121.762 ; 
      RECT 38.108 117.666 38.448 122.04 ; 
      RECT 37.532 117.666 37.636 122.04 ; 
      RECT 37.1 117.666 37.204 122.04 ; 
      RECT 36.668 117.666 36.772 122.04 ; 
      RECT 36.236 117.666 36.34 122.04 ; 
      RECT 35.804 117.666 35.908 122.04 ; 
      RECT 35.372 117.666 35.476 122.04 ; 
      RECT 34.94 117.666 35.044 122.04 ; 
      RECT 34.508 117.666 34.612 122.04 ; 
      RECT 34.076 117.666 34.18 122.04 ; 
      RECT 33.644 117.666 33.748 122.04 ; 
      RECT 33.212 117.666 33.316 122.04 ; 
      RECT 32.78 117.666 32.884 122.04 ; 
      RECT 32.348 117.666 32.452 122.04 ; 
      RECT 31.916 117.666 32.02 122.04 ; 
      RECT 31.484 117.666 31.588 122.04 ; 
      RECT 31.052 117.666 31.156 122.04 ; 
      RECT 30.62 117.666 30.724 122.04 ; 
      RECT 30.188 117.666 30.292 122.04 ; 
      RECT 29.756 117.666 29.86 122.04 ; 
      RECT 29.324 117.666 29.428 122.04 ; 
      RECT 28.892 117.666 28.996 122.04 ; 
      RECT 28.46 117.666 28.564 122.04 ; 
      RECT 28.028 117.666 28.132 122.04 ; 
      RECT 27.596 117.666 27.7 122.04 ; 
      RECT 27.164 117.666 27.268 122.04 ; 
      RECT 26.732 117.666 26.836 122.04 ; 
      RECT 26.3 117.666 26.404 122.04 ; 
      RECT 25.868 117.666 25.972 122.04 ; 
      RECT 25.436 117.666 25.54 122.04 ; 
      RECT 25.004 117.666 25.108 122.04 ; 
      RECT 24.572 117.666 24.676 122.04 ; 
      RECT 24.14 117.666 24.244 122.04 ; 
      RECT 23.708 117.666 23.812 122.04 ; 
      RECT 22.856 117.666 23.164 122.04 ; 
      RECT 15.284 117.666 15.592 122.04 ; 
      RECT 14.636 117.666 14.74 122.04 ; 
      RECT 14.204 117.666 14.308 122.04 ; 
      RECT 13.772 117.666 13.876 122.04 ; 
      RECT 13.34 117.666 13.444 122.04 ; 
      RECT 12.908 117.666 13.012 122.04 ; 
      RECT 12.476 117.666 12.58 122.04 ; 
      RECT 12.044 117.666 12.148 122.04 ; 
      RECT 11.612 117.666 11.716 122.04 ; 
      RECT 11.18 117.666 11.284 122.04 ; 
      RECT 10.748 117.666 10.852 122.04 ; 
      RECT 10.316 117.666 10.42 122.04 ; 
      RECT 9.884 117.666 9.988 122.04 ; 
      RECT 9.452 117.666 9.556 122.04 ; 
      RECT 9.02 117.666 9.124 122.04 ; 
      RECT 8.588 117.666 8.692 122.04 ; 
      RECT 8.156 117.666 8.26 122.04 ; 
      RECT 7.724 117.666 7.828 122.04 ; 
      RECT 7.292 117.666 7.396 122.04 ; 
      RECT 6.86 117.666 6.964 122.04 ; 
      RECT 6.428 117.666 6.532 122.04 ; 
      RECT 5.996 117.666 6.1 122.04 ; 
      RECT 5.564 117.666 5.668 122.04 ; 
      RECT 5.132 117.666 5.236 122.04 ; 
      RECT 4.7 117.666 4.804 122.04 ; 
      RECT 4.268 117.666 4.372 122.04 ; 
      RECT 3.836 117.666 3.94 122.04 ; 
      RECT 3.404 117.666 3.508 122.04 ; 
      RECT 2.972 117.666 3.076 122.04 ; 
      RECT 2.54 117.666 2.644 122.04 ; 
      RECT 2.108 117.666 2.212 122.04 ; 
      RECT 1.676 117.666 1.78 122.04 ; 
      RECT 1.244 117.666 1.348 122.04 ; 
      RECT 0.812 117.666 0.916 122.04 ; 
      RECT 0 117.666 0.34 122.04 ; 
      RECT 20.72 121.986 21.232 126.36 ; 
      RECT 20.664 124.648 21.232 125.938 ; 
      RECT 20.072 123.556 20.32 126.36 ; 
      RECT 20.016 124.794 20.32 125.408 ; 
      RECT 20.072 121.986 20.176 126.36 ; 
      RECT 20.072 122.47 20.232 123.428 ; 
      RECT 20.072 121.986 20.32 122.342 ; 
      RECT 18.884 123.788 19.708 126.36 ; 
      RECT 19.604 121.986 19.708 126.36 ; 
      RECT 18.884 124.896 19.764 125.928 ; 
      RECT 18.884 121.986 19.276 126.36 ; 
      RECT 17.216 121.986 17.548 126.36 ; 
      RECT 17.216 122.34 17.604 126.082 ; 
      RECT 38.108 121.986 38.448 126.36 ; 
      RECT 37.532 121.986 37.636 126.36 ; 
      RECT 37.1 121.986 37.204 126.36 ; 
      RECT 36.668 121.986 36.772 126.36 ; 
      RECT 36.236 121.986 36.34 126.36 ; 
      RECT 35.804 121.986 35.908 126.36 ; 
      RECT 35.372 121.986 35.476 126.36 ; 
      RECT 34.94 121.986 35.044 126.36 ; 
      RECT 34.508 121.986 34.612 126.36 ; 
      RECT 34.076 121.986 34.18 126.36 ; 
      RECT 33.644 121.986 33.748 126.36 ; 
      RECT 33.212 121.986 33.316 126.36 ; 
      RECT 32.78 121.986 32.884 126.36 ; 
      RECT 32.348 121.986 32.452 126.36 ; 
      RECT 31.916 121.986 32.02 126.36 ; 
      RECT 31.484 121.986 31.588 126.36 ; 
      RECT 31.052 121.986 31.156 126.36 ; 
      RECT 30.62 121.986 30.724 126.36 ; 
      RECT 30.188 121.986 30.292 126.36 ; 
      RECT 29.756 121.986 29.86 126.36 ; 
      RECT 29.324 121.986 29.428 126.36 ; 
      RECT 28.892 121.986 28.996 126.36 ; 
      RECT 28.46 121.986 28.564 126.36 ; 
      RECT 28.028 121.986 28.132 126.36 ; 
      RECT 27.596 121.986 27.7 126.36 ; 
      RECT 27.164 121.986 27.268 126.36 ; 
      RECT 26.732 121.986 26.836 126.36 ; 
      RECT 26.3 121.986 26.404 126.36 ; 
      RECT 25.868 121.986 25.972 126.36 ; 
      RECT 25.436 121.986 25.54 126.36 ; 
      RECT 25.004 121.986 25.108 126.36 ; 
      RECT 24.572 121.986 24.676 126.36 ; 
      RECT 24.14 121.986 24.244 126.36 ; 
      RECT 23.708 121.986 23.812 126.36 ; 
      RECT 22.856 121.986 23.164 126.36 ; 
      RECT 15.284 121.986 15.592 126.36 ; 
      RECT 14.636 121.986 14.74 126.36 ; 
      RECT 14.204 121.986 14.308 126.36 ; 
      RECT 13.772 121.986 13.876 126.36 ; 
      RECT 13.34 121.986 13.444 126.36 ; 
      RECT 12.908 121.986 13.012 126.36 ; 
      RECT 12.476 121.986 12.58 126.36 ; 
      RECT 12.044 121.986 12.148 126.36 ; 
      RECT 11.612 121.986 11.716 126.36 ; 
      RECT 11.18 121.986 11.284 126.36 ; 
      RECT 10.748 121.986 10.852 126.36 ; 
      RECT 10.316 121.986 10.42 126.36 ; 
      RECT 9.884 121.986 9.988 126.36 ; 
      RECT 9.452 121.986 9.556 126.36 ; 
      RECT 9.02 121.986 9.124 126.36 ; 
      RECT 8.588 121.986 8.692 126.36 ; 
      RECT 8.156 121.986 8.26 126.36 ; 
      RECT 7.724 121.986 7.828 126.36 ; 
      RECT 7.292 121.986 7.396 126.36 ; 
      RECT 6.86 121.986 6.964 126.36 ; 
      RECT 6.428 121.986 6.532 126.36 ; 
      RECT 5.996 121.986 6.1 126.36 ; 
      RECT 5.564 121.986 5.668 126.36 ; 
      RECT 5.132 121.986 5.236 126.36 ; 
      RECT 4.7 121.986 4.804 126.36 ; 
      RECT 4.268 121.986 4.372 126.36 ; 
      RECT 3.836 121.986 3.94 126.36 ; 
      RECT 3.404 121.986 3.508 126.36 ; 
      RECT 2.972 121.986 3.076 126.36 ; 
      RECT 2.54 121.986 2.644 126.36 ; 
      RECT 2.108 121.986 2.212 126.36 ; 
      RECT 1.676 121.986 1.78 126.36 ; 
      RECT 1.244 121.986 1.348 126.36 ; 
      RECT 0.812 121.986 0.916 126.36 ; 
      RECT 0 121.986 0.34 126.36 ; 
      RECT 20.72 126.306 21.232 130.68 ; 
      RECT 20.664 128.968 21.232 130.258 ; 
      RECT 20.072 127.876 20.32 130.68 ; 
      RECT 20.016 129.114 20.32 129.728 ; 
      RECT 20.072 126.306 20.176 130.68 ; 
      RECT 20.072 126.79 20.232 127.748 ; 
      RECT 20.072 126.306 20.32 126.662 ; 
      RECT 18.884 128.108 19.708 130.68 ; 
      RECT 19.604 126.306 19.708 130.68 ; 
      RECT 18.884 129.216 19.764 130.248 ; 
      RECT 18.884 126.306 19.276 130.68 ; 
      RECT 17.216 126.306 17.548 130.68 ; 
      RECT 17.216 126.66 17.604 130.402 ; 
      RECT 38.108 126.306 38.448 130.68 ; 
      RECT 37.532 126.306 37.636 130.68 ; 
      RECT 37.1 126.306 37.204 130.68 ; 
      RECT 36.668 126.306 36.772 130.68 ; 
      RECT 36.236 126.306 36.34 130.68 ; 
      RECT 35.804 126.306 35.908 130.68 ; 
      RECT 35.372 126.306 35.476 130.68 ; 
      RECT 34.94 126.306 35.044 130.68 ; 
      RECT 34.508 126.306 34.612 130.68 ; 
      RECT 34.076 126.306 34.18 130.68 ; 
      RECT 33.644 126.306 33.748 130.68 ; 
      RECT 33.212 126.306 33.316 130.68 ; 
      RECT 32.78 126.306 32.884 130.68 ; 
      RECT 32.348 126.306 32.452 130.68 ; 
      RECT 31.916 126.306 32.02 130.68 ; 
      RECT 31.484 126.306 31.588 130.68 ; 
      RECT 31.052 126.306 31.156 130.68 ; 
      RECT 30.62 126.306 30.724 130.68 ; 
      RECT 30.188 126.306 30.292 130.68 ; 
      RECT 29.756 126.306 29.86 130.68 ; 
      RECT 29.324 126.306 29.428 130.68 ; 
      RECT 28.892 126.306 28.996 130.68 ; 
      RECT 28.46 126.306 28.564 130.68 ; 
      RECT 28.028 126.306 28.132 130.68 ; 
      RECT 27.596 126.306 27.7 130.68 ; 
      RECT 27.164 126.306 27.268 130.68 ; 
      RECT 26.732 126.306 26.836 130.68 ; 
      RECT 26.3 126.306 26.404 130.68 ; 
      RECT 25.868 126.306 25.972 130.68 ; 
      RECT 25.436 126.306 25.54 130.68 ; 
      RECT 25.004 126.306 25.108 130.68 ; 
      RECT 24.572 126.306 24.676 130.68 ; 
      RECT 24.14 126.306 24.244 130.68 ; 
      RECT 23.708 126.306 23.812 130.68 ; 
      RECT 22.856 126.306 23.164 130.68 ; 
      RECT 15.284 126.306 15.592 130.68 ; 
      RECT 14.636 126.306 14.74 130.68 ; 
      RECT 14.204 126.306 14.308 130.68 ; 
      RECT 13.772 126.306 13.876 130.68 ; 
      RECT 13.34 126.306 13.444 130.68 ; 
      RECT 12.908 126.306 13.012 130.68 ; 
      RECT 12.476 126.306 12.58 130.68 ; 
      RECT 12.044 126.306 12.148 130.68 ; 
      RECT 11.612 126.306 11.716 130.68 ; 
      RECT 11.18 126.306 11.284 130.68 ; 
      RECT 10.748 126.306 10.852 130.68 ; 
      RECT 10.316 126.306 10.42 130.68 ; 
      RECT 9.884 126.306 9.988 130.68 ; 
      RECT 9.452 126.306 9.556 130.68 ; 
      RECT 9.02 126.306 9.124 130.68 ; 
      RECT 8.588 126.306 8.692 130.68 ; 
      RECT 8.156 126.306 8.26 130.68 ; 
      RECT 7.724 126.306 7.828 130.68 ; 
      RECT 7.292 126.306 7.396 130.68 ; 
      RECT 6.86 126.306 6.964 130.68 ; 
      RECT 6.428 126.306 6.532 130.68 ; 
      RECT 5.996 126.306 6.1 130.68 ; 
      RECT 5.564 126.306 5.668 130.68 ; 
      RECT 5.132 126.306 5.236 130.68 ; 
      RECT 4.7 126.306 4.804 130.68 ; 
      RECT 4.268 126.306 4.372 130.68 ; 
      RECT 3.836 126.306 3.94 130.68 ; 
      RECT 3.404 126.306 3.508 130.68 ; 
      RECT 2.972 126.306 3.076 130.68 ; 
      RECT 2.54 126.306 2.644 130.68 ; 
      RECT 2.108 126.306 2.212 130.68 ; 
      RECT 1.676 126.306 1.78 130.68 ; 
      RECT 1.244 126.306 1.348 130.68 ; 
      RECT 0.812 126.306 0.916 130.68 ; 
      RECT 0 126.306 0.34 130.68 ; 
      RECT 20.72 130.626 21.232 135 ; 
      RECT 20.664 133.288 21.232 134.578 ; 
      RECT 20.072 132.196 20.32 135 ; 
      RECT 20.016 133.434 20.32 134.048 ; 
      RECT 20.072 130.626 20.176 135 ; 
      RECT 20.072 131.11 20.232 132.068 ; 
      RECT 20.072 130.626 20.32 130.982 ; 
      RECT 18.884 132.428 19.708 135 ; 
      RECT 19.604 130.626 19.708 135 ; 
      RECT 18.884 133.536 19.764 134.568 ; 
      RECT 18.884 130.626 19.276 135 ; 
      RECT 17.216 130.626 17.548 135 ; 
      RECT 17.216 130.98 17.604 134.722 ; 
      RECT 38.108 130.626 38.448 135 ; 
      RECT 37.532 130.626 37.636 135 ; 
      RECT 37.1 130.626 37.204 135 ; 
      RECT 36.668 130.626 36.772 135 ; 
      RECT 36.236 130.626 36.34 135 ; 
      RECT 35.804 130.626 35.908 135 ; 
      RECT 35.372 130.626 35.476 135 ; 
      RECT 34.94 130.626 35.044 135 ; 
      RECT 34.508 130.626 34.612 135 ; 
      RECT 34.076 130.626 34.18 135 ; 
      RECT 33.644 130.626 33.748 135 ; 
      RECT 33.212 130.626 33.316 135 ; 
      RECT 32.78 130.626 32.884 135 ; 
      RECT 32.348 130.626 32.452 135 ; 
      RECT 31.916 130.626 32.02 135 ; 
      RECT 31.484 130.626 31.588 135 ; 
      RECT 31.052 130.626 31.156 135 ; 
      RECT 30.62 130.626 30.724 135 ; 
      RECT 30.188 130.626 30.292 135 ; 
      RECT 29.756 130.626 29.86 135 ; 
      RECT 29.324 130.626 29.428 135 ; 
      RECT 28.892 130.626 28.996 135 ; 
      RECT 28.46 130.626 28.564 135 ; 
      RECT 28.028 130.626 28.132 135 ; 
      RECT 27.596 130.626 27.7 135 ; 
      RECT 27.164 130.626 27.268 135 ; 
      RECT 26.732 130.626 26.836 135 ; 
      RECT 26.3 130.626 26.404 135 ; 
      RECT 25.868 130.626 25.972 135 ; 
      RECT 25.436 130.626 25.54 135 ; 
      RECT 25.004 130.626 25.108 135 ; 
      RECT 24.572 130.626 24.676 135 ; 
      RECT 24.14 130.626 24.244 135 ; 
      RECT 23.708 130.626 23.812 135 ; 
      RECT 22.856 130.626 23.164 135 ; 
      RECT 15.284 130.626 15.592 135 ; 
      RECT 14.636 130.626 14.74 135 ; 
      RECT 14.204 130.626 14.308 135 ; 
      RECT 13.772 130.626 13.876 135 ; 
      RECT 13.34 130.626 13.444 135 ; 
      RECT 12.908 130.626 13.012 135 ; 
      RECT 12.476 130.626 12.58 135 ; 
      RECT 12.044 130.626 12.148 135 ; 
      RECT 11.612 130.626 11.716 135 ; 
      RECT 11.18 130.626 11.284 135 ; 
      RECT 10.748 130.626 10.852 135 ; 
      RECT 10.316 130.626 10.42 135 ; 
      RECT 9.884 130.626 9.988 135 ; 
      RECT 9.452 130.626 9.556 135 ; 
      RECT 9.02 130.626 9.124 135 ; 
      RECT 8.588 130.626 8.692 135 ; 
      RECT 8.156 130.626 8.26 135 ; 
      RECT 7.724 130.626 7.828 135 ; 
      RECT 7.292 130.626 7.396 135 ; 
      RECT 6.86 130.626 6.964 135 ; 
      RECT 6.428 130.626 6.532 135 ; 
      RECT 5.996 130.626 6.1 135 ; 
      RECT 5.564 130.626 5.668 135 ; 
      RECT 5.132 130.626 5.236 135 ; 
      RECT 4.7 130.626 4.804 135 ; 
      RECT 4.268 130.626 4.372 135 ; 
      RECT 3.836 130.626 3.94 135 ; 
      RECT 3.404 130.626 3.508 135 ; 
      RECT 2.972 130.626 3.076 135 ; 
      RECT 2.54 130.626 2.644 135 ; 
      RECT 2.108 130.626 2.212 135 ; 
      RECT 1.676 130.626 1.78 135 ; 
      RECT 1.244 130.626 1.348 135 ; 
      RECT 0.812 130.626 0.916 135 ; 
      RECT 0 130.626 0.34 135 ; 
      RECT 20.72 134.946 21.232 139.32 ; 
      RECT 20.664 137.608 21.232 138.898 ; 
      RECT 20.072 136.516 20.32 139.32 ; 
      RECT 20.016 137.754 20.32 138.368 ; 
      RECT 20.072 134.946 20.176 139.32 ; 
      RECT 20.072 135.43 20.232 136.388 ; 
      RECT 20.072 134.946 20.32 135.302 ; 
      RECT 18.884 136.748 19.708 139.32 ; 
      RECT 19.604 134.946 19.708 139.32 ; 
      RECT 18.884 137.856 19.764 138.888 ; 
      RECT 18.884 134.946 19.276 139.32 ; 
      RECT 17.216 134.946 17.548 139.32 ; 
      RECT 17.216 135.3 17.604 139.042 ; 
      RECT 38.108 134.946 38.448 139.32 ; 
      RECT 37.532 134.946 37.636 139.32 ; 
      RECT 37.1 134.946 37.204 139.32 ; 
      RECT 36.668 134.946 36.772 139.32 ; 
      RECT 36.236 134.946 36.34 139.32 ; 
      RECT 35.804 134.946 35.908 139.32 ; 
      RECT 35.372 134.946 35.476 139.32 ; 
      RECT 34.94 134.946 35.044 139.32 ; 
      RECT 34.508 134.946 34.612 139.32 ; 
      RECT 34.076 134.946 34.18 139.32 ; 
      RECT 33.644 134.946 33.748 139.32 ; 
      RECT 33.212 134.946 33.316 139.32 ; 
      RECT 32.78 134.946 32.884 139.32 ; 
      RECT 32.348 134.946 32.452 139.32 ; 
      RECT 31.916 134.946 32.02 139.32 ; 
      RECT 31.484 134.946 31.588 139.32 ; 
      RECT 31.052 134.946 31.156 139.32 ; 
      RECT 30.62 134.946 30.724 139.32 ; 
      RECT 30.188 134.946 30.292 139.32 ; 
      RECT 29.756 134.946 29.86 139.32 ; 
      RECT 29.324 134.946 29.428 139.32 ; 
      RECT 28.892 134.946 28.996 139.32 ; 
      RECT 28.46 134.946 28.564 139.32 ; 
      RECT 28.028 134.946 28.132 139.32 ; 
      RECT 27.596 134.946 27.7 139.32 ; 
      RECT 27.164 134.946 27.268 139.32 ; 
      RECT 26.732 134.946 26.836 139.32 ; 
      RECT 26.3 134.946 26.404 139.32 ; 
      RECT 25.868 134.946 25.972 139.32 ; 
      RECT 25.436 134.946 25.54 139.32 ; 
      RECT 25.004 134.946 25.108 139.32 ; 
      RECT 24.572 134.946 24.676 139.32 ; 
      RECT 24.14 134.946 24.244 139.32 ; 
      RECT 23.708 134.946 23.812 139.32 ; 
      RECT 22.856 134.946 23.164 139.32 ; 
      RECT 15.284 134.946 15.592 139.32 ; 
      RECT 14.636 134.946 14.74 139.32 ; 
      RECT 14.204 134.946 14.308 139.32 ; 
      RECT 13.772 134.946 13.876 139.32 ; 
      RECT 13.34 134.946 13.444 139.32 ; 
      RECT 12.908 134.946 13.012 139.32 ; 
      RECT 12.476 134.946 12.58 139.32 ; 
      RECT 12.044 134.946 12.148 139.32 ; 
      RECT 11.612 134.946 11.716 139.32 ; 
      RECT 11.18 134.946 11.284 139.32 ; 
      RECT 10.748 134.946 10.852 139.32 ; 
      RECT 10.316 134.946 10.42 139.32 ; 
      RECT 9.884 134.946 9.988 139.32 ; 
      RECT 9.452 134.946 9.556 139.32 ; 
      RECT 9.02 134.946 9.124 139.32 ; 
      RECT 8.588 134.946 8.692 139.32 ; 
      RECT 8.156 134.946 8.26 139.32 ; 
      RECT 7.724 134.946 7.828 139.32 ; 
      RECT 7.292 134.946 7.396 139.32 ; 
      RECT 6.86 134.946 6.964 139.32 ; 
      RECT 6.428 134.946 6.532 139.32 ; 
      RECT 5.996 134.946 6.1 139.32 ; 
      RECT 5.564 134.946 5.668 139.32 ; 
      RECT 5.132 134.946 5.236 139.32 ; 
      RECT 4.7 134.946 4.804 139.32 ; 
      RECT 4.268 134.946 4.372 139.32 ; 
      RECT 3.836 134.946 3.94 139.32 ; 
      RECT 3.404 134.946 3.508 139.32 ; 
      RECT 2.972 134.946 3.076 139.32 ; 
      RECT 2.54 134.946 2.644 139.32 ; 
      RECT 2.108 134.946 2.212 139.32 ; 
      RECT 1.676 134.946 1.78 139.32 ; 
      RECT 1.244 134.946 1.348 139.32 ; 
      RECT 0.812 134.946 0.916 139.32 ; 
      RECT 0 134.946 0.34 139.32 ; 
      RECT 20.72 139.266 21.232 143.64 ; 
      RECT 20.664 141.928 21.232 143.218 ; 
      RECT 20.072 140.836 20.32 143.64 ; 
      RECT 20.016 142.074 20.32 142.688 ; 
      RECT 20.072 139.266 20.176 143.64 ; 
      RECT 20.072 139.75 20.232 140.708 ; 
      RECT 20.072 139.266 20.32 139.622 ; 
      RECT 18.884 141.068 19.708 143.64 ; 
      RECT 19.604 139.266 19.708 143.64 ; 
      RECT 18.884 142.176 19.764 143.208 ; 
      RECT 18.884 139.266 19.276 143.64 ; 
      RECT 17.216 139.266 17.548 143.64 ; 
      RECT 17.216 139.62 17.604 143.362 ; 
      RECT 38.108 139.266 38.448 143.64 ; 
      RECT 37.532 139.266 37.636 143.64 ; 
      RECT 37.1 139.266 37.204 143.64 ; 
      RECT 36.668 139.266 36.772 143.64 ; 
      RECT 36.236 139.266 36.34 143.64 ; 
      RECT 35.804 139.266 35.908 143.64 ; 
      RECT 35.372 139.266 35.476 143.64 ; 
      RECT 34.94 139.266 35.044 143.64 ; 
      RECT 34.508 139.266 34.612 143.64 ; 
      RECT 34.076 139.266 34.18 143.64 ; 
      RECT 33.644 139.266 33.748 143.64 ; 
      RECT 33.212 139.266 33.316 143.64 ; 
      RECT 32.78 139.266 32.884 143.64 ; 
      RECT 32.348 139.266 32.452 143.64 ; 
      RECT 31.916 139.266 32.02 143.64 ; 
      RECT 31.484 139.266 31.588 143.64 ; 
      RECT 31.052 139.266 31.156 143.64 ; 
      RECT 30.62 139.266 30.724 143.64 ; 
      RECT 30.188 139.266 30.292 143.64 ; 
      RECT 29.756 139.266 29.86 143.64 ; 
      RECT 29.324 139.266 29.428 143.64 ; 
      RECT 28.892 139.266 28.996 143.64 ; 
      RECT 28.46 139.266 28.564 143.64 ; 
      RECT 28.028 139.266 28.132 143.64 ; 
      RECT 27.596 139.266 27.7 143.64 ; 
      RECT 27.164 139.266 27.268 143.64 ; 
      RECT 26.732 139.266 26.836 143.64 ; 
      RECT 26.3 139.266 26.404 143.64 ; 
      RECT 25.868 139.266 25.972 143.64 ; 
      RECT 25.436 139.266 25.54 143.64 ; 
      RECT 25.004 139.266 25.108 143.64 ; 
      RECT 24.572 139.266 24.676 143.64 ; 
      RECT 24.14 139.266 24.244 143.64 ; 
      RECT 23.708 139.266 23.812 143.64 ; 
      RECT 22.856 139.266 23.164 143.64 ; 
      RECT 15.284 139.266 15.592 143.64 ; 
      RECT 14.636 139.266 14.74 143.64 ; 
      RECT 14.204 139.266 14.308 143.64 ; 
      RECT 13.772 139.266 13.876 143.64 ; 
      RECT 13.34 139.266 13.444 143.64 ; 
      RECT 12.908 139.266 13.012 143.64 ; 
      RECT 12.476 139.266 12.58 143.64 ; 
      RECT 12.044 139.266 12.148 143.64 ; 
      RECT 11.612 139.266 11.716 143.64 ; 
      RECT 11.18 139.266 11.284 143.64 ; 
      RECT 10.748 139.266 10.852 143.64 ; 
      RECT 10.316 139.266 10.42 143.64 ; 
      RECT 9.884 139.266 9.988 143.64 ; 
      RECT 9.452 139.266 9.556 143.64 ; 
      RECT 9.02 139.266 9.124 143.64 ; 
      RECT 8.588 139.266 8.692 143.64 ; 
      RECT 8.156 139.266 8.26 143.64 ; 
      RECT 7.724 139.266 7.828 143.64 ; 
      RECT 7.292 139.266 7.396 143.64 ; 
      RECT 6.86 139.266 6.964 143.64 ; 
      RECT 6.428 139.266 6.532 143.64 ; 
      RECT 5.996 139.266 6.1 143.64 ; 
      RECT 5.564 139.266 5.668 143.64 ; 
      RECT 5.132 139.266 5.236 143.64 ; 
      RECT 4.7 139.266 4.804 143.64 ; 
      RECT 4.268 139.266 4.372 143.64 ; 
      RECT 3.836 139.266 3.94 143.64 ; 
      RECT 3.404 139.266 3.508 143.64 ; 
      RECT 2.972 139.266 3.076 143.64 ; 
      RECT 2.54 139.266 2.644 143.64 ; 
      RECT 2.108 139.266 2.212 143.64 ; 
      RECT 1.676 139.266 1.78 143.64 ; 
      RECT 1.244 139.266 1.348 143.64 ; 
      RECT 0.812 139.266 0.916 143.64 ; 
      RECT 0 139.266 0.34 143.64 ; 
      RECT 20.72 143.586 21.232 147.96 ; 
      RECT 20.664 146.248 21.232 147.538 ; 
      RECT 20.072 145.156 20.32 147.96 ; 
      RECT 20.016 146.394 20.32 147.008 ; 
      RECT 20.072 143.586 20.176 147.96 ; 
      RECT 20.072 144.07 20.232 145.028 ; 
      RECT 20.072 143.586 20.32 143.942 ; 
      RECT 18.884 145.388 19.708 147.96 ; 
      RECT 19.604 143.586 19.708 147.96 ; 
      RECT 18.884 146.496 19.764 147.528 ; 
      RECT 18.884 143.586 19.276 147.96 ; 
      RECT 17.216 143.586 17.548 147.96 ; 
      RECT 17.216 143.94 17.604 147.682 ; 
      RECT 38.108 143.586 38.448 147.96 ; 
      RECT 37.532 143.586 37.636 147.96 ; 
      RECT 37.1 143.586 37.204 147.96 ; 
      RECT 36.668 143.586 36.772 147.96 ; 
      RECT 36.236 143.586 36.34 147.96 ; 
      RECT 35.804 143.586 35.908 147.96 ; 
      RECT 35.372 143.586 35.476 147.96 ; 
      RECT 34.94 143.586 35.044 147.96 ; 
      RECT 34.508 143.586 34.612 147.96 ; 
      RECT 34.076 143.586 34.18 147.96 ; 
      RECT 33.644 143.586 33.748 147.96 ; 
      RECT 33.212 143.586 33.316 147.96 ; 
      RECT 32.78 143.586 32.884 147.96 ; 
      RECT 32.348 143.586 32.452 147.96 ; 
      RECT 31.916 143.586 32.02 147.96 ; 
      RECT 31.484 143.586 31.588 147.96 ; 
      RECT 31.052 143.586 31.156 147.96 ; 
      RECT 30.62 143.586 30.724 147.96 ; 
      RECT 30.188 143.586 30.292 147.96 ; 
      RECT 29.756 143.586 29.86 147.96 ; 
      RECT 29.324 143.586 29.428 147.96 ; 
      RECT 28.892 143.586 28.996 147.96 ; 
      RECT 28.46 143.586 28.564 147.96 ; 
      RECT 28.028 143.586 28.132 147.96 ; 
      RECT 27.596 143.586 27.7 147.96 ; 
      RECT 27.164 143.586 27.268 147.96 ; 
      RECT 26.732 143.586 26.836 147.96 ; 
      RECT 26.3 143.586 26.404 147.96 ; 
      RECT 25.868 143.586 25.972 147.96 ; 
      RECT 25.436 143.586 25.54 147.96 ; 
      RECT 25.004 143.586 25.108 147.96 ; 
      RECT 24.572 143.586 24.676 147.96 ; 
      RECT 24.14 143.586 24.244 147.96 ; 
      RECT 23.708 143.586 23.812 147.96 ; 
      RECT 22.856 143.586 23.164 147.96 ; 
      RECT 15.284 143.586 15.592 147.96 ; 
      RECT 14.636 143.586 14.74 147.96 ; 
      RECT 14.204 143.586 14.308 147.96 ; 
      RECT 13.772 143.586 13.876 147.96 ; 
      RECT 13.34 143.586 13.444 147.96 ; 
      RECT 12.908 143.586 13.012 147.96 ; 
      RECT 12.476 143.586 12.58 147.96 ; 
      RECT 12.044 143.586 12.148 147.96 ; 
      RECT 11.612 143.586 11.716 147.96 ; 
      RECT 11.18 143.586 11.284 147.96 ; 
      RECT 10.748 143.586 10.852 147.96 ; 
      RECT 10.316 143.586 10.42 147.96 ; 
      RECT 9.884 143.586 9.988 147.96 ; 
      RECT 9.452 143.586 9.556 147.96 ; 
      RECT 9.02 143.586 9.124 147.96 ; 
      RECT 8.588 143.586 8.692 147.96 ; 
      RECT 8.156 143.586 8.26 147.96 ; 
      RECT 7.724 143.586 7.828 147.96 ; 
      RECT 7.292 143.586 7.396 147.96 ; 
      RECT 6.86 143.586 6.964 147.96 ; 
      RECT 6.428 143.586 6.532 147.96 ; 
      RECT 5.996 143.586 6.1 147.96 ; 
      RECT 5.564 143.586 5.668 147.96 ; 
      RECT 5.132 143.586 5.236 147.96 ; 
      RECT 4.7 143.586 4.804 147.96 ; 
      RECT 4.268 143.586 4.372 147.96 ; 
      RECT 3.836 143.586 3.94 147.96 ; 
      RECT 3.404 143.586 3.508 147.96 ; 
      RECT 2.972 143.586 3.076 147.96 ; 
      RECT 2.54 143.586 2.644 147.96 ; 
      RECT 2.108 143.586 2.212 147.96 ; 
      RECT 1.676 143.586 1.78 147.96 ; 
      RECT 1.244 143.586 1.348 147.96 ; 
      RECT 0.812 143.586 0.916 147.96 ; 
      RECT 0 143.586 0.34 147.96 ; 
      RECT 20.72 147.906 21.232 152.28 ; 
      RECT 20.664 150.568 21.232 151.858 ; 
      RECT 20.072 149.476 20.32 152.28 ; 
      RECT 20.016 150.714 20.32 151.328 ; 
      RECT 20.072 147.906 20.176 152.28 ; 
      RECT 20.072 148.39 20.232 149.348 ; 
      RECT 20.072 147.906 20.32 148.262 ; 
      RECT 18.884 149.708 19.708 152.28 ; 
      RECT 19.604 147.906 19.708 152.28 ; 
      RECT 18.884 150.816 19.764 151.848 ; 
      RECT 18.884 147.906 19.276 152.28 ; 
      RECT 17.216 147.906 17.548 152.28 ; 
      RECT 17.216 148.26 17.604 152.002 ; 
      RECT 38.108 147.906 38.448 152.28 ; 
      RECT 37.532 147.906 37.636 152.28 ; 
      RECT 37.1 147.906 37.204 152.28 ; 
      RECT 36.668 147.906 36.772 152.28 ; 
      RECT 36.236 147.906 36.34 152.28 ; 
      RECT 35.804 147.906 35.908 152.28 ; 
      RECT 35.372 147.906 35.476 152.28 ; 
      RECT 34.94 147.906 35.044 152.28 ; 
      RECT 34.508 147.906 34.612 152.28 ; 
      RECT 34.076 147.906 34.18 152.28 ; 
      RECT 33.644 147.906 33.748 152.28 ; 
      RECT 33.212 147.906 33.316 152.28 ; 
      RECT 32.78 147.906 32.884 152.28 ; 
      RECT 32.348 147.906 32.452 152.28 ; 
      RECT 31.916 147.906 32.02 152.28 ; 
      RECT 31.484 147.906 31.588 152.28 ; 
      RECT 31.052 147.906 31.156 152.28 ; 
      RECT 30.62 147.906 30.724 152.28 ; 
      RECT 30.188 147.906 30.292 152.28 ; 
      RECT 29.756 147.906 29.86 152.28 ; 
      RECT 29.324 147.906 29.428 152.28 ; 
      RECT 28.892 147.906 28.996 152.28 ; 
      RECT 28.46 147.906 28.564 152.28 ; 
      RECT 28.028 147.906 28.132 152.28 ; 
      RECT 27.596 147.906 27.7 152.28 ; 
      RECT 27.164 147.906 27.268 152.28 ; 
      RECT 26.732 147.906 26.836 152.28 ; 
      RECT 26.3 147.906 26.404 152.28 ; 
      RECT 25.868 147.906 25.972 152.28 ; 
      RECT 25.436 147.906 25.54 152.28 ; 
      RECT 25.004 147.906 25.108 152.28 ; 
      RECT 24.572 147.906 24.676 152.28 ; 
      RECT 24.14 147.906 24.244 152.28 ; 
      RECT 23.708 147.906 23.812 152.28 ; 
      RECT 22.856 147.906 23.164 152.28 ; 
      RECT 15.284 147.906 15.592 152.28 ; 
      RECT 14.636 147.906 14.74 152.28 ; 
      RECT 14.204 147.906 14.308 152.28 ; 
      RECT 13.772 147.906 13.876 152.28 ; 
      RECT 13.34 147.906 13.444 152.28 ; 
      RECT 12.908 147.906 13.012 152.28 ; 
      RECT 12.476 147.906 12.58 152.28 ; 
      RECT 12.044 147.906 12.148 152.28 ; 
      RECT 11.612 147.906 11.716 152.28 ; 
      RECT 11.18 147.906 11.284 152.28 ; 
      RECT 10.748 147.906 10.852 152.28 ; 
      RECT 10.316 147.906 10.42 152.28 ; 
      RECT 9.884 147.906 9.988 152.28 ; 
      RECT 9.452 147.906 9.556 152.28 ; 
      RECT 9.02 147.906 9.124 152.28 ; 
      RECT 8.588 147.906 8.692 152.28 ; 
      RECT 8.156 147.906 8.26 152.28 ; 
      RECT 7.724 147.906 7.828 152.28 ; 
      RECT 7.292 147.906 7.396 152.28 ; 
      RECT 6.86 147.906 6.964 152.28 ; 
      RECT 6.428 147.906 6.532 152.28 ; 
      RECT 5.996 147.906 6.1 152.28 ; 
      RECT 5.564 147.906 5.668 152.28 ; 
      RECT 5.132 147.906 5.236 152.28 ; 
      RECT 4.7 147.906 4.804 152.28 ; 
      RECT 4.268 147.906 4.372 152.28 ; 
      RECT 3.836 147.906 3.94 152.28 ; 
      RECT 3.404 147.906 3.508 152.28 ; 
      RECT 2.972 147.906 3.076 152.28 ; 
      RECT 2.54 147.906 2.644 152.28 ; 
      RECT 2.108 147.906 2.212 152.28 ; 
      RECT 1.676 147.906 1.78 152.28 ; 
      RECT 1.244 147.906 1.348 152.28 ; 
      RECT 0.812 147.906 0.916 152.28 ; 
      RECT 0 147.906 0.34 152.28 ; 
      RECT 20.72 152.226 21.232 156.6 ; 
      RECT 20.664 154.888 21.232 156.178 ; 
      RECT 20.072 153.796 20.32 156.6 ; 
      RECT 20.016 155.034 20.32 155.648 ; 
      RECT 20.072 152.226 20.176 156.6 ; 
      RECT 20.072 152.71 20.232 153.668 ; 
      RECT 20.072 152.226 20.32 152.582 ; 
      RECT 18.884 154.028 19.708 156.6 ; 
      RECT 19.604 152.226 19.708 156.6 ; 
      RECT 18.884 155.136 19.764 156.168 ; 
      RECT 18.884 152.226 19.276 156.6 ; 
      RECT 17.216 152.226 17.548 156.6 ; 
      RECT 17.216 152.58 17.604 156.322 ; 
      RECT 38.108 152.226 38.448 156.6 ; 
      RECT 37.532 152.226 37.636 156.6 ; 
      RECT 37.1 152.226 37.204 156.6 ; 
      RECT 36.668 152.226 36.772 156.6 ; 
      RECT 36.236 152.226 36.34 156.6 ; 
      RECT 35.804 152.226 35.908 156.6 ; 
      RECT 35.372 152.226 35.476 156.6 ; 
      RECT 34.94 152.226 35.044 156.6 ; 
      RECT 34.508 152.226 34.612 156.6 ; 
      RECT 34.076 152.226 34.18 156.6 ; 
      RECT 33.644 152.226 33.748 156.6 ; 
      RECT 33.212 152.226 33.316 156.6 ; 
      RECT 32.78 152.226 32.884 156.6 ; 
      RECT 32.348 152.226 32.452 156.6 ; 
      RECT 31.916 152.226 32.02 156.6 ; 
      RECT 31.484 152.226 31.588 156.6 ; 
      RECT 31.052 152.226 31.156 156.6 ; 
      RECT 30.62 152.226 30.724 156.6 ; 
      RECT 30.188 152.226 30.292 156.6 ; 
      RECT 29.756 152.226 29.86 156.6 ; 
      RECT 29.324 152.226 29.428 156.6 ; 
      RECT 28.892 152.226 28.996 156.6 ; 
      RECT 28.46 152.226 28.564 156.6 ; 
      RECT 28.028 152.226 28.132 156.6 ; 
      RECT 27.596 152.226 27.7 156.6 ; 
      RECT 27.164 152.226 27.268 156.6 ; 
      RECT 26.732 152.226 26.836 156.6 ; 
      RECT 26.3 152.226 26.404 156.6 ; 
      RECT 25.868 152.226 25.972 156.6 ; 
      RECT 25.436 152.226 25.54 156.6 ; 
      RECT 25.004 152.226 25.108 156.6 ; 
      RECT 24.572 152.226 24.676 156.6 ; 
      RECT 24.14 152.226 24.244 156.6 ; 
      RECT 23.708 152.226 23.812 156.6 ; 
      RECT 22.856 152.226 23.164 156.6 ; 
      RECT 15.284 152.226 15.592 156.6 ; 
      RECT 14.636 152.226 14.74 156.6 ; 
      RECT 14.204 152.226 14.308 156.6 ; 
      RECT 13.772 152.226 13.876 156.6 ; 
      RECT 13.34 152.226 13.444 156.6 ; 
      RECT 12.908 152.226 13.012 156.6 ; 
      RECT 12.476 152.226 12.58 156.6 ; 
      RECT 12.044 152.226 12.148 156.6 ; 
      RECT 11.612 152.226 11.716 156.6 ; 
      RECT 11.18 152.226 11.284 156.6 ; 
      RECT 10.748 152.226 10.852 156.6 ; 
      RECT 10.316 152.226 10.42 156.6 ; 
      RECT 9.884 152.226 9.988 156.6 ; 
      RECT 9.452 152.226 9.556 156.6 ; 
      RECT 9.02 152.226 9.124 156.6 ; 
      RECT 8.588 152.226 8.692 156.6 ; 
      RECT 8.156 152.226 8.26 156.6 ; 
      RECT 7.724 152.226 7.828 156.6 ; 
      RECT 7.292 152.226 7.396 156.6 ; 
      RECT 6.86 152.226 6.964 156.6 ; 
      RECT 6.428 152.226 6.532 156.6 ; 
      RECT 5.996 152.226 6.1 156.6 ; 
      RECT 5.564 152.226 5.668 156.6 ; 
      RECT 5.132 152.226 5.236 156.6 ; 
      RECT 4.7 152.226 4.804 156.6 ; 
      RECT 4.268 152.226 4.372 156.6 ; 
      RECT 3.836 152.226 3.94 156.6 ; 
      RECT 3.404 152.226 3.508 156.6 ; 
      RECT 2.972 152.226 3.076 156.6 ; 
      RECT 2.54 152.226 2.644 156.6 ; 
      RECT 2.108 152.226 2.212 156.6 ; 
      RECT 1.676 152.226 1.78 156.6 ; 
      RECT 1.244 152.226 1.348 156.6 ; 
      RECT 0.812 152.226 0.916 156.6 ; 
      RECT 0 152.226 0.34 156.6 ; 
      RECT 20.72 156.546 21.232 160.92 ; 
      RECT 20.664 159.208 21.232 160.498 ; 
      RECT 20.072 158.116 20.32 160.92 ; 
      RECT 20.016 159.354 20.32 159.968 ; 
      RECT 20.072 156.546 20.176 160.92 ; 
      RECT 20.072 157.03 20.232 157.988 ; 
      RECT 20.072 156.546 20.32 156.902 ; 
      RECT 18.884 158.348 19.708 160.92 ; 
      RECT 19.604 156.546 19.708 160.92 ; 
      RECT 18.884 159.456 19.764 160.488 ; 
      RECT 18.884 156.546 19.276 160.92 ; 
      RECT 17.216 156.546 17.548 160.92 ; 
      RECT 17.216 156.9 17.604 160.642 ; 
      RECT 38.108 156.546 38.448 160.92 ; 
      RECT 37.532 156.546 37.636 160.92 ; 
      RECT 37.1 156.546 37.204 160.92 ; 
      RECT 36.668 156.546 36.772 160.92 ; 
      RECT 36.236 156.546 36.34 160.92 ; 
      RECT 35.804 156.546 35.908 160.92 ; 
      RECT 35.372 156.546 35.476 160.92 ; 
      RECT 34.94 156.546 35.044 160.92 ; 
      RECT 34.508 156.546 34.612 160.92 ; 
      RECT 34.076 156.546 34.18 160.92 ; 
      RECT 33.644 156.546 33.748 160.92 ; 
      RECT 33.212 156.546 33.316 160.92 ; 
      RECT 32.78 156.546 32.884 160.92 ; 
      RECT 32.348 156.546 32.452 160.92 ; 
      RECT 31.916 156.546 32.02 160.92 ; 
      RECT 31.484 156.546 31.588 160.92 ; 
      RECT 31.052 156.546 31.156 160.92 ; 
      RECT 30.62 156.546 30.724 160.92 ; 
      RECT 30.188 156.546 30.292 160.92 ; 
      RECT 29.756 156.546 29.86 160.92 ; 
      RECT 29.324 156.546 29.428 160.92 ; 
      RECT 28.892 156.546 28.996 160.92 ; 
      RECT 28.46 156.546 28.564 160.92 ; 
      RECT 28.028 156.546 28.132 160.92 ; 
      RECT 27.596 156.546 27.7 160.92 ; 
      RECT 27.164 156.546 27.268 160.92 ; 
      RECT 26.732 156.546 26.836 160.92 ; 
      RECT 26.3 156.546 26.404 160.92 ; 
      RECT 25.868 156.546 25.972 160.92 ; 
      RECT 25.436 156.546 25.54 160.92 ; 
      RECT 25.004 156.546 25.108 160.92 ; 
      RECT 24.572 156.546 24.676 160.92 ; 
      RECT 24.14 156.546 24.244 160.92 ; 
      RECT 23.708 156.546 23.812 160.92 ; 
      RECT 22.856 156.546 23.164 160.92 ; 
      RECT 15.284 156.546 15.592 160.92 ; 
      RECT 14.636 156.546 14.74 160.92 ; 
      RECT 14.204 156.546 14.308 160.92 ; 
      RECT 13.772 156.546 13.876 160.92 ; 
      RECT 13.34 156.546 13.444 160.92 ; 
      RECT 12.908 156.546 13.012 160.92 ; 
      RECT 12.476 156.546 12.58 160.92 ; 
      RECT 12.044 156.546 12.148 160.92 ; 
      RECT 11.612 156.546 11.716 160.92 ; 
      RECT 11.18 156.546 11.284 160.92 ; 
      RECT 10.748 156.546 10.852 160.92 ; 
      RECT 10.316 156.546 10.42 160.92 ; 
      RECT 9.884 156.546 9.988 160.92 ; 
      RECT 9.452 156.546 9.556 160.92 ; 
      RECT 9.02 156.546 9.124 160.92 ; 
      RECT 8.588 156.546 8.692 160.92 ; 
      RECT 8.156 156.546 8.26 160.92 ; 
      RECT 7.724 156.546 7.828 160.92 ; 
      RECT 7.292 156.546 7.396 160.92 ; 
      RECT 6.86 156.546 6.964 160.92 ; 
      RECT 6.428 156.546 6.532 160.92 ; 
      RECT 5.996 156.546 6.1 160.92 ; 
      RECT 5.564 156.546 5.668 160.92 ; 
      RECT 5.132 156.546 5.236 160.92 ; 
      RECT 4.7 156.546 4.804 160.92 ; 
      RECT 4.268 156.546 4.372 160.92 ; 
      RECT 3.836 156.546 3.94 160.92 ; 
      RECT 3.404 156.546 3.508 160.92 ; 
      RECT 2.972 156.546 3.076 160.92 ; 
      RECT 2.54 156.546 2.644 160.92 ; 
      RECT 2.108 156.546 2.212 160.92 ; 
      RECT 1.676 156.546 1.78 160.92 ; 
      RECT 1.244 156.546 1.348 160.92 ; 
      RECT 0.812 156.546 0.916 160.92 ; 
      RECT 0 156.546 0.34 160.92 ; 
      RECT 20.72 160.866 21.232 165.24 ; 
      RECT 20.664 163.528 21.232 164.818 ; 
      RECT 20.072 162.436 20.32 165.24 ; 
      RECT 20.016 163.674 20.32 164.288 ; 
      RECT 20.072 160.866 20.176 165.24 ; 
      RECT 20.072 161.35 20.232 162.308 ; 
      RECT 20.072 160.866 20.32 161.222 ; 
      RECT 18.884 162.668 19.708 165.24 ; 
      RECT 19.604 160.866 19.708 165.24 ; 
      RECT 18.884 163.776 19.764 164.808 ; 
      RECT 18.884 160.866 19.276 165.24 ; 
      RECT 17.216 160.866 17.548 165.24 ; 
      RECT 17.216 161.22 17.604 164.962 ; 
      RECT 38.108 160.866 38.448 165.24 ; 
      RECT 37.532 160.866 37.636 165.24 ; 
      RECT 37.1 160.866 37.204 165.24 ; 
      RECT 36.668 160.866 36.772 165.24 ; 
      RECT 36.236 160.866 36.34 165.24 ; 
      RECT 35.804 160.866 35.908 165.24 ; 
      RECT 35.372 160.866 35.476 165.24 ; 
      RECT 34.94 160.866 35.044 165.24 ; 
      RECT 34.508 160.866 34.612 165.24 ; 
      RECT 34.076 160.866 34.18 165.24 ; 
      RECT 33.644 160.866 33.748 165.24 ; 
      RECT 33.212 160.866 33.316 165.24 ; 
      RECT 32.78 160.866 32.884 165.24 ; 
      RECT 32.348 160.866 32.452 165.24 ; 
      RECT 31.916 160.866 32.02 165.24 ; 
      RECT 31.484 160.866 31.588 165.24 ; 
      RECT 31.052 160.866 31.156 165.24 ; 
      RECT 30.62 160.866 30.724 165.24 ; 
      RECT 30.188 160.866 30.292 165.24 ; 
      RECT 29.756 160.866 29.86 165.24 ; 
      RECT 29.324 160.866 29.428 165.24 ; 
      RECT 28.892 160.866 28.996 165.24 ; 
      RECT 28.46 160.866 28.564 165.24 ; 
      RECT 28.028 160.866 28.132 165.24 ; 
      RECT 27.596 160.866 27.7 165.24 ; 
      RECT 27.164 160.866 27.268 165.24 ; 
      RECT 26.732 160.866 26.836 165.24 ; 
      RECT 26.3 160.866 26.404 165.24 ; 
      RECT 25.868 160.866 25.972 165.24 ; 
      RECT 25.436 160.866 25.54 165.24 ; 
      RECT 25.004 160.866 25.108 165.24 ; 
      RECT 24.572 160.866 24.676 165.24 ; 
      RECT 24.14 160.866 24.244 165.24 ; 
      RECT 23.708 160.866 23.812 165.24 ; 
      RECT 22.856 160.866 23.164 165.24 ; 
      RECT 15.284 160.866 15.592 165.24 ; 
      RECT 14.636 160.866 14.74 165.24 ; 
      RECT 14.204 160.866 14.308 165.24 ; 
      RECT 13.772 160.866 13.876 165.24 ; 
      RECT 13.34 160.866 13.444 165.24 ; 
      RECT 12.908 160.866 13.012 165.24 ; 
      RECT 12.476 160.866 12.58 165.24 ; 
      RECT 12.044 160.866 12.148 165.24 ; 
      RECT 11.612 160.866 11.716 165.24 ; 
      RECT 11.18 160.866 11.284 165.24 ; 
      RECT 10.748 160.866 10.852 165.24 ; 
      RECT 10.316 160.866 10.42 165.24 ; 
      RECT 9.884 160.866 9.988 165.24 ; 
      RECT 9.452 160.866 9.556 165.24 ; 
      RECT 9.02 160.866 9.124 165.24 ; 
      RECT 8.588 160.866 8.692 165.24 ; 
      RECT 8.156 160.866 8.26 165.24 ; 
      RECT 7.724 160.866 7.828 165.24 ; 
      RECT 7.292 160.866 7.396 165.24 ; 
      RECT 6.86 160.866 6.964 165.24 ; 
      RECT 6.428 160.866 6.532 165.24 ; 
      RECT 5.996 160.866 6.1 165.24 ; 
      RECT 5.564 160.866 5.668 165.24 ; 
      RECT 5.132 160.866 5.236 165.24 ; 
      RECT 4.7 160.866 4.804 165.24 ; 
      RECT 4.268 160.866 4.372 165.24 ; 
      RECT 3.836 160.866 3.94 165.24 ; 
      RECT 3.404 160.866 3.508 165.24 ; 
      RECT 2.972 160.866 3.076 165.24 ; 
      RECT 2.54 160.866 2.644 165.24 ; 
      RECT 2.108 160.866 2.212 165.24 ; 
      RECT 1.676 160.866 1.78 165.24 ; 
      RECT 1.244 160.866 1.348 165.24 ; 
      RECT 0.812 160.866 0.916 165.24 ; 
      RECT 0 160.866 0.34 165.24 ; 
      RECT 20.72 165.186 21.232 169.56 ; 
      RECT 20.664 167.848 21.232 169.138 ; 
      RECT 20.072 166.756 20.32 169.56 ; 
      RECT 20.016 167.994 20.32 168.608 ; 
      RECT 20.072 165.186 20.176 169.56 ; 
      RECT 20.072 165.67 20.232 166.628 ; 
      RECT 20.072 165.186 20.32 165.542 ; 
      RECT 18.884 166.988 19.708 169.56 ; 
      RECT 19.604 165.186 19.708 169.56 ; 
      RECT 18.884 168.096 19.764 169.128 ; 
      RECT 18.884 165.186 19.276 169.56 ; 
      RECT 17.216 165.186 17.548 169.56 ; 
      RECT 17.216 165.54 17.604 169.282 ; 
      RECT 38.108 165.186 38.448 169.56 ; 
      RECT 37.532 165.186 37.636 169.56 ; 
      RECT 37.1 165.186 37.204 169.56 ; 
      RECT 36.668 165.186 36.772 169.56 ; 
      RECT 36.236 165.186 36.34 169.56 ; 
      RECT 35.804 165.186 35.908 169.56 ; 
      RECT 35.372 165.186 35.476 169.56 ; 
      RECT 34.94 165.186 35.044 169.56 ; 
      RECT 34.508 165.186 34.612 169.56 ; 
      RECT 34.076 165.186 34.18 169.56 ; 
      RECT 33.644 165.186 33.748 169.56 ; 
      RECT 33.212 165.186 33.316 169.56 ; 
      RECT 32.78 165.186 32.884 169.56 ; 
      RECT 32.348 165.186 32.452 169.56 ; 
      RECT 31.916 165.186 32.02 169.56 ; 
      RECT 31.484 165.186 31.588 169.56 ; 
      RECT 31.052 165.186 31.156 169.56 ; 
      RECT 30.62 165.186 30.724 169.56 ; 
      RECT 30.188 165.186 30.292 169.56 ; 
      RECT 29.756 165.186 29.86 169.56 ; 
      RECT 29.324 165.186 29.428 169.56 ; 
      RECT 28.892 165.186 28.996 169.56 ; 
      RECT 28.46 165.186 28.564 169.56 ; 
      RECT 28.028 165.186 28.132 169.56 ; 
      RECT 27.596 165.186 27.7 169.56 ; 
      RECT 27.164 165.186 27.268 169.56 ; 
      RECT 26.732 165.186 26.836 169.56 ; 
      RECT 26.3 165.186 26.404 169.56 ; 
      RECT 25.868 165.186 25.972 169.56 ; 
      RECT 25.436 165.186 25.54 169.56 ; 
      RECT 25.004 165.186 25.108 169.56 ; 
      RECT 24.572 165.186 24.676 169.56 ; 
      RECT 24.14 165.186 24.244 169.56 ; 
      RECT 23.708 165.186 23.812 169.56 ; 
      RECT 22.856 165.186 23.164 169.56 ; 
      RECT 15.284 165.186 15.592 169.56 ; 
      RECT 14.636 165.186 14.74 169.56 ; 
      RECT 14.204 165.186 14.308 169.56 ; 
      RECT 13.772 165.186 13.876 169.56 ; 
      RECT 13.34 165.186 13.444 169.56 ; 
      RECT 12.908 165.186 13.012 169.56 ; 
      RECT 12.476 165.186 12.58 169.56 ; 
      RECT 12.044 165.186 12.148 169.56 ; 
      RECT 11.612 165.186 11.716 169.56 ; 
      RECT 11.18 165.186 11.284 169.56 ; 
      RECT 10.748 165.186 10.852 169.56 ; 
      RECT 10.316 165.186 10.42 169.56 ; 
      RECT 9.884 165.186 9.988 169.56 ; 
      RECT 9.452 165.186 9.556 169.56 ; 
      RECT 9.02 165.186 9.124 169.56 ; 
      RECT 8.588 165.186 8.692 169.56 ; 
      RECT 8.156 165.186 8.26 169.56 ; 
      RECT 7.724 165.186 7.828 169.56 ; 
      RECT 7.292 165.186 7.396 169.56 ; 
      RECT 6.86 165.186 6.964 169.56 ; 
      RECT 6.428 165.186 6.532 169.56 ; 
      RECT 5.996 165.186 6.1 169.56 ; 
      RECT 5.564 165.186 5.668 169.56 ; 
      RECT 5.132 165.186 5.236 169.56 ; 
      RECT 4.7 165.186 4.804 169.56 ; 
      RECT 4.268 165.186 4.372 169.56 ; 
      RECT 3.836 165.186 3.94 169.56 ; 
      RECT 3.404 165.186 3.508 169.56 ; 
      RECT 2.972 165.186 3.076 169.56 ; 
      RECT 2.54 165.186 2.644 169.56 ; 
      RECT 2.108 165.186 2.212 169.56 ; 
      RECT 1.676 165.186 1.78 169.56 ; 
      RECT 1.244 165.186 1.348 169.56 ; 
      RECT 0.812 165.186 0.916 169.56 ; 
      RECT 0 165.186 0.34 169.56 ; 
      RECT 20.72 169.506 21.232 173.88 ; 
      RECT 20.664 172.168 21.232 173.458 ; 
      RECT 20.072 171.076 20.32 173.88 ; 
      RECT 20.016 172.314 20.32 172.928 ; 
      RECT 20.072 169.506 20.176 173.88 ; 
      RECT 20.072 169.99 20.232 170.948 ; 
      RECT 20.072 169.506 20.32 169.862 ; 
      RECT 18.884 171.308 19.708 173.88 ; 
      RECT 19.604 169.506 19.708 173.88 ; 
      RECT 18.884 172.416 19.764 173.448 ; 
      RECT 18.884 169.506 19.276 173.88 ; 
      RECT 17.216 169.506 17.548 173.88 ; 
      RECT 17.216 169.86 17.604 173.602 ; 
      RECT 38.108 169.506 38.448 173.88 ; 
      RECT 37.532 169.506 37.636 173.88 ; 
      RECT 37.1 169.506 37.204 173.88 ; 
      RECT 36.668 169.506 36.772 173.88 ; 
      RECT 36.236 169.506 36.34 173.88 ; 
      RECT 35.804 169.506 35.908 173.88 ; 
      RECT 35.372 169.506 35.476 173.88 ; 
      RECT 34.94 169.506 35.044 173.88 ; 
      RECT 34.508 169.506 34.612 173.88 ; 
      RECT 34.076 169.506 34.18 173.88 ; 
      RECT 33.644 169.506 33.748 173.88 ; 
      RECT 33.212 169.506 33.316 173.88 ; 
      RECT 32.78 169.506 32.884 173.88 ; 
      RECT 32.348 169.506 32.452 173.88 ; 
      RECT 31.916 169.506 32.02 173.88 ; 
      RECT 31.484 169.506 31.588 173.88 ; 
      RECT 31.052 169.506 31.156 173.88 ; 
      RECT 30.62 169.506 30.724 173.88 ; 
      RECT 30.188 169.506 30.292 173.88 ; 
      RECT 29.756 169.506 29.86 173.88 ; 
      RECT 29.324 169.506 29.428 173.88 ; 
      RECT 28.892 169.506 28.996 173.88 ; 
      RECT 28.46 169.506 28.564 173.88 ; 
      RECT 28.028 169.506 28.132 173.88 ; 
      RECT 27.596 169.506 27.7 173.88 ; 
      RECT 27.164 169.506 27.268 173.88 ; 
      RECT 26.732 169.506 26.836 173.88 ; 
      RECT 26.3 169.506 26.404 173.88 ; 
      RECT 25.868 169.506 25.972 173.88 ; 
      RECT 25.436 169.506 25.54 173.88 ; 
      RECT 25.004 169.506 25.108 173.88 ; 
      RECT 24.572 169.506 24.676 173.88 ; 
      RECT 24.14 169.506 24.244 173.88 ; 
      RECT 23.708 169.506 23.812 173.88 ; 
      RECT 22.856 169.506 23.164 173.88 ; 
      RECT 15.284 169.506 15.592 173.88 ; 
      RECT 14.636 169.506 14.74 173.88 ; 
      RECT 14.204 169.506 14.308 173.88 ; 
      RECT 13.772 169.506 13.876 173.88 ; 
      RECT 13.34 169.506 13.444 173.88 ; 
      RECT 12.908 169.506 13.012 173.88 ; 
      RECT 12.476 169.506 12.58 173.88 ; 
      RECT 12.044 169.506 12.148 173.88 ; 
      RECT 11.612 169.506 11.716 173.88 ; 
      RECT 11.18 169.506 11.284 173.88 ; 
      RECT 10.748 169.506 10.852 173.88 ; 
      RECT 10.316 169.506 10.42 173.88 ; 
      RECT 9.884 169.506 9.988 173.88 ; 
      RECT 9.452 169.506 9.556 173.88 ; 
      RECT 9.02 169.506 9.124 173.88 ; 
      RECT 8.588 169.506 8.692 173.88 ; 
      RECT 8.156 169.506 8.26 173.88 ; 
      RECT 7.724 169.506 7.828 173.88 ; 
      RECT 7.292 169.506 7.396 173.88 ; 
      RECT 6.86 169.506 6.964 173.88 ; 
      RECT 6.428 169.506 6.532 173.88 ; 
      RECT 5.996 169.506 6.1 173.88 ; 
      RECT 5.564 169.506 5.668 173.88 ; 
      RECT 5.132 169.506 5.236 173.88 ; 
      RECT 4.7 169.506 4.804 173.88 ; 
      RECT 4.268 169.506 4.372 173.88 ; 
      RECT 3.836 169.506 3.94 173.88 ; 
      RECT 3.404 169.506 3.508 173.88 ; 
      RECT 2.972 169.506 3.076 173.88 ; 
      RECT 2.54 169.506 2.644 173.88 ; 
      RECT 2.108 169.506 2.212 173.88 ; 
      RECT 1.676 169.506 1.78 173.88 ; 
      RECT 1.244 169.506 1.348 173.88 ; 
      RECT 0.812 169.506 0.916 173.88 ; 
      RECT 0 169.506 0.34 173.88 ; 
      RECT 0 207.216 38.448 208.386 ; 
      RECT 38.108 173.772 38.448 208.386 ; 
      RECT 18.164 206.622 38.448 208.386 ; 
      RECT 0 206.622 17.548 208.386 ; 
      RECT 23.708 179.788 37.636 208.386 ; 
      RECT 29.54 173.772 37.636 208.386 ; 
      RECT 18.164 206.516 23.38 208.386 ; 
      RECT 20.72 206.512 23.38 208.386 ; 
      RECT 15.068 180.22 17.548 208.386 ; 
      RECT 15.284 176.836 17.548 208.386 ; 
      RECT 0.812 179.008 14.74 208.386 ; 
      RECT 13.556 173.772 14.74 208.386 ; 
      RECT 0 173.772 0.34 208.386 ; 
      RECT 18.164 206.504 20.32 208.386 ; 
      RECT 20.072 205.42 20.32 208.386 ; 
      RECT 20.72 205.42 23.164 208.386 ; 
      RECT 18.164 205.42 19.708 208.386 ; 
      RECT 23.652 188.944 37.636 206.384 ; 
      RECT 0.812 188.944 14.796 206.384 ; 
      RECT 23.652 188.944 37.692 206.366 ; 
      RECT 0.756 188.944 14.796 206.366 ; 
      RECT 20.756 176.836 23.164 208.386 ; 
      RECT 18.884 176.512 19.564 208.386 ; 
      RECT 19.316 173.772 19.564 208.386 ; 
      RECT 16.148 176.108 17.692 204.82 ; 
      RECT 15.068 204.652 17.748 204.8 ; 
      RECT 20.7 200.356 23.164 204.788 ; 
      RECT 18.828 203.596 19.564 204.5 ; 
      RECT 18.884 201.292 19.62 202.34 ; 
      RECT 15.068 200.5 17.748 202.34 ; 
      RECT 18.828 198.34 19.564 200.18 ; 
      RECT 20.7 190.204 23.164 199.532 ; 
      RECT 15.068 192.796 17.748 197.372 ; 
      RECT 18.884 191.716 19.62 196.94 ; 
      RECT 18.828 194.02 19.62 195.86 ; 
      RECT 18.828 181.06 19.564 193.7 ; 
      RECT 18.828 181.06 19.62 191.54 ; 
      RECT 15.068 190.636 17.748 191.54 ; 
      RECT 20.9 174.478 23.38 188.816 ; 
      RECT 20.7 178.9 23.38 186.044 ; 
      RECT 15.068 182.788 17.748 184.268 ; 
      RECT 18.884 179.98 19.62 180.74 ; 
      RECT 15.284 179.836 17.748 180.596 ; 
      RECT 18.828 179.404 19.564 179.948 ; 
      RECT 18.884 178.9 19.62 179.804 ; 
      RECT 24.356 179.02 37.636 208.386 ; 
      RECT 28.676 179.008 37.636 208.386 ; 
      RECT 23.708 173.772 24.028 208.386 ; 
      RECT 15.068 176.512 15.82 179.768 ; 
      RECT 23.708 173.772 24.892 179.384 ; 
      RECT 23.708 178.24 28.348 179.384 ; 
      RECT 28.676 173.772 29.212 208.386 ; 
      RECT 10.1 177.484 13.228 208.386 ; 
      RECT 0.812 173.772 9.772 208.386 ; 
      RECT 23.708 178.24 29.212 178.616 ; 
      RECT 27.812 173.772 37.636 178.604 ; 
      RECT 12.692 173.772 14.74 178.604 ; 
      RECT 18.828 178.324 19.62 178.58 ; 
      RECT 18.828 177.82 19.564 178.58 ; 
      RECT 26.948 176.704 37.636 178.604 ; 
      RECT 23.708 176.836 26.62 179.384 ; 
      RECT 18.884 176.74 19.62 177.788 ; 
      RECT 0.812 176.704 12.364 178.604 ; 
      RECT 11.828 173.772 12.364 208.386 ; 
      RECT 26.084 173.772 27.484 177.26 ; 
      RECT 23.708 176.512 25.756 179.384 ; 
      RECT 25.22 173.772 25.756 208.386 ; 
      RECT 10.964 176.512 12.364 208.386 ; 
      RECT 0.812 173.772 10.636 178.604 ; 
      RECT 18.884 173.772 18.988 208.386 ; 
      RECT 15.428 173.772 15.82 208.386 ; 
      RECT 10.964 173.772 11.5 208.386 ; 
      RECT 25.22 173.772 27.484 176.312 ; 
      RECT 20.756 173.772 23.164 176.312 ; 
      RECT 15.428 173.772 17.548 176.312 ; 
      RECT 11.828 173.772 14.74 176.312 ; 
      RECT 25.22 173.772 37.636 176.3 ; 
      RECT 0.812 173.772 11.5 176.3 ; 
      RECT 20.7 175.66 23.38 176.276 ; 
      RECT 15.428 175.66 17.604 176.312 ; 
      RECT 23.708 173.772 37.636 175.244 ; 
      RECT 18.884 173.772 19.564 175.244 ; 
      RECT 15.068 173.772 17.548 175.244 ; 
      RECT 0.812 173.772 14.74 175.244 ; 
      RECT 18.164 173.772 19.564 174.832 ; 
      RECT 20.72 173.772 23.164 174.432 ; 
      RECT 18.164 173.772 19.708 174.432 ; 
      RECT 20.72 173.772 23.38 173.856 ; 
      RECT 25.236 173.666 25.308 208.386 ; 
      RECT 24.804 173.666 24.876 208.386 ; 
      RECT 11.844 173.666 11.916 208.386 ; 
      RECT 11.412 173.666 11.484 208.386 ; 
      RECT 20.072 173.772 20.32 174.432 ; 
        RECT 20.72 206.334 21.232 210.708 ; 
        RECT 20.664 208.996 21.232 210.286 ; 
        RECT 20.072 207.904 20.32 210.708 ; 
        RECT 20.016 209.142 20.32 209.756 ; 
        RECT 20.072 206.334 20.176 210.708 ; 
        RECT 20.072 206.818 20.232 207.776 ; 
        RECT 20.072 206.334 20.32 206.69 ; 
        RECT 18.884 208.136 19.708 210.708 ; 
        RECT 19.604 206.334 19.708 210.708 ; 
        RECT 18.884 209.244 19.764 210.276 ; 
        RECT 18.884 206.334 19.276 210.708 ; 
        RECT 17.216 206.334 17.548 210.708 ; 
        RECT 17.216 206.688 17.604 210.43 ; 
        RECT 38.108 206.334 38.448 210.708 ; 
        RECT 37.532 206.334 37.636 210.708 ; 
        RECT 37.1 206.334 37.204 210.708 ; 
        RECT 36.668 206.334 36.772 210.708 ; 
        RECT 36.236 206.334 36.34 210.708 ; 
        RECT 35.804 206.334 35.908 210.708 ; 
        RECT 35.372 206.334 35.476 210.708 ; 
        RECT 34.94 206.334 35.044 210.708 ; 
        RECT 34.508 206.334 34.612 210.708 ; 
        RECT 34.076 206.334 34.18 210.708 ; 
        RECT 33.644 206.334 33.748 210.708 ; 
        RECT 33.212 206.334 33.316 210.708 ; 
        RECT 32.78 206.334 32.884 210.708 ; 
        RECT 32.348 206.334 32.452 210.708 ; 
        RECT 31.916 206.334 32.02 210.708 ; 
        RECT 31.484 206.334 31.588 210.708 ; 
        RECT 31.052 206.334 31.156 210.708 ; 
        RECT 30.62 206.334 30.724 210.708 ; 
        RECT 30.188 206.334 30.292 210.708 ; 
        RECT 29.756 206.334 29.86 210.708 ; 
        RECT 29.324 206.334 29.428 210.708 ; 
        RECT 28.892 206.334 28.996 210.708 ; 
        RECT 28.46 206.334 28.564 210.708 ; 
        RECT 28.028 206.334 28.132 210.708 ; 
        RECT 27.596 206.334 27.7 210.708 ; 
        RECT 27.164 206.334 27.268 210.708 ; 
        RECT 26.732 206.334 26.836 210.708 ; 
        RECT 26.3 206.334 26.404 210.708 ; 
        RECT 25.868 206.334 25.972 210.708 ; 
        RECT 25.436 206.334 25.54 210.708 ; 
        RECT 25.004 206.334 25.108 210.708 ; 
        RECT 24.572 206.334 24.676 210.708 ; 
        RECT 24.14 206.334 24.244 210.708 ; 
        RECT 23.708 206.334 23.812 210.708 ; 
        RECT 22.856 206.334 23.164 210.708 ; 
        RECT 15.284 206.334 15.592 210.708 ; 
        RECT 14.636 206.334 14.74 210.708 ; 
        RECT 14.204 206.334 14.308 210.708 ; 
        RECT 13.772 206.334 13.876 210.708 ; 
        RECT 13.34 206.334 13.444 210.708 ; 
        RECT 12.908 206.334 13.012 210.708 ; 
        RECT 12.476 206.334 12.58 210.708 ; 
        RECT 12.044 206.334 12.148 210.708 ; 
        RECT 11.612 206.334 11.716 210.708 ; 
        RECT 11.18 206.334 11.284 210.708 ; 
        RECT 10.748 206.334 10.852 210.708 ; 
        RECT 10.316 206.334 10.42 210.708 ; 
        RECT 9.884 206.334 9.988 210.708 ; 
        RECT 9.452 206.334 9.556 210.708 ; 
        RECT 9.02 206.334 9.124 210.708 ; 
        RECT 8.588 206.334 8.692 210.708 ; 
        RECT 8.156 206.334 8.26 210.708 ; 
        RECT 7.724 206.334 7.828 210.708 ; 
        RECT 7.292 206.334 7.396 210.708 ; 
        RECT 6.86 206.334 6.964 210.708 ; 
        RECT 6.428 206.334 6.532 210.708 ; 
        RECT 5.996 206.334 6.1 210.708 ; 
        RECT 5.564 206.334 5.668 210.708 ; 
        RECT 5.132 206.334 5.236 210.708 ; 
        RECT 4.7 206.334 4.804 210.708 ; 
        RECT 4.268 206.334 4.372 210.708 ; 
        RECT 3.836 206.334 3.94 210.708 ; 
        RECT 3.404 206.334 3.508 210.708 ; 
        RECT 2.972 206.334 3.076 210.708 ; 
        RECT 2.54 206.334 2.644 210.708 ; 
        RECT 2.108 206.334 2.212 210.708 ; 
        RECT 1.676 206.334 1.78 210.708 ; 
        RECT 1.244 206.334 1.348 210.708 ; 
        RECT 0.812 206.334 0.916 210.708 ; 
        RECT 0 206.334 0.34 210.708 ; 
        RECT 20.72 210.654 21.232 215.028 ; 
        RECT 20.664 213.316 21.232 214.606 ; 
        RECT 20.072 212.224 20.32 215.028 ; 
        RECT 20.016 213.462 20.32 214.076 ; 
        RECT 20.072 210.654 20.176 215.028 ; 
        RECT 20.072 211.138 20.232 212.096 ; 
        RECT 20.072 210.654 20.32 211.01 ; 
        RECT 18.884 212.456 19.708 215.028 ; 
        RECT 19.604 210.654 19.708 215.028 ; 
        RECT 18.884 213.564 19.764 214.596 ; 
        RECT 18.884 210.654 19.276 215.028 ; 
        RECT 17.216 210.654 17.548 215.028 ; 
        RECT 17.216 211.008 17.604 214.75 ; 
        RECT 38.108 210.654 38.448 215.028 ; 
        RECT 37.532 210.654 37.636 215.028 ; 
        RECT 37.1 210.654 37.204 215.028 ; 
        RECT 36.668 210.654 36.772 215.028 ; 
        RECT 36.236 210.654 36.34 215.028 ; 
        RECT 35.804 210.654 35.908 215.028 ; 
        RECT 35.372 210.654 35.476 215.028 ; 
        RECT 34.94 210.654 35.044 215.028 ; 
        RECT 34.508 210.654 34.612 215.028 ; 
        RECT 34.076 210.654 34.18 215.028 ; 
        RECT 33.644 210.654 33.748 215.028 ; 
        RECT 33.212 210.654 33.316 215.028 ; 
        RECT 32.78 210.654 32.884 215.028 ; 
        RECT 32.348 210.654 32.452 215.028 ; 
        RECT 31.916 210.654 32.02 215.028 ; 
        RECT 31.484 210.654 31.588 215.028 ; 
        RECT 31.052 210.654 31.156 215.028 ; 
        RECT 30.62 210.654 30.724 215.028 ; 
        RECT 30.188 210.654 30.292 215.028 ; 
        RECT 29.756 210.654 29.86 215.028 ; 
        RECT 29.324 210.654 29.428 215.028 ; 
        RECT 28.892 210.654 28.996 215.028 ; 
        RECT 28.46 210.654 28.564 215.028 ; 
        RECT 28.028 210.654 28.132 215.028 ; 
        RECT 27.596 210.654 27.7 215.028 ; 
        RECT 27.164 210.654 27.268 215.028 ; 
        RECT 26.732 210.654 26.836 215.028 ; 
        RECT 26.3 210.654 26.404 215.028 ; 
        RECT 25.868 210.654 25.972 215.028 ; 
        RECT 25.436 210.654 25.54 215.028 ; 
        RECT 25.004 210.654 25.108 215.028 ; 
        RECT 24.572 210.654 24.676 215.028 ; 
        RECT 24.14 210.654 24.244 215.028 ; 
        RECT 23.708 210.654 23.812 215.028 ; 
        RECT 22.856 210.654 23.164 215.028 ; 
        RECT 15.284 210.654 15.592 215.028 ; 
        RECT 14.636 210.654 14.74 215.028 ; 
        RECT 14.204 210.654 14.308 215.028 ; 
        RECT 13.772 210.654 13.876 215.028 ; 
        RECT 13.34 210.654 13.444 215.028 ; 
        RECT 12.908 210.654 13.012 215.028 ; 
        RECT 12.476 210.654 12.58 215.028 ; 
        RECT 12.044 210.654 12.148 215.028 ; 
        RECT 11.612 210.654 11.716 215.028 ; 
        RECT 11.18 210.654 11.284 215.028 ; 
        RECT 10.748 210.654 10.852 215.028 ; 
        RECT 10.316 210.654 10.42 215.028 ; 
        RECT 9.884 210.654 9.988 215.028 ; 
        RECT 9.452 210.654 9.556 215.028 ; 
        RECT 9.02 210.654 9.124 215.028 ; 
        RECT 8.588 210.654 8.692 215.028 ; 
        RECT 8.156 210.654 8.26 215.028 ; 
        RECT 7.724 210.654 7.828 215.028 ; 
        RECT 7.292 210.654 7.396 215.028 ; 
        RECT 6.86 210.654 6.964 215.028 ; 
        RECT 6.428 210.654 6.532 215.028 ; 
        RECT 5.996 210.654 6.1 215.028 ; 
        RECT 5.564 210.654 5.668 215.028 ; 
        RECT 5.132 210.654 5.236 215.028 ; 
        RECT 4.7 210.654 4.804 215.028 ; 
        RECT 4.268 210.654 4.372 215.028 ; 
        RECT 3.836 210.654 3.94 215.028 ; 
        RECT 3.404 210.654 3.508 215.028 ; 
        RECT 2.972 210.654 3.076 215.028 ; 
        RECT 2.54 210.654 2.644 215.028 ; 
        RECT 2.108 210.654 2.212 215.028 ; 
        RECT 1.676 210.654 1.78 215.028 ; 
        RECT 1.244 210.654 1.348 215.028 ; 
        RECT 0.812 210.654 0.916 215.028 ; 
        RECT 0 210.654 0.34 215.028 ; 
        RECT 20.72 214.974 21.232 219.348 ; 
        RECT 20.664 217.636 21.232 218.926 ; 
        RECT 20.072 216.544 20.32 219.348 ; 
        RECT 20.016 217.782 20.32 218.396 ; 
        RECT 20.072 214.974 20.176 219.348 ; 
        RECT 20.072 215.458 20.232 216.416 ; 
        RECT 20.072 214.974 20.32 215.33 ; 
        RECT 18.884 216.776 19.708 219.348 ; 
        RECT 19.604 214.974 19.708 219.348 ; 
        RECT 18.884 217.884 19.764 218.916 ; 
        RECT 18.884 214.974 19.276 219.348 ; 
        RECT 17.216 214.974 17.548 219.348 ; 
        RECT 17.216 215.328 17.604 219.07 ; 
        RECT 38.108 214.974 38.448 219.348 ; 
        RECT 37.532 214.974 37.636 219.348 ; 
        RECT 37.1 214.974 37.204 219.348 ; 
        RECT 36.668 214.974 36.772 219.348 ; 
        RECT 36.236 214.974 36.34 219.348 ; 
        RECT 35.804 214.974 35.908 219.348 ; 
        RECT 35.372 214.974 35.476 219.348 ; 
        RECT 34.94 214.974 35.044 219.348 ; 
        RECT 34.508 214.974 34.612 219.348 ; 
        RECT 34.076 214.974 34.18 219.348 ; 
        RECT 33.644 214.974 33.748 219.348 ; 
        RECT 33.212 214.974 33.316 219.348 ; 
        RECT 32.78 214.974 32.884 219.348 ; 
        RECT 32.348 214.974 32.452 219.348 ; 
        RECT 31.916 214.974 32.02 219.348 ; 
        RECT 31.484 214.974 31.588 219.348 ; 
        RECT 31.052 214.974 31.156 219.348 ; 
        RECT 30.62 214.974 30.724 219.348 ; 
        RECT 30.188 214.974 30.292 219.348 ; 
        RECT 29.756 214.974 29.86 219.348 ; 
        RECT 29.324 214.974 29.428 219.348 ; 
        RECT 28.892 214.974 28.996 219.348 ; 
        RECT 28.46 214.974 28.564 219.348 ; 
        RECT 28.028 214.974 28.132 219.348 ; 
        RECT 27.596 214.974 27.7 219.348 ; 
        RECT 27.164 214.974 27.268 219.348 ; 
        RECT 26.732 214.974 26.836 219.348 ; 
        RECT 26.3 214.974 26.404 219.348 ; 
        RECT 25.868 214.974 25.972 219.348 ; 
        RECT 25.436 214.974 25.54 219.348 ; 
        RECT 25.004 214.974 25.108 219.348 ; 
        RECT 24.572 214.974 24.676 219.348 ; 
        RECT 24.14 214.974 24.244 219.348 ; 
        RECT 23.708 214.974 23.812 219.348 ; 
        RECT 22.856 214.974 23.164 219.348 ; 
        RECT 15.284 214.974 15.592 219.348 ; 
        RECT 14.636 214.974 14.74 219.348 ; 
        RECT 14.204 214.974 14.308 219.348 ; 
        RECT 13.772 214.974 13.876 219.348 ; 
        RECT 13.34 214.974 13.444 219.348 ; 
        RECT 12.908 214.974 13.012 219.348 ; 
        RECT 12.476 214.974 12.58 219.348 ; 
        RECT 12.044 214.974 12.148 219.348 ; 
        RECT 11.612 214.974 11.716 219.348 ; 
        RECT 11.18 214.974 11.284 219.348 ; 
        RECT 10.748 214.974 10.852 219.348 ; 
        RECT 10.316 214.974 10.42 219.348 ; 
        RECT 9.884 214.974 9.988 219.348 ; 
        RECT 9.452 214.974 9.556 219.348 ; 
        RECT 9.02 214.974 9.124 219.348 ; 
        RECT 8.588 214.974 8.692 219.348 ; 
        RECT 8.156 214.974 8.26 219.348 ; 
        RECT 7.724 214.974 7.828 219.348 ; 
        RECT 7.292 214.974 7.396 219.348 ; 
        RECT 6.86 214.974 6.964 219.348 ; 
        RECT 6.428 214.974 6.532 219.348 ; 
        RECT 5.996 214.974 6.1 219.348 ; 
        RECT 5.564 214.974 5.668 219.348 ; 
        RECT 5.132 214.974 5.236 219.348 ; 
        RECT 4.7 214.974 4.804 219.348 ; 
        RECT 4.268 214.974 4.372 219.348 ; 
        RECT 3.836 214.974 3.94 219.348 ; 
        RECT 3.404 214.974 3.508 219.348 ; 
        RECT 2.972 214.974 3.076 219.348 ; 
        RECT 2.54 214.974 2.644 219.348 ; 
        RECT 2.108 214.974 2.212 219.348 ; 
        RECT 1.676 214.974 1.78 219.348 ; 
        RECT 1.244 214.974 1.348 219.348 ; 
        RECT 0.812 214.974 0.916 219.348 ; 
        RECT 0 214.974 0.34 219.348 ; 
        RECT 20.72 219.294 21.232 223.668 ; 
        RECT 20.664 221.956 21.232 223.246 ; 
        RECT 20.072 220.864 20.32 223.668 ; 
        RECT 20.016 222.102 20.32 222.716 ; 
        RECT 20.072 219.294 20.176 223.668 ; 
        RECT 20.072 219.778 20.232 220.736 ; 
        RECT 20.072 219.294 20.32 219.65 ; 
        RECT 18.884 221.096 19.708 223.668 ; 
        RECT 19.604 219.294 19.708 223.668 ; 
        RECT 18.884 222.204 19.764 223.236 ; 
        RECT 18.884 219.294 19.276 223.668 ; 
        RECT 17.216 219.294 17.548 223.668 ; 
        RECT 17.216 219.648 17.604 223.39 ; 
        RECT 38.108 219.294 38.448 223.668 ; 
        RECT 37.532 219.294 37.636 223.668 ; 
        RECT 37.1 219.294 37.204 223.668 ; 
        RECT 36.668 219.294 36.772 223.668 ; 
        RECT 36.236 219.294 36.34 223.668 ; 
        RECT 35.804 219.294 35.908 223.668 ; 
        RECT 35.372 219.294 35.476 223.668 ; 
        RECT 34.94 219.294 35.044 223.668 ; 
        RECT 34.508 219.294 34.612 223.668 ; 
        RECT 34.076 219.294 34.18 223.668 ; 
        RECT 33.644 219.294 33.748 223.668 ; 
        RECT 33.212 219.294 33.316 223.668 ; 
        RECT 32.78 219.294 32.884 223.668 ; 
        RECT 32.348 219.294 32.452 223.668 ; 
        RECT 31.916 219.294 32.02 223.668 ; 
        RECT 31.484 219.294 31.588 223.668 ; 
        RECT 31.052 219.294 31.156 223.668 ; 
        RECT 30.62 219.294 30.724 223.668 ; 
        RECT 30.188 219.294 30.292 223.668 ; 
        RECT 29.756 219.294 29.86 223.668 ; 
        RECT 29.324 219.294 29.428 223.668 ; 
        RECT 28.892 219.294 28.996 223.668 ; 
        RECT 28.46 219.294 28.564 223.668 ; 
        RECT 28.028 219.294 28.132 223.668 ; 
        RECT 27.596 219.294 27.7 223.668 ; 
        RECT 27.164 219.294 27.268 223.668 ; 
        RECT 26.732 219.294 26.836 223.668 ; 
        RECT 26.3 219.294 26.404 223.668 ; 
        RECT 25.868 219.294 25.972 223.668 ; 
        RECT 25.436 219.294 25.54 223.668 ; 
        RECT 25.004 219.294 25.108 223.668 ; 
        RECT 24.572 219.294 24.676 223.668 ; 
        RECT 24.14 219.294 24.244 223.668 ; 
        RECT 23.708 219.294 23.812 223.668 ; 
        RECT 22.856 219.294 23.164 223.668 ; 
        RECT 15.284 219.294 15.592 223.668 ; 
        RECT 14.636 219.294 14.74 223.668 ; 
        RECT 14.204 219.294 14.308 223.668 ; 
        RECT 13.772 219.294 13.876 223.668 ; 
        RECT 13.34 219.294 13.444 223.668 ; 
        RECT 12.908 219.294 13.012 223.668 ; 
        RECT 12.476 219.294 12.58 223.668 ; 
        RECT 12.044 219.294 12.148 223.668 ; 
        RECT 11.612 219.294 11.716 223.668 ; 
        RECT 11.18 219.294 11.284 223.668 ; 
        RECT 10.748 219.294 10.852 223.668 ; 
        RECT 10.316 219.294 10.42 223.668 ; 
        RECT 9.884 219.294 9.988 223.668 ; 
        RECT 9.452 219.294 9.556 223.668 ; 
        RECT 9.02 219.294 9.124 223.668 ; 
        RECT 8.588 219.294 8.692 223.668 ; 
        RECT 8.156 219.294 8.26 223.668 ; 
        RECT 7.724 219.294 7.828 223.668 ; 
        RECT 7.292 219.294 7.396 223.668 ; 
        RECT 6.86 219.294 6.964 223.668 ; 
        RECT 6.428 219.294 6.532 223.668 ; 
        RECT 5.996 219.294 6.1 223.668 ; 
        RECT 5.564 219.294 5.668 223.668 ; 
        RECT 5.132 219.294 5.236 223.668 ; 
        RECT 4.7 219.294 4.804 223.668 ; 
        RECT 4.268 219.294 4.372 223.668 ; 
        RECT 3.836 219.294 3.94 223.668 ; 
        RECT 3.404 219.294 3.508 223.668 ; 
        RECT 2.972 219.294 3.076 223.668 ; 
        RECT 2.54 219.294 2.644 223.668 ; 
        RECT 2.108 219.294 2.212 223.668 ; 
        RECT 1.676 219.294 1.78 223.668 ; 
        RECT 1.244 219.294 1.348 223.668 ; 
        RECT 0.812 219.294 0.916 223.668 ; 
        RECT 0 219.294 0.34 223.668 ; 
        RECT 20.72 223.614 21.232 227.988 ; 
        RECT 20.664 226.276 21.232 227.566 ; 
        RECT 20.072 225.184 20.32 227.988 ; 
        RECT 20.016 226.422 20.32 227.036 ; 
        RECT 20.072 223.614 20.176 227.988 ; 
        RECT 20.072 224.098 20.232 225.056 ; 
        RECT 20.072 223.614 20.32 223.97 ; 
        RECT 18.884 225.416 19.708 227.988 ; 
        RECT 19.604 223.614 19.708 227.988 ; 
        RECT 18.884 226.524 19.764 227.556 ; 
        RECT 18.884 223.614 19.276 227.988 ; 
        RECT 17.216 223.614 17.548 227.988 ; 
        RECT 17.216 223.968 17.604 227.71 ; 
        RECT 38.108 223.614 38.448 227.988 ; 
        RECT 37.532 223.614 37.636 227.988 ; 
        RECT 37.1 223.614 37.204 227.988 ; 
        RECT 36.668 223.614 36.772 227.988 ; 
        RECT 36.236 223.614 36.34 227.988 ; 
        RECT 35.804 223.614 35.908 227.988 ; 
        RECT 35.372 223.614 35.476 227.988 ; 
        RECT 34.94 223.614 35.044 227.988 ; 
        RECT 34.508 223.614 34.612 227.988 ; 
        RECT 34.076 223.614 34.18 227.988 ; 
        RECT 33.644 223.614 33.748 227.988 ; 
        RECT 33.212 223.614 33.316 227.988 ; 
        RECT 32.78 223.614 32.884 227.988 ; 
        RECT 32.348 223.614 32.452 227.988 ; 
        RECT 31.916 223.614 32.02 227.988 ; 
        RECT 31.484 223.614 31.588 227.988 ; 
        RECT 31.052 223.614 31.156 227.988 ; 
        RECT 30.62 223.614 30.724 227.988 ; 
        RECT 30.188 223.614 30.292 227.988 ; 
        RECT 29.756 223.614 29.86 227.988 ; 
        RECT 29.324 223.614 29.428 227.988 ; 
        RECT 28.892 223.614 28.996 227.988 ; 
        RECT 28.46 223.614 28.564 227.988 ; 
        RECT 28.028 223.614 28.132 227.988 ; 
        RECT 27.596 223.614 27.7 227.988 ; 
        RECT 27.164 223.614 27.268 227.988 ; 
        RECT 26.732 223.614 26.836 227.988 ; 
        RECT 26.3 223.614 26.404 227.988 ; 
        RECT 25.868 223.614 25.972 227.988 ; 
        RECT 25.436 223.614 25.54 227.988 ; 
        RECT 25.004 223.614 25.108 227.988 ; 
        RECT 24.572 223.614 24.676 227.988 ; 
        RECT 24.14 223.614 24.244 227.988 ; 
        RECT 23.708 223.614 23.812 227.988 ; 
        RECT 22.856 223.614 23.164 227.988 ; 
        RECT 15.284 223.614 15.592 227.988 ; 
        RECT 14.636 223.614 14.74 227.988 ; 
        RECT 14.204 223.614 14.308 227.988 ; 
        RECT 13.772 223.614 13.876 227.988 ; 
        RECT 13.34 223.614 13.444 227.988 ; 
        RECT 12.908 223.614 13.012 227.988 ; 
        RECT 12.476 223.614 12.58 227.988 ; 
        RECT 12.044 223.614 12.148 227.988 ; 
        RECT 11.612 223.614 11.716 227.988 ; 
        RECT 11.18 223.614 11.284 227.988 ; 
        RECT 10.748 223.614 10.852 227.988 ; 
        RECT 10.316 223.614 10.42 227.988 ; 
        RECT 9.884 223.614 9.988 227.988 ; 
        RECT 9.452 223.614 9.556 227.988 ; 
        RECT 9.02 223.614 9.124 227.988 ; 
        RECT 8.588 223.614 8.692 227.988 ; 
        RECT 8.156 223.614 8.26 227.988 ; 
        RECT 7.724 223.614 7.828 227.988 ; 
        RECT 7.292 223.614 7.396 227.988 ; 
        RECT 6.86 223.614 6.964 227.988 ; 
        RECT 6.428 223.614 6.532 227.988 ; 
        RECT 5.996 223.614 6.1 227.988 ; 
        RECT 5.564 223.614 5.668 227.988 ; 
        RECT 5.132 223.614 5.236 227.988 ; 
        RECT 4.7 223.614 4.804 227.988 ; 
        RECT 4.268 223.614 4.372 227.988 ; 
        RECT 3.836 223.614 3.94 227.988 ; 
        RECT 3.404 223.614 3.508 227.988 ; 
        RECT 2.972 223.614 3.076 227.988 ; 
        RECT 2.54 223.614 2.644 227.988 ; 
        RECT 2.108 223.614 2.212 227.988 ; 
        RECT 1.676 223.614 1.78 227.988 ; 
        RECT 1.244 223.614 1.348 227.988 ; 
        RECT 0.812 223.614 0.916 227.988 ; 
        RECT 0 223.614 0.34 227.988 ; 
        RECT 20.72 227.934 21.232 232.308 ; 
        RECT 20.664 230.596 21.232 231.886 ; 
        RECT 20.072 229.504 20.32 232.308 ; 
        RECT 20.016 230.742 20.32 231.356 ; 
        RECT 20.072 227.934 20.176 232.308 ; 
        RECT 20.072 228.418 20.232 229.376 ; 
        RECT 20.072 227.934 20.32 228.29 ; 
        RECT 18.884 229.736 19.708 232.308 ; 
        RECT 19.604 227.934 19.708 232.308 ; 
        RECT 18.884 230.844 19.764 231.876 ; 
        RECT 18.884 227.934 19.276 232.308 ; 
        RECT 17.216 227.934 17.548 232.308 ; 
        RECT 17.216 228.288 17.604 232.03 ; 
        RECT 38.108 227.934 38.448 232.308 ; 
        RECT 37.532 227.934 37.636 232.308 ; 
        RECT 37.1 227.934 37.204 232.308 ; 
        RECT 36.668 227.934 36.772 232.308 ; 
        RECT 36.236 227.934 36.34 232.308 ; 
        RECT 35.804 227.934 35.908 232.308 ; 
        RECT 35.372 227.934 35.476 232.308 ; 
        RECT 34.94 227.934 35.044 232.308 ; 
        RECT 34.508 227.934 34.612 232.308 ; 
        RECT 34.076 227.934 34.18 232.308 ; 
        RECT 33.644 227.934 33.748 232.308 ; 
        RECT 33.212 227.934 33.316 232.308 ; 
        RECT 32.78 227.934 32.884 232.308 ; 
        RECT 32.348 227.934 32.452 232.308 ; 
        RECT 31.916 227.934 32.02 232.308 ; 
        RECT 31.484 227.934 31.588 232.308 ; 
        RECT 31.052 227.934 31.156 232.308 ; 
        RECT 30.62 227.934 30.724 232.308 ; 
        RECT 30.188 227.934 30.292 232.308 ; 
        RECT 29.756 227.934 29.86 232.308 ; 
        RECT 29.324 227.934 29.428 232.308 ; 
        RECT 28.892 227.934 28.996 232.308 ; 
        RECT 28.46 227.934 28.564 232.308 ; 
        RECT 28.028 227.934 28.132 232.308 ; 
        RECT 27.596 227.934 27.7 232.308 ; 
        RECT 27.164 227.934 27.268 232.308 ; 
        RECT 26.732 227.934 26.836 232.308 ; 
        RECT 26.3 227.934 26.404 232.308 ; 
        RECT 25.868 227.934 25.972 232.308 ; 
        RECT 25.436 227.934 25.54 232.308 ; 
        RECT 25.004 227.934 25.108 232.308 ; 
        RECT 24.572 227.934 24.676 232.308 ; 
        RECT 24.14 227.934 24.244 232.308 ; 
        RECT 23.708 227.934 23.812 232.308 ; 
        RECT 22.856 227.934 23.164 232.308 ; 
        RECT 15.284 227.934 15.592 232.308 ; 
        RECT 14.636 227.934 14.74 232.308 ; 
        RECT 14.204 227.934 14.308 232.308 ; 
        RECT 13.772 227.934 13.876 232.308 ; 
        RECT 13.34 227.934 13.444 232.308 ; 
        RECT 12.908 227.934 13.012 232.308 ; 
        RECT 12.476 227.934 12.58 232.308 ; 
        RECT 12.044 227.934 12.148 232.308 ; 
        RECT 11.612 227.934 11.716 232.308 ; 
        RECT 11.18 227.934 11.284 232.308 ; 
        RECT 10.748 227.934 10.852 232.308 ; 
        RECT 10.316 227.934 10.42 232.308 ; 
        RECT 9.884 227.934 9.988 232.308 ; 
        RECT 9.452 227.934 9.556 232.308 ; 
        RECT 9.02 227.934 9.124 232.308 ; 
        RECT 8.588 227.934 8.692 232.308 ; 
        RECT 8.156 227.934 8.26 232.308 ; 
        RECT 7.724 227.934 7.828 232.308 ; 
        RECT 7.292 227.934 7.396 232.308 ; 
        RECT 6.86 227.934 6.964 232.308 ; 
        RECT 6.428 227.934 6.532 232.308 ; 
        RECT 5.996 227.934 6.1 232.308 ; 
        RECT 5.564 227.934 5.668 232.308 ; 
        RECT 5.132 227.934 5.236 232.308 ; 
        RECT 4.7 227.934 4.804 232.308 ; 
        RECT 4.268 227.934 4.372 232.308 ; 
        RECT 3.836 227.934 3.94 232.308 ; 
        RECT 3.404 227.934 3.508 232.308 ; 
        RECT 2.972 227.934 3.076 232.308 ; 
        RECT 2.54 227.934 2.644 232.308 ; 
        RECT 2.108 227.934 2.212 232.308 ; 
        RECT 1.676 227.934 1.78 232.308 ; 
        RECT 1.244 227.934 1.348 232.308 ; 
        RECT 0.812 227.934 0.916 232.308 ; 
        RECT 0 227.934 0.34 232.308 ; 
        RECT 20.72 232.254 21.232 236.628 ; 
        RECT 20.664 234.916 21.232 236.206 ; 
        RECT 20.072 233.824 20.32 236.628 ; 
        RECT 20.016 235.062 20.32 235.676 ; 
        RECT 20.072 232.254 20.176 236.628 ; 
        RECT 20.072 232.738 20.232 233.696 ; 
        RECT 20.072 232.254 20.32 232.61 ; 
        RECT 18.884 234.056 19.708 236.628 ; 
        RECT 19.604 232.254 19.708 236.628 ; 
        RECT 18.884 235.164 19.764 236.196 ; 
        RECT 18.884 232.254 19.276 236.628 ; 
        RECT 17.216 232.254 17.548 236.628 ; 
        RECT 17.216 232.608 17.604 236.35 ; 
        RECT 38.108 232.254 38.448 236.628 ; 
        RECT 37.532 232.254 37.636 236.628 ; 
        RECT 37.1 232.254 37.204 236.628 ; 
        RECT 36.668 232.254 36.772 236.628 ; 
        RECT 36.236 232.254 36.34 236.628 ; 
        RECT 35.804 232.254 35.908 236.628 ; 
        RECT 35.372 232.254 35.476 236.628 ; 
        RECT 34.94 232.254 35.044 236.628 ; 
        RECT 34.508 232.254 34.612 236.628 ; 
        RECT 34.076 232.254 34.18 236.628 ; 
        RECT 33.644 232.254 33.748 236.628 ; 
        RECT 33.212 232.254 33.316 236.628 ; 
        RECT 32.78 232.254 32.884 236.628 ; 
        RECT 32.348 232.254 32.452 236.628 ; 
        RECT 31.916 232.254 32.02 236.628 ; 
        RECT 31.484 232.254 31.588 236.628 ; 
        RECT 31.052 232.254 31.156 236.628 ; 
        RECT 30.62 232.254 30.724 236.628 ; 
        RECT 30.188 232.254 30.292 236.628 ; 
        RECT 29.756 232.254 29.86 236.628 ; 
        RECT 29.324 232.254 29.428 236.628 ; 
        RECT 28.892 232.254 28.996 236.628 ; 
        RECT 28.46 232.254 28.564 236.628 ; 
        RECT 28.028 232.254 28.132 236.628 ; 
        RECT 27.596 232.254 27.7 236.628 ; 
        RECT 27.164 232.254 27.268 236.628 ; 
        RECT 26.732 232.254 26.836 236.628 ; 
        RECT 26.3 232.254 26.404 236.628 ; 
        RECT 25.868 232.254 25.972 236.628 ; 
        RECT 25.436 232.254 25.54 236.628 ; 
        RECT 25.004 232.254 25.108 236.628 ; 
        RECT 24.572 232.254 24.676 236.628 ; 
        RECT 24.14 232.254 24.244 236.628 ; 
        RECT 23.708 232.254 23.812 236.628 ; 
        RECT 22.856 232.254 23.164 236.628 ; 
        RECT 15.284 232.254 15.592 236.628 ; 
        RECT 14.636 232.254 14.74 236.628 ; 
        RECT 14.204 232.254 14.308 236.628 ; 
        RECT 13.772 232.254 13.876 236.628 ; 
        RECT 13.34 232.254 13.444 236.628 ; 
        RECT 12.908 232.254 13.012 236.628 ; 
        RECT 12.476 232.254 12.58 236.628 ; 
        RECT 12.044 232.254 12.148 236.628 ; 
        RECT 11.612 232.254 11.716 236.628 ; 
        RECT 11.18 232.254 11.284 236.628 ; 
        RECT 10.748 232.254 10.852 236.628 ; 
        RECT 10.316 232.254 10.42 236.628 ; 
        RECT 9.884 232.254 9.988 236.628 ; 
        RECT 9.452 232.254 9.556 236.628 ; 
        RECT 9.02 232.254 9.124 236.628 ; 
        RECT 8.588 232.254 8.692 236.628 ; 
        RECT 8.156 232.254 8.26 236.628 ; 
        RECT 7.724 232.254 7.828 236.628 ; 
        RECT 7.292 232.254 7.396 236.628 ; 
        RECT 6.86 232.254 6.964 236.628 ; 
        RECT 6.428 232.254 6.532 236.628 ; 
        RECT 5.996 232.254 6.1 236.628 ; 
        RECT 5.564 232.254 5.668 236.628 ; 
        RECT 5.132 232.254 5.236 236.628 ; 
        RECT 4.7 232.254 4.804 236.628 ; 
        RECT 4.268 232.254 4.372 236.628 ; 
        RECT 3.836 232.254 3.94 236.628 ; 
        RECT 3.404 232.254 3.508 236.628 ; 
        RECT 2.972 232.254 3.076 236.628 ; 
        RECT 2.54 232.254 2.644 236.628 ; 
        RECT 2.108 232.254 2.212 236.628 ; 
        RECT 1.676 232.254 1.78 236.628 ; 
        RECT 1.244 232.254 1.348 236.628 ; 
        RECT 0.812 232.254 0.916 236.628 ; 
        RECT 0 232.254 0.34 236.628 ; 
        RECT 20.72 236.574 21.232 240.948 ; 
        RECT 20.664 239.236 21.232 240.526 ; 
        RECT 20.072 238.144 20.32 240.948 ; 
        RECT 20.016 239.382 20.32 239.996 ; 
        RECT 20.072 236.574 20.176 240.948 ; 
        RECT 20.072 237.058 20.232 238.016 ; 
        RECT 20.072 236.574 20.32 236.93 ; 
        RECT 18.884 238.376 19.708 240.948 ; 
        RECT 19.604 236.574 19.708 240.948 ; 
        RECT 18.884 239.484 19.764 240.516 ; 
        RECT 18.884 236.574 19.276 240.948 ; 
        RECT 17.216 236.574 17.548 240.948 ; 
        RECT 17.216 236.928 17.604 240.67 ; 
        RECT 38.108 236.574 38.448 240.948 ; 
        RECT 37.532 236.574 37.636 240.948 ; 
        RECT 37.1 236.574 37.204 240.948 ; 
        RECT 36.668 236.574 36.772 240.948 ; 
        RECT 36.236 236.574 36.34 240.948 ; 
        RECT 35.804 236.574 35.908 240.948 ; 
        RECT 35.372 236.574 35.476 240.948 ; 
        RECT 34.94 236.574 35.044 240.948 ; 
        RECT 34.508 236.574 34.612 240.948 ; 
        RECT 34.076 236.574 34.18 240.948 ; 
        RECT 33.644 236.574 33.748 240.948 ; 
        RECT 33.212 236.574 33.316 240.948 ; 
        RECT 32.78 236.574 32.884 240.948 ; 
        RECT 32.348 236.574 32.452 240.948 ; 
        RECT 31.916 236.574 32.02 240.948 ; 
        RECT 31.484 236.574 31.588 240.948 ; 
        RECT 31.052 236.574 31.156 240.948 ; 
        RECT 30.62 236.574 30.724 240.948 ; 
        RECT 30.188 236.574 30.292 240.948 ; 
        RECT 29.756 236.574 29.86 240.948 ; 
        RECT 29.324 236.574 29.428 240.948 ; 
        RECT 28.892 236.574 28.996 240.948 ; 
        RECT 28.46 236.574 28.564 240.948 ; 
        RECT 28.028 236.574 28.132 240.948 ; 
        RECT 27.596 236.574 27.7 240.948 ; 
        RECT 27.164 236.574 27.268 240.948 ; 
        RECT 26.732 236.574 26.836 240.948 ; 
        RECT 26.3 236.574 26.404 240.948 ; 
        RECT 25.868 236.574 25.972 240.948 ; 
        RECT 25.436 236.574 25.54 240.948 ; 
        RECT 25.004 236.574 25.108 240.948 ; 
        RECT 24.572 236.574 24.676 240.948 ; 
        RECT 24.14 236.574 24.244 240.948 ; 
        RECT 23.708 236.574 23.812 240.948 ; 
        RECT 22.856 236.574 23.164 240.948 ; 
        RECT 15.284 236.574 15.592 240.948 ; 
        RECT 14.636 236.574 14.74 240.948 ; 
        RECT 14.204 236.574 14.308 240.948 ; 
        RECT 13.772 236.574 13.876 240.948 ; 
        RECT 13.34 236.574 13.444 240.948 ; 
        RECT 12.908 236.574 13.012 240.948 ; 
        RECT 12.476 236.574 12.58 240.948 ; 
        RECT 12.044 236.574 12.148 240.948 ; 
        RECT 11.612 236.574 11.716 240.948 ; 
        RECT 11.18 236.574 11.284 240.948 ; 
        RECT 10.748 236.574 10.852 240.948 ; 
        RECT 10.316 236.574 10.42 240.948 ; 
        RECT 9.884 236.574 9.988 240.948 ; 
        RECT 9.452 236.574 9.556 240.948 ; 
        RECT 9.02 236.574 9.124 240.948 ; 
        RECT 8.588 236.574 8.692 240.948 ; 
        RECT 8.156 236.574 8.26 240.948 ; 
        RECT 7.724 236.574 7.828 240.948 ; 
        RECT 7.292 236.574 7.396 240.948 ; 
        RECT 6.86 236.574 6.964 240.948 ; 
        RECT 6.428 236.574 6.532 240.948 ; 
        RECT 5.996 236.574 6.1 240.948 ; 
        RECT 5.564 236.574 5.668 240.948 ; 
        RECT 5.132 236.574 5.236 240.948 ; 
        RECT 4.7 236.574 4.804 240.948 ; 
        RECT 4.268 236.574 4.372 240.948 ; 
        RECT 3.836 236.574 3.94 240.948 ; 
        RECT 3.404 236.574 3.508 240.948 ; 
        RECT 2.972 236.574 3.076 240.948 ; 
        RECT 2.54 236.574 2.644 240.948 ; 
        RECT 2.108 236.574 2.212 240.948 ; 
        RECT 1.676 236.574 1.78 240.948 ; 
        RECT 1.244 236.574 1.348 240.948 ; 
        RECT 0.812 236.574 0.916 240.948 ; 
        RECT 0 236.574 0.34 240.948 ; 
        RECT 20.72 240.894 21.232 245.268 ; 
        RECT 20.664 243.556 21.232 244.846 ; 
        RECT 20.072 242.464 20.32 245.268 ; 
        RECT 20.016 243.702 20.32 244.316 ; 
        RECT 20.072 240.894 20.176 245.268 ; 
        RECT 20.072 241.378 20.232 242.336 ; 
        RECT 20.072 240.894 20.32 241.25 ; 
        RECT 18.884 242.696 19.708 245.268 ; 
        RECT 19.604 240.894 19.708 245.268 ; 
        RECT 18.884 243.804 19.764 244.836 ; 
        RECT 18.884 240.894 19.276 245.268 ; 
        RECT 17.216 240.894 17.548 245.268 ; 
        RECT 17.216 241.248 17.604 244.99 ; 
        RECT 38.108 240.894 38.448 245.268 ; 
        RECT 37.532 240.894 37.636 245.268 ; 
        RECT 37.1 240.894 37.204 245.268 ; 
        RECT 36.668 240.894 36.772 245.268 ; 
        RECT 36.236 240.894 36.34 245.268 ; 
        RECT 35.804 240.894 35.908 245.268 ; 
        RECT 35.372 240.894 35.476 245.268 ; 
        RECT 34.94 240.894 35.044 245.268 ; 
        RECT 34.508 240.894 34.612 245.268 ; 
        RECT 34.076 240.894 34.18 245.268 ; 
        RECT 33.644 240.894 33.748 245.268 ; 
        RECT 33.212 240.894 33.316 245.268 ; 
        RECT 32.78 240.894 32.884 245.268 ; 
        RECT 32.348 240.894 32.452 245.268 ; 
        RECT 31.916 240.894 32.02 245.268 ; 
        RECT 31.484 240.894 31.588 245.268 ; 
        RECT 31.052 240.894 31.156 245.268 ; 
        RECT 30.62 240.894 30.724 245.268 ; 
        RECT 30.188 240.894 30.292 245.268 ; 
        RECT 29.756 240.894 29.86 245.268 ; 
        RECT 29.324 240.894 29.428 245.268 ; 
        RECT 28.892 240.894 28.996 245.268 ; 
        RECT 28.46 240.894 28.564 245.268 ; 
        RECT 28.028 240.894 28.132 245.268 ; 
        RECT 27.596 240.894 27.7 245.268 ; 
        RECT 27.164 240.894 27.268 245.268 ; 
        RECT 26.732 240.894 26.836 245.268 ; 
        RECT 26.3 240.894 26.404 245.268 ; 
        RECT 25.868 240.894 25.972 245.268 ; 
        RECT 25.436 240.894 25.54 245.268 ; 
        RECT 25.004 240.894 25.108 245.268 ; 
        RECT 24.572 240.894 24.676 245.268 ; 
        RECT 24.14 240.894 24.244 245.268 ; 
        RECT 23.708 240.894 23.812 245.268 ; 
        RECT 22.856 240.894 23.164 245.268 ; 
        RECT 15.284 240.894 15.592 245.268 ; 
        RECT 14.636 240.894 14.74 245.268 ; 
        RECT 14.204 240.894 14.308 245.268 ; 
        RECT 13.772 240.894 13.876 245.268 ; 
        RECT 13.34 240.894 13.444 245.268 ; 
        RECT 12.908 240.894 13.012 245.268 ; 
        RECT 12.476 240.894 12.58 245.268 ; 
        RECT 12.044 240.894 12.148 245.268 ; 
        RECT 11.612 240.894 11.716 245.268 ; 
        RECT 11.18 240.894 11.284 245.268 ; 
        RECT 10.748 240.894 10.852 245.268 ; 
        RECT 10.316 240.894 10.42 245.268 ; 
        RECT 9.884 240.894 9.988 245.268 ; 
        RECT 9.452 240.894 9.556 245.268 ; 
        RECT 9.02 240.894 9.124 245.268 ; 
        RECT 8.588 240.894 8.692 245.268 ; 
        RECT 8.156 240.894 8.26 245.268 ; 
        RECT 7.724 240.894 7.828 245.268 ; 
        RECT 7.292 240.894 7.396 245.268 ; 
        RECT 6.86 240.894 6.964 245.268 ; 
        RECT 6.428 240.894 6.532 245.268 ; 
        RECT 5.996 240.894 6.1 245.268 ; 
        RECT 5.564 240.894 5.668 245.268 ; 
        RECT 5.132 240.894 5.236 245.268 ; 
        RECT 4.7 240.894 4.804 245.268 ; 
        RECT 4.268 240.894 4.372 245.268 ; 
        RECT 3.836 240.894 3.94 245.268 ; 
        RECT 3.404 240.894 3.508 245.268 ; 
        RECT 2.972 240.894 3.076 245.268 ; 
        RECT 2.54 240.894 2.644 245.268 ; 
        RECT 2.108 240.894 2.212 245.268 ; 
        RECT 1.676 240.894 1.78 245.268 ; 
        RECT 1.244 240.894 1.348 245.268 ; 
        RECT 0.812 240.894 0.916 245.268 ; 
        RECT 0 240.894 0.34 245.268 ; 
        RECT 20.72 245.214 21.232 249.588 ; 
        RECT 20.664 247.876 21.232 249.166 ; 
        RECT 20.072 246.784 20.32 249.588 ; 
        RECT 20.016 248.022 20.32 248.636 ; 
        RECT 20.072 245.214 20.176 249.588 ; 
        RECT 20.072 245.698 20.232 246.656 ; 
        RECT 20.072 245.214 20.32 245.57 ; 
        RECT 18.884 247.016 19.708 249.588 ; 
        RECT 19.604 245.214 19.708 249.588 ; 
        RECT 18.884 248.124 19.764 249.156 ; 
        RECT 18.884 245.214 19.276 249.588 ; 
        RECT 17.216 245.214 17.548 249.588 ; 
        RECT 17.216 245.568 17.604 249.31 ; 
        RECT 38.108 245.214 38.448 249.588 ; 
        RECT 37.532 245.214 37.636 249.588 ; 
        RECT 37.1 245.214 37.204 249.588 ; 
        RECT 36.668 245.214 36.772 249.588 ; 
        RECT 36.236 245.214 36.34 249.588 ; 
        RECT 35.804 245.214 35.908 249.588 ; 
        RECT 35.372 245.214 35.476 249.588 ; 
        RECT 34.94 245.214 35.044 249.588 ; 
        RECT 34.508 245.214 34.612 249.588 ; 
        RECT 34.076 245.214 34.18 249.588 ; 
        RECT 33.644 245.214 33.748 249.588 ; 
        RECT 33.212 245.214 33.316 249.588 ; 
        RECT 32.78 245.214 32.884 249.588 ; 
        RECT 32.348 245.214 32.452 249.588 ; 
        RECT 31.916 245.214 32.02 249.588 ; 
        RECT 31.484 245.214 31.588 249.588 ; 
        RECT 31.052 245.214 31.156 249.588 ; 
        RECT 30.62 245.214 30.724 249.588 ; 
        RECT 30.188 245.214 30.292 249.588 ; 
        RECT 29.756 245.214 29.86 249.588 ; 
        RECT 29.324 245.214 29.428 249.588 ; 
        RECT 28.892 245.214 28.996 249.588 ; 
        RECT 28.46 245.214 28.564 249.588 ; 
        RECT 28.028 245.214 28.132 249.588 ; 
        RECT 27.596 245.214 27.7 249.588 ; 
        RECT 27.164 245.214 27.268 249.588 ; 
        RECT 26.732 245.214 26.836 249.588 ; 
        RECT 26.3 245.214 26.404 249.588 ; 
        RECT 25.868 245.214 25.972 249.588 ; 
        RECT 25.436 245.214 25.54 249.588 ; 
        RECT 25.004 245.214 25.108 249.588 ; 
        RECT 24.572 245.214 24.676 249.588 ; 
        RECT 24.14 245.214 24.244 249.588 ; 
        RECT 23.708 245.214 23.812 249.588 ; 
        RECT 22.856 245.214 23.164 249.588 ; 
        RECT 15.284 245.214 15.592 249.588 ; 
        RECT 14.636 245.214 14.74 249.588 ; 
        RECT 14.204 245.214 14.308 249.588 ; 
        RECT 13.772 245.214 13.876 249.588 ; 
        RECT 13.34 245.214 13.444 249.588 ; 
        RECT 12.908 245.214 13.012 249.588 ; 
        RECT 12.476 245.214 12.58 249.588 ; 
        RECT 12.044 245.214 12.148 249.588 ; 
        RECT 11.612 245.214 11.716 249.588 ; 
        RECT 11.18 245.214 11.284 249.588 ; 
        RECT 10.748 245.214 10.852 249.588 ; 
        RECT 10.316 245.214 10.42 249.588 ; 
        RECT 9.884 245.214 9.988 249.588 ; 
        RECT 9.452 245.214 9.556 249.588 ; 
        RECT 9.02 245.214 9.124 249.588 ; 
        RECT 8.588 245.214 8.692 249.588 ; 
        RECT 8.156 245.214 8.26 249.588 ; 
        RECT 7.724 245.214 7.828 249.588 ; 
        RECT 7.292 245.214 7.396 249.588 ; 
        RECT 6.86 245.214 6.964 249.588 ; 
        RECT 6.428 245.214 6.532 249.588 ; 
        RECT 5.996 245.214 6.1 249.588 ; 
        RECT 5.564 245.214 5.668 249.588 ; 
        RECT 5.132 245.214 5.236 249.588 ; 
        RECT 4.7 245.214 4.804 249.588 ; 
        RECT 4.268 245.214 4.372 249.588 ; 
        RECT 3.836 245.214 3.94 249.588 ; 
        RECT 3.404 245.214 3.508 249.588 ; 
        RECT 2.972 245.214 3.076 249.588 ; 
        RECT 2.54 245.214 2.644 249.588 ; 
        RECT 2.108 245.214 2.212 249.588 ; 
        RECT 1.676 245.214 1.78 249.588 ; 
        RECT 1.244 245.214 1.348 249.588 ; 
        RECT 0.812 245.214 0.916 249.588 ; 
        RECT 0 245.214 0.34 249.588 ; 
        RECT 20.72 249.534 21.232 253.908 ; 
        RECT 20.664 252.196 21.232 253.486 ; 
        RECT 20.072 251.104 20.32 253.908 ; 
        RECT 20.016 252.342 20.32 252.956 ; 
        RECT 20.072 249.534 20.176 253.908 ; 
        RECT 20.072 250.018 20.232 250.976 ; 
        RECT 20.072 249.534 20.32 249.89 ; 
        RECT 18.884 251.336 19.708 253.908 ; 
        RECT 19.604 249.534 19.708 253.908 ; 
        RECT 18.884 252.444 19.764 253.476 ; 
        RECT 18.884 249.534 19.276 253.908 ; 
        RECT 17.216 249.534 17.548 253.908 ; 
        RECT 17.216 249.888 17.604 253.63 ; 
        RECT 38.108 249.534 38.448 253.908 ; 
        RECT 37.532 249.534 37.636 253.908 ; 
        RECT 37.1 249.534 37.204 253.908 ; 
        RECT 36.668 249.534 36.772 253.908 ; 
        RECT 36.236 249.534 36.34 253.908 ; 
        RECT 35.804 249.534 35.908 253.908 ; 
        RECT 35.372 249.534 35.476 253.908 ; 
        RECT 34.94 249.534 35.044 253.908 ; 
        RECT 34.508 249.534 34.612 253.908 ; 
        RECT 34.076 249.534 34.18 253.908 ; 
        RECT 33.644 249.534 33.748 253.908 ; 
        RECT 33.212 249.534 33.316 253.908 ; 
        RECT 32.78 249.534 32.884 253.908 ; 
        RECT 32.348 249.534 32.452 253.908 ; 
        RECT 31.916 249.534 32.02 253.908 ; 
        RECT 31.484 249.534 31.588 253.908 ; 
        RECT 31.052 249.534 31.156 253.908 ; 
        RECT 30.62 249.534 30.724 253.908 ; 
        RECT 30.188 249.534 30.292 253.908 ; 
        RECT 29.756 249.534 29.86 253.908 ; 
        RECT 29.324 249.534 29.428 253.908 ; 
        RECT 28.892 249.534 28.996 253.908 ; 
        RECT 28.46 249.534 28.564 253.908 ; 
        RECT 28.028 249.534 28.132 253.908 ; 
        RECT 27.596 249.534 27.7 253.908 ; 
        RECT 27.164 249.534 27.268 253.908 ; 
        RECT 26.732 249.534 26.836 253.908 ; 
        RECT 26.3 249.534 26.404 253.908 ; 
        RECT 25.868 249.534 25.972 253.908 ; 
        RECT 25.436 249.534 25.54 253.908 ; 
        RECT 25.004 249.534 25.108 253.908 ; 
        RECT 24.572 249.534 24.676 253.908 ; 
        RECT 24.14 249.534 24.244 253.908 ; 
        RECT 23.708 249.534 23.812 253.908 ; 
        RECT 22.856 249.534 23.164 253.908 ; 
        RECT 15.284 249.534 15.592 253.908 ; 
        RECT 14.636 249.534 14.74 253.908 ; 
        RECT 14.204 249.534 14.308 253.908 ; 
        RECT 13.772 249.534 13.876 253.908 ; 
        RECT 13.34 249.534 13.444 253.908 ; 
        RECT 12.908 249.534 13.012 253.908 ; 
        RECT 12.476 249.534 12.58 253.908 ; 
        RECT 12.044 249.534 12.148 253.908 ; 
        RECT 11.612 249.534 11.716 253.908 ; 
        RECT 11.18 249.534 11.284 253.908 ; 
        RECT 10.748 249.534 10.852 253.908 ; 
        RECT 10.316 249.534 10.42 253.908 ; 
        RECT 9.884 249.534 9.988 253.908 ; 
        RECT 9.452 249.534 9.556 253.908 ; 
        RECT 9.02 249.534 9.124 253.908 ; 
        RECT 8.588 249.534 8.692 253.908 ; 
        RECT 8.156 249.534 8.26 253.908 ; 
        RECT 7.724 249.534 7.828 253.908 ; 
        RECT 7.292 249.534 7.396 253.908 ; 
        RECT 6.86 249.534 6.964 253.908 ; 
        RECT 6.428 249.534 6.532 253.908 ; 
        RECT 5.996 249.534 6.1 253.908 ; 
        RECT 5.564 249.534 5.668 253.908 ; 
        RECT 5.132 249.534 5.236 253.908 ; 
        RECT 4.7 249.534 4.804 253.908 ; 
        RECT 4.268 249.534 4.372 253.908 ; 
        RECT 3.836 249.534 3.94 253.908 ; 
        RECT 3.404 249.534 3.508 253.908 ; 
        RECT 2.972 249.534 3.076 253.908 ; 
        RECT 2.54 249.534 2.644 253.908 ; 
        RECT 2.108 249.534 2.212 253.908 ; 
        RECT 1.676 249.534 1.78 253.908 ; 
        RECT 1.244 249.534 1.348 253.908 ; 
        RECT 0.812 249.534 0.916 253.908 ; 
        RECT 0 249.534 0.34 253.908 ; 
        RECT 20.72 253.854 21.232 258.228 ; 
        RECT 20.664 256.516 21.232 257.806 ; 
        RECT 20.072 255.424 20.32 258.228 ; 
        RECT 20.016 256.662 20.32 257.276 ; 
        RECT 20.072 253.854 20.176 258.228 ; 
        RECT 20.072 254.338 20.232 255.296 ; 
        RECT 20.072 253.854 20.32 254.21 ; 
        RECT 18.884 255.656 19.708 258.228 ; 
        RECT 19.604 253.854 19.708 258.228 ; 
        RECT 18.884 256.764 19.764 257.796 ; 
        RECT 18.884 253.854 19.276 258.228 ; 
        RECT 17.216 253.854 17.548 258.228 ; 
        RECT 17.216 254.208 17.604 257.95 ; 
        RECT 38.108 253.854 38.448 258.228 ; 
        RECT 37.532 253.854 37.636 258.228 ; 
        RECT 37.1 253.854 37.204 258.228 ; 
        RECT 36.668 253.854 36.772 258.228 ; 
        RECT 36.236 253.854 36.34 258.228 ; 
        RECT 35.804 253.854 35.908 258.228 ; 
        RECT 35.372 253.854 35.476 258.228 ; 
        RECT 34.94 253.854 35.044 258.228 ; 
        RECT 34.508 253.854 34.612 258.228 ; 
        RECT 34.076 253.854 34.18 258.228 ; 
        RECT 33.644 253.854 33.748 258.228 ; 
        RECT 33.212 253.854 33.316 258.228 ; 
        RECT 32.78 253.854 32.884 258.228 ; 
        RECT 32.348 253.854 32.452 258.228 ; 
        RECT 31.916 253.854 32.02 258.228 ; 
        RECT 31.484 253.854 31.588 258.228 ; 
        RECT 31.052 253.854 31.156 258.228 ; 
        RECT 30.62 253.854 30.724 258.228 ; 
        RECT 30.188 253.854 30.292 258.228 ; 
        RECT 29.756 253.854 29.86 258.228 ; 
        RECT 29.324 253.854 29.428 258.228 ; 
        RECT 28.892 253.854 28.996 258.228 ; 
        RECT 28.46 253.854 28.564 258.228 ; 
        RECT 28.028 253.854 28.132 258.228 ; 
        RECT 27.596 253.854 27.7 258.228 ; 
        RECT 27.164 253.854 27.268 258.228 ; 
        RECT 26.732 253.854 26.836 258.228 ; 
        RECT 26.3 253.854 26.404 258.228 ; 
        RECT 25.868 253.854 25.972 258.228 ; 
        RECT 25.436 253.854 25.54 258.228 ; 
        RECT 25.004 253.854 25.108 258.228 ; 
        RECT 24.572 253.854 24.676 258.228 ; 
        RECT 24.14 253.854 24.244 258.228 ; 
        RECT 23.708 253.854 23.812 258.228 ; 
        RECT 22.856 253.854 23.164 258.228 ; 
        RECT 15.284 253.854 15.592 258.228 ; 
        RECT 14.636 253.854 14.74 258.228 ; 
        RECT 14.204 253.854 14.308 258.228 ; 
        RECT 13.772 253.854 13.876 258.228 ; 
        RECT 13.34 253.854 13.444 258.228 ; 
        RECT 12.908 253.854 13.012 258.228 ; 
        RECT 12.476 253.854 12.58 258.228 ; 
        RECT 12.044 253.854 12.148 258.228 ; 
        RECT 11.612 253.854 11.716 258.228 ; 
        RECT 11.18 253.854 11.284 258.228 ; 
        RECT 10.748 253.854 10.852 258.228 ; 
        RECT 10.316 253.854 10.42 258.228 ; 
        RECT 9.884 253.854 9.988 258.228 ; 
        RECT 9.452 253.854 9.556 258.228 ; 
        RECT 9.02 253.854 9.124 258.228 ; 
        RECT 8.588 253.854 8.692 258.228 ; 
        RECT 8.156 253.854 8.26 258.228 ; 
        RECT 7.724 253.854 7.828 258.228 ; 
        RECT 7.292 253.854 7.396 258.228 ; 
        RECT 6.86 253.854 6.964 258.228 ; 
        RECT 6.428 253.854 6.532 258.228 ; 
        RECT 5.996 253.854 6.1 258.228 ; 
        RECT 5.564 253.854 5.668 258.228 ; 
        RECT 5.132 253.854 5.236 258.228 ; 
        RECT 4.7 253.854 4.804 258.228 ; 
        RECT 4.268 253.854 4.372 258.228 ; 
        RECT 3.836 253.854 3.94 258.228 ; 
        RECT 3.404 253.854 3.508 258.228 ; 
        RECT 2.972 253.854 3.076 258.228 ; 
        RECT 2.54 253.854 2.644 258.228 ; 
        RECT 2.108 253.854 2.212 258.228 ; 
        RECT 1.676 253.854 1.78 258.228 ; 
        RECT 1.244 253.854 1.348 258.228 ; 
        RECT 0.812 253.854 0.916 258.228 ; 
        RECT 0 253.854 0.34 258.228 ; 
        RECT 20.72 258.174 21.232 262.548 ; 
        RECT 20.664 260.836 21.232 262.126 ; 
        RECT 20.072 259.744 20.32 262.548 ; 
        RECT 20.016 260.982 20.32 261.596 ; 
        RECT 20.072 258.174 20.176 262.548 ; 
        RECT 20.072 258.658 20.232 259.616 ; 
        RECT 20.072 258.174 20.32 258.53 ; 
        RECT 18.884 259.976 19.708 262.548 ; 
        RECT 19.604 258.174 19.708 262.548 ; 
        RECT 18.884 261.084 19.764 262.116 ; 
        RECT 18.884 258.174 19.276 262.548 ; 
        RECT 17.216 258.174 17.548 262.548 ; 
        RECT 17.216 258.528 17.604 262.27 ; 
        RECT 38.108 258.174 38.448 262.548 ; 
        RECT 37.532 258.174 37.636 262.548 ; 
        RECT 37.1 258.174 37.204 262.548 ; 
        RECT 36.668 258.174 36.772 262.548 ; 
        RECT 36.236 258.174 36.34 262.548 ; 
        RECT 35.804 258.174 35.908 262.548 ; 
        RECT 35.372 258.174 35.476 262.548 ; 
        RECT 34.94 258.174 35.044 262.548 ; 
        RECT 34.508 258.174 34.612 262.548 ; 
        RECT 34.076 258.174 34.18 262.548 ; 
        RECT 33.644 258.174 33.748 262.548 ; 
        RECT 33.212 258.174 33.316 262.548 ; 
        RECT 32.78 258.174 32.884 262.548 ; 
        RECT 32.348 258.174 32.452 262.548 ; 
        RECT 31.916 258.174 32.02 262.548 ; 
        RECT 31.484 258.174 31.588 262.548 ; 
        RECT 31.052 258.174 31.156 262.548 ; 
        RECT 30.62 258.174 30.724 262.548 ; 
        RECT 30.188 258.174 30.292 262.548 ; 
        RECT 29.756 258.174 29.86 262.548 ; 
        RECT 29.324 258.174 29.428 262.548 ; 
        RECT 28.892 258.174 28.996 262.548 ; 
        RECT 28.46 258.174 28.564 262.548 ; 
        RECT 28.028 258.174 28.132 262.548 ; 
        RECT 27.596 258.174 27.7 262.548 ; 
        RECT 27.164 258.174 27.268 262.548 ; 
        RECT 26.732 258.174 26.836 262.548 ; 
        RECT 26.3 258.174 26.404 262.548 ; 
        RECT 25.868 258.174 25.972 262.548 ; 
        RECT 25.436 258.174 25.54 262.548 ; 
        RECT 25.004 258.174 25.108 262.548 ; 
        RECT 24.572 258.174 24.676 262.548 ; 
        RECT 24.14 258.174 24.244 262.548 ; 
        RECT 23.708 258.174 23.812 262.548 ; 
        RECT 22.856 258.174 23.164 262.548 ; 
        RECT 15.284 258.174 15.592 262.548 ; 
        RECT 14.636 258.174 14.74 262.548 ; 
        RECT 14.204 258.174 14.308 262.548 ; 
        RECT 13.772 258.174 13.876 262.548 ; 
        RECT 13.34 258.174 13.444 262.548 ; 
        RECT 12.908 258.174 13.012 262.548 ; 
        RECT 12.476 258.174 12.58 262.548 ; 
        RECT 12.044 258.174 12.148 262.548 ; 
        RECT 11.612 258.174 11.716 262.548 ; 
        RECT 11.18 258.174 11.284 262.548 ; 
        RECT 10.748 258.174 10.852 262.548 ; 
        RECT 10.316 258.174 10.42 262.548 ; 
        RECT 9.884 258.174 9.988 262.548 ; 
        RECT 9.452 258.174 9.556 262.548 ; 
        RECT 9.02 258.174 9.124 262.548 ; 
        RECT 8.588 258.174 8.692 262.548 ; 
        RECT 8.156 258.174 8.26 262.548 ; 
        RECT 7.724 258.174 7.828 262.548 ; 
        RECT 7.292 258.174 7.396 262.548 ; 
        RECT 6.86 258.174 6.964 262.548 ; 
        RECT 6.428 258.174 6.532 262.548 ; 
        RECT 5.996 258.174 6.1 262.548 ; 
        RECT 5.564 258.174 5.668 262.548 ; 
        RECT 5.132 258.174 5.236 262.548 ; 
        RECT 4.7 258.174 4.804 262.548 ; 
        RECT 4.268 258.174 4.372 262.548 ; 
        RECT 3.836 258.174 3.94 262.548 ; 
        RECT 3.404 258.174 3.508 262.548 ; 
        RECT 2.972 258.174 3.076 262.548 ; 
        RECT 2.54 258.174 2.644 262.548 ; 
        RECT 2.108 258.174 2.212 262.548 ; 
        RECT 1.676 258.174 1.78 262.548 ; 
        RECT 1.244 258.174 1.348 262.548 ; 
        RECT 0.812 258.174 0.916 262.548 ; 
        RECT 0 258.174 0.34 262.548 ; 
        RECT 20.72 262.494 21.232 266.868 ; 
        RECT 20.664 265.156 21.232 266.446 ; 
        RECT 20.072 264.064 20.32 266.868 ; 
        RECT 20.016 265.302 20.32 265.916 ; 
        RECT 20.072 262.494 20.176 266.868 ; 
        RECT 20.072 262.978 20.232 263.936 ; 
        RECT 20.072 262.494 20.32 262.85 ; 
        RECT 18.884 264.296 19.708 266.868 ; 
        RECT 19.604 262.494 19.708 266.868 ; 
        RECT 18.884 265.404 19.764 266.436 ; 
        RECT 18.884 262.494 19.276 266.868 ; 
        RECT 17.216 262.494 17.548 266.868 ; 
        RECT 17.216 262.848 17.604 266.59 ; 
        RECT 38.108 262.494 38.448 266.868 ; 
        RECT 37.532 262.494 37.636 266.868 ; 
        RECT 37.1 262.494 37.204 266.868 ; 
        RECT 36.668 262.494 36.772 266.868 ; 
        RECT 36.236 262.494 36.34 266.868 ; 
        RECT 35.804 262.494 35.908 266.868 ; 
        RECT 35.372 262.494 35.476 266.868 ; 
        RECT 34.94 262.494 35.044 266.868 ; 
        RECT 34.508 262.494 34.612 266.868 ; 
        RECT 34.076 262.494 34.18 266.868 ; 
        RECT 33.644 262.494 33.748 266.868 ; 
        RECT 33.212 262.494 33.316 266.868 ; 
        RECT 32.78 262.494 32.884 266.868 ; 
        RECT 32.348 262.494 32.452 266.868 ; 
        RECT 31.916 262.494 32.02 266.868 ; 
        RECT 31.484 262.494 31.588 266.868 ; 
        RECT 31.052 262.494 31.156 266.868 ; 
        RECT 30.62 262.494 30.724 266.868 ; 
        RECT 30.188 262.494 30.292 266.868 ; 
        RECT 29.756 262.494 29.86 266.868 ; 
        RECT 29.324 262.494 29.428 266.868 ; 
        RECT 28.892 262.494 28.996 266.868 ; 
        RECT 28.46 262.494 28.564 266.868 ; 
        RECT 28.028 262.494 28.132 266.868 ; 
        RECT 27.596 262.494 27.7 266.868 ; 
        RECT 27.164 262.494 27.268 266.868 ; 
        RECT 26.732 262.494 26.836 266.868 ; 
        RECT 26.3 262.494 26.404 266.868 ; 
        RECT 25.868 262.494 25.972 266.868 ; 
        RECT 25.436 262.494 25.54 266.868 ; 
        RECT 25.004 262.494 25.108 266.868 ; 
        RECT 24.572 262.494 24.676 266.868 ; 
        RECT 24.14 262.494 24.244 266.868 ; 
        RECT 23.708 262.494 23.812 266.868 ; 
        RECT 22.856 262.494 23.164 266.868 ; 
        RECT 15.284 262.494 15.592 266.868 ; 
        RECT 14.636 262.494 14.74 266.868 ; 
        RECT 14.204 262.494 14.308 266.868 ; 
        RECT 13.772 262.494 13.876 266.868 ; 
        RECT 13.34 262.494 13.444 266.868 ; 
        RECT 12.908 262.494 13.012 266.868 ; 
        RECT 12.476 262.494 12.58 266.868 ; 
        RECT 12.044 262.494 12.148 266.868 ; 
        RECT 11.612 262.494 11.716 266.868 ; 
        RECT 11.18 262.494 11.284 266.868 ; 
        RECT 10.748 262.494 10.852 266.868 ; 
        RECT 10.316 262.494 10.42 266.868 ; 
        RECT 9.884 262.494 9.988 266.868 ; 
        RECT 9.452 262.494 9.556 266.868 ; 
        RECT 9.02 262.494 9.124 266.868 ; 
        RECT 8.588 262.494 8.692 266.868 ; 
        RECT 8.156 262.494 8.26 266.868 ; 
        RECT 7.724 262.494 7.828 266.868 ; 
        RECT 7.292 262.494 7.396 266.868 ; 
        RECT 6.86 262.494 6.964 266.868 ; 
        RECT 6.428 262.494 6.532 266.868 ; 
        RECT 5.996 262.494 6.1 266.868 ; 
        RECT 5.564 262.494 5.668 266.868 ; 
        RECT 5.132 262.494 5.236 266.868 ; 
        RECT 4.7 262.494 4.804 266.868 ; 
        RECT 4.268 262.494 4.372 266.868 ; 
        RECT 3.836 262.494 3.94 266.868 ; 
        RECT 3.404 262.494 3.508 266.868 ; 
        RECT 2.972 262.494 3.076 266.868 ; 
        RECT 2.54 262.494 2.644 266.868 ; 
        RECT 2.108 262.494 2.212 266.868 ; 
        RECT 1.676 262.494 1.78 266.868 ; 
        RECT 1.244 262.494 1.348 266.868 ; 
        RECT 0.812 262.494 0.916 266.868 ; 
        RECT 0 262.494 0.34 266.868 ; 
        RECT 20.72 266.814 21.232 271.188 ; 
        RECT 20.664 269.476 21.232 270.766 ; 
        RECT 20.072 268.384 20.32 271.188 ; 
        RECT 20.016 269.622 20.32 270.236 ; 
        RECT 20.072 266.814 20.176 271.188 ; 
        RECT 20.072 267.298 20.232 268.256 ; 
        RECT 20.072 266.814 20.32 267.17 ; 
        RECT 18.884 268.616 19.708 271.188 ; 
        RECT 19.604 266.814 19.708 271.188 ; 
        RECT 18.884 269.724 19.764 270.756 ; 
        RECT 18.884 266.814 19.276 271.188 ; 
        RECT 17.216 266.814 17.548 271.188 ; 
        RECT 17.216 267.168 17.604 270.91 ; 
        RECT 38.108 266.814 38.448 271.188 ; 
        RECT 37.532 266.814 37.636 271.188 ; 
        RECT 37.1 266.814 37.204 271.188 ; 
        RECT 36.668 266.814 36.772 271.188 ; 
        RECT 36.236 266.814 36.34 271.188 ; 
        RECT 35.804 266.814 35.908 271.188 ; 
        RECT 35.372 266.814 35.476 271.188 ; 
        RECT 34.94 266.814 35.044 271.188 ; 
        RECT 34.508 266.814 34.612 271.188 ; 
        RECT 34.076 266.814 34.18 271.188 ; 
        RECT 33.644 266.814 33.748 271.188 ; 
        RECT 33.212 266.814 33.316 271.188 ; 
        RECT 32.78 266.814 32.884 271.188 ; 
        RECT 32.348 266.814 32.452 271.188 ; 
        RECT 31.916 266.814 32.02 271.188 ; 
        RECT 31.484 266.814 31.588 271.188 ; 
        RECT 31.052 266.814 31.156 271.188 ; 
        RECT 30.62 266.814 30.724 271.188 ; 
        RECT 30.188 266.814 30.292 271.188 ; 
        RECT 29.756 266.814 29.86 271.188 ; 
        RECT 29.324 266.814 29.428 271.188 ; 
        RECT 28.892 266.814 28.996 271.188 ; 
        RECT 28.46 266.814 28.564 271.188 ; 
        RECT 28.028 266.814 28.132 271.188 ; 
        RECT 27.596 266.814 27.7 271.188 ; 
        RECT 27.164 266.814 27.268 271.188 ; 
        RECT 26.732 266.814 26.836 271.188 ; 
        RECT 26.3 266.814 26.404 271.188 ; 
        RECT 25.868 266.814 25.972 271.188 ; 
        RECT 25.436 266.814 25.54 271.188 ; 
        RECT 25.004 266.814 25.108 271.188 ; 
        RECT 24.572 266.814 24.676 271.188 ; 
        RECT 24.14 266.814 24.244 271.188 ; 
        RECT 23.708 266.814 23.812 271.188 ; 
        RECT 22.856 266.814 23.164 271.188 ; 
        RECT 15.284 266.814 15.592 271.188 ; 
        RECT 14.636 266.814 14.74 271.188 ; 
        RECT 14.204 266.814 14.308 271.188 ; 
        RECT 13.772 266.814 13.876 271.188 ; 
        RECT 13.34 266.814 13.444 271.188 ; 
        RECT 12.908 266.814 13.012 271.188 ; 
        RECT 12.476 266.814 12.58 271.188 ; 
        RECT 12.044 266.814 12.148 271.188 ; 
        RECT 11.612 266.814 11.716 271.188 ; 
        RECT 11.18 266.814 11.284 271.188 ; 
        RECT 10.748 266.814 10.852 271.188 ; 
        RECT 10.316 266.814 10.42 271.188 ; 
        RECT 9.884 266.814 9.988 271.188 ; 
        RECT 9.452 266.814 9.556 271.188 ; 
        RECT 9.02 266.814 9.124 271.188 ; 
        RECT 8.588 266.814 8.692 271.188 ; 
        RECT 8.156 266.814 8.26 271.188 ; 
        RECT 7.724 266.814 7.828 271.188 ; 
        RECT 7.292 266.814 7.396 271.188 ; 
        RECT 6.86 266.814 6.964 271.188 ; 
        RECT 6.428 266.814 6.532 271.188 ; 
        RECT 5.996 266.814 6.1 271.188 ; 
        RECT 5.564 266.814 5.668 271.188 ; 
        RECT 5.132 266.814 5.236 271.188 ; 
        RECT 4.7 266.814 4.804 271.188 ; 
        RECT 4.268 266.814 4.372 271.188 ; 
        RECT 3.836 266.814 3.94 271.188 ; 
        RECT 3.404 266.814 3.508 271.188 ; 
        RECT 2.972 266.814 3.076 271.188 ; 
        RECT 2.54 266.814 2.644 271.188 ; 
        RECT 2.108 266.814 2.212 271.188 ; 
        RECT 1.676 266.814 1.78 271.188 ; 
        RECT 1.244 266.814 1.348 271.188 ; 
        RECT 0.812 266.814 0.916 271.188 ; 
        RECT 0 266.814 0.34 271.188 ; 
        RECT 20.72 271.134 21.232 275.508 ; 
        RECT 20.664 273.796 21.232 275.086 ; 
        RECT 20.072 272.704 20.32 275.508 ; 
        RECT 20.016 273.942 20.32 274.556 ; 
        RECT 20.072 271.134 20.176 275.508 ; 
        RECT 20.072 271.618 20.232 272.576 ; 
        RECT 20.072 271.134 20.32 271.49 ; 
        RECT 18.884 272.936 19.708 275.508 ; 
        RECT 19.604 271.134 19.708 275.508 ; 
        RECT 18.884 274.044 19.764 275.076 ; 
        RECT 18.884 271.134 19.276 275.508 ; 
        RECT 17.216 271.134 17.548 275.508 ; 
        RECT 17.216 271.488 17.604 275.23 ; 
        RECT 38.108 271.134 38.448 275.508 ; 
        RECT 37.532 271.134 37.636 275.508 ; 
        RECT 37.1 271.134 37.204 275.508 ; 
        RECT 36.668 271.134 36.772 275.508 ; 
        RECT 36.236 271.134 36.34 275.508 ; 
        RECT 35.804 271.134 35.908 275.508 ; 
        RECT 35.372 271.134 35.476 275.508 ; 
        RECT 34.94 271.134 35.044 275.508 ; 
        RECT 34.508 271.134 34.612 275.508 ; 
        RECT 34.076 271.134 34.18 275.508 ; 
        RECT 33.644 271.134 33.748 275.508 ; 
        RECT 33.212 271.134 33.316 275.508 ; 
        RECT 32.78 271.134 32.884 275.508 ; 
        RECT 32.348 271.134 32.452 275.508 ; 
        RECT 31.916 271.134 32.02 275.508 ; 
        RECT 31.484 271.134 31.588 275.508 ; 
        RECT 31.052 271.134 31.156 275.508 ; 
        RECT 30.62 271.134 30.724 275.508 ; 
        RECT 30.188 271.134 30.292 275.508 ; 
        RECT 29.756 271.134 29.86 275.508 ; 
        RECT 29.324 271.134 29.428 275.508 ; 
        RECT 28.892 271.134 28.996 275.508 ; 
        RECT 28.46 271.134 28.564 275.508 ; 
        RECT 28.028 271.134 28.132 275.508 ; 
        RECT 27.596 271.134 27.7 275.508 ; 
        RECT 27.164 271.134 27.268 275.508 ; 
        RECT 26.732 271.134 26.836 275.508 ; 
        RECT 26.3 271.134 26.404 275.508 ; 
        RECT 25.868 271.134 25.972 275.508 ; 
        RECT 25.436 271.134 25.54 275.508 ; 
        RECT 25.004 271.134 25.108 275.508 ; 
        RECT 24.572 271.134 24.676 275.508 ; 
        RECT 24.14 271.134 24.244 275.508 ; 
        RECT 23.708 271.134 23.812 275.508 ; 
        RECT 22.856 271.134 23.164 275.508 ; 
        RECT 15.284 271.134 15.592 275.508 ; 
        RECT 14.636 271.134 14.74 275.508 ; 
        RECT 14.204 271.134 14.308 275.508 ; 
        RECT 13.772 271.134 13.876 275.508 ; 
        RECT 13.34 271.134 13.444 275.508 ; 
        RECT 12.908 271.134 13.012 275.508 ; 
        RECT 12.476 271.134 12.58 275.508 ; 
        RECT 12.044 271.134 12.148 275.508 ; 
        RECT 11.612 271.134 11.716 275.508 ; 
        RECT 11.18 271.134 11.284 275.508 ; 
        RECT 10.748 271.134 10.852 275.508 ; 
        RECT 10.316 271.134 10.42 275.508 ; 
        RECT 9.884 271.134 9.988 275.508 ; 
        RECT 9.452 271.134 9.556 275.508 ; 
        RECT 9.02 271.134 9.124 275.508 ; 
        RECT 8.588 271.134 8.692 275.508 ; 
        RECT 8.156 271.134 8.26 275.508 ; 
        RECT 7.724 271.134 7.828 275.508 ; 
        RECT 7.292 271.134 7.396 275.508 ; 
        RECT 6.86 271.134 6.964 275.508 ; 
        RECT 6.428 271.134 6.532 275.508 ; 
        RECT 5.996 271.134 6.1 275.508 ; 
        RECT 5.564 271.134 5.668 275.508 ; 
        RECT 5.132 271.134 5.236 275.508 ; 
        RECT 4.7 271.134 4.804 275.508 ; 
        RECT 4.268 271.134 4.372 275.508 ; 
        RECT 3.836 271.134 3.94 275.508 ; 
        RECT 3.404 271.134 3.508 275.508 ; 
        RECT 2.972 271.134 3.076 275.508 ; 
        RECT 2.54 271.134 2.644 275.508 ; 
        RECT 2.108 271.134 2.212 275.508 ; 
        RECT 1.676 271.134 1.78 275.508 ; 
        RECT 1.244 271.134 1.348 275.508 ; 
        RECT 0.812 271.134 0.916 275.508 ; 
        RECT 0 271.134 0.34 275.508 ; 
        RECT 20.72 275.454 21.232 279.828 ; 
        RECT 20.664 278.116 21.232 279.406 ; 
        RECT 20.072 277.024 20.32 279.828 ; 
        RECT 20.016 278.262 20.32 278.876 ; 
        RECT 20.072 275.454 20.176 279.828 ; 
        RECT 20.072 275.938 20.232 276.896 ; 
        RECT 20.072 275.454 20.32 275.81 ; 
        RECT 18.884 277.256 19.708 279.828 ; 
        RECT 19.604 275.454 19.708 279.828 ; 
        RECT 18.884 278.364 19.764 279.396 ; 
        RECT 18.884 275.454 19.276 279.828 ; 
        RECT 17.216 275.454 17.548 279.828 ; 
        RECT 17.216 275.808 17.604 279.55 ; 
        RECT 38.108 275.454 38.448 279.828 ; 
        RECT 37.532 275.454 37.636 279.828 ; 
        RECT 37.1 275.454 37.204 279.828 ; 
        RECT 36.668 275.454 36.772 279.828 ; 
        RECT 36.236 275.454 36.34 279.828 ; 
        RECT 35.804 275.454 35.908 279.828 ; 
        RECT 35.372 275.454 35.476 279.828 ; 
        RECT 34.94 275.454 35.044 279.828 ; 
        RECT 34.508 275.454 34.612 279.828 ; 
        RECT 34.076 275.454 34.18 279.828 ; 
        RECT 33.644 275.454 33.748 279.828 ; 
        RECT 33.212 275.454 33.316 279.828 ; 
        RECT 32.78 275.454 32.884 279.828 ; 
        RECT 32.348 275.454 32.452 279.828 ; 
        RECT 31.916 275.454 32.02 279.828 ; 
        RECT 31.484 275.454 31.588 279.828 ; 
        RECT 31.052 275.454 31.156 279.828 ; 
        RECT 30.62 275.454 30.724 279.828 ; 
        RECT 30.188 275.454 30.292 279.828 ; 
        RECT 29.756 275.454 29.86 279.828 ; 
        RECT 29.324 275.454 29.428 279.828 ; 
        RECT 28.892 275.454 28.996 279.828 ; 
        RECT 28.46 275.454 28.564 279.828 ; 
        RECT 28.028 275.454 28.132 279.828 ; 
        RECT 27.596 275.454 27.7 279.828 ; 
        RECT 27.164 275.454 27.268 279.828 ; 
        RECT 26.732 275.454 26.836 279.828 ; 
        RECT 26.3 275.454 26.404 279.828 ; 
        RECT 25.868 275.454 25.972 279.828 ; 
        RECT 25.436 275.454 25.54 279.828 ; 
        RECT 25.004 275.454 25.108 279.828 ; 
        RECT 24.572 275.454 24.676 279.828 ; 
        RECT 24.14 275.454 24.244 279.828 ; 
        RECT 23.708 275.454 23.812 279.828 ; 
        RECT 22.856 275.454 23.164 279.828 ; 
        RECT 15.284 275.454 15.592 279.828 ; 
        RECT 14.636 275.454 14.74 279.828 ; 
        RECT 14.204 275.454 14.308 279.828 ; 
        RECT 13.772 275.454 13.876 279.828 ; 
        RECT 13.34 275.454 13.444 279.828 ; 
        RECT 12.908 275.454 13.012 279.828 ; 
        RECT 12.476 275.454 12.58 279.828 ; 
        RECT 12.044 275.454 12.148 279.828 ; 
        RECT 11.612 275.454 11.716 279.828 ; 
        RECT 11.18 275.454 11.284 279.828 ; 
        RECT 10.748 275.454 10.852 279.828 ; 
        RECT 10.316 275.454 10.42 279.828 ; 
        RECT 9.884 275.454 9.988 279.828 ; 
        RECT 9.452 275.454 9.556 279.828 ; 
        RECT 9.02 275.454 9.124 279.828 ; 
        RECT 8.588 275.454 8.692 279.828 ; 
        RECT 8.156 275.454 8.26 279.828 ; 
        RECT 7.724 275.454 7.828 279.828 ; 
        RECT 7.292 275.454 7.396 279.828 ; 
        RECT 6.86 275.454 6.964 279.828 ; 
        RECT 6.428 275.454 6.532 279.828 ; 
        RECT 5.996 275.454 6.1 279.828 ; 
        RECT 5.564 275.454 5.668 279.828 ; 
        RECT 5.132 275.454 5.236 279.828 ; 
        RECT 4.7 275.454 4.804 279.828 ; 
        RECT 4.268 275.454 4.372 279.828 ; 
        RECT 3.836 275.454 3.94 279.828 ; 
        RECT 3.404 275.454 3.508 279.828 ; 
        RECT 2.972 275.454 3.076 279.828 ; 
        RECT 2.54 275.454 2.644 279.828 ; 
        RECT 2.108 275.454 2.212 279.828 ; 
        RECT 1.676 275.454 1.78 279.828 ; 
        RECT 1.244 275.454 1.348 279.828 ; 
        RECT 0.812 275.454 0.916 279.828 ; 
        RECT 0 275.454 0.34 279.828 ; 
        RECT 20.72 279.774 21.232 284.148 ; 
        RECT 20.664 282.436 21.232 283.726 ; 
        RECT 20.072 281.344 20.32 284.148 ; 
        RECT 20.016 282.582 20.32 283.196 ; 
        RECT 20.072 279.774 20.176 284.148 ; 
        RECT 20.072 280.258 20.232 281.216 ; 
        RECT 20.072 279.774 20.32 280.13 ; 
        RECT 18.884 281.576 19.708 284.148 ; 
        RECT 19.604 279.774 19.708 284.148 ; 
        RECT 18.884 282.684 19.764 283.716 ; 
        RECT 18.884 279.774 19.276 284.148 ; 
        RECT 17.216 279.774 17.548 284.148 ; 
        RECT 17.216 280.128 17.604 283.87 ; 
        RECT 38.108 279.774 38.448 284.148 ; 
        RECT 37.532 279.774 37.636 284.148 ; 
        RECT 37.1 279.774 37.204 284.148 ; 
        RECT 36.668 279.774 36.772 284.148 ; 
        RECT 36.236 279.774 36.34 284.148 ; 
        RECT 35.804 279.774 35.908 284.148 ; 
        RECT 35.372 279.774 35.476 284.148 ; 
        RECT 34.94 279.774 35.044 284.148 ; 
        RECT 34.508 279.774 34.612 284.148 ; 
        RECT 34.076 279.774 34.18 284.148 ; 
        RECT 33.644 279.774 33.748 284.148 ; 
        RECT 33.212 279.774 33.316 284.148 ; 
        RECT 32.78 279.774 32.884 284.148 ; 
        RECT 32.348 279.774 32.452 284.148 ; 
        RECT 31.916 279.774 32.02 284.148 ; 
        RECT 31.484 279.774 31.588 284.148 ; 
        RECT 31.052 279.774 31.156 284.148 ; 
        RECT 30.62 279.774 30.724 284.148 ; 
        RECT 30.188 279.774 30.292 284.148 ; 
        RECT 29.756 279.774 29.86 284.148 ; 
        RECT 29.324 279.774 29.428 284.148 ; 
        RECT 28.892 279.774 28.996 284.148 ; 
        RECT 28.46 279.774 28.564 284.148 ; 
        RECT 28.028 279.774 28.132 284.148 ; 
        RECT 27.596 279.774 27.7 284.148 ; 
        RECT 27.164 279.774 27.268 284.148 ; 
        RECT 26.732 279.774 26.836 284.148 ; 
        RECT 26.3 279.774 26.404 284.148 ; 
        RECT 25.868 279.774 25.972 284.148 ; 
        RECT 25.436 279.774 25.54 284.148 ; 
        RECT 25.004 279.774 25.108 284.148 ; 
        RECT 24.572 279.774 24.676 284.148 ; 
        RECT 24.14 279.774 24.244 284.148 ; 
        RECT 23.708 279.774 23.812 284.148 ; 
        RECT 22.856 279.774 23.164 284.148 ; 
        RECT 15.284 279.774 15.592 284.148 ; 
        RECT 14.636 279.774 14.74 284.148 ; 
        RECT 14.204 279.774 14.308 284.148 ; 
        RECT 13.772 279.774 13.876 284.148 ; 
        RECT 13.34 279.774 13.444 284.148 ; 
        RECT 12.908 279.774 13.012 284.148 ; 
        RECT 12.476 279.774 12.58 284.148 ; 
        RECT 12.044 279.774 12.148 284.148 ; 
        RECT 11.612 279.774 11.716 284.148 ; 
        RECT 11.18 279.774 11.284 284.148 ; 
        RECT 10.748 279.774 10.852 284.148 ; 
        RECT 10.316 279.774 10.42 284.148 ; 
        RECT 9.884 279.774 9.988 284.148 ; 
        RECT 9.452 279.774 9.556 284.148 ; 
        RECT 9.02 279.774 9.124 284.148 ; 
        RECT 8.588 279.774 8.692 284.148 ; 
        RECT 8.156 279.774 8.26 284.148 ; 
        RECT 7.724 279.774 7.828 284.148 ; 
        RECT 7.292 279.774 7.396 284.148 ; 
        RECT 6.86 279.774 6.964 284.148 ; 
        RECT 6.428 279.774 6.532 284.148 ; 
        RECT 5.996 279.774 6.1 284.148 ; 
        RECT 5.564 279.774 5.668 284.148 ; 
        RECT 5.132 279.774 5.236 284.148 ; 
        RECT 4.7 279.774 4.804 284.148 ; 
        RECT 4.268 279.774 4.372 284.148 ; 
        RECT 3.836 279.774 3.94 284.148 ; 
        RECT 3.404 279.774 3.508 284.148 ; 
        RECT 2.972 279.774 3.076 284.148 ; 
        RECT 2.54 279.774 2.644 284.148 ; 
        RECT 2.108 279.774 2.212 284.148 ; 
        RECT 1.676 279.774 1.78 284.148 ; 
        RECT 1.244 279.774 1.348 284.148 ; 
        RECT 0.812 279.774 0.916 284.148 ; 
        RECT 0 279.774 0.34 284.148 ; 
        RECT 20.72 284.094 21.232 288.468 ; 
        RECT 20.664 286.756 21.232 288.046 ; 
        RECT 20.072 285.664 20.32 288.468 ; 
        RECT 20.016 286.902 20.32 287.516 ; 
        RECT 20.072 284.094 20.176 288.468 ; 
        RECT 20.072 284.578 20.232 285.536 ; 
        RECT 20.072 284.094 20.32 284.45 ; 
        RECT 18.884 285.896 19.708 288.468 ; 
        RECT 19.604 284.094 19.708 288.468 ; 
        RECT 18.884 287.004 19.764 288.036 ; 
        RECT 18.884 284.094 19.276 288.468 ; 
        RECT 17.216 284.094 17.548 288.468 ; 
        RECT 17.216 284.448 17.604 288.19 ; 
        RECT 38.108 284.094 38.448 288.468 ; 
        RECT 37.532 284.094 37.636 288.468 ; 
        RECT 37.1 284.094 37.204 288.468 ; 
        RECT 36.668 284.094 36.772 288.468 ; 
        RECT 36.236 284.094 36.34 288.468 ; 
        RECT 35.804 284.094 35.908 288.468 ; 
        RECT 35.372 284.094 35.476 288.468 ; 
        RECT 34.94 284.094 35.044 288.468 ; 
        RECT 34.508 284.094 34.612 288.468 ; 
        RECT 34.076 284.094 34.18 288.468 ; 
        RECT 33.644 284.094 33.748 288.468 ; 
        RECT 33.212 284.094 33.316 288.468 ; 
        RECT 32.78 284.094 32.884 288.468 ; 
        RECT 32.348 284.094 32.452 288.468 ; 
        RECT 31.916 284.094 32.02 288.468 ; 
        RECT 31.484 284.094 31.588 288.468 ; 
        RECT 31.052 284.094 31.156 288.468 ; 
        RECT 30.62 284.094 30.724 288.468 ; 
        RECT 30.188 284.094 30.292 288.468 ; 
        RECT 29.756 284.094 29.86 288.468 ; 
        RECT 29.324 284.094 29.428 288.468 ; 
        RECT 28.892 284.094 28.996 288.468 ; 
        RECT 28.46 284.094 28.564 288.468 ; 
        RECT 28.028 284.094 28.132 288.468 ; 
        RECT 27.596 284.094 27.7 288.468 ; 
        RECT 27.164 284.094 27.268 288.468 ; 
        RECT 26.732 284.094 26.836 288.468 ; 
        RECT 26.3 284.094 26.404 288.468 ; 
        RECT 25.868 284.094 25.972 288.468 ; 
        RECT 25.436 284.094 25.54 288.468 ; 
        RECT 25.004 284.094 25.108 288.468 ; 
        RECT 24.572 284.094 24.676 288.468 ; 
        RECT 24.14 284.094 24.244 288.468 ; 
        RECT 23.708 284.094 23.812 288.468 ; 
        RECT 22.856 284.094 23.164 288.468 ; 
        RECT 15.284 284.094 15.592 288.468 ; 
        RECT 14.636 284.094 14.74 288.468 ; 
        RECT 14.204 284.094 14.308 288.468 ; 
        RECT 13.772 284.094 13.876 288.468 ; 
        RECT 13.34 284.094 13.444 288.468 ; 
        RECT 12.908 284.094 13.012 288.468 ; 
        RECT 12.476 284.094 12.58 288.468 ; 
        RECT 12.044 284.094 12.148 288.468 ; 
        RECT 11.612 284.094 11.716 288.468 ; 
        RECT 11.18 284.094 11.284 288.468 ; 
        RECT 10.748 284.094 10.852 288.468 ; 
        RECT 10.316 284.094 10.42 288.468 ; 
        RECT 9.884 284.094 9.988 288.468 ; 
        RECT 9.452 284.094 9.556 288.468 ; 
        RECT 9.02 284.094 9.124 288.468 ; 
        RECT 8.588 284.094 8.692 288.468 ; 
        RECT 8.156 284.094 8.26 288.468 ; 
        RECT 7.724 284.094 7.828 288.468 ; 
        RECT 7.292 284.094 7.396 288.468 ; 
        RECT 6.86 284.094 6.964 288.468 ; 
        RECT 6.428 284.094 6.532 288.468 ; 
        RECT 5.996 284.094 6.1 288.468 ; 
        RECT 5.564 284.094 5.668 288.468 ; 
        RECT 5.132 284.094 5.236 288.468 ; 
        RECT 4.7 284.094 4.804 288.468 ; 
        RECT 4.268 284.094 4.372 288.468 ; 
        RECT 3.836 284.094 3.94 288.468 ; 
        RECT 3.404 284.094 3.508 288.468 ; 
        RECT 2.972 284.094 3.076 288.468 ; 
        RECT 2.54 284.094 2.644 288.468 ; 
        RECT 2.108 284.094 2.212 288.468 ; 
        RECT 1.676 284.094 1.78 288.468 ; 
        RECT 1.244 284.094 1.348 288.468 ; 
        RECT 0.812 284.094 0.916 288.468 ; 
        RECT 0 284.094 0.34 288.468 ; 
        RECT 20.72 288.414 21.232 292.788 ; 
        RECT 20.664 291.076 21.232 292.366 ; 
        RECT 20.072 289.984 20.32 292.788 ; 
        RECT 20.016 291.222 20.32 291.836 ; 
        RECT 20.072 288.414 20.176 292.788 ; 
        RECT 20.072 288.898 20.232 289.856 ; 
        RECT 20.072 288.414 20.32 288.77 ; 
        RECT 18.884 290.216 19.708 292.788 ; 
        RECT 19.604 288.414 19.708 292.788 ; 
        RECT 18.884 291.324 19.764 292.356 ; 
        RECT 18.884 288.414 19.276 292.788 ; 
        RECT 17.216 288.414 17.548 292.788 ; 
        RECT 17.216 288.768 17.604 292.51 ; 
        RECT 38.108 288.414 38.448 292.788 ; 
        RECT 37.532 288.414 37.636 292.788 ; 
        RECT 37.1 288.414 37.204 292.788 ; 
        RECT 36.668 288.414 36.772 292.788 ; 
        RECT 36.236 288.414 36.34 292.788 ; 
        RECT 35.804 288.414 35.908 292.788 ; 
        RECT 35.372 288.414 35.476 292.788 ; 
        RECT 34.94 288.414 35.044 292.788 ; 
        RECT 34.508 288.414 34.612 292.788 ; 
        RECT 34.076 288.414 34.18 292.788 ; 
        RECT 33.644 288.414 33.748 292.788 ; 
        RECT 33.212 288.414 33.316 292.788 ; 
        RECT 32.78 288.414 32.884 292.788 ; 
        RECT 32.348 288.414 32.452 292.788 ; 
        RECT 31.916 288.414 32.02 292.788 ; 
        RECT 31.484 288.414 31.588 292.788 ; 
        RECT 31.052 288.414 31.156 292.788 ; 
        RECT 30.62 288.414 30.724 292.788 ; 
        RECT 30.188 288.414 30.292 292.788 ; 
        RECT 29.756 288.414 29.86 292.788 ; 
        RECT 29.324 288.414 29.428 292.788 ; 
        RECT 28.892 288.414 28.996 292.788 ; 
        RECT 28.46 288.414 28.564 292.788 ; 
        RECT 28.028 288.414 28.132 292.788 ; 
        RECT 27.596 288.414 27.7 292.788 ; 
        RECT 27.164 288.414 27.268 292.788 ; 
        RECT 26.732 288.414 26.836 292.788 ; 
        RECT 26.3 288.414 26.404 292.788 ; 
        RECT 25.868 288.414 25.972 292.788 ; 
        RECT 25.436 288.414 25.54 292.788 ; 
        RECT 25.004 288.414 25.108 292.788 ; 
        RECT 24.572 288.414 24.676 292.788 ; 
        RECT 24.14 288.414 24.244 292.788 ; 
        RECT 23.708 288.414 23.812 292.788 ; 
        RECT 22.856 288.414 23.164 292.788 ; 
        RECT 15.284 288.414 15.592 292.788 ; 
        RECT 14.636 288.414 14.74 292.788 ; 
        RECT 14.204 288.414 14.308 292.788 ; 
        RECT 13.772 288.414 13.876 292.788 ; 
        RECT 13.34 288.414 13.444 292.788 ; 
        RECT 12.908 288.414 13.012 292.788 ; 
        RECT 12.476 288.414 12.58 292.788 ; 
        RECT 12.044 288.414 12.148 292.788 ; 
        RECT 11.612 288.414 11.716 292.788 ; 
        RECT 11.18 288.414 11.284 292.788 ; 
        RECT 10.748 288.414 10.852 292.788 ; 
        RECT 10.316 288.414 10.42 292.788 ; 
        RECT 9.884 288.414 9.988 292.788 ; 
        RECT 9.452 288.414 9.556 292.788 ; 
        RECT 9.02 288.414 9.124 292.788 ; 
        RECT 8.588 288.414 8.692 292.788 ; 
        RECT 8.156 288.414 8.26 292.788 ; 
        RECT 7.724 288.414 7.828 292.788 ; 
        RECT 7.292 288.414 7.396 292.788 ; 
        RECT 6.86 288.414 6.964 292.788 ; 
        RECT 6.428 288.414 6.532 292.788 ; 
        RECT 5.996 288.414 6.1 292.788 ; 
        RECT 5.564 288.414 5.668 292.788 ; 
        RECT 5.132 288.414 5.236 292.788 ; 
        RECT 4.7 288.414 4.804 292.788 ; 
        RECT 4.268 288.414 4.372 292.788 ; 
        RECT 3.836 288.414 3.94 292.788 ; 
        RECT 3.404 288.414 3.508 292.788 ; 
        RECT 2.972 288.414 3.076 292.788 ; 
        RECT 2.54 288.414 2.644 292.788 ; 
        RECT 2.108 288.414 2.212 292.788 ; 
        RECT 1.676 288.414 1.78 292.788 ; 
        RECT 1.244 288.414 1.348 292.788 ; 
        RECT 0.812 288.414 0.916 292.788 ; 
        RECT 0 288.414 0.34 292.788 ; 
        RECT 20.72 292.734 21.232 297.108 ; 
        RECT 20.664 295.396 21.232 296.686 ; 
        RECT 20.072 294.304 20.32 297.108 ; 
        RECT 20.016 295.542 20.32 296.156 ; 
        RECT 20.072 292.734 20.176 297.108 ; 
        RECT 20.072 293.218 20.232 294.176 ; 
        RECT 20.072 292.734 20.32 293.09 ; 
        RECT 18.884 294.536 19.708 297.108 ; 
        RECT 19.604 292.734 19.708 297.108 ; 
        RECT 18.884 295.644 19.764 296.676 ; 
        RECT 18.884 292.734 19.276 297.108 ; 
        RECT 17.216 292.734 17.548 297.108 ; 
        RECT 17.216 293.088 17.604 296.83 ; 
        RECT 38.108 292.734 38.448 297.108 ; 
        RECT 37.532 292.734 37.636 297.108 ; 
        RECT 37.1 292.734 37.204 297.108 ; 
        RECT 36.668 292.734 36.772 297.108 ; 
        RECT 36.236 292.734 36.34 297.108 ; 
        RECT 35.804 292.734 35.908 297.108 ; 
        RECT 35.372 292.734 35.476 297.108 ; 
        RECT 34.94 292.734 35.044 297.108 ; 
        RECT 34.508 292.734 34.612 297.108 ; 
        RECT 34.076 292.734 34.18 297.108 ; 
        RECT 33.644 292.734 33.748 297.108 ; 
        RECT 33.212 292.734 33.316 297.108 ; 
        RECT 32.78 292.734 32.884 297.108 ; 
        RECT 32.348 292.734 32.452 297.108 ; 
        RECT 31.916 292.734 32.02 297.108 ; 
        RECT 31.484 292.734 31.588 297.108 ; 
        RECT 31.052 292.734 31.156 297.108 ; 
        RECT 30.62 292.734 30.724 297.108 ; 
        RECT 30.188 292.734 30.292 297.108 ; 
        RECT 29.756 292.734 29.86 297.108 ; 
        RECT 29.324 292.734 29.428 297.108 ; 
        RECT 28.892 292.734 28.996 297.108 ; 
        RECT 28.46 292.734 28.564 297.108 ; 
        RECT 28.028 292.734 28.132 297.108 ; 
        RECT 27.596 292.734 27.7 297.108 ; 
        RECT 27.164 292.734 27.268 297.108 ; 
        RECT 26.732 292.734 26.836 297.108 ; 
        RECT 26.3 292.734 26.404 297.108 ; 
        RECT 25.868 292.734 25.972 297.108 ; 
        RECT 25.436 292.734 25.54 297.108 ; 
        RECT 25.004 292.734 25.108 297.108 ; 
        RECT 24.572 292.734 24.676 297.108 ; 
        RECT 24.14 292.734 24.244 297.108 ; 
        RECT 23.708 292.734 23.812 297.108 ; 
        RECT 22.856 292.734 23.164 297.108 ; 
        RECT 15.284 292.734 15.592 297.108 ; 
        RECT 14.636 292.734 14.74 297.108 ; 
        RECT 14.204 292.734 14.308 297.108 ; 
        RECT 13.772 292.734 13.876 297.108 ; 
        RECT 13.34 292.734 13.444 297.108 ; 
        RECT 12.908 292.734 13.012 297.108 ; 
        RECT 12.476 292.734 12.58 297.108 ; 
        RECT 12.044 292.734 12.148 297.108 ; 
        RECT 11.612 292.734 11.716 297.108 ; 
        RECT 11.18 292.734 11.284 297.108 ; 
        RECT 10.748 292.734 10.852 297.108 ; 
        RECT 10.316 292.734 10.42 297.108 ; 
        RECT 9.884 292.734 9.988 297.108 ; 
        RECT 9.452 292.734 9.556 297.108 ; 
        RECT 9.02 292.734 9.124 297.108 ; 
        RECT 8.588 292.734 8.692 297.108 ; 
        RECT 8.156 292.734 8.26 297.108 ; 
        RECT 7.724 292.734 7.828 297.108 ; 
        RECT 7.292 292.734 7.396 297.108 ; 
        RECT 6.86 292.734 6.964 297.108 ; 
        RECT 6.428 292.734 6.532 297.108 ; 
        RECT 5.996 292.734 6.1 297.108 ; 
        RECT 5.564 292.734 5.668 297.108 ; 
        RECT 5.132 292.734 5.236 297.108 ; 
        RECT 4.7 292.734 4.804 297.108 ; 
        RECT 4.268 292.734 4.372 297.108 ; 
        RECT 3.836 292.734 3.94 297.108 ; 
        RECT 3.404 292.734 3.508 297.108 ; 
        RECT 2.972 292.734 3.076 297.108 ; 
        RECT 2.54 292.734 2.644 297.108 ; 
        RECT 2.108 292.734 2.212 297.108 ; 
        RECT 1.676 292.734 1.78 297.108 ; 
        RECT 1.244 292.734 1.348 297.108 ; 
        RECT 0.812 292.734 0.916 297.108 ; 
        RECT 0 292.734 0.34 297.108 ; 
        RECT 20.72 297.054 21.232 301.428 ; 
        RECT 20.664 299.716 21.232 301.006 ; 
        RECT 20.072 298.624 20.32 301.428 ; 
        RECT 20.016 299.862 20.32 300.476 ; 
        RECT 20.072 297.054 20.176 301.428 ; 
        RECT 20.072 297.538 20.232 298.496 ; 
        RECT 20.072 297.054 20.32 297.41 ; 
        RECT 18.884 298.856 19.708 301.428 ; 
        RECT 19.604 297.054 19.708 301.428 ; 
        RECT 18.884 299.964 19.764 300.996 ; 
        RECT 18.884 297.054 19.276 301.428 ; 
        RECT 17.216 297.054 17.548 301.428 ; 
        RECT 17.216 297.408 17.604 301.15 ; 
        RECT 38.108 297.054 38.448 301.428 ; 
        RECT 37.532 297.054 37.636 301.428 ; 
        RECT 37.1 297.054 37.204 301.428 ; 
        RECT 36.668 297.054 36.772 301.428 ; 
        RECT 36.236 297.054 36.34 301.428 ; 
        RECT 35.804 297.054 35.908 301.428 ; 
        RECT 35.372 297.054 35.476 301.428 ; 
        RECT 34.94 297.054 35.044 301.428 ; 
        RECT 34.508 297.054 34.612 301.428 ; 
        RECT 34.076 297.054 34.18 301.428 ; 
        RECT 33.644 297.054 33.748 301.428 ; 
        RECT 33.212 297.054 33.316 301.428 ; 
        RECT 32.78 297.054 32.884 301.428 ; 
        RECT 32.348 297.054 32.452 301.428 ; 
        RECT 31.916 297.054 32.02 301.428 ; 
        RECT 31.484 297.054 31.588 301.428 ; 
        RECT 31.052 297.054 31.156 301.428 ; 
        RECT 30.62 297.054 30.724 301.428 ; 
        RECT 30.188 297.054 30.292 301.428 ; 
        RECT 29.756 297.054 29.86 301.428 ; 
        RECT 29.324 297.054 29.428 301.428 ; 
        RECT 28.892 297.054 28.996 301.428 ; 
        RECT 28.46 297.054 28.564 301.428 ; 
        RECT 28.028 297.054 28.132 301.428 ; 
        RECT 27.596 297.054 27.7 301.428 ; 
        RECT 27.164 297.054 27.268 301.428 ; 
        RECT 26.732 297.054 26.836 301.428 ; 
        RECT 26.3 297.054 26.404 301.428 ; 
        RECT 25.868 297.054 25.972 301.428 ; 
        RECT 25.436 297.054 25.54 301.428 ; 
        RECT 25.004 297.054 25.108 301.428 ; 
        RECT 24.572 297.054 24.676 301.428 ; 
        RECT 24.14 297.054 24.244 301.428 ; 
        RECT 23.708 297.054 23.812 301.428 ; 
        RECT 22.856 297.054 23.164 301.428 ; 
        RECT 15.284 297.054 15.592 301.428 ; 
        RECT 14.636 297.054 14.74 301.428 ; 
        RECT 14.204 297.054 14.308 301.428 ; 
        RECT 13.772 297.054 13.876 301.428 ; 
        RECT 13.34 297.054 13.444 301.428 ; 
        RECT 12.908 297.054 13.012 301.428 ; 
        RECT 12.476 297.054 12.58 301.428 ; 
        RECT 12.044 297.054 12.148 301.428 ; 
        RECT 11.612 297.054 11.716 301.428 ; 
        RECT 11.18 297.054 11.284 301.428 ; 
        RECT 10.748 297.054 10.852 301.428 ; 
        RECT 10.316 297.054 10.42 301.428 ; 
        RECT 9.884 297.054 9.988 301.428 ; 
        RECT 9.452 297.054 9.556 301.428 ; 
        RECT 9.02 297.054 9.124 301.428 ; 
        RECT 8.588 297.054 8.692 301.428 ; 
        RECT 8.156 297.054 8.26 301.428 ; 
        RECT 7.724 297.054 7.828 301.428 ; 
        RECT 7.292 297.054 7.396 301.428 ; 
        RECT 6.86 297.054 6.964 301.428 ; 
        RECT 6.428 297.054 6.532 301.428 ; 
        RECT 5.996 297.054 6.1 301.428 ; 
        RECT 5.564 297.054 5.668 301.428 ; 
        RECT 5.132 297.054 5.236 301.428 ; 
        RECT 4.7 297.054 4.804 301.428 ; 
        RECT 4.268 297.054 4.372 301.428 ; 
        RECT 3.836 297.054 3.94 301.428 ; 
        RECT 3.404 297.054 3.508 301.428 ; 
        RECT 2.972 297.054 3.076 301.428 ; 
        RECT 2.54 297.054 2.644 301.428 ; 
        RECT 2.108 297.054 2.212 301.428 ; 
        RECT 1.676 297.054 1.78 301.428 ; 
        RECT 1.244 297.054 1.348 301.428 ; 
        RECT 0.812 297.054 0.916 301.428 ; 
        RECT 0 297.054 0.34 301.428 ; 
        RECT 20.72 301.374 21.232 305.748 ; 
        RECT 20.664 304.036 21.232 305.326 ; 
        RECT 20.072 302.944 20.32 305.748 ; 
        RECT 20.016 304.182 20.32 304.796 ; 
        RECT 20.072 301.374 20.176 305.748 ; 
        RECT 20.072 301.858 20.232 302.816 ; 
        RECT 20.072 301.374 20.32 301.73 ; 
        RECT 18.884 303.176 19.708 305.748 ; 
        RECT 19.604 301.374 19.708 305.748 ; 
        RECT 18.884 304.284 19.764 305.316 ; 
        RECT 18.884 301.374 19.276 305.748 ; 
        RECT 17.216 301.374 17.548 305.748 ; 
        RECT 17.216 301.728 17.604 305.47 ; 
        RECT 38.108 301.374 38.448 305.748 ; 
        RECT 37.532 301.374 37.636 305.748 ; 
        RECT 37.1 301.374 37.204 305.748 ; 
        RECT 36.668 301.374 36.772 305.748 ; 
        RECT 36.236 301.374 36.34 305.748 ; 
        RECT 35.804 301.374 35.908 305.748 ; 
        RECT 35.372 301.374 35.476 305.748 ; 
        RECT 34.94 301.374 35.044 305.748 ; 
        RECT 34.508 301.374 34.612 305.748 ; 
        RECT 34.076 301.374 34.18 305.748 ; 
        RECT 33.644 301.374 33.748 305.748 ; 
        RECT 33.212 301.374 33.316 305.748 ; 
        RECT 32.78 301.374 32.884 305.748 ; 
        RECT 32.348 301.374 32.452 305.748 ; 
        RECT 31.916 301.374 32.02 305.748 ; 
        RECT 31.484 301.374 31.588 305.748 ; 
        RECT 31.052 301.374 31.156 305.748 ; 
        RECT 30.62 301.374 30.724 305.748 ; 
        RECT 30.188 301.374 30.292 305.748 ; 
        RECT 29.756 301.374 29.86 305.748 ; 
        RECT 29.324 301.374 29.428 305.748 ; 
        RECT 28.892 301.374 28.996 305.748 ; 
        RECT 28.46 301.374 28.564 305.748 ; 
        RECT 28.028 301.374 28.132 305.748 ; 
        RECT 27.596 301.374 27.7 305.748 ; 
        RECT 27.164 301.374 27.268 305.748 ; 
        RECT 26.732 301.374 26.836 305.748 ; 
        RECT 26.3 301.374 26.404 305.748 ; 
        RECT 25.868 301.374 25.972 305.748 ; 
        RECT 25.436 301.374 25.54 305.748 ; 
        RECT 25.004 301.374 25.108 305.748 ; 
        RECT 24.572 301.374 24.676 305.748 ; 
        RECT 24.14 301.374 24.244 305.748 ; 
        RECT 23.708 301.374 23.812 305.748 ; 
        RECT 22.856 301.374 23.164 305.748 ; 
        RECT 15.284 301.374 15.592 305.748 ; 
        RECT 14.636 301.374 14.74 305.748 ; 
        RECT 14.204 301.374 14.308 305.748 ; 
        RECT 13.772 301.374 13.876 305.748 ; 
        RECT 13.34 301.374 13.444 305.748 ; 
        RECT 12.908 301.374 13.012 305.748 ; 
        RECT 12.476 301.374 12.58 305.748 ; 
        RECT 12.044 301.374 12.148 305.748 ; 
        RECT 11.612 301.374 11.716 305.748 ; 
        RECT 11.18 301.374 11.284 305.748 ; 
        RECT 10.748 301.374 10.852 305.748 ; 
        RECT 10.316 301.374 10.42 305.748 ; 
        RECT 9.884 301.374 9.988 305.748 ; 
        RECT 9.452 301.374 9.556 305.748 ; 
        RECT 9.02 301.374 9.124 305.748 ; 
        RECT 8.588 301.374 8.692 305.748 ; 
        RECT 8.156 301.374 8.26 305.748 ; 
        RECT 7.724 301.374 7.828 305.748 ; 
        RECT 7.292 301.374 7.396 305.748 ; 
        RECT 6.86 301.374 6.964 305.748 ; 
        RECT 6.428 301.374 6.532 305.748 ; 
        RECT 5.996 301.374 6.1 305.748 ; 
        RECT 5.564 301.374 5.668 305.748 ; 
        RECT 5.132 301.374 5.236 305.748 ; 
        RECT 4.7 301.374 4.804 305.748 ; 
        RECT 4.268 301.374 4.372 305.748 ; 
        RECT 3.836 301.374 3.94 305.748 ; 
        RECT 3.404 301.374 3.508 305.748 ; 
        RECT 2.972 301.374 3.076 305.748 ; 
        RECT 2.54 301.374 2.644 305.748 ; 
        RECT 2.108 301.374 2.212 305.748 ; 
        RECT 1.676 301.374 1.78 305.748 ; 
        RECT 1.244 301.374 1.348 305.748 ; 
        RECT 0.812 301.374 0.916 305.748 ; 
        RECT 0 301.374 0.34 305.748 ; 
        RECT 20.72 305.694 21.232 310.068 ; 
        RECT 20.664 308.356 21.232 309.646 ; 
        RECT 20.072 307.264 20.32 310.068 ; 
        RECT 20.016 308.502 20.32 309.116 ; 
        RECT 20.072 305.694 20.176 310.068 ; 
        RECT 20.072 306.178 20.232 307.136 ; 
        RECT 20.072 305.694 20.32 306.05 ; 
        RECT 18.884 307.496 19.708 310.068 ; 
        RECT 19.604 305.694 19.708 310.068 ; 
        RECT 18.884 308.604 19.764 309.636 ; 
        RECT 18.884 305.694 19.276 310.068 ; 
        RECT 17.216 305.694 17.548 310.068 ; 
        RECT 17.216 306.048 17.604 309.79 ; 
        RECT 38.108 305.694 38.448 310.068 ; 
        RECT 37.532 305.694 37.636 310.068 ; 
        RECT 37.1 305.694 37.204 310.068 ; 
        RECT 36.668 305.694 36.772 310.068 ; 
        RECT 36.236 305.694 36.34 310.068 ; 
        RECT 35.804 305.694 35.908 310.068 ; 
        RECT 35.372 305.694 35.476 310.068 ; 
        RECT 34.94 305.694 35.044 310.068 ; 
        RECT 34.508 305.694 34.612 310.068 ; 
        RECT 34.076 305.694 34.18 310.068 ; 
        RECT 33.644 305.694 33.748 310.068 ; 
        RECT 33.212 305.694 33.316 310.068 ; 
        RECT 32.78 305.694 32.884 310.068 ; 
        RECT 32.348 305.694 32.452 310.068 ; 
        RECT 31.916 305.694 32.02 310.068 ; 
        RECT 31.484 305.694 31.588 310.068 ; 
        RECT 31.052 305.694 31.156 310.068 ; 
        RECT 30.62 305.694 30.724 310.068 ; 
        RECT 30.188 305.694 30.292 310.068 ; 
        RECT 29.756 305.694 29.86 310.068 ; 
        RECT 29.324 305.694 29.428 310.068 ; 
        RECT 28.892 305.694 28.996 310.068 ; 
        RECT 28.46 305.694 28.564 310.068 ; 
        RECT 28.028 305.694 28.132 310.068 ; 
        RECT 27.596 305.694 27.7 310.068 ; 
        RECT 27.164 305.694 27.268 310.068 ; 
        RECT 26.732 305.694 26.836 310.068 ; 
        RECT 26.3 305.694 26.404 310.068 ; 
        RECT 25.868 305.694 25.972 310.068 ; 
        RECT 25.436 305.694 25.54 310.068 ; 
        RECT 25.004 305.694 25.108 310.068 ; 
        RECT 24.572 305.694 24.676 310.068 ; 
        RECT 24.14 305.694 24.244 310.068 ; 
        RECT 23.708 305.694 23.812 310.068 ; 
        RECT 22.856 305.694 23.164 310.068 ; 
        RECT 15.284 305.694 15.592 310.068 ; 
        RECT 14.636 305.694 14.74 310.068 ; 
        RECT 14.204 305.694 14.308 310.068 ; 
        RECT 13.772 305.694 13.876 310.068 ; 
        RECT 13.34 305.694 13.444 310.068 ; 
        RECT 12.908 305.694 13.012 310.068 ; 
        RECT 12.476 305.694 12.58 310.068 ; 
        RECT 12.044 305.694 12.148 310.068 ; 
        RECT 11.612 305.694 11.716 310.068 ; 
        RECT 11.18 305.694 11.284 310.068 ; 
        RECT 10.748 305.694 10.852 310.068 ; 
        RECT 10.316 305.694 10.42 310.068 ; 
        RECT 9.884 305.694 9.988 310.068 ; 
        RECT 9.452 305.694 9.556 310.068 ; 
        RECT 9.02 305.694 9.124 310.068 ; 
        RECT 8.588 305.694 8.692 310.068 ; 
        RECT 8.156 305.694 8.26 310.068 ; 
        RECT 7.724 305.694 7.828 310.068 ; 
        RECT 7.292 305.694 7.396 310.068 ; 
        RECT 6.86 305.694 6.964 310.068 ; 
        RECT 6.428 305.694 6.532 310.068 ; 
        RECT 5.996 305.694 6.1 310.068 ; 
        RECT 5.564 305.694 5.668 310.068 ; 
        RECT 5.132 305.694 5.236 310.068 ; 
        RECT 4.7 305.694 4.804 310.068 ; 
        RECT 4.268 305.694 4.372 310.068 ; 
        RECT 3.836 305.694 3.94 310.068 ; 
        RECT 3.404 305.694 3.508 310.068 ; 
        RECT 2.972 305.694 3.076 310.068 ; 
        RECT 2.54 305.694 2.644 310.068 ; 
        RECT 2.108 305.694 2.212 310.068 ; 
        RECT 1.676 305.694 1.78 310.068 ; 
        RECT 1.244 305.694 1.348 310.068 ; 
        RECT 0.812 305.694 0.916 310.068 ; 
        RECT 0 305.694 0.34 310.068 ; 
        RECT 20.72 310.014 21.232 314.388 ; 
        RECT 20.664 312.676 21.232 313.966 ; 
        RECT 20.072 311.584 20.32 314.388 ; 
        RECT 20.016 312.822 20.32 313.436 ; 
        RECT 20.072 310.014 20.176 314.388 ; 
        RECT 20.072 310.498 20.232 311.456 ; 
        RECT 20.072 310.014 20.32 310.37 ; 
        RECT 18.884 311.816 19.708 314.388 ; 
        RECT 19.604 310.014 19.708 314.388 ; 
        RECT 18.884 312.924 19.764 313.956 ; 
        RECT 18.884 310.014 19.276 314.388 ; 
        RECT 17.216 310.014 17.548 314.388 ; 
        RECT 17.216 310.368 17.604 314.11 ; 
        RECT 38.108 310.014 38.448 314.388 ; 
        RECT 37.532 310.014 37.636 314.388 ; 
        RECT 37.1 310.014 37.204 314.388 ; 
        RECT 36.668 310.014 36.772 314.388 ; 
        RECT 36.236 310.014 36.34 314.388 ; 
        RECT 35.804 310.014 35.908 314.388 ; 
        RECT 35.372 310.014 35.476 314.388 ; 
        RECT 34.94 310.014 35.044 314.388 ; 
        RECT 34.508 310.014 34.612 314.388 ; 
        RECT 34.076 310.014 34.18 314.388 ; 
        RECT 33.644 310.014 33.748 314.388 ; 
        RECT 33.212 310.014 33.316 314.388 ; 
        RECT 32.78 310.014 32.884 314.388 ; 
        RECT 32.348 310.014 32.452 314.388 ; 
        RECT 31.916 310.014 32.02 314.388 ; 
        RECT 31.484 310.014 31.588 314.388 ; 
        RECT 31.052 310.014 31.156 314.388 ; 
        RECT 30.62 310.014 30.724 314.388 ; 
        RECT 30.188 310.014 30.292 314.388 ; 
        RECT 29.756 310.014 29.86 314.388 ; 
        RECT 29.324 310.014 29.428 314.388 ; 
        RECT 28.892 310.014 28.996 314.388 ; 
        RECT 28.46 310.014 28.564 314.388 ; 
        RECT 28.028 310.014 28.132 314.388 ; 
        RECT 27.596 310.014 27.7 314.388 ; 
        RECT 27.164 310.014 27.268 314.388 ; 
        RECT 26.732 310.014 26.836 314.388 ; 
        RECT 26.3 310.014 26.404 314.388 ; 
        RECT 25.868 310.014 25.972 314.388 ; 
        RECT 25.436 310.014 25.54 314.388 ; 
        RECT 25.004 310.014 25.108 314.388 ; 
        RECT 24.572 310.014 24.676 314.388 ; 
        RECT 24.14 310.014 24.244 314.388 ; 
        RECT 23.708 310.014 23.812 314.388 ; 
        RECT 22.856 310.014 23.164 314.388 ; 
        RECT 15.284 310.014 15.592 314.388 ; 
        RECT 14.636 310.014 14.74 314.388 ; 
        RECT 14.204 310.014 14.308 314.388 ; 
        RECT 13.772 310.014 13.876 314.388 ; 
        RECT 13.34 310.014 13.444 314.388 ; 
        RECT 12.908 310.014 13.012 314.388 ; 
        RECT 12.476 310.014 12.58 314.388 ; 
        RECT 12.044 310.014 12.148 314.388 ; 
        RECT 11.612 310.014 11.716 314.388 ; 
        RECT 11.18 310.014 11.284 314.388 ; 
        RECT 10.748 310.014 10.852 314.388 ; 
        RECT 10.316 310.014 10.42 314.388 ; 
        RECT 9.884 310.014 9.988 314.388 ; 
        RECT 9.452 310.014 9.556 314.388 ; 
        RECT 9.02 310.014 9.124 314.388 ; 
        RECT 8.588 310.014 8.692 314.388 ; 
        RECT 8.156 310.014 8.26 314.388 ; 
        RECT 7.724 310.014 7.828 314.388 ; 
        RECT 7.292 310.014 7.396 314.388 ; 
        RECT 6.86 310.014 6.964 314.388 ; 
        RECT 6.428 310.014 6.532 314.388 ; 
        RECT 5.996 310.014 6.1 314.388 ; 
        RECT 5.564 310.014 5.668 314.388 ; 
        RECT 5.132 310.014 5.236 314.388 ; 
        RECT 4.7 310.014 4.804 314.388 ; 
        RECT 4.268 310.014 4.372 314.388 ; 
        RECT 3.836 310.014 3.94 314.388 ; 
        RECT 3.404 310.014 3.508 314.388 ; 
        RECT 2.972 310.014 3.076 314.388 ; 
        RECT 2.54 310.014 2.644 314.388 ; 
        RECT 2.108 310.014 2.212 314.388 ; 
        RECT 1.676 310.014 1.78 314.388 ; 
        RECT 1.244 310.014 1.348 314.388 ; 
        RECT 0.812 310.014 0.916 314.388 ; 
        RECT 0 310.014 0.34 314.388 ; 
        RECT 20.72 314.334 21.232 318.708 ; 
        RECT 20.664 316.996 21.232 318.286 ; 
        RECT 20.072 315.904 20.32 318.708 ; 
        RECT 20.016 317.142 20.32 317.756 ; 
        RECT 20.072 314.334 20.176 318.708 ; 
        RECT 20.072 314.818 20.232 315.776 ; 
        RECT 20.072 314.334 20.32 314.69 ; 
        RECT 18.884 316.136 19.708 318.708 ; 
        RECT 19.604 314.334 19.708 318.708 ; 
        RECT 18.884 317.244 19.764 318.276 ; 
        RECT 18.884 314.334 19.276 318.708 ; 
        RECT 17.216 314.334 17.548 318.708 ; 
        RECT 17.216 314.688 17.604 318.43 ; 
        RECT 38.108 314.334 38.448 318.708 ; 
        RECT 37.532 314.334 37.636 318.708 ; 
        RECT 37.1 314.334 37.204 318.708 ; 
        RECT 36.668 314.334 36.772 318.708 ; 
        RECT 36.236 314.334 36.34 318.708 ; 
        RECT 35.804 314.334 35.908 318.708 ; 
        RECT 35.372 314.334 35.476 318.708 ; 
        RECT 34.94 314.334 35.044 318.708 ; 
        RECT 34.508 314.334 34.612 318.708 ; 
        RECT 34.076 314.334 34.18 318.708 ; 
        RECT 33.644 314.334 33.748 318.708 ; 
        RECT 33.212 314.334 33.316 318.708 ; 
        RECT 32.78 314.334 32.884 318.708 ; 
        RECT 32.348 314.334 32.452 318.708 ; 
        RECT 31.916 314.334 32.02 318.708 ; 
        RECT 31.484 314.334 31.588 318.708 ; 
        RECT 31.052 314.334 31.156 318.708 ; 
        RECT 30.62 314.334 30.724 318.708 ; 
        RECT 30.188 314.334 30.292 318.708 ; 
        RECT 29.756 314.334 29.86 318.708 ; 
        RECT 29.324 314.334 29.428 318.708 ; 
        RECT 28.892 314.334 28.996 318.708 ; 
        RECT 28.46 314.334 28.564 318.708 ; 
        RECT 28.028 314.334 28.132 318.708 ; 
        RECT 27.596 314.334 27.7 318.708 ; 
        RECT 27.164 314.334 27.268 318.708 ; 
        RECT 26.732 314.334 26.836 318.708 ; 
        RECT 26.3 314.334 26.404 318.708 ; 
        RECT 25.868 314.334 25.972 318.708 ; 
        RECT 25.436 314.334 25.54 318.708 ; 
        RECT 25.004 314.334 25.108 318.708 ; 
        RECT 24.572 314.334 24.676 318.708 ; 
        RECT 24.14 314.334 24.244 318.708 ; 
        RECT 23.708 314.334 23.812 318.708 ; 
        RECT 22.856 314.334 23.164 318.708 ; 
        RECT 15.284 314.334 15.592 318.708 ; 
        RECT 14.636 314.334 14.74 318.708 ; 
        RECT 14.204 314.334 14.308 318.708 ; 
        RECT 13.772 314.334 13.876 318.708 ; 
        RECT 13.34 314.334 13.444 318.708 ; 
        RECT 12.908 314.334 13.012 318.708 ; 
        RECT 12.476 314.334 12.58 318.708 ; 
        RECT 12.044 314.334 12.148 318.708 ; 
        RECT 11.612 314.334 11.716 318.708 ; 
        RECT 11.18 314.334 11.284 318.708 ; 
        RECT 10.748 314.334 10.852 318.708 ; 
        RECT 10.316 314.334 10.42 318.708 ; 
        RECT 9.884 314.334 9.988 318.708 ; 
        RECT 9.452 314.334 9.556 318.708 ; 
        RECT 9.02 314.334 9.124 318.708 ; 
        RECT 8.588 314.334 8.692 318.708 ; 
        RECT 8.156 314.334 8.26 318.708 ; 
        RECT 7.724 314.334 7.828 318.708 ; 
        RECT 7.292 314.334 7.396 318.708 ; 
        RECT 6.86 314.334 6.964 318.708 ; 
        RECT 6.428 314.334 6.532 318.708 ; 
        RECT 5.996 314.334 6.1 318.708 ; 
        RECT 5.564 314.334 5.668 318.708 ; 
        RECT 5.132 314.334 5.236 318.708 ; 
        RECT 4.7 314.334 4.804 318.708 ; 
        RECT 4.268 314.334 4.372 318.708 ; 
        RECT 3.836 314.334 3.94 318.708 ; 
        RECT 3.404 314.334 3.508 318.708 ; 
        RECT 2.972 314.334 3.076 318.708 ; 
        RECT 2.54 314.334 2.644 318.708 ; 
        RECT 2.108 314.334 2.212 318.708 ; 
        RECT 1.676 314.334 1.78 318.708 ; 
        RECT 1.244 314.334 1.348 318.708 ; 
        RECT 0.812 314.334 0.916 318.708 ; 
        RECT 0 314.334 0.34 318.708 ; 
        RECT 20.72 318.654 21.232 323.028 ; 
        RECT 20.664 321.316 21.232 322.606 ; 
        RECT 20.072 320.224 20.32 323.028 ; 
        RECT 20.016 321.462 20.32 322.076 ; 
        RECT 20.072 318.654 20.176 323.028 ; 
        RECT 20.072 319.138 20.232 320.096 ; 
        RECT 20.072 318.654 20.32 319.01 ; 
        RECT 18.884 320.456 19.708 323.028 ; 
        RECT 19.604 318.654 19.708 323.028 ; 
        RECT 18.884 321.564 19.764 322.596 ; 
        RECT 18.884 318.654 19.276 323.028 ; 
        RECT 17.216 318.654 17.548 323.028 ; 
        RECT 17.216 319.008 17.604 322.75 ; 
        RECT 38.108 318.654 38.448 323.028 ; 
        RECT 37.532 318.654 37.636 323.028 ; 
        RECT 37.1 318.654 37.204 323.028 ; 
        RECT 36.668 318.654 36.772 323.028 ; 
        RECT 36.236 318.654 36.34 323.028 ; 
        RECT 35.804 318.654 35.908 323.028 ; 
        RECT 35.372 318.654 35.476 323.028 ; 
        RECT 34.94 318.654 35.044 323.028 ; 
        RECT 34.508 318.654 34.612 323.028 ; 
        RECT 34.076 318.654 34.18 323.028 ; 
        RECT 33.644 318.654 33.748 323.028 ; 
        RECT 33.212 318.654 33.316 323.028 ; 
        RECT 32.78 318.654 32.884 323.028 ; 
        RECT 32.348 318.654 32.452 323.028 ; 
        RECT 31.916 318.654 32.02 323.028 ; 
        RECT 31.484 318.654 31.588 323.028 ; 
        RECT 31.052 318.654 31.156 323.028 ; 
        RECT 30.62 318.654 30.724 323.028 ; 
        RECT 30.188 318.654 30.292 323.028 ; 
        RECT 29.756 318.654 29.86 323.028 ; 
        RECT 29.324 318.654 29.428 323.028 ; 
        RECT 28.892 318.654 28.996 323.028 ; 
        RECT 28.46 318.654 28.564 323.028 ; 
        RECT 28.028 318.654 28.132 323.028 ; 
        RECT 27.596 318.654 27.7 323.028 ; 
        RECT 27.164 318.654 27.268 323.028 ; 
        RECT 26.732 318.654 26.836 323.028 ; 
        RECT 26.3 318.654 26.404 323.028 ; 
        RECT 25.868 318.654 25.972 323.028 ; 
        RECT 25.436 318.654 25.54 323.028 ; 
        RECT 25.004 318.654 25.108 323.028 ; 
        RECT 24.572 318.654 24.676 323.028 ; 
        RECT 24.14 318.654 24.244 323.028 ; 
        RECT 23.708 318.654 23.812 323.028 ; 
        RECT 22.856 318.654 23.164 323.028 ; 
        RECT 15.284 318.654 15.592 323.028 ; 
        RECT 14.636 318.654 14.74 323.028 ; 
        RECT 14.204 318.654 14.308 323.028 ; 
        RECT 13.772 318.654 13.876 323.028 ; 
        RECT 13.34 318.654 13.444 323.028 ; 
        RECT 12.908 318.654 13.012 323.028 ; 
        RECT 12.476 318.654 12.58 323.028 ; 
        RECT 12.044 318.654 12.148 323.028 ; 
        RECT 11.612 318.654 11.716 323.028 ; 
        RECT 11.18 318.654 11.284 323.028 ; 
        RECT 10.748 318.654 10.852 323.028 ; 
        RECT 10.316 318.654 10.42 323.028 ; 
        RECT 9.884 318.654 9.988 323.028 ; 
        RECT 9.452 318.654 9.556 323.028 ; 
        RECT 9.02 318.654 9.124 323.028 ; 
        RECT 8.588 318.654 8.692 323.028 ; 
        RECT 8.156 318.654 8.26 323.028 ; 
        RECT 7.724 318.654 7.828 323.028 ; 
        RECT 7.292 318.654 7.396 323.028 ; 
        RECT 6.86 318.654 6.964 323.028 ; 
        RECT 6.428 318.654 6.532 323.028 ; 
        RECT 5.996 318.654 6.1 323.028 ; 
        RECT 5.564 318.654 5.668 323.028 ; 
        RECT 5.132 318.654 5.236 323.028 ; 
        RECT 4.7 318.654 4.804 323.028 ; 
        RECT 4.268 318.654 4.372 323.028 ; 
        RECT 3.836 318.654 3.94 323.028 ; 
        RECT 3.404 318.654 3.508 323.028 ; 
        RECT 2.972 318.654 3.076 323.028 ; 
        RECT 2.54 318.654 2.644 323.028 ; 
        RECT 2.108 318.654 2.212 323.028 ; 
        RECT 1.676 318.654 1.78 323.028 ; 
        RECT 1.244 318.654 1.348 323.028 ; 
        RECT 0.812 318.654 0.916 323.028 ; 
        RECT 0 318.654 0.34 323.028 ; 
        RECT 20.72 322.974 21.232 327.348 ; 
        RECT 20.664 325.636 21.232 326.926 ; 
        RECT 20.072 324.544 20.32 327.348 ; 
        RECT 20.016 325.782 20.32 326.396 ; 
        RECT 20.072 322.974 20.176 327.348 ; 
        RECT 20.072 323.458 20.232 324.416 ; 
        RECT 20.072 322.974 20.32 323.33 ; 
        RECT 18.884 324.776 19.708 327.348 ; 
        RECT 19.604 322.974 19.708 327.348 ; 
        RECT 18.884 325.884 19.764 326.916 ; 
        RECT 18.884 322.974 19.276 327.348 ; 
        RECT 17.216 322.974 17.548 327.348 ; 
        RECT 17.216 323.328 17.604 327.07 ; 
        RECT 38.108 322.974 38.448 327.348 ; 
        RECT 37.532 322.974 37.636 327.348 ; 
        RECT 37.1 322.974 37.204 327.348 ; 
        RECT 36.668 322.974 36.772 327.348 ; 
        RECT 36.236 322.974 36.34 327.348 ; 
        RECT 35.804 322.974 35.908 327.348 ; 
        RECT 35.372 322.974 35.476 327.348 ; 
        RECT 34.94 322.974 35.044 327.348 ; 
        RECT 34.508 322.974 34.612 327.348 ; 
        RECT 34.076 322.974 34.18 327.348 ; 
        RECT 33.644 322.974 33.748 327.348 ; 
        RECT 33.212 322.974 33.316 327.348 ; 
        RECT 32.78 322.974 32.884 327.348 ; 
        RECT 32.348 322.974 32.452 327.348 ; 
        RECT 31.916 322.974 32.02 327.348 ; 
        RECT 31.484 322.974 31.588 327.348 ; 
        RECT 31.052 322.974 31.156 327.348 ; 
        RECT 30.62 322.974 30.724 327.348 ; 
        RECT 30.188 322.974 30.292 327.348 ; 
        RECT 29.756 322.974 29.86 327.348 ; 
        RECT 29.324 322.974 29.428 327.348 ; 
        RECT 28.892 322.974 28.996 327.348 ; 
        RECT 28.46 322.974 28.564 327.348 ; 
        RECT 28.028 322.974 28.132 327.348 ; 
        RECT 27.596 322.974 27.7 327.348 ; 
        RECT 27.164 322.974 27.268 327.348 ; 
        RECT 26.732 322.974 26.836 327.348 ; 
        RECT 26.3 322.974 26.404 327.348 ; 
        RECT 25.868 322.974 25.972 327.348 ; 
        RECT 25.436 322.974 25.54 327.348 ; 
        RECT 25.004 322.974 25.108 327.348 ; 
        RECT 24.572 322.974 24.676 327.348 ; 
        RECT 24.14 322.974 24.244 327.348 ; 
        RECT 23.708 322.974 23.812 327.348 ; 
        RECT 22.856 322.974 23.164 327.348 ; 
        RECT 15.284 322.974 15.592 327.348 ; 
        RECT 14.636 322.974 14.74 327.348 ; 
        RECT 14.204 322.974 14.308 327.348 ; 
        RECT 13.772 322.974 13.876 327.348 ; 
        RECT 13.34 322.974 13.444 327.348 ; 
        RECT 12.908 322.974 13.012 327.348 ; 
        RECT 12.476 322.974 12.58 327.348 ; 
        RECT 12.044 322.974 12.148 327.348 ; 
        RECT 11.612 322.974 11.716 327.348 ; 
        RECT 11.18 322.974 11.284 327.348 ; 
        RECT 10.748 322.974 10.852 327.348 ; 
        RECT 10.316 322.974 10.42 327.348 ; 
        RECT 9.884 322.974 9.988 327.348 ; 
        RECT 9.452 322.974 9.556 327.348 ; 
        RECT 9.02 322.974 9.124 327.348 ; 
        RECT 8.588 322.974 8.692 327.348 ; 
        RECT 8.156 322.974 8.26 327.348 ; 
        RECT 7.724 322.974 7.828 327.348 ; 
        RECT 7.292 322.974 7.396 327.348 ; 
        RECT 6.86 322.974 6.964 327.348 ; 
        RECT 6.428 322.974 6.532 327.348 ; 
        RECT 5.996 322.974 6.1 327.348 ; 
        RECT 5.564 322.974 5.668 327.348 ; 
        RECT 5.132 322.974 5.236 327.348 ; 
        RECT 4.7 322.974 4.804 327.348 ; 
        RECT 4.268 322.974 4.372 327.348 ; 
        RECT 3.836 322.974 3.94 327.348 ; 
        RECT 3.404 322.974 3.508 327.348 ; 
        RECT 2.972 322.974 3.076 327.348 ; 
        RECT 2.54 322.974 2.644 327.348 ; 
        RECT 2.108 322.974 2.212 327.348 ; 
        RECT 1.676 322.974 1.78 327.348 ; 
        RECT 1.244 322.974 1.348 327.348 ; 
        RECT 0.812 322.974 0.916 327.348 ; 
        RECT 0 322.974 0.34 327.348 ; 
        RECT 20.72 327.294 21.232 331.668 ; 
        RECT 20.664 329.956 21.232 331.246 ; 
        RECT 20.072 328.864 20.32 331.668 ; 
        RECT 20.016 330.102 20.32 330.716 ; 
        RECT 20.072 327.294 20.176 331.668 ; 
        RECT 20.072 327.778 20.232 328.736 ; 
        RECT 20.072 327.294 20.32 327.65 ; 
        RECT 18.884 329.096 19.708 331.668 ; 
        RECT 19.604 327.294 19.708 331.668 ; 
        RECT 18.884 330.204 19.764 331.236 ; 
        RECT 18.884 327.294 19.276 331.668 ; 
        RECT 17.216 327.294 17.548 331.668 ; 
        RECT 17.216 327.648 17.604 331.39 ; 
        RECT 38.108 327.294 38.448 331.668 ; 
        RECT 37.532 327.294 37.636 331.668 ; 
        RECT 37.1 327.294 37.204 331.668 ; 
        RECT 36.668 327.294 36.772 331.668 ; 
        RECT 36.236 327.294 36.34 331.668 ; 
        RECT 35.804 327.294 35.908 331.668 ; 
        RECT 35.372 327.294 35.476 331.668 ; 
        RECT 34.94 327.294 35.044 331.668 ; 
        RECT 34.508 327.294 34.612 331.668 ; 
        RECT 34.076 327.294 34.18 331.668 ; 
        RECT 33.644 327.294 33.748 331.668 ; 
        RECT 33.212 327.294 33.316 331.668 ; 
        RECT 32.78 327.294 32.884 331.668 ; 
        RECT 32.348 327.294 32.452 331.668 ; 
        RECT 31.916 327.294 32.02 331.668 ; 
        RECT 31.484 327.294 31.588 331.668 ; 
        RECT 31.052 327.294 31.156 331.668 ; 
        RECT 30.62 327.294 30.724 331.668 ; 
        RECT 30.188 327.294 30.292 331.668 ; 
        RECT 29.756 327.294 29.86 331.668 ; 
        RECT 29.324 327.294 29.428 331.668 ; 
        RECT 28.892 327.294 28.996 331.668 ; 
        RECT 28.46 327.294 28.564 331.668 ; 
        RECT 28.028 327.294 28.132 331.668 ; 
        RECT 27.596 327.294 27.7 331.668 ; 
        RECT 27.164 327.294 27.268 331.668 ; 
        RECT 26.732 327.294 26.836 331.668 ; 
        RECT 26.3 327.294 26.404 331.668 ; 
        RECT 25.868 327.294 25.972 331.668 ; 
        RECT 25.436 327.294 25.54 331.668 ; 
        RECT 25.004 327.294 25.108 331.668 ; 
        RECT 24.572 327.294 24.676 331.668 ; 
        RECT 24.14 327.294 24.244 331.668 ; 
        RECT 23.708 327.294 23.812 331.668 ; 
        RECT 22.856 327.294 23.164 331.668 ; 
        RECT 15.284 327.294 15.592 331.668 ; 
        RECT 14.636 327.294 14.74 331.668 ; 
        RECT 14.204 327.294 14.308 331.668 ; 
        RECT 13.772 327.294 13.876 331.668 ; 
        RECT 13.34 327.294 13.444 331.668 ; 
        RECT 12.908 327.294 13.012 331.668 ; 
        RECT 12.476 327.294 12.58 331.668 ; 
        RECT 12.044 327.294 12.148 331.668 ; 
        RECT 11.612 327.294 11.716 331.668 ; 
        RECT 11.18 327.294 11.284 331.668 ; 
        RECT 10.748 327.294 10.852 331.668 ; 
        RECT 10.316 327.294 10.42 331.668 ; 
        RECT 9.884 327.294 9.988 331.668 ; 
        RECT 9.452 327.294 9.556 331.668 ; 
        RECT 9.02 327.294 9.124 331.668 ; 
        RECT 8.588 327.294 8.692 331.668 ; 
        RECT 8.156 327.294 8.26 331.668 ; 
        RECT 7.724 327.294 7.828 331.668 ; 
        RECT 7.292 327.294 7.396 331.668 ; 
        RECT 6.86 327.294 6.964 331.668 ; 
        RECT 6.428 327.294 6.532 331.668 ; 
        RECT 5.996 327.294 6.1 331.668 ; 
        RECT 5.564 327.294 5.668 331.668 ; 
        RECT 5.132 327.294 5.236 331.668 ; 
        RECT 4.7 327.294 4.804 331.668 ; 
        RECT 4.268 327.294 4.372 331.668 ; 
        RECT 3.836 327.294 3.94 331.668 ; 
        RECT 3.404 327.294 3.508 331.668 ; 
        RECT 2.972 327.294 3.076 331.668 ; 
        RECT 2.54 327.294 2.644 331.668 ; 
        RECT 2.108 327.294 2.212 331.668 ; 
        RECT 1.676 327.294 1.78 331.668 ; 
        RECT 1.244 327.294 1.348 331.668 ; 
        RECT 0.812 327.294 0.916 331.668 ; 
        RECT 0 327.294 0.34 331.668 ; 
        RECT 20.72 331.614 21.232 335.988 ; 
        RECT 20.664 334.276 21.232 335.566 ; 
        RECT 20.072 333.184 20.32 335.988 ; 
        RECT 20.016 334.422 20.32 335.036 ; 
        RECT 20.072 331.614 20.176 335.988 ; 
        RECT 20.072 332.098 20.232 333.056 ; 
        RECT 20.072 331.614 20.32 331.97 ; 
        RECT 18.884 333.416 19.708 335.988 ; 
        RECT 19.604 331.614 19.708 335.988 ; 
        RECT 18.884 334.524 19.764 335.556 ; 
        RECT 18.884 331.614 19.276 335.988 ; 
        RECT 17.216 331.614 17.548 335.988 ; 
        RECT 17.216 331.968 17.604 335.71 ; 
        RECT 38.108 331.614 38.448 335.988 ; 
        RECT 37.532 331.614 37.636 335.988 ; 
        RECT 37.1 331.614 37.204 335.988 ; 
        RECT 36.668 331.614 36.772 335.988 ; 
        RECT 36.236 331.614 36.34 335.988 ; 
        RECT 35.804 331.614 35.908 335.988 ; 
        RECT 35.372 331.614 35.476 335.988 ; 
        RECT 34.94 331.614 35.044 335.988 ; 
        RECT 34.508 331.614 34.612 335.988 ; 
        RECT 34.076 331.614 34.18 335.988 ; 
        RECT 33.644 331.614 33.748 335.988 ; 
        RECT 33.212 331.614 33.316 335.988 ; 
        RECT 32.78 331.614 32.884 335.988 ; 
        RECT 32.348 331.614 32.452 335.988 ; 
        RECT 31.916 331.614 32.02 335.988 ; 
        RECT 31.484 331.614 31.588 335.988 ; 
        RECT 31.052 331.614 31.156 335.988 ; 
        RECT 30.62 331.614 30.724 335.988 ; 
        RECT 30.188 331.614 30.292 335.988 ; 
        RECT 29.756 331.614 29.86 335.988 ; 
        RECT 29.324 331.614 29.428 335.988 ; 
        RECT 28.892 331.614 28.996 335.988 ; 
        RECT 28.46 331.614 28.564 335.988 ; 
        RECT 28.028 331.614 28.132 335.988 ; 
        RECT 27.596 331.614 27.7 335.988 ; 
        RECT 27.164 331.614 27.268 335.988 ; 
        RECT 26.732 331.614 26.836 335.988 ; 
        RECT 26.3 331.614 26.404 335.988 ; 
        RECT 25.868 331.614 25.972 335.988 ; 
        RECT 25.436 331.614 25.54 335.988 ; 
        RECT 25.004 331.614 25.108 335.988 ; 
        RECT 24.572 331.614 24.676 335.988 ; 
        RECT 24.14 331.614 24.244 335.988 ; 
        RECT 23.708 331.614 23.812 335.988 ; 
        RECT 22.856 331.614 23.164 335.988 ; 
        RECT 15.284 331.614 15.592 335.988 ; 
        RECT 14.636 331.614 14.74 335.988 ; 
        RECT 14.204 331.614 14.308 335.988 ; 
        RECT 13.772 331.614 13.876 335.988 ; 
        RECT 13.34 331.614 13.444 335.988 ; 
        RECT 12.908 331.614 13.012 335.988 ; 
        RECT 12.476 331.614 12.58 335.988 ; 
        RECT 12.044 331.614 12.148 335.988 ; 
        RECT 11.612 331.614 11.716 335.988 ; 
        RECT 11.18 331.614 11.284 335.988 ; 
        RECT 10.748 331.614 10.852 335.988 ; 
        RECT 10.316 331.614 10.42 335.988 ; 
        RECT 9.884 331.614 9.988 335.988 ; 
        RECT 9.452 331.614 9.556 335.988 ; 
        RECT 9.02 331.614 9.124 335.988 ; 
        RECT 8.588 331.614 8.692 335.988 ; 
        RECT 8.156 331.614 8.26 335.988 ; 
        RECT 7.724 331.614 7.828 335.988 ; 
        RECT 7.292 331.614 7.396 335.988 ; 
        RECT 6.86 331.614 6.964 335.988 ; 
        RECT 6.428 331.614 6.532 335.988 ; 
        RECT 5.996 331.614 6.1 335.988 ; 
        RECT 5.564 331.614 5.668 335.988 ; 
        RECT 5.132 331.614 5.236 335.988 ; 
        RECT 4.7 331.614 4.804 335.988 ; 
        RECT 4.268 331.614 4.372 335.988 ; 
        RECT 3.836 331.614 3.94 335.988 ; 
        RECT 3.404 331.614 3.508 335.988 ; 
        RECT 2.972 331.614 3.076 335.988 ; 
        RECT 2.54 331.614 2.644 335.988 ; 
        RECT 2.108 331.614 2.212 335.988 ; 
        RECT 1.676 331.614 1.78 335.988 ; 
        RECT 1.244 331.614 1.348 335.988 ; 
        RECT 0.812 331.614 0.916 335.988 ; 
        RECT 0 331.614 0.34 335.988 ; 
        RECT 20.72 335.934 21.232 340.308 ; 
        RECT 20.664 338.596 21.232 339.886 ; 
        RECT 20.072 337.504 20.32 340.308 ; 
        RECT 20.016 338.742 20.32 339.356 ; 
        RECT 20.072 335.934 20.176 340.308 ; 
        RECT 20.072 336.418 20.232 337.376 ; 
        RECT 20.072 335.934 20.32 336.29 ; 
        RECT 18.884 337.736 19.708 340.308 ; 
        RECT 19.604 335.934 19.708 340.308 ; 
        RECT 18.884 338.844 19.764 339.876 ; 
        RECT 18.884 335.934 19.276 340.308 ; 
        RECT 17.216 335.934 17.548 340.308 ; 
        RECT 17.216 336.288 17.604 340.03 ; 
        RECT 38.108 335.934 38.448 340.308 ; 
        RECT 37.532 335.934 37.636 340.308 ; 
        RECT 37.1 335.934 37.204 340.308 ; 
        RECT 36.668 335.934 36.772 340.308 ; 
        RECT 36.236 335.934 36.34 340.308 ; 
        RECT 35.804 335.934 35.908 340.308 ; 
        RECT 35.372 335.934 35.476 340.308 ; 
        RECT 34.94 335.934 35.044 340.308 ; 
        RECT 34.508 335.934 34.612 340.308 ; 
        RECT 34.076 335.934 34.18 340.308 ; 
        RECT 33.644 335.934 33.748 340.308 ; 
        RECT 33.212 335.934 33.316 340.308 ; 
        RECT 32.78 335.934 32.884 340.308 ; 
        RECT 32.348 335.934 32.452 340.308 ; 
        RECT 31.916 335.934 32.02 340.308 ; 
        RECT 31.484 335.934 31.588 340.308 ; 
        RECT 31.052 335.934 31.156 340.308 ; 
        RECT 30.62 335.934 30.724 340.308 ; 
        RECT 30.188 335.934 30.292 340.308 ; 
        RECT 29.756 335.934 29.86 340.308 ; 
        RECT 29.324 335.934 29.428 340.308 ; 
        RECT 28.892 335.934 28.996 340.308 ; 
        RECT 28.46 335.934 28.564 340.308 ; 
        RECT 28.028 335.934 28.132 340.308 ; 
        RECT 27.596 335.934 27.7 340.308 ; 
        RECT 27.164 335.934 27.268 340.308 ; 
        RECT 26.732 335.934 26.836 340.308 ; 
        RECT 26.3 335.934 26.404 340.308 ; 
        RECT 25.868 335.934 25.972 340.308 ; 
        RECT 25.436 335.934 25.54 340.308 ; 
        RECT 25.004 335.934 25.108 340.308 ; 
        RECT 24.572 335.934 24.676 340.308 ; 
        RECT 24.14 335.934 24.244 340.308 ; 
        RECT 23.708 335.934 23.812 340.308 ; 
        RECT 22.856 335.934 23.164 340.308 ; 
        RECT 15.284 335.934 15.592 340.308 ; 
        RECT 14.636 335.934 14.74 340.308 ; 
        RECT 14.204 335.934 14.308 340.308 ; 
        RECT 13.772 335.934 13.876 340.308 ; 
        RECT 13.34 335.934 13.444 340.308 ; 
        RECT 12.908 335.934 13.012 340.308 ; 
        RECT 12.476 335.934 12.58 340.308 ; 
        RECT 12.044 335.934 12.148 340.308 ; 
        RECT 11.612 335.934 11.716 340.308 ; 
        RECT 11.18 335.934 11.284 340.308 ; 
        RECT 10.748 335.934 10.852 340.308 ; 
        RECT 10.316 335.934 10.42 340.308 ; 
        RECT 9.884 335.934 9.988 340.308 ; 
        RECT 9.452 335.934 9.556 340.308 ; 
        RECT 9.02 335.934 9.124 340.308 ; 
        RECT 8.588 335.934 8.692 340.308 ; 
        RECT 8.156 335.934 8.26 340.308 ; 
        RECT 7.724 335.934 7.828 340.308 ; 
        RECT 7.292 335.934 7.396 340.308 ; 
        RECT 6.86 335.934 6.964 340.308 ; 
        RECT 6.428 335.934 6.532 340.308 ; 
        RECT 5.996 335.934 6.1 340.308 ; 
        RECT 5.564 335.934 5.668 340.308 ; 
        RECT 5.132 335.934 5.236 340.308 ; 
        RECT 4.7 335.934 4.804 340.308 ; 
        RECT 4.268 335.934 4.372 340.308 ; 
        RECT 3.836 335.934 3.94 340.308 ; 
        RECT 3.404 335.934 3.508 340.308 ; 
        RECT 2.972 335.934 3.076 340.308 ; 
        RECT 2.54 335.934 2.644 340.308 ; 
        RECT 2.108 335.934 2.212 340.308 ; 
        RECT 1.676 335.934 1.78 340.308 ; 
        RECT 1.244 335.934 1.348 340.308 ; 
        RECT 0.812 335.934 0.916 340.308 ; 
        RECT 0 335.934 0.34 340.308 ; 
        RECT 20.72 340.254 21.232 344.628 ; 
        RECT 20.664 342.916 21.232 344.206 ; 
        RECT 20.072 341.824 20.32 344.628 ; 
        RECT 20.016 343.062 20.32 343.676 ; 
        RECT 20.072 340.254 20.176 344.628 ; 
        RECT 20.072 340.738 20.232 341.696 ; 
        RECT 20.072 340.254 20.32 340.61 ; 
        RECT 18.884 342.056 19.708 344.628 ; 
        RECT 19.604 340.254 19.708 344.628 ; 
        RECT 18.884 343.164 19.764 344.196 ; 
        RECT 18.884 340.254 19.276 344.628 ; 
        RECT 17.216 340.254 17.548 344.628 ; 
        RECT 17.216 340.608 17.604 344.35 ; 
        RECT 38.108 340.254 38.448 344.628 ; 
        RECT 37.532 340.254 37.636 344.628 ; 
        RECT 37.1 340.254 37.204 344.628 ; 
        RECT 36.668 340.254 36.772 344.628 ; 
        RECT 36.236 340.254 36.34 344.628 ; 
        RECT 35.804 340.254 35.908 344.628 ; 
        RECT 35.372 340.254 35.476 344.628 ; 
        RECT 34.94 340.254 35.044 344.628 ; 
        RECT 34.508 340.254 34.612 344.628 ; 
        RECT 34.076 340.254 34.18 344.628 ; 
        RECT 33.644 340.254 33.748 344.628 ; 
        RECT 33.212 340.254 33.316 344.628 ; 
        RECT 32.78 340.254 32.884 344.628 ; 
        RECT 32.348 340.254 32.452 344.628 ; 
        RECT 31.916 340.254 32.02 344.628 ; 
        RECT 31.484 340.254 31.588 344.628 ; 
        RECT 31.052 340.254 31.156 344.628 ; 
        RECT 30.62 340.254 30.724 344.628 ; 
        RECT 30.188 340.254 30.292 344.628 ; 
        RECT 29.756 340.254 29.86 344.628 ; 
        RECT 29.324 340.254 29.428 344.628 ; 
        RECT 28.892 340.254 28.996 344.628 ; 
        RECT 28.46 340.254 28.564 344.628 ; 
        RECT 28.028 340.254 28.132 344.628 ; 
        RECT 27.596 340.254 27.7 344.628 ; 
        RECT 27.164 340.254 27.268 344.628 ; 
        RECT 26.732 340.254 26.836 344.628 ; 
        RECT 26.3 340.254 26.404 344.628 ; 
        RECT 25.868 340.254 25.972 344.628 ; 
        RECT 25.436 340.254 25.54 344.628 ; 
        RECT 25.004 340.254 25.108 344.628 ; 
        RECT 24.572 340.254 24.676 344.628 ; 
        RECT 24.14 340.254 24.244 344.628 ; 
        RECT 23.708 340.254 23.812 344.628 ; 
        RECT 22.856 340.254 23.164 344.628 ; 
        RECT 15.284 340.254 15.592 344.628 ; 
        RECT 14.636 340.254 14.74 344.628 ; 
        RECT 14.204 340.254 14.308 344.628 ; 
        RECT 13.772 340.254 13.876 344.628 ; 
        RECT 13.34 340.254 13.444 344.628 ; 
        RECT 12.908 340.254 13.012 344.628 ; 
        RECT 12.476 340.254 12.58 344.628 ; 
        RECT 12.044 340.254 12.148 344.628 ; 
        RECT 11.612 340.254 11.716 344.628 ; 
        RECT 11.18 340.254 11.284 344.628 ; 
        RECT 10.748 340.254 10.852 344.628 ; 
        RECT 10.316 340.254 10.42 344.628 ; 
        RECT 9.884 340.254 9.988 344.628 ; 
        RECT 9.452 340.254 9.556 344.628 ; 
        RECT 9.02 340.254 9.124 344.628 ; 
        RECT 8.588 340.254 8.692 344.628 ; 
        RECT 8.156 340.254 8.26 344.628 ; 
        RECT 7.724 340.254 7.828 344.628 ; 
        RECT 7.292 340.254 7.396 344.628 ; 
        RECT 6.86 340.254 6.964 344.628 ; 
        RECT 6.428 340.254 6.532 344.628 ; 
        RECT 5.996 340.254 6.1 344.628 ; 
        RECT 5.564 340.254 5.668 344.628 ; 
        RECT 5.132 340.254 5.236 344.628 ; 
        RECT 4.7 340.254 4.804 344.628 ; 
        RECT 4.268 340.254 4.372 344.628 ; 
        RECT 3.836 340.254 3.94 344.628 ; 
        RECT 3.404 340.254 3.508 344.628 ; 
        RECT 2.972 340.254 3.076 344.628 ; 
        RECT 2.54 340.254 2.644 344.628 ; 
        RECT 2.108 340.254 2.212 344.628 ; 
        RECT 1.676 340.254 1.78 344.628 ; 
        RECT 1.244 340.254 1.348 344.628 ; 
        RECT 0.812 340.254 0.916 344.628 ; 
        RECT 0 340.254 0.34 344.628 ; 
        RECT 20.72 344.574 21.232 348.948 ; 
        RECT 20.664 347.236 21.232 348.526 ; 
        RECT 20.072 346.144 20.32 348.948 ; 
        RECT 20.016 347.382 20.32 347.996 ; 
        RECT 20.072 344.574 20.176 348.948 ; 
        RECT 20.072 345.058 20.232 346.016 ; 
        RECT 20.072 344.574 20.32 344.93 ; 
        RECT 18.884 346.376 19.708 348.948 ; 
        RECT 19.604 344.574 19.708 348.948 ; 
        RECT 18.884 347.484 19.764 348.516 ; 
        RECT 18.884 344.574 19.276 348.948 ; 
        RECT 17.216 344.574 17.548 348.948 ; 
        RECT 17.216 344.928 17.604 348.67 ; 
        RECT 38.108 344.574 38.448 348.948 ; 
        RECT 37.532 344.574 37.636 348.948 ; 
        RECT 37.1 344.574 37.204 348.948 ; 
        RECT 36.668 344.574 36.772 348.948 ; 
        RECT 36.236 344.574 36.34 348.948 ; 
        RECT 35.804 344.574 35.908 348.948 ; 
        RECT 35.372 344.574 35.476 348.948 ; 
        RECT 34.94 344.574 35.044 348.948 ; 
        RECT 34.508 344.574 34.612 348.948 ; 
        RECT 34.076 344.574 34.18 348.948 ; 
        RECT 33.644 344.574 33.748 348.948 ; 
        RECT 33.212 344.574 33.316 348.948 ; 
        RECT 32.78 344.574 32.884 348.948 ; 
        RECT 32.348 344.574 32.452 348.948 ; 
        RECT 31.916 344.574 32.02 348.948 ; 
        RECT 31.484 344.574 31.588 348.948 ; 
        RECT 31.052 344.574 31.156 348.948 ; 
        RECT 30.62 344.574 30.724 348.948 ; 
        RECT 30.188 344.574 30.292 348.948 ; 
        RECT 29.756 344.574 29.86 348.948 ; 
        RECT 29.324 344.574 29.428 348.948 ; 
        RECT 28.892 344.574 28.996 348.948 ; 
        RECT 28.46 344.574 28.564 348.948 ; 
        RECT 28.028 344.574 28.132 348.948 ; 
        RECT 27.596 344.574 27.7 348.948 ; 
        RECT 27.164 344.574 27.268 348.948 ; 
        RECT 26.732 344.574 26.836 348.948 ; 
        RECT 26.3 344.574 26.404 348.948 ; 
        RECT 25.868 344.574 25.972 348.948 ; 
        RECT 25.436 344.574 25.54 348.948 ; 
        RECT 25.004 344.574 25.108 348.948 ; 
        RECT 24.572 344.574 24.676 348.948 ; 
        RECT 24.14 344.574 24.244 348.948 ; 
        RECT 23.708 344.574 23.812 348.948 ; 
        RECT 22.856 344.574 23.164 348.948 ; 
        RECT 15.284 344.574 15.592 348.948 ; 
        RECT 14.636 344.574 14.74 348.948 ; 
        RECT 14.204 344.574 14.308 348.948 ; 
        RECT 13.772 344.574 13.876 348.948 ; 
        RECT 13.34 344.574 13.444 348.948 ; 
        RECT 12.908 344.574 13.012 348.948 ; 
        RECT 12.476 344.574 12.58 348.948 ; 
        RECT 12.044 344.574 12.148 348.948 ; 
        RECT 11.612 344.574 11.716 348.948 ; 
        RECT 11.18 344.574 11.284 348.948 ; 
        RECT 10.748 344.574 10.852 348.948 ; 
        RECT 10.316 344.574 10.42 348.948 ; 
        RECT 9.884 344.574 9.988 348.948 ; 
        RECT 9.452 344.574 9.556 348.948 ; 
        RECT 9.02 344.574 9.124 348.948 ; 
        RECT 8.588 344.574 8.692 348.948 ; 
        RECT 8.156 344.574 8.26 348.948 ; 
        RECT 7.724 344.574 7.828 348.948 ; 
        RECT 7.292 344.574 7.396 348.948 ; 
        RECT 6.86 344.574 6.964 348.948 ; 
        RECT 6.428 344.574 6.532 348.948 ; 
        RECT 5.996 344.574 6.1 348.948 ; 
        RECT 5.564 344.574 5.668 348.948 ; 
        RECT 5.132 344.574 5.236 348.948 ; 
        RECT 4.7 344.574 4.804 348.948 ; 
        RECT 4.268 344.574 4.372 348.948 ; 
        RECT 3.836 344.574 3.94 348.948 ; 
        RECT 3.404 344.574 3.508 348.948 ; 
        RECT 2.972 344.574 3.076 348.948 ; 
        RECT 2.54 344.574 2.644 348.948 ; 
        RECT 2.108 344.574 2.212 348.948 ; 
        RECT 1.676 344.574 1.78 348.948 ; 
        RECT 1.244 344.574 1.348 348.948 ; 
        RECT 0.812 344.574 0.916 348.948 ; 
        RECT 0 344.574 0.34 348.948 ; 
        RECT 20.72 348.894 21.232 353.268 ; 
        RECT 20.664 351.556 21.232 352.846 ; 
        RECT 20.072 350.464 20.32 353.268 ; 
        RECT 20.016 351.702 20.32 352.316 ; 
        RECT 20.072 348.894 20.176 353.268 ; 
        RECT 20.072 349.378 20.232 350.336 ; 
        RECT 20.072 348.894 20.32 349.25 ; 
        RECT 18.884 350.696 19.708 353.268 ; 
        RECT 19.604 348.894 19.708 353.268 ; 
        RECT 18.884 351.804 19.764 352.836 ; 
        RECT 18.884 348.894 19.276 353.268 ; 
        RECT 17.216 348.894 17.548 353.268 ; 
        RECT 17.216 349.248 17.604 352.99 ; 
        RECT 38.108 348.894 38.448 353.268 ; 
        RECT 37.532 348.894 37.636 353.268 ; 
        RECT 37.1 348.894 37.204 353.268 ; 
        RECT 36.668 348.894 36.772 353.268 ; 
        RECT 36.236 348.894 36.34 353.268 ; 
        RECT 35.804 348.894 35.908 353.268 ; 
        RECT 35.372 348.894 35.476 353.268 ; 
        RECT 34.94 348.894 35.044 353.268 ; 
        RECT 34.508 348.894 34.612 353.268 ; 
        RECT 34.076 348.894 34.18 353.268 ; 
        RECT 33.644 348.894 33.748 353.268 ; 
        RECT 33.212 348.894 33.316 353.268 ; 
        RECT 32.78 348.894 32.884 353.268 ; 
        RECT 32.348 348.894 32.452 353.268 ; 
        RECT 31.916 348.894 32.02 353.268 ; 
        RECT 31.484 348.894 31.588 353.268 ; 
        RECT 31.052 348.894 31.156 353.268 ; 
        RECT 30.62 348.894 30.724 353.268 ; 
        RECT 30.188 348.894 30.292 353.268 ; 
        RECT 29.756 348.894 29.86 353.268 ; 
        RECT 29.324 348.894 29.428 353.268 ; 
        RECT 28.892 348.894 28.996 353.268 ; 
        RECT 28.46 348.894 28.564 353.268 ; 
        RECT 28.028 348.894 28.132 353.268 ; 
        RECT 27.596 348.894 27.7 353.268 ; 
        RECT 27.164 348.894 27.268 353.268 ; 
        RECT 26.732 348.894 26.836 353.268 ; 
        RECT 26.3 348.894 26.404 353.268 ; 
        RECT 25.868 348.894 25.972 353.268 ; 
        RECT 25.436 348.894 25.54 353.268 ; 
        RECT 25.004 348.894 25.108 353.268 ; 
        RECT 24.572 348.894 24.676 353.268 ; 
        RECT 24.14 348.894 24.244 353.268 ; 
        RECT 23.708 348.894 23.812 353.268 ; 
        RECT 22.856 348.894 23.164 353.268 ; 
        RECT 15.284 348.894 15.592 353.268 ; 
        RECT 14.636 348.894 14.74 353.268 ; 
        RECT 14.204 348.894 14.308 353.268 ; 
        RECT 13.772 348.894 13.876 353.268 ; 
        RECT 13.34 348.894 13.444 353.268 ; 
        RECT 12.908 348.894 13.012 353.268 ; 
        RECT 12.476 348.894 12.58 353.268 ; 
        RECT 12.044 348.894 12.148 353.268 ; 
        RECT 11.612 348.894 11.716 353.268 ; 
        RECT 11.18 348.894 11.284 353.268 ; 
        RECT 10.748 348.894 10.852 353.268 ; 
        RECT 10.316 348.894 10.42 353.268 ; 
        RECT 9.884 348.894 9.988 353.268 ; 
        RECT 9.452 348.894 9.556 353.268 ; 
        RECT 9.02 348.894 9.124 353.268 ; 
        RECT 8.588 348.894 8.692 353.268 ; 
        RECT 8.156 348.894 8.26 353.268 ; 
        RECT 7.724 348.894 7.828 353.268 ; 
        RECT 7.292 348.894 7.396 353.268 ; 
        RECT 6.86 348.894 6.964 353.268 ; 
        RECT 6.428 348.894 6.532 353.268 ; 
        RECT 5.996 348.894 6.1 353.268 ; 
        RECT 5.564 348.894 5.668 353.268 ; 
        RECT 5.132 348.894 5.236 353.268 ; 
        RECT 4.7 348.894 4.804 353.268 ; 
        RECT 4.268 348.894 4.372 353.268 ; 
        RECT 3.836 348.894 3.94 353.268 ; 
        RECT 3.404 348.894 3.508 353.268 ; 
        RECT 2.972 348.894 3.076 353.268 ; 
        RECT 2.54 348.894 2.644 353.268 ; 
        RECT 2.108 348.894 2.212 353.268 ; 
        RECT 1.676 348.894 1.78 353.268 ; 
        RECT 1.244 348.894 1.348 353.268 ; 
        RECT 0.812 348.894 0.916 353.268 ; 
        RECT 0 348.894 0.34 353.268 ; 
        RECT 20.72 353.214 21.232 357.588 ; 
        RECT 20.664 355.876 21.232 357.166 ; 
        RECT 20.072 354.784 20.32 357.588 ; 
        RECT 20.016 356.022 20.32 356.636 ; 
        RECT 20.072 353.214 20.176 357.588 ; 
        RECT 20.072 353.698 20.232 354.656 ; 
        RECT 20.072 353.214 20.32 353.57 ; 
        RECT 18.884 355.016 19.708 357.588 ; 
        RECT 19.604 353.214 19.708 357.588 ; 
        RECT 18.884 356.124 19.764 357.156 ; 
        RECT 18.884 353.214 19.276 357.588 ; 
        RECT 17.216 353.214 17.548 357.588 ; 
        RECT 17.216 353.568 17.604 357.31 ; 
        RECT 38.108 353.214 38.448 357.588 ; 
        RECT 37.532 353.214 37.636 357.588 ; 
        RECT 37.1 353.214 37.204 357.588 ; 
        RECT 36.668 353.214 36.772 357.588 ; 
        RECT 36.236 353.214 36.34 357.588 ; 
        RECT 35.804 353.214 35.908 357.588 ; 
        RECT 35.372 353.214 35.476 357.588 ; 
        RECT 34.94 353.214 35.044 357.588 ; 
        RECT 34.508 353.214 34.612 357.588 ; 
        RECT 34.076 353.214 34.18 357.588 ; 
        RECT 33.644 353.214 33.748 357.588 ; 
        RECT 33.212 353.214 33.316 357.588 ; 
        RECT 32.78 353.214 32.884 357.588 ; 
        RECT 32.348 353.214 32.452 357.588 ; 
        RECT 31.916 353.214 32.02 357.588 ; 
        RECT 31.484 353.214 31.588 357.588 ; 
        RECT 31.052 353.214 31.156 357.588 ; 
        RECT 30.62 353.214 30.724 357.588 ; 
        RECT 30.188 353.214 30.292 357.588 ; 
        RECT 29.756 353.214 29.86 357.588 ; 
        RECT 29.324 353.214 29.428 357.588 ; 
        RECT 28.892 353.214 28.996 357.588 ; 
        RECT 28.46 353.214 28.564 357.588 ; 
        RECT 28.028 353.214 28.132 357.588 ; 
        RECT 27.596 353.214 27.7 357.588 ; 
        RECT 27.164 353.214 27.268 357.588 ; 
        RECT 26.732 353.214 26.836 357.588 ; 
        RECT 26.3 353.214 26.404 357.588 ; 
        RECT 25.868 353.214 25.972 357.588 ; 
        RECT 25.436 353.214 25.54 357.588 ; 
        RECT 25.004 353.214 25.108 357.588 ; 
        RECT 24.572 353.214 24.676 357.588 ; 
        RECT 24.14 353.214 24.244 357.588 ; 
        RECT 23.708 353.214 23.812 357.588 ; 
        RECT 22.856 353.214 23.164 357.588 ; 
        RECT 15.284 353.214 15.592 357.588 ; 
        RECT 14.636 353.214 14.74 357.588 ; 
        RECT 14.204 353.214 14.308 357.588 ; 
        RECT 13.772 353.214 13.876 357.588 ; 
        RECT 13.34 353.214 13.444 357.588 ; 
        RECT 12.908 353.214 13.012 357.588 ; 
        RECT 12.476 353.214 12.58 357.588 ; 
        RECT 12.044 353.214 12.148 357.588 ; 
        RECT 11.612 353.214 11.716 357.588 ; 
        RECT 11.18 353.214 11.284 357.588 ; 
        RECT 10.748 353.214 10.852 357.588 ; 
        RECT 10.316 353.214 10.42 357.588 ; 
        RECT 9.884 353.214 9.988 357.588 ; 
        RECT 9.452 353.214 9.556 357.588 ; 
        RECT 9.02 353.214 9.124 357.588 ; 
        RECT 8.588 353.214 8.692 357.588 ; 
        RECT 8.156 353.214 8.26 357.588 ; 
        RECT 7.724 353.214 7.828 357.588 ; 
        RECT 7.292 353.214 7.396 357.588 ; 
        RECT 6.86 353.214 6.964 357.588 ; 
        RECT 6.428 353.214 6.532 357.588 ; 
        RECT 5.996 353.214 6.1 357.588 ; 
        RECT 5.564 353.214 5.668 357.588 ; 
        RECT 5.132 353.214 5.236 357.588 ; 
        RECT 4.7 353.214 4.804 357.588 ; 
        RECT 4.268 353.214 4.372 357.588 ; 
        RECT 3.836 353.214 3.94 357.588 ; 
        RECT 3.404 353.214 3.508 357.588 ; 
        RECT 2.972 353.214 3.076 357.588 ; 
        RECT 2.54 353.214 2.644 357.588 ; 
        RECT 2.108 353.214 2.212 357.588 ; 
        RECT 1.676 353.214 1.78 357.588 ; 
        RECT 1.244 353.214 1.348 357.588 ; 
        RECT 0.812 353.214 0.916 357.588 ; 
        RECT 0 353.214 0.34 357.588 ; 
        RECT 20.72 357.534 21.232 361.908 ; 
        RECT 20.664 360.196 21.232 361.486 ; 
        RECT 20.072 359.104 20.32 361.908 ; 
        RECT 20.016 360.342 20.32 360.956 ; 
        RECT 20.072 357.534 20.176 361.908 ; 
        RECT 20.072 358.018 20.232 358.976 ; 
        RECT 20.072 357.534 20.32 357.89 ; 
        RECT 18.884 359.336 19.708 361.908 ; 
        RECT 19.604 357.534 19.708 361.908 ; 
        RECT 18.884 360.444 19.764 361.476 ; 
        RECT 18.884 357.534 19.276 361.908 ; 
        RECT 17.216 357.534 17.548 361.908 ; 
        RECT 17.216 357.888 17.604 361.63 ; 
        RECT 38.108 357.534 38.448 361.908 ; 
        RECT 37.532 357.534 37.636 361.908 ; 
        RECT 37.1 357.534 37.204 361.908 ; 
        RECT 36.668 357.534 36.772 361.908 ; 
        RECT 36.236 357.534 36.34 361.908 ; 
        RECT 35.804 357.534 35.908 361.908 ; 
        RECT 35.372 357.534 35.476 361.908 ; 
        RECT 34.94 357.534 35.044 361.908 ; 
        RECT 34.508 357.534 34.612 361.908 ; 
        RECT 34.076 357.534 34.18 361.908 ; 
        RECT 33.644 357.534 33.748 361.908 ; 
        RECT 33.212 357.534 33.316 361.908 ; 
        RECT 32.78 357.534 32.884 361.908 ; 
        RECT 32.348 357.534 32.452 361.908 ; 
        RECT 31.916 357.534 32.02 361.908 ; 
        RECT 31.484 357.534 31.588 361.908 ; 
        RECT 31.052 357.534 31.156 361.908 ; 
        RECT 30.62 357.534 30.724 361.908 ; 
        RECT 30.188 357.534 30.292 361.908 ; 
        RECT 29.756 357.534 29.86 361.908 ; 
        RECT 29.324 357.534 29.428 361.908 ; 
        RECT 28.892 357.534 28.996 361.908 ; 
        RECT 28.46 357.534 28.564 361.908 ; 
        RECT 28.028 357.534 28.132 361.908 ; 
        RECT 27.596 357.534 27.7 361.908 ; 
        RECT 27.164 357.534 27.268 361.908 ; 
        RECT 26.732 357.534 26.836 361.908 ; 
        RECT 26.3 357.534 26.404 361.908 ; 
        RECT 25.868 357.534 25.972 361.908 ; 
        RECT 25.436 357.534 25.54 361.908 ; 
        RECT 25.004 357.534 25.108 361.908 ; 
        RECT 24.572 357.534 24.676 361.908 ; 
        RECT 24.14 357.534 24.244 361.908 ; 
        RECT 23.708 357.534 23.812 361.908 ; 
        RECT 22.856 357.534 23.164 361.908 ; 
        RECT 15.284 357.534 15.592 361.908 ; 
        RECT 14.636 357.534 14.74 361.908 ; 
        RECT 14.204 357.534 14.308 361.908 ; 
        RECT 13.772 357.534 13.876 361.908 ; 
        RECT 13.34 357.534 13.444 361.908 ; 
        RECT 12.908 357.534 13.012 361.908 ; 
        RECT 12.476 357.534 12.58 361.908 ; 
        RECT 12.044 357.534 12.148 361.908 ; 
        RECT 11.612 357.534 11.716 361.908 ; 
        RECT 11.18 357.534 11.284 361.908 ; 
        RECT 10.748 357.534 10.852 361.908 ; 
        RECT 10.316 357.534 10.42 361.908 ; 
        RECT 9.884 357.534 9.988 361.908 ; 
        RECT 9.452 357.534 9.556 361.908 ; 
        RECT 9.02 357.534 9.124 361.908 ; 
        RECT 8.588 357.534 8.692 361.908 ; 
        RECT 8.156 357.534 8.26 361.908 ; 
        RECT 7.724 357.534 7.828 361.908 ; 
        RECT 7.292 357.534 7.396 361.908 ; 
        RECT 6.86 357.534 6.964 361.908 ; 
        RECT 6.428 357.534 6.532 361.908 ; 
        RECT 5.996 357.534 6.1 361.908 ; 
        RECT 5.564 357.534 5.668 361.908 ; 
        RECT 5.132 357.534 5.236 361.908 ; 
        RECT 4.7 357.534 4.804 361.908 ; 
        RECT 4.268 357.534 4.372 361.908 ; 
        RECT 3.836 357.534 3.94 361.908 ; 
        RECT 3.404 357.534 3.508 361.908 ; 
        RECT 2.972 357.534 3.076 361.908 ; 
        RECT 2.54 357.534 2.644 361.908 ; 
        RECT 2.108 357.534 2.212 361.908 ; 
        RECT 1.676 357.534 1.78 361.908 ; 
        RECT 1.244 357.534 1.348 361.908 ; 
        RECT 0.812 357.534 0.916 361.908 ; 
        RECT 0 357.534 0.34 361.908 ; 
        RECT 20.72 361.854 21.232 366.228 ; 
        RECT 20.664 364.516 21.232 365.806 ; 
        RECT 20.072 363.424 20.32 366.228 ; 
        RECT 20.016 364.662 20.32 365.276 ; 
        RECT 20.072 361.854 20.176 366.228 ; 
        RECT 20.072 362.338 20.232 363.296 ; 
        RECT 20.072 361.854 20.32 362.21 ; 
        RECT 18.884 363.656 19.708 366.228 ; 
        RECT 19.604 361.854 19.708 366.228 ; 
        RECT 18.884 364.764 19.764 365.796 ; 
        RECT 18.884 361.854 19.276 366.228 ; 
        RECT 17.216 361.854 17.548 366.228 ; 
        RECT 17.216 362.208 17.604 365.95 ; 
        RECT 38.108 361.854 38.448 366.228 ; 
        RECT 37.532 361.854 37.636 366.228 ; 
        RECT 37.1 361.854 37.204 366.228 ; 
        RECT 36.668 361.854 36.772 366.228 ; 
        RECT 36.236 361.854 36.34 366.228 ; 
        RECT 35.804 361.854 35.908 366.228 ; 
        RECT 35.372 361.854 35.476 366.228 ; 
        RECT 34.94 361.854 35.044 366.228 ; 
        RECT 34.508 361.854 34.612 366.228 ; 
        RECT 34.076 361.854 34.18 366.228 ; 
        RECT 33.644 361.854 33.748 366.228 ; 
        RECT 33.212 361.854 33.316 366.228 ; 
        RECT 32.78 361.854 32.884 366.228 ; 
        RECT 32.348 361.854 32.452 366.228 ; 
        RECT 31.916 361.854 32.02 366.228 ; 
        RECT 31.484 361.854 31.588 366.228 ; 
        RECT 31.052 361.854 31.156 366.228 ; 
        RECT 30.62 361.854 30.724 366.228 ; 
        RECT 30.188 361.854 30.292 366.228 ; 
        RECT 29.756 361.854 29.86 366.228 ; 
        RECT 29.324 361.854 29.428 366.228 ; 
        RECT 28.892 361.854 28.996 366.228 ; 
        RECT 28.46 361.854 28.564 366.228 ; 
        RECT 28.028 361.854 28.132 366.228 ; 
        RECT 27.596 361.854 27.7 366.228 ; 
        RECT 27.164 361.854 27.268 366.228 ; 
        RECT 26.732 361.854 26.836 366.228 ; 
        RECT 26.3 361.854 26.404 366.228 ; 
        RECT 25.868 361.854 25.972 366.228 ; 
        RECT 25.436 361.854 25.54 366.228 ; 
        RECT 25.004 361.854 25.108 366.228 ; 
        RECT 24.572 361.854 24.676 366.228 ; 
        RECT 24.14 361.854 24.244 366.228 ; 
        RECT 23.708 361.854 23.812 366.228 ; 
        RECT 22.856 361.854 23.164 366.228 ; 
        RECT 15.284 361.854 15.592 366.228 ; 
        RECT 14.636 361.854 14.74 366.228 ; 
        RECT 14.204 361.854 14.308 366.228 ; 
        RECT 13.772 361.854 13.876 366.228 ; 
        RECT 13.34 361.854 13.444 366.228 ; 
        RECT 12.908 361.854 13.012 366.228 ; 
        RECT 12.476 361.854 12.58 366.228 ; 
        RECT 12.044 361.854 12.148 366.228 ; 
        RECT 11.612 361.854 11.716 366.228 ; 
        RECT 11.18 361.854 11.284 366.228 ; 
        RECT 10.748 361.854 10.852 366.228 ; 
        RECT 10.316 361.854 10.42 366.228 ; 
        RECT 9.884 361.854 9.988 366.228 ; 
        RECT 9.452 361.854 9.556 366.228 ; 
        RECT 9.02 361.854 9.124 366.228 ; 
        RECT 8.588 361.854 8.692 366.228 ; 
        RECT 8.156 361.854 8.26 366.228 ; 
        RECT 7.724 361.854 7.828 366.228 ; 
        RECT 7.292 361.854 7.396 366.228 ; 
        RECT 6.86 361.854 6.964 366.228 ; 
        RECT 6.428 361.854 6.532 366.228 ; 
        RECT 5.996 361.854 6.1 366.228 ; 
        RECT 5.564 361.854 5.668 366.228 ; 
        RECT 5.132 361.854 5.236 366.228 ; 
        RECT 4.7 361.854 4.804 366.228 ; 
        RECT 4.268 361.854 4.372 366.228 ; 
        RECT 3.836 361.854 3.94 366.228 ; 
        RECT 3.404 361.854 3.508 366.228 ; 
        RECT 2.972 361.854 3.076 366.228 ; 
        RECT 2.54 361.854 2.644 366.228 ; 
        RECT 2.108 361.854 2.212 366.228 ; 
        RECT 1.676 361.854 1.78 366.228 ; 
        RECT 1.244 361.854 1.348 366.228 ; 
        RECT 0.812 361.854 0.916 366.228 ; 
        RECT 0 361.854 0.34 366.228 ; 
        RECT 20.72 366.174 21.232 370.548 ; 
        RECT 20.664 368.836 21.232 370.126 ; 
        RECT 20.072 367.744 20.32 370.548 ; 
        RECT 20.016 368.982 20.32 369.596 ; 
        RECT 20.072 366.174 20.176 370.548 ; 
        RECT 20.072 366.658 20.232 367.616 ; 
        RECT 20.072 366.174 20.32 366.53 ; 
        RECT 18.884 367.976 19.708 370.548 ; 
        RECT 19.604 366.174 19.708 370.548 ; 
        RECT 18.884 369.084 19.764 370.116 ; 
        RECT 18.884 366.174 19.276 370.548 ; 
        RECT 17.216 366.174 17.548 370.548 ; 
        RECT 17.216 366.528 17.604 370.27 ; 
        RECT 38.108 366.174 38.448 370.548 ; 
        RECT 37.532 366.174 37.636 370.548 ; 
        RECT 37.1 366.174 37.204 370.548 ; 
        RECT 36.668 366.174 36.772 370.548 ; 
        RECT 36.236 366.174 36.34 370.548 ; 
        RECT 35.804 366.174 35.908 370.548 ; 
        RECT 35.372 366.174 35.476 370.548 ; 
        RECT 34.94 366.174 35.044 370.548 ; 
        RECT 34.508 366.174 34.612 370.548 ; 
        RECT 34.076 366.174 34.18 370.548 ; 
        RECT 33.644 366.174 33.748 370.548 ; 
        RECT 33.212 366.174 33.316 370.548 ; 
        RECT 32.78 366.174 32.884 370.548 ; 
        RECT 32.348 366.174 32.452 370.548 ; 
        RECT 31.916 366.174 32.02 370.548 ; 
        RECT 31.484 366.174 31.588 370.548 ; 
        RECT 31.052 366.174 31.156 370.548 ; 
        RECT 30.62 366.174 30.724 370.548 ; 
        RECT 30.188 366.174 30.292 370.548 ; 
        RECT 29.756 366.174 29.86 370.548 ; 
        RECT 29.324 366.174 29.428 370.548 ; 
        RECT 28.892 366.174 28.996 370.548 ; 
        RECT 28.46 366.174 28.564 370.548 ; 
        RECT 28.028 366.174 28.132 370.548 ; 
        RECT 27.596 366.174 27.7 370.548 ; 
        RECT 27.164 366.174 27.268 370.548 ; 
        RECT 26.732 366.174 26.836 370.548 ; 
        RECT 26.3 366.174 26.404 370.548 ; 
        RECT 25.868 366.174 25.972 370.548 ; 
        RECT 25.436 366.174 25.54 370.548 ; 
        RECT 25.004 366.174 25.108 370.548 ; 
        RECT 24.572 366.174 24.676 370.548 ; 
        RECT 24.14 366.174 24.244 370.548 ; 
        RECT 23.708 366.174 23.812 370.548 ; 
        RECT 22.856 366.174 23.164 370.548 ; 
        RECT 15.284 366.174 15.592 370.548 ; 
        RECT 14.636 366.174 14.74 370.548 ; 
        RECT 14.204 366.174 14.308 370.548 ; 
        RECT 13.772 366.174 13.876 370.548 ; 
        RECT 13.34 366.174 13.444 370.548 ; 
        RECT 12.908 366.174 13.012 370.548 ; 
        RECT 12.476 366.174 12.58 370.548 ; 
        RECT 12.044 366.174 12.148 370.548 ; 
        RECT 11.612 366.174 11.716 370.548 ; 
        RECT 11.18 366.174 11.284 370.548 ; 
        RECT 10.748 366.174 10.852 370.548 ; 
        RECT 10.316 366.174 10.42 370.548 ; 
        RECT 9.884 366.174 9.988 370.548 ; 
        RECT 9.452 366.174 9.556 370.548 ; 
        RECT 9.02 366.174 9.124 370.548 ; 
        RECT 8.588 366.174 8.692 370.548 ; 
        RECT 8.156 366.174 8.26 370.548 ; 
        RECT 7.724 366.174 7.828 370.548 ; 
        RECT 7.292 366.174 7.396 370.548 ; 
        RECT 6.86 366.174 6.964 370.548 ; 
        RECT 6.428 366.174 6.532 370.548 ; 
        RECT 5.996 366.174 6.1 370.548 ; 
        RECT 5.564 366.174 5.668 370.548 ; 
        RECT 5.132 366.174 5.236 370.548 ; 
        RECT 4.7 366.174 4.804 370.548 ; 
        RECT 4.268 366.174 4.372 370.548 ; 
        RECT 3.836 366.174 3.94 370.548 ; 
        RECT 3.404 366.174 3.508 370.548 ; 
        RECT 2.972 366.174 3.076 370.548 ; 
        RECT 2.54 366.174 2.644 370.548 ; 
        RECT 2.108 366.174 2.212 370.548 ; 
        RECT 1.676 366.174 1.78 370.548 ; 
        RECT 1.244 366.174 1.348 370.548 ; 
        RECT 0.812 366.174 0.916 370.548 ; 
        RECT 0 366.174 0.34 370.548 ; 
        RECT 20.72 370.494 21.232 374.868 ; 
        RECT 20.664 373.156 21.232 374.446 ; 
        RECT 20.072 372.064 20.32 374.868 ; 
        RECT 20.016 373.302 20.32 373.916 ; 
        RECT 20.072 370.494 20.176 374.868 ; 
        RECT 20.072 370.978 20.232 371.936 ; 
        RECT 20.072 370.494 20.32 370.85 ; 
        RECT 18.884 372.296 19.708 374.868 ; 
        RECT 19.604 370.494 19.708 374.868 ; 
        RECT 18.884 373.404 19.764 374.436 ; 
        RECT 18.884 370.494 19.276 374.868 ; 
        RECT 17.216 370.494 17.548 374.868 ; 
        RECT 17.216 370.848 17.604 374.59 ; 
        RECT 38.108 370.494 38.448 374.868 ; 
        RECT 37.532 370.494 37.636 374.868 ; 
        RECT 37.1 370.494 37.204 374.868 ; 
        RECT 36.668 370.494 36.772 374.868 ; 
        RECT 36.236 370.494 36.34 374.868 ; 
        RECT 35.804 370.494 35.908 374.868 ; 
        RECT 35.372 370.494 35.476 374.868 ; 
        RECT 34.94 370.494 35.044 374.868 ; 
        RECT 34.508 370.494 34.612 374.868 ; 
        RECT 34.076 370.494 34.18 374.868 ; 
        RECT 33.644 370.494 33.748 374.868 ; 
        RECT 33.212 370.494 33.316 374.868 ; 
        RECT 32.78 370.494 32.884 374.868 ; 
        RECT 32.348 370.494 32.452 374.868 ; 
        RECT 31.916 370.494 32.02 374.868 ; 
        RECT 31.484 370.494 31.588 374.868 ; 
        RECT 31.052 370.494 31.156 374.868 ; 
        RECT 30.62 370.494 30.724 374.868 ; 
        RECT 30.188 370.494 30.292 374.868 ; 
        RECT 29.756 370.494 29.86 374.868 ; 
        RECT 29.324 370.494 29.428 374.868 ; 
        RECT 28.892 370.494 28.996 374.868 ; 
        RECT 28.46 370.494 28.564 374.868 ; 
        RECT 28.028 370.494 28.132 374.868 ; 
        RECT 27.596 370.494 27.7 374.868 ; 
        RECT 27.164 370.494 27.268 374.868 ; 
        RECT 26.732 370.494 26.836 374.868 ; 
        RECT 26.3 370.494 26.404 374.868 ; 
        RECT 25.868 370.494 25.972 374.868 ; 
        RECT 25.436 370.494 25.54 374.868 ; 
        RECT 25.004 370.494 25.108 374.868 ; 
        RECT 24.572 370.494 24.676 374.868 ; 
        RECT 24.14 370.494 24.244 374.868 ; 
        RECT 23.708 370.494 23.812 374.868 ; 
        RECT 22.856 370.494 23.164 374.868 ; 
        RECT 15.284 370.494 15.592 374.868 ; 
        RECT 14.636 370.494 14.74 374.868 ; 
        RECT 14.204 370.494 14.308 374.868 ; 
        RECT 13.772 370.494 13.876 374.868 ; 
        RECT 13.34 370.494 13.444 374.868 ; 
        RECT 12.908 370.494 13.012 374.868 ; 
        RECT 12.476 370.494 12.58 374.868 ; 
        RECT 12.044 370.494 12.148 374.868 ; 
        RECT 11.612 370.494 11.716 374.868 ; 
        RECT 11.18 370.494 11.284 374.868 ; 
        RECT 10.748 370.494 10.852 374.868 ; 
        RECT 10.316 370.494 10.42 374.868 ; 
        RECT 9.884 370.494 9.988 374.868 ; 
        RECT 9.452 370.494 9.556 374.868 ; 
        RECT 9.02 370.494 9.124 374.868 ; 
        RECT 8.588 370.494 8.692 374.868 ; 
        RECT 8.156 370.494 8.26 374.868 ; 
        RECT 7.724 370.494 7.828 374.868 ; 
        RECT 7.292 370.494 7.396 374.868 ; 
        RECT 6.86 370.494 6.964 374.868 ; 
        RECT 6.428 370.494 6.532 374.868 ; 
        RECT 5.996 370.494 6.1 374.868 ; 
        RECT 5.564 370.494 5.668 374.868 ; 
        RECT 5.132 370.494 5.236 374.868 ; 
        RECT 4.7 370.494 4.804 374.868 ; 
        RECT 4.268 370.494 4.372 374.868 ; 
        RECT 3.836 370.494 3.94 374.868 ; 
        RECT 3.404 370.494 3.508 374.868 ; 
        RECT 2.972 370.494 3.076 374.868 ; 
        RECT 2.54 370.494 2.644 374.868 ; 
        RECT 2.108 370.494 2.212 374.868 ; 
        RECT 1.676 370.494 1.78 374.868 ; 
        RECT 1.244 370.494 1.348 374.868 ; 
        RECT 0.812 370.494 0.916 374.868 ; 
        RECT 0 370.494 0.34 374.868 ; 
        RECT 20.72 374.814 21.232 379.188 ; 
        RECT 20.664 377.476 21.232 378.766 ; 
        RECT 20.072 376.384 20.32 379.188 ; 
        RECT 20.016 377.622 20.32 378.236 ; 
        RECT 20.072 374.814 20.176 379.188 ; 
        RECT 20.072 375.298 20.232 376.256 ; 
        RECT 20.072 374.814 20.32 375.17 ; 
        RECT 18.884 376.616 19.708 379.188 ; 
        RECT 19.604 374.814 19.708 379.188 ; 
        RECT 18.884 377.724 19.764 378.756 ; 
        RECT 18.884 374.814 19.276 379.188 ; 
        RECT 17.216 374.814 17.548 379.188 ; 
        RECT 17.216 375.168 17.604 378.91 ; 
        RECT 38.108 374.814 38.448 379.188 ; 
        RECT 37.532 374.814 37.636 379.188 ; 
        RECT 37.1 374.814 37.204 379.188 ; 
        RECT 36.668 374.814 36.772 379.188 ; 
        RECT 36.236 374.814 36.34 379.188 ; 
        RECT 35.804 374.814 35.908 379.188 ; 
        RECT 35.372 374.814 35.476 379.188 ; 
        RECT 34.94 374.814 35.044 379.188 ; 
        RECT 34.508 374.814 34.612 379.188 ; 
        RECT 34.076 374.814 34.18 379.188 ; 
        RECT 33.644 374.814 33.748 379.188 ; 
        RECT 33.212 374.814 33.316 379.188 ; 
        RECT 32.78 374.814 32.884 379.188 ; 
        RECT 32.348 374.814 32.452 379.188 ; 
        RECT 31.916 374.814 32.02 379.188 ; 
        RECT 31.484 374.814 31.588 379.188 ; 
        RECT 31.052 374.814 31.156 379.188 ; 
        RECT 30.62 374.814 30.724 379.188 ; 
        RECT 30.188 374.814 30.292 379.188 ; 
        RECT 29.756 374.814 29.86 379.188 ; 
        RECT 29.324 374.814 29.428 379.188 ; 
        RECT 28.892 374.814 28.996 379.188 ; 
        RECT 28.46 374.814 28.564 379.188 ; 
        RECT 28.028 374.814 28.132 379.188 ; 
        RECT 27.596 374.814 27.7 379.188 ; 
        RECT 27.164 374.814 27.268 379.188 ; 
        RECT 26.732 374.814 26.836 379.188 ; 
        RECT 26.3 374.814 26.404 379.188 ; 
        RECT 25.868 374.814 25.972 379.188 ; 
        RECT 25.436 374.814 25.54 379.188 ; 
        RECT 25.004 374.814 25.108 379.188 ; 
        RECT 24.572 374.814 24.676 379.188 ; 
        RECT 24.14 374.814 24.244 379.188 ; 
        RECT 23.708 374.814 23.812 379.188 ; 
        RECT 22.856 374.814 23.164 379.188 ; 
        RECT 15.284 374.814 15.592 379.188 ; 
        RECT 14.636 374.814 14.74 379.188 ; 
        RECT 14.204 374.814 14.308 379.188 ; 
        RECT 13.772 374.814 13.876 379.188 ; 
        RECT 13.34 374.814 13.444 379.188 ; 
        RECT 12.908 374.814 13.012 379.188 ; 
        RECT 12.476 374.814 12.58 379.188 ; 
        RECT 12.044 374.814 12.148 379.188 ; 
        RECT 11.612 374.814 11.716 379.188 ; 
        RECT 11.18 374.814 11.284 379.188 ; 
        RECT 10.748 374.814 10.852 379.188 ; 
        RECT 10.316 374.814 10.42 379.188 ; 
        RECT 9.884 374.814 9.988 379.188 ; 
        RECT 9.452 374.814 9.556 379.188 ; 
        RECT 9.02 374.814 9.124 379.188 ; 
        RECT 8.588 374.814 8.692 379.188 ; 
        RECT 8.156 374.814 8.26 379.188 ; 
        RECT 7.724 374.814 7.828 379.188 ; 
        RECT 7.292 374.814 7.396 379.188 ; 
        RECT 6.86 374.814 6.964 379.188 ; 
        RECT 6.428 374.814 6.532 379.188 ; 
        RECT 5.996 374.814 6.1 379.188 ; 
        RECT 5.564 374.814 5.668 379.188 ; 
        RECT 5.132 374.814 5.236 379.188 ; 
        RECT 4.7 374.814 4.804 379.188 ; 
        RECT 4.268 374.814 4.372 379.188 ; 
        RECT 3.836 374.814 3.94 379.188 ; 
        RECT 3.404 374.814 3.508 379.188 ; 
        RECT 2.972 374.814 3.076 379.188 ; 
        RECT 2.54 374.814 2.644 379.188 ; 
        RECT 2.108 374.814 2.212 379.188 ; 
        RECT 1.676 374.814 1.78 379.188 ; 
        RECT 1.244 374.814 1.348 379.188 ; 
        RECT 0.812 374.814 0.916 379.188 ; 
        RECT 0 374.814 0.34 379.188 ; 
  LAYER V3 ; 
      RECT 0 4.88 38.448 5.4 ; 
      RECT 37.98 1.026 38.448 5.4 ; 
      RECT 23.364 4.496 37.908 5.4 ; 
      RECT 18.036 4.496 23.292 5.4 ; 
      RECT 15.156 1.026 17.676 5.4 ; 
      RECT 0.54 4.496 15.084 5.4 ; 
      RECT 0 1.026 0.468 5.4 ; 
      RECT 37.836 1.026 38.448 4.688 ; 
      RECT 23.58 1.026 37.764 5.4 ; 
      RECT 20.592 1.026 23.508 4.688 ; 
      RECT 19.944 1.808 20.448 5.4 ; 
      RECT 14.94 1.424 19.836 4.688 ; 
      RECT 0.684 1.026 14.868 5.4 ; 
      RECT 0 1.026 0.612 4.688 ; 
      RECT 20.376 1.026 38.448 4.304 ; 
      RECT 0 1.424 20.304 4.304 ; 
      RECT 19.476 1.026 38.448 1.712 ; 
      RECT 0 1.026 19.404 4.304 ; 
      RECT 0 1.026 38.448 1.328 ; 
      RECT 0 9.2 38.448 9.72 ; 
      RECT 37.98 5.346 38.448 9.72 ; 
      RECT 23.364 8.816 37.908 9.72 ; 
      RECT 18.036 8.816 23.292 9.72 ; 
      RECT 15.156 5.346 17.676 9.72 ; 
      RECT 0.54 8.816 15.084 9.72 ; 
      RECT 0 5.346 0.468 9.72 ; 
      RECT 37.836 5.346 38.448 9.008 ; 
      RECT 23.58 5.346 37.764 9.72 ; 
      RECT 20.592 5.346 23.508 9.008 ; 
      RECT 19.944 6.128 20.448 9.72 ; 
      RECT 14.94 5.744 19.836 9.008 ; 
      RECT 0.684 5.346 14.868 9.72 ; 
      RECT 0 5.346 0.612 9.008 ; 
      RECT 20.376 5.346 38.448 8.624 ; 
      RECT 0 5.744 20.304 8.624 ; 
      RECT 19.476 5.346 38.448 6.032 ; 
      RECT 0 5.346 19.404 8.624 ; 
      RECT 0 5.346 38.448 5.648 ; 
      RECT 0 13.52 38.448 14.04 ; 
      RECT 37.98 9.666 38.448 14.04 ; 
      RECT 23.364 13.136 37.908 14.04 ; 
      RECT 18.036 13.136 23.292 14.04 ; 
      RECT 15.156 9.666 17.676 14.04 ; 
      RECT 0.54 13.136 15.084 14.04 ; 
      RECT 0 9.666 0.468 14.04 ; 
      RECT 37.836 9.666 38.448 13.328 ; 
      RECT 23.58 9.666 37.764 14.04 ; 
      RECT 20.592 9.666 23.508 13.328 ; 
      RECT 19.944 10.448 20.448 14.04 ; 
      RECT 14.94 10.064 19.836 13.328 ; 
      RECT 0.684 9.666 14.868 14.04 ; 
      RECT 0 9.666 0.612 13.328 ; 
      RECT 20.376 9.666 38.448 12.944 ; 
      RECT 0 10.064 20.304 12.944 ; 
      RECT 19.476 9.666 38.448 10.352 ; 
      RECT 0 9.666 19.404 12.944 ; 
      RECT 0 9.666 38.448 9.968 ; 
      RECT 0 17.84 38.448 18.36 ; 
      RECT 37.98 13.986 38.448 18.36 ; 
      RECT 23.364 17.456 37.908 18.36 ; 
      RECT 18.036 17.456 23.292 18.36 ; 
      RECT 15.156 13.986 17.676 18.36 ; 
      RECT 0.54 17.456 15.084 18.36 ; 
      RECT 0 13.986 0.468 18.36 ; 
      RECT 37.836 13.986 38.448 17.648 ; 
      RECT 23.58 13.986 37.764 18.36 ; 
      RECT 20.592 13.986 23.508 17.648 ; 
      RECT 19.944 14.768 20.448 18.36 ; 
      RECT 14.94 14.384 19.836 17.648 ; 
      RECT 0.684 13.986 14.868 18.36 ; 
      RECT 0 13.986 0.612 17.648 ; 
      RECT 20.376 13.986 38.448 17.264 ; 
      RECT 0 14.384 20.304 17.264 ; 
      RECT 19.476 13.986 38.448 14.672 ; 
      RECT 0 13.986 19.404 17.264 ; 
      RECT 0 13.986 38.448 14.288 ; 
      RECT 0 22.16 38.448 22.68 ; 
      RECT 37.98 18.306 38.448 22.68 ; 
      RECT 23.364 21.776 37.908 22.68 ; 
      RECT 18.036 21.776 23.292 22.68 ; 
      RECT 15.156 18.306 17.676 22.68 ; 
      RECT 0.54 21.776 15.084 22.68 ; 
      RECT 0 18.306 0.468 22.68 ; 
      RECT 37.836 18.306 38.448 21.968 ; 
      RECT 23.58 18.306 37.764 22.68 ; 
      RECT 20.592 18.306 23.508 21.968 ; 
      RECT 19.944 19.088 20.448 22.68 ; 
      RECT 14.94 18.704 19.836 21.968 ; 
      RECT 0.684 18.306 14.868 22.68 ; 
      RECT 0 18.306 0.612 21.968 ; 
      RECT 20.376 18.306 38.448 21.584 ; 
      RECT 0 18.704 20.304 21.584 ; 
      RECT 19.476 18.306 38.448 18.992 ; 
      RECT 0 18.306 19.404 21.584 ; 
      RECT 0 18.306 38.448 18.608 ; 
      RECT 0 26.48 38.448 27 ; 
      RECT 37.98 22.626 38.448 27 ; 
      RECT 23.364 26.096 37.908 27 ; 
      RECT 18.036 26.096 23.292 27 ; 
      RECT 15.156 22.626 17.676 27 ; 
      RECT 0.54 26.096 15.084 27 ; 
      RECT 0 22.626 0.468 27 ; 
      RECT 37.836 22.626 38.448 26.288 ; 
      RECT 23.58 22.626 37.764 27 ; 
      RECT 20.592 22.626 23.508 26.288 ; 
      RECT 19.944 23.408 20.448 27 ; 
      RECT 14.94 23.024 19.836 26.288 ; 
      RECT 0.684 22.626 14.868 27 ; 
      RECT 0 22.626 0.612 26.288 ; 
      RECT 20.376 22.626 38.448 25.904 ; 
      RECT 0 23.024 20.304 25.904 ; 
      RECT 19.476 22.626 38.448 23.312 ; 
      RECT 0 22.626 19.404 25.904 ; 
      RECT 0 22.626 38.448 22.928 ; 
      RECT 0 30.8 38.448 31.32 ; 
      RECT 37.98 26.946 38.448 31.32 ; 
      RECT 23.364 30.416 37.908 31.32 ; 
      RECT 18.036 30.416 23.292 31.32 ; 
      RECT 15.156 26.946 17.676 31.32 ; 
      RECT 0.54 30.416 15.084 31.32 ; 
      RECT 0 26.946 0.468 31.32 ; 
      RECT 37.836 26.946 38.448 30.608 ; 
      RECT 23.58 26.946 37.764 31.32 ; 
      RECT 20.592 26.946 23.508 30.608 ; 
      RECT 19.944 27.728 20.448 31.32 ; 
      RECT 14.94 27.344 19.836 30.608 ; 
      RECT 0.684 26.946 14.868 31.32 ; 
      RECT 0 26.946 0.612 30.608 ; 
      RECT 20.376 26.946 38.448 30.224 ; 
      RECT 0 27.344 20.304 30.224 ; 
      RECT 19.476 26.946 38.448 27.632 ; 
      RECT 0 26.946 19.404 30.224 ; 
      RECT 0 26.946 38.448 27.248 ; 
      RECT 0 35.12 38.448 35.64 ; 
      RECT 37.98 31.266 38.448 35.64 ; 
      RECT 23.364 34.736 37.908 35.64 ; 
      RECT 18.036 34.736 23.292 35.64 ; 
      RECT 15.156 31.266 17.676 35.64 ; 
      RECT 0.54 34.736 15.084 35.64 ; 
      RECT 0 31.266 0.468 35.64 ; 
      RECT 37.836 31.266 38.448 34.928 ; 
      RECT 23.58 31.266 37.764 35.64 ; 
      RECT 20.592 31.266 23.508 34.928 ; 
      RECT 19.944 32.048 20.448 35.64 ; 
      RECT 14.94 31.664 19.836 34.928 ; 
      RECT 0.684 31.266 14.868 35.64 ; 
      RECT 0 31.266 0.612 34.928 ; 
      RECT 20.376 31.266 38.448 34.544 ; 
      RECT 0 31.664 20.304 34.544 ; 
      RECT 19.476 31.266 38.448 31.952 ; 
      RECT 0 31.266 19.404 34.544 ; 
      RECT 0 31.266 38.448 31.568 ; 
      RECT 0 39.44 38.448 39.96 ; 
      RECT 37.98 35.586 38.448 39.96 ; 
      RECT 23.364 39.056 37.908 39.96 ; 
      RECT 18.036 39.056 23.292 39.96 ; 
      RECT 15.156 35.586 17.676 39.96 ; 
      RECT 0.54 39.056 15.084 39.96 ; 
      RECT 0 35.586 0.468 39.96 ; 
      RECT 37.836 35.586 38.448 39.248 ; 
      RECT 23.58 35.586 37.764 39.96 ; 
      RECT 20.592 35.586 23.508 39.248 ; 
      RECT 19.944 36.368 20.448 39.96 ; 
      RECT 14.94 35.984 19.836 39.248 ; 
      RECT 0.684 35.586 14.868 39.96 ; 
      RECT 0 35.586 0.612 39.248 ; 
      RECT 20.376 35.586 38.448 38.864 ; 
      RECT 0 35.984 20.304 38.864 ; 
      RECT 19.476 35.586 38.448 36.272 ; 
      RECT 0 35.586 19.404 38.864 ; 
      RECT 0 35.586 38.448 35.888 ; 
      RECT 0 43.76 38.448 44.28 ; 
      RECT 37.98 39.906 38.448 44.28 ; 
      RECT 23.364 43.376 37.908 44.28 ; 
      RECT 18.036 43.376 23.292 44.28 ; 
      RECT 15.156 39.906 17.676 44.28 ; 
      RECT 0.54 43.376 15.084 44.28 ; 
      RECT 0 39.906 0.468 44.28 ; 
      RECT 37.836 39.906 38.448 43.568 ; 
      RECT 23.58 39.906 37.764 44.28 ; 
      RECT 20.592 39.906 23.508 43.568 ; 
      RECT 19.944 40.688 20.448 44.28 ; 
      RECT 14.94 40.304 19.836 43.568 ; 
      RECT 0.684 39.906 14.868 44.28 ; 
      RECT 0 39.906 0.612 43.568 ; 
      RECT 20.376 39.906 38.448 43.184 ; 
      RECT 0 40.304 20.304 43.184 ; 
      RECT 19.476 39.906 38.448 40.592 ; 
      RECT 0 39.906 19.404 43.184 ; 
      RECT 0 39.906 38.448 40.208 ; 
      RECT 0 48.08 38.448 48.6 ; 
      RECT 37.98 44.226 38.448 48.6 ; 
      RECT 23.364 47.696 37.908 48.6 ; 
      RECT 18.036 47.696 23.292 48.6 ; 
      RECT 15.156 44.226 17.676 48.6 ; 
      RECT 0.54 47.696 15.084 48.6 ; 
      RECT 0 44.226 0.468 48.6 ; 
      RECT 37.836 44.226 38.448 47.888 ; 
      RECT 23.58 44.226 37.764 48.6 ; 
      RECT 20.592 44.226 23.508 47.888 ; 
      RECT 19.944 45.008 20.448 48.6 ; 
      RECT 14.94 44.624 19.836 47.888 ; 
      RECT 0.684 44.226 14.868 48.6 ; 
      RECT 0 44.226 0.612 47.888 ; 
      RECT 20.376 44.226 38.448 47.504 ; 
      RECT 0 44.624 20.304 47.504 ; 
      RECT 19.476 44.226 38.448 44.912 ; 
      RECT 0 44.226 19.404 47.504 ; 
      RECT 0 44.226 38.448 44.528 ; 
      RECT 0 52.4 38.448 52.92 ; 
      RECT 37.98 48.546 38.448 52.92 ; 
      RECT 23.364 52.016 37.908 52.92 ; 
      RECT 18.036 52.016 23.292 52.92 ; 
      RECT 15.156 48.546 17.676 52.92 ; 
      RECT 0.54 52.016 15.084 52.92 ; 
      RECT 0 48.546 0.468 52.92 ; 
      RECT 37.836 48.546 38.448 52.208 ; 
      RECT 23.58 48.546 37.764 52.92 ; 
      RECT 20.592 48.546 23.508 52.208 ; 
      RECT 19.944 49.328 20.448 52.92 ; 
      RECT 14.94 48.944 19.836 52.208 ; 
      RECT 0.684 48.546 14.868 52.92 ; 
      RECT 0 48.546 0.612 52.208 ; 
      RECT 20.376 48.546 38.448 51.824 ; 
      RECT 0 48.944 20.304 51.824 ; 
      RECT 19.476 48.546 38.448 49.232 ; 
      RECT 0 48.546 19.404 51.824 ; 
      RECT 0 48.546 38.448 48.848 ; 
      RECT 0 56.72 38.448 57.24 ; 
      RECT 37.98 52.866 38.448 57.24 ; 
      RECT 23.364 56.336 37.908 57.24 ; 
      RECT 18.036 56.336 23.292 57.24 ; 
      RECT 15.156 52.866 17.676 57.24 ; 
      RECT 0.54 56.336 15.084 57.24 ; 
      RECT 0 52.866 0.468 57.24 ; 
      RECT 37.836 52.866 38.448 56.528 ; 
      RECT 23.58 52.866 37.764 57.24 ; 
      RECT 20.592 52.866 23.508 56.528 ; 
      RECT 19.944 53.648 20.448 57.24 ; 
      RECT 14.94 53.264 19.836 56.528 ; 
      RECT 0.684 52.866 14.868 57.24 ; 
      RECT 0 52.866 0.612 56.528 ; 
      RECT 20.376 52.866 38.448 56.144 ; 
      RECT 0 53.264 20.304 56.144 ; 
      RECT 19.476 52.866 38.448 53.552 ; 
      RECT 0 52.866 19.404 56.144 ; 
      RECT 0 52.866 38.448 53.168 ; 
      RECT 0 61.04 38.448 61.56 ; 
      RECT 37.98 57.186 38.448 61.56 ; 
      RECT 23.364 60.656 37.908 61.56 ; 
      RECT 18.036 60.656 23.292 61.56 ; 
      RECT 15.156 57.186 17.676 61.56 ; 
      RECT 0.54 60.656 15.084 61.56 ; 
      RECT 0 57.186 0.468 61.56 ; 
      RECT 37.836 57.186 38.448 60.848 ; 
      RECT 23.58 57.186 37.764 61.56 ; 
      RECT 20.592 57.186 23.508 60.848 ; 
      RECT 19.944 57.968 20.448 61.56 ; 
      RECT 14.94 57.584 19.836 60.848 ; 
      RECT 0.684 57.186 14.868 61.56 ; 
      RECT 0 57.186 0.612 60.848 ; 
      RECT 20.376 57.186 38.448 60.464 ; 
      RECT 0 57.584 20.304 60.464 ; 
      RECT 19.476 57.186 38.448 57.872 ; 
      RECT 0 57.186 19.404 60.464 ; 
      RECT 0 57.186 38.448 57.488 ; 
      RECT 0 65.36 38.448 65.88 ; 
      RECT 37.98 61.506 38.448 65.88 ; 
      RECT 23.364 64.976 37.908 65.88 ; 
      RECT 18.036 64.976 23.292 65.88 ; 
      RECT 15.156 61.506 17.676 65.88 ; 
      RECT 0.54 64.976 15.084 65.88 ; 
      RECT 0 61.506 0.468 65.88 ; 
      RECT 37.836 61.506 38.448 65.168 ; 
      RECT 23.58 61.506 37.764 65.88 ; 
      RECT 20.592 61.506 23.508 65.168 ; 
      RECT 19.944 62.288 20.448 65.88 ; 
      RECT 14.94 61.904 19.836 65.168 ; 
      RECT 0.684 61.506 14.868 65.88 ; 
      RECT 0 61.506 0.612 65.168 ; 
      RECT 20.376 61.506 38.448 64.784 ; 
      RECT 0 61.904 20.304 64.784 ; 
      RECT 19.476 61.506 38.448 62.192 ; 
      RECT 0 61.506 19.404 64.784 ; 
      RECT 0 61.506 38.448 61.808 ; 
      RECT 0 69.68 38.448 70.2 ; 
      RECT 37.98 65.826 38.448 70.2 ; 
      RECT 23.364 69.296 37.908 70.2 ; 
      RECT 18.036 69.296 23.292 70.2 ; 
      RECT 15.156 65.826 17.676 70.2 ; 
      RECT 0.54 69.296 15.084 70.2 ; 
      RECT 0 65.826 0.468 70.2 ; 
      RECT 37.836 65.826 38.448 69.488 ; 
      RECT 23.58 65.826 37.764 70.2 ; 
      RECT 20.592 65.826 23.508 69.488 ; 
      RECT 19.944 66.608 20.448 70.2 ; 
      RECT 14.94 66.224 19.836 69.488 ; 
      RECT 0.684 65.826 14.868 70.2 ; 
      RECT 0 65.826 0.612 69.488 ; 
      RECT 20.376 65.826 38.448 69.104 ; 
      RECT 0 66.224 20.304 69.104 ; 
      RECT 19.476 65.826 38.448 66.512 ; 
      RECT 0 65.826 19.404 69.104 ; 
      RECT 0 65.826 38.448 66.128 ; 
      RECT 0 74 38.448 74.52 ; 
      RECT 37.98 70.146 38.448 74.52 ; 
      RECT 23.364 73.616 37.908 74.52 ; 
      RECT 18.036 73.616 23.292 74.52 ; 
      RECT 15.156 70.146 17.676 74.52 ; 
      RECT 0.54 73.616 15.084 74.52 ; 
      RECT 0 70.146 0.468 74.52 ; 
      RECT 37.836 70.146 38.448 73.808 ; 
      RECT 23.58 70.146 37.764 74.52 ; 
      RECT 20.592 70.146 23.508 73.808 ; 
      RECT 19.944 70.928 20.448 74.52 ; 
      RECT 14.94 70.544 19.836 73.808 ; 
      RECT 0.684 70.146 14.868 74.52 ; 
      RECT 0 70.146 0.612 73.808 ; 
      RECT 20.376 70.146 38.448 73.424 ; 
      RECT 0 70.544 20.304 73.424 ; 
      RECT 19.476 70.146 38.448 70.832 ; 
      RECT 0 70.146 19.404 73.424 ; 
      RECT 0 70.146 38.448 70.448 ; 
      RECT 0 78.32 38.448 78.84 ; 
      RECT 37.98 74.466 38.448 78.84 ; 
      RECT 23.364 77.936 37.908 78.84 ; 
      RECT 18.036 77.936 23.292 78.84 ; 
      RECT 15.156 74.466 17.676 78.84 ; 
      RECT 0.54 77.936 15.084 78.84 ; 
      RECT 0 74.466 0.468 78.84 ; 
      RECT 37.836 74.466 38.448 78.128 ; 
      RECT 23.58 74.466 37.764 78.84 ; 
      RECT 20.592 74.466 23.508 78.128 ; 
      RECT 19.944 75.248 20.448 78.84 ; 
      RECT 14.94 74.864 19.836 78.128 ; 
      RECT 0.684 74.466 14.868 78.84 ; 
      RECT 0 74.466 0.612 78.128 ; 
      RECT 20.376 74.466 38.448 77.744 ; 
      RECT 0 74.864 20.304 77.744 ; 
      RECT 19.476 74.466 38.448 75.152 ; 
      RECT 0 74.466 19.404 77.744 ; 
      RECT 0 74.466 38.448 74.768 ; 
      RECT 0 82.64 38.448 83.16 ; 
      RECT 37.98 78.786 38.448 83.16 ; 
      RECT 23.364 82.256 37.908 83.16 ; 
      RECT 18.036 82.256 23.292 83.16 ; 
      RECT 15.156 78.786 17.676 83.16 ; 
      RECT 0.54 82.256 15.084 83.16 ; 
      RECT 0 78.786 0.468 83.16 ; 
      RECT 37.836 78.786 38.448 82.448 ; 
      RECT 23.58 78.786 37.764 83.16 ; 
      RECT 20.592 78.786 23.508 82.448 ; 
      RECT 19.944 79.568 20.448 83.16 ; 
      RECT 14.94 79.184 19.836 82.448 ; 
      RECT 0.684 78.786 14.868 83.16 ; 
      RECT 0 78.786 0.612 82.448 ; 
      RECT 20.376 78.786 38.448 82.064 ; 
      RECT 0 79.184 20.304 82.064 ; 
      RECT 19.476 78.786 38.448 79.472 ; 
      RECT 0 78.786 19.404 82.064 ; 
      RECT 0 78.786 38.448 79.088 ; 
      RECT 0 86.96 38.448 87.48 ; 
      RECT 37.98 83.106 38.448 87.48 ; 
      RECT 23.364 86.576 37.908 87.48 ; 
      RECT 18.036 86.576 23.292 87.48 ; 
      RECT 15.156 83.106 17.676 87.48 ; 
      RECT 0.54 86.576 15.084 87.48 ; 
      RECT 0 83.106 0.468 87.48 ; 
      RECT 37.836 83.106 38.448 86.768 ; 
      RECT 23.58 83.106 37.764 87.48 ; 
      RECT 20.592 83.106 23.508 86.768 ; 
      RECT 19.944 83.888 20.448 87.48 ; 
      RECT 14.94 83.504 19.836 86.768 ; 
      RECT 0.684 83.106 14.868 87.48 ; 
      RECT 0 83.106 0.612 86.768 ; 
      RECT 20.376 83.106 38.448 86.384 ; 
      RECT 0 83.504 20.304 86.384 ; 
      RECT 19.476 83.106 38.448 83.792 ; 
      RECT 0 83.106 19.404 86.384 ; 
      RECT 0 83.106 38.448 83.408 ; 
      RECT 0 91.28 38.448 91.8 ; 
      RECT 37.98 87.426 38.448 91.8 ; 
      RECT 23.364 90.896 37.908 91.8 ; 
      RECT 18.036 90.896 23.292 91.8 ; 
      RECT 15.156 87.426 17.676 91.8 ; 
      RECT 0.54 90.896 15.084 91.8 ; 
      RECT 0 87.426 0.468 91.8 ; 
      RECT 37.836 87.426 38.448 91.088 ; 
      RECT 23.58 87.426 37.764 91.8 ; 
      RECT 20.592 87.426 23.508 91.088 ; 
      RECT 19.944 88.208 20.448 91.8 ; 
      RECT 14.94 87.824 19.836 91.088 ; 
      RECT 0.684 87.426 14.868 91.8 ; 
      RECT 0 87.426 0.612 91.088 ; 
      RECT 20.376 87.426 38.448 90.704 ; 
      RECT 0 87.824 20.304 90.704 ; 
      RECT 19.476 87.426 38.448 88.112 ; 
      RECT 0 87.426 19.404 90.704 ; 
      RECT 0 87.426 38.448 87.728 ; 
      RECT 0 95.6 38.448 96.12 ; 
      RECT 37.98 91.746 38.448 96.12 ; 
      RECT 23.364 95.216 37.908 96.12 ; 
      RECT 18.036 95.216 23.292 96.12 ; 
      RECT 15.156 91.746 17.676 96.12 ; 
      RECT 0.54 95.216 15.084 96.12 ; 
      RECT 0 91.746 0.468 96.12 ; 
      RECT 37.836 91.746 38.448 95.408 ; 
      RECT 23.58 91.746 37.764 96.12 ; 
      RECT 20.592 91.746 23.508 95.408 ; 
      RECT 19.944 92.528 20.448 96.12 ; 
      RECT 14.94 92.144 19.836 95.408 ; 
      RECT 0.684 91.746 14.868 96.12 ; 
      RECT 0 91.746 0.612 95.408 ; 
      RECT 20.376 91.746 38.448 95.024 ; 
      RECT 0 92.144 20.304 95.024 ; 
      RECT 19.476 91.746 38.448 92.432 ; 
      RECT 0 91.746 19.404 95.024 ; 
      RECT 0 91.746 38.448 92.048 ; 
      RECT 0 99.92 38.448 100.44 ; 
      RECT 37.98 96.066 38.448 100.44 ; 
      RECT 23.364 99.536 37.908 100.44 ; 
      RECT 18.036 99.536 23.292 100.44 ; 
      RECT 15.156 96.066 17.676 100.44 ; 
      RECT 0.54 99.536 15.084 100.44 ; 
      RECT 0 96.066 0.468 100.44 ; 
      RECT 37.836 96.066 38.448 99.728 ; 
      RECT 23.58 96.066 37.764 100.44 ; 
      RECT 20.592 96.066 23.508 99.728 ; 
      RECT 19.944 96.848 20.448 100.44 ; 
      RECT 14.94 96.464 19.836 99.728 ; 
      RECT 0.684 96.066 14.868 100.44 ; 
      RECT 0 96.066 0.612 99.728 ; 
      RECT 20.376 96.066 38.448 99.344 ; 
      RECT 0 96.464 20.304 99.344 ; 
      RECT 19.476 96.066 38.448 96.752 ; 
      RECT 0 96.066 19.404 99.344 ; 
      RECT 0 96.066 38.448 96.368 ; 
      RECT 0 104.24 38.448 104.76 ; 
      RECT 37.98 100.386 38.448 104.76 ; 
      RECT 23.364 103.856 37.908 104.76 ; 
      RECT 18.036 103.856 23.292 104.76 ; 
      RECT 15.156 100.386 17.676 104.76 ; 
      RECT 0.54 103.856 15.084 104.76 ; 
      RECT 0 100.386 0.468 104.76 ; 
      RECT 37.836 100.386 38.448 104.048 ; 
      RECT 23.58 100.386 37.764 104.76 ; 
      RECT 20.592 100.386 23.508 104.048 ; 
      RECT 19.944 101.168 20.448 104.76 ; 
      RECT 14.94 100.784 19.836 104.048 ; 
      RECT 0.684 100.386 14.868 104.76 ; 
      RECT 0 100.386 0.612 104.048 ; 
      RECT 20.376 100.386 38.448 103.664 ; 
      RECT 0 100.784 20.304 103.664 ; 
      RECT 19.476 100.386 38.448 101.072 ; 
      RECT 0 100.386 19.404 103.664 ; 
      RECT 0 100.386 38.448 100.688 ; 
      RECT 0 108.56 38.448 109.08 ; 
      RECT 37.98 104.706 38.448 109.08 ; 
      RECT 23.364 108.176 37.908 109.08 ; 
      RECT 18.036 108.176 23.292 109.08 ; 
      RECT 15.156 104.706 17.676 109.08 ; 
      RECT 0.54 108.176 15.084 109.08 ; 
      RECT 0 104.706 0.468 109.08 ; 
      RECT 37.836 104.706 38.448 108.368 ; 
      RECT 23.58 104.706 37.764 109.08 ; 
      RECT 20.592 104.706 23.508 108.368 ; 
      RECT 19.944 105.488 20.448 109.08 ; 
      RECT 14.94 105.104 19.836 108.368 ; 
      RECT 0.684 104.706 14.868 109.08 ; 
      RECT 0 104.706 0.612 108.368 ; 
      RECT 20.376 104.706 38.448 107.984 ; 
      RECT 0 105.104 20.304 107.984 ; 
      RECT 19.476 104.706 38.448 105.392 ; 
      RECT 0 104.706 19.404 107.984 ; 
      RECT 0 104.706 38.448 105.008 ; 
      RECT 0 112.88 38.448 113.4 ; 
      RECT 37.98 109.026 38.448 113.4 ; 
      RECT 23.364 112.496 37.908 113.4 ; 
      RECT 18.036 112.496 23.292 113.4 ; 
      RECT 15.156 109.026 17.676 113.4 ; 
      RECT 0.54 112.496 15.084 113.4 ; 
      RECT 0 109.026 0.468 113.4 ; 
      RECT 37.836 109.026 38.448 112.688 ; 
      RECT 23.58 109.026 37.764 113.4 ; 
      RECT 20.592 109.026 23.508 112.688 ; 
      RECT 19.944 109.808 20.448 113.4 ; 
      RECT 14.94 109.424 19.836 112.688 ; 
      RECT 0.684 109.026 14.868 113.4 ; 
      RECT 0 109.026 0.612 112.688 ; 
      RECT 20.376 109.026 38.448 112.304 ; 
      RECT 0 109.424 20.304 112.304 ; 
      RECT 19.476 109.026 38.448 109.712 ; 
      RECT 0 109.026 19.404 112.304 ; 
      RECT 0 109.026 38.448 109.328 ; 
      RECT 0 117.2 38.448 117.72 ; 
      RECT 37.98 113.346 38.448 117.72 ; 
      RECT 23.364 116.816 37.908 117.72 ; 
      RECT 18.036 116.816 23.292 117.72 ; 
      RECT 15.156 113.346 17.676 117.72 ; 
      RECT 0.54 116.816 15.084 117.72 ; 
      RECT 0 113.346 0.468 117.72 ; 
      RECT 37.836 113.346 38.448 117.008 ; 
      RECT 23.58 113.346 37.764 117.72 ; 
      RECT 20.592 113.346 23.508 117.008 ; 
      RECT 19.944 114.128 20.448 117.72 ; 
      RECT 14.94 113.744 19.836 117.008 ; 
      RECT 0.684 113.346 14.868 117.72 ; 
      RECT 0 113.346 0.612 117.008 ; 
      RECT 20.376 113.346 38.448 116.624 ; 
      RECT 0 113.744 20.304 116.624 ; 
      RECT 19.476 113.346 38.448 114.032 ; 
      RECT 0 113.346 19.404 116.624 ; 
      RECT 0 113.346 38.448 113.648 ; 
      RECT 0 121.52 38.448 122.04 ; 
      RECT 37.98 117.666 38.448 122.04 ; 
      RECT 23.364 121.136 37.908 122.04 ; 
      RECT 18.036 121.136 23.292 122.04 ; 
      RECT 15.156 117.666 17.676 122.04 ; 
      RECT 0.54 121.136 15.084 122.04 ; 
      RECT 0 117.666 0.468 122.04 ; 
      RECT 37.836 117.666 38.448 121.328 ; 
      RECT 23.58 117.666 37.764 122.04 ; 
      RECT 20.592 117.666 23.508 121.328 ; 
      RECT 19.944 118.448 20.448 122.04 ; 
      RECT 14.94 118.064 19.836 121.328 ; 
      RECT 0.684 117.666 14.868 122.04 ; 
      RECT 0 117.666 0.612 121.328 ; 
      RECT 20.376 117.666 38.448 120.944 ; 
      RECT 0 118.064 20.304 120.944 ; 
      RECT 19.476 117.666 38.448 118.352 ; 
      RECT 0 117.666 19.404 120.944 ; 
      RECT 0 117.666 38.448 117.968 ; 
      RECT 0 125.84 38.448 126.36 ; 
      RECT 37.98 121.986 38.448 126.36 ; 
      RECT 23.364 125.456 37.908 126.36 ; 
      RECT 18.036 125.456 23.292 126.36 ; 
      RECT 15.156 121.986 17.676 126.36 ; 
      RECT 0.54 125.456 15.084 126.36 ; 
      RECT 0 121.986 0.468 126.36 ; 
      RECT 37.836 121.986 38.448 125.648 ; 
      RECT 23.58 121.986 37.764 126.36 ; 
      RECT 20.592 121.986 23.508 125.648 ; 
      RECT 19.944 122.768 20.448 126.36 ; 
      RECT 14.94 122.384 19.836 125.648 ; 
      RECT 0.684 121.986 14.868 126.36 ; 
      RECT 0 121.986 0.612 125.648 ; 
      RECT 20.376 121.986 38.448 125.264 ; 
      RECT 0 122.384 20.304 125.264 ; 
      RECT 19.476 121.986 38.448 122.672 ; 
      RECT 0 121.986 19.404 125.264 ; 
      RECT 0 121.986 38.448 122.288 ; 
      RECT 0 130.16 38.448 130.68 ; 
      RECT 37.98 126.306 38.448 130.68 ; 
      RECT 23.364 129.776 37.908 130.68 ; 
      RECT 18.036 129.776 23.292 130.68 ; 
      RECT 15.156 126.306 17.676 130.68 ; 
      RECT 0.54 129.776 15.084 130.68 ; 
      RECT 0 126.306 0.468 130.68 ; 
      RECT 37.836 126.306 38.448 129.968 ; 
      RECT 23.58 126.306 37.764 130.68 ; 
      RECT 20.592 126.306 23.508 129.968 ; 
      RECT 19.944 127.088 20.448 130.68 ; 
      RECT 14.94 126.704 19.836 129.968 ; 
      RECT 0.684 126.306 14.868 130.68 ; 
      RECT 0 126.306 0.612 129.968 ; 
      RECT 20.376 126.306 38.448 129.584 ; 
      RECT 0 126.704 20.304 129.584 ; 
      RECT 19.476 126.306 38.448 126.992 ; 
      RECT 0 126.306 19.404 129.584 ; 
      RECT 0 126.306 38.448 126.608 ; 
      RECT 0 134.48 38.448 135 ; 
      RECT 37.98 130.626 38.448 135 ; 
      RECT 23.364 134.096 37.908 135 ; 
      RECT 18.036 134.096 23.292 135 ; 
      RECT 15.156 130.626 17.676 135 ; 
      RECT 0.54 134.096 15.084 135 ; 
      RECT 0 130.626 0.468 135 ; 
      RECT 37.836 130.626 38.448 134.288 ; 
      RECT 23.58 130.626 37.764 135 ; 
      RECT 20.592 130.626 23.508 134.288 ; 
      RECT 19.944 131.408 20.448 135 ; 
      RECT 14.94 131.024 19.836 134.288 ; 
      RECT 0.684 130.626 14.868 135 ; 
      RECT 0 130.626 0.612 134.288 ; 
      RECT 20.376 130.626 38.448 133.904 ; 
      RECT 0 131.024 20.304 133.904 ; 
      RECT 19.476 130.626 38.448 131.312 ; 
      RECT 0 130.626 19.404 133.904 ; 
      RECT 0 130.626 38.448 130.928 ; 
      RECT 0 138.8 38.448 139.32 ; 
      RECT 37.98 134.946 38.448 139.32 ; 
      RECT 23.364 138.416 37.908 139.32 ; 
      RECT 18.036 138.416 23.292 139.32 ; 
      RECT 15.156 134.946 17.676 139.32 ; 
      RECT 0.54 138.416 15.084 139.32 ; 
      RECT 0 134.946 0.468 139.32 ; 
      RECT 37.836 134.946 38.448 138.608 ; 
      RECT 23.58 134.946 37.764 139.32 ; 
      RECT 20.592 134.946 23.508 138.608 ; 
      RECT 19.944 135.728 20.448 139.32 ; 
      RECT 14.94 135.344 19.836 138.608 ; 
      RECT 0.684 134.946 14.868 139.32 ; 
      RECT 0 134.946 0.612 138.608 ; 
      RECT 20.376 134.946 38.448 138.224 ; 
      RECT 0 135.344 20.304 138.224 ; 
      RECT 19.476 134.946 38.448 135.632 ; 
      RECT 0 134.946 19.404 138.224 ; 
      RECT 0 134.946 38.448 135.248 ; 
      RECT 0 143.12 38.448 143.64 ; 
      RECT 37.98 139.266 38.448 143.64 ; 
      RECT 23.364 142.736 37.908 143.64 ; 
      RECT 18.036 142.736 23.292 143.64 ; 
      RECT 15.156 139.266 17.676 143.64 ; 
      RECT 0.54 142.736 15.084 143.64 ; 
      RECT 0 139.266 0.468 143.64 ; 
      RECT 37.836 139.266 38.448 142.928 ; 
      RECT 23.58 139.266 37.764 143.64 ; 
      RECT 20.592 139.266 23.508 142.928 ; 
      RECT 19.944 140.048 20.448 143.64 ; 
      RECT 14.94 139.664 19.836 142.928 ; 
      RECT 0.684 139.266 14.868 143.64 ; 
      RECT 0 139.266 0.612 142.928 ; 
      RECT 20.376 139.266 38.448 142.544 ; 
      RECT 0 139.664 20.304 142.544 ; 
      RECT 19.476 139.266 38.448 139.952 ; 
      RECT 0 139.266 19.404 142.544 ; 
      RECT 0 139.266 38.448 139.568 ; 
      RECT 0 147.44 38.448 147.96 ; 
      RECT 37.98 143.586 38.448 147.96 ; 
      RECT 23.364 147.056 37.908 147.96 ; 
      RECT 18.036 147.056 23.292 147.96 ; 
      RECT 15.156 143.586 17.676 147.96 ; 
      RECT 0.54 147.056 15.084 147.96 ; 
      RECT 0 143.586 0.468 147.96 ; 
      RECT 37.836 143.586 38.448 147.248 ; 
      RECT 23.58 143.586 37.764 147.96 ; 
      RECT 20.592 143.586 23.508 147.248 ; 
      RECT 19.944 144.368 20.448 147.96 ; 
      RECT 14.94 143.984 19.836 147.248 ; 
      RECT 0.684 143.586 14.868 147.96 ; 
      RECT 0 143.586 0.612 147.248 ; 
      RECT 20.376 143.586 38.448 146.864 ; 
      RECT 0 143.984 20.304 146.864 ; 
      RECT 19.476 143.586 38.448 144.272 ; 
      RECT 0 143.586 19.404 146.864 ; 
      RECT 0 143.586 38.448 143.888 ; 
      RECT 0 151.76 38.448 152.28 ; 
      RECT 37.98 147.906 38.448 152.28 ; 
      RECT 23.364 151.376 37.908 152.28 ; 
      RECT 18.036 151.376 23.292 152.28 ; 
      RECT 15.156 147.906 17.676 152.28 ; 
      RECT 0.54 151.376 15.084 152.28 ; 
      RECT 0 147.906 0.468 152.28 ; 
      RECT 37.836 147.906 38.448 151.568 ; 
      RECT 23.58 147.906 37.764 152.28 ; 
      RECT 20.592 147.906 23.508 151.568 ; 
      RECT 19.944 148.688 20.448 152.28 ; 
      RECT 14.94 148.304 19.836 151.568 ; 
      RECT 0.684 147.906 14.868 152.28 ; 
      RECT 0 147.906 0.612 151.568 ; 
      RECT 20.376 147.906 38.448 151.184 ; 
      RECT 0 148.304 20.304 151.184 ; 
      RECT 19.476 147.906 38.448 148.592 ; 
      RECT 0 147.906 19.404 151.184 ; 
      RECT 0 147.906 38.448 148.208 ; 
      RECT 0 156.08 38.448 156.6 ; 
      RECT 37.98 152.226 38.448 156.6 ; 
      RECT 23.364 155.696 37.908 156.6 ; 
      RECT 18.036 155.696 23.292 156.6 ; 
      RECT 15.156 152.226 17.676 156.6 ; 
      RECT 0.54 155.696 15.084 156.6 ; 
      RECT 0 152.226 0.468 156.6 ; 
      RECT 37.836 152.226 38.448 155.888 ; 
      RECT 23.58 152.226 37.764 156.6 ; 
      RECT 20.592 152.226 23.508 155.888 ; 
      RECT 19.944 153.008 20.448 156.6 ; 
      RECT 14.94 152.624 19.836 155.888 ; 
      RECT 0.684 152.226 14.868 156.6 ; 
      RECT 0 152.226 0.612 155.888 ; 
      RECT 20.376 152.226 38.448 155.504 ; 
      RECT 0 152.624 20.304 155.504 ; 
      RECT 19.476 152.226 38.448 152.912 ; 
      RECT 0 152.226 19.404 155.504 ; 
      RECT 0 152.226 38.448 152.528 ; 
      RECT 0 160.4 38.448 160.92 ; 
      RECT 37.98 156.546 38.448 160.92 ; 
      RECT 23.364 160.016 37.908 160.92 ; 
      RECT 18.036 160.016 23.292 160.92 ; 
      RECT 15.156 156.546 17.676 160.92 ; 
      RECT 0.54 160.016 15.084 160.92 ; 
      RECT 0 156.546 0.468 160.92 ; 
      RECT 37.836 156.546 38.448 160.208 ; 
      RECT 23.58 156.546 37.764 160.92 ; 
      RECT 20.592 156.546 23.508 160.208 ; 
      RECT 19.944 157.328 20.448 160.92 ; 
      RECT 14.94 156.944 19.836 160.208 ; 
      RECT 0.684 156.546 14.868 160.92 ; 
      RECT 0 156.546 0.612 160.208 ; 
      RECT 20.376 156.546 38.448 159.824 ; 
      RECT 0 156.944 20.304 159.824 ; 
      RECT 19.476 156.546 38.448 157.232 ; 
      RECT 0 156.546 19.404 159.824 ; 
      RECT 0 156.546 38.448 156.848 ; 
      RECT 0 164.72 38.448 165.24 ; 
      RECT 37.98 160.866 38.448 165.24 ; 
      RECT 23.364 164.336 37.908 165.24 ; 
      RECT 18.036 164.336 23.292 165.24 ; 
      RECT 15.156 160.866 17.676 165.24 ; 
      RECT 0.54 164.336 15.084 165.24 ; 
      RECT 0 160.866 0.468 165.24 ; 
      RECT 37.836 160.866 38.448 164.528 ; 
      RECT 23.58 160.866 37.764 165.24 ; 
      RECT 20.592 160.866 23.508 164.528 ; 
      RECT 19.944 161.648 20.448 165.24 ; 
      RECT 14.94 161.264 19.836 164.528 ; 
      RECT 0.684 160.866 14.868 165.24 ; 
      RECT 0 160.866 0.612 164.528 ; 
      RECT 20.376 160.866 38.448 164.144 ; 
      RECT 0 161.264 20.304 164.144 ; 
      RECT 19.476 160.866 38.448 161.552 ; 
      RECT 0 160.866 19.404 164.144 ; 
      RECT 0 160.866 38.448 161.168 ; 
      RECT 0 169.04 38.448 169.56 ; 
      RECT 37.98 165.186 38.448 169.56 ; 
      RECT 23.364 168.656 37.908 169.56 ; 
      RECT 18.036 168.656 23.292 169.56 ; 
      RECT 15.156 165.186 17.676 169.56 ; 
      RECT 0.54 168.656 15.084 169.56 ; 
      RECT 0 165.186 0.468 169.56 ; 
      RECT 37.836 165.186 38.448 168.848 ; 
      RECT 23.58 165.186 37.764 169.56 ; 
      RECT 20.592 165.186 23.508 168.848 ; 
      RECT 19.944 165.968 20.448 169.56 ; 
      RECT 14.94 165.584 19.836 168.848 ; 
      RECT 0.684 165.186 14.868 169.56 ; 
      RECT 0 165.186 0.612 168.848 ; 
      RECT 20.376 165.186 38.448 168.464 ; 
      RECT 0 165.584 20.304 168.464 ; 
      RECT 19.476 165.186 38.448 165.872 ; 
      RECT 0 165.186 19.404 168.464 ; 
      RECT 0 165.186 38.448 165.488 ; 
      RECT 0 173.36 38.448 173.88 ; 
      RECT 37.98 169.506 38.448 173.88 ; 
      RECT 23.364 172.976 37.908 173.88 ; 
      RECT 18.036 172.976 23.292 173.88 ; 
      RECT 15.156 169.506 17.676 173.88 ; 
      RECT 0.54 172.976 15.084 173.88 ; 
      RECT 0 169.506 0.468 173.88 ; 
      RECT 37.836 169.506 38.448 173.168 ; 
      RECT 23.58 169.506 37.764 173.88 ; 
      RECT 20.592 169.506 23.508 173.168 ; 
      RECT 19.944 170.288 20.448 173.88 ; 
      RECT 14.94 169.904 19.836 173.168 ; 
      RECT 0.684 169.506 14.868 173.88 ; 
      RECT 0 169.506 0.612 173.168 ; 
      RECT 20.376 169.506 38.448 172.784 ; 
      RECT 0 169.904 20.304 172.784 ; 
      RECT 19.476 169.506 38.448 170.192 ; 
      RECT 0 169.506 19.404 172.784 ; 
      RECT 0 169.506 38.448 169.808 ; 
      RECT 0 203.052 38.448 208.386 ; 
      RECT 29.412 173.772 38.448 208.386 ; 
      RECT 20.612 189.228 38.448 208.386 ; 
      RECT 24.228 178.86 38.448 208.386 ; 
      RECT 20.404 173.772 20.54 208.386 ; 
      RECT 20.196 173.772 20.332 208.386 ; 
      RECT 19.988 173.772 20.124 208.386 ; 
      RECT 19.78 173.772 19.916 208.386 ; 
      RECT 0 201.324 19.708 208.386 ; 
      RECT 18.74 190.38 38.448 202.188 ; 
      RECT 18.532 173.772 18.668 208.386 ; 
      RECT 18.324 173.772 18.46 208.386 ; 
      RECT 18.116 173.772 18.252 208.386 ; 
      RECT 17.908 173.772 18.044 208.386 ; 
      RECT 0 180.012 17.836 208.386 ; 
      RECT 0 188.652 19.708 200.46 ; 
      RECT 18.74 177.708 23.292 189.516 ; 
      RECT 23.364 179.628 38.448 208.386 ; 
      RECT 20.772 174.092 24.156 189.132 ; 
      RECT 16.02 175.98 19.116 187.788 ; 
      RECT 15.156 176.556 17.836 208.386 ; 
      RECT 0 178.86 15.084 208.386 ; 
      RECT 13.428 173.772 15.228 179.916 ; 
      RECT 28.548 173.772 29.34 208.386 ; 
      RECT 13.428 178.092 28.476 179.532 ; 
      RECT 9.972 176.556 13.356 208.386 ; 
      RECT 0 177.708 9.9 208.386 ; 
      RECT 27.684 173.772 38.448 178.764 ; 
      RECT 26.82 176.556 38.448 178.764 ; 
      RECT 0 177.708 26.748 178.764 ; 
      RECT 25.956 173.772 27.612 177.996 ; 
      RECT 20.612 176.556 38.448 177.996 ; 
      RECT 0.684 176.556 19.708 178.764 ; 
      RECT 18.74 176.364 19.708 208.386 ; 
      RECT 0 175.98 0.612 208.386 ; 
      RECT 19.188 173.772 20.7 176.844 ; 
      RECT 20.772 176.364 25.884 179.532 ; 
      RECT 12.564 176.364 15.948 178.764 ; 
      RECT 10.836 176.364 12.492 208.386 ; 
      RECT 0 175.98 10.764 176.844 ; 
      RECT 25.092 173.772 38.448 176.46 ; 
      RECT 19.188 174.092 25.02 176.46 ; 
      RECT 15.3 175.98 19.116 176.46 ; 
      RECT 11.7 173.772 15.228 176.46 ; 
      RECT 0 175.98 11.628 176.46 ; 
      RECT 23.364 173.772 38.448 176.268 ; 
      RECT 18.74 174.092 38.448 176.268 ; 
      RECT 0.54 173.772 17.836 176.268 ; 
      RECT 0 173.772 0.468 208.386 ; 
      RECT 0 173.772 23.292 175.116 ; 
      RECT 0 173.772 38.448 173.996 ; 
        RECT 0 210.188 38.448 210.708 ; 
        RECT 37.98 206.334 38.448 210.708 ; 
        RECT 23.364 209.804 37.908 210.708 ; 
        RECT 18.036 209.804 23.292 210.708 ; 
        RECT 15.156 206.334 17.676 210.708 ; 
        RECT 0.54 209.804 15.084 210.708 ; 
        RECT 0 206.334 0.468 210.708 ; 
        RECT 37.836 206.334 38.448 209.996 ; 
        RECT 23.58 206.334 37.764 210.708 ; 
        RECT 20.592 206.334 23.508 209.996 ; 
        RECT 19.944 207.116 20.448 210.708 ; 
        RECT 14.94 206.732 19.836 209.996 ; 
        RECT 0.684 206.334 14.868 210.708 ; 
        RECT 0 206.334 0.612 209.996 ; 
        RECT 20.376 206.334 38.448 209.612 ; 
        RECT 0 206.732 20.304 209.612 ; 
        RECT 19.476 206.334 38.448 207.02 ; 
        RECT 0 206.334 19.404 209.612 ; 
        RECT 0 206.334 38.448 206.636 ; 
        RECT 0 214.508 38.448 215.028 ; 
        RECT 37.98 210.654 38.448 215.028 ; 
        RECT 23.364 214.124 37.908 215.028 ; 
        RECT 18.036 214.124 23.292 215.028 ; 
        RECT 15.156 210.654 17.676 215.028 ; 
        RECT 0.54 214.124 15.084 215.028 ; 
        RECT 0 210.654 0.468 215.028 ; 
        RECT 37.836 210.654 38.448 214.316 ; 
        RECT 23.58 210.654 37.764 215.028 ; 
        RECT 20.592 210.654 23.508 214.316 ; 
        RECT 19.944 211.436 20.448 215.028 ; 
        RECT 14.94 211.052 19.836 214.316 ; 
        RECT 0.684 210.654 14.868 215.028 ; 
        RECT 0 210.654 0.612 214.316 ; 
        RECT 20.376 210.654 38.448 213.932 ; 
        RECT 0 211.052 20.304 213.932 ; 
        RECT 19.476 210.654 38.448 211.34 ; 
        RECT 0 210.654 19.404 213.932 ; 
        RECT 0 210.654 38.448 210.956 ; 
        RECT 0 218.828 38.448 219.348 ; 
        RECT 37.98 214.974 38.448 219.348 ; 
        RECT 23.364 218.444 37.908 219.348 ; 
        RECT 18.036 218.444 23.292 219.348 ; 
        RECT 15.156 214.974 17.676 219.348 ; 
        RECT 0.54 218.444 15.084 219.348 ; 
        RECT 0 214.974 0.468 219.348 ; 
        RECT 37.836 214.974 38.448 218.636 ; 
        RECT 23.58 214.974 37.764 219.348 ; 
        RECT 20.592 214.974 23.508 218.636 ; 
        RECT 19.944 215.756 20.448 219.348 ; 
        RECT 14.94 215.372 19.836 218.636 ; 
        RECT 0.684 214.974 14.868 219.348 ; 
        RECT 0 214.974 0.612 218.636 ; 
        RECT 20.376 214.974 38.448 218.252 ; 
        RECT 0 215.372 20.304 218.252 ; 
        RECT 19.476 214.974 38.448 215.66 ; 
        RECT 0 214.974 19.404 218.252 ; 
        RECT 0 214.974 38.448 215.276 ; 
        RECT 0 223.148 38.448 223.668 ; 
        RECT 37.98 219.294 38.448 223.668 ; 
        RECT 23.364 222.764 37.908 223.668 ; 
        RECT 18.036 222.764 23.292 223.668 ; 
        RECT 15.156 219.294 17.676 223.668 ; 
        RECT 0.54 222.764 15.084 223.668 ; 
        RECT 0 219.294 0.468 223.668 ; 
        RECT 37.836 219.294 38.448 222.956 ; 
        RECT 23.58 219.294 37.764 223.668 ; 
        RECT 20.592 219.294 23.508 222.956 ; 
        RECT 19.944 220.076 20.448 223.668 ; 
        RECT 14.94 219.692 19.836 222.956 ; 
        RECT 0.684 219.294 14.868 223.668 ; 
        RECT 0 219.294 0.612 222.956 ; 
        RECT 20.376 219.294 38.448 222.572 ; 
        RECT 0 219.692 20.304 222.572 ; 
        RECT 19.476 219.294 38.448 219.98 ; 
        RECT 0 219.294 19.404 222.572 ; 
        RECT 0 219.294 38.448 219.596 ; 
        RECT 0 227.468 38.448 227.988 ; 
        RECT 37.98 223.614 38.448 227.988 ; 
        RECT 23.364 227.084 37.908 227.988 ; 
        RECT 18.036 227.084 23.292 227.988 ; 
        RECT 15.156 223.614 17.676 227.988 ; 
        RECT 0.54 227.084 15.084 227.988 ; 
        RECT 0 223.614 0.468 227.988 ; 
        RECT 37.836 223.614 38.448 227.276 ; 
        RECT 23.58 223.614 37.764 227.988 ; 
        RECT 20.592 223.614 23.508 227.276 ; 
        RECT 19.944 224.396 20.448 227.988 ; 
        RECT 14.94 224.012 19.836 227.276 ; 
        RECT 0.684 223.614 14.868 227.988 ; 
        RECT 0 223.614 0.612 227.276 ; 
        RECT 20.376 223.614 38.448 226.892 ; 
        RECT 0 224.012 20.304 226.892 ; 
        RECT 19.476 223.614 38.448 224.3 ; 
        RECT 0 223.614 19.404 226.892 ; 
        RECT 0 223.614 38.448 223.916 ; 
        RECT 0 231.788 38.448 232.308 ; 
        RECT 37.98 227.934 38.448 232.308 ; 
        RECT 23.364 231.404 37.908 232.308 ; 
        RECT 18.036 231.404 23.292 232.308 ; 
        RECT 15.156 227.934 17.676 232.308 ; 
        RECT 0.54 231.404 15.084 232.308 ; 
        RECT 0 227.934 0.468 232.308 ; 
        RECT 37.836 227.934 38.448 231.596 ; 
        RECT 23.58 227.934 37.764 232.308 ; 
        RECT 20.592 227.934 23.508 231.596 ; 
        RECT 19.944 228.716 20.448 232.308 ; 
        RECT 14.94 228.332 19.836 231.596 ; 
        RECT 0.684 227.934 14.868 232.308 ; 
        RECT 0 227.934 0.612 231.596 ; 
        RECT 20.376 227.934 38.448 231.212 ; 
        RECT 0 228.332 20.304 231.212 ; 
        RECT 19.476 227.934 38.448 228.62 ; 
        RECT 0 227.934 19.404 231.212 ; 
        RECT 0 227.934 38.448 228.236 ; 
        RECT 0 236.108 38.448 236.628 ; 
        RECT 37.98 232.254 38.448 236.628 ; 
        RECT 23.364 235.724 37.908 236.628 ; 
        RECT 18.036 235.724 23.292 236.628 ; 
        RECT 15.156 232.254 17.676 236.628 ; 
        RECT 0.54 235.724 15.084 236.628 ; 
        RECT 0 232.254 0.468 236.628 ; 
        RECT 37.836 232.254 38.448 235.916 ; 
        RECT 23.58 232.254 37.764 236.628 ; 
        RECT 20.592 232.254 23.508 235.916 ; 
        RECT 19.944 233.036 20.448 236.628 ; 
        RECT 14.94 232.652 19.836 235.916 ; 
        RECT 0.684 232.254 14.868 236.628 ; 
        RECT 0 232.254 0.612 235.916 ; 
        RECT 20.376 232.254 38.448 235.532 ; 
        RECT 0 232.652 20.304 235.532 ; 
        RECT 19.476 232.254 38.448 232.94 ; 
        RECT 0 232.254 19.404 235.532 ; 
        RECT 0 232.254 38.448 232.556 ; 
        RECT 0 240.428 38.448 240.948 ; 
        RECT 37.98 236.574 38.448 240.948 ; 
        RECT 23.364 240.044 37.908 240.948 ; 
        RECT 18.036 240.044 23.292 240.948 ; 
        RECT 15.156 236.574 17.676 240.948 ; 
        RECT 0.54 240.044 15.084 240.948 ; 
        RECT 0 236.574 0.468 240.948 ; 
        RECT 37.836 236.574 38.448 240.236 ; 
        RECT 23.58 236.574 37.764 240.948 ; 
        RECT 20.592 236.574 23.508 240.236 ; 
        RECT 19.944 237.356 20.448 240.948 ; 
        RECT 14.94 236.972 19.836 240.236 ; 
        RECT 0.684 236.574 14.868 240.948 ; 
        RECT 0 236.574 0.612 240.236 ; 
        RECT 20.376 236.574 38.448 239.852 ; 
        RECT 0 236.972 20.304 239.852 ; 
        RECT 19.476 236.574 38.448 237.26 ; 
        RECT 0 236.574 19.404 239.852 ; 
        RECT 0 236.574 38.448 236.876 ; 
        RECT 0 244.748 38.448 245.268 ; 
        RECT 37.98 240.894 38.448 245.268 ; 
        RECT 23.364 244.364 37.908 245.268 ; 
        RECT 18.036 244.364 23.292 245.268 ; 
        RECT 15.156 240.894 17.676 245.268 ; 
        RECT 0.54 244.364 15.084 245.268 ; 
        RECT 0 240.894 0.468 245.268 ; 
        RECT 37.836 240.894 38.448 244.556 ; 
        RECT 23.58 240.894 37.764 245.268 ; 
        RECT 20.592 240.894 23.508 244.556 ; 
        RECT 19.944 241.676 20.448 245.268 ; 
        RECT 14.94 241.292 19.836 244.556 ; 
        RECT 0.684 240.894 14.868 245.268 ; 
        RECT 0 240.894 0.612 244.556 ; 
        RECT 20.376 240.894 38.448 244.172 ; 
        RECT 0 241.292 20.304 244.172 ; 
        RECT 19.476 240.894 38.448 241.58 ; 
        RECT 0 240.894 19.404 244.172 ; 
        RECT 0 240.894 38.448 241.196 ; 
        RECT 0 249.068 38.448 249.588 ; 
        RECT 37.98 245.214 38.448 249.588 ; 
        RECT 23.364 248.684 37.908 249.588 ; 
        RECT 18.036 248.684 23.292 249.588 ; 
        RECT 15.156 245.214 17.676 249.588 ; 
        RECT 0.54 248.684 15.084 249.588 ; 
        RECT 0 245.214 0.468 249.588 ; 
        RECT 37.836 245.214 38.448 248.876 ; 
        RECT 23.58 245.214 37.764 249.588 ; 
        RECT 20.592 245.214 23.508 248.876 ; 
        RECT 19.944 245.996 20.448 249.588 ; 
        RECT 14.94 245.612 19.836 248.876 ; 
        RECT 0.684 245.214 14.868 249.588 ; 
        RECT 0 245.214 0.612 248.876 ; 
        RECT 20.376 245.214 38.448 248.492 ; 
        RECT 0 245.612 20.304 248.492 ; 
        RECT 19.476 245.214 38.448 245.9 ; 
        RECT 0 245.214 19.404 248.492 ; 
        RECT 0 245.214 38.448 245.516 ; 
        RECT 0 253.388 38.448 253.908 ; 
        RECT 37.98 249.534 38.448 253.908 ; 
        RECT 23.364 253.004 37.908 253.908 ; 
        RECT 18.036 253.004 23.292 253.908 ; 
        RECT 15.156 249.534 17.676 253.908 ; 
        RECT 0.54 253.004 15.084 253.908 ; 
        RECT 0 249.534 0.468 253.908 ; 
        RECT 37.836 249.534 38.448 253.196 ; 
        RECT 23.58 249.534 37.764 253.908 ; 
        RECT 20.592 249.534 23.508 253.196 ; 
        RECT 19.944 250.316 20.448 253.908 ; 
        RECT 14.94 249.932 19.836 253.196 ; 
        RECT 0.684 249.534 14.868 253.908 ; 
        RECT 0 249.534 0.612 253.196 ; 
        RECT 20.376 249.534 38.448 252.812 ; 
        RECT 0 249.932 20.304 252.812 ; 
        RECT 19.476 249.534 38.448 250.22 ; 
        RECT 0 249.534 19.404 252.812 ; 
        RECT 0 249.534 38.448 249.836 ; 
        RECT 0 257.708 38.448 258.228 ; 
        RECT 37.98 253.854 38.448 258.228 ; 
        RECT 23.364 257.324 37.908 258.228 ; 
        RECT 18.036 257.324 23.292 258.228 ; 
        RECT 15.156 253.854 17.676 258.228 ; 
        RECT 0.54 257.324 15.084 258.228 ; 
        RECT 0 253.854 0.468 258.228 ; 
        RECT 37.836 253.854 38.448 257.516 ; 
        RECT 23.58 253.854 37.764 258.228 ; 
        RECT 20.592 253.854 23.508 257.516 ; 
        RECT 19.944 254.636 20.448 258.228 ; 
        RECT 14.94 254.252 19.836 257.516 ; 
        RECT 0.684 253.854 14.868 258.228 ; 
        RECT 0 253.854 0.612 257.516 ; 
        RECT 20.376 253.854 38.448 257.132 ; 
        RECT 0 254.252 20.304 257.132 ; 
        RECT 19.476 253.854 38.448 254.54 ; 
        RECT 0 253.854 19.404 257.132 ; 
        RECT 0 253.854 38.448 254.156 ; 
        RECT 0 262.028 38.448 262.548 ; 
        RECT 37.98 258.174 38.448 262.548 ; 
        RECT 23.364 261.644 37.908 262.548 ; 
        RECT 18.036 261.644 23.292 262.548 ; 
        RECT 15.156 258.174 17.676 262.548 ; 
        RECT 0.54 261.644 15.084 262.548 ; 
        RECT 0 258.174 0.468 262.548 ; 
        RECT 37.836 258.174 38.448 261.836 ; 
        RECT 23.58 258.174 37.764 262.548 ; 
        RECT 20.592 258.174 23.508 261.836 ; 
        RECT 19.944 258.956 20.448 262.548 ; 
        RECT 14.94 258.572 19.836 261.836 ; 
        RECT 0.684 258.174 14.868 262.548 ; 
        RECT 0 258.174 0.612 261.836 ; 
        RECT 20.376 258.174 38.448 261.452 ; 
        RECT 0 258.572 20.304 261.452 ; 
        RECT 19.476 258.174 38.448 258.86 ; 
        RECT 0 258.174 19.404 261.452 ; 
        RECT 0 258.174 38.448 258.476 ; 
        RECT 0 266.348 38.448 266.868 ; 
        RECT 37.98 262.494 38.448 266.868 ; 
        RECT 23.364 265.964 37.908 266.868 ; 
        RECT 18.036 265.964 23.292 266.868 ; 
        RECT 15.156 262.494 17.676 266.868 ; 
        RECT 0.54 265.964 15.084 266.868 ; 
        RECT 0 262.494 0.468 266.868 ; 
        RECT 37.836 262.494 38.448 266.156 ; 
        RECT 23.58 262.494 37.764 266.868 ; 
        RECT 20.592 262.494 23.508 266.156 ; 
        RECT 19.944 263.276 20.448 266.868 ; 
        RECT 14.94 262.892 19.836 266.156 ; 
        RECT 0.684 262.494 14.868 266.868 ; 
        RECT 0 262.494 0.612 266.156 ; 
        RECT 20.376 262.494 38.448 265.772 ; 
        RECT 0 262.892 20.304 265.772 ; 
        RECT 19.476 262.494 38.448 263.18 ; 
        RECT 0 262.494 19.404 265.772 ; 
        RECT 0 262.494 38.448 262.796 ; 
        RECT 0 270.668 38.448 271.188 ; 
        RECT 37.98 266.814 38.448 271.188 ; 
        RECT 23.364 270.284 37.908 271.188 ; 
        RECT 18.036 270.284 23.292 271.188 ; 
        RECT 15.156 266.814 17.676 271.188 ; 
        RECT 0.54 270.284 15.084 271.188 ; 
        RECT 0 266.814 0.468 271.188 ; 
        RECT 37.836 266.814 38.448 270.476 ; 
        RECT 23.58 266.814 37.764 271.188 ; 
        RECT 20.592 266.814 23.508 270.476 ; 
        RECT 19.944 267.596 20.448 271.188 ; 
        RECT 14.94 267.212 19.836 270.476 ; 
        RECT 0.684 266.814 14.868 271.188 ; 
        RECT 0 266.814 0.612 270.476 ; 
        RECT 20.376 266.814 38.448 270.092 ; 
        RECT 0 267.212 20.304 270.092 ; 
        RECT 19.476 266.814 38.448 267.5 ; 
        RECT 0 266.814 19.404 270.092 ; 
        RECT 0 266.814 38.448 267.116 ; 
        RECT 0 274.988 38.448 275.508 ; 
        RECT 37.98 271.134 38.448 275.508 ; 
        RECT 23.364 274.604 37.908 275.508 ; 
        RECT 18.036 274.604 23.292 275.508 ; 
        RECT 15.156 271.134 17.676 275.508 ; 
        RECT 0.54 274.604 15.084 275.508 ; 
        RECT 0 271.134 0.468 275.508 ; 
        RECT 37.836 271.134 38.448 274.796 ; 
        RECT 23.58 271.134 37.764 275.508 ; 
        RECT 20.592 271.134 23.508 274.796 ; 
        RECT 19.944 271.916 20.448 275.508 ; 
        RECT 14.94 271.532 19.836 274.796 ; 
        RECT 0.684 271.134 14.868 275.508 ; 
        RECT 0 271.134 0.612 274.796 ; 
        RECT 20.376 271.134 38.448 274.412 ; 
        RECT 0 271.532 20.304 274.412 ; 
        RECT 19.476 271.134 38.448 271.82 ; 
        RECT 0 271.134 19.404 274.412 ; 
        RECT 0 271.134 38.448 271.436 ; 
        RECT 0 279.308 38.448 279.828 ; 
        RECT 37.98 275.454 38.448 279.828 ; 
        RECT 23.364 278.924 37.908 279.828 ; 
        RECT 18.036 278.924 23.292 279.828 ; 
        RECT 15.156 275.454 17.676 279.828 ; 
        RECT 0.54 278.924 15.084 279.828 ; 
        RECT 0 275.454 0.468 279.828 ; 
        RECT 37.836 275.454 38.448 279.116 ; 
        RECT 23.58 275.454 37.764 279.828 ; 
        RECT 20.592 275.454 23.508 279.116 ; 
        RECT 19.944 276.236 20.448 279.828 ; 
        RECT 14.94 275.852 19.836 279.116 ; 
        RECT 0.684 275.454 14.868 279.828 ; 
        RECT 0 275.454 0.612 279.116 ; 
        RECT 20.376 275.454 38.448 278.732 ; 
        RECT 0 275.852 20.304 278.732 ; 
        RECT 19.476 275.454 38.448 276.14 ; 
        RECT 0 275.454 19.404 278.732 ; 
        RECT 0 275.454 38.448 275.756 ; 
        RECT 0 283.628 38.448 284.148 ; 
        RECT 37.98 279.774 38.448 284.148 ; 
        RECT 23.364 283.244 37.908 284.148 ; 
        RECT 18.036 283.244 23.292 284.148 ; 
        RECT 15.156 279.774 17.676 284.148 ; 
        RECT 0.54 283.244 15.084 284.148 ; 
        RECT 0 279.774 0.468 284.148 ; 
        RECT 37.836 279.774 38.448 283.436 ; 
        RECT 23.58 279.774 37.764 284.148 ; 
        RECT 20.592 279.774 23.508 283.436 ; 
        RECT 19.944 280.556 20.448 284.148 ; 
        RECT 14.94 280.172 19.836 283.436 ; 
        RECT 0.684 279.774 14.868 284.148 ; 
        RECT 0 279.774 0.612 283.436 ; 
        RECT 20.376 279.774 38.448 283.052 ; 
        RECT 0 280.172 20.304 283.052 ; 
        RECT 19.476 279.774 38.448 280.46 ; 
        RECT 0 279.774 19.404 283.052 ; 
        RECT 0 279.774 38.448 280.076 ; 
        RECT 0 287.948 38.448 288.468 ; 
        RECT 37.98 284.094 38.448 288.468 ; 
        RECT 23.364 287.564 37.908 288.468 ; 
        RECT 18.036 287.564 23.292 288.468 ; 
        RECT 15.156 284.094 17.676 288.468 ; 
        RECT 0.54 287.564 15.084 288.468 ; 
        RECT 0 284.094 0.468 288.468 ; 
        RECT 37.836 284.094 38.448 287.756 ; 
        RECT 23.58 284.094 37.764 288.468 ; 
        RECT 20.592 284.094 23.508 287.756 ; 
        RECT 19.944 284.876 20.448 288.468 ; 
        RECT 14.94 284.492 19.836 287.756 ; 
        RECT 0.684 284.094 14.868 288.468 ; 
        RECT 0 284.094 0.612 287.756 ; 
        RECT 20.376 284.094 38.448 287.372 ; 
        RECT 0 284.492 20.304 287.372 ; 
        RECT 19.476 284.094 38.448 284.78 ; 
        RECT 0 284.094 19.404 287.372 ; 
        RECT 0 284.094 38.448 284.396 ; 
        RECT 0 292.268 38.448 292.788 ; 
        RECT 37.98 288.414 38.448 292.788 ; 
        RECT 23.364 291.884 37.908 292.788 ; 
        RECT 18.036 291.884 23.292 292.788 ; 
        RECT 15.156 288.414 17.676 292.788 ; 
        RECT 0.54 291.884 15.084 292.788 ; 
        RECT 0 288.414 0.468 292.788 ; 
        RECT 37.836 288.414 38.448 292.076 ; 
        RECT 23.58 288.414 37.764 292.788 ; 
        RECT 20.592 288.414 23.508 292.076 ; 
        RECT 19.944 289.196 20.448 292.788 ; 
        RECT 14.94 288.812 19.836 292.076 ; 
        RECT 0.684 288.414 14.868 292.788 ; 
        RECT 0 288.414 0.612 292.076 ; 
        RECT 20.376 288.414 38.448 291.692 ; 
        RECT 0 288.812 20.304 291.692 ; 
        RECT 19.476 288.414 38.448 289.1 ; 
        RECT 0 288.414 19.404 291.692 ; 
        RECT 0 288.414 38.448 288.716 ; 
        RECT 0 296.588 38.448 297.108 ; 
        RECT 37.98 292.734 38.448 297.108 ; 
        RECT 23.364 296.204 37.908 297.108 ; 
        RECT 18.036 296.204 23.292 297.108 ; 
        RECT 15.156 292.734 17.676 297.108 ; 
        RECT 0.54 296.204 15.084 297.108 ; 
        RECT 0 292.734 0.468 297.108 ; 
        RECT 37.836 292.734 38.448 296.396 ; 
        RECT 23.58 292.734 37.764 297.108 ; 
        RECT 20.592 292.734 23.508 296.396 ; 
        RECT 19.944 293.516 20.448 297.108 ; 
        RECT 14.94 293.132 19.836 296.396 ; 
        RECT 0.684 292.734 14.868 297.108 ; 
        RECT 0 292.734 0.612 296.396 ; 
        RECT 20.376 292.734 38.448 296.012 ; 
        RECT 0 293.132 20.304 296.012 ; 
        RECT 19.476 292.734 38.448 293.42 ; 
        RECT 0 292.734 19.404 296.012 ; 
        RECT 0 292.734 38.448 293.036 ; 
        RECT 0 300.908 38.448 301.428 ; 
        RECT 37.98 297.054 38.448 301.428 ; 
        RECT 23.364 300.524 37.908 301.428 ; 
        RECT 18.036 300.524 23.292 301.428 ; 
        RECT 15.156 297.054 17.676 301.428 ; 
        RECT 0.54 300.524 15.084 301.428 ; 
        RECT 0 297.054 0.468 301.428 ; 
        RECT 37.836 297.054 38.448 300.716 ; 
        RECT 23.58 297.054 37.764 301.428 ; 
        RECT 20.592 297.054 23.508 300.716 ; 
        RECT 19.944 297.836 20.448 301.428 ; 
        RECT 14.94 297.452 19.836 300.716 ; 
        RECT 0.684 297.054 14.868 301.428 ; 
        RECT 0 297.054 0.612 300.716 ; 
        RECT 20.376 297.054 38.448 300.332 ; 
        RECT 0 297.452 20.304 300.332 ; 
        RECT 19.476 297.054 38.448 297.74 ; 
        RECT 0 297.054 19.404 300.332 ; 
        RECT 0 297.054 38.448 297.356 ; 
        RECT 0 305.228 38.448 305.748 ; 
        RECT 37.98 301.374 38.448 305.748 ; 
        RECT 23.364 304.844 37.908 305.748 ; 
        RECT 18.036 304.844 23.292 305.748 ; 
        RECT 15.156 301.374 17.676 305.748 ; 
        RECT 0.54 304.844 15.084 305.748 ; 
        RECT 0 301.374 0.468 305.748 ; 
        RECT 37.836 301.374 38.448 305.036 ; 
        RECT 23.58 301.374 37.764 305.748 ; 
        RECT 20.592 301.374 23.508 305.036 ; 
        RECT 19.944 302.156 20.448 305.748 ; 
        RECT 14.94 301.772 19.836 305.036 ; 
        RECT 0.684 301.374 14.868 305.748 ; 
        RECT 0 301.374 0.612 305.036 ; 
        RECT 20.376 301.374 38.448 304.652 ; 
        RECT 0 301.772 20.304 304.652 ; 
        RECT 19.476 301.374 38.448 302.06 ; 
        RECT 0 301.374 19.404 304.652 ; 
        RECT 0 301.374 38.448 301.676 ; 
        RECT 0 309.548 38.448 310.068 ; 
        RECT 37.98 305.694 38.448 310.068 ; 
        RECT 23.364 309.164 37.908 310.068 ; 
        RECT 18.036 309.164 23.292 310.068 ; 
        RECT 15.156 305.694 17.676 310.068 ; 
        RECT 0.54 309.164 15.084 310.068 ; 
        RECT 0 305.694 0.468 310.068 ; 
        RECT 37.836 305.694 38.448 309.356 ; 
        RECT 23.58 305.694 37.764 310.068 ; 
        RECT 20.592 305.694 23.508 309.356 ; 
        RECT 19.944 306.476 20.448 310.068 ; 
        RECT 14.94 306.092 19.836 309.356 ; 
        RECT 0.684 305.694 14.868 310.068 ; 
        RECT 0 305.694 0.612 309.356 ; 
        RECT 20.376 305.694 38.448 308.972 ; 
        RECT 0 306.092 20.304 308.972 ; 
        RECT 19.476 305.694 38.448 306.38 ; 
        RECT 0 305.694 19.404 308.972 ; 
        RECT 0 305.694 38.448 305.996 ; 
        RECT 0 313.868 38.448 314.388 ; 
        RECT 37.98 310.014 38.448 314.388 ; 
        RECT 23.364 313.484 37.908 314.388 ; 
        RECT 18.036 313.484 23.292 314.388 ; 
        RECT 15.156 310.014 17.676 314.388 ; 
        RECT 0.54 313.484 15.084 314.388 ; 
        RECT 0 310.014 0.468 314.388 ; 
        RECT 37.836 310.014 38.448 313.676 ; 
        RECT 23.58 310.014 37.764 314.388 ; 
        RECT 20.592 310.014 23.508 313.676 ; 
        RECT 19.944 310.796 20.448 314.388 ; 
        RECT 14.94 310.412 19.836 313.676 ; 
        RECT 0.684 310.014 14.868 314.388 ; 
        RECT 0 310.014 0.612 313.676 ; 
        RECT 20.376 310.014 38.448 313.292 ; 
        RECT 0 310.412 20.304 313.292 ; 
        RECT 19.476 310.014 38.448 310.7 ; 
        RECT 0 310.014 19.404 313.292 ; 
        RECT 0 310.014 38.448 310.316 ; 
        RECT 0 318.188 38.448 318.708 ; 
        RECT 37.98 314.334 38.448 318.708 ; 
        RECT 23.364 317.804 37.908 318.708 ; 
        RECT 18.036 317.804 23.292 318.708 ; 
        RECT 15.156 314.334 17.676 318.708 ; 
        RECT 0.54 317.804 15.084 318.708 ; 
        RECT 0 314.334 0.468 318.708 ; 
        RECT 37.836 314.334 38.448 317.996 ; 
        RECT 23.58 314.334 37.764 318.708 ; 
        RECT 20.592 314.334 23.508 317.996 ; 
        RECT 19.944 315.116 20.448 318.708 ; 
        RECT 14.94 314.732 19.836 317.996 ; 
        RECT 0.684 314.334 14.868 318.708 ; 
        RECT 0 314.334 0.612 317.996 ; 
        RECT 20.376 314.334 38.448 317.612 ; 
        RECT 0 314.732 20.304 317.612 ; 
        RECT 19.476 314.334 38.448 315.02 ; 
        RECT 0 314.334 19.404 317.612 ; 
        RECT 0 314.334 38.448 314.636 ; 
        RECT 0 322.508 38.448 323.028 ; 
        RECT 37.98 318.654 38.448 323.028 ; 
        RECT 23.364 322.124 37.908 323.028 ; 
        RECT 18.036 322.124 23.292 323.028 ; 
        RECT 15.156 318.654 17.676 323.028 ; 
        RECT 0.54 322.124 15.084 323.028 ; 
        RECT 0 318.654 0.468 323.028 ; 
        RECT 37.836 318.654 38.448 322.316 ; 
        RECT 23.58 318.654 37.764 323.028 ; 
        RECT 20.592 318.654 23.508 322.316 ; 
        RECT 19.944 319.436 20.448 323.028 ; 
        RECT 14.94 319.052 19.836 322.316 ; 
        RECT 0.684 318.654 14.868 323.028 ; 
        RECT 0 318.654 0.612 322.316 ; 
        RECT 20.376 318.654 38.448 321.932 ; 
        RECT 0 319.052 20.304 321.932 ; 
        RECT 19.476 318.654 38.448 319.34 ; 
        RECT 0 318.654 19.404 321.932 ; 
        RECT 0 318.654 38.448 318.956 ; 
        RECT 0 326.828 38.448 327.348 ; 
        RECT 37.98 322.974 38.448 327.348 ; 
        RECT 23.364 326.444 37.908 327.348 ; 
        RECT 18.036 326.444 23.292 327.348 ; 
        RECT 15.156 322.974 17.676 327.348 ; 
        RECT 0.54 326.444 15.084 327.348 ; 
        RECT 0 322.974 0.468 327.348 ; 
        RECT 37.836 322.974 38.448 326.636 ; 
        RECT 23.58 322.974 37.764 327.348 ; 
        RECT 20.592 322.974 23.508 326.636 ; 
        RECT 19.944 323.756 20.448 327.348 ; 
        RECT 14.94 323.372 19.836 326.636 ; 
        RECT 0.684 322.974 14.868 327.348 ; 
        RECT 0 322.974 0.612 326.636 ; 
        RECT 20.376 322.974 38.448 326.252 ; 
        RECT 0 323.372 20.304 326.252 ; 
        RECT 19.476 322.974 38.448 323.66 ; 
        RECT 0 322.974 19.404 326.252 ; 
        RECT 0 322.974 38.448 323.276 ; 
        RECT 0 331.148 38.448 331.668 ; 
        RECT 37.98 327.294 38.448 331.668 ; 
        RECT 23.364 330.764 37.908 331.668 ; 
        RECT 18.036 330.764 23.292 331.668 ; 
        RECT 15.156 327.294 17.676 331.668 ; 
        RECT 0.54 330.764 15.084 331.668 ; 
        RECT 0 327.294 0.468 331.668 ; 
        RECT 37.836 327.294 38.448 330.956 ; 
        RECT 23.58 327.294 37.764 331.668 ; 
        RECT 20.592 327.294 23.508 330.956 ; 
        RECT 19.944 328.076 20.448 331.668 ; 
        RECT 14.94 327.692 19.836 330.956 ; 
        RECT 0.684 327.294 14.868 331.668 ; 
        RECT 0 327.294 0.612 330.956 ; 
        RECT 20.376 327.294 38.448 330.572 ; 
        RECT 0 327.692 20.304 330.572 ; 
        RECT 19.476 327.294 38.448 327.98 ; 
        RECT 0 327.294 19.404 330.572 ; 
        RECT 0 327.294 38.448 327.596 ; 
        RECT 0 335.468 38.448 335.988 ; 
        RECT 37.98 331.614 38.448 335.988 ; 
        RECT 23.364 335.084 37.908 335.988 ; 
        RECT 18.036 335.084 23.292 335.988 ; 
        RECT 15.156 331.614 17.676 335.988 ; 
        RECT 0.54 335.084 15.084 335.988 ; 
        RECT 0 331.614 0.468 335.988 ; 
        RECT 37.836 331.614 38.448 335.276 ; 
        RECT 23.58 331.614 37.764 335.988 ; 
        RECT 20.592 331.614 23.508 335.276 ; 
        RECT 19.944 332.396 20.448 335.988 ; 
        RECT 14.94 332.012 19.836 335.276 ; 
        RECT 0.684 331.614 14.868 335.988 ; 
        RECT 0 331.614 0.612 335.276 ; 
        RECT 20.376 331.614 38.448 334.892 ; 
        RECT 0 332.012 20.304 334.892 ; 
        RECT 19.476 331.614 38.448 332.3 ; 
        RECT 0 331.614 19.404 334.892 ; 
        RECT 0 331.614 38.448 331.916 ; 
        RECT 0 339.788 38.448 340.308 ; 
        RECT 37.98 335.934 38.448 340.308 ; 
        RECT 23.364 339.404 37.908 340.308 ; 
        RECT 18.036 339.404 23.292 340.308 ; 
        RECT 15.156 335.934 17.676 340.308 ; 
        RECT 0.54 339.404 15.084 340.308 ; 
        RECT 0 335.934 0.468 340.308 ; 
        RECT 37.836 335.934 38.448 339.596 ; 
        RECT 23.58 335.934 37.764 340.308 ; 
        RECT 20.592 335.934 23.508 339.596 ; 
        RECT 19.944 336.716 20.448 340.308 ; 
        RECT 14.94 336.332 19.836 339.596 ; 
        RECT 0.684 335.934 14.868 340.308 ; 
        RECT 0 335.934 0.612 339.596 ; 
        RECT 20.376 335.934 38.448 339.212 ; 
        RECT 0 336.332 20.304 339.212 ; 
        RECT 19.476 335.934 38.448 336.62 ; 
        RECT 0 335.934 19.404 339.212 ; 
        RECT 0 335.934 38.448 336.236 ; 
        RECT 0 344.108 38.448 344.628 ; 
        RECT 37.98 340.254 38.448 344.628 ; 
        RECT 23.364 343.724 37.908 344.628 ; 
        RECT 18.036 343.724 23.292 344.628 ; 
        RECT 15.156 340.254 17.676 344.628 ; 
        RECT 0.54 343.724 15.084 344.628 ; 
        RECT 0 340.254 0.468 344.628 ; 
        RECT 37.836 340.254 38.448 343.916 ; 
        RECT 23.58 340.254 37.764 344.628 ; 
        RECT 20.592 340.254 23.508 343.916 ; 
        RECT 19.944 341.036 20.448 344.628 ; 
        RECT 14.94 340.652 19.836 343.916 ; 
        RECT 0.684 340.254 14.868 344.628 ; 
        RECT 0 340.254 0.612 343.916 ; 
        RECT 20.376 340.254 38.448 343.532 ; 
        RECT 0 340.652 20.304 343.532 ; 
        RECT 19.476 340.254 38.448 340.94 ; 
        RECT 0 340.254 19.404 343.532 ; 
        RECT 0 340.254 38.448 340.556 ; 
        RECT 0 348.428 38.448 348.948 ; 
        RECT 37.98 344.574 38.448 348.948 ; 
        RECT 23.364 348.044 37.908 348.948 ; 
        RECT 18.036 348.044 23.292 348.948 ; 
        RECT 15.156 344.574 17.676 348.948 ; 
        RECT 0.54 348.044 15.084 348.948 ; 
        RECT 0 344.574 0.468 348.948 ; 
        RECT 37.836 344.574 38.448 348.236 ; 
        RECT 23.58 344.574 37.764 348.948 ; 
        RECT 20.592 344.574 23.508 348.236 ; 
        RECT 19.944 345.356 20.448 348.948 ; 
        RECT 14.94 344.972 19.836 348.236 ; 
        RECT 0.684 344.574 14.868 348.948 ; 
        RECT 0 344.574 0.612 348.236 ; 
        RECT 20.376 344.574 38.448 347.852 ; 
        RECT 0 344.972 20.304 347.852 ; 
        RECT 19.476 344.574 38.448 345.26 ; 
        RECT 0 344.574 19.404 347.852 ; 
        RECT 0 344.574 38.448 344.876 ; 
        RECT 0 352.748 38.448 353.268 ; 
        RECT 37.98 348.894 38.448 353.268 ; 
        RECT 23.364 352.364 37.908 353.268 ; 
        RECT 18.036 352.364 23.292 353.268 ; 
        RECT 15.156 348.894 17.676 353.268 ; 
        RECT 0.54 352.364 15.084 353.268 ; 
        RECT 0 348.894 0.468 353.268 ; 
        RECT 37.836 348.894 38.448 352.556 ; 
        RECT 23.58 348.894 37.764 353.268 ; 
        RECT 20.592 348.894 23.508 352.556 ; 
        RECT 19.944 349.676 20.448 353.268 ; 
        RECT 14.94 349.292 19.836 352.556 ; 
        RECT 0.684 348.894 14.868 353.268 ; 
        RECT 0 348.894 0.612 352.556 ; 
        RECT 20.376 348.894 38.448 352.172 ; 
        RECT 0 349.292 20.304 352.172 ; 
        RECT 19.476 348.894 38.448 349.58 ; 
        RECT 0 348.894 19.404 352.172 ; 
        RECT 0 348.894 38.448 349.196 ; 
        RECT 0 357.068 38.448 357.588 ; 
        RECT 37.98 353.214 38.448 357.588 ; 
        RECT 23.364 356.684 37.908 357.588 ; 
        RECT 18.036 356.684 23.292 357.588 ; 
        RECT 15.156 353.214 17.676 357.588 ; 
        RECT 0.54 356.684 15.084 357.588 ; 
        RECT 0 353.214 0.468 357.588 ; 
        RECT 37.836 353.214 38.448 356.876 ; 
        RECT 23.58 353.214 37.764 357.588 ; 
        RECT 20.592 353.214 23.508 356.876 ; 
        RECT 19.944 353.996 20.448 357.588 ; 
        RECT 14.94 353.612 19.836 356.876 ; 
        RECT 0.684 353.214 14.868 357.588 ; 
        RECT 0 353.214 0.612 356.876 ; 
        RECT 20.376 353.214 38.448 356.492 ; 
        RECT 0 353.612 20.304 356.492 ; 
        RECT 19.476 353.214 38.448 353.9 ; 
        RECT 0 353.214 19.404 356.492 ; 
        RECT 0 353.214 38.448 353.516 ; 
        RECT 0 361.388 38.448 361.908 ; 
        RECT 37.98 357.534 38.448 361.908 ; 
        RECT 23.364 361.004 37.908 361.908 ; 
        RECT 18.036 361.004 23.292 361.908 ; 
        RECT 15.156 357.534 17.676 361.908 ; 
        RECT 0.54 361.004 15.084 361.908 ; 
        RECT 0 357.534 0.468 361.908 ; 
        RECT 37.836 357.534 38.448 361.196 ; 
        RECT 23.58 357.534 37.764 361.908 ; 
        RECT 20.592 357.534 23.508 361.196 ; 
        RECT 19.944 358.316 20.448 361.908 ; 
        RECT 14.94 357.932 19.836 361.196 ; 
        RECT 0.684 357.534 14.868 361.908 ; 
        RECT 0 357.534 0.612 361.196 ; 
        RECT 20.376 357.534 38.448 360.812 ; 
        RECT 0 357.932 20.304 360.812 ; 
        RECT 19.476 357.534 38.448 358.22 ; 
        RECT 0 357.534 19.404 360.812 ; 
        RECT 0 357.534 38.448 357.836 ; 
        RECT 0 365.708 38.448 366.228 ; 
        RECT 37.98 361.854 38.448 366.228 ; 
        RECT 23.364 365.324 37.908 366.228 ; 
        RECT 18.036 365.324 23.292 366.228 ; 
        RECT 15.156 361.854 17.676 366.228 ; 
        RECT 0.54 365.324 15.084 366.228 ; 
        RECT 0 361.854 0.468 366.228 ; 
        RECT 37.836 361.854 38.448 365.516 ; 
        RECT 23.58 361.854 37.764 366.228 ; 
        RECT 20.592 361.854 23.508 365.516 ; 
        RECT 19.944 362.636 20.448 366.228 ; 
        RECT 14.94 362.252 19.836 365.516 ; 
        RECT 0.684 361.854 14.868 366.228 ; 
        RECT 0 361.854 0.612 365.516 ; 
        RECT 20.376 361.854 38.448 365.132 ; 
        RECT 0 362.252 20.304 365.132 ; 
        RECT 19.476 361.854 38.448 362.54 ; 
        RECT 0 361.854 19.404 365.132 ; 
        RECT 0 361.854 38.448 362.156 ; 
        RECT 0 370.028 38.448 370.548 ; 
        RECT 37.98 366.174 38.448 370.548 ; 
        RECT 23.364 369.644 37.908 370.548 ; 
        RECT 18.036 369.644 23.292 370.548 ; 
        RECT 15.156 366.174 17.676 370.548 ; 
        RECT 0.54 369.644 15.084 370.548 ; 
        RECT 0 366.174 0.468 370.548 ; 
        RECT 37.836 366.174 38.448 369.836 ; 
        RECT 23.58 366.174 37.764 370.548 ; 
        RECT 20.592 366.174 23.508 369.836 ; 
        RECT 19.944 366.956 20.448 370.548 ; 
        RECT 14.94 366.572 19.836 369.836 ; 
        RECT 0.684 366.174 14.868 370.548 ; 
        RECT 0 366.174 0.612 369.836 ; 
        RECT 20.376 366.174 38.448 369.452 ; 
        RECT 0 366.572 20.304 369.452 ; 
        RECT 19.476 366.174 38.448 366.86 ; 
        RECT 0 366.174 19.404 369.452 ; 
        RECT 0 366.174 38.448 366.476 ; 
        RECT 0 374.348 38.448 374.868 ; 
        RECT 37.98 370.494 38.448 374.868 ; 
        RECT 23.364 373.964 37.908 374.868 ; 
        RECT 18.036 373.964 23.292 374.868 ; 
        RECT 15.156 370.494 17.676 374.868 ; 
        RECT 0.54 373.964 15.084 374.868 ; 
        RECT 0 370.494 0.468 374.868 ; 
        RECT 37.836 370.494 38.448 374.156 ; 
        RECT 23.58 370.494 37.764 374.868 ; 
        RECT 20.592 370.494 23.508 374.156 ; 
        RECT 19.944 371.276 20.448 374.868 ; 
        RECT 14.94 370.892 19.836 374.156 ; 
        RECT 0.684 370.494 14.868 374.868 ; 
        RECT 0 370.494 0.612 374.156 ; 
        RECT 20.376 370.494 38.448 373.772 ; 
        RECT 0 370.892 20.304 373.772 ; 
        RECT 19.476 370.494 38.448 371.18 ; 
        RECT 0 370.494 19.404 373.772 ; 
        RECT 0 370.494 38.448 370.796 ; 
        RECT 0 378.668 38.448 379.188 ; 
        RECT 37.98 374.814 38.448 379.188 ; 
        RECT 23.364 378.284 37.908 379.188 ; 
        RECT 18.036 378.284 23.292 379.188 ; 
        RECT 15.156 374.814 17.676 379.188 ; 
        RECT 0.54 378.284 15.084 379.188 ; 
        RECT 0 374.814 0.468 379.188 ; 
        RECT 37.836 374.814 38.448 378.476 ; 
        RECT 23.58 374.814 37.764 379.188 ; 
        RECT 20.592 374.814 23.508 378.476 ; 
        RECT 19.944 375.596 20.448 379.188 ; 
        RECT 14.94 375.212 19.836 378.476 ; 
        RECT 0.684 374.814 14.868 379.188 ; 
        RECT 0 374.814 0.612 378.476 ; 
        RECT 20.376 374.814 38.448 378.092 ; 
        RECT 0 375.212 20.304 378.092 ; 
        RECT 19.476 374.814 38.448 375.5 ; 
        RECT 0 374.814 19.404 378.092 ; 
        RECT 0 374.814 38.448 375.116 ; 
  LAYER M4 ; 
      RECT 6.428 180.624 32.01 180.72 ; 
      RECT 6.428 181.776 32.01 181.872 ; 
      RECT 6.428 183.312 32.01 183.408 ; 
      RECT 6.428 183.696 32.01 183.792 ; 
      RECT 6.428 185.04 32.01 185.136 ; 
      RECT 29.996 176.46 30.332 176.556 ; 
      RECT 29.276 178.188 29.744 178.284 ; 
      RECT 29.276 180.816 29.744 180.912 ; 
      RECT 29.276 181.968 29.744 182.064 ; 
      RECT 26.714 178.188 28.992 178.284 ; 
      RECT 26.972 181.296 27.404 181.392 ; 
      RECT 21.628 182.796 26 182.892 ; 
      RECT 24.38 181.068 24.716 181.164 ; 
      RECT 21.244 185.868 24.716 185.964 ; 
      RECT 24.38 186.252 24.716 186.348 ; 
      RECT 23.668 179.148 24.004 179.244 ; 
      RECT 23.516 184.524 23.852 184.62 ; 
      RECT 22.804 178.764 23.14 178.86 ; 
      RECT 21.948 173.612 23 173.708 ; 
      RECT 21.948 208.172 23 208.268 ; 
      RECT 22.012 184.716 22.988 184.812 ; 
      RECT 22.652 185.292 22.988 185.388 ; 
      RECT 16.828 186.252 22.988 186.348 ; 
      RECT 22.652 187.404 22.988 187.5 ; 
      RECT 21.716 207.788 22.768 207.884 ; 
      RECT 21.712 173.228 22.764 173.324 ; 
      RECT 21.56 172.844 22.612 172.94 ; 
      RECT 21.56 207.02 22.612 207.116 ; 
      RECT 22.22 189.132 22.556 189.228 ; 
      RECT 19.132 190.668 22.556 190.764 ; 
      RECT 20.668 199.692 22.556 199.788 ; 
      RECT 22.22 200.076 22.556 200.172 ; 
      RECT 21.368 172.46 22.42 172.556 ; 
      RECT 21.368 206.636 22.42 206.732 ; 
      RECT 20.476 196.044 22.256 196.14 ; 
      RECT 21.192 172.076 22.244 172.172 ; 
      RECT 21.192 207.98 22.244 208.076 ; 
      RECT 20.996 173.42 22.048 173.516 ; 
      RECT 20.996 207.596 22.048 207.692 ; 
      RECT 21.52 185.292 22.004 185.388 ; 
      RECT 21.436 193.74 21.968 193.836 ; 
      RECT 20.808 173.036 21.86 173.132 ; 
      RECT 20.808 207.212 21.86 207.308 ; 
      RECT 20.668 171.884 21.72 171.98 ; 
      RECT 20.668 206.828 21.72 206.924 ; 
      RECT 17.404 200.076 21.68 200.172 ; 
      RECT 21.344 204.684 21.68 204.78 ; 
      RECT 20.444 171.308 21.496 171.404 ; 
      RECT 20.444 206.444 21.496 206.54 ; 
      RECT 21.052 189.132 21.392 189.228 ; 
      RECT 16.636 191.436 21.104 191.532 ; 
      RECT 19.216 182.796 21.044 182.892 ; 
      RECT 18.524 174.188 19.592 174.284 ; 
      RECT 18.524 205.868 19.592 205.964 ; 
      RECT 19.072 188.94 19.508 189.036 ; 
      RECT 18.432 173.804 19.4 173.9 ; 
      RECT 18.432 208.364 19.4 208.46 ; 
      RECT 18.208 171.884 19.176 171.98 ; 
      RECT 18.324 208.748 19.176 208.844 ; 
      RECT 18.788 187.404 19.124 187.5 ; 
      RECT 17.992 172.268 18.984 172.364 ; 
      RECT 17.992 208.172 18.984 208.268 ; 
      RECT 17.056 197.772 18.74 197.868 ; 
      RECT 16.928 173.612 17.996 173.708 ; 
      RECT 16.928 208.748 17.996 208.844 ; 
      RECT 17.488 192.012 17.972 192.108 ; 
      RECT 17.456 204.684 17.792 204.78 ; 
      RECT 16.792 173.228 17.78 173.324 ; 
      RECT 16.524 207.02 17.78 207.116 ; 
      RECT 16.688 172.844 17.608 172.94 ; 
      RECT 16.64 208.364 17.608 208.46 ; 
      RECT 16.476 172.46 17.396 172.556 ; 
      RECT 17.06 198.348 17.396 198.444 ; 
      RECT 16.276 206.636 17.396 206.732 ; 
      RECT 16.296 172.076 17.216 172.172 ; 
      RECT 16.296 207.98 17.216 208.076 ; 
      RECT 12.448 187.404 17.204 187.5 ; 
      RECT 16.144 173.036 17.064 173.132 ; 
      RECT 16.144 207.596 17.064 207.692 ; 
      RECT 16.072 172.652 16.844 172.748 ; 
      RECT 16.072 207.212 16.844 207.308 ; 
      RECT 15.876 172.268 16.648 172.364 ; 
      RECT 15.876 206.828 16.648 206.924 ; 
      RECT 15.892 191.052 16.628 191.148 ; 
      RECT 15.668 171.884 16.44 171.98 ; 
      RECT 15.668 206.444 16.44 206.54 ; 
      RECT 13.732 180.3 16.436 180.396 ; 
      RECT 15.892 191.436 16.228 191.532 ; 
      RECT 14.816 173.996 15.868 174.092 ; 
      RECT 15.032 189.132 15.48 189.228 ; 
      RECT 13.58 181.068 13.916 181.164 ; 
  LAYER V4 ; 
      RECT 30.192 176.46 30.288 176.556 ; 
      RECT 30.192 180.624 30.288 180.72 ; 
      RECT 29.52 178.188 29.616 178.284 ; 
      RECT 29.52 180.816 29.616 180.912 ; 
      RECT 29.52 181.968 29.616 182.064 ; 
      RECT 27.024 178.188 27.12 178.284 ; 
      RECT 27.024 181.296 27.12 181.392 ; 
      RECT 24.576 181.068 24.672 181.164 ; 
      RECT 24.576 181.776 24.672 181.872 ; 
      RECT 24.576 185.868 24.672 185.964 ; 
      RECT 24.576 186.252 24.672 186.348 ; 
      RECT 23.712 179.148 23.808 179.244 ; 
      RECT 23.712 183.312 23.808 183.408 ; 
      RECT 23.712 184.524 23.808 184.62 ; 
      RECT 23.712 185.04 23.808 185.136 ; 
      RECT 22.848 178.764 22.944 178.86 ; 
      RECT 22.848 183.696 22.944 183.792 ; 
      RECT 22.848 184.716 22.944 184.812 ; 
      RECT 22.848 185.292 22.944 185.388 ; 
      RECT 22.848 186.252 22.944 186.348 ; 
      RECT 22.848 187.404 22.944 187.5 ; 
      RECT 22.416 189.132 22.512 189.228 ; 
      RECT 22.416 190.668 22.512 190.764 ; 
      RECT 22.416 199.692 22.512 199.788 ; 
      RECT 22.416 200.076 22.512 200.172 ; 
      RECT 22.056 173.612 22.152 173.708 ; 
      RECT 22.056 184.716 22.152 184.812 ; 
      RECT 22.056 208.172 22.152 208.268 ; 
      RECT 21.864 173.228 21.96 173.324 ; 
      RECT 21.864 185.292 21.96 185.388 ; 
      RECT 21.864 207.788 21.96 207.884 ; 
      RECT 21.672 172.844 21.768 172.94 ; 
      RECT 21.672 182.796 21.768 182.892 ; 
      RECT 21.672 207.02 21.768 207.116 ; 
      RECT 21.48 172.46 21.576 172.556 ; 
      RECT 21.48 193.74 21.576 193.836 ; 
      RECT 21.48 204.684 21.576 204.78 ; 
      RECT 21.48 206.636 21.576 206.732 ; 
      RECT 21.288 172.076 21.384 172.172 ; 
      RECT 21.288 185.868 21.384 185.964 ; 
      RECT 21.288 207.98 21.384 208.076 ; 
      RECT 21.096 173.42 21.192 173.516 ; 
      RECT 21.096 189.132 21.192 189.228 ; 
      RECT 21.096 207.596 21.192 207.692 ; 
      RECT 20.904 173.036 21 173.132 ; 
      RECT 20.904 182.796 21 182.892 ; 
      RECT 20.904 207.212 21 207.308 ; 
      RECT 20.712 171.884 20.808 171.98 ; 
      RECT 20.712 199.692 20.808 199.788 ; 
      RECT 20.712 206.828 20.808 206.924 ; 
      RECT 20.52 171.308 20.616 171.404 ; 
      RECT 20.52 196.044 20.616 196.14 ; 
      RECT 20.52 206.444 20.616 206.54 ; 
      RECT 19.368 174.188 19.464 174.284 ; 
      RECT 19.368 188.94 19.464 189.036 ; 
      RECT 19.368 205.868 19.464 205.964 ; 
      RECT 19.176 173.804 19.272 173.9 ; 
      RECT 19.176 190.668 19.272 190.764 ; 
      RECT 19.176 208.364 19.272 208.46 ; 
      RECT 18.984 171.884 19.08 171.98 ; 
      RECT 18.984 187.404 19.08 187.5 ; 
      RECT 18.984 208.748 19.08 208.844 ; 
      RECT 18.6 172.268 18.696 172.364 ; 
      RECT 18.6 197.772 18.696 197.868 ; 
      RECT 18.6 208.172 18.696 208.268 ; 
      RECT 17.832 173.612 17.928 173.708 ; 
      RECT 17.832 192.012 17.928 192.108 ; 
      RECT 17.832 208.748 17.928 208.844 ; 
      RECT 17.64 173.228 17.736 173.324 ; 
      RECT 17.64 204.684 17.736 204.78 ; 
      RECT 17.64 207.02 17.736 207.116 ; 
      RECT 17.448 172.844 17.544 172.94 ; 
      RECT 17.448 200.076 17.544 200.172 ; 
      RECT 17.448 208.364 17.544 208.46 ; 
      RECT 17.256 172.46 17.352 172.556 ; 
      RECT 17.256 198.348 17.352 198.444 ; 
      RECT 17.256 206.636 17.352 206.732 ; 
      RECT 17.064 172.076 17.16 172.172 ; 
      RECT 17.064 187.404 17.16 187.5 ; 
      RECT 17.064 207.98 17.16 208.076 ; 
      RECT 16.872 173.036 16.968 173.132 ; 
      RECT 16.872 186.252 16.968 186.348 ; 
      RECT 16.872 207.596 16.968 207.692 ; 
      RECT 16.68 172.652 16.776 172.748 ; 
      RECT 16.68 191.436 16.776 191.532 ; 
      RECT 16.68 207.212 16.776 207.308 ; 
      RECT 16.488 172.268 16.584 172.364 ; 
      RECT 16.488 191.052 16.584 191.148 ; 
      RECT 16.488 206.828 16.584 206.924 ; 
      RECT 16.296 171.884 16.392 171.98 ; 
      RECT 16.296 180.3 16.392 180.396 ; 
      RECT 16.296 206.444 16.392 206.54 ; 
      RECT 15.936 191.052 16.032 191.148 ; 
      RECT 15.936 191.436 16.032 191.532 ; 
      RECT 15.268 173.996 15.364 174.092 ; 
      RECT 15.268 189.132 15.364 189.228 ; 
      RECT 13.776 180.3 13.872 180.396 ; 
      RECT 13.776 181.068 13.872 181.164 ; 
  LAYER M5 ; 
      RECT 30.192 176.416 30.288 180.764 ; 
      RECT 29.52 178.134 29.616 182.264 ; 
      RECT 27.024 178.11 27.12 181.44 ; 
      RECT 24.576 181.024 24.672 181.916 ; 
      RECT 24.576 185.824 24.672 186.392 ; 
      RECT 23.712 179.104 23.808 183.452 ; 
      RECT 23.712 184.48 23.808 185.18 ; 
      RECT 22.848 178.72 22.944 183.836 ; 
      RECT 22.848 184.672 22.944 185.432 ; 
      RECT 22.848 186.208 22.944 187.544 ; 
      RECT 22.416 189.088 22.512 190.808 ; 
      RECT 22.416 199.648 22.512 200.216 ; 
      RECT 22.056 174.96 22.152 205.292 ; 
      RECT 21.864 174.96 21.96 205.292 ; 
      RECT 21.672 174.96 21.768 205.292 ; 
      RECT 21.48 174.96 21.576 205.292 ; 
      RECT 21.288 174.96 21.384 205.292 ; 
      RECT 21.096 174.96 21.192 205.292 ; 
      RECT 20.904 174.96 21 205.292 ; 
      RECT 20.712 174.96 20.808 205.292 ; 
      RECT 20.52 174.96 20.616 205.292 ; 
      RECT 19.368 173.912 19.464 206.044 ; 
      RECT 19.176 171.828 19.272 209.144 ; 
      RECT 18.984 171.704 19.08 209.14 ; 
      RECT 18.6 171.888 18.696 209.144 ; 
      RECT 17.832 171.884 17.928 208.956 ; 
      RECT 17.64 171.884 17.736 208.956 ; 
      RECT 17.448 171.884 17.544 208.956 ; 
      RECT 17.256 171.884 17.352 208.956 ; 
      RECT 17.064 171.884 17.16 208.956 ; 
      RECT 16.872 171.768 16.968 208.956 ; 
      RECT 16.68 171.592 16.776 208.96 ; 
      RECT 16.488 171.444 16.584 208.964 ; 
      RECT 16.296 171.204 16.392 208.964 ; 
      RECT 15.936 191.008 16.032 191.576 ; 
      RECT 15.268 173.924 15.364 189.3 ; 
      RECT 13.776 180.256 13.872 181.208 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 38.016 380.016 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 38.016 380.016 ; 
  END 
END srambank_64x4x80_6t122 
