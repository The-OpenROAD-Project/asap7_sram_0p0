VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_64x4x80_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_64x4x80_6t122 0 0 ;
  SIZE 9.612 BY 95.04 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1010 1.1720 9.5090 1.2200 ;
        RECT 0.1010 2.2520 9.5090 2.3000 ;
        RECT 0.1010 3.3320 9.5090 3.3800 ;
        RECT 0.1010 4.4120 9.5090 4.4600 ;
        RECT 0.1010 5.4920 9.5090 5.5400 ;
        RECT 0.1010 6.5720 9.5090 6.6200 ;
        RECT 0.1010 7.6520 9.5090 7.7000 ;
        RECT 0.1010 8.7320 9.5090 8.7800 ;
        RECT 0.1010 9.8120 9.5090 9.8600 ;
        RECT 0.1010 10.8920 9.5090 10.9400 ;
        RECT 0.1010 11.9720 9.5090 12.0200 ;
        RECT 0.1010 13.0520 9.5090 13.1000 ;
        RECT 0.1010 14.1320 9.5090 14.1800 ;
        RECT 0.1010 15.2120 9.5090 15.2600 ;
        RECT 0.1010 16.2920 9.5090 16.3400 ;
        RECT 0.1010 17.3720 9.5090 17.4200 ;
        RECT 0.1010 18.4520 9.5090 18.5000 ;
        RECT 0.1010 19.5320 9.5090 19.5800 ;
        RECT 0.1010 20.6120 9.5090 20.6600 ;
        RECT 0.1010 21.6920 9.5090 21.7400 ;
        RECT 0.1010 22.7720 9.5090 22.8200 ;
        RECT 0.1010 23.8520 9.5090 23.9000 ;
        RECT 0.1010 24.9320 9.5090 24.9800 ;
        RECT 0.1010 26.0120 9.5090 26.0600 ;
        RECT 0.1010 27.0920 9.5090 27.1400 ;
        RECT 0.1010 28.1720 9.5090 28.2200 ;
        RECT 0.1010 29.2520 9.5090 29.3000 ;
        RECT 0.1010 30.3320 9.5090 30.3800 ;
        RECT 0.1010 31.4120 9.5090 31.4600 ;
        RECT 0.1010 32.4920 9.5090 32.5400 ;
        RECT 0.1010 33.5720 9.5090 33.6200 ;
        RECT 0.1010 34.6520 9.5090 34.7000 ;
        RECT 0.1010 35.7320 9.5090 35.7800 ;
        RECT 0.1010 36.8120 9.5090 36.8600 ;
        RECT 0.1010 37.8920 9.5090 37.9400 ;
        RECT 0.1010 38.9720 9.5090 39.0200 ;
        RECT 0.1010 40.0520 9.5090 40.1000 ;
        RECT 0.1010 41.1320 9.5090 41.1800 ;
        RECT 0.1010 42.2120 9.5090 42.2600 ;
        RECT 0.1010 43.2920 9.5090 43.3400 ;
        RECT 0.1080 43.7790 9.5040 43.9950 ;
        RECT 5.6100 43.4990 5.8730 43.5230 ;
        RECT 5.7410 47.2830 5.8530 47.3070 ;
        RECT 3.9420 46.9470 5.6700 47.1630 ;
        RECT 3.9420 50.1150 5.6700 50.3310 ;
        RECT 0.1010 52.4990 9.5090 52.5470 ;
        RECT 0.1010 53.5790 9.5090 53.6270 ;
        RECT 0.1010 54.6590 9.5090 54.7070 ;
        RECT 0.1010 55.7390 9.5090 55.7870 ;
        RECT 0.1010 56.8190 9.5090 56.8670 ;
        RECT 0.1010 57.8990 9.5090 57.9470 ;
        RECT 0.1010 58.9790 9.5090 59.0270 ;
        RECT 0.1010 60.0590 9.5090 60.1070 ;
        RECT 0.1010 61.1390 9.5090 61.1870 ;
        RECT 0.1010 62.2190 9.5090 62.2670 ;
        RECT 0.1010 63.2990 9.5090 63.3470 ;
        RECT 0.1010 64.3790 9.5090 64.4270 ;
        RECT 0.1010 65.4590 9.5090 65.5070 ;
        RECT 0.1010 66.5390 9.5090 66.5870 ;
        RECT 0.1010 67.6190 9.5090 67.6670 ;
        RECT 0.1010 68.6990 9.5090 68.7470 ;
        RECT 0.1010 69.7790 9.5090 69.8270 ;
        RECT 0.1010 70.8590 9.5090 70.9070 ;
        RECT 0.1010 71.9390 9.5090 71.9870 ;
        RECT 0.1010 73.0190 9.5090 73.0670 ;
        RECT 0.1010 74.0990 9.5090 74.1470 ;
        RECT 0.1010 75.1790 9.5090 75.2270 ;
        RECT 0.1010 76.2590 9.5090 76.3070 ;
        RECT 0.1010 77.3390 9.5090 77.3870 ;
        RECT 0.1010 78.4190 9.5090 78.4670 ;
        RECT 0.1010 79.4990 9.5090 79.5470 ;
        RECT 0.1010 80.5790 9.5090 80.6270 ;
        RECT 0.1010 81.6590 9.5090 81.7070 ;
        RECT 0.1010 82.7390 9.5090 82.7870 ;
        RECT 0.1010 83.8190 9.5090 83.8670 ;
        RECT 0.1010 84.8990 9.5090 84.9470 ;
        RECT 0.1010 85.9790 9.5090 86.0270 ;
        RECT 0.1010 87.0590 9.5090 87.1070 ;
        RECT 0.1010 88.1390 9.5090 88.1870 ;
        RECT 0.1010 89.2190 9.5090 89.2670 ;
        RECT 0.1010 90.2990 9.5090 90.3470 ;
        RECT 0.1010 91.3790 9.5090 91.4270 ;
        RECT 0.1010 92.4590 9.5090 92.5070 ;
        RECT 0.1010 93.5390 9.5090 93.5870 ;
        RECT 0.1010 94.6190 9.5090 94.6670 ;
      LAYER M3  ;
        RECT 9.4770 0.2165 9.4950 1.3765 ;
        RECT 5.8230 0.2170 5.8410 1.3760 ;
        RECT 4.4190 0.2530 4.5090 1.3670 ;
        RECT 3.7710 0.2170 3.7890 1.3760 ;
        RECT 0.1170 0.2165 0.1350 1.3765 ;
        RECT 9.4770 1.2965 9.4950 2.4565 ;
        RECT 5.8230 1.2970 5.8410 2.4560 ;
        RECT 4.4190 1.3330 4.5090 2.4470 ;
        RECT 3.7710 1.2970 3.7890 2.4560 ;
        RECT 0.1170 1.2965 0.1350 2.4565 ;
        RECT 9.4770 2.3765 9.4950 3.5365 ;
        RECT 5.8230 2.3770 5.8410 3.5360 ;
        RECT 4.4190 2.4130 4.5090 3.5270 ;
        RECT 3.7710 2.3770 3.7890 3.5360 ;
        RECT 0.1170 2.3765 0.1350 3.5365 ;
        RECT 9.4770 3.4565 9.4950 4.6165 ;
        RECT 5.8230 3.4570 5.8410 4.6160 ;
        RECT 4.4190 3.4930 4.5090 4.6070 ;
        RECT 3.7710 3.4570 3.7890 4.6160 ;
        RECT 0.1170 3.4565 0.1350 4.6165 ;
        RECT 9.4770 4.5365 9.4950 5.6965 ;
        RECT 5.8230 4.5370 5.8410 5.6960 ;
        RECT 4.4190 4.5730 4.5090 5.6870 ;
        RECT 3.7710 4.5370 3.7890 5.6960 ;
        RECT 0.1170 4.5365 0.1350 5.6965 ;
        RECT 9.4770 5.6165 9.4950 6.7765 ;
        RECT 5.8230 5.6170 5.8410 6.7760 ;
        RECT 4.4190 5.6530 4.5090 6.7670 ;
        RECT 3.7710 5.6170 3.7890 6.7760 ;
        RECT 0.1170 5.6165 0.1350 6.7765 ;
        RECT 9.4770 6.6965 9.4950 7.8565 ;
        RECT 5.8230 6.6970 5.8410 7.8560 ;
        RECT 4.4190 6.7330 4.5090 7.8470 ;
        RECT 3.7710 6.6970 3.7890 7.8560 ;
        RECT 0.1170 6.6965 0.1350 7.8565 ;
        RECT 9.4770 7.7765 9.4950 8.9365 ;
        RECT 5.8230 7.7770 5.8410 8.9360 ;
        RECT 4.4190 7.8130 4.5090 8.9270 ;
        RECT 3.7710 7.7770 3.7890 8.9360 ;
        RECT 0.1170 7.7765 0.1350 8.9365 ;
        RECT 9.4770 8.8565 9.4950 10.0165 ;
        RECT 5.8230 8.8570 5.8410 10.0160 ;
        RECT 4.4190 8.8930 4.5090 10.0070 ;
        RECT 3.7710 8.8570 3.7890 10.0160 ;
        RECT 0.1170 8.8565 0.1350 10.0165 ;
        RECT 9.4770 9.9365 9.4950 11.0965 ;
        RECT 5.8230 9.9370 5.8410 11.0960 ;
        RECT 4.4190 9.9730 4.5090 11.0870 ;
        RECT 3.7710 9.9370 3.7890 11.0960 ;
        RECT 0.1170 9.9365 0.1350 11.0965 ;
        RECT 9.4770 11.0165 9.4950 12.1765 ;
        RECT 5.8230 11.0170 5.8410 12.1760 ;
        RECT 4.4190 11.0530 4.5090 12.1670 ;
        RECT 3.7710 11.0170 3.7890 12.1760 ;
        RECT 0.1170 11.0165 0.1350 12.1765 ;
        RECT 9.4770 12.0965 9.4950 13.2565 ;
        RECT 5.8230 12.0970 5.8410 13.2560 ;
        RECT 4.4190 12.1330 4.5090 13.2470 ;
        RECT 3.7710 12.0970 3.7890 13.2560 ;
        RECT 0.1170 12.0965 0.1350 13.2565 ;
        RECT 9.4770 13.1765 9.4950 14.3365 ;
        RECT 5.8230 13.1770 5.8410 14.3360 ;
        RECT 4.4190 13.2130 4.5090 14.3270 ;
        RECT 3.7710 13.1770 3.7890 14.3360 ;
        RECT 0.1170 13.1765 0.1350 14.3365 ;
        RECT 9.4770 14.2565 9.4950 15.4165 ;
        RECT 5.8230 14.2570 5.8410 15.4160 ;
        RECT 4.4190 14.2930 4.5090 15.4070 ;
        RECT 3.7710 14.2570 3.7890 15.4160 ;
        RECT 0.1170 14.2565 0.1350 15.4165 ;
        RECT 9.4770 15.3365 9.4950 16.4965 ;
        RECT 5.8230 15.3370 5.8410 16.4960 ;
        RECT 4.4190 15.3730 4.5090 16.4870 ;
        RECT 3.7710 15.3370 3.7890 16.4960 ;
        RECT 0.1170 15.3365 0.1350 16.4965 ;
        RECT 9.4770 16.4165 9.4950 17.5765 ;
        RECT 5.8230 16.4170 5.8410 17.5760 ;
        RECT 4.4190 16.4530 4.5090 17.5670 ;
        RECT 3.7710 16.4170 3.7890 17.5760 ;
        RECT 0.1170 16.4165 0.1350 17.5765 ;
        RECT 9.4770 17.4965 9.4950 18.6565 ;
        RECT 5.8230 17.4970 5.8410 18.6560 ;
        RECT 4.4190 17.5330 4.5090 18.6470 ;
        RECT 3.7710 17.4970 3.7890 18.6560 ;
        RECT 0.1170 17.4965 0.1350 18.6565 ;
        RECT 9.4770 18.5765 9.4950 19.7365 ;
        RECT 5.8230 18.5770 5.8410 19.7360 ;
        RECT 4.4190 18.6130 4.5090 19.7270 ;
        RECT 3.7710 18.5770 3.7890 19.7360 ;
        RECT 0.1170 18.5765 0.1350 19.7365 ;
        RECT 9.4770 19.6565 9.4950 20.8165 ;
        RECT 5.8230 19.6570 5.8410 20.8160 ;
        RECT 4.4190 19.6930 4.5090 20.8070 ;
        RECT 3.7710 19.6570 3.7890 20.8160 ;
        RECT 0.1170 19.6565 0.1350 20.8165 ;
        RECT 9.4770 20.7365 9.4950 21.8965 ;
        RECT 5.8230 20.7370 5.8410 21.8960 ;
        RECT 4.4190 20.7730 4.5090 21.8870 ;
        RECT 3.7710 20.7370 3.7890 21.8960 ;
        RECT 0.1170 20.7365 0.1350 21.8965 ;
        RECT 9.4770 21.8165 9.4950 22.9765 ;
        RECT 5.8230 21.8170 5.8410 22.9760 ;
        RECT 4.4190 21.8530 4.5090 22.9670 ;
        RECT 3.7710 21.8170 3.7890 22.9760 ;
        RECT 0.1170 21.8165 0.1350 22.9765 ;
        RECT 9.4770 22.8965 9.4950 24.0565 ;
        RECT 5.8230 22.8970 5.8410 24.0560 ;
        RECT 4.4190 22.9330 4.5090 24.0470 ;
        RECT 3.7710 22.8970 3.7890 24.0560 ;
        RECT 0.1170 22.8965 0.1350 24.0565 ;
        RECT 9.4770 23.9765 9.4950 25.1365 ;
        RECT 5.8230 23.9770 5.8410 25.1360 ;
        RECT 4.4190 24.0130 4.5090 25.1270 ;
        RECT 3.7710 23.9770 3.7890 25.1360 ;
        RECT 0.1170 23.9765 0.1350 25.1365 ;
        RECT 9.4770 25.0565 9.4950 26.2165 ;
        RECT 5.8230 25.0570 5.8410 26.2160 ;
        RECT 4.4190 25.0930 4.5090 26.2070 ;
        RECT 3.7710 25.0570 3.7890 26.2160 ;
        RECT 0.1170 25.0565 0.1350 26.2165 ;
        RECT 9.4770 26.1365 9.4950 27.2965 ;
        RECT 5.8230 26.1370 5.8410 27.2960 ;
        RECT 4.4190 26.1730 4.5090 27.2870 ;
        RECT 3.7710 26.1370 3.7890 27.2960 ;
        RECT 0.1170 26.1365 0.1350 27.2965 ;
        RECT 9.4770 27.2165 9.4950 28.3765 ;
        RECT 5.8230 27.2170 5.8410 28.3760 ;
        RECT 4.4190 27.2530 4.5090 28.3670 ;
        RECT 3.7710 27.2170 3.7890 28.3760 ;
        RECT 0.1170 27.2165 0.1350 28.3765 ;
        RECT 9.4770 28.2965 9.4950 29.4565 ;
        RECT 5.8230 28.2970 5.8410 29.4560 ;
        RECT 4.4190 28.3330 4.5090 29.4470 ;
        RECT 3.7710 28.2970 3.7890 29.4560 ;
        RECT 0.1170 28.2965 0.1350 29.4565 ;
        RECT 9.4770 29.3765 9.4950 30.5365 ;
        RECT 5.8230 29.3770 5.8410 30.5360 ;
        RECT 4.4190 29.4130 4.5090 30.5270 ;
        RECT 3.7710 29.3770 3.7890 30.5360 ;
        RECT 0.1170 29.3765 0.1350 30.5365 ;
        RECT 9.4770 30.4565 9.4950 31.6165 ;
        RECT 5.8230 30.4570 5.8410 31.6160 ;
        RECT 4.4190 30.4930 4.5090 31.6070 ;
        RECT 3.7710 30.4570 3.7890 31.6160 ;
        RECT 0.1170 30.4565 0.1350 31.6165 ;
        RECT 9.4770 31.5365 9.4950 32.6965 ;
        RECT 5.8230 31.5370 5.8410 32.6960 ;
        RECT 4.4190 31.5730 4.5090 32.6870 ;
        RECT 3.7710 31.5370 3.7890 32.6960 ;
        RECT 0.1170 31.5365 0.1350 32.6965 ;
        RECT 9.4770 32.6165 9.4950 33.7765 ;
        RECT 5.8230 32.6170 5.8410 33.7760 ;
        RECT 4.4190 32.6530 4.5090 33.7670 ;
        RECT 3.7710 32.6170 3.7890 33.7760 ;
        RECT 0.1170 32.6165 0.1350 33.7765 ;
        RECT 9.4770 33.6965 9.4950 34.8565 ;
        RECT 5.8230 33.6970 5.8410 34.8560 ;
        RECT 4.4190 33.7330 4.5090 34.8470 ;
        RECT 3.7710 33.6970 3.7890 34.8560 ;
        RECT 0.1170 33.6965 0.1350 34.8565 ;
        RECT 9.4770 34.7765 9.4950 35.9365 ;
        RECT 5.8230 34.7770 5.8410 35.9360 ;
        RECT 4.4190 34.8130 4.5090 35.9270 ;
        RECT 3.7710 34.7770 3.7890 35.9360 ;
        RECT 0.1170 34.7765 0.1350 35.9365 ;
        RECT 9.4770 35.8565 9.4950 37.0165 ;
        RECT 5.8230 35.8570 5.8410 37.0160 ;
        RECT 4.4190 35.8930 4.5090 37.0070 ;
        RECT 3.7710 35.8570 3.7890 37.0160 ;
        RECT 0.1170 35.8565 0.1350 37.0165 ;
        RECT 9.4770 36.9365 9.4950 38.0965 ;
        RECT 5.8230 36.9370 5.8410 38.0960 ;
        RECT 4.4190 36.9730 4.5090 38.0870 ;
        RECT 3.7710 36.9370 3.7890 38.0960 ;
        RECT 0.1170 36.9365 0.1350 38.0965 ;
        RECT 9.4770 38.0165 9.4950 39.1765 ;
        RECT 5.8230 38.0170 5.8410 39.1760 ;
        RECT 4.4190 38.0530 4.5090 39.1670 ;
        RECT 3.7710 38.0170 3.7890 39.1760 ;
        RECT 0.1170 38.0165 0.1350 39.1765 ;
        RECT 9.4770 39.0965 9.4950 40.2565 ;
        RECT 5.8230 39.0970 5.8410 40.2560 ;
        RECT 4.4190 39.1330 4.5090 40.2470 ;
        RECT 3.7710 39.0970 3.7890 40.2560 ;
        RECT 0.1170 39.0965 0.1350 40.2565 ;
        RECT 9.4770 40.1765 9.4950 41.3365 ;
        RECT 5.8230 40.1770 5.8410 41.3360 ;
        RECT 4.4190 40.2130 4.5090 41.3270 ;
        RECT 3.7710 40.1770 3.7890 41.3360 ;
        RECT 0.1170 40.1765 0.1350 41.3365 ;
        RECT 9.4770 41.2565 9.4950 42.4165 ;
        RECT 5.8230 41.2570 5.8410 42.4160 ;
        RECT 4.4190 41.2930 4.5090 42.4070 ;
        RECT 3.7710 41.2570 3.7890 42.4160 ;
        RECT 0.1170 41.2565 0.1350 42.4165 ;
        RECT 9.4770 42.3365 9.4950 43.4965 ;
        RECT 5.8230 42.3370 5.8410 43.4960 ;
        RECT 4.4190 42.3730 4.5090 43.4870 ;
        RECT 3.7710 42.3370 3.7890 43.4960 ;
        RECT 0.1170 42.3365 0.1350 43.4965 ;
        RECT 9.4770 43.4165 9.4950 51.6235 ;
        RECT 5.8230 43.4960 5.8410 43.5875 ;
        RECT 5.8230 47.2360 5.8410 51.5960 ;
        RECT 4.4550 43.7400 4.6890 51.3230 ;
        RECT 4.4190 51.2370 4.5090 51.7720 ;
        RECT 4.4190 43.4600 4.5090 43.9950 ;
        RECT 0.1170 43.4165 0.1350 51.6235 ;
        RECT 9.4770 51.5435 9.4950 52.7035 ;
        RECT 5.8230 51.5440 5.8410 52.7030 ;
        RECT 4.4190 51.5800 4.5090 52.6940 ;
        RECT 3.7710 51.5440 3.7890 52.7030 ;
        RECT 0.1170 51.5435 0.1350 52.7035 ;
        RECT 9.4770 52.6235 9.4950 53.7835 ;
        RECT 5.8230 52.6240 5.8410 53.7830 ;
        RECT 4.4190 52.6600 4.5090 53.7740 ;
        RECT 3.7710 52.6240 3.7890 53.7830 ;
        RECT 0.1170 52.6235 0.1350 53.7835 ;
        RECT 9.4770 53.7035 9.4950 54.8635 ;
        RECT 5.8230 53.7040 5.8410 54.8630 ;
        RECT 4.4190 53.7400 4.5090 54.8540 ;
        RECT 3.7710 53.7040 3.7890 54.8630 ;
        RECT 0.1170 53.7035 0.1350 54.8635 ;
        RECT 9.4770 54.7835 9.4950 55.9435 ;
        RECT 5.8230 54.7840 5.8410 55.9430 ;
        RECT 4.4190 54.8200 4.5090 55.9340 ;
        RECT 3.7710 54.7840 3.7890 55.9430 ;
        RECT 0.1170 54.7835 0.1350 55.9435 ;
        RECT 9.4770 55.8635 9.4950 57.0235 ;
        RECT 5.8230 55.8640 5.8410 57.0230 ;
        RECT 4.4190 55.9000 4.5090 57.0140 ;
        RECT 3.7710 55.8640 3.7890 57.0230 ;
        RECT 0.1170 55.8635 0.1350 57.0235 ;
        RECT 9.4770 56.9435 9.4950 58.1035 ;
        RECT 5.8230 56.9440 5.8410 58.1030 ;
        RECT 4.4190 56.9800 4.5090 58.0940 ;
        RECT 3.7710 56.9440 3.7890 58.1030 ;
        RECT 0.1170 56.9435 0.1350 58.1035 ;
        RECT 9.4770 58.0235 9.4950 59.1835 ;
        RECT 5.8230 58.0240 5.8410 59.1830 ;
        RECT 4.4190 58.0600 4.5090 59.1740 ;
        RECT 3.7710 58.0240 3.7890 59.1830 ;
        RECT 0.1170 58.0235 0.1350 59.1835 ;
        RECT 9.4770 59.1035 9.4950 60.2635 ;
        RECT 5.8230 59.1040 5.8410 60.2630 ;
        RECT 4.4190 59.1400 4.5090 60.2540 ;
        RECT 3.7710 59.1040 3.7890 60.2630 ;
        RECT 0.1170 59.1035 0.1350 60.2635 ;
        RECT 9.4770 60.1835 9.4950 61.3435 ;
        RECT 5.8230 60.1840 5.8410 61.3430 ;
        RECT 4.4190 60.2200 4.5090 61.3340 ;
        RECT 3.7710 60.1840 3.7890 61.3430 ;
        RECT 0.1170 60.1835 0.1350 61.3435 ;
        RECT 9.4770 61.2635 9.4950 62.4235 ;
        RECT 5.8230 61.2640 5.8410 62.4230 ;
        RECT 4.4190 61.3000 4.5090 62.4140 ;
        RECT 3.7710 61.2640 3.7890 62.4230 ;
        RECT 0.1170 61.2635 0.1350 62.4235 ;
        RECT 9.4770 62.3435 9.4950 63.5035 ;
        RECT 5.8230 62.3440 5.8410 63.5030 ;
        RECT 4.4190 62.3800 4.5090 63.4940 ;
        RECT 3.7710 62.3440 3.7890 63.5030 ;
        RECT 0.1170 62.3435 0.1350 63.5035 ;
        RECT 9.4770 63.4235 9.4950 64.5835 ;
        RECT 5.8230 63.4240 5.8410 64.5830 ;
        RECT 4.4190 63.4600 4.5090 64.5740 ;
        RECT 3.7710 63.4240 3.7890 64.5830 ;
        RECT 0.1170 63.4235 0.1350 64.5835 ;
        RECT 9.4770 64.5035 9.4950 65.6635 ;
        RECT 5.8230 64.5040 5.8410 65.6630 ;
        RECT 4.4190 64.5400 4.5090 65.6540 ;
        RECT 3.7710 64.5040 3.7890 65.6630 ;
        RECT 0.1170 64.5035 0.1350 65.6635 ;
        RECT 9.4770 65.5835 9.4950 66.7435 ;
        RECT 5.8230 65.5840 5.8410 66.7430 ;
        RECT 4.4190 65.6200 4.5090 66.7340 ;
        RECT 3.7710 65.5840 3.7890 66.7430 ;
        RECT 0.1170 65.5835 0.1350 66.7435 ;
        RECT 9.4770 66.6635 9.4950 67.8235 ;
        RECT 5.8230 66.6640 5.8410 67.8230 ;
        RECT 4.4190 66.7000 4.5090 67.8140 ;
        RECT 3.7710 66.6640 3.7890 67.8230 ;
        RECT 0.1170 66.6635 0.1350 67.8235 ;
        RECT 9.4770 67.7435 9.4950 68.9035 ;
        RECT 5.8230 67.7440 5.8410 68.9030 ;
        RECT 4.4190 67.7800 4.5090 68.8940 ;
        RECT 3.7710 67.7440 3.7890 68.9030 ;
        RECT 0.1170 67.7435 0.1350 68.9035 ;
        RECT 9.4770 68.8235 9.4950 69.9835 ;
        RECT 5.8230 68.8240 5.8410 69.9830 ;
        RECT 4.4190 68.8600 4.5090 69.9740 ;
        RECT 3.7710 68.8240 3.7890 69.9830 ;
        RECT 0.1170 68.8235 0.1350 69.9835 ;
        RECT 9.4770 69.9035 9.4950 71.0635 ;
        RECT 5.8230 69.9040 5.8410 71.0630 ;
        RECT 4.4190 69.9400 4.5090 71.0540 ;
        RECT 3.7710 69.9040 3.7890 71.0630 ;
        RECT 0.1170 69.9035 0.1350 71.0635 ;
        RECT 9.4770 70.9835 9.4950 72.1435 ;
        RECT 5.8230 70.9840 5.8410 72.1430 ;
        RECT 4.4190 71.0200 4.5090 72.1340 ;
        RECT 3.7710 70.9840 3.7890 72.1430 ;
        RECT 0.1170 70.9835 0.1350 72.1435 ;
        RECT 9.4770 72.0635 9.4950 73.2235 ;
        RECT 5.8230 72.0640 5.8410 73.2230 ;
        RECT 4.4190 72.1000 4.5090 73.2140 ;
        RECT 3.7710 72.0640 3.7890 73.2230 ;
        RECT 0.1170 72.0635 0.1350 73.2235 ;
        RECT 9.4770 73.1435 9.4950 74.3035 ;
        RECT 5.8230 73.1440 5.8410 74.3030 ;
        RECT 4.4190 73.1800 4.5090 74.2940 ;
        RECT 3.7710 73.1440 3.7890 74.3030 ;
        RECT 0.1170 73.1435 0.1350 74.3035 ;
        RECT 9.4770 74.2235 9.4950 75.3835 ;
        RECT 5.8230 74.2240 5.8410 75.3830 ;
        RECT 4.4190 74.2600 4.5090 75.3740 ;
        RECT 3.7710 74.2240 3.7890 75.3830 ;
        RECT 0.1170 74.2235 0.1350 75.3835 ;
        RECT 9.4770 75.3035 9.4950 76.4635 ;
        RECT 5.8230 75.3040 5.8410 76.4630 ;
        RECT 4.4190 75.3400 4.5090 76.4540 ;
        RECT 3.7710 75.3040 3.7890 76.4630 ;
        RECT 0.1170 75.3035 0.1350 76.4635 ;
        RECT 9.4770 76.3835 9.4950 77.5435 ;
        RECT 5.8230 76.3840 5.8410 77.5430 ;
        RECT 4.4190 76.4200 4.5090 77.5340 ;
        RECT 3.7710 76.3840 3.7890 77.5430 ;
        RECT 0.1170 76.3835 0.1350 77.5435 ;
        RECT 9.4770 77.4635 9.4950 78.6235 ;
        RECT 5.8230 77.4640 5.8410 78.6230 ;
        RECT 4.4190 77.5000 4.5090 78.6140 ;
        RECT 3.7710 77.4640 3.7890 78.6230 ;
        RECT 0.1170 77.4635 0.1350 78.6235 ;
        RECT 9.4770 78.5435 9.4950 79.7035 ;
        RECT 5.8230 78.5440 5.8410 79.7030 ;
        RECT 4.4190 78.5800 4.5090 79.6940 ;
        RECT 3.7710 78.5440 3.7890 79.7030 ;
        RECT 0.1170 78.5435 0.1350 79.7035 ;
        RECT 9.4770 79.6235 9.4950 80.7835 ;
        RECT 5.8230 79.6240 5.8410 80.7830 ;
        RECT 4.4190 79.6600 4.5090 80.7740 ;
        RECT 3.7710 79.6240 3.7890 80.7830 ;
        RECT 0.1170 79.6235 0.1350 80.7835 ;
        RECT 9.4770 80.7035 9.4950 81.8635 ;
        RECT 5.8230 80.7040 5.8410 81.8630 ;
        RECT 4.4190 80.7400 4.5090 81.8540 ;
        RECT 3.7710 80.7040 3.7890 81.8630 ;
        RECT 0.1170 80.7035 0.1350 81.8635 ;
        RECT 9.4770 81.7835 9.4950 82.9435 ;
        RECT 5.8230 81.7840 5.8410 82.9430 ;
        RECT 4.4190 81.8200 4.5090 82.9340 ;
        RECT 3.7710 81.7840 3.7890 82.9430 ;
        RECT 0.1170 81.7835 0.1350 82.9435 ;
        RECT 9.4770 82.8635 9.4950 84.0235 ;
        RECT 5.8230 82.8640 5.8410 84.0230 ;
        RECT 4.4190 82.9000 4.5090 84.0140 ;
        RECT 3.7710 82.8640 3.7890 84.0230 ;
        RECT 0.1170 82.8635 0.1350 84.0235 ;
        RECT 9.4770 83.9435 9.4950 85.1035 ;
        RECT 5.8230 83.9440 5.8410 85.1030 ;
        RECT 4.4190 83.9800 4.5090 85.0940 ;
        RECT 3.7710 83.9440 3.7890 85.1030 ;
        RECT 0.1170 83.9435 0.1350 85.1035 ;
        RECT 9.4770 85.0235 9.4950 86.1835 ;
        RECT 5.8230 85.0240 5.8410 86.1830 ;
        RECT 4.4190 85.0600 4.5090 86.1740 ;
        RECT 3.7710 85.0240 3.7890 86.1830 ;
        RECT 0.1170 85.0235 0.1350 86.1835 ;
        RECT 9.4770 86.1035 9.4950 87.2635 ;
        RECT 5.8230 86.1040 5.8410 87.2630 ;
        RECT 4.4190 86.1400 4.5090 87.2540 ;
        RECT 3.7710 86.1040 3.7890 87.2630 ;
        RECT 0.1170 86.1035 0.1350 87.2635 ;
        RECT 9.4770 87.1835 9.4950 88.3435 ;
        RECT 5.8230 87.1840 5.8410 88.3430 ;
        RECT 4.4190 87.2200 4.5090 88.3340 ;
        RECT 3.7710 87.1840 3.7890 88.3430 ;
        RECT 0.1170 87.1835 0.1350 88.3435 ;
        RECT 9.4770 88.2635 9.4950 89.4235 ;
        RECT 5.8230 88.2640 5.8410 89.4230 ;
        RECT 4.4190 88.3000 4.5090 89.4140 ;
        RECT 3.7710 88.2640 3.7890 89.4230 ;
        RECT 0.1170 88.2635 0.1350 89.4235 ;
        RECT 9.4770 89.3435 9.4950 90.5035 ;
        RECT 5.8230 89.3440 5.8410 90.5030 ;
        RECT 4.4190 89.3800 4.5090 90.4940 ;
        RECT 3.7710 89.3440 3.7890 90.5030 ;
        RECT 0.1170 89.3435 0.1350 90.5035 ;
        RECT 9.4770 90.4235 9.4950 91.5835 ;
        RECT 5.8230 90.4240 5.8410 91.5830 ;
        RECT 4.4190 90.4600 4.5090 91.5740 ;
        RECT 3.7710 90.4240 3.7890 91.5830 ;
        RECT 0.1170 90.4235 0.1350 91.5835 ;
        RECT 9.4770 91.5035 9.4950 92.6635 ;
        RECT 5.8230 91.5040 5.8410 92.6630 ;
        RECT 4.4190 91.5400 4.5090 92.6540 ;
        RECT 3.7710 91.5040 3.7890 92.6630 ;
        RECT 0.1170 91.5035 0.1350 92.6635 ;
        RECT 9.4770 92.5835 9.4950 93.7435 ;
        RECT 5.8230 92.5840 5.8410 93.7430 ;
        RECT 4.4190 92.6200 4.5090 93.7340 ;
        RECT 3.7710 92.5840 3.7890 93.7430 ;
        RECT 0.1170 92.5835 0.1350 93.7435 ;
        RECT 9.4770 93.6635 9.4950 94.8235 ;
        RECT 5.8230 93.6640 5.8410 94.8230 ;
        RECT 4.4190 93.7000 4.5090 94.8140 ;
        RECT 3.7710 93.6640 3.7890 94.8230 ;
        RECT 0.1170 93.6635 0.1350 94.8235 ;
      LAYER V3  ;
        RECT 0.1170 1.1720 0.1350 1.2200 ;
        RECT 3.7710 1.1720 3.7890 1.2200 ;
        RECT 4.4190 1.1720 4.5090 1.2200 ;
        RECT 5.8230 1.1720 5.8410 1.2200 ;
        RECT 9.4770 1.1720 9.4950 1.2200 ;
        RECT 0.1170 2.2520 0.1350 2.3000 ;
        RECT 3.7710 2.2520 3.7890 2.3000 ;
        RECT 4.4190 2.2520 4.5090 2.3000 ;
        RECT 5.8230 2.2520 5.8410 2.3000 ;
        RECT 9.4770 2.2520 9.4950 2.3000 ;
        RECT 0.1170 3.3320 0.1350 3.3800 ;
        RECT 3.7710 3.3320 3.7890 3.3800 ;
        RECT 4.4190 3.3320 4.5090 3.3800 ;
        RECT 5.8230 3.3320 5.8410 3.3800 ;
        RECT 9.4770 3.3320 9.4950 3.3800 ;
        RECT 0.1170 4.4120 0.1350 4.4600 ;
        RECT 3.7710 4.4120 3.7890 4.4600 ;
        RECT 4.4190 4.4120 4.5090 4.4600 ;
        RECT 5.8230 4.4120 5.8410 4.4600 ;
        RECT 9.4770 4.4120 9.4950 4.4600 ;
        RECT 0.1170 5.4920 0.1350 5.5400 ;
        RECT 3.7710 5.4920 3.7890 5.5400 ;
        RECT 4.4190 5.4920 4.5090 5.5400 ;
        RECT 5.8230 5.4920 5.8410 5.5400 ;
        RECT 9.4770 5.4920 9.4950 5.5400 ;
        RECT 0.1170 6.5720 0.1350 6.6200 ;
        RECT 3.7710 6.5720 3.7890 6.6200 ;
        RECT 4.4190 6.5720 4.5090 6.6200 ;
        RECT 5.8230 6.5720 5.8410 6.6200 ;
        RECT 9.4770 6.5720 9.4950 6.6200 ;
        RECT 0.1170 7.6520 0.1350 7.7000 ;
        RECT 3.7710 7.6520 3.7890 7.7000 ;
        RECT 4.4190 7.6520 4.5090 7.7000 ;
        RECT 5.8230 7.6520 5.8410 7.7000 ;
        RECT 9.4770 7.6520 9.4950 7.7000 ;
        RECT 0.1170 8.7320 0.1350 8.7800 ;
        RECT 3.7710 8.7320 3.7890 8.7800 ;
        RECT 4.4190 8.7320 4.5090 8.7800 ;
        RECT 5.8230 8.7320 5.8410 8.7800 ;
        RECT 9.4770 8.7320 9.4950 8.7800 ;
        RECT 0.1170 9.8120 0.1350 9.8600 ;
        RECT 3.7710 9.8120 3.7890 9.8600 ;
        RECT 4.4190 9.8120 4.5090 9.8600 ;
        RECT 5.8230 9.8120 5.8410 9.8600 ;
        RECT 9.4770 9.8120 9.4950 9.8600 ;
        RECT 0.1170 10.8920 0.1350 10.9400 ;
        RECT 3.7710 10.8920 3.7890 10.9400 ;
        RECT 4.4190 10.8920 4.5090 10.9400 ;
        RECT 5.8230 10.8920 5.8410 10.9400 ;
        RECT 9.4770 10.8920 9.4950 10.9400 ;
        RECT 0.1170 11.9720 0.1350 12.0200 ;
        RECT 3.7710 11.9720 3.7890 12.0200 ;
        RECT 4.4190 11.9720 4.5090 12.0200 ;
        RECT 5.8230 11.9720 5.8410 12.0200 ;
        RECT 9.4770 11.9720 9.4950 12.0200 ;
        RECT 0.1170 13.0520 0.1350 13.1000 ;
        RECT 3.7710 13.0520 3.7890 13.1000 ;
        RECT 4.4190 13.0520 4.5090 13.1000 ;
        RECT 5.8230 13.0520 5.8410 13.1000 ;
        RECT 9.4770 13.0520 9.4950 13.1000 ;
        RECT 0.1170 14.1320 0.1350 14.1800 ;
        RECT 3.7710 14.1320 3.7890 14.1800 ;
        RECT 4.4190 14.1320 4.5090 14.1800 ;
        RECT 5.8230 14.1320 5.8410 14.1800 ;
        RECT 9.4770 14.1320 9.4950 14.1800 ;
        RECT 0.1170 15.2120 0.1350 15.2600 ;
        RECT 3.7710 15.2120 3.7890 15.2600 ;
        RECT 4.4190 15.2120 4.5090 15.2600 ;
        RECT 5.8230 15.2120 5.8410 15.2600 ;
        RECT 9.4770 15.2120 9.4950 15.2600 ;
        RECT 0.1170 16.2920 0.1350 16.3400 ;
        RECT 3.7710 16.2920 3.7890 16.3400 ;
        RECT 4.4190 16.2920 4.5090 16.3400 ;
        RECT 5.8230 16.2920 5.8410 16.3400 ;
        RECT 9.4770 16.2920 9.4950 16.3400 ;
        RECT 0.1170 17.3720 0.1350 17.4200 ;
        RECT 3.7710 17.3720 3.7890 17.4200 ;
        RECT 4.4190 17.3720 4.5090 17.4200 ;
        RECT 5.8230 17.3720 5.8410 17.4200 ;
        RECT 9.4770 17.3720 9.4950 17.4200 ;
        RECT 0.1170 18.4520 0.1350 18.5000 ;
        RECT 3.7710 18.4520 3.7890 18.5000 ;
        RECT 4.4190 18.4520 4.5090 18.5000 ;
        RECT 5.8230 18.4520 5.8410 18.5000 ;
        RECT 9.4770 18.4520 9.4950 18.5000 ;
        RECT 0.1170 19.5320 0.1350 19.5800 ;
        RECT 3.7710 19.5320 3.7890 19.5800 ;
        RECT 4.4190 19.5320 4.5090 19.5800 ;
        RECT 5.8230 19.5320 5.8410 19.5800 ;
        RECT 9.4770 19.5320 9.4950 19.5800 ;
        RECT 0.1170 20.6120 0.1350 20.6600 ;
        RECT 3.7710 20.6120 3.7890 20.6600 ;
        RECT 4.4190 20.6120 4.5090 20.6600 ;
        RECT 5.8230 20.6120 5.8410 20.6600 ;
        RECT 9.4770 20.6120 9.4950 20.6600 ;
        RECT 0.1170 21.6920 0.1350 21.7400 ;
        RECT 3.7710 21.6920 3.7890 21.7400 ;
        RECT 4.4190 21.6920 4.5090 21.7400 ;
        RECT 5.8230 21.6920 5.8410 21.7400 ;
        RECT 9.4770 21.6920 9.4950 21.7400 ;
        RECT 0.1170 22.7720 0.1350 22.8200 ;
        RECT 3.7710 22.7720 3.7890 22.8200 ;
        RECT 4.4190 22.7720 4.5090 22.8200 ;
        RECT 5.8230 22.7720 5.8410 22.8200 ;
        RECT 9.4770 22.7720 9.4950 22.8200 ;
        RECT 0.1170 23.8520 0.1350 23.9000 ;
        RECT 3.7710 23.8520 3.7890 23.9000 ;
        RECT 4.4190 23.8520 4.5090 23.9000 ;
        RECT 5.8230 23.8520 5.8410 23.9000 ;
        RECT 9.4770 23.8520 9.4950 23.9000 ;
        RECT 0.1170 24.9320 0.1350 24.9800 ;
        RECT 3.7710 24.9320 3.7890 24.9800 ;
        RECT 4.4190 24.9320 4.5090 24.9800 ;
        RECT 5.8230 24.9320 5.8410 24.9800 ;
        RECT 9.4770 24.9320 9.4950 24.9800 ;
        RECT 0.1170 26.0120 0.1350 26.0600 ;
        RECT 3.7710 26.0120 3.7890 26.0600 ;
        RECT 4.4190 26.0120 4.5090 26.0600 ;
        RECT 5.8230 26.0120 5.8410 26.0600 ;
        RECT 9.4770 26.0120 9.4950 26.0600 ;
        RECT 0.1170 27.0920 0.1350 27.1400 ;
        RECT 3.7710 27.0920 3.7890 27.1400 ;
        RECT 4.4190 27.0920 4.5090 27.1400 ;
        RECT 5.8230 27.0920 5.8410 27.1400 ;
        RECT 9.4770 27.0920 9.4950 27.1400 ;
        RECT 0.1170 28.1720 0.1350 28.2200 ;
        RECT 3.7710 28.1720 3.7890 28.2200 ;
        RECT 4.4190 28.1720 4.5090 28.2200 ;
        RECT 5.8230 28.1720 5.8410 28.2200 ;
        RECT 9.4770 28.1720 9.4950 28.2200 ;
        RECT 0.1170 29.2520 0.1350 29.3000 ;
        RECT 3.7710 29.2520 3.7890 29.3000 ;
        RECT 4.4190 29.2520 4.5090 29.3000 ;
        RECT 5.8230 29.2520 5.8410 29.3000 ;
        RECT 9.4770 29.2520 9.4950 29.3000 ;
        RECT 0.1170 30.3320 0.1350 30.3800 ;
        RECT 3.7710 30.3320 3.7890 30.3800 ;
        RECT 4.4190 30.3320 4.5090 30.3800 ;
        RECT 5.8230 30.3320 5.8410 30.3800 ;
        RECT 9.4770 30.3320 9.4950 30.3800 ;
        RECT 0.1170 31.4120 0.1350 31.4600 ;
        RECT 3.7710 31.4120 3.7890 31.4600 ;
        RECT 4.4190 31.4120 4.5090 31.4600 ;
        RECT 5.8230 31.4120 5.8410 31.4600 ;
        RECT 9.4770 31.4120 9.4950 31.4600 ;
        RECT 0.1170 32.4920 0.1350 32.5400 ;
        RECT 3.7710 32.4920 3.7890 32.5400 ;
        RECT 4.4190 32.4920 4.5090 32.5400 ;
        RECT 5.8230 32.4920 5.8410 32.5400 ;
        RECT 9.4770 32.4920 9.4950 32.5400 ;
        RECT 0.1170 33.5720 0.1350 33.6200 ;
        RECT 3.7710 33.5720 3.7890 33.6200 ;
        RECT 4.4190 33.5720 4.5090 33.6200 ;
        RECT 5.8230 33.5720 5.8410 33.6200 ;
        RECT 9.4770 33.5720 9.4950 33.6200 ;
        RECT 0.1170 34.6520 0.1350 34.7000 ;
        RECT 3.7710 34.6520 3.7890 34.7000 ;
        RECT 4.4190 34.6520 4.5090 34.7000 ;
        RECT 5.8230 34.6520 5.8410 34.7000 ;
        RECT 9.4770 34.6520 9.4950 34.7000 ;
        RECT 0.1170 35.7320 0.1350 35.7800 ;
        RECT 3.7710 35.7320 3.7890 35.7800 ;
        RECT 4.4190 35.7320 4.5090 35.7800 ;
        RECT 5.8230 35.7320 5.8410 35.7800 ;
        RECT 9.4770 35.7320 9.4950 35.7800 ;
        RECT 0.1170 36.8120 0.1350 36.8600 ;
        RECT 3.7710 36.8120 3.7890 36.8600 ;
        RECT 4.4190 36.8120 4.5090 36.8600 ;
        RECT 5.8230 36.8120 5.8410 36.8600 ;
        RECT 9.4770 36.8120 9.4950 36.8600 ;
        RECT 0.1170 37.8920 0.1350 37.9400 ;
        RECT 3.7710 37.8920 3.7890 37.9400 ;
        RECT 4.4190 37.8920 4.5090 37.9400 ;
        RECT 5.8230 37.8920 5.8410 37.9400 ;
        RECT 9.4770 37.8920 9.4950 37.9400 ;
        RECT 0.1170 38.9720 0.1350 39.0200 ;
        RECT 3.7710 38.9720 3.7890 39.0200 ;
        RECT 4.4190 38.9720 4.5090 39.0200 ;
        RECT 5.8230 38.9720 5.8410 39.0200 ;
        RECT 9.4770 38.9720 9.4950 39.0200 ;
        RECT 0.1170 40.0520 0.1350 40.1000 ;
        RECT 3.7710 40.0520 3.7890 40.1000 ;
        RECT 4.4190 40.0520 4.5090 40.1000 ;
        RECT 5.8230 40.0520 5.8410 40.1000 ;
        RECT 9.4770 40.0520 9.4950 40.1000 ;
        RECT 0.1170 41.1320 0.1350 41.1800 ;
        RECT 3.7710 41.1320 3.7890 41.1800 ;
        RECT 4.4190 41.1320 4.5090 41.1800 ;
        RECT 5.8230 41.1320 5.8410 41.1800 ;
        RECT 9.4770 41.1320 9.4950 41.1800 ;
        RECT 0.1170 42.2120 0.1350 42.2600 ;
        RECT 3.7710 42.2120 3.7890 42.2600 ;
        RECT 4.4190 42.2120 4.5090 42.2600 ;
        RECT 5.8230 42.2120 5.8410 42.2600 ;
        RECT 9.4770 42.2120 9.4950 42.2600 ;
        RECT 0.1170 43.2920 0.1350 43.3400 ;
        RECT 3.7710 43.2920 3.7890 43.3400 ;
        RECT 4.4190 43.2920 4.5090 43.3400 ;
        RECT 5.8230 43.2920 5.8410 43.3400 ;
        RECT 9.4770 43.2920 9.4950 43.3400 ;
        RECT 0.1170 43.7790 0.1350 43.9950 ;
        RECT 4.4590 50.1150 4.4770 50.3310 ;
        RECT 4.4590 46.9470 4.4770 47.1630 ;
        RECT 4.4590 43.7790 4.4770 43.9950 ;
        RECT 4.5110 50.1150 4.5290 50.3310 ;
        RECT 4.5110 46.9470 4.5290 47.1630 ;
        RECT 4.5110 43.7790 4.5290 43.9950 ;
        RECT 4.5630 50.1150 4.5810 50.3310 ;
        RECT 4.5630 46.9470 4.5810 47.1630 ;
        RECT 4.5630 43.7790 4.5810 43.9950 ;
        RECT 4.6150 50.1150 4.6330 50.3310 ;
        RECT 4.6150 46.9470 4.6330 47.1630 ;
        RECT 4.6150 43.7790 4.6330 43.9950 ;
        RECT 4.6670 50.1150 4.6850 50.3310 ;
        RECT 4.6670 46.9470 4.6850 47.1630 ;
        RECT 4.6670 43.7790 4.6850 43.9950 ;
        RECT 5.8230 47.2830 5.8410 47.3070 ;
        RECT 5.8230 43.4990 5.8410 43.5230 ;
        RECT 0.1170 52.4990 0.1350 52.5470 ;
        RECT 3.7710 52.4990 3.7890 52.5470 ;
        RECT 4.4190 52.4990 4.5090 52.5470 ;
        RECT 5.8230 52.4990 5.8410 52.5470 ;
        RECT 9.4770 52.4990 9.4950 52.5470 ;
        RECT 0.1170 53.5790 0.1350 53.6270 ;
        RECT 3.7710 53.5790 3.7890 53.6270 ;
        RECT 4.4190 53.5790 4.5090 53.6270 ;
        RECT 5.8230 53.5790 5.8410 53.6270 ;
        RECT 9.4770 53.5790 9.4950 53.6270 ;
        RECT 0.1170 54.6590 0.1350 54.7070 ;
        RECT 3.7710 54.6590 3.7890 54.7070 ;
        RECT 4.4190 54.6590 4.5090 54.7070 ;
        RECT 5.8230 54.6590 5.8410 54.7070 ;
        RECT 9.4770 54.6590 9.4950 54.7070 ;
        RECT 0.1170 55.7390 0.1350 55.7870 ;
        RECT 3.7710 55.7390 3.7890 55.7870 ;
        RECT 4.4190 55.7390 4.5090 55.7870 ;
        RECT 5.8230 55.7390 5.8410 55.7870 ;
        RECT 9.4770 55.7390 9.4950 55.7870 ;
        RECT 0.1170 56.8190 0.1350 56.8670 ;
        RECT 3.7710 56.8190 3.7890 56.8670 ;
        RECT 4.4190 56.8190 4.5090 56.8670 ;
        RECT 5.8230 56.8190 5.8410 56.8670 ;
        RECT 9.4770 56.8190 9.4950 56.8670 ;
        RECT 0.1170 57.8990 0.1350 57.9470 ;
        RECT 3.7710 57.8990 3.7890 57.9470 ;
        RECT 4.4190 57.8990 4.5090 57.9470 ;
        RECT 5.8230 57.8990 5.8410 57.9470 ;
        RECT 9.4770 57.8990 9.4950 57.9470 ;
        RECT 0.1170 58.9790 0.1350 59.0270 ;
        RECT 3.7710 58.9790 3.7890 59.0270 ;
        RECT 4.4190 58.9790 4.5090 59.0270 ;
        RECT 5.8230 58.9790 5.8410 59.0270 ;
        RECT 9.4770 58.9790 9.4950 59.0270 ;
        RECT 0.1170 60.0590 0.1350 60.1070 ;
        RECT 3.7710 60.0590 3.7890 60.1070 ;
        RECT 4.4190 60.0590 4.5090 60.1070 ;
        RECT 5.8230 60.0590 5.8410 60.1070 ;
        RECT 9.4770 60.0590 9.4950 60.1070 ;
        RECT 0.1170 61.1390 0.1350 61.1870 ;
        RECT 3.7710 61.1390 3.7890 61.1870 ;
        RECT 4.4190 61.1390 4.5090 61.1870 ;
        RECT 5.8230 61.1390 5.8410 61.1870 ;
        RECT 9.4770 61.1390 9.4950 61.1870 ;
        RECT 0.1170 62.2190 0.1350 62.2670 ;
        RECT 3.7710 62.2190 3.7890 62.2670 ;
        RECT 4.4190 62.2190 4.5090 62.2670 ;
        RECT 5.8230 62.2190 5.8410 62.2670 ;
        RECT 9.4770 62.2190 9.4950 62.2670 ;
        RECT 0.1170 63.2990 0.1350 63.3470 ;
        RECT 3.7710 63.2990 3.7890 63.3470 ;
        RECT 4.4190 63.2990 4.5090 63.3470 ;
        RECT 5.8230 63.2990 5.8410 63.3470 ;
        RECT 9.4770 63.2990 9.4950 63.3470 ;
        RECT 0.1170 64.3790 0.1350 64.4270 ;
        RECT 3.7710 64.3790 3.7890 64.4270 ;
        RECT 4.4190 64.3790 4.5090 64.4270 ;
        RECT 5.8230 64.3790 5.8410 64.4270 ;
        RECT 9.4770 64.3790 9.4950 64.4270 ;
        RECT 0.1170 65.4590 0.1350 65.5070 ;
        RECT 3.7710 65.4590 3.7890 65.5070 ;
        RECT 4.4190 65.4590 4.5090 65.5070 ;
        RECT 5.8230 65.4590 5.8410 65.5070 ;
        RECT 9.4770 65.4590 9.4950 65.5070 ;
        RECT 0.1170 66.5390 0.1350 66.5870 ;
        RECT 3.7710 66.5390 3.7890 66.5870 ;
        RECT 4.4190 66.5390 4.5090 66.5870 ;
        RECT 5.8230 66.5390 5.8410 66.5870 ;
        RECT 9.4770 66.5390 9.4950 66.5870 ;
        RECT 0.1170 67.6190 0.1350 67.6670 ;
        RECT 3.7710 67.6190 3.7890 67.6670 ;
        RECT 4.4190 67.6190 4.5090 67.6670 ;
        RECT 5.8230 67.6190 5.8410 67.6670 ;
        RECT 9.4770 67.6190 9.4950 67.6670 ;
        RECT 0.1170 68.6990 0.1350 68.7470 ;
        RECT 3.7710 68.6990 3.7890 68.7470 ;
        RECT 4.4190 68.6990 4.5090 68.7470 ;
        RECT 5.8230 68.6990 5.8410 68.7470 ;
        RECT 9.4770 68.6990 9.4950 68.7470 ;
        RECT 0.1170 69.7790 0.1350 69.8270 ;
        RECT 3.7710 69.7790 3.7890 69.8270 ;
        RECT 4.4190 69.7790 4.5090 69.8270 ;
        RECT 5.8230 69.7790 5.8410 69.8270 ;
        RECT 9.4770 69.7790 9.4950 69.8270 ;
        RECT 0.1170 70.8590 0.1350 70.9070 ;
        RECT 3.7710 70.8590 3.7890 70.9070 ;
        RECT 4.4190 70.8590 4.5090 70.9070 ;
        RECT 5.8230 70.8590 5.8410 70.9070 ;
        RECT 9.4770 70.8590 9.4950 70.9070 ;
        RECT 0.1170 71.9390 0.1350 71.9870 ;
        RECT 3.7710 71.9390 3.7890 71.9870 ;
        RECT 4.4190 71.9390 4.5090 71.9870 ;
        RECT 5.8230 71.9390 5.8410 71.9870 ;
        RECT 9.4770 71.9390 9.4950 71.9870 ;
        RECT 0.1170 73.0190 0.1350 73.0670 ;
        RECT 3.7710 73.0190 3.7890 73.0670 ;
        RECT 4.4190 73.0190 4.5090 73.0670 ;
        RECT 5.8230 73.0190 5.8410 73.0670 ;
        RECT 9.4770 73.0190 9.4950 73.0670 ;
        RECT 0.1170 74.0990 0.1350 74.1470 ;
        RECT 3.7710 74.0990 3.7890 74.1470 ;
        RECT 4.4190 74.0990 4.5090 74.1470 ;
        RECT 5.8230 74.0990 5.8410 74.1470 ;
        RECT 9.4770 74.0990 9.4950 74.1470 ;
        RECT 0.1170 75.1790 0.1350 75.2270 ;
        RECT 3.7710 75.1790 3.7890 75.2270 ;
        RECT 4.4190 75.1790 4.5090 75.2270 ;
        RECT 5.8230 75.1790 5.8410 75.2270 ;
        RECT 9.4770 75.1790 9.4950 75.2270 ;
        RECT 0.1170 76.2590 0.1350 76.3070 ;
        RECT 3.7710 76.2590 3.7890 76.3070 ;
        RECT 4.4190 76.2590 4.5090 76.3070 ;
        RECT 5.8230 76.2590 5.8410 76.3070 ;
        RECT 9.4770 76.2590 9.4950 76.3070 ;
        RECT 0.1170 77.3390 0.1350 77.3870 ;
        RECT 3.7710 77.3390 3.7890 77.3870 ;
        RECT 4.4190 77.3390 4.5090 77.3870 ;
        RECT 5.8230 77.3390 5.8410 77.3870 ;
        RECT 9.4770 77.3390 9.4950 77.3870 ;
        RECT 0.1170 78.4190 0.1350 78.4670 ;
        RECT 3.7710 78.4190 3.7890 78.4670 ;
        RECT 4.4190 78.4190 4.5090 78.4670 ;
        RECT 5.8230 78.4190 5.8410 78.4670 ;
        RECT 9.4770 78.4190 9.4950 78.4670 ;
        RECT 0.1170 79.4990 0.1350 79.5470 ;
        RECT 3.7710 79.4990 3.7890 79.5470 ;
        RECT 4.4190 79.4990 4.5090 79.5470 ;
        RECT 5.8230 79.4990 5.8410 79.5470 ;
        RECT 9.4770 79.4990 9.4950 79.5470 ;
        RECT 0.1170 80.5790 0.1350 80.6270 ;
        RECT 3.7710 80.5790 3.7890 80.6270 ;
        RECT 4.4190 80.5790 4.5090 80.6270 ;
        RECT 5.8230 80.5790 5.8410 80.6270 ;
        RECT 9.4770 80.5790 9.4950 80.6270 ;
        RECT 0.1170 81.6590 0.1350 81.7070 ;
        RECT 3.7710 81.6590 3.7890 81.7070 ;
        RECT 4.4190 81.6590 4.5090 81.7070 ;
        RECT 5.8230 81.6590 5.8410 81.7070 ;
        RECT 9.4770 81.6590 9.4950 81.7070 ;
        RECT 0.1170 82.7390 0.1350 82.7870 ;
        RECT 3.7710 82.7390 3.7890 82.7870 ;
        RECT 4.4190 82.7390 4.5090 82.7870 ;
        RECT 5.8230 82.7390 5.8410 82.7870 ;
        RECT 9.4770 82.7390 9.4950 82.7870 ;
        RECT 0.1170 83.8190 0.1350 83.8670 ;
        RECT 3.7710 83.8190 3.7890 83.8670 ;
        RECT 4.4190 83.8190 4.5090 83.8670 ;
        RECT 5.8230 83.8190 5.8410 83.8670 ;
        RECT 9.4770 83.8190 9.4950 83.8670 ;
        RECT 0.1170 84.8990 0.1350 84.9470 ;
        RECT 3.7710 84.8990 3.7890 84.9470 ;
        RECT 4.4190 84.8990 4.5090 84.9470 ;
        RECT 5.8230 84.8990 5.8410 84.9470 ;
        RECT 9.4770 84.8990 9.4950 84.9470 ;
        RECT 0.1170 85.9790 0.1350 86.0270 ;
        RECT 3.7710 85.9790 3.7890 86.0270 ;
        RECT 4.4190 85.9790 4.5090 86.0270 ;
        RECT 5.8230 85.9790 5.8410 86.0270 ;
        RECT 9.4770 85.9790 9.4950 86.0270 ;
        RECT 0.1170 87.0590 0.1350 87.1070 ;
        RECT 3.7710 87.0590 3.7890 87.1070 ;
        RECT 4.4190 87.0590 4.5090 87.1070 ;
        RECT 5.8230 87.0590 5.8410 87.1070 ;
        RECT 9.4770 87.0590 9.4950 87.1070 ;
        RECT 0.1170 88.1390 0.1350 88.1870 ;
        RECT 3.7710 88.1390 3.7890 88.1870 ;
        RECT 4.4190 88.1390 4.5090 88.1870 ;
        RECT 5.8230 88.1390 5.8410 88.1870 ;
        RECT 9.4770 88.1390 9.4950 88.1870 ;
        RECT 0.1170 89.2190 0.1350 89.2670 ;
        RECT 3.7710 89.2190 3.7890 89.2670 ;
        RECT 4.4190 89.2190 4.5090 89.2670 ;
        RECT 5.8230 89.2190 5.8410 89.2670 ;
        RECT 9.4770 89.2190 9.4950 89.2670 ;
        RECT 0.1170 90.2990 0.1350 90.3470 ;
        RECT 3.7710 90.2990 3.7890 90.3470 ;
        RECT 4.4190 90.2990 4.5090 90.3470 ;
        RECT 5.8230 90.2990 5.8410 90.3470 ;
        RECT 9.4770 90.2990 9.4950 90.3470 ;
        RECT 0.1170 91.3790 0.1350 91.4270 ;
        RECT 3.7710 91.3790 3.7890 91.4270 ;
        RECT 4.4190 91.3790 4.5090 91.4270 ;
        RECT 5.8230 91.3790 5.8410 91.4270 ;
        RECT 9.4770 91.3790 9.4950 91.4270 ;
        RECT 0.1170 92.4590 0.1350 92.5070 ;
        RECT 3.7710 92.4590 3.7890 92.5070 ;
        RECT 4.4190 92.4590 4.5090 92.5070 ;
        RECT 5.8230 92.4590 5.8410 92.5070 ;
        RECT 9.4770 92.4590 9.4950 92.5070 ;
        RECT 0.1170 93.5390 0.1350 93.5870 ;
        RECT 3.7710 93.5390 3.7890 93.5870 ;
        RECT 4.4190 93.5390 4.5090 93.5870 ;
        RECT 5.8230 93.5390 5.8410 93.5870 ;
        RECT 9.4770 93.5390 9.4950 93.5870 ;
        RECT 0.1170 94.6190 0.1350 94.6670 ;
        RECT 3.7710 94.6190 3.7890 94.6670 ;
        RECT 4.4190 94.6190 4.5090 94.6670 ;
        RECT 5.8230 94.6190 5.8410 94.6670 ;
        RECT 9.4770 94.6190 9.4950 94.6670 ;
      LAYER M5  ;
        RECT 5.7590 43.4810 5.7830 47.3250 ;
      LAYER V4  ;
        RECT 5.7590 47.2830 5.7830 47.3070 ;
        RECT 5.7590 43.4990 5.7830 43.5230 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1010 1.0760 9.5040 1.1240 ;
        RECT 0.1010 2.1560 9.5040 2.2040 ;
        RECT 0.1010 3.2360 9.5040 3.2840 ;
        RECT 0.1010 4.3160 9.5040 4.3640 ;
        RECT 0.1010 5.3960 9.5040 5.4440 ;
        RECT 0.1010 6.4760 9.5040 6.5240 ;
        RECT 0.1010 7.5560 9.5040 7.6040 ;
        RECT 0.1010 8.6360 9.5040 8.6840 ;
        RECT 0.1010 9.7160 9.5040 9.7640 ;
        RECT 0.1010 10.7960 9.5040 10.8440 ;
        RECT 0.1010 11.8760 9.5040 11.9240 ;
        RECT 0.1010 12.9560 9.5040 13.0040 ;
        RECT 0.1010 14.0360 9.5040 14.0840 ;
        RECT 0.1010 15.1160 9.5040 15.1640 ;
        RECT 0.1010 16.1960 9.5040 16.2440 ;
        RECT 0.1010 17.2760 9.5040 17.3240 ;
        RECT 0.1010 18.3560 9.5040 18.4040 ;
        RECT 0.1010 19.4360 9.5040 19.4840 ;
        RECT 0.1010 20.5160 9.5040 20.5640 ;
        RECT 0.1010 21.5960 9.5040 21.6440 ;
        RECT 0.1010 22.6760 9.5040 22.7240 ;
        RECT 0.1010 23.7560 9.5040 23.8040 ;
        RECT 0.1010 24.8360 9.5040 24.8840 ;
        RECT 0.1010 25.9160 9.5040 25.9640 ;
        RECT 0.1010 26.9960 9.5040 27.0440 ;
        RECT 0.1010 28.0760 9.5040 28.1240 ;
        RECT 0.1010 29.1560 9.5040 29.2040 ;
        RECT 0.1010 30.2360 9.5040 30.2840 ;
        RECT 0.1010 31.3160 9.5040 31.3640 ;
        RECT 0.1010 32.3960 9.5040 32.4440 ;
        RECT 0.1010 33.4760 9.5040 33.5240 ;
        RECT 0.1010 34.5560 9.5040 34.6040 ;
        RECT 0.1010 35.6360 9.5040 35.6840 ;
        RECT 0.1010 36.7160 9.5040 36.7640 ;
        RECT 0.1010 37.7960 9.5040 37.8440 ;
        RECT 0.1010 38.8760 9.5040 38.9240 ;
        RECT 0.1010 39.9560 9.5040 40.0040 ;
        RECT 0.1010 41.0360 9.5040 41.0840 ;
        RECT 0.1010 42.1160 9.5040 42.1640 ;
        RECT 0.1010 43.1960 9.5040 43.2440 ;
        RECT 0.1080 44.2110 9.5040 44.4270 ;
        RECT 3.9420 47.3790 5.6700 47.5950 ;
        RECT 3.9420 50.5470 5.6700 50.7630 ;
        RECT 0.1010 52.4030 9.5040 52.4510 ;
        RECT 0.1010 53.4830 9.5040 53.5310 ;
        RECT 0.1010 54.5630 9.5040 54.6110 ;
        RECT 0.1010 55.6430 9.5040 55.6910 ;
        RECT 0.1010 56.7230 9.5040 56.7710 ;
        RECT 0.1010 57.8030 9.5040 57.8510 ;
        RECT 0.1010 58.8830 9.5040 58.9310 ;
        RECT 0.1010 59.9630 9.5040 60.0110 ;
        RECT 0.1010 61.0430 9.5040 61.0910 ;
        RECT 0.1010 62.1230 9.5040 62.1710 ;
        RECT 0.1010 63.2030 9.5040 63.2510 ;
        RECT 0.1010 64.2830 9.5040 64.3310 ;
        RECT 0.1010 65.3630 9.5040 65.4110 ;
        RECT 0.1010 66.4430 9.5040 66.4910 ;
        RECT 0.1010 67.5230 9.5040 67.5710 ;
        RECT 0.1010 68.6030 9.5040 68.6510 ;
        RECT 0.1010 69.6830 9.5040 69.7310 ;
        RECT 0.1010 70.7630 9.5040 70.8110 ;
        RECT 0.1010 71.8430 9.5040 71.8910 ;
        RECT 0.1010 72.9230 9.5040 72.9710 ;
        RECT 0.1010 74.0030 9.5040 74.0510 ;
        RECT 0.1010 75.0830 9.5040 75.1310 ;
        RECT 0.1010 76.1630 9.5040 76.2110 ;
        RECT 0.1010 77.2430 9.5040 77.2910 ;
        RECT 0.1010 78.3230 9.5040 78.3710 ;
        RECT 0.1010 79.4030 9.5040 79.4510 ;
        RECT 0.1010 80.4830 9.5040 80.5310 ;
        RECT 0.1010 81.5630 9.5040 81.6110 ;
        RECT 0.1010 82.6430 9.5040 82.6910 ;
        RECT 0.1010 83.7230 9.5040 83.7710 ;
        RECT 0.1010 84.8030 9.5040 84.8510 ;
        RECT 0.1010 85.8830 9.5040 85.9310 ;
        RECT 0.1010 86.9630 9.5040 87.0110 ;
        RECT 0.1010 88.0430 9.5040 88.0910 ;
        RECT 0.1010 89.1230 9.5040 89.1710 ;
        RECT 0.1010 90.2030 9.5040 90.2510 ;
        RECT 0.1010 91.2830 9.5040 91.3310 ;
        RECT 0.1010 92.3630 9.5040 92.4110 ;
        RECT 0.1010 93.4430 9.5040 93.4910 ;
        RECT 0.1010 94.5230 9.5040 94.5710 ;
      LAYER M3  ;
        RECT 9.4410 0.2165 9.4590 1.3765 ;
        RECT 5.8770 0.2165 5.8950 1.3765 ;
        RECT 5.1120 0.2530 5.1480 1.3670 ;
        RECT 4.9590 0.2530 4.9860 1.3670 ;
        RECT 3.7170 0.2165 3.7350 1.3765 ;
        RECT 0.1530 0.2165 0.1710 1.3765 ;
        RECT 9.4410 1.2965 9.4590 2.4565 ;
        RECT 5.8770 1.2965 5.8950 2.4565 ;
        RECT 5.1120 1.3330 5.1480 2.4470 ;
        RECT 4.9590 1.3330 4.9860 2.4470 ;
        RECT 3.7170 1.2965 3.7350 2.4565 ;
        RECT 0.1530 1.2965 0.1710 2.4565 ;
        RECT 9.4410 2.3765 9.4590 3.5365 ;
        RECT 5.8770 2.3765 5.8950 3.5365 ;
        RECT 5.1120 2.4130 5.1480 3.5270 ;
        RECT 4.9590 2.4130 4.9860 3.5270 ;
        RECT 3.7170 2.3765 3.7350 3.5365 ;
        RECT 0.1530 2.3765 0.1710 3.5365 ;
        RECT 9.4410 3.4565 9.4590 4.6165 ;
        RECT 5.8770 3.4565 5.8950 4.6165 ;
        RECT 5.1120 3.4930 5.1480 4.6070 ;
        RECT 4.9590 3.4930 4.9860 4.6070 ;
        RECT 3.7170 3.4565 3.7350 4.6165 ;
        RECT 0.1530 3.4565 0.1710 4.6165 ;
        RECT 9.4410 4.5365 9.4590 5.6965 ;
        RECT 5.8770 4.5365 5.8950 5.6965 ;
        RECT 5.1120 4.5730 5.1480 5.6870 ;
        RECT 4.9590 4.5730 4.9860 5.6870 ;
        RECT 3.7170 4.5365 3.7350 5.6965 ;
        RECT 0.1530 4.5365 0.1710 5.6965 ;
        RECT 9.4410 5.6165 9.4590 6.7765 ;
        RECT 5.8770 5.6165 5.8950 6.7765 ;
        RECT 5.1120 5.6530 5.1480 6.7670 ;
        RECT 4.9590 5.6530 4.9860 6.7670 ;
        RECT 3.7170 5.6165 3.7350 6.7765 ;
        RECT 0.1530 5.6165 0.1710 6.7765 ;
        RECT 9.4410 6.6965 9.4590 7.8565 ;
        RECT 5.8770 6.6965 5.8950 7.8565 ;
        RECT 5.1120 6.7330 5.1480 7.8470 ;
        RECT 4.9590 6.7330 4.9860 7.8470 ;
        RECT 3.7170 6.6965 3.7350 7.8565 ;
        RECT 0.1530 6.6965 0.1710 7.8565 ;
        RECT 9.4410 7.7765 9.4590 8.9365 ;
        RECT 5.8770 7.7765 5.8950 8.9365 ;
        RECT 5.1120 7.8130 5.1480 8.9270 ;
        RECT 4.9590 7.8130 4.9860 8.9270 ;
        RECT 3.7170 7.7765 3.7350 8.9365 ;
        RECT 0.1530 7.7765 0.1710 8.9365 ;
        RECT 9.4410 8.8565 9.4590 10.0165 ;
        RECT 5.8770 8.8565 5.8950 10.0165 ;
        RECT 5.1120 8.8930 5.1480 10.0070 ;
        RECT 4.9590 8.8930 4.9860 10.0070 ;
        RECT 3.7170 8.8565 3.7350 10.0165 ;
        RECT 0.1530 8.8565 0.1710 10.0165 ;
        RECT 9.4410 9.9365 9.4590 11.0965 ;
        RECT 5.8770 9.9365 5.8950 11.0965 ;
        RECT 5.1120 9.9730 5.1480 11.0870 ;
        RECT 4.9590 9.9730 4.9860 11.0870 ;
        RECT 3.7170 9.9365 3.7350 11.0965 ;
        RECT 0.1530 9.9365 0.1710 11.0965 ;
        RECT 9.4410 11.0165 9.4590 12.1765 ;
        RECT 5.8770 11.0165 5.8950 12.1765 ;
        RECT 5.1120 11.0530 5.1480 12.1670 ;
        RECT 4.9590 11.0530 4.9860 12.1670 ;
        RECT 3.7170 11.0165 3.7350 12.1765 ;
        RECT 0.1530 11.0165 0.1710 12.1765 ;
        RECT 9.4410 12.0965 9.4590 13.2565 ;
        RECT 5.8770 12.0965 5.8950 13.2565 ;
        RECT 5.1120 12.1330 5.1480 13.2470 ;
        RECT 4.9590 12.1330 4.9860 13.2470 ;
        RECT 3.7170 12.0965 3.7350 13.2565 ;
        RECT 0.1530 12.0965 0.1710 13.2565 ;
        RECT 9.4410 13.1765 9.4590 14.3365 ;
        RECT 5.8770 13.1765 5.8950 14.3365 ;
        RECT 5.1120 13.2130 5.1480 14.3270 ;
        RECT 4.9590 13.2130 4.9860 14.3270 ;
        RECT 3.7170 13.1765 3.7350 14.3365 ;
        RECT 0.1530 13.1765 0.1710 14.3365 ;
        RECT 9.4410 14.2565 9.4590 15.4165 ;
        RECT 5.8770 14.2565 5.8950 15.4165 ;
        RECT 5.1120 14.2930 5.1480 15.4070 ;
        RECT 4.9590 14.2930 4.9860 15.4070 ;
        RECT 3.7170 14.2565 3.7350 15.4165 ;
        RECT 0.1530 14.2565 0.1710 15.4165 ;
        RECT 9.4410 15.3365 9.4590 16.4965 ;
        RECT 5.8770 15.3365 5.8950 16.4965 ;
        RECT 5.1120 15.3730 5.1480 16.4870 ;
        RECT 4.9590 15.3730 4.9860 16.4870 ;
        RECT 3.7170 15.3365 3.7350 16.4965 ;
        RECT 0.1530 15.3365 0.1710 16.4965 ;
        RECT 9.4410 16.4165 9.4590 17.5765 ;
        RECT 5.8770 16.4165 5.8950 17.5765 ;
        RECT 5.1120 16.4530 5.1480 17.5670 ;
        RECT 4.9590 16.4530 4.9860 17.5670 ;
        RECT 3.7170 16.4165 3.7350 17.5765 ;
        RECT 0.1530 16.4165 0.1710 17.5765 ;
        RECT 9.4410 17.4965 9.4590 18.6565 ;
        RECT 5.8770 17.4965 5.8950 18.6565 ;
        RECT 5.1120 17.5330 5.1480 18.6470 ;
        RECT 4.9590 17.5330 4.9860 18.6470 ;
        RECT 3.7170 17.4965 3.7350 18.6565 ;
        RECT 0.1530 17.4965 0.1710 18.6565 ;
        RECT 9.4410 18.5765 9.4590 19.7365 ;
        RECT 5.8770 18.5765 5.8950 19.7365 ;
        RECT 5.1120 18.6130 5.1480 19.7270 ;
        RECT 4.9590 18.6130 4.9860 19.7270 ;
        RECT 3.7170 18.5765 3.7350 19.7365 ;
        RECT 0.1530 18.5765 0.1710 19.7365 ;
        RECT 9.4410 19.6565 9.4590 20.8165 ;
        RECT 5.8770 19.6565 5.8950 20.8165 ;
        RECT 5.1120 19.6930 5.1480 20.8070 ;
        RECT 4.9590 19.6930 4.9860 20.8070 ;
        RECT 3.7170 19.6565 3.7350 20.8165 ;
        RECT 0.1530 19.6565 0.1710 20.8165 ;
        RECT 9.4410 20.7365 9.4590 21.8965 ;
        RECT 5.8770 20.7365 5.8950 21.8965 ;
        RECT 5.1120 20.7730 5.1480 21.8870 ;
        RECT 4.9590 20.7730 4.9860 21.8870 ;
        RECT 3.7170 20.7365 3.7350 21.8965 ;
        RECT 0.1530 20.7365 0.1710 21.8965 ;
        RECT 9.4410 21.8165 9.4590 22.9765 ;
        RECT 5.8770 21.8165 5.8950 22.9765 ;
        RECT 5.1120 21.8530 5.1480 22.9670 ;
        RECT 4.9590 21.8530 4.9860 22.9670 ;
        RECT 3.7170 21.8165 3.7350 22.9765 ;
        RECT 0.1530 21.8165 0.1710 22.9765 ;
        RECT 9.4410 22.8965 9.4590 24.0565 ;
        RECT 5.8770 22.8965 5.8950 24.0565 ;
        RECT 5.1120 22.9330 5.1480 24.0470 ;
        RECT 4.9590 22.9330 4.9860 24.0470 ;
        RECT 3.7170 22.8965 3.7350 24.0565 ;
        RECT 0.1530 22.8965 0.1710 24.0565 ;
        RECT 9.4410 23.9765 9.4590 25.1365 ;
        RECT 5.8770 23.9765 5.8950 25.1365 ;
        RECT 5.1120 24.0130 5.1480 25.1270 ;
        RECT 4.9590 24.0130 4.9860 25.1270 ;
        RECT 3.7170 23.9765 3.7350 25.1365 ;
        RECT 0.1530 23.9765 0.1710 25.1365 ;
        RECT 9.4410 25.0565 9.4590 26.2165 ;
        RECT 5.8770 25.0565 5.8950 26.2165 ;
        RECT 5.1120 25.0930 5.1480 26.2070 ;
        RECT 4.9590 25.0930 4.9860 26.2070 ;
        RECT 3.7170 25.0565 3.7350 26.2165 ;
        RECT 0.1530 25.0565 0.1710 26.2165 ;
        RECT 9.4410 26.1365 9.4590 27.2965 ;
        RECT 5.8770 26.1365 5.8950 27.2965 ;
        RECT 5.1120 26.1730 5.1480 27.2870 ;
        RECT 4.9590 26.1730 4.9860 27.2870 ;
        RECT 3.7170 26.1365 3.7350 27.2965 ;
        RECT 0.1530 26.1365 0.1710 27.2965 ;
        RECT 9.4410 27.2165 9.4590 28.3765 ;
        RECT 5.8770 27.2165 5.8950 28.3765 ;
        RECT 5.1120 27.2530 5.1480 28.3670 ;
        RECT 4.9590 27.2530 4.9860 28.3670 ;
        RECT 3.7170 27.2165 3.7350 28.3765 ;
        RECT 0.1530 27.2165 0.1710 28.3765 ;
        RECT 9.4410 28.2965 9.4590 29.4565 ;
        RECT 5.8770 28.2965 5.8950 29.4565 ;
        RECT 5.1120 28.3330 5.1480 29.4470 ;
        RECT 4.9590 28.3330 4.9860 29.4470 ;
        RECT 3.7170 28.2965 3.7350 29.4565 ;
        RECT 0.1530 28.2965 0.1710 29.4565 ;
        RECT 9.4410 29.3765 9.4590 30.5365 ;
        RECT 5.8770 29.3765 5.8950 30.5365 ;
        RECT 5.1120 29.4130 5.1480 30.5270 ;
        RECT 4.9590 29.4130 4.9860 30.5270 ;
        RECT 3.7170 29.3765 3.7350 30.5365 ;
        RECT 0.1530 29.3765 0.1710 30.5365 ;
        RECT 9.4410 30.4565 9.4590 31.6165 ;
        RECT 5.8770 30.4565 5.8950 31.6165 ;
        RECT 5.1120 30.4930 5.1480 31.6070 ;
        RECT 4.9590 30.4930 4.9860 31.6070 ;
        RECT 3.7170 30.4565 3.7350 31.6165 ;
        RECT 0.1530 30.4565 0.1710 31.6165 ;
        RECT 9.4410 31.5365 9.4590 32.6965 ;
        RECT 5.8770 31.5365 5.8950 32.6965 ;
        RECT 5.1120 31.5730 5.1480 32.6870 ;
        RECT 4.9590 31.5730 4.9860 32.6870 ;
        RECT 3.7170 31.5365 3.7350 32.6965 ;
        RECT 0.1530 31.5365 0.1710 32.6965 ;
        RECT 9.4410 32.6165 9.4590 33.7765 ;
        RECT 5.8770 32.6165 5.8950 33.7765 ;
        RECT 5.1120 32.6530 5.1480 33.7670 ;
        RECT 4.9590 32.6530 4.9860 33.7670 ;
        RECT 3.7170 32.6165 3.7350 33.7765 ;
        RECT 0.1530 32.6165 0.1710 33.7765 ;
        RECT 9.4410 33.6965 9.4590 34.8565 ;
        RECT 5.8770 33.6965 5.8950 34.8565 ;
        RECT 5.1120 33.7330 5.1480 34.8470 ;
        RECT 4.9590 33.7330 4.9860 34.8470 ;
        RECT 3.7170 33.6965 3.7350 34.8565 ;
        RECT 0.1530 33.6965 0.1710 34.8565 ;
        RECT 9.4410 34.7765 9.4590 35.9365 ;
        RECT 5.8770 34.7765 5.8950 35.9365 ;
        RECT 5.1120 34.8130 5.1480 35.9270 ;
        RECT 4.9590 34.8130 4.9860 35.9270 ;
        RECT 3.7170 34.7765 3.7350 35.9365 ;
        RECT 0.1530 34.7765 0.1710 35.9365 ;
        RECT 9.4410 35.8565 9.4590 37.0165 ;
        RECT 5.8770 35.8565 5.8950 37.0165 ;
        RECT 5.1120 35.8930 5.1480 37.0070 ;
        RECT 4.9590 35.8930 4.9860 37.0070 ;
        RECT 3.7170 35.8565 3.7350 37.0165 ;
        RECT 0.1530 35.8565 0.1710 37.0165 ;
        RECT 9.4410 36.9365 9.4590 38.0965 ;
        RECT 5.8770 36.9365 5.8950 38.0965 ;
        RECT 5.1120 36.9730 5.1480 38.0870 ;
        RECT 4.9590 36.9730 4.9860 38.0870 ;
        RECT 3.7170 36.9365 3.7350 38.0965 ;
        RECT 0.1530 36.9365 0.1710 38.0965 ;
        RECT 9.4410 38.0165 9.4590 39.1765 ;
        RECT 5.8770 38.0165 5.8950 39.1765 ;
        RECT 5.1120 38.0530 5.1480 39.1670 ;
        RECT 4.9590 38.0530 4.9860 39.1670 ;
        RECT 3.7170 38.0165 3.7350 39.1765 ;
        RECT 0.1530 38.0165 0.1710 39.1765 ;
        RECT 9.4410 39.0965 9.4590 40.2565 ;
        RECT 5.8770 39.0965 5.8950 40.2565 ;
        RECT 5.1120 39.1330 5.1480 40.2470 ;
        RECT 4.9590 39.1330 4.9860 40.2470 ;
        RECT 3.7170 39.0965 3.7350 40.2565 ;
        RECT 0.1530 39.0965 0.1710 40.2565 ;
        RECT 9.4410 40.1765 9.4590 41.3365 ;
        RECT 5.8770 40.1765 5.8950 41.3365 ;
        RECT 5.1120 40.2130 5.1480 41.3270 ;
        RECT 4.9590 40.2130 4.9860 41.3270 ;
        RECT 3.7170 40.1765 3.7350 41.3365 ;
        RECT 0.1530 40.1765 0.1710 41.3365 ;
        RECT 9.4410 41.2565 9.4590 42.4165 ;
        RECT 5.8770 41.2565 5.8950 42.4165 ;
        RECT 5.1120 41.2930 5.1480 42.4070 ;
        RECT 4.9590 41.2930 4.9860 42.4070 ;
        RECT 3.7170 41.2565 3.7350 42.4165 ;
        RECT 0.1530 41.2565 0.1710 42.4165 ;
        RECT 9.4410 42.3365 9.4590 43.4965 ;
        RECT 5.8770 42.3365 5.8950 43.4965 ;
        RECT 5.1120 42.3730 5.1480 43.4870 ;
        RECT 4.9590 42.3730 4.9860 43.4870 ;
        RECT 3.7170 42.3365 3.7350 43.4965 ;
        RECT 0.1530 42.3365 0.1710 43.4965 ;
        RECT 9.4410 43.4165 9.4590 51.6235 ;
        RECT 5.8770 43.4165 5.8950 51.6235 ;
        RECT 4.9230 43.6400 5.1570 51.3230 ;
        RECT 5.1120 43.4600 5.1480 51.5970 ;
        RECT 4.9590 43.4600 4.9860 51.5940 ;
        RECT 3.7170 43.4165 3.7350 51.6235 ;
        RECT 0.1530 43.4165 0.1710 51.6235 ;
        RECT 9.4410 51.5435 9.4590 52.7035 ;
        RECT 5.8770 51.5435 5.8950 52.7035 ;
        RECT 5.1120 51.5800 5.1480 52.6940 ;
        RECT 4.9590 51.5800 4.9860 52.6940 ;
        RECT 3.7170 51.5435 3.7350 52.7035 ;
        RECT 0.1530 51.5435 0.1710 52.7035 ;
        RECT 9.4410 52.6235 9.4590 53.7835 ;
        RECT 5.8770 52.6235 5.8950 53.7835 ;
        RECT 5.1120 52.6600 5.1480 53.7740 ;
        RECT 4.9590 52.6600 4.9860 53.7740 ;
        RECT 3.7170 52.6235 3.7350 53.7835 ;
        RECT 0.1530 52.6235 0.1710 53.7835 ;
        RECT 9.4410 53.7035 9.4590 54.8635 ;
        RECT 5.8770 53.7035 5.8950 54.8635 ;
        RECT 5.1120 53.7400 5.1480 54.8540 ;
        RECT 4.9590 53.7400 4.9860 54.8540 ;
        RECT 3.7170 53.7035 3.7350 54.8635 ;
        RECT 0.1530 53.7035 0.1710 54.8635 ;
        RECT 9.4410 54.7835 9.4590 55.9435 ;
        RECT 5.8770 54.7835 5.8950 55.9435 ;
        RECT 5.1120 54.8200 5.1480 55.9340 ;
        RECT 4.9590 54.8200 4.9860 55.9340 ;
        RECT 3.7170 54.7835 3.7350 55.9435 ;
        RECT 0.1530 54.7835 0.1710 55.9435 ;
        RECT 9.4410 55.8635 9.4590 57.0235 ;
        RECT 5.8770 55.8635 5.8950 57.0235 ;
        RECT 5.1120 55.9000 5.1480 57.0140 ;
        RECT 4.9590 55.9000 4.9860 57.0140 ;
        RECT 3.7170 55.8635 3.7350 57.0235 ;
        RECT 0.1530 55.8635 0.1710 57.0235 ;
        RECT 9.4410 56.9435 9.4590 58.1035 ;
        RECT 5.8770 56.9435 5.8950 58.1035 ;
        RECT 5.1120 56.9800 5.1480 58.0940 ;
        RECT 4.9590 56.9800 4.9860 58.0940 ;
        RECT 3.7170 56.9435 3.7350 58.1035 ;
        RECT 0.1530 56.9435 0.1710 58.1035 ;
        RECT 9.4410 58.0235 9.4590 59.1835 ;
        RECT 5.8770 58.0235 5.8950 59.1835 ;
        RECT 5.1120 58.0600 5.1480 59.1740 ;
        RECT 4.9590 58.0600 4.9860 59.1740 ;
        RECT 3.7170 58.0235 3.7350 59.1835 ;
        RECT 0.1530 58.0235 0.1710 59.1835 ;
        RECT 9.4410 59.1035 9.4590 60.2635 ;
        RECT 5.8770 59.1035 5.8950 60.2635 ;
        RECT 5.1120 59.1400 5.1480 60.2540 ;
        RECT 4.9590 59.1400 4.9860 60.2540 ;
        RECT 3.7170 59.1035 3.7350 60.2635 ;
        RECT 0.1530 59.1035 0.1710 60.2635 ;
        RECT 9.4410 60.1835 9.4590 61.3435 ;
        RECT 5.8770 60.1835 5.8950 61.3435 ;
        RECT 5.1120 60.2200 5.1480 61.3340 ;
        RECT 4.9590 60.2200 4.9860 61.3340 ;
        RECT 3.7170 60.1835 3.7350 61.3435 ;
        RECT 0.1530 60.1835 0.1710 61.3435 ;
        RECT 9.4410 61.2635 9.4590 62.4235 ;
        RECT 5.8770 61.2635 5.8950 62.4235 ;
        RECT 5.1120 61.3000 5.1480 62.4140 ;
        RECT 4.9590 61.3000 4.9860 62.4140 ;
        RECT 3.7170 61.2635 3.7350 62.4235 ;
        RECT 0.1530 61.2635 0.1710 62.4235 ;
        RECT 9.4410 62.3435 9.4590 63.5035 ;
        RECT 5.8770 62.3435 5.8950 63.5035 ;
        RECT 5.1120 62.3800 5.1480 63.4940 ;
        RECT 4.9590 62.3800 4.9860 63.4940 ;
        RECT 3.7170 62.3435 3.7350 63.5035 ;
        RECT 0.1530 62.3435 0.1710 63.5035 ;
        RECT 9.4410 63.4235 9.4590 64.5835 ;
        RECT 5.8770 63.4235 5.8950 64.5835 ;
        RECT 5.1120 63.4600 5.1480 64.5740 ;
        RECT 4.9590 63.4600 4.9860 64.5740 ;
        RECT 3.7170 63.4235 3.7350 64.5835 ;
        RECT 0.1530 63.4235 0.1710 64.5835 ;
        RECT 9.4410 64.5035 9.4590 65.6635 ;
        RECT 5.8770 64.5035 5.8950 65.6635 ;
        RECT 5.1120 64.5400 5.1480 65.6540 ;
        RECT 4.9590 64.5400 4.9860 65.6540 ;
        RECT 3.7170 64.5035 3.7350 65.6635 ;
        RECT 0.1530 64.5035 0.1710 65.6635 ;
        RECT 9.4410 65.5835 9.4590 66.7435 ;
        RECT 5.8770 65.5835 5.8950 66.7435 ;
        RECT 5.1120 65.6200 5.1480 66.7340 ;
        RECT 4.9590 65.6200 4.9860 66.7340 ;
        RECT 3.7170 65.5835 3.7350 66.7435 ;
        RECT 0.1530 65.5835 0.1710 66.7435 ;
        RECT 9.4410 66.6635 9.4590 67.8235 ;
        RECT 5.8770 66.6635 5.8950 67.8235 ;
        RECT 5.1120 66.7000 5.1480 67.8140 ;
        RECT 4.9590 66.7000 4.9860 67.8140 ;
        RECT 3.7170 66.6635 3.7350 67.8235 ;
        RECT 0.1530 66.6635 0.1710 67.8235 ;
        RECT 9.4410 67.7435 9.4590 68.9035 ;
        RECT 5.8770 67.7435 5.8950 68.9035 ;
        RECT 5.1120 67.7800 5.1480 68.8940 ;
        RECT 4.9590 67.7800 4.9860 68.8940 ;
        RECT 3.7170 67.7435 3.7350 68.9035 ;
        RECT 0.1530 67.7435 0.1710 68.9035 ;
        RECT 9.4410 68.8235 9.4590 69.9835 ;
        RECT 5.8770 68.8235 5.8950 69.9835 ;
        RECT 5.1120 68.8600 5.1480 69.9740 ;
        RECT 4.9590 68.8600 4.9860 69.9740 ;
        RECT 3.7170 68.8235 3.7350 69.9835 ;
        RECT 0.1530 68.8235 0.1710 69.9835 ;
        RECT 9.4410 69.9035 9.4590 71.0635 ;
        RECT 5.8770 69.9035 5.8950 71.0635 ;
        RECT 5.1120 69.9400 5.1480 71.0540 ;
        RECT 4.9590 69.9400 4.9860 71.0540 ;
        RECT 3.7170 69.9035 3.7350 71.0635 ;
        RECT 0.1530 69.9035 0.1710 71.0635 ;
        RECT 9.4410 70.9835 9.4590 72.1435 ;
        RECT 5.8770 70.9835 5.8950 72.1435 ;
        RECT 5.1120 71.0200 5.1480 72.1340 ;
        RECT 4.9590 71.0200 4.9860 72.1340 ;
        RECT 3.7170 70.9835 3.7350 72.1435 ;
        RECT 0.1530 70.9835 0.1710 72.1435 ;
        RECT 9.4410 72.0635 9.4590 73.2235 ;
        RECT 5.8770 72.0635 5.8950 73.2235 ;
        RECT 5.1120 72.1000 5.1480 73.2140 ;
        RECT 4.9590 72.1000 4.9860 73.2140 ;
        RECT 3.7170 72.0635 3.7350 73.2235 ;
        RECT 0.1530 72.0635 0.1710 73.2235 ;
        RECT 9.4410 73.1435 9.4590 74.3035 ;
        RECT 5.8770 73.1435 5.8950 74.3035 ;
        RECT 5.1120 73.1800 5.1480 74.2940 ;
        RECT 4.9590 73.1800 4.9860 74.2940 ;
        RECT 3.7170 73.1435 3.7350 74.3035 ;
        RECT 0.1530 73.1435 0.1710 74.3035 ;
        RECT 9.4410 74.2235 9.4590 75.3835 ;
        RECT 5.8770 74.2235 5.8950 75.3835 ;
        RECT 5.1120 74.2600 5.1480 75.3740 ;
        RECT 4.9590 74.2600 4.9860 75.3740 ;
        RECT 3.7170 74.2235 3.7350 75.3835 ;
        RECT 0.1530 74.2235 0.1710 75.3835 ;
        RECT 9.4410 75.3035 9.4590 76.4635 ;
        RECT 5.8770 75.3035 5.8950 76.4635 ;
        RECT 5.1120 75.3400 5.1480 76.4540 ;
        RECT 4.9590 75.3400 4.9860 76.4540 ;
        RECT 3.7170 75.3035 3.7350 76.4635 ;
        RECT 0.1530 75.3035 0.1710 76.4635 ;
        RECT 9.4410 76.3835 9.4590 77.5435 ;
        RECT 5.8770 76.3835 5.8950 77.5435 ;
        RECT 5.1120 76.4200 5.1480 77.5340 ;
        RECT 4.9590 76.4200 4.9860 77.5340 ;
        RECT 3.7170 76.3835 3.7350 77.5435 ;
        RECT 0.1530 76.3835 0.1710 77.5435 ;
        RECT 9.4410 77.4635 9.4590 78.6235 ;
        RECT 5.8770 77.4635 5.8950 78.6235 ;
        RECT 5.1120 77.5000 5.1480 78.6140 ;
        RECT 4.9590 77.5000 4.9860 78.6140 ;
        RECT 3.7170 77.4635 3.7350 78.6235 ;
        RECT 0.1530 77.4635 0.1710 78.6235 ;
        RECT 9.4410 78.5435 9.4590 79.7035 ;
        RECT 5.8770 78.5435 5.8950 79.7035 ;
        RECT 5.1120 78.5800 5.1480 79.6940 ;
        RECT 4.9590 78.5800 4.9860 79.6940 ;
        RECT 3.7170 78.5435 3.7350 79.7035 ;
        RECT 0.1530 78.5435 0.1710 79.7035 ;
        RECT 9.4410 79.6235 9.4590 80.7835 ;
        RECT 5.8770 79.6235 5.8950 80.7835 ;
        RECT 5.1120 79.6600 5.1480 80.7740 ;
        RECT 4.9590 79.6600 4.9860 80.7740 ;
        RECT 3.7170 79.6235 3.7350 80.7835 ;
        RECT 0.1530 79.6235 0.1710 80.7835 ;
        RECT 9.4410 80.7035 9.4590 81.8635 ;
        RECT 5.8770 80.7035 5.8950 81.8635 ;
        RECT 5.1120 80.7400 5.1480 81.8540 ;
        RECT 4.9590 80.7400 4.9860 81.8540 ;
        RECT 3.7170 80.7035 3.7350 81.8635 ;
        RECT 0.1530 80.7035 0.1710 81.8635 ;
        RECT 9.4410 81.7835 9.4590 82.9435 ;
        RECT 5.8770 81.7835 5.8950 82.9435 ;
        RECT 5.1120 81.8200 5.1480 82.9340 ;
        RECT 4.9590 81.8200 4.9860 82.9340 ;
        RECT 3.7170 81.7835 3.7350 82.9435 ;
        RECT 0.1530 81.7835 0.1710 82.9435 ;
        RECT 9.4410 82.8635 9.4590 84.0235 ;
        RECT 5.8770 82.8635 5.8950 84.0235 ;
        RECT 5.1120 82.9000 5.1480 84.0140 ;
        RECT 4.9590 82.9000 4.9860 84.0140 ;
        RECT 3.7170 82.8635 3.7350 84.0235 ;
        RECT 0.1530 82.8635 0.1710 84.0235 ;
        RECT 9.4410 83.9435 9.4590 85.1035 ;
        RECT 5.8770 83.9435 5.8950 85.1035 ;
        RECT 5.1120 83.9800 5.1480 85.0940 ;
        RECT 4.9590 83.9800 4.9860 85.0940 ;
        RECT 3.7170 83.9435 3.7350 85.1035 ;
        RECT 0.1530 83.9435 0.1710 85.1035 ;
        RECT 9.4410 85.0235 9.4590 86.1835 ;
        RECT 5.8770 85.0235 5.8950 86.1835 ;
        RECT 5.1120 85.0600 5.1480 86.1740 ;
        RECT 4.9590 85.0600 4.9860 86.1740 ;
        RECT 3.7170 85.0235 3.7350 86.1835 ;
        RECT 0.1530 85.0235 0.1710 86.1835 ;
        RECT 9.4410 86.1035 9.4590 87.2635 ;
        RECT 5.8770 86.1035 5.8950 87.2635 ;
        RECT 5.1120 86.1400 5.1480 87.2540 ;
        RECT 4.9590 86.1400 4.9860 87.2540 ;
        RECT 3.7170 86.1035 3.7350 87.2635 ;
        RECT 0.1530 86.1035 0.1710 87.2635 ;
        RECT 9.4410 87.1835 9.4590 88.3435 ;
        RECT 5.8770 87.1835 5.8950 88.3435 ;
        RECT 5.1120 87.2200 5.1480 88.3340 ;
        RECT 4.9590 87.2200 4.9860 88.3340 ;
        RECT 3.7170 87.1835 3.7350 88.3435 ;
        RECT 0.1530 87.1835 0.1710 88.3435 ;
        RECT 9.4410 88.2635 9.4590 89.4235 ;
        RECT 5.8770 88.2635 5.8950 89.4235 ;
        RECT 5.1120 88.3000 5.1480 89.4140 ;
        RECT 4.9590 88.3000 4.9860 89.4140 ;
        RECT 3.7170 88.2635 3.7350 89.4235 ;
        RECT 0.1530 88.2635 0.1710 89.4235 ;
        RECT 9.4410 89.3435 9.4590 90.5035 ;
        RECT 5.8770 89.3435 5.8950 90.5035 ;
        RECT 5.1120 89.3800 5.1480 90.4940 ;
        RECT 4.9590 89.3800 4.9860 90.4940 ;
        RECT 3.7170 89.3435 3.7350 90.5035 ;
        RECT 0.1530 89.3435 0.1710 90.5035 ;
        RECT 9.4410 90.4235 9.4590 91.5835 ;
        RECT 5.8770 90.4235 5.8950 91.5835 ;
        RECT 5.1120 90.4600 5.1480 91.5740 ;
        RECT 4.9590 90.4600 4.9860 91.5740 ;
        RECT 3.7170 90.4235 3.7350 91.5835 ;
        RECT 0.1530 90.4235 0.1710 91.5835 ;
        RECT 9.4410 91.5035 9.4590 92.6635 ;
        RECT 5.8770 91.5035 5.8950 92.6635 ;
        RECT 5.1120 91.5400 5.1480 92.6540 ;
        RECT 4.9590 91.5400 4.9860 92.6540 ;
        RECT 3.7170 91.5035 3.7350 92.6635 ;
        RECT 0.1530 91.5035 0.1710 92.6635 ;
        RECT 9.4410 92.5835 9.4590 93.7435 ;
        RECT 5.8770 92.5835 5.8950 93.7435 ;
        RECT 5.1120 92.6200 5.1480 93.7340 ;
        RECT 4.9590 92.6200 4.9860 93.7340 ;
        RECT 3.7170 92.5835 3.7350 93.7435 ;
        RECT 0.1530 92.5835 0.1710 93.7435 ;
        RECT 9.4410 93.6635 9.4590 94.8235 ;
        RECT 5.8770 93.6635 5.8950 94.8235 ;
        RECT 5.1120 93.7000 5.1480 94.8140 ;
        RECT 4.9590 93.7000 4.9860 94.8140 ;
        RECT 3.7170 93.6635 3.7350 94.8235 ;
        RECT 0.1530 93.6635 0.1710 94.8235 ;
      LAYER V3  ;
        RECT 0.1530 1.0760 0.1710 1.1240 ;
        RECT 3.7170 1.0760 3.7350 1.1240 ;
        RECT 4.9590 1.0760 4.9860 1.1240 ;
        RECT 5.1120 1.0760 5.1480 1.1240 ;
        RECT 5.8770 1.0760 5.8950 1.1240 ;
        RECT 9.4410 1.0760 9.4590 1.1240 ;
        RECT 0.1530 2.1560 0.1710 2.2040 ;
        RECT 3.7170 2.1560 3.7350 2.2040 ;
        RECT 4.9590 2.1560 4.9860 2.2040 ;
        RECT 5.1120 2.1560 5.1480 2.2040 ;
        RECT 5.8770 2.1560 5.8950 2.2040 ;
        RECT 9.4410 2.1560 9.4590 2.2040 ;
        RECT 0.1530 3.2360 0.1710 3.2840 ;
        RECT 3.7170 3.2360 3.7350 3.2840 ;
        RECT 4.9590 3.2360 4.9860 3.2840 ;
        RECT 5.1120 3.2360 5.1480 3.2840 ;
        RECT 5.8770 3.2360 5.8950 3.2840 ;
        RECT 9.4410 3.2360 9.4590 3.2840 ;
        RECT 0.1530 4.3160 0.1710 4.3640 ;
        RECT 3.7170 4.3160 3.7350 4.3640 ;
        RECT 4.9590 4.3160 4.9860 4.3640 ;
        RECT 5.1120 4.3160 5.1480 4.3640 ;
        RECT 5.8770 4.3160 5.8950 4.3640 ;
        RECT 9.4410 4.3160 9.4590 4.3640 ;
        RECT 0.1530 5.3960 0.1710 5.4440 ;
        RECT 3.7170 5.3960 3.7350 5.4440 ;
        RECT 4.9590 5.3960 4.9860 5.4440 ;
        RECT 5.1120 5.3960 5.1480 5.4440 ;
        RECT 5.8770 5.3960 5.8950 5.4440 ;
        RECT 9.4410 5.3960 9.4590 5.4440 ;
        RECT 0.1530 6.4760 0.1710 6.5240 ;
        RECT 3.7170 6.4760 3.7350 6.5240 ;
        RECT 4.9590 6.4760 4.9860 6.5240 ;
        RECT 5.1120 6.4760 5.1480 6.5240 ;
        RECT 5.8770 6.4760 5.8950 6.5240 ;
        RECT 9.4410 6.4760 9.4590 6.5240 ;
        RECT 0.1530 7.5560 0.1710 7.6040 ;
        RECT 3.7170 7.5560 3.7350 7.6040 ;
        RECT 4.9590 7.5560 4.9860 7.6040 ;
        RECT 5.1120 7.5560 5.1480 7.6040 ;
        RECT 5.8770 7.5560 5.8950 7.6040 ;
        RECT 9.4410 7.5560 9.4590 7.6040 ;
        RECT 0.1530 8.6360 0.1710 8.6840 ;
        RECT 3.7170 8.6360 3.7350 8.6840 ;
        RECT 4.9590 8.6360 4.9860 8.6840 ;
        RECT 5.1120 8.6360 5.1480 8.6840 ;
        RECT 5.8770 8.6360 5.8950 8.6840 ;
        RECT 9.4410 8.6360 9.4590 8.6840 ;
        RECT 0.1530 9.7160 0.1710 9.7640 ;
        RECT 3.7170 9.7160 3.7350 9.7640 ;
        RECT 4.9590 9.7160 4.9860 9.7640 ;
        RECT 5.1120 9.7160 5.1480 9.7640 ;
        RECT 5.8770 9.7160 5.8950 9.7640 ;
        RECT 9.4410 9.7160 9.4590 9.7640 ;
        RECT 0.1530 10.7960 0.1710 10.8440 ;
        RECT 3.7170 10.7960 3.7350 10.8440 ;
        RECT 4.9590 10.7960 4.9860 10.8440 ;
        RECT 5.1120 10.7960 5.1480 10.8440 ;
        RECT 5.8770 10.7960 5.8950 10.8440 ;
        RECT 9.4410 10.7960 9.4590 10.8440 ;
        RECT 0.1530 11.8760 0.1710 11.9240 ;
        RECT 3.7170 11.8760 3.7350 11.9240 ;
        RECT 4.9590 11.8760 4.9860 11.9240 ;
        RECT 5.1120 11.8760 5.1480 11.9240 ;
        RECT 5.8770 11.8760 5.8950 11.9240 ;
        RECT 9.4410 11.8760 9.4590 11.9240 ;
        RECT 0.1530 12.9560 0.1710 13.0040 ;
        RECT 3.7170 12.9560 3.7350 13.0040 ;
        RECT 4.9590 12.9560 4.9860 13.0040 ;
        RECT 5.1120 12.9560 5.1480 13.0040 ;
        RECT 5.8770 12.9560 5.8950 13.0040 ;
        RECT 9.4410 12.9560 9.4590 13.0040 ;
        RECT 0.1530 14.0360 0.1710 14.0840 ;
        RECT 3.7170 14.0360 3.7350 14.0840 ;
        RECT 4.9590 14.0360 4.9860 14.0840 ;
        RECT 5.1120 14.0360 5.1480 14.0840 ;
        RECT 5.8770 14.0360 5.8950 14.0840 ;
        RECT 9.4410 14.0360 9.4590 14.0840 ;
        RECT 0.1530 15.1160 0.1710 15.1640 ;
        RECT 3.7170 15.1160 3.7350 15.1640 ;
        RECT 4.9590 15.1160 4.9860 15.1640 ;
        RECT 5.1120 15.1160 5.1480 15.1640 ;
        RECT 5.8770 15.1160 5.8950 15.1640 ;
        RECT 9.4410 15.1160 9.4590 15.1640 ;
        RECT 0.1530 16.1960 0.1710 16.2440 ;
        RECT 3.7170 16.1960 3.7350 16.2440 ;
        RECT 4.9590 16.1960 4.9860 16.2440 ;
        RECT 5.1120 16.1960 5.1480 16.2440 ;
        RECT 5.8770 16.1960 5.8950 16.2440 ;
        RECT 9.4410 16.1960 9.4590 16.2440 ;
        RECT 0.1530 17.2760 0.1710 17.3240 ;
        RECT 3.7170 17.2760 3.7350 17.3240 ;
        RECT 4.9590 17.2760 4.9860 17.3240 ;
        RECT 5.1120 17.2760 5.1480 17.3240 ;
        RECT 5.8770 17.2760 5.8950 17.3240 ;
        RECT 9.4410 17.2760 9.4590 17.3240 ;
        RECT 0.1530 18.3560 0.1710 18.4040 ;
        RECT 3.7170 18.3560 3.7350 18.4040 ;
        RECT 4.9590 18.3560 4.9860 18.4040 ;
        RECT 5.1120 18.3560 5.1480 18.4040 ;
        RECT 5.8770 18.3560 5.8950 18.4040 ;
        RECT 9.4410 18.3560 9.4590 18.4040 ;
        RECT 0.1530 19.4360 0.1710 19.4840 ;
        RECT 3.7170 19.4360 3.7350 19.4840 ;
        RECT 4.9590 19.4360 4.9860 19.4840 ;
        RECT 5.1120 19.4360 5.1480 19.4840 ;
        RECT 5.8770 19.4360 5.8950 19.4840 ;
        RECT 9.4410 19.4360 9.4590 19.4840 ;
        RECT 0.1530 20.5160 0.1710 20.5640 ;
        RECT 3.7170 20.5160 3.7350 20.5640 ;
        RECT 4.9590 20.5160 4.9860 20.5640 ;
        RECT 5.1120 20.5160 5.1480 20.5640 ;
        RECT 5.8770 20.5160 5.8950 20.5640 ;
        RECT 9.4410 20.5160 9.4590 20.5640 ;
        RECT 0.1530 21.5960 0.1710 21.6440 ;
        RECT 3.7170 21.5960 3.7350 21.6440 ;
        RECT 4.9590 21.5960 4.9860 21.6440 ;
        RECT 5.1120 21.5960 5.1480 21.6440 ;
        RECT 5.8770 21.5960 5.8950 21.6440 ;
        RECT 9.4410 21.5960 9.4590 21.6440 ;
        RECT 0.1530 22.6760 0.1710 22.7240 ;
        RECT 3.7170 22.6760 3.7350 22.7240 ;
        RECT 4.9590 22.6760 4.9860 22.7240 ;
        RECT 5.1120 22.6760 5.1480 22.7240 ;
        RECT 5.8770 22.6760 5.8950 22.7240 ;
        RECT 9.4410 22.6760 9.4590 22.7240 ;
        RECT 0.1530 23.7560 0.1710 23.8040 ;
        RECT 3.7170 23.7560 3.7350 23.8040 ;
        RECT 4.9590 23.7560 4.9860 23.8040 ;
        RECT 5.1120 23.7560 5.1480 23.8040 ;
        RECT 5.8770 23.7560 5.8950 23.8040 ;
        RECT 9.4410 23.7560 9.4590 23.8040 ;
        RECT 0.1530 24.8360 0.1710 24.8840 ;
        RECT 3.7170 24.8360 3.7350 24.8840 ;
        RECT 4.9590 24.8360 4.9860 24.8840 ;
        RECT 5.1120 24.8360 5.1480 24.8840 ;
        RECT 5.8770 24.8360 5.8950 24.8840 ;
        RECT 9.4410 24.8360 9.4590 24.8840 ;
        RECT 0.1530 25.9160 0.1710 25.9640 ;
        RECT 3.7170 25.9160 3.7350 25.9640 ;
        RECT 4.9590 25.9160 4.9860 25.9640 ;
        RECT 5.1120 25.9160 5.1480 25.9640 ;
        RECT 5.8770 25.9160 5.8950 25.9640 ;
        RECT 9.4410 25.9160 9.4590 25.9640 ;
        RECT 0.1530 26.9960 0.1710 27.0440 ;
        RECT 3.7170 26.9960 3.7350 27.0440 ;
        RECT 4.9590 26.9960 4.9860 27.0440 ;
        RECT 5.1120 26.9960 5.1480 27.0440 ;
        RECT 5.8770 26.9960 5.8950 27.0440 ;
        RECT 9.4410 26.9960 9.4590 27.0440 ;
        RECT 0.1530 28.0760 0.1710 28.1240 ;
        RECT 3.7170 28.0760 3.7350 28.1240 ;
        RECT 4.9590 28.0760 4.9860 28.1240 ;
        RECT 5.1120 28.0760 5.1480 28.1240 ;
        RECT 5.8770 28.0760 5.8950 28.1240 ;
        RECT 9.4410 28.0760 9.4590 28.1240 ;
        RECT 0.1530 29.1560 0.1710 29.2040 ;
        RECT 3.7170 29.1560 3.7350 29.2040 ;
        RECT 4.9590 29.1560 4.9860 29.2040 ;
        RECT 5.1120 29.1560 5.1480 29.2040 ;
        RECT 5.8770 29.1560 5.8950 29.2040 ;
        RECT 9.4410 29.1560 9.4590 29.2040 ;
        RECT 0.1530 30.2360 0.1710 30.2840 ;
        RECT 3.7170 30.2360 3.7350 30.2840 ;
        RECT 4.9590 30.2360 4.9860 30.2840 ;
        RECT 5.1120 30.2360 5.1480 30.2840 ;
        RECT 5.8770 30.2360 5.8950 30.2840 ;
        RECT 9.4410 30.2360 9.4590 30.2840 ;
        RECT 0.1530 31.3160 0.1710 31.3640 ;
        RECT 3.7170 31.3160 3.7350 31.3640 ;
        RECT 4.9590 31.3160 4.9860 31.3640 ;
        RECT 5.1120 31.3160 5.1480 31.3640 ;
        RECT 5.8770 31.3160 5.8950 31.3640 ;
        RECT 9.4410 31.3160 9.4590 31.3640 ;
        RECT 0.1530 32.3960 0.1710 32.4440 ;
        RECT 3.7170 32.3960 3.7350 32.4440 ;
        RECT 4.9590 32.3960 4.9860 32.4440 ;
        RECT 5.1120 32.3960 5.1480 32.4440 ;
        RECT 5.8770 32.3960 5.8950 32.4440 ;
        RECT 9.4410 32.3960 9.4590 32.4440 ;
        RECT 0.1530 33.4760 0.1710 33.5240 ;
        RECT 3.7170 33.4760 3.7350 33.5240 ;
        RECT 4.9590 33.4760 4.9860 33.5240 ;
        RECT 5.1120 33.4760 5.1480 33.5240 ;
        RECT 5.8770 33.4760 5.8950 33.5240 ;
        RECT 9.4410 33.4760 9.4590 33.5240 ;
        RECT 0.1530 34.5560 0.1710 34.6040 ;
        RECT 3.7170 34.5560 3.7350 34.6040 ;
        RECT 4.9590 34.5560 4.9860 34.6040 ;
        RECT 5.1120 34.5560 5.1480 34.6040 ;
        RECT 5.8770 34.5560 5.8950 34.6040 ;
        RECT 9.4410 34.5560 9.4590 34.6040 ;
        RECT 0.1530 35.6360 0.1710 35.6840 ;
        RECT 3.7170 35.6360 3.7350 35.6840 ;
        RECT 4.9590 35.6360 4.9860 35.6840 ;
        RECT 5.1120 35.6360 5.1480 35.6840 ;
        RECT 5.8770 35.6360 5.8950 35.6840 ;
        RECT 9.4410 35.6360 9.4590 35.6840 ;
        RECT 0.1530 36.7160 0.1710 36.7640 ;
        RECT 3.7170 36.7160 3.7350 36.7640 ;
        RECT 4.9590 36.7160 4.9860 36.7640 ;
        RECT 5.1120 36.7160 5.1480 36.7640 ;
        RECT 5.8770 36.7160 5.8950 36.7640 ;
        RECT 9.4410 36.7160 9.4590 36.7640 ;
        RECT 0.1530 37.7960 0.1710 37.8440 ;
        RECT 3.7170 37.7960 3.7350 37.8440 ;
        RECT 4.9590 37.7960 4.9860 37.8440 ;
        RECT 5.1120 37.7960 5.1480 37.8440 ;
        RECT 5.8770 37.7960 5.8950 37.8440 ;
        RECT 9.4410 37.7960 9.4590 37.8440 ;
        RECT 0.1530 38.8760 0.1710 38.9240 ;
        RECT 3.7170 38.8760 3.7350 38.9240 ;
        RECT 4.9590 38.8760 4.9860 38.9240 ;
        RECT 5.1120 38.8760 5.1480 38.9240 ;
        RECT 5.8770 38.8760 5.8950 38.9240 ;
        RECT 9.4410 38.8760 9.4590 38.9240 ;
        RECT 0.1530 39.9560 0.1710 40.0040 ;
        RECT 3.7170 39.9560 3.7350 40.0040 ;
        RECT 4.9590 39.9560 4.9860 40.0040 ;
        RECT 5.1120 39.9560 5.1480 40.0040 ;
        RECT 5.8770 39.9560 5.8950 40.0040 ;
        RECT 9.4410 39.9560 9.4590 40.0040 ;
        RECT 0.1530 41.0360 0.1710 41.0840 ;
        RECT 3.7170 41.0360 3.7350 41.0840 ;
        RECT 4.9590 41.0360 4.9860 41.0840 ;
        RECT 5.1120 41.0360 5.1480 41.0840 ;
        RECT 5.8770 41.0360 5.8950 41.0840 ;
        RECT 9.4410 41.0360 9.4590 41.0840 ;
        RECT 0.1530 42.1160 0.1710 42.1640 ;
        RECT 3.7170 42.1160 3.7350 42.1640 ;
        RECT 4.9590 42.1160 4.9860 42.1640 ;
        RECT 5.1120 42.1160 5.1480 42.1640 ;
        RECT 5.8770 42.1160 5.8950 42.1640 ;
        RECT 9.4410 42.1160 9.4590 42.1640 ;
        RECT 0.1530 43.1960 0.1710 43.2440 ;
        RECT 3.7170 43.1960 3.7350 43.2440 ;
        RECT 4.9590 43.1960 4.9860 43.2440 ;
        RECT 5.1120 43.1960 5.1480 43.2440 ;
        RECT 5.8770 43.1960 5.8950 43.2440 ;
        RECT 9.4410 43.1960 9.4590 43.2440 ;
        RECT 0.1530 44.2110 0.1710 44.4270 ;
        RECT 4.9270 50.5470 4.9450 50.7630 ;
        RECT 4.9270 47.3790 4.9450 47.5950 ;
        RECT 4.9270 44.2110 4.9450 44.4270 ;
        RECT 4.9790 50.5470 4.9970 50.7630 ;
        RECT 4.9790 47.3790 4.9970 47.5950 ;
        RECT 4.9790 44.2110 4.9970 44.4270 ;
        RECT 5.0310 50.5470 5.0490 50.7630 ;
        RECT 5.0310 47.3790 5.0490 47.5950 ;
        RECT 5.0310 44.2110 5.0490 44.4270 ;
        RECT 5.0830 50.5470 5.1010 50.7630 ;
        RECT 5.0830 47.3790 5.1010 47.5950 ;
        RECT 5.0830 44.2110 5.1010 44.4270 ;
        RECT 5.1350 50.5470 5.1530 50.7630 ;
        RECT 5.1350 47.3790 5.1530 47.5950 ;
        RECT 5.1350 44.2110 5.1530 44.4270 ;
        RECT 0.1530 52.4030 0.1710 52.4510 ;
        RECT 3.7170 52.4030 3.7350 52.4510 ;
        RECT 4.9590 52.4030 4.9860 52.4510 ;
        RECT 5.1120 52.4030 5.1480 52.4510 ;
        RECT 5.8770 52.4030 5.8950 52.4510 ;
        RECT 9.4410 52.4030 9.4590 52.4510 ;
        RECT 0.1530 53.4830 0.1710 53.5310 ;
        RECT 3.7170 53.4830 3.7350 53.5310 ;
        RECT 4.9590 53.4830 4.9860 53.5310 ;
        RECT 5.1120 53.4830 5.1480 53.5310 ;
        RECT 5.8770 53.4830 5.8950 53.5310 ;
        RECT 9.4410 53.4830 9.4590 53.5310 ;
        RECT 0.1530 54.5630 0.1710 54.6110 ;
        RECT 3.7170 54.5630 3.7350 54.6110 ;
        RECT 4.9590 54.5630 4.9860 54.6110 ;
        RECT 5.1120 54.5630 5.1480 54.6110 ;
        RECT 5.8770 54.5630 5.8950 54.6110 ;
        RECT 9.4410 54.5630 9.4590 54.6110 ;
        RECT 0.1530 55.6430 0.1710 55.6910 ;
        RECT 3.7170 55.6430 3.7350 55.6910 ;
        RECT 4.9590 55.6430 4.9860 55.6910 ;
        RECT 5.1120 55.6430 5.1480 55.6910 ;
        RECT 5.8770 55.6430 5.8950 55.6910 ;
        RECT 9.4410 55.6430 9.4590 55.6910 ;
        RECT 0.1530 56.7230 0.1710 56.7710 ;
        RECT 3.7170 56.7230 3.7350 56.7710 ;
        RECT 4.9590 56.7230 4.9860 56.7710 ;
        RECT 5.1120 56.7230 5.1480 56.7710 ;
        RECT 5.8770 56.7230 5.8950 56.7710 ;
        RECT 9.4410 56.7230 9.4590 56.7710 ;
        RECT 0.1530 57.8030 0.1710 57.8510 ;
        RECT 3.7170 57.8030 3.7350 57.8510 ;
        RECT 4.9590 57.8030 4.9860 57.8510 ;
        RECT 5.1120 57.8030 5.1480 57.8510 ;
        RECT 5.8770 57.8030 5.8950 57.8510 ;
        RECT 9.4410 57.8030 9.4590 57.8510 ;
        RECT 0.1530 58.8830 0.1710 58.9310 ;
        RECT 3.7170 58.8830 3.7350 58.9310 ;
        RECT 4.9590 58.8830 4.9860 58.9310 ;
        RECT 5.1120 58.8830 5.1480 58.9310 ;
        RECT 5.8770 58.8830 5.8950 58.9310 ;
        RECT 9.4410 58.8830 9.4590 58.9310 ;
        RECT 0.1530 59.9630 0.1710 60.0110 ;
        RECT 3.7170 59.9630 3.7350 60.0110 ;
        RECT 4.9590 59.9630 4.9860 60.0110 ;
        RECT 5.1120 59.9630 5.1480 60.0110 ;
        RECT 5.8770 59.9630 5.8950 60.0110 ;
        RECT 9.4410 59.9630 9.4590 60.0110 ;
        RECT 0.1530 61.0430 0.1710 61.0910 ;
        RECT 3.7170 61.0430 3.7350 61.0910 ;
        RECT 4.9590 61.0430 4.9860 61.0910 ;
        RECT 5.1120 61.0430 5.1480 61.0910 ;
        RECT 5.8770 61.0430 5.8950 61.0910 ;
        RECT 9.4410 61.0430 9.4590 61.0910 ;
        RECT 0.1530 62.1230 0.1710 62.1710 ;
        RECT 3.7170 62.1230 3.7350 62.1710 ;
        RECT 4.9590 62.1230 4.9860 62.1710 ;
        RECT 5.1120 62.1230 5.1480 62.1710 ;
        RECT 5.8770 62.1230 5.8950 62.1710 ;
        RECT 9.4410 62.1230 9.4590 62.1710 ;
        RECT 0.1530 63.2030 0.1710 63.2510 ;
        RECT 3.7170 63.2030 3.7350 63.2510 ;
        RECT 4.9590 63.2030 4.9860 63.2510 ;
        RECT 5.1120 63.2030 5.1480 63.2510 ;
        RECT 5.8770 63.2030 5.8950 63.2510 ;
        RECT 9.4410 63.2030 9.4590 63.2510 ;
        RECT 0.1530 64.2830 0.1710 64.3310 ;
        RECT 3.7170 64.2830 3.7350 64.3310 ;
        RECT 4.9590 64.2830 4.9860 64.3310 ;
        RECT 5.1120 64.2830 5.1480 64.3310 ;
        RECT 5.8770 64.2830 5.8950 64.3310 ;
        RECT 9.4410 64.2830 9.4590 64.3310 ;
        RECT 0.1530 65.3630 0.1710 65.4110 ;
        RECT 3.7170 65.3630 3.7350 65.4110 ;
        RECT 4.9590 65.3630 4.9860 65.4110 ;
        RECT 5.1120 65.3630 5.1480 65.4110 ;
        RECT 5.8770 65.3630 5.8950 65.4110 ;
        RECT 9.4410 65.3630 9.4590 65.4110 ;
        RECT 0.1530 66.4430 0.1710 66.4910 ;
        RECT 3.7170 66.4430 3.7350 66.4910 ;
        RECT 4.9590 66.4430 4.9860 66.4910 ;
        RECT 5.1120 66.4430 5.1480 66.4910 ;
        RECT 5.8770 66.4430 5.8950 66.4910 ;
        RECT 9.4410 66.4430 9.4590 66.4910 ;
        RECT 0.1530 67.5230 0.1710 67.5710 ;
        RECT 3.7170 67.5230 3.7350 67.5710 ;
        RECT 4.9590 67.5230 4.9860 67.5710 ;
        RECT 5.1120 67.5230 5.1480 67.5710 ;
        RECT 5.8770 67.5230 5.8950 67.5710 ;
        RECT 9.4410 67.5230 9.4590 67.5710 ;
        RECT 0.1530 68.6030 0.1710 68.6510 ;
        RECT 3.7170 68.6030 3.7350 68.6510 ;
        RECT 4.9590 68.6030 4.9860 68.6510 ;
        RECT 5.1120 68.6030 5.1480 68.6510 ;
        RECT 5.8770 68.6030 5.8950 68.6510 ;
        RECT 9.4410 68.6030 9.4590 68.6510 ;
        RECT 0.1530 69.6830 0.1710 69.7310 ;
        RECT 3.7170 69.6830 3.7350 69.7310 ;
        RECT 4.9590 69.6830 4.9860 69.7310 ;
        RECT 5.1120 69.6830 5.1480 69.7310 ;
        RECT 5.8770 69.6830 5.8950 69.7310 ;
        RECT 9.4410 69.6830 9.4590 69.7310 ;
        RECT 0.1530 70.7630 0.1710 70.8110 ;
        RECT 3.7170 70.7630 3.7350 70.8110 ;
        RECT 4.9590 70.7630 4.9860 70.8110 ;
        RECT 5.1120 70.7630 5.1480 70.8110 ;
        RECT 5.8770 70.7630 5.8950 70.8110 ;
        RECT 9.4410 70.7630 9.4590 70.8110 ;
        RECT 0.1530 71.8430 0.1710 71.8910 ;
        RECT 3.7170 71.8430 3.7350 71.8910 ;
        RECT 4.9590 71.8430 4.9860 71.8910 ;
        RECT 5.1120 71.8430 5.1480 71.8910 ;
        RECT 5.8770 71.8430 5.8950 71.8910 ;
        RECT 9.4410 71.8430 9.4590 71.8910 ;
        RECT 0.1530 72.9230 0.1710 72.9710 ;
        RECT 3.7170 72.9230 3.7350 72.9710 ;
        RECT 4.9590 72.9230 4.9860 72.9710 ;
        RECT 5.1120 72.9230 5.1480 72.9710 ;
        RECT 5.8770 72.9230 5.8950 72.9710 ;
        RECT 9.4410 72.9230 9.4590 72.9710 ;
        RECT 0.1530 74.0030 0.1710 74.0510 ;
        RECT 3.7170 74.0030 3.7350 74.0510 ;
        RECT 4.9590 74.0030 4.9860 74.0510 ;
        RECT 5.1120 74.0030 5.1480 74.0510 ;
        RECT 5.8770 74.0030 5.8950 74.0510 ;
        RECT 9.4410 74.0030 9.4590 74.0510 ;
        RECT 0.1530 75.0830 0.1710 75.1310 ;
        RECT 3.7170 75.0830 3.7350 75.1310 ;
        RECT 4.9590 75.0830 4.9860 75.1310 ;
        RECT 5.1120 75.0830 5.1480 75.1310 ;
        RECT 5.8770 75.0830 5.8950 75.1310 ;
        RECT 9.4410 75.0830 9.4590 75.1310 ;
        RECT 0.1530 76.1630 0.1710 76.2110 ;
        RECT 3.7170 76.1630 3.7350 76.2110 ;
        RECT 4.9590 76.1630 4.9860 76.2110 ;
        RECT 5.1120 76.1630 5.1480 76.2110 ;
        RECT 5.8770 76.1630 5.8950 76.2110 ;
        RECT 9.4410 76.1630 9.4590 76.2110 ;
        RECT 0.1530 77.2430 0.1710 77.2910 ;
        RECT 3.7170 77.2430 3.7350 77.2910 ;
        RECT 4.9590 77.2430 4.9860 77.2910 ;
        RECT 5.1120 77.2430 5.1480 77.2910 ;
        RECT 5.8770 77.2430 5.8950 77.2910 ;
        RECT 9.4410 77.2430 9.4590 77.2910 ;
        RECT 0.1530 78.3230 0.1710 78.3710 ;
        RECT 3.7170 78.3230 3.7350 78.3710 ;
        RECT 4.9590 78.3230 4.9860 78.3710 ;
        RECT 5.1120 78.3230 5.1480 78.3710 ;
        RECT 5.8770 78.3230 5.8950 78.3710 ;
        RECT 9.4410 78.3230 9.4590 78.3710 ;
        RECT 0.1530 79.4030 0.1710 79.4510 ;
        RECT 3.7170 79.4030 3.7350 79.4510 ;
        RECT 4.9590 79.4030 4.9860 79.4510 ;
        RECT 5.1120 79.4030 5.1480 79.4510 ;
        RECT 5.8770 79.4030 5.8950 79.4510 ;
        RECT 9.4410 79.4030 9.4590 79.4510 ;
        RECT 0.1530 80.4830 0.1710 80.5310 ;
        RECT 3.7170 80.4830 3.7350 80.5310 ;
        RECT 4.9590 80.4830 4.9860 80.5310 ;
        RECT 5.1120 80.4830 5.1480 80.5310 ;
        RECT 5.8770 80.4830 5.8950 80.5310 ;
        RECT 9.4410 80.4830 9.4590 80.5310 ;
        RECT 0.1530 81.5630 0.1710 81.6110 ;
        RECT 3.7170 81.5630 3.7350 81.6110 ;
        RECT 4.9590 81.5630 4.9860 81.6110 ;
        RECT 5.1120 81.5630 5.1480 81.6110 ;
        RECT 5.8770 81.5630 5.8950 81.6110 ;
        RECT 9.4410 81.5630 9.4590 81.6110 ;
        RECT 0.1530 82.6430 0.1710 82.6910 ;
        RECT 3.7170 82.6430 3.7350 82.6910 ;
        RECT 4.9590 82.6430 4.9860 82.6910 ;
        RECT 5.1120 82.6430 5.1480 82.6910 ;
        RECT 5.8770 82.6430 5.8950 82.6910 ;
        RECT 9.4410 82.6430 9.4590 82.6910 ;
        RECT 0.1530 83.7230 0.1710 83.7710 ;
        RECT 3.7170 83.7230 3.7350 83.7710 ;
        RECT 4.9590 83.7230 4.9860 83.7710 ;
        RECT 5.1120 83.7230 5.1480 83.7710 ;
        RECT 5.8770 83.7230 5.8950 83.7710 ;
        RECT 9.4410 83.7230 9.4590 83.7710 ;
        RECT 0.1530 84.8030 0.1710 84.8510 ;
        RECT 3.7170 84.8030 3.7350 84.8510 ;
        RECT 4.9590 84.8030 4.9860 84.8510 ;
        RECT 5.1120 84.8030 5.1480 84.8510 ;
        RECT 5.8770 84.8030 5.8950 84.8510 ;
        RECT 9.4410 84.8030 9.4590 84.8510 ;
        RECT 0.1530 85.8830 0.1710 85.9310 ;
        RECT 3.7170 85.8830 3.7350 85.9310 ;
        RECT 4.9590 85.8830 4.9860 85.9310 ;
        RECT 5.1120 85.8830 5.1480 85.9310 ;
        RECT 5.8770 85.8830 5.8950 85.9310 ;
        RECT 9.4410 85.8830 9.4590 85.9310 ;
        RECT 0.1530 86.9630 0.1710 87.0110 ;
        RECT 3.7170 86.9630 3.7350 87.0110 ;
        RECT 4.9590 86.9630 4.9860 87.0110 ;
        RECT 5.1120 86.9630 5.1480 87.0110 ;
        RECT 5.8770 86.9630 5.8950 87.0110 ;
        RECT 9.4410 86.9630 9.4590 87.0110 ;
        RECT 0.1530 88.0430 0.1710 88.0910 ;
        RECT 3.7170 88.0430 3.7350 88.0910 ;
        RECT 4.9590 88.0430 4.9860 88.0910 ;
        RECT 5.1120 88.0430 5.1480 88.0910 ;
        RECT 5.8770 88.0430 5.8950 88.0910 ;
        RECT 9.4410 88.0430 9.4590 88.0910 ;
        RECT 0.1530 89.1230 0.1710 89.1710 ;
        RECT 3.7170 89.1230 3.7350 89.1710 ;
        RECT 4.9590 89.1230 4.9860 89.1710 ;
        RECT 5.1120 89.1230 5.1480 89.1710 ;
        RECT 5.8770 89.1230 5.8950 89.1710 ;
        RECT 9.4410 89.1230 9.4590 89.1710 ;
        RECT 0.1530 90.2030 0.1710 90.2510 ;
        RECT 3.7170 90.2030 3.7350 90.2510 ;
        RECT 4.9590 90.2030 4.9860 90.2510 ;
        RECT 5.1120 90.2030 5.1480 90.2510 ;
        RECT 5.8770 90.2030 5.8950 90.2510 ;
        RECT 9.4410 90.2030 9.4590 90.2510 ;
        RECT 0.1530 91.2830 0.1710 91.3310 ;
        RECT 3.7170 91.2830 3.7350 91.3310 ;
        RECT 4.9590 91.2830 4.9860 91.3310 ;
        RECT 5.1120 91.2830 5.1480 91.3310 ;
        RECT 5.8770 91.2830 5.8950 91.3310 ;
        RECT 9.4410 91.2830 9.4590 91.3310 ;
        RECT 0.1530 92.3630 0.1710 92.4110 ;
        RECT 3.7170 92.3630 3.7350 92.4110 ;
        RECT 4.9590 92.3630 4.9860 92.4110 ;
        RECT 5.1120 92.3630 5.1480 92.4110 ;
        RECT 5.8770 92.3630 5.8950 92.4110 ;
        RECT 9.4410 92.3630 9.4590 92.4110 ;
        RECT 0.1530 93.4430 0.1710 93.4910 ;
        RECT 3.7170 93.4430 3.7350 93.4910 ;
        RECT 4.9590 93.4430 4.9860 93.4910 ;
        RECT 5.1120 93.4430 5.1480 93.4910 ;
        RECT 5.8770 93.4430 5.8950 93.4910 ;
        RECT 9.4410 93.4430 9.4590 93.4910 ;
        RECT 0.1530 94.5230 0.1710 94.5710 ;
        RECT 3.7170 94.5230 3.7350 94.5710 ;
        RECT 4.9590 94.5230 4.9860 94.5710 ;
        RECT 5.1120 94.5230 5.1480 94.5710 ;
        RECT 5.8770 94.5230 5.8950 94.5710 ;
        RECT 9.4410 94.5230 9.4590 94.5710 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.3350 44.6830 7.3530 44.7200 ;
      LAYER M4  ;
        RECT 7.2830 44.6910 7.3670 44.7150 ;
      LAYER M5  ;
        RECT 7.3320 43.7400 7.3560 46.9800 ;
      LAYER V3  ;
        RECT 7.3350 44.6910 7.3530 44.7150 ;
      LAYER V4  ;
        RECT 7.3320 44.6910 7.3560 44.7150 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.1190 44.6860 7.1370 44.7230 ;
      LAYER M4  ;
        RECT 7.0670 44.6910 7.1510 44.7150 ;
      LAYER M5  ;
        RECT 7.1160 43.7400 7.1400 46.9800 ;
      LAYER V3  ;
        RECT 7.1190 44.6910 7.1370 44.7150 ;
      LAYER V4  ;
        RECT 7.1160 44.6910 7.1400 44.7150 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.9030 44.1070 6.9210 44.1440 ;
      LAYER M4  ;
        RECT 6.8510 44.1150 6.9350 44.1390 ;
      LAYER M5  ;
        RECT 6.9000 43.7400 6.9240 46.9800 ;
      LAYER V3  ;
        RECT 6.9030 44.1150 6.9210 44.1390 ;
      LAYER V4  ;
        RECT 6.9000 44.1150 6.9240 44.1390 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.6870 44.3470 6.7050 44.5280 ;
      LAYER M4  ;
        RECT 6.6350 44.4990 6.7190 44.5230 ;
      LAYER M5  ;
        RECT 6.6840 43.7400 6.7080 46.9800 ;
      LAYER V3  ;
        RECT 6.6870 44.4990 6.7050 44.5230 ;
      LAYER V4  ;
        RECT 6.6840 44.4990 6.7080 44.5230 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.4710 44.1100 6.4890 44.1770 ;
      LAYER M4  ;
        RECT 6.4190 44.1150 6.5030 44.1390 ;
      LAYER M5  ;
        RECT 6.4680 43.7400 6.4920 46.9800 ;
      LAYER V3  ;
        RECT 6.4710 44.1150 6.4890 44.1390 ;
      LAYER V4  ;
        RECT 6.4680 44.1150 6.4920 44.1390 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.2550 43.8430 6.2730 44.0960 ;
      LAYER M4  ;
        RECT 6.2030 44.0670 6.2870 44.0910 ;
      LAYER M5  ;
        RECT 6.2520 43.7400 6.2760 46.9800 ;
      LAYER V3  ;
        RECT 6.2550 44.0670 6.2730 44.0910 ;
      LAYER V4  ;
        RECT 6.2520 44.0670 6.2760 44.0910 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.0390 44.8780 6.0570 44.9150 ;
      LAYER M4  ;
        RECT 5.9870 44.8830 6.0710 44.9070 ;
      LAYER M5  ;
        RECT 6.0360 43.7400 6.0600 46.9800 ;
      LAYER V3  ;
        RECT 6.0390 44.8830 6.0570 44.9070 ;
      LAYER V4  ;
        RECT 6.0360 44.8830 6.0600 44.9070 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 5.1750 44.1100 5.1930 44.1770 ;
      LAYER M4  ;
        RECT 4.8910 44.1150 5.2040 44.1390 ;
      LAYER M5  ;
        RECT 4.9020 43.7400 4.9260 46.9800 ;
      LAYER V3  ;
        RECT 5.1750 44.1150 5.1930 44.1390 ;
      LAYER V4  ;
        RECT 4.9020 44.1150 4.9260 44.1390 ;
    END
  END ADDRESS[7]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 4.7790 43.8430 4.7970 44.0960 ;
      LAYER M4  ;
        RECT 4.5670 44.0670 4.8080 44.0910 ;
      LAYER M5  ;
        RECT 4.5780 43.7400 4.6020 46.9800 ;
      LAYER V3  ;
        RECT 4.7790 44.0670 4.7970 44.0910 ;
      LAYER V4  ;
        RECT 4.5780 44.0670 4.6020 44.0910 ;
    END
  END banksel
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.9870 44.1100 4.0050 44.1770 ;
      LAYER M4  ;
        RECT 3.9350 44.1150 4.0190 44.1390 ;
      LAYER M5  ;
        RECT 3.9840 43.7400 4.0080 46.9800 ;
      LAYER V3  ;
        RECT 3.9870 44.1150 4.0050 44.1390 ;
      LAYER V4  ;
        RECT 3.9840 44.1150 4.0080 44.1390 ;
    END
  END write
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.7710 44.9740 3.7890 45.0230 ;
      LAYER M4  ;
        RECT 3.7190 44.9790 3.8030 45.0030 ;
      LAYER M5  ;
        RECT 3.7680 43.7400 3.7920 46.9800 ;
      LAYER V3  ;
        RECT 3.7710 44.9790 3.7890 45.0030 ;
      LAYER V4  ;
        RECT 3.7680 44.9790 3.7920 45.0030 ;
    END
  END clk
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.8070 43.8430 3.8250 44.0960 ;
      LAYER M4  ;
        RECT 3.5410 44.0670 3.8360 44.0910 ;
      LAYER M5  ;
        RECT 3.5520 43.7400 3.5760 46.9800 ;
      LAYER V3  ;
        RECT 3.8070 44.0670 3.8250 44.0910 ;
      LAYER V4  ;
        RECT 3.5520 44.0670 3.5760 44.0910 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.3390 44.6830 3.3570 44.7200 ;
      LAYER M4  ;
        RECT 3.2870 44.6910 3.3710 44.7150 ;
      LAYER M5  ;
        RECT 3.3360 43.7400 3.3600 46.9800 ;
      LAYER V3  ;
        RECT 3.3390 44.6910 3.3570 44.7150 ;
      LAYER V4  ;
        RECT 3.3360 44.6910 3.3600 44.7150 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.1230 44.1100 3.1410 44.3390 ;
      LAYER M4  ;
        RECT 3.0710 44.1150 3.1550 44.1390 ;
      LAYER M5  ;
        RECT 3.1200 43.7400 3.1440 46.9800 ;
      LAYER V3  ;
        RECT 3.1230 44.1150 3.1410 44.1390 ;
      LAYER V4  ;
        RECT 3.1200 44.1150 3.1440 44.1390 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.9070 43.8430 2.9250 44.0960 ;
      LAYER M4  ;
        RECT 2.8550 44.0670 2.9390 44.0910 ;
      LAYER M5  ;
        RECT 2.9040 43.7400 2.9280 46.9800 ;
      LAYER V3  ;
        RECT 2.9070 44.0670 2.9250 44.0910 ;
      LAYER V4  ;
        RECT 2.9040 44.0670 2.9280 44.0910 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.6910 44.1070 2.7090 44.1440 ;
      LAYER M4  ;
        RECT 2.6390 44.1150 2.7230 44.1390 ;
      LAYER M5  ;
        RECT 2.6880 43.7400 2.7120 46.9800 ;
      LAYER V3  ;
        RECT 2.6910 44.1150 2.7090 44.1390 ;
      LAYER V4  ;
        RECT 2.6880 44.1150 2.7120 44.1390 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.4750 44.6830 2.4930 44.7200 ;
      LAYER M4  ;
        RECT 2.4230 44.6910 2.5070 44.7150 ;
      LAYER M5  ;
        RECT 2.4720 43.7400 2.4960 46.9800 ;
      LAYER V3  ;
        RECT 2.4750 44.6910 2.4930 44.7150 ;
      LAYER V4  ;
        RECT 2.4720 44.6910 2.4960 44.7150 ;
    END
  END sdel[4]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 0.4280 5.1360 0.4520 ;
      LAYER M3  ;
        RECT 5.0760 0.3775 5.0940 0.6170 ;
      LAYER V3  ;
        RECT 5.0760 0.4280 5.0940 0.4520 ;
    END
  END dataout[0]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 0.3320 5.2040 0.3560 ;
      LAYER M3  ;
        RECT 4.8510 0.2700 4.8690 0.6750 ;
      LAYER V3  ;
        RECT 4.8510 0.3320 4.8690 0.3560 ;
    END
  END wd[0]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 1.5080 5.1360 1.5320 ;
      LAYER M3  ;
        RECT 5.0760 1.4575 5.0940 1.6970 ;
      LAYER V3  ;
        RECT 5.0760 1.5080 5.0940 1.5320 ;
    END
  END dataout[1]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 1.4120 5.2040 1.4360 ;
      LAYER M3  ;
        RECT 4.8510 1.3500 4.8690 1.7550 ;
      LAYER V3  ;
        RECT 4.8510 1.4120 4.8690 1.4360 ;
    END
  END wd[1]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 2.5880 5.1360 2.6120 ;
      LAYER M3  ;
        RECT 5.0760 2.5375 5.0940 2.7770 ;
      LAYER V3  ;
        RECT 5.0760 2.5880 5.0940 2.6120 ;
    END
  END dataout[2]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 2.4920 5.2040 2.5160 ;
      LAYER M3  ;
        RECT 4.8510 2.4300 4.8690 2.8350 ;
      LAYER V3  ;
        RECT 4.8510 2.4920 4.8690 2.5160 ;
    END
  END wd[2]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 3.6680 5.1360 3.6920 ;
      LAYER M3  ;
        RECT 5.0760 3.6175 5.0940 3.8570 ;
      LAYER V3  ;
        RECT 5.0760 3.6680 5.0940 3.6920 ;
    END
  END dataout[3]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 3.5720 5.2040 3.5960 ;
      LAYER M3  ;
        RECT 4.8510 3.5100 4.8690 3.9150 ;
      LAYER V3  ;
        RECT 4.8510 3.5720 4.8690 3.5960 ;
    END
  END wd[3]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 4.7480 5.1360 4.7720 ;
      LAYER M3  ;
        RECT 5.0760 4.6975 5.0940 4.9370 ;
      LAYER V3  ;
        RECT 5.0760 4.7480 5.0940 4.7720 ;
    END
  END dataout[4]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 4.6520 5.2040 4.6760 ;
      LAYER M3  ;
        RECT 4.8510 4.5900 4.8690 4.9950 ;
      LAYER V3  ;
        RECT 4.8510 4.6520 4.8690 4.6760 ;
    END
  END wd[4]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 5.8280 5.1360 5.8520 ;
      LAYER M3  ;
        RECT 5.0760 5.7775 5.0940 6.0170 ;
      LAYER V3  ;
        RECT 5.0760 5.8280 5.0940 5.8520 ;
    END
  END dataout[5]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 5.7320 5.2040 5.7560 ;
      LAYER M3  ;
        RECT 4.8510 5.6700 4.8690 6.0750 ;
      LAYER V3  ;
        RECT 4.8510 5.7320 4.8690 5.7560 ;
    END
  END wd[5]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 6.9080 5.1360 6.9320 ;
      LAYER M3  ;
        RECT 5.0760 6.8575 5.0940 7.0970 ;
      LAYER V3  ;
        RECT 5.0760 6.9080 5.0940 6.9320 ;
    END
  END dataout[6]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 6.8120 5.2040 6.8360 ;
      LAYER M3  ;
        RECT 4.8510 6.7500 4.8690 7.1550 ;
      LAYER V3  ;
        RECT 4.8510 6.8120 4.8690 6.8360 ;
    END
  END wd[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 7.9880 5.1360 8.0120 ;
      LAYER M3  ;
        RECT 5.0760 7.9375 5.0940 8.1770 ;
      LAYER V3  ;
        RECT 5.0760 7.9880 5.0940 8.0120 ;
    END
  END dataout[7]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 7.8920 5.2040 7.9160 ;
      LAYER M3  ;
        RECT 4.8510 7.8300 4.8690 8.2350 ;
      LAYER V3  ;
        RECT 4.8510 7.8920 4.8690 7.9160 ;
    END
  END wd[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 9.0680 5.1360 9.0920 ;
      LAYER M3  ;
        RECT 5.0760 9.0175 5.0940 9.2570 ;
      LAYER V3  ;
        RECT 5.0760 9.0680 5.0940 9.0920 ;
    END
  END dataout[8]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 8.9720 5.2040 8.9960 ;
      LAYER M3  ;
        RECT 4.8510 8.9100 4.8690 9.3150 ;
      LAYER V3  ;
        RECT 4.8510 8.9720 4.8690 8.9960 ;
    END
  END wd[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 10.1480 5.1360 10.1720 ;
      LAYER M3  ;
        RECT 5.0760 10.0975 5.0940 10.3370 ;
      LAYER V3  ;
        RECT 5.0760 10.1480 5.0940 10.1720 ;
    END
  END dataout[9]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 10.0520 5.2040 10.0760 ;
      LAYER M3  ;
        RECT 4.8510 9.9900 4.8690 10.3950 ;
      LAYER V3  ;
        RECT 4.8510 10.0520 4.8690 10.0760 ;
    END
  END wd[9]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 11.2280 5.1360 11.2520 ;
      LAYER M3  ;
        RECT 5.0760 11.1775 5.0940 11.4170 ;
      LAYER V3  ;
        RECT 5.0760 11.2280 5.0940 11.2520 ;
    END
  END dataout[10]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 11.1320 5.2040 11.1560 ;
      LAYER M3  ;
        RECT 4.8510 11.0700 4.8690 11.4750 ;
      LAYER V3  ;
        RECT 4.8510 11.1320 4.8690 11.1560 ;
    END
  END wd[10]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 12.3080 5.1360 12.3320 ;
      LAYER M3  ;
        RECT 5.0760 12.2575 5.0940 12.4970 ;
      LAYER V3  ;
        RECT 5.0760 12.3080 5.0940 12.3320 ;
    END
  END dataout[11]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 12.2120 5.2040 12.2360 ;
      LAYER M3  ;
        RECT 4.8510 12.1500 4.8690 12.5550 ;
      LAYER V3  ;
        RECT 4.8510 12.2120 4.8690 12.2360 ;
    END
  END wd[11]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 13.3880 5.1360 13.4120 ;
      LAYER M3  ;
        RECT 5.0760 13.3375 5.0940 13.5770 ;
      LAYER V3  ;
        RECT 5.0760 13.3880 5.0940 13.4120 ;
    END
  END dataout[12]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 13.2920 5.2040 13.3160 ;
      LAYER M3  ;
        RECT 4.8510 13.2300 4.8690 13.6350 ;
      LAYER V3  ;
        RECT 4.8510 13.2920 4.8690 13.3160 ;
    END
  END wd[12]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 14.4680 5.1360 14.4920 ;
      LAYER M3  ;
        RECT 5.0760 14.4175 5.0940 14.6570 ;
      LAYER V3  ;
        RECT 5.0760 14.4680 5.0940 14.4920 ;
    END
  END dataout[13]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 14.3720 5.2040 14.3960 ;
      LAYER M3  ;
        RECT 4.8510 14.3100 4.8690 14.7150 ;
      LAYER V3  ;
        RECT 4.8510 14.3720 4.8690 14.3960 ;
    END
  END wd[13]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 15.5480 5.1360 15.5720 ;
      LAYER M3  ;
        RECT 5.0760 15.4975 5.0940 15.7370 ;
      LAYER V3  ;
        RECT 5.0760 15.5480 5.0940 15.5720 ;
    END
  END dataout[14]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 15.4520 5.2040 15.4760 ;
      LAYER M3  ;
        RECT 4.8510 15.3900 4.8690 15.7950 ;
      LAYER V3  ;
        RECT 4.8510 15.4520 4.8690 15.4760 ;
    END
  END wd[14]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 16.6280 5.1360 16.6520 ;
      LAYER M3  ;
        RECT 5.0760 16.5775 5.0940 16.8170 ;
      LAYER V3  ;
        RECT 5.0760 16.6280 5.0940 16.6520 ;
    END
  END dataout[15]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 16.5320 5.2040 16.5560 ;
      LAYER M3  ;
        RECT 4.8510 16.4700 4.8690 16.8750 ;
      LAYER V3  ;
        RECT 4.8510 16.5320 4.8690 16.5560 ;
    END
  END wd[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 17.7080 5.1360 17.7320 ;
      LAYER M3  ;
        RECT 5.0760 17.6575 5.0940 17.8970 ;
      LAYER V3  ;
        RECT 5.0760 17.7080 5.0940 17.7320 ;
    END
  END dataout[16]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 17.6120 5.2040 17.6360 ;
      LAYER M3  ;
        RECT 4.8510 17.5500 4.8690 17.9550 ;
      LAYER V3  ;
        RECT 4.8510 17.6120 4.8690 17.6360 ;
    END
  END wd[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 18.7880 5.1360 18.8120 ;
      LAYER M3  ;
        RECT 5.0760 18.7375 5.0940 18.9770 ;
      LAYER V3  ;
        RECT 5.0760 18.7880 5.0940 18.8120 ;
    END
  END dataout[17]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 18.6920 5.2040 18.7160 ;
      LAYER M3  ;
        RECT 4.8510 18.6300 4.8690 19.0350 ;
      LAYER V3  ;
        RECT 4.8510 18.6920 4.8690 18.7160 ;
    END
  END wd[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 19.8680 5.1360 19.8920 ;
      LAYER M3  ;
        RECT 5.0760 19.8175 5.0940 20.0570 ;
      LAYER V3  ;
        RECT 5.0760 19.8680 5.0940 19.8920 ;
    END
  END dataout[18]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 19.7720 5.2040 19.7960 ;
      LAYER M3  ;
        RECT 4.8510 19.7100 4.8690 20.1150 ;
      LAYER V3  ;
        RECT 4.8510 19.7720 4.8690 19.7960 ;
    END
  END wd[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 20.9480 5.1360 20.9720 ;
      LAYER M3  ;
        RECT 5.0760 20.8975 5.0940 21.1370 ;
      LAYER V3  ;
        RECT 5.0760 20.9480 5.0940 20.9720 ;
    END
  END dataout[19]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 20.8520 5.2040 20.8760 ;
      LAYER M3  ;
        RECT 4.8510 20.7900 4.8690 21.1950 ;
      LAYER V3  ;
        RECT 4.8510 20.8520 4.8690 20.8760 ;
    END
  END wd[19]
  PIN dataout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 22.0280 5.1360 22.0520 ;
      LAYER M3  ;
        RECT 5.0760 21.9775 5.0940 22.2170 ;
      LAYER V3  ;
        RECT 5.0760 22.0280 5.0940 22.0520 ;
    END
  END dataout[20]
  PIN wd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 21.9320 5.2040 21.9560 ;
      LAYER M3  ;
        RECT 4.8510 21.8700 4.8690 22.2750 ;
      LAYER V3  ;
        RECT 4.8510 21.9320 4.8690 21.9560 ;
    END
  END wd[20]
  PIN dataout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 23.1080 5.1360 23.1320 ;
      LAYER M3  ;
        RECT 5.0760 23.0575 5.0940 23.2970 ;
      LAYER V3  ;
        RECT 5.0760 23.1080 5.0940 23.1320 ;
    END
  END dataout[21]
  PIN wd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 23.0120 5.2040 23.0360 ;
      LAYER M3  ;
        RECT 4.8510 22.9500 4.8690 23.3550 ;
      LAYER V3  ;
        RECT 4.8510 23.0120 4.8690 23.0360 ;
    END
  END wd[21]
  PIN dataout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 24.1880 5.1360 24.2120 ;
      LAYER M3  ;
        RECT 5.0760 24.1375 5.0940 24.3770 ;
      LAYER V3  ;
        RECT 5.0760 24.1880 5.0940 24.2120 ;
    END
  END dataout[22]
  PIN wd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 24.0920 5.2040 24.1160 ;
      LAYER M3  ;
        RECT 4.8510 24.0300 4.8690 24.4350 ;
      LAYER V3  ;
        RECT 4.8510 24.0920 4.8690 24.1160 ;
    END
  END wd[22]
  PIN dataout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 25.2680 5.1360 25.2920 ;
      LAYER M3  ;
        RECT 5.0760 25.2175 5.0940 25.4570 ;
      LAYER V3  ;
        RECT 5.0760 25.2680 5.0940 25.2920 ;
    END
  END dataout[23]
  PIN wd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 25.1720 5.2040 25.1960 ;
      LAYER M3  ;
        RECT 4.8510 25.1100 4.8690 25.5150 ;
      LAYER V3  ;
        RECT 4.8510 25.1720 4.8690 25.1960 ;
    END
  END wd[23]
  PIN dataout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 26.3480 5.1360 26.3720 ;
      LAYER M3  ;
        RECT 5.0760 26.2975 5.0940 26.5370 ;
      LAYER V3  ;
        RECT 5.0760 26.3480 5.0940 26.3720 ;
    END
  END dataout[24]
  PIN wd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 26.2520 5.2040 26.2760 ;
      LAYER M3  ;
        RECT 4.8510 26.1900 4.8690 26.5950 ;
      LAYER V3  ;
        RECT 4.8510 26.2520 4.8690 26.2760 ;
    END
  END wd[24]
  PIN dataout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 27.4280 5.1360 27.4520 ;
      LAYER M3  ;
        RECT 5.0760 27.3775 5.0940 27.6170 ;
      LAYER V3  ;
        RECT 5.0760 27.4280 5.0940 27.4520 ;
    END
  END dataout[25]
  PIN wd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 27.3320 5.2040 27.3560 ;
      LAYER M3  ;
        RECT 4.8510 27.2700 4.8690 27.6750 ;
      LAYER V3  ;
        RECT 4.8510 27.3320 4.8690 27.3560 ;
    END
  END wd[25]
  PIN dataout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 28.5080 5.1360 28.5320 ;
      LAYER M3  ;
        RECT 5.0760 28.4575 5.0940 28.6970 ;
      LAYER V3  ;
        RECT 5.0760 28.5080 5.0940 28.5320 ;
    END
  END dataout[26]
  PIN wd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 28.4120 5.2040 28.4360 ;
      LAYER M3  ;
        RECT 4.8510 28.3500 4.8690 28.7550 ;
      LAYER V3  ;
        RECT 4.8510 28.4120 4.8690 28.4360 ;
    END
  END wd[26]
  PIN dataout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 29.5880 5.1360 29.6120 ;
      LAYER M3  ;
        RECT 5.0760 29.5375 5.0940 29.7770 ;
      LAYER V3  ;
        RECT 5.0760 29.5880 5.0940 29.6120 ;
    END
  END dataout[27]
  PIN wd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 29.4920 5.2040 29.5160 ;
      LAYER M3  ;
        RECT 4.8510 29.4300 4.8690 29.8350 ;
      LAYER V3  ;
        RECT 4.8510 29.4920 4.8690 29.5160 ;
    END
  END wd[27]
  PIN dataout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 30.6680 5.1360 30.6920 ;
      LAYER M3  ;
        RECT 5.0760 30.6175 5.0940 30.8570 ;
      LAYER V3  ;
        RECT 5.0760 30.6680 5.0940 30.6920 ;
    END
  END dataout[28]
  PIN wd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 30.5720 5.2040 30.5960 ;
      LAYER M3  ;
        RECT 4.8510 30.5100 4.8690 30.9150 ;
      LAYER V3  ;
        RECT 4.8510 30.5720 4.8690 30.5960 ;
    END
  END wd[28]
  PIN dataout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 31.7480 5.1360 31.7720 ;
      LAYER M3  ;
        RECT 5.0760 31.6975 5.0940 31.9370 ;
      LAYER V3  ;
        RECT 5.0760 31.7480 5.0940 31.7720 ;
    END
  END dataout[29]
  PIN wd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 31.6520 5.2040 31.6760 ;
      LAYER M3  ;
        RECT 4.8510 31.5900 4.8690 31.9950 ;
      LAYER V3  ;
        RECT 4.8510 31.6520 4.8690 31.6760 ;
    END
  END wd[29]
  PIN dataout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 32.8280 5.1360 32.8520 ;
      LAYER M3  ;
        RECT 5.0760 32.7775 5.0940 33.0170 ;
      LAYER V3  ;
        RECT 5.0760 32.8280 5.0940 32.8520 ;
    END
  END dataout[30]
  PIN wd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 32.7320 5.2040 32.7560 ;
      LAYER M3  ;
        RECT 4.8510 32.6700 4.8690 33.0750 ;
      LAYER V3  ;
        RECT 4.8510 32.7320 4.8690 32.7560 ;
    END
  END wd[30]
  PIN dataout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 33.9080 5.1360 33.9320 ;
      LAYER M3  ;
        RECT 5.0760 33.8575 5.0940 34.0970 ;
      LAYER V3  ;
        RECT 5.0760 33.9080 5.0940 33.9320 ;
    END
  END dataout[31]
  PIN wd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 33.8120 5.2040 33.8360 ;
      LAYER M3  ;
        RECT 4.8510 33.7500 4.8690 34.1550 ;
      LAYER V3  ;
        RECT 4.8510 33.8120 4.8690 33.8360 ;
    END
  END wd[31]
  PIN dataout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 34.9880 5.1360 35.0120 ;
      LAYER M3  ;
        RECT 5.0760 34.9375 5.0940 35.1770 ;
      LAYER V3  ;
        RECT 5.0760 34.9880 5.0940 35.0120 ;
    END
  END dataout[32]
  PIN wd[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 34.8920 5.2040 34.9160 ;
      LAYER M3  ;
        RECT 4.8510 34.8300 4.8690 35.2350 ;
      LAYER V3  ;
        RECT 4.8510 34.8920 4.8690 34.9160 ;
    END
  END wd[32]
  PIN dataout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 36.0680 5.1360 36.0920 ;
      LAYER M3  ;
        RECT 5.0760 36.0175 5.0940 36.2570 ;
      LAYER V3  ;
        RECT 5.0760 36.0680 5.0940 36.0920 ;
    END
  END dataout[33]
  PIN wd[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 35.9720 5.2040 35.9960 ;
      LAYER M3  ;
        RECT 4.8510 35.9100 4.8690 36.3150 ;
      LAYER V3  ;
        RECT 4.8510 35.9720 4.8690 35.9960 ;
    END
  END wd[33]
  PIN dataout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 37.1480 5.1360 37.1720 ;
      LAYER M3  ;
        RECT 5.0760 37.0975 5.0940 37.3370 ;
      LAYER V3  ;
        RECT 5.0760 37.1480 5.0940 37.1720 ;
    END
  END dataout[34]
  PIN wd[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 37.0520 5.2040 37.0760 ;
      LAYER M3  ;
        RECT 4.8510 36.9900 4.8690 37.3950 ;
      LAYER V3  ;
        RECT 4.8510 37.0520 4.8690 37.0760 ;
    END
  END wd[34]
  PIN dataout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 38.2280 5.1360 38.2520 ;
      LAYER M3  ;
        RECT 5.0760 38.1775 5.0940 38.4170 ;
      LAYER V3  ;
        RECT 5.0760 38.2280 5.0940 38.2520 ;
    END
  END dataout[35]
  PIN wd[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 38.1320 5.2040 38.1560 ;
      LAYER M3  ;
        RECT 4.8510 38.0700 4.8690 38.4750 ;
      LAYER V3  ;
        RECT 4.8510 38.1320 4.8690 38.1560 ;
    END
  END wd[35]
  PIN dataout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 39.3080 5.1360 39.3320 ;
      LAYER M3  ;
        RECT 5.0760 39.2575 5.0940 39.4970 ;
      LAYER V3  ;
        RECT 5.0760 39.3080 5.0940 39.3320 ;
    END
  END dataout[36]
  PIN wd[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 39.2120 5.2040 39.2360 ;
      LAYER M3  ;
        RECT 4.8510 39.1500 4.8690 39.5550 ;
      LAYER V3  ;
        RECT 4.8510 39.2120 4.8690 39.2360 ;
    END
  END wd[36]
  PIN dataout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 40.3880 5.1360 40.4120 ;
      LAYER M3  ;
        RECT 5.0760 40.3375 5.0940 40.5770 ;
      LAYER V3  ;
        RECT 5.0760 40.3880 5.0940 40.4120 ;
    END
  END dataout[37]
  PIN wd[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 40.2920 5.2040 40.3160 ;
      LAYER M3  ;
        RECT 4.8510 40.2300 4.8690 40.6350 ;
      LAYER V3  ;
        RECT 4.8510 40.2920 4.8690 40.3160 ;
    END
  END wd[37]
  PIN dataout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 41.4680 5.1360 41.4920 ;
      LAYER M3  ;
        RECT 5.0760 41.4175 5.0940 41.6570 ;
      LAYER V3  ;
        RECT 5.0760 41.4680 5.0940 41.4920 ;
    END
  END dataout[38]
  PIN wd[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 41.3720 5.2040 41.3960 ;
      LAYER M3  ;
        RECT 4.8510 41.3100 4.8690 41.7150 ;
      LAYER V3  ;
        RECT 4.8510 41.3720 4.8690 41.3960 ;
    END
  END wd[38]
  PIN dataout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 42.5480 5.1360 42.5720 ;
      LAYER M3  ;
        RECT 5.0760 42.4975 5.0940 42.7370 ;
      LAYER V3  ;
        RECT 5.0760 42.5480 5.0940 42.5720 ;
    END
  END dataout[39]
  PIN wd[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 42.4520 5.2040 42.4760 ;
      LAYER M3  ;
        RECT 4.8510 42.3900 4.8690 42.7950 ;
      LAYER V3  ;
        RECT 4.8510 42.4520 4.8690 42.4760 ;
    END
  END wd[39]
  PIN dataout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 51.7550 5.1360 51.7790 ;
      LAYER M3  ;
        RECT 5.0760 51.7045 5.0940 51.9440 ;
      LAYER V3  ;
        RECT 5.0760 51.7550 5.0940 51.7790 ;
    END
  END dataout[40]
  PIN wd[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 51.6590 5.2040 51.6830 ;
      LAYER M3  ;
        RECT 4.8510 51.5970 4.8690 52.0020 ;
      LAYER V3  ;
        RECT 4.8510 51.6590 4.8690 51.6830 ;
    END
  END wd[40]
  PIN dataout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 52.8350 5.1360 52.8590 ;
      LAYER M3  ;
        RECT 5.0760 52.7845 5.0940 53.0240 ;
      LAYER V3  ;
        RECT 5.0760 52.8350 5.0940 52.8590 ;
    END
  END dataout[41]
  PIN wd[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 52.7390 5.2040 52.7630 ;
      LAYER M3  ;
        RECT 4.8510 52.6770 4.8690 53.0820 ;
      LAYER V3  ;
        RECT 4.8510 52.7390 4.8690 52.7630 ;
    END
  END wd[41]
  PIN dataout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 53.9150 5.1360 53.9390 ;
      LAYER M3  ;
        RECT 5.0760 53.8645 5.0940 54.1040 ;
      LAYER V3  ;
        RECT 5.0760 53.9150 5.0940 53.9390 ;
    END
  END dataout[42]
  PIN wd[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 53.8190 5.2040 53.8430 ;
      LAYER M3  ;
        RECT 4.8510 53.7570 4.8690 54.1620 ;
      LAYER V3  ;
        RECT 4.8510 53.8190 4.8690 53.8430 ;
    END
  END wd[42]
  PIN dataout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 54.9950 5.1360 55.0190 ;
      LAYER M3  ;
        RECT 5.0760 54.9445 5.0940 55.1840 ;
      LAYER V3  ;
        RECT 5.0760 54.9950 5.0940 55.0190 ;
    END
  END dataout[43]
  PIN wd[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 54.8990 5.2040 54.9230 ;
      LAYER M3  ;
        RECT 4.8510 54.8370 4.8690 55.2420 ;
      LAYER V3  ;
        RECT 4.8510 54.8990 4.8690 54.9230 ;
    END
  END wd[43]
  PIN dataout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 56.0750 5.1360 56.0990 ;
      LAYER M3  ;
        RECT 5.0760 56.0245 5.0940 56.2640 ;
      LAYER V3  ;
        RECT 5.0760 56.0750 5.0940 56.0990 ;
    END
  END dataout[44]
  PIN wd[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 55.9790 5.2040 56.0030 ;
      LAYER M3  ;
        RECT 4.8510 55.9170 4.8690 56.3220 ;
      LAYER V3  ;
        RECT 4.8510 55.9790 4.8690 56.0030 ;
    END
  END wd[44]
  PIN dataout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 57.1550 5.1360 57.1790 ;
      LAYER M3  ;
        RECT 5.0760 57.1045 5.0940 57.3440 ;
      LAYER V3  ;
        RECT 5.0760 57.1550 5.0940 57.1790 ;
    END
  END dataout[45]
  PIN wd[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 57.0590 5.2040 57.0830 ;
      LAYER M3  ;
        RECT 4.8510 56.9970 4.8690 57.4020 ;
      LAYER V3  ;
        RECT 4.8510 57.0590 4.8690 57.0830 ;
    END
  END wd[45]
  PIN dataout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 58.2350 5.1360 58.2590 ;
      LAYER M3  ;
        RECT 5.0760 58.1845 5.0940 58.4240 ;
      LAYER V3  ;
        RECT 5.0760 58.2350 5.0940 58.2590 ;
    END
  END dataout[46]
  PIN wd[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 58.1390 5.2040 58.1630 ;
      LAYER M3  ;
        RECT 4.8510 58.0770 4.8690 58.4820 ;
      LAYER V3  ;
        RECT 4.8510 58.1390 4.8690 58.1630 ;
    END
  END wd[46]
  PIN dataout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 59.3150 5.1360 59.3390 ;
      LAYER M3  ;
        RECT 5.0760 59.2645 5.0940 59.5040 ;
      LAYER V3  ;
        RECT 5.0760 59.3150 5.0940 59.3390 ;
    END
  END dataout[47]
  PIN wd[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 59.2190 5.2040 59.2430 ;
      LAYER M3  ;
        RECT 4.8510 59.1570 4.8690 59.5620 ;
      LAYER V3  ;
        RECT 4.8510 59.2190 4.8690 59.2430 ;
    END
  END wd[47]
  PIN dataout[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 60.3950 5.1360 60.4190 ;
      LAYER M3  ;
        RECT 5.0760 60.3445 5.0940 60.5840 ;
      LAYER V3  ;
        RECT 5.0760 60.3950 5.0940 60.4190 ;
    END
  END dataout[48]
  PIN wd[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 60.2990 5.2040 60.3230 ;
      LAYER M3  ;
        RECT 4.8510 60.2370 4.8690 60.6420 ;
      LAYER V3  ;
        RECT 4.8510 60.2990 4.8690 60.3230 ;
    END
  END wd[48]
  PIN dataout[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 61.4750 5.1360 61.4990 ;
      LAYER M3  ;
        RECT 5.0760 61.4245 5.0940 61.6640 ;
      LAYER V3  ;
        RECT 5.0760 61.4750 5.0940 61.4990 ;
    END
  END dataout[49]
  PIN wd[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 61.3790 5.2040 61.4030 ;
      LAYER M3  ;
        RECT 4.8510 61.3170 4.8690 61.7220 ;
      LAYER V3  ;
        RECT 4.8510 61.3790 4.8690 61.4030 ;
    END
  END wd[49]
  PIN dataout[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 62.5550 5.1360 62.5790 ;
      LAYER M3  ;
        RECT 5.0760 62.5045 5.0940 62.7440 ;
      LAYER V3  ;
        RECT 5.0760 62.5550 5.0940 62.5790 ;
    END
  END dataout[50]
  PIN wd[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 62.4590 5.2040 62.4830 ;
      LAYER M3  ;
        RECT 4.8510 62.3970 4.8690 62.8020 ;
      LAYER V3  ;
        RECT 4.8510 62.4590 4.8690 62.4830 ;
    END
  END wd[50]
  PIN dataout[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 63.6350 5.1360 63.6590 ;
      LAYER M3  ;
        RECT 5.0760 63.5845 5.0940 63.8240 ;
      LAYER V3  ;
        RECT 5.0760 63.6350 5.0940 63.6590 ;
    END
  END dataout[51]
  PIN wd[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 63.5390 5.2040 63.5630 ;
      LAYER M3  ;
        RECT 4.8510 63.4770 4.8690 63.8820 ;
      LAYER V3  ;
        RECT 4.8510 63.5390 4.8690 63.5630 ;
    END
  END wd[51]
  PIN dataout[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 64.7150 5.1360 64.7390 ;
      LAYER M3  ;
        RECT 5.0760 64.6645 5.0940 64.9040 ;
      LAYER V3  ;
        RECT 5.0760 64.7150 5.0940 64.7390 ;
    END
  END dataout[52]
  PIN wd[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 64.6190 5.2040 64.6430 ;
      LAYER M3  ;
        RECT 4.8510 64.5570 4.8690 64.9620 ;
      LAYER V3  ;
        RECT 4.8510 64.6190 4.8690 64.6430 ;
    END
  END wd[52]
  PIN dataout[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 65.7950 5.1360 65.8190 ;
      LAYER M3  ;
        RECT 5.0760 65.7445 5.0940 65.9840 ;
      LAYER V3  ;
        RECT 5.0760 65.7950 5.0940 65.8190 ;
    END
  END dataout[53]
  PIN wd[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 65.6990 5.2040 65.7230 ;
      LAYER M3  ;
        RECT 4.8510 65.6370 4.8690 66.0420 ;
      LAYER V3  ;
        RECT 4.8510 65.6990 4.8690 65.7230 ;
    END
  END wd[53]
  PIN dataout[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 66.8750 5.1360 66.8990 ;
      LAYER M3  ;
        RECT 5.0760 66.8245 5.0940 67.0640 ;
      LAYER V3  ;
        RECT 5.0760 66.8750 5.0940 66.8990 ;
    END
  END dataout[54]
  PIN wd[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 66.7790 5.2040 66.8030 ;
      LAYER M3  ;
        RECT 4.8510 66.7170 4.8690 67.1220 ;
      LAYER V3  ;
        RECT 4.8510 66.7790 4.8690 66.8030 ;
    END
  END wd[54]
  PIN dataout[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 67.9550 5.1360 67.9790 ;
      LAYER M3  ;
        RECT 5.0760 67.9045 5.0940 68.1440 ;
      LAYER V3  ;
        RECT 5.0760 67.9550 5.0940 67.9790 ;
    END
  END dataout[55]
  PIN wd[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 67.8590 5.2040 67.8830 ;
      LAYER M3  ;
        RECT 4.8510 67.7970 4.8690 68.2020 ;
      LAYER V3  ;
        RECT 4.8510 67.8590 4.8690 67.8830 ;
    END
  END wd[55]
  PIN dataout[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 69.0350 5.1360 69.0590 ;
      LAYER M3  ;
        RECT 5.0760 68.9845 5.0940 69.2240 ;
      LAYER V3  ;
        RECT 5.0760 69.0350 5.0940 69.0590 ;
    END
  END dataout[56]
  PIN wd[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 68.9390 5.2040 68.9630 ;
      LAYER M3  ;
        RECT 4.8510 68.8770 4.8690 69.2820 ;
      LAYER V3  ;
        RECT 4.8510 68.9390 4.8690 68.9630 ;
    END
  END wd[56]
  PIN dataout[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 70.1150 5.1360 70.1390 ;
      LAYER M3  ;
        RECT 5.0760 70.0645 5.0940 70.3040 ;
      LAYER V3  ;
        RECT 5.0760 70.1150 5.0940 70.1390 ;
    END
  END dataout[57]
  PIN wd[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 70.0190 5.2040 70.0430 ;
      LAYER M3  ;
        RECT 4.8510 69.9570 4.8690 70.3620 ;
      LAYER V3  ;
        RECT 4.8510 70.0190 4.8690 70.0430 ;
    END
  END wd[57]
  PIN dataout[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 71.1950 5.1360 71.2190 ;
      LAYER M3  ;
        RECT 5.0760 71.1445 5.0940 71.3840 ;
      LAYER V3  ;
        RECT 5.0760 71.1950 5.0940 71.2190 ;
    END
  END dataout[58]
  PIN wd[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 71.0990 5.2040 71.1230 ;
      LAYER M3  ;
        RECT 4.8510 71.0370 4.8690 71.4420 ;
      LAYER V3  ;
        RECT 4.8510 71.0990 4.8690 71.1230 ;
    END
  END wd[58]
  PIN dataout[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 72.2750 5.1360 72.2990 ;
      LAYER M3  ;
        RECT 5.0760 72.2245 5.0940 72.4640 ;
      LAYER V3  ;
        RECT 5.0760 72.2750 5.0940 72.2990 ;
    END
  END dataout[59]
  PIN wd[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 72.1790 5.2040 72.2030 ;
      LAYER M3  ;
        RECT 4.8510 72.1170 4.8690 72.5220 ;
      LAYER V3  ;
        RECT 4.8510 72.1790 4.8690 72.2030 ;
    END
  END wd[59]
  PIN dataout[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 73.3550 5.1360 73.3790 ;
      LAYER M3  ;
        RECT 5.0760 73.3045 5.0940 73.5440 ;
      LAYER V3  ;
        RECT 5.0760 73.3550 5.0940 73.3790 ;
    END
  END dataout[60]
  PIN wd[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 73.2590 5.2040 73.2830 ;
      LAYER M3  ;
        RECT 4.8510 73.1970 4.8690 73.6020 ;
      LAYER V3  ;
        RECT 4.8510 73.2590 4.8690 73.2830 ;
    END
  END wd[60]
  PIN dataout[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 74.4350 5.1360 74.4590 ;
      LAYER M3  ;
        RECT 5.0760 74.3845 5.0940 74.6240 ;
      LAYER V3  ;
        RECT 5.0760 74.4350 5.0940 74.4590 ;
    END
  END dataout[61]
  PIN wd[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 74.3390 5.2040 74.3630 ;
      LAYER M3  ;
        RECT 4.8510 74.2770 4.8690 74.6820 ;
      LAYER V3  ;
        RECT 4.8510 74.3390 4.8690 74.3630 ;
    END
  END wd[61]
  PIN dataout[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 75.5150 5.1360 75.5390 ;
      LAYER M3  ;
        RECT 5.0760 75.4645 5.0940 75.7040 ;
      LAYER V3  ;
        RECT 5.0760 75.5150 5.0940 75.5390 ;
    END
  END dataout[62]
  PIN wd[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 75.4190 5.2040 75.4430 ;
      LAYER M3  ;
        RECT 4.8510 75.3570 4.8690 75.7620 ;
      LAYER V3  ;
        RECT 4.8510 75.4190 4.8690 75.4430 ;
    END
  END wd[62]
  PIN dataout[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 76.5950 5.1360 76.6190 ;
      LAYER M3  ;
        RECT 5.0760 76.5445 5.0940 76.7840 ;
      LAYER V3  ;
        RECT 5.0760 76.5950 5.0940 76.6190 ;
    END
  END dataout[63]
  PIN wd[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 76.4990 5.2040 76.5230 ;
      LAYER M3  ;
        RECT 4.8510 76.4370 4.8690 76.8420 ;
      LAYER V3  ;
        RECT 4.8510 76.4990 4.8690 76.5230 ;
    END
  END wd[63]
  PIN dataout[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 77.6750 5.1360 77.6990 ;
      LAYER M3  ;
        RECT 5.0760 77.6245 5.0940 77.8640 ;
      LAYER V3  ;
        RECT 5.0760 77.6750 5.0940 77.6990 ;
    END
  END dataout[64]
  PIN wd[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 77.5790 5.2040 77.6030 ;
      LAYER M3  ;
        RECT 4.8510 77.5170 4.8690 77.9220 ;
      LAYER V3  ;
        RECT 4.8510 77.5790 4.8690 77.6030 ;
    END
  END wd[64]
  PIN dataout[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 78.7550 5.1360 78.7790 ;
      LAYER M3  ;
        RECT 5.0760 78.7045 5.0940 78.9440 ;
      LAYER V3  ;
        RECT 5.0760 78.7550 5.0940 78.7790 ;
    END
  END dataout[65]
  PIN wd[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 78.6590 5.2040 78.6830 ;
      LAYER M3  ;
        RECT 4.8510 78.5970 4.8690 79.0020 ;
      LAYER V3  ;
        RECT 4.8510 78.6590 4.8690 78.6830 ;
    END
  END wd[65]
  PIN dataout[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 79.8350 5.1360 79.8590 ;
      LAYER M3  ;
        RECT 5.0760 79.7845 5.0940 80.0240 ;
      LAYER V3  ;
        RECT 5.0760 79.8350 5.0940 79.8590 ;
    END
  END dataout[66]
  PIN wd[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 79.7390 5.2040 79.7630 ;
      LAYER M3  ;
        RECT 4.8510 79.6770 4.8690 80.0820 ;
      LAYER V3  ;
        RECT 4.8510 79.7390 4.8690 79.7630 ;
    END
  END wd[66]
  PIN dataout[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 80.9150 5.1360 80.9390 ;
      LAYER M3  ;
        RECT 5.0760 80.8645 5.0940 81.1040 ;
      LAYER V3  ;
        RECT 5.0760 80.9150 5.0940 80.9390 ;
    END
  END dataout[67]
  PIN wd[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 80.8190 5.2040 80.8430 ;
      LAYER M3  ;
        RECT 4.8510 80.7570 4.8690 81.1620 ;
      LAYER V3  ;
        RECT 4.8510 80.8190 4.8690 80.8430 ;
    END
  END wd[67]
  PIN dataout[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 81.9950 5.1360 82.0190 ;
      LAYER M3  ;
        RECT 5.0760 81.9445 5.0940 82.1840 ;
      LAYER V3  ;
        RECT 5.0760 81.9950 5.0940 82.0190 ;
    END
  END dataout[68]
  PIN wd[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 81.8990 5.2040 81.9230 ;
      LAYER M3  ;
        RECT 4.8510 81.8370 4.8690 82.2420 ;
      LAYER V3  ;
        RECT 4.8510 81.8990 4.8690 81.9230 ;
    END
  END wd[68]
  PIN dataout[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 83.0750 5.1360 83.0990 ;
      LAYER M3  ;
        RECT 5.0760 83.0245 5.0940 83.2640 ;
      LAYER V3  ;
        RECT 5.0760 83.0750 5.0940 83.0990 ;
    END
  END dataout[69]
  PIN wd[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 82.9790 5.2040 83.0030 ;
      LAYER M3  ;
        RECT 4.8510 82.9170 4.8690 83.3220 ;
      LAYER V3  ;
        RECT 4.8510 82.9790 4.8690 83.0030 ;
    END
  END wd[69]
  PIN dataout[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 84.1550 5.1360 84.1790 ;
      LAYER M3  ;
        RECT 5.0760 84.1045 5.0940 84.3440 ;
      LAYER V3  ;
        RECT 5.0760 84.1550 5.0940 84.1790 ;
    END
  END dataout[70]
  PIN wd[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 84.0590 5.2040 84.0830 ;
      LAYER M3  ;
        RECT 4.8510 83.9970 4.8690 84.4020 ;
      LAYER V3  ;
        RECT 4.8510 84.0590 4.8690 84.0830 ;
    END
  END wd[70]
  PIN dataout[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 85.2350 5.1360 85.2590 ;
      LAYER M3  ;
        RECT 5.0760 85.1845 5.0940 85.4240 ;
      LAYER V3  ;
        RECT 5.0760 85.2350 5.0940 85.2590 ;
    END
  END dataout[71]
  PIN wd[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 85.1390 5.2040 85.1630 ;
      LAYER M3  ;
        RECT 4.8510 85.0770 4.8690 85.4820 ;
      LAYER V3  ;
        RECT 4.8510 85.1390 4.8690 85.1630 ;
    END
  END wd[71]
  PIN dataout[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 86.3150 5.1360 86.3390 ;
      LAYER M3  ;
        RECT 5.0760 86.2645 5.0940 86.5040 ;
      LAYER V3  ;
        RECT 5.0760 86.3150 5.0940 86.3390 ;
    END
  END dataout[72]
  PIN wd[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 86.2190 5.2040 86.2430 ;
      LAYER M3  ;
        RECT 4.8510 86.1570 4.8690 86.5620 ;
      LAYER V3  ;
        RECT 4.8510 86.2190 4.8690 86.2430 ;
    END
  END wd[72]
  PIN dataout[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 87.3950 5.1360 87.4190 ;
      LAYER M3  ;
        RECT 5.0760 87.3445 5.0940 87.5840 ;
      LAYER V3  ;
        RECT 5.0760 87.3950 5.0940 87.4190 ;
    END
  END dataout[73]
  PIN wd[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 87.2990 5.2040 87.3230 ;
      LAYER M3  ;
        RECT 4.8510 87.2370 4.8690 87.6420 ;
      LAYER V3  ;
        RECT 4.8510 87.2990 4.8690 87.3230 ;
    END
  END wd[73]
  PIN dataout[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 88.4750 5.1360 88.4990 ;
      LAYER M3  ;
        RECT 5.0760 88.4245 5.0940 88.6640 ;
      LAYER V3  ;
        RECT 5.0760 88.4750 5.0940 88.4990 ;
    END
  END dataout[74]
  PIN wd[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 88.3790 5.2040 88.4030 ;
      LAYER M3  ;
        RECT 4.8510 88.3170 4.8690 88.7220 ;
      LAYER V3  ;
        RECT 4.8510 88.3790 4.8690 88.4030 ;
    END
  END wd[74]
  PIN dataout[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 89.5550 5.1360 89.5790 ;
      LAYER M3  ;
        RECT 5.0760 89.5045 5.0940 89.7440 ;
      LAYER V3  ;
        RECT 5.0760 89.5550 5.0940 89.5790 ;
    END
  END dataout[75]
  PIN wd[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 89.4590 5.2040 89.4830 ;
      LAYER M3  ;
        RECT 4.8510 89.3970 4.8690 89.8020 ;
      LAYER V3  ;
        RECT 4.8510 89.4590 4.8690 89.4830 ;
    END
  END wd[75]
  PIN dataout[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 90.6350 5.1360 90.6590 ;
      LAYER M3  ;
        RECT 5.0760 90.5845 5.0940 90.8240 ;
      LAYER V3  ;
        RECT 5.0760 90.6350 5.0940 90.6590 ;
    END
  END dataout[76]
  PIN wd[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 90.5390 5.2040 90.5630 ;
      LAYER M3  ;
        RECT 4.8510 90.4770 4.8690 90.8820 ;
      LAYER V3  ;
        RECT 4.8510 90.5390 4.8690 90.5630 ;
    END
  END wd[76]
  PIN dataout[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 91.7150 5.1360 91.7390 ;
      LAYER M3  ;
        RECT 5.0760 91.6645 5.0940 91.9040 ;
      LAYER V3  ;
        RECT 5.0760 91.7150 5.0940 91.7390 ;
    END
  END dataout[77]
  PIN wd[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 91.6190 5.2040 91.6430 ;
      LAYER M3  ;
        RECT 4.8510 91.5570 4.8690 91.9620 ;
      LAYER V3  ;
        RECT 4.8510 91.6190 4.8690 91.6430 ;
    END
  END wd[77]
  PIN dataout[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 92.7950 5.1360 92.8190 ;
      LAYER M3  ;
        RECT 5.0760 92.7445 5.0940 92.9840 ;
      LAYER V3  ;
        RECT 5.0760 92.7950 5.0940 92.8190 ;
    END
  END dataout[78]
  PIN wd[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 92.6990 5.2040 92.7230 ;
      LAYER M3  ;
        RECT 4.8510 92.6370 4.8690 93.0420 ;
      LAYER V3  ;
        RECT 4.8510 92.6990 4.8690 92.7230 ;
    END
  END wd[78]
  PIN dataout[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 93.8750 5.1360 93.8990 ;
      LAYER M3  ;
        RECT 5.0760 93.8245 5.0940 94.0640 ;
      LAYER V3  ;
        RECT 5.0760 93.8750 5.0940 93.8990 ;
    END
  END dataout[79]
  PIN wd[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 93.7790 5.2040 93.8030 ;
      LAYER M3  ;
        RECT 4.8510 93.7170 4.8690 94.1220 ;
      LAYER V3  ;
        RECT 4.8510 93.7790 4.8690 93.8030 ;
    END
  END wd[79]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5365 9.6120 18.6300 ;
      RECT 0.0000 18.6165 9.6120 19.7100 ;
      RECT 0.0000 19.6965 9.6120 20.7900 ;
      RECT 0.0000 20.7765 9.6120 21.8700 ;
      RECT 0.0000 21.8565 9.6120 22.9500 ;
      RECT 0.0000 22.9365 9.6120 24.0300 ;
      RECT 0.0000 24.0165 9.6120 25.1100 ;
      RECT 0.0000 25.0965 9.6120 26.1900 ;
      RECT 0.0000 26.1765 9.6120 27.2700 ;
      RECT 0.0000 27.2565 9.6120 28.3500 ;
      RECT 0.0000 28.3365 9.6120 29.4300 ;
      RECT 0.0000 29.4165 9.6120 30.5100 ;
      RECT 0.0000 30.4965 9.6120 31.5900 ;
      RECT 0.0000 31.5765 9.6120 32.6700 ;
      RECT 0.0000 32.6565 9.6120 33.7500 ;
      RECT 0.0000 33.7365 9.6120 34.8300 ;
      RECT 0.0000 34.8165 9.6120 35.9100 ;
      RECT 0.0000 35.8965 9.6120 36.9900 ;
      RECT 0.0000 36.9765 9.6120 38.0700 ;
      RECT 0.0000 38.0565 9.6120 39.1500 ;
      RECT 0.0000 39.1365 9.6120 40.2300 ;
      RECT 0.0000 40.2165 9.6120 41.3100 ;
      RECT 0.0000 41.2965 9.6120 42.3900 ;
      RECT 0.0000 42.3765 9.6120 43.4700 ;
      RECT 0.0000 43.4430 9.6120 52.0965 ;
        RECT 0.0000 51.5835 9.6120 52.6770 ;
        RECT 0.0000 52.6635 9.6120 53.7570 ;
        RECT 0.0000 53.7435 9.6120 54.8370 ;
        RECT 0.0000 54.8235 9.6120 55.9170 ;
        RECT 0.0000 55.9035 9.6120 56.9970 ;
        RECT 0.0000 56.9835 9.6120 58.0770 ;
        RECT 0.0000 58.0635 9.6120 59.1570 ;
        RECT 0.0000 59.1435 9.6120 60.2370 ;
        RECT 0.0000 60.2235 9.6120 61.3170 ;
        RECT 0.0000 61.3035 9.6120 62.3970 ;
        RECT 0.0000 62.3835 9.6120 63.4770 ;
        RECT 0.0000 63.4635 9.6120 64.5570 ;
        RECT 0.0000 64.5435 9.6120 65.6370 ;
        RECT 0.0000 65.6235 9.6120 66.7170 ;
        RECT 0.0000 66.7035 9.6120 67.7970 ;
        RECT 0.0000 67.7835 9.6120 68.8770 ;
        RECT 0.0000 68.8635 9.6120 69.9570 ;
        RECT 0.0000 69.9435 9.6120 71.0370 ;
        RECT 0.0000 71.0235 9.6120 72.1170 ;
        RECT 0.0000 72.1035 9.6120 73.1970 ;
        RECT 0.0000 73.1835 9.6120 74.2770 ;
        RECT 0.0000 74.2635 9.6120 75.3570 ;
        RECT 0.0000 75.3435 9.6120 76.4370 ;
        RECT 0.0000 76.4235 9.6120 77.5170 ;
        RECT 0.0000 77.5035 9.6120 78.5970 ;
        RECT 0.0000 78.5835 9.6120 79.6770 ;
        RECT 0.0000 79.6635 9.6120 80.7570 ;
        RECT 0.0000 80.7435 9.6120 81.8370 ;
        RECT 0.0000 81.8235 9.6120 82.9170 ;
        RECT 0.0000 82.9035 9.6120 83.9970 ;
        RECT 0.0000 83.9835 9.6120 85.0770 ;
        RECT 0.0000 85.0635 9.6120 86.1570 ;
        RECT 0.0000 86.1435 9.6120 87.2370 ;
        RECT 0.0000 87.2235 9.6120 88.3170 ;
        RECT 0.0000 88.3035 9.6120 89.3970 ;
        RECT 0.0000 89.3835 9.6120 90.4770 ;
        RECT 0.0000 90.4635 9.6120 91.5570 ;
        RECT 0.0000 91.5435 9.6120 92.6370 ;
        RECT 0.0000 92.6235 9.6120 93.7170 ;
        RECT 0.0000 93.7035 9.6120 94.7970 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5365 9.6120 18.6300 ;
      RECT 0.0000 18.6165 9.6120 19.7100 ;
      RECT 0.0000 19.6965 9.6120 20.7900 ;
      RECT 0.0000 20.7765 9.6120 21.8700 ;
      RECT 0.0000 21.8565 9.6120 22.9500 ;
      RECT 0.0000 22.9365 9.6120 24.0300 ;
      RECT 0.0000 24.0165 9.6120 25.1100 ;
      RECT 0.0000 25.0965 9.6120 26.1900 ;
      RECT 0.0000 26.1765 9.6120 27.2700 ;
      RECT 0.0000 27.2565 9.6120 28.3500 ;
      RECT 0.0000 28.3365 9.6120 29.4300 ;
      RECT 0.0000 29.4165 9.6120 30.5100 ;
      RECT 0.0000 30.4965 9.6120 31.5900 ;
      RECT 0.0000 31.5765 9.6120 32.6700 ;
      RECT 0.0000 32.6565 9.6120 33.7500 ;
      RECT 0.0000 33.7365 9.6120 34.8300 ;
      RECT 0.0000 34.8165 9.6120 35.9100 ;
      RECT 0.0000 35.8965 9.6120 36.9900 ;
      RECT 0.0000 36.9765 9.6120 38.0700 ;
      RECT 0.0000 38.0565 9.6120 39.1500 ;
      RECT 0.0000 39.1365 9.6120 40.2300 ;
      RECT 0.0000 40.2165 9.6120 41.3100 ;
      RECT 0.0000 41.2965 9.6120 42.3900 ;
      RECT 0.0000 42.3765 9.6120 43.4700 ;
      RECT 0.0000 43.4430 9.6120 52.0965 ;
        RECT 0.0000 51.5835 9.6120 52.6770 ;
        RECT 0.0000 52.6635 9.6120 53.7570 ;
        RECT 0.0000 53.7435 9.6120 54.8370 ;
        RECT 0.0000 54.8235 9.6120 55.9170 ;
        RECT 0.0000 55.9035 9.6120 56.9970 ;
        RECT 0.0000 56.9835 9.6120 58.0770 ;
        RECT 0.0000 58.0635 9.6120 59.1570 ;
        RECT 0.0000 59.1435 9.6120 60.2370 ;
        RECT 0.0000 60.2235 9.6120 61.3170 ;
        RECT 0.0000 61.3035 9.6120 62.3970 ;
        RECT 0.0000 62.3835 9.6120 63.4770 ;
        RECT 0.0000 63.4635 9.6120 64.5570 ;
        RECT 0.0000 64.5435 9.6120 65.6370 ;
        RECT 0.0000 65.6235 9.6120 66.7170 ;
        RECT 0.0000 66.7035 9.6120 67.7970 ;
        RECT 0.0000 67.7835 9.6120 68.8770 ;
        RECT 0.0000 68.8635 9.6120 69.9570 ;
        RECT 0.0000 69.9435 9.6120 71.0370 ;
        RECT 0.0000 71.0235 9.6120 72.1170 ;
        RECT 0.0000 72.1035 9.6120 73.1970 ;
        RECT 0.0000 73.1835 9.6120 74.2770 ;
        RECT 0.0000 74.2635 9.6120 75.3570 ;
        RECT 0.0000 75.3435 9.6120 76.4370 ;
        RECT 0.0000 76.4235 9.6120 77.5170 ;
        RECT 0.0000 77.5035 9.6120 78.5970 ;
        RECT 0.0000 78.5835 9.6120 79.6770 ;
        RECT 0.0000 79.6635 9.6120 80.7570 ;
        RECT 0.0000 80.7435 9.6120 81.8370 ;
        RECT 0.0000 81.8235 9.6120 82.9170 ;
        RECT 0.0000 82.9035 9.6120 83.9970 ;
        RECT 0.0000 83.9835 9.6120 85.0770 ;
        RECT 0.0000 85.0635 9.6120 86.1570 ;
        RECT 0.0000 86.1435 9.6120 87.2370 ;
        RECT 0.0000 87.2235 9.6120 88.3170 ;
        RECT 0.0000 88.3035 9.6120 89.3970 ;
        RECT 0.0000 89.3835 9.6120 90.4770 ;
        RECT 0.0000 90.4635 9.6120 91.5570 ;
        RECT 0.0000 91.5435 9.6120 92.6370 ;
        RECT 0.0000 92.6235 9.6120 93.7170 ;
        RECT 0.0000 93.7035 9.6120 94.7970 ;
  LAYER V1  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5365 9.6120 18.6300 ;
      RECT 0.0000 18.6165 9.6120 19.7100 ;
      RECT 0.0000 19.6965 9.6120 20.7900 ;
      RECT 0.0000 20.7765 9.6120 21.8700 ;
      RECT 0.0000 21.8565 9.6120 22.9500 ;
      RECT 0.0000 22.9365 9.6120 24.0300 ;
      RECT 0.0000 24.0165 9.6120 25.1100 ;
      RECT 0.0000 25.0965 9.6120 26.1900 ;
      RECT 0.0000 26.1765 9.6120 27.2700 ;
      RECT 0.0000 27.2565 9.6120 28.3500 ;
      RECT 0.0000 28.3365 9.6120 29.4300 ;
      RECT 0.0000 29.4165 9.6120 30.5100 ;
      RECT 0.0000 30.4965 9.6120 31.5900 ;
      RECT 0.0000 31.5765 9.6120 32.6700 ;
      RECT 0.0000 32.6565 9.6120 33.7500 ;
      RECT 0.0000 33.7365 9.6120 34.8300 ;
      RECT 0.0000 34.8165 9.6120 35.9100 ;
      RECT 0.0000 35.8965 9.6120 36.9900 ;
      RECT 0.0000 36.9765 9.6120 38.0700 ;
      RECT 0.0000 38.0565 9.6120 39.1500 ;
      RECT 0.0000 39.1365 9.6120 40.2300 ;
      RECT 0.0000 40.2165 9.6120 41.3100 ;
      RECT 0.0000 41.2965 9.6120 42.3900 ;
      RECT 0.0000 42.3765 9.6120 43.4700 ;
      RECT 0.0000 43.4430 9.6120 52.0965 ;
        RECT 0.0000 51.5835 9.6120 52.6770 ;
        RECT 0.0000 52.6635 9.6120 53.7570 ;
        RECT 0.0000 53.7435 9.6120 54.8370 ;
        RECT 0.0000 54.8235 9.6120 55.9170 ;
        RECT 0.0000 55.9035 9.6120 56.9970 ;
        RECT 0.0000 56.9835 9.6120 58.0770 ;
        RECT 0.0000 58.0635 9.6120 59.1570 ;
        RECT 0.0000 59.1435 9.6120 60.2370 ;
        RECT 0.0000 60.2235 9.6120 61.3170 ;
        RECT 0.0000 61.3035 9.6120 62.3970 ;
        RECT 0.0000 62.3835 9.6120 63.4770 ;
        RECT 0.0000 63.4635 9.6120 64.5570 ;
        RECT 0.0000 64.5435 9.6120 65.6370 ;
        RECT 0.0000 65.6235 9.6120 66.7170 ;
        RECT 0.0000 66.7035 9.6120 67.7970 ;
        RECT 0.0000 67.7835 9.6120 68.8770 ;
        RECT 0.0000 68.8635 9.6120 69.9570 ;
        RECT 0.0000 69.9435 9.6120 71.0370 ;
        RECT 0.0000 71.0235 9.6120 72.1170 ;
        RECT 0.0000 72.1035 9.6120 73.1970 ;
        RECT 0.0000 73.1835 9.6120 74.2770 ;
        RECT 0.0000 74.2635 9.6120 75.3570 ;
        RECT 0.0000 75.3435 9.6120 76.4370 ;
        RECT 0.0000 76.4235 9.6120 77.5170 ;
        RECT 0.0000 77.5035 9.6120 78.5970 ;
        RECT 0.0000 78.5835 9.6120 79.6770 ;
        RECT 0.0000 79.6635 9.6120 80.7570 ;
        RECT 0.0000 80.7435 9.6120 81.8370 ;
        RECT 0.0000 81.8235 9.6120 82.9170 ;
        RECT 0.0000 82.9035 9.6120 83.9970 ;
        RECT 0.0000 83.9835 9.6120 85.0770 ;
        RECT 0.0000 85.0635 9.6120 86.1570 ;
        RECT 0.0000 86.1435 9.6120 87.2370 ;
        RECT 0.0000 87.2235 9.6120 88.3170 ;
        RECT 0.0000 88.3035 9.6120 89.3970 ;
        RECT 0.0000 89.3835 9.6120 90.4770 ;
        RECT 0.0000 90.4635 9.6120 91.5570 ;
        RECT 0.0000 91.5435 9.6120 92.6370 ;
        RECT 0.0000 92.6235 9.6120 93.7170 ;
        RECT 0.0000 93.7035 9.6120 94.7970 ;
  LAYER V2  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8965 9.6120 9.9900 ;
      RECT 0.0000 9.9765 9.6120 11.0700 ;
      RECT 0.0000 11.0565 9.6120 12.1500 ;
      RECT 0.0000 12.1365 9.6120 13.2300 ;
      RECT 0.0000 13.2165 9.6120 14.3100 ;
      RECT 0.0000 14.2965 9.6120 15.3900 ;
      RECT 0.0000 15.3765 9.6120 16.4700 ;
      RECT 0.0000 16.4565 9.6120 17.5500 ;
      RECT 0.0000 17.5365 9.6120 18.6300 ;
      RECT 0.0000 18.6165 9.6120 19.7100 ;
      RECT 0.0000 19.6965 9.6120 20.7900 ;
      RECT 0.0000 20.7765 9.6120 21.8700 ;
      RECT 0.0000 21.8565 9.6120 22.9500 ;
      RECT 0.0000 22.9365 9.6120 24.0300 ;
      RECT 0.0000 24.0165 9.6120 25.1100 ;
      RECT 0.0000 25.0965 9.6120 26.1900 ;
      RECT 0.0000 26.1765 9.6120 27.2700 ;
      RECT 0.0000 27.2565 9.6120 28.3500 ;
      RECT 0.0000 28.3365 9.6120 29.4300 ;
      RECT 0.0000 29.4165 9.6120 30.5100 ;
      RECT 0.0000 30.4965 9.6120 31.5900 ;
      RECT 0.0000 31.5765 9.6120 32.6700 ;
      RECT 0.0000 32.6565 9.6120 33.7500 ;
      RECT 0.0000 33.7365 9.6120 34.8300 ;
      RECT 0.0000 34.8165 9.6120 35.9100 ;
      RECT 0.0000 35.8965 9.6120 36.9900 ;
      RECT 0.0000 36.9765 9.6120 38.0700 ;
      RECT 0.0000 38.0565 9.6120 39.1500 ;
      RECT 0.0000 39.1365 9.6120 40.2300 ;
      RECT 0.0000 40.2165 9.6120 41.3100 ;
      RECT 0.0000 41.2965 9.6120 42.3900 ;
      RECT 0.0000 42.3765 9.6120 43.4700 ;
      RECT 0.0000 43.4430 9.6120 52.0965 ;
        RECT 0.0000 51.5835 9.6120 52.6770 ;
        RECT 0.0000 52.6635 9.6120 53.7570 ;
        RECT 0.0000 53.7435 9.6120 54.8370 ;
        RECT 0.0000 54.8235 9.6120 55.9170 ;
        RECT 0.0000 55.9035 9.6120 56.9970 ;
        RECT 0.0000 56.9835 9.6120 58.0770 ;
        RECT 0.0000 58.0635 9.6120 59.1570 ;
        RECT 0.0000 59.1435 9.6120 60.2370 ;
        RECT 0.0000 60.2235 9.6120 61.3170 ;
        RECT 0.0000 61.3035 9.6120 62.3970 ;
        RECT 0.0000 62.3835 9.6120 63.4770 ;
        RECT 0.0000 63.4635 9.6120 64.5570 ;
        RECT 0.0000 64.5435 9.6120 65.6370 ;
        RECT 0.0000 65.6235 9.6120 66.7170 ;
        RECT 0.0000 66.7035 9.6120 67.7970 ;
        RECT 0.0000 67.7835 9.6120 68.8770 ;
        RECT 0.0000 68.8635 9.6120 69.9570 ;
        RECT 0.0000 69.9435 9.6120 71.0370 ;
        RECT 0.0000 71.0235 9.6120 72.1170 ;
        RECT 0.0000 72.1035 9.6120 73.1970 ;
        RECT 0.0000 73.1835 9.6120 74.2770 ;
        RECT 0.0000 74.2635 9.6120 75.3570 ;
        RECT 0.0000 75.3435 9.6120 76.4370 ;
        RECT 0.0000 76.4235 9.6120 77.5170 ;
        RECT 0.0000 77.5035 9.6120 78.5970 ;
        RECT 0.0000 78.5835 9.6120 79.6770 ;
        RECT 0.0000 79.6635 9.6120 80.7570 ;
        RECT 0.0000 80.7435 9.6120 81.8370 ;
        RECT 0.0000 81.8235 9.6120 82.9170 ;
        RECT 0.0000 82.9035 9.6120 83.9970 ;
        RECT 0.0000 83.9835 9.6120 85.0770 ;
        RECT 0.0000 85.0635 9.6120 86.1570 ;
        RECT 0.0000 86.1435 9.6120 87.2370 ;
        RECT 0.0000 87.2235 9.6120 88.3170 ;
        RECT 0.0000 88.3035 9.6120 89.3970 ;
        RECT 0.0000 89.3835 9.6120 90.4770 ;
        RECT 0.0000 90.4635 9.6120 91.5570 ;
        RECT 0.0000 91.5435 9.6120 92.6370 ;
        RECT 0.0000 92.6235 9.6120 93.7170 ;
        RECT 0.0000 93.7035 9.6120 94.7970 ;
  LAYER M3  ;
      RECT 5.2380 0.3450 5.2560 1.2805 ;
      RECT 5.2020 0.3450 5.2200 1.2805 ;
      RECT 5.1660 0.9220 5.1840 1.2445 ;
      RECT 5.0490 1.1190 5.0670 1.2285 ;
      RECT 5.0400 0.3775 5.0580 0.6170 ;
      RECT 5.0040 0.9585 5.0220 1.1120 ;
      RECT 4.9230 0.9840 4.9410 1.2420 ;
      RECT 4.3830 0.3450 4.4010 1.2805 ;
      RECT 4.3470 0.3450 4.3650 1.2805 ;
      RECT 4.3110 0.5260 4.3290 1.0940 ;
      RECT 5.2380 1.4250 5.2560 2.3605 ;
      RECT 5.2020 1.4250 5.2200 2.3605 ;
      RECT 5.1660 2.0020 5.1840 2.3245 ;
      RECT 5.0490 2.1990 5.0670 2.3085 ;
      RECT 5.0400 1.4575 5.0580 1.6970 ;
      RECT 5.0040 2.0385 5.0220 2.1920 ;
      RECT 4.9230 2.0640 4.9410 2.3220 ;
      RECT 4.3830 1.4250 4.4010 2.3605 ;
      RECT 4.3470 1.4250 4.3650 2.3605 ;
      RECT 4.3110 1.6060 4.3290 2.1740 ;
      RECT 5.2380 2.5050 5.2560 3.4405 ;
      RECT 5.2020 2.5050 5.2200 3.4405 ;
      RECT 5.1660 3.0820 5.1840 3.4045 ;
      RECT 5.0490 3.2790 5.0670 3.3885 ;
      RECT 5.0400 2.5375 5.0580 2.7770 ;
      RECT 5.0040 3.1185 5.0220 3.2720 ;
      RECT 4.9230 3.1440 4.9410 3.4020 ;
      RECT 4.3830 2.5050 4.4010 3.4405 ;
      RECT 4.3470 2.5050 4.3650 3.4405 ;
      RECT 4.3110 2.6860 4.3290 3.2540 ;
      RECT 5.2380 3.5850 5.2560 4.5205 ;
      RECT 5.2020 3.5850 5.2200 4.5205 ;
      RECT 5.1660 4.1620 5.1840 4.4845 ;
      RECT 5.0490 4.3590 5.0670 4.4685 ;
      RECT 5.0400 3.6175 5.0580 3.8570 ;
      RECT 5.0040 4.1985 5.0220 4.3520 ;
      RECT 4.9230 4.2240 4.9410 4.4820 ;
      RECT 4.3830 3.5850 4.4010 4.5205 ;
      RECT 4.3470 3.5850 4.3650 4.5205 ;
      RECT 4.3110 3.7660 4.3290 4.3340 ;
      RECT 5.2380 4.6650 5.2560 5.6005 ;
      RECT 5.2020 4.6650 5.2200 5.6005 ;
      RECT 5.1660 5.2420 5.1840 5.5645 ;
      RECT 5.0490 5.4390 5.0670 5.5485 ;
      RECT 5.0400 4.6975 5.0580 4.9370 ;
      RECT 5.0040 5.2785 5.0220 5.4320 ;
      RECT 4.9230 5.3040 4.9410 5.5620 ;
      RECT 4.3830 4.6650 4.4010 5.6005 ;
      RECT 4.3470 4.6650 4.3650 5.6005 ;
      RECT 4.3110 4.8460 4.3290 5.4140 ;
      RECT 5.2380 5.7450 5.2560 6.6805 ;
      RECT 5.2020 5.7450 5.2200 6.6805 ;
      RECT 5.1660 6.3220 5.1840 6.6445 ;
      RECT 5.0490 6.5190 5.0670 6.6285 ;
      RECT 5.0400 5.7775 5.0580 6.0170 ;
      RECT 5.0040 6.3585 5.0220 6.5120 ;
      RECT 4.9230 6.3840 4.9410 6.6420 ;
      RECT 4.3830 5.7450 4.4010 6.6805 ;
      RECT 4.3470 5.7450 4.3650 6.6805 ;
      RECT 4.3110 5.9260 4.3290 6.4940 ;
      RECT 5.2380 6.8250 5.2560 7.7605 ;
      RECT 5.2020 6.8250 5.2200 7.7605 ;
      RECT 5.1660 7.4020 5.1840 7.7245 ;
      RECT 5.0490 7.5990 5.0670 7.7085 ;
      RECT 5.0400 6.8575 5.0580 7.0970 ;
      RECT 5.0040 7.4385 5.0220 7.5920 ;
      RECT 4.9230 7.4640 4.9410 7.7220 ;
      RECT 4.3830 6.8250 4.4010 7.7605 ;
      RECT 4.3470 6.8250 4.3650 7.7605 ;
      RECT 4.3110 7.0060 4.3290 7.5740 ;
      RECT 5.2380 7.9050 5.2560 8.8405 ;
      RECT 5.2020 7.9050 5.2200 8.8405 ;
      RECT 5.1660 8.4820 5.1840 8.8045 ;
      RECT 5.0490 8.6790 5.0670 8.7885 ;
      RECT 5.0400 7.9375 5.0580 8.1770 ;
      RECT 5.0040 8.5185 5.0220 8.6720 ;
      RECT 4.9230 8.5440 4.9410 8.8020 ;
      RECT 4.3830 7.9050 4.4010 8.8405 ;
      RECT 4.3470 7.9050 4.3650 8.8405 ;
      RECT 4.3110 8.0860 4.3290 8.6540 ;
      RECT 5.2380 8.9850 5.2560 9.9205 ;
      RECT 5.2020 8.9850 5.2200 9.9205 ;
      RECT 5.1660 9.5620 5.1840 9.8845 ;
      RECT 5.0490 9.7590 5.0670 9.8685 ;
      RECT 5.0400 9.0175 5.0580 9.2570 ;
      RECT 5.0040 9.5985 5.0220 9.7520 ;
      RECT 4.9230 9.6240 4.9410 9.8820 ;
      RECT 4.3830 8.9850 4.4010 9.9205 ;
      RECT 4.3470 8.9850 4.3650 9.9205 ;
      RECT 4.3110 9.1660 4.3290 9.7340 ;
      RECT 5.2380 10.0650 5.2560 11.0005 ;
      RECT 5.2020 10.0650 5.2200 11.0005 ;
      RECT 5.1660 10.6420 5.1840 10.9645 ;
      RECT 5.0490 10.8390 5.0670 10.9485 ;
      RECT 5.0400 10.0975 5.0580 10.3370 ;
      RECT 5.0040 10.6785 5.0220 10.8320 ;
      RECT 4.9230 10.7040 4.9410 10.9620 ;
      RECT 4.3830 10.0650 4.4010 11.0005 ;
      RECT 4.3470 10.0650 4.3650 11.0005 ;
      RECT 4.3110 10.2460 4.3290 10.8140 ;
      RECT 5.2380 11.1450 5.2560 12.0805 ;
      RECT 5.2020 11.1450 5.2200 12.0805 ;
      RECT 5.1660 11.7220 5.1840 12.0445 ;
      RECT 5.0490 11.9190 5.0670 12.0285 ;
      RECT 5.0400 11.1775 5.0580 11.4170 ;
      RECT 5.0040 11.7585 5.0220 11.9120 ;
      RECT 4.9230 11.7840 4.9410 12.0420 ;
      RECT 4.3830 11.1450 4.4010 12.0805 ;
      RECT 4.3470 11.1450 4.3650 12.0805 ;
      RECT 4.3110 11.3260 4.3290 11.8940 ;
      RECT 5.2380 12.2250 5.2560 13.1605 ;
      RECT 5.2020 12.2250 5.2200 13.1605 ;
      RECT 5.1660 12.8020 5.1840 13.1245 ;
      RECT 5.0490 12.9990 5.0670 13.1085 ;
      RECT 5.0400 12.2575 5.0580 12.4970 ;
      RECT 5.0040 12.8385 5.0220 12.9920 ;
      RECT 4.9230 12.8640 4.9410 13.1220 ;
      RECT 4.3830 12.2250 4.4010 13.1605 ;
      RECT 4.3470 12.2250 4.3650 13.1605 ;
      RECT 4.3110 12.4060 4.3290 12.9740 ;
      RECT 5.2380 13.3050 5.2560 14.2405 ;
      RECT 5.2020 13.3050 5.2200 14.2405 ;
      RECT 5.1660 13.8820 5.1840 14.2045 ;
      RECT 5.0490 14.0790 5.0670 14.1885 ;
      RECT 5.0400 13.3375 5.0580 13.5770 ;
      RECT 5.0040 13.9185 5.0220 14.0720 ;
      RECT 4.9230 13.9440 4.9410 14.2020 ;
      RECT 4.3830 13.3050 4.4010 14.2405 ;
      RECT 4.3470 13.3050 4.3650 14.2405 ;
      RECT 4.3110 13.4860 4.3290 14.0540 ;
      RECT 5.2380 14.3850 5.2560 15.3205 ;
      RECT 5.2020 14.3850 5.2200 15.3205 ;
      RECT 5.1660 14.9620 5.1840 15.2845 ;
      RECT 5.0490 15.1590 5.0670 15.2685 ;
      RECT 5.0400 14.4175 5.0580 14.6570 ;
      RECT 5.0040 14.9985 5.0220 15.1520 ;
      RECT 4.9230 15.0240 4.9410 15.2820 ;
      RECT 4.3830 14.3850 4.4010 15.3205 ;
      RECT 4.3470 14.3850 4.3650 15.3205 ;
      RECT 4.3110 14.5660 4.3290 15.1340 ;
      RECT 5.2380 15.4650 5.2560 16.4005 ;
      RECT 5.2020 15.4650 5.2200 16.4005 ;
      RECT 5.1660 16.0420 5.1840 16.3645 ;
      RECT 5.0490 16.2390 5.0670 16.3485 ;
      RECT 5.0400 15.4975 5.0580 15.7370 ;
      RECT 5.0040 16.0785 5.0220 16.2320 ;
      RECT 4.9230 16.1040 4.9410 16.3620 ;
      RECT 4.3830 15.4650 4.4010 16.4005 ;
      RECT 4.3470 15.4650 4.3650 16.4005 ;
      RECT 4.3110 15.6460 4.3290 16.2140 ;
      RECT 5.2380 16.5450 5.2560 17.4805 ;
      RECT 5.2020 16.5450 5.2200 17.4805 ;
      RECT 5.1660 17.1220 5.1840 17.4445 ;
      RECT 5.0490 17.3190 5.0670 17.4285 ;
      RECT 5.0400 16.5775 5.0580 16.8170 ;
      RECT 5.0040 17.1585 5.0220 17.3120 ;
      RECT 4.9230 17.1840 4.9410 17.4420 ;
      RECT 4.3830 16.5450 4.4010 17.4805 ;
      RECT 4.3470 16.5450 4.3650 17.4805 ;
      RECT 4.3110 16.7260 4.3290 17.2940 ;
      RECT 5.2380 17.6250 5.2560 18.5605 ;
      RECT 5.2020 17.6250 5.2200 18.5605 ;
      RECT 5.1660 18.2020 5.1840 18.5245 ;
      RECT 5.0490 18.3990 5.0670 18.5085 ;
      RECT 5.0400 17.6575 5.0580 17.8970 ;
      RECT 5.0040 18.2385 5.0220 18.3920 ;
      RECT 4.9230 18.2640 4.9410 18.5220 ;
      RECT 4.3830 17.6250 4.4010 18.5605 ;
      RECT 4.3470 17.6250 4.3650 18.5605 ;
      RECT 4.3110 17.8060 4.3290 18.3740 ;
      RECT 5.2380 18.7050 5.2560 19.6405 ;
      RECT 5.2020 18.7050 5.2200 19.6405 ;
      RECT 5.1660 19.2820 5.1840 19.6045 ;
      RECT 5.0490 19.4790 5.0670 19.5885 ;
      RECT 5.0400 18.7375 5.0580 18.9770 ;
      RECT 5.0040 19.3185 5.0220 19.4720 ;
      RECT 4.9230 19.3440 4.9410 19.6020 ;
      RECT 4.3830 18.7050 4.4010 19.6405 ;
      RECT 4.3470 18.7050 4.3650 19.6405 ;
      RECT 4.3110 18.8860 4.3290 19.4540 ;
      RECT 5.2380 19.7850 5.2560 20.7205 ;
      RECT 5.2020 19.7850 5.2200 20.7205 ;
      RECT 5.1660 20.3620 5.1840 20.6845 ;
      RECT 5.0490 20.5590 5.0670 20.6685 ;
      RECT 5.0400 19.8175 5.0580 20.0570 ;
      RECT 5.0040 20.3985 5.0220 20.5520 ;
      RECT 4.9230 20.4240 4.9410 20.6820 ;
      RECT 4.3830 19.7850 4.4010 20.7205 ;
      RECT 4.3470 19.7850 4.3650 20.7205 ;
      RECT 4.3110 19.9660 4.3290 20.5340 ;
      RECT 5.2380 20.8650 5.2560 21.8005 ;
      RECT 5.2020 20.8650 5.2200 21.8005 ;
      RECT 5.1660 21.4420 5.1840 21.7645 ;
      RECT 5.0490 21.6390 5.0670 21.7485 ;
      RECT 5.0400 20.8975 5.0580 21.1370 ;
      RECT 5.0040 21.4785 5.0220 21.6320 ;
      RECT 4.9230 21.5040 4.9410 21.7620 ;
      RECT 4.3830 20.8650 4.4010 21.8005 ;
      RECT 4.3470 20.8650 4.3650 21.8005 ;
      RECT 4.3110 21.0460 4.3290 21.6140 ;
      RECT 5.2380 21.9450 5.2560 22.8805 ;
      RECT 5.2020 21.9450 5.2200 22.8805 ;
      RECT 5.1660 22.5220 5.1840 22.8445 ;
      RECT 5.0490 22.7190 5.0670 22.8285 ;
      RECT 5.0400 21.9775 5.0580 22.2170 ;
      RECT 5.0040 22.5585 5.0220 22.7120 ;
      RECT 4.9230 22.5840 4.9410 22.8420 ;
      RECT 4.3830 21.9450 4.4010 22.8805 ;
      RECT 4.3470 21.9450 4.3650 22.8805 ;
      RECT 4.3110 22.1260 4.3290 22.6940 ;
      RECT 5.2380 23.0250 5.2560 23.9605 ;
      RECT 5.2020 23.0250 5.2200 23.9605 ;
      RECT 5.1660 23.6020 5.1840 23.9245 ;
      RECT 5.0490 23.7990 5.0670 23.9085 ;
      RECT 5.0400 23.0575 5.0580 23.2970 ;
      RECT 5.0040 23.6385 5.0220 23.7920 ;
      RECT 4.9230 23.6640 4.9410 23.9220 ;
      RECT 4.3830 23.0250 4.4010 23.9605 ;
      RECT 4.3470 23.0250 4.3650 23.9605 ;
      RECT 4.3110 23.2060 4.3290 23.7740 ;
      RECT 5.2380 24.1050 5.2560 25.0405 ;
      RECT 5.2020 24.1050 5.2200 25.0405 ;
      RECT 5.1660 24.6820 5.1840 25.0045 ;
      RECT 5.0490 24.8790 5.0670 24.9885 ;
      RECT 5.0400 24.1375 5.0580 24.3770 ;
      RECT 5.0040 24.7185 5.0220 24.8720 ;
      RECT 4.9230 24.7440 4.9410 25.0020 ;
      RECT 4.3830 24.1050 4.4010 25.0405 ;
      RECT 4.3470 24.1050 4.3650 25.0405 ;
      RECT 4.3110 24.2860 4.3290 24.8540 ;
      RECT 5.2380 25.1850 5.2560 26.1205 ;
      RECT 5.2020 25.1850 5.2200 26.1205 ;
      RECT 5.1660 25.7620 5.1840 26.0845 ;
      RECT 5.0490 25.9590 5.0670 26.0685 ;
      RECT 5.0400 25.2175 5.0580 25.4570 ;
      RECT 5.0040 25.7985 5.0220 25.9520 ;
      RECT 4.9230 25.8240 4.9410 26.0820 ;
      RECT 4.3830 25.1850 4.4010 26.1205 ;
      RECT 4.3470 25.1850 4.3650 26.1205 ;
      RECT 4.3110 25.3660 4.3290 25.9340 ;
      RECT 5.2380 26.2650 5.2560 27.2005 ;
      RECT 5.2020 26.2650 5.2200 27.2005 ;
      RECT 5.1660 26.8420 5.1840 27.1645 ;
      RECT 5.0490 27.0390 5.0670 27.1485 ;
      RECT 5.0400 26.2975 5.0580 26.5370 ;
      RECT 5.0040 26.8785 5.0220 27.0320 ;
      RECT 4.9230 26.9040 4.9410 27.1620 ;
      RECT 4.3830 26.2650 4.4010 27.2005 ;
      RECT 4.3470 26.2650 4.3650 27.2005 ;
      RECT 4.3110 26.4460 4.3290 27.0140 ;
      RECT 5.2380 27.3450 5.2560 28.2805 ;
      RECT 5.2020 27.3450 5.2200 28.2805 ;
      RECT 5.1660 27.9220 5.1840 28.2445 ;
      RECT 5.0490 28.1190 5.0670 28.2285 ;
      RECT 5.0400 27.3775 5.0580 27.6170 ;
      RECT 5.0040 27.9585 5.0220 28.1120 ;
      RECT 4.9230 27.9840 4.9410 28.2420 ;
      RECT 4.3830 27.3450 4.4010 28.2805 ;
      RECT 4.3470 27.3450 4.3650 28.2805 ;
      RECT 4.3110 27.5260 4.3290 28.0940 ;
      RECT 5.2380 28.4250 5.2560 29.3605 ;
      RECT 5.2020 28.4250 5.2200 29.3605 ;
      RECT 5.1660 29.0020 5.1840 29.3245 ;
      RECT 5.0490 29.1990 5.0670 29.3085 ;
      RECT 5.0400 28.4575 5.0580 28.6970 ;
      RECT 5.0040 29.0385 5.0220 29.1920 ;
      RECT 4.9230 29.0640 4.9410 29.3220 ;
      RECT 4.3830 28.4250 4.4010 29.3605 ;
      RECT 4.3470 28.4250 4.3650 29.3605 ;
      RECT 4.3110 28.6060 4.3290 29.1740 ;
      RECT 5.2380 29.5050 5.2560 30.4405 ;
      RECT 5.2020 29.5050 5.2200 30.4405 ;
      RECT 5.1660 30.0820 5.1840 30.4045 ;
      RECT 5.0490 30.2790 5.0670 30.3885 ;
      RECT 5.0400 29.5375 5.0580 29.7770 ;
      RECT 5.0040 30.1185 5.0220 30.2720 ;
      RECT 4.9230 30.1440 4.9410 30.4020 ;
      RECT 4.3830 29.5050 4.4010 30.4405 ;
      RECT 4.3470 29.5050 4.3650 30.4405 ;
      RECT 4.3110 29.6860 4.3290 30.2540 ;
      RECT 5.2380 30.5850 5.2560 31.5205 ;
      RECT 5.2020 30.5850 5.2200 31.5205 ;
      RECT 5.1660 31.1620 5.1840 31.4845 ;
      RECT 5.0490 31.3590 5.0670 31.4685 ;
      RECT 5.0400 30.6175 5.0580 30.8570 ;
      RECT 5.0040 31.1985 5.0220 31.3520 ;
      RECT 4.9230 31.2240 4.9410 31.4820 ;
      RECT 4.3830 30.5850 4.4010 31.5205 ;
      RECT 4.3470 30.5850 4.3650 31.5205 ;
      RECT 4.3110 30.7660 4.3290 31.3340 ;
      RECT 5.2380 31.6650 5.2560 32.6005 ;
      RECT 5.2020 31.6650 5.2200 32.6005 ;
      RECT 5.1660 32.2420 5.1840 32.5645 ;
      RECT 5.0490 32.4390 5.0670 32.5485 ;
      RECT 5.0400 31.6975 5.0580 31.9370 ;
      RECT 5.0040 32.2785 5.0220 32.4320 ;
      RECT 4.9230 32.3040 4.9410 32.5620 ;
      RECT 4.3830 31.6650 4.4010 32.6005 ;
      RECT 4.3470 31.6650 4.3650 32.6005 ;
      RECT 4.3110 31.8460 4.3290 32.4140 ;
      RECT 5.2380 32.7450 5.2560 33.6805 ;
      RECT 5.2020 32.7450 5.2200 33.6805 ;
      RECT 5.1660 33.3220 5.1840 33.6445 ;
      RECT 5.0490 33.5190 5.0670 33.6285 ;
      RECT 5.0400 32.7775 5.0580 33.0170 ;
      RECT 5.0040 33.3585 5.0220 33.5120 ;
      RECT 4.9230 33.3840 4.9410 33.6420 ;
      RECT 4.3830 32.7450 4.4010 33.6805 ;
      RECT 4.3470 32.7450 4.3650 33.6805 ;
      RECT 4.3110 32.9260 4.3290 33.4940 ;
      RECT 5.2380 33.8250 5.2560 34.7605 ;
      RECT 5.2020 33.8250 5.2200 34.7605 ;
      RECT 5.1660 34.4020 5.1840 34.7245 ;
      RECT 5.0490 34.5990 5.0670 34.7085 ;
      RECT 5.0400 33.8575 5.0580 34.0970 ;
      RECT 5.0040 34.4385 5.0220 34.5920 ;
      RECT 4.9230 34.4640 4.9410 34.7220 ;
      RECT 4.3830 33.8250 4.4010 34.7605 ;
      RECT 4.3470 33.8250 4.3650 34.7605 ;
      RECT 4.3110 34.0060 4.3290 34.5740 ;
      RECT 5.2380 34.9050 5.2560 35.8405 ;
      RECT 5.2020 34.9050 5.2200 35.8405 ;
      RECT 5.1660 35.4820 5.1840 35.8045 ;
      RECT 5.0490 35.6790 5.0670 35.7885 ;
      RECT 5.0400 34.9375 5.0580 35.1770 ;
      RECT 5.0040 35.5185 5.0220 35.6720 ;
      RECT 4.9230 35.5440 4.9410 35.8020 ;
      RECT 4.3830 34.9050 4.4010 35.8405 ;
      RECT 4.3470 34.9050 4.3650 35.8405 ;
      RECT 4.3110 35.0860 4.3290 35.6540 ;
      RECT 5.2380 35.9850 5.2560 36.9205 ;
      RECT 5.2020 35.9850 5.2200 36.9205 ;
      RECT 5.1660 36.5620 5.1840 36.8845 ;
      RECT 5.0490 36.7590 5.0670 36.8685 ;
      RECT 5.0400 36.0175 5.0580 36.2570 ;
      RECT 5.0040 36.5985 5.0220 36.7520 ;
      RECT 4.9230 36.6240 4.9410 36.8820 ;
      RECT 4.3830 35.9850 4.4010 36.9205 ;
      RECT 4.3470 35.9850 4.3650 36.9205 ;
      RECT 4.3110 36.1660 4.3290 36.7340 ;
      RECT 5.2380 37.0650 5.2560 38.0005 ;
      RECT 5.2020 37.0650 5.2200 38.0005 ;
      RECT 5.1660 37.6420 5.1840 37.9645 ;
      RECT 5.0490 37.8390 5.0670 37.9485 ;
      RECT 5.0400 37.0975 5.0580 37.3370 ;
      RECT 5.0040 37.6785 5.0220 37.8320 ;
      RECT 4.9230 37.7040 4.9410 37.9620 ;
      RECT 4.3830 37.0650 4.4010 38.0005 ;
      RECT 4.3470 37.0650 4.3650 38.0005 ;
      RECT 4.3110 37.2460 4.3290 37.8140 ;
      RECT 5.2380 38.1450 5.2560 39.0805 ;
      RECT 5.2020 38.1450 5.2200 39.0805 ;
      RECT 5.1660 38.7220 5.1840 39.0445 ;
      RECT 5.0490 38.9190 5.0670 39.0285 ;
      RECT 5.0400 38.1775 5.0580 38.4170 ;
      RECT 5.0040 38.7585 5.0220 38.9120 ;
      RECT 4.9230 38.7840 4.9410 39.0420 ;
      RECT 4.3830 38.1450 4.4010 39.0805 ;
      RECT 4.3470 38.1450 4.3650 39.0805 ;
      RECT 4.3110 38.3260 4.3290 38.8940 ;
      RECT 5.2380 39.2250 5.2560 40.1605 ;
      RECT 5.2020 39.2250 5.2200 40.1605 ;
      RECT 5.1660 39.8020 5.1840 40.1245 ;
      RECT 5.0490 39.9990 5.0670 40.1085 ;
      RECT 5.0400 39.2575 5.0580 39.4970 ;
      RECT 5.0040 39.8385 5.0220 39.9920 ;
      RECT 4.9230 39.8640 4.9410 40.1220 ;
      RECT 4.3830 39.2250 4.4010 40.1605 ;
      RECT 4.3470 39.2250 4.3650 40.1605 ;
      RECT 4.3110 39.4060 4.3290 39.9740 ;
      RECT 5.2380 40.3050 5.2560 41.2405 ;
      RECT 5.2020 40.3050 5.2200 41.2405 ;
      RECT 5.1660 40.8820 5.1840 41.2045 ;
      RECT 5.0490 41.0790 5.0670 41.1885 ;
      RECT 5.0400 40.3375 5.0580 40.5770 ;
      RECT 5.0040 40.9185 5.0220 41.0720 ;
      RECT 4.9230 40.9440 4.9410 41.2020 ;
      RECT 4.3830 40.3050 4.4010 41.2405 ;
      RECT 4.3470 40.3050 4.3650 41.2405 ;
      RECT 4.3110 40.4860 4.3290 41.0540 ;
      RECT 5.2380 41.3850 5.2560 42.3205 ;
      RECT 5.2020 41.3850 5.2200 42.3205 ;
      RECT 5.1660 41.9620 5.1840 42.2845 ;
      RECT 5.0490 42.1590 5.0670 42.2685 ;
      RECT 5.0400 41.4175 5.0580 41.6570 ;
      RECT 5.0040 41.9985 5.0220 42.1520 ;
      RECT 4.9230 42.0240 4.9410 42.2820 ;
      RECT 4.3830 41.3850 4.4010 42.3205 ;
      RECT 4.3470 41.3850 4.3650 42.3205 ;
      RECT 4.3110 41.5660 4.3290 42.1340 ;
      RECT 5.2380 42.4650 5.2560 43.4005 ;
      RECT 5.2020 42.4650 5.2200 43.4005 ;
      RECT 5.1660 43.0420 5.1840 43.3645 ;
      RECT 5.0490 43.2390 5.0670 43.3485 ;
      RECT 5.0400 42.4975 5.0580 42.7370 ;
      RECT 5.0040 43.0785 5.0220 43.2320 ;
      RECT 4.9230 43.1040 4.9410 43.3620 ;
      RECT 4.3830 42.4650 4.4010 43.4005 ;
      RECT 4.3470 42.4650 4.3650 43.4005 ;
      RECT 4.3110 42.6460 4.3290 43.2140 ;
      RECT 9.4050 47.2360 9.4230 51.5915 ;
      RECT 9.3690 45.9210 9.3870 45.9900 ;
      RECT 9.3690 47.7290 9.3870 48.1935 ;
      RECT 9.3330 43.4165 9.3510 51.6235 ;
      RECT 9.2970 47.1860 9.3150 47.9585 ;
      RECT 9.2970 48.0097 9.3150 48.5010 ;
      RECT 9.2970 48.5510 9.3150 48.9225 ;
      RECT 9.2970 48.9855 9.3150 49.7970 ;
      RECT 9.2610 47.2715 9.2790 47.9135 ;
      RECT 9.2610 48.5910 9.2790 49.1230 ;
      RECT 9.2250 43.4165 9.2430 43.7665 ;
      RECT 9.1170 43.4165 9.1350 43.7665 ;
      RECT 9.0090 43.4165 9.0270 43.7665 ;
      RECT 8.9010 43.4165 8.9190 43.7665 ;
      RECT 8.7930 43.4165 8.8110 43.7665 ;
      RECT 8.6850 43.4165 8.7030 43.7665 ;
      RECT 8.5770 43.4165 8.5950 43.7665 ;
      RECT 8.4690 43.4165 8.4870 43.7665 ;
      RECT 8.3610 43.4165 8.3790 43.7665 ;
      RECT 8.2530 43.4165 8.2710 43.7665 ;
      RECT 8.1450 43.4165 8.1630 43.7665 ;
      RECT 8.0370 43.4165 8.0550 43.7665 ;
      RECT 7.9290 43.4165 7.9470 43.7665 ;
      RECT 7.8210 43.4165 7.8390 43.7665 ;
      RECT 7.7130 43.4165 7.7310 43.7665 ;
      RECT 7.6050 43.4165 7.6230 43.7665 ;
      RECT 7.4970 43.4165 7.5150 43.7665 ;
      RECT 7.3890 43.4165 7.4070 43.7665 ;
      RECT 7.2810 43.4165 7.2990 43.7665 ;
      RECT 7.1730 43.4165 7.1910 43.7665 ;
      RECT 7.0650 43.4165 7.0830 43.7665 ;
      RECT 6.9570 43.4165 6.9750 43.7665 ;
      RECT 6.8490 43.4165 6.8670 43.7665 ;
      RECT 6.7410 43.4165 6.7590 43.7665 ;
      RECT 6.6330 43.4165 6.6510 43.7665 ;
      RECT 6.5250 43.4165 6.5430 43.7665 ;
      RECT 6.4170 43.4165 6.4350 43.7665 ;
      RECT 6.3090 43.4165 6.3270 43.7665 ;
      RECT 6.2010 43.4165 6.2190 43.7665 ;
      RECT 6.0930 43.4165 6.1110 43.7665 ;
      RECT 6.0570 47.2050 6.0750 47.9097 ;
      RECT 6.0570 48.6520 6.0750 49.8330 ;
      RECT 6.0390 44.0770 6.0570 44.7530 ;
      RECT 6.0390 45.4990 6.0570 45.7970 ;
      RECT 6.0210 47.2685 6.0390 47.9585 ;
      RECT 6.0210 48.0095 6.0390 49.0010 ;
      RECT 6.0210 49.0310 6.0390 49.8150 ;
      RECT 5.9850 43.4165 6.0030 51.6235 ;
      RECT 5.9490 47.5410 5.9670 47.6240 ;
      RECT 5.9310 44.1850 5.9490 44.8160 ;
      RECT 5.9310 45.2290 5.9490 45.4190 ;
      RECT 5.9310 46.1110 5.9490 46.1600 ;
      RECT 5.9130 47.2360 5.9310 51.5960 ;
      RECT 5.8230 43.8070 5.8410 44.6090 ;
      RECT 5.8230 45.1570 5.8410 45.7250 ;
      RECT 5.7870 45.2290 5.8050 45.5990 ;
      RECT 5.7510 44.5810 5.7690 44.7170 ;
      RECT 5.7510 45.5710 5.7690 45.7970 ;
      RECT 5.7510 46.8130 5.7690 46.8770 ;
      RECT 5.7150 44.6830 5.7330 44.7200 ;
      RECT 5.7150 46.3090 5.7330 46.3520 ;
      RECT 5.7150 46.8430 5.7330 46.8800 ;
      RECT 5.6790 44.9950 5.6970 45.4910 ;
      RECT 5.6790 45.5350 5.6970 45.7250 ;
      RECT 5.6790 46.4950 5.6970 46.8050 ;
      RECT 5.6430 48.7750 5.6610 49.5050 ;
      RECT 5.6430 49.8550 5.6610 50.5850 ;
      RECT 5.3190 44.6170 5.3370 44.9150 ;
      RECT 5.3190 45.8050 5.3370 45.8690 ;
      RECT 5.3190 46.0750 5.3370 46.5350 ;
      RECT 5.3190 47.2750 5.3370 47.3120 ;
      RECT 5.3190 49.3150 5.3370 49.6130 ;
      RECT 5.2830 44.6890 5.3010 45.1940 ;
      RECT 5.2830 45.4630 5.3010 46.2650 ;
      RECT 5.2830 47.3080 5.3010 47.5790 ;
      RECT 5.2830 47.6590 5.3010 47.8850 ;
      RECT 5.2470 44.6170 5.2650 45.2930 ;
      RECT 5.2470 45.3910 5.2650 45.7250 ;
      RECT 5.2470 45.9310 5.2650 46.0670 ;
      RECT 5.2470 46.6150 5.2650 47.4170 ;
      RECT 5.2470 47.8510 5.2650 47.8880 ;
      RECT 5.2470 50.0170 5.2650 50.3510 ;
      RECT 5.2110 44.8510 5.2290 44.9870 ;
      RECT 5.2110 46.7410 5.2290 47.7230 ;
      RECT 5.2110 48.1630 5.2290 48.4610 ;
      RECT 5.2110 49.8550 5.2290 50.1170 ;
      RECT 5.1750 43.9150 5.1930 44.0690 ;
      RECT 5.1750 44.7250 5.1930 46.5110 ;
      RECT 5.1750 47.5510 5.1930 49.8830 ;
      RECT 5.1750 50.0890 5.1930 51.1970 ;
      RECT 4.8870 44.1850 4.9050 44.4470 ;
      RECT 4.8870 44.5810 4.9050 44.6450 ;
      RECT 4.8870 44.7250 4.9050 44.9510 ;
      RECT 4.8870 44.9950 4.9050 45.1850 ;
      RECT 4.8870 45.2650 4.9050 47.8850 ;
      RECT 4.8870 47.9290 4.9050 49.2350 ;
      RECT 4.8870 50.3230 4.9050 50.5850 ;
      RECT 4.8510 45.1840 4.8690 45.4550 ;
      RECT 4.8510 45.5350 4.8690 46.3730 ;
      RECT 4.8510 46.5430 4.8690 47.3810 ;
      RECT 4.8510 47.4250 4.8690 48.6950 ;
      RECT 4.8510 48.9010 4.8690 49.0730 ;
      RECT 4.8510 49.7830 4.8690 50.8550 ;
      RECT 4.8150 45.2650 4.8330 45.5360 ;
      RECT 4.8150 45.6910 4.8330 45.7280 ;
      RECT 4.8150 46.4710 4.8330 47.4530 ;
      RECT 4.8150 47.6950 4.8330 48.1550 ;
      RECT 4.8150 48.5050 4.8330 49.2440 ;
      RECT 4.7790 44.3830 4.7970 45.4550 ;
      RECT 4.7790 47.0470 4.7970 47.2640 ;
      RECT 4.7790 48.4330 4.7970 48.7310 ;
      RECT 4.7430 45.0310 4.7610 45.4910 ;
      RECT 4.7430 46.6150 4.7610 46.8050 ;
      RECT 4.7430 46.8460 4.7610 46.8830 ;
      RECT 4.7430 47.1190 4.7610 47.4530 ;
      RECT 4.7430 47.5870 4.7610 48.9290 ;
      RECT 4.7430 49.0360 4.7610 50.1530 ;
      RECT 4.7070 44.4550 4.7250 44.6450 ;
      RECT 4.7070 44.8510 4.7250 44.9870 ;
      RECT 4.7070 45.2650 4.7250 48.4250 ;
      RECT 4.7070 48.5050 4.7250 48.9650 ;
      RECT 4.7070 49.5850 4.7250 50.0450 ;
      RECT 4.7070 50.8990 4.7250 51.1250 ;
      RECT 4.6710 43.4430 4.6890 43.5970 ;
      RECT 4.6710 51.4540 4.6890 51.6080 ;
      RECT 4.6350 43.4430 4.6530 43.4930 ;
      RECT 4.5630 43.4430 4.5810 43.5145 ;
      RECT 4.5630 51.5235 4.5810 51.6235 ;
      RECT 4.4190 44.9590 4.4370 45.1490 ;
      RECT 4.4190 45.6970 4.4370 46.0670 ;
      RECT 4.4190 47.6590 4.4370 47.8850 ;
      RECT 4.4190 48.1990 4.4370 49.3430 ;
      RECT 4.4190 50.1250 4.4370 50.5850 ;
      RECT 4.4190 51.1630 4.4370 51.2000 ;
      RECT 4.3830 43.9150 4.4010 44.4110 ;
      RECT 4.3830 47.9950 4.4010 48.0320 ;
      RECT 4.3830 49.0720 4.4010 49.8830 ;
      RECT 4.3470 44.3830 4.3650 44.6450 ;
      RECT 4.3470 44.9230 4.3650 45.2570 ;
      RECT 4.3470 45.4630 4.3650 45.5630 ;
      RECT 4.3470 46.3450 4.3650 49.1090 ;
      RECT 4.3470 49.2430 4.3650 49.4690 ;
      RECT 4.3110 44.0410 4.3290 45.1850 ;
      RECT 4.3110 48.7750 4.3290 48.9650 ;
      RECT 4.3110 49.5790 4.3290 49.6160 ;
      RECT 4.3110 49.8550 4.3290 50.6570 ;
      RECT 4.2750 44.9950 4.2930 45.9950 ;
      RECT 4.2750 49.4350 4.2930 49.4720 ;
      RECT 4.2390 44.1850 4.2570 44.2130 ;
      RECT 3.9150 44.5810 3.9330 44.9870 ;
      RECT 3.8430 44.6170 3.8610 45.2210 ;
      RECT 3.8070 44.4550 3.8250 44.5190 ;
      RECT 3.7710 43.4960 3.7890 43.5470 ;
      RECT 3.7710 46.6150 3.7890 46.8050 ;
      RECT 3.7710 47.2360 3.7890 51.5960 ;
      RECT 3.6810 47.2360 3.6990 51.5960 ;
      RECT 3.6630 43.9150 3.6810 44.1050 ;
      RECT 3.6630 44.6890 3.6810 46.9490 ;
      RECT 3.6450 47.5410 3.6630 47.6240 ;
      RECT 3.6090 43.4165 3.6270 51.6235 ;
      RECT 3.5730 47.2685 3.5910 47.9585 ;
      RECT 3.5730 48.0095 3.5910 49.0010 ;
      RECT 3.5730 49.0310 3.5910 49.8150 ;
      RECT 3.5550 43.9150 3.5730 44.4110 ;
      RECT 3.5550 45.1930 3.5730 45.7610 ;
      RECT 3.5550 46.0750 3.5730 46.8050 ;
      RECT 3.5370 47.2050 3.5550 47.9097 ;
      RECT 3.5370 48.6520 3.5550 49.8330 ;
      RECT 3.5010 43.4165 3.5190 43.7665 ;
      RECT 3.3930 43.4165 3.4110 43.7665 ;
      RECT 3.2850 43.4165 3.3030 43.7665 ;
      RECT 3.1770 43.4165 3.1950 43.7665 ;
      RECT 3.0690 43.4165 3.0870 43.7665 ;
      RECT 2.9610 43.4165 2.9790 43.7665 ;
      RECT 2.8530 43.4165 2.8710 43.7665 ;
      RECT 2.7450 43.4165 2.7630 43.7665 ;
      RECT 2.6370 43.4165 2.6550 43.7665 ;
      RECT 2.5290 43.4165 2.5470 43.7665 ;
      RECT 2.4210 43.4165 2.4390 43.7665 ;
      RECT 2.3130 43.4165 2.3310 43.7665 ;
      RECT 2.2050 43.4165 2.2230 43.7665 ;
      RECT 2.0970 43.4165 2.1150 43.7665 ;
      RECT 1.9890 43.4165 2.0070 43.7665 ;
      RECT 1.8810 43.4165 1.8990 43.7665 ;
      RECT 1.7730 43.4165 1.7910 43.7665 ;
      RECT 1.6650 43.4165 1.6830 43.7665 ;
      RECT 1.5570 43.4165 1.5750 43.7665 ;
      RECT 1.4490 43.4165 1.4670 43.7665 ;
      RECT 1.3410 43.4165 1.3590 43.7665 ;
      RECT 1.2330 43.4165 1.2510 43.7665 ;
      RECT 1.1250 43.4165 1.1430 43.7665 ;
      RECT 1.0170 43.4165 1.0350 43.7665 ;
      RECT 0.9090 43.4165 0.9270 43.7665 ;
      RECT 0.8010 43.4165 0.8190 43.7665 ;
      RECT 0.6930 43.4165 0.7110 43.7665 ;
      RECT 0.5850 43.4165 0.6030 43.7665 ;
      RECT 0.4770 43.4165 0.4950 43.7665 ;
      RECT 0.3690 43.4165 0.3870 43.7665 ;
      RECT 0.3330 47.2715 0.3510 47.9135 ;
      RECT 0.3330 48.5910 0.3510 49.1230 ;
      RECT 0.3150 44.4550 0.3330 44.6810 ;
      RECT 0.2970 47.1860 0.3150 47.9585 ;
      RECT 0.2970 48.0097 0.3150 48.5010 ;
      RECT 0.2970 48.5510 0.3150 48.9225 ;
      RECT 0.2970 48.9855 0.3150 49.7970 ;
      RECT 0.2610 43.4165 0.2790 51.6235 ;
      RECT 0.2250 45.9210 0.2430 45.9900 ;
      RECT 0.2250 47.7290 0.2430 48.1935 ;
      RECT 0.1890 47.2360 0.2070 51.5915 ;
        RECT 5.2380 51.6720 5.2560 52.6075 ;
        RECT 5.2020 51.6720 5.2200 52.6075 ;
        RECT 5.1660 52.2490 5.1840 52.5715 ;
        RECT 5.0490 52.4460 5.0670 52.5555 ;
        RECT 5.0400 51.7045 5.0580 51.9440 ;
        RECT 5.0040 52.2855 5.0220 52.4390 ;
        RECT 4.9230 52.3110 4.9410 52.5690 ;
        RECT 4.3830 51.6720 4.4010 52.6075 ;
        RECT 4.3470 51.6720 4.3650 52.6075 ;
        RECT 4.3110 51.8530 4.3290 52.4210 ;
        RECT 5.2380 52.7520 5.2560 53.6875 ;
        RECT 5.2020 52.7520 5.2200 53.6875 ;
        RECT 5.1660 53.3290 5.1840 53.6515 ;
        RECT 5.0490 53.5260 5.0670 53.6355 ;
        RECT 5.0400 52.7845 5.0580 53.0240 ;
        RECT 5.0040 53.3655 5.0220 53.5190 ;
        RECT 4.9230 53.3910 4.9410 53.6490 ;
        RECT 4.3830 52.7520 4.4010 53.6875 ;
        RECT 4.3470 52.7520 4.3650 53.6875 ;
        RECT 4.3110 52.9330 4.3290 53.5010 ;
        RECT 5.2380 53.8320 5.2560 54.7675 ;
        RECT 5.2020 53.8320 5.2200 54.7675 ;
        RECT 5.1660 54.4090 5.1840 54.7315 ;
        RECT 5.0490 54.6060 5.0670 54.7155 ;
        RECT 5.0400 53.8645 5.0580 54.1040 ;
        RECT 5.0040 54.4455 5.0220 54.5990 ;
        RECT 4.9230 54.4710 4.9410 54.7290 ;
        RECT 4.3830 53.8320 4.4010 54.7675 ;
        RECT 4.3470 53.8320 4.3650 54.7675 ;
        RECT 4.3110 54.0130 4.3290 54.5810 ;
        RECT 5.2380 54.9120 5.2560 55.8475 ;
        RECT 5.2020 54.9120 5.2200 55.8475 ;
        RECT 5.1660 55.4890 5.1840 55.8115 ;
        RECT 5.0490 55.6860 5.0670 55.7955 ;
        RECT 5.0400 54.9445 5.0580 55.1840 ;
        RECT 5.0040 55.5255 5.0220 55.6790 ;
        RECT 4.9230 55.5510 4.9410 55.8090 ;
        RECT 4.3830 54.9120 4.4010 55.8475 ;
        RECT 4.3470 54.9120 4.3650 55.8475 ;
        RECT 4.3110 55.0930 4.3290 55.6610 ;
        RECT 5.2380 55.9920 5.2560 56.9275 ;
        RECT 5.2020 55.9920 5.2200 56.9275 ;
        RECT 5.1660 56.5690 5.1840 56.8915 ;
        RECT 5.0490 56.7660 5.0670 56.8755 ;
        RECT 5.0400 56.0245 5.0580 56.2640 ;
        RECT 5.0040 56.6055 5.0220 56.7590 ;
        RECT 4.9230 56.6310 4.9410 56.8890 ;
        RECT 4.3830 55.9920 4.4010 56.9275 ;
        RECT 4.3470 55.9920 4.3650 56.9275 ;
        RECT 4.3110 56.1730 4.3290 56.7410 ;
        RECT 5.2380 57.0720 5.2560 58.0075 ;
        RECT 5.2020 57.0720 5.2200 58.0075 ;
        RECT 5.1660 57.6490 5.1840 57.9715 ;
        RECT 5.0490 57.8460 5.0670 57.9555 ;
        RECT 5.0400 57.1045 5.0580 57.3440 ;
        RECT 5.0040 57.6855 5.0220 57.8390 ;
        RECT 4.9230 57.7110 4.9410 57.9690 ;
        RECT 4.3830 57.0720 4.4010 58.0075 ;
        RECT 4.3470 57.0720 4.3650 58.0075 ;
        RECT 4.3110 57.2530 4.3290 57.8210 ;
        RECT 5.2380 58.1520 5.2560 59.0875 ;
        RECT 5.2020 58.1520 5.2200 59.0875 ;
        RECT 5.1660 58.7290 5.1840 59.0515 ;
        RECT 5.0490 58.9260 5.0670 59.0355 ;
        RECT 5.0400 58.1845 5.0580 58.4240 ;
        RECT 5.0040 58.7655 5.0220 58.9190 ;
        RECT 4.9230 58.7910 4.9410 59.0490 ;
        RECT 4.3830 58.1520 4.4010 59.0875 ;
        RECT 4.3470 58.1520 4.3650 59.0875 ;
        RECT 4.3110 58.3330 4.3290 58.9010 ;
        RECT 5.2380 59.2320 5.2560 60.1675 ;
        RECT 5.2020 59.2320 5.2200 60.1675 ;
        RECT 5.1660 59.8090 5.1840 60.1315 ;
        RECT 5.0490 60.0060 5.0670 60.1155 ;
        RECT 5.0400 59.2645 5.0580 59.5040 ;
        RECT 5.0040 59.8455 5.0220 59.9990 ;
        RECT 4.9230 59.8710 4.9410 60.1290 ;
        RECT 4.3830 59.2320 4.4010 60.1675 ;
        RECT 4.3470 59.2320 4.3650 60.1675 ;
        RECT 4.3110 59.4130 4.3290 59.9810 ;
        RECT 5.2380 60.3120 5.2560 61.2475 ;
        RECT 5.2020 60.3120 5.2200 61.2475 ;
        RECT 5.1660 60.8890 5.1840 61.2115 ;
        RECT 5.0490 61.0860 5.0670 61.1955 ;
        RECT 5.0400 60.3445 5.0580 60.5840 ;
        RECT 5.0040 60.9255 5.0220 61.0790 ;
        RECT 4.9230 60.9510 4.9410 61.2090 ;
        RECT 4.3830 60.3120 4.4010 61.2475 ;
        RECT 4.3470 60.3120 4.3650 61.2475 ;
        RECT 4.3110 60.4930 4.3290 61.0610 ;
        RECT 5.2380 61.3920 5.2560 62.3275 ;
        RECT 5.2020 61.3920 5.2200 62.3275 ;
        RECT 5.1660 61.9690 5.1840 62.2915 ;
        RECT 5.0490 62.1660 5.0670 62.2755 ;
        RECT 5.0400 61.4245 5.0580 61.6640 ;
        RECT 5.0040 62.0055 5.0220 62.1590 ;
        RECT 4.9230 62.0310 4.9410 62.2890 ;
        RECT 4.3830 61.3920 4.4010 62.3275 ;
        RECT 4.3470 61.3920 4.3650 62.3275 ;
        RECT 4.3110 61.5730 4.3290 62.1410 ;
        RECT 5.2380 62.4720 5.2560 63.4075 ;
        RECT 5.2020 62.4720 5.2200 63.4075 ;
        RECT 5.1660 63.0490 5.1840 63.3715 ;
        RECT 5.0490 63.2460 5.0670 63.3555 ;
        RECT 5.0400 62.5045 5.0580 62.7440 ;
        RECT 5.0040 63.0855 5.0220 63.2390 ;
        RECT 4.9230 63.1110 4.9410 63.3690 ;
        RECT 4.3830 62.4720 4.4010 63.4075 ;
        RECT 4.3470 62.4720 4.3650 63.4075 ;
        RECT 4.3110 62.6530 4.3290 63.2210 ;
        RECT 5.2380 63.5520 5.2560 64.4875 ;
        RECT 5.2020 63.5520 5.2200 64.4875 ;
        RECT 5.1660 64.1290 5.1840 64.4515 ;
        RECT 5.0490 64.3260 5.0670 64.4355 ;
        RECT 5.0400 63.5845 5.0580 63.8240 ;
        RECT 5.0040 64.1655 5.0220 64.3190 ;
        RECT 4.9230 64.1910 4.9410 64.4490 ;
        RECT 4.3830 63.5520 4.4010 64.4875 ;
        RECT 4.3470 63.5520 4.3650 64.4875 ;
        RECT 4.3110 63.7330 4.3290 64.3010 ;
        RECT 5.2380 64.6320 5.2560 65.5675 ;
        RECT 5.2020 64.6320 5.2200 65.5675 ;
        RECT 5.1660 65.2090 5.1840 65.5315 ;
        RECT 5.0490 65.4060 5.0670 65.5155 ;
        RECT 5.0400 64.6645 5.0580 64.9040 ;
        RECT 5.0040 65.2455 5.0220 65.3990 ;
        RECT 4.9230 65.2710 4.9410 65.5290 ;
        RECT 4.3830 64.6320 4.4010 65.5675 ;
        RECT 4.3470 64.6320 4.3650 65.5675 ;
        RECT 4.3110 64.8130 4.3290 65.3810 ;
        RECT 5.2380 65.7120 5.2560 66.6475 ;
        RECT 5.2020 65.7120 5.2200 66.6475 ;
        RECT 5.1660 66.2890 5.1840 66.6115 ;
        RECT 5.0490 66.4860 5.0670 66.5955 ;
        RECT 5.0400 65.7445 5.0580 65.9840 ;
        RECT 5.0040 66.3255 5.0220 66.4790 ;
        RECT 4.9230 66.3510 4.9410 66.6090 ;
        RECT 4.3830 65.7120 4.4010 66.6475 ;
        RECT 4.3470 65.7120 4.3650 66.6475 ;
        RECT 4.3110 65.8930 4.3290 66.4610 ;
        RECT 5.2380 66.7920 5.2560 67.7275 ;
        RECT 5.2020 66.7920 5.2200 67.7275 ;
        RECT 5.1660 67.3690 5.1840 67.6915 ;
        RECT 5.0490 67.5660 5.0670 67.6755 ;
        RECT 5.0400 66.8245 5.0580 67.0640 ;
        RECT 5.0040 67.4055 5.0220 67.5590 ;
        RECT 4.9230 67.4310 4.9410 67.6890 ;
        RECT 4.3830 66.7920 4.4010 67.7275 ;
        RECT 4.3470 66.7920 4.3650 67.7275 ;
        RECT 4.3110 66.9730 4.3290 67.5410 ;
        RECT 5.2380 67.8720 5.2560 68.8075 ;
        RECT 5.2020 67.8720 5.2200 68.8075 ;
        RECT 5.1660 68.4490 5.1840 68.7715 ;
        RECT 5.0490 68.6460 5.0670 68.7555 ;
        RECT 5.0400 67.9045 5.0580 68.1440 ;
        RECT 5.0040 68.4855 5.0220 68.6390 ;
        RECT 4.9230 68.5110 4.9410 68.7690 ;
        RECT 4.3830 67.8720 4.4010 68.8075 ;
        RECT 4.3470 67.8720 4.3650 68.8075 ;
        RECT 4.3110 68.0530 4.3290 68.6210 ;
        RECT 5.2380 68.9520 5.2560 69.8875 ;
        RECT 5.2020 68.9520 5.2200 69.8875 ;
        RECT 5.1660 69.5290 5.1840 69.8515 ;
        RECT 5.0490 69.7260 5.0670 69.8355 ;
        RECT 5.0400 68.9845 5.0580 69.2240 ;
        RECT 5.0040 69.5655 5.0220 69.7190 ;
        RECT 4.9230 69.5910 4.9410 69.8490 ;
        RECT 4.3830 68.9520 4.4010 69.8875 ;
        RECT 4.3470 68.9520 4.3650 69.8875 ;
        RECT 4.3110 69.1330 4.3290 69.7010 ;
        RECT 5.2380 70.0320 5.2560 70.9675 ;
        RECT 5.2020 70.0320 5.2200 70.9675 ;
        RECT 5.1660 70.6090 5.1840 70.9315 ;
        RECT 5.0490 70.8060 5.0670 70.9155 ;
        RECT 5.0400 70.0645 5.0580 70.3040 ;
        RECT 5.0040 70.6455 5.0220 70.7990 ;
        RECT 4.9230 70.6710 4.9410 70.9290 ;
        RECT 4.3830 70.0320 4.4010 70.9675 ;
        RECT 4.3470 70.0320 4.3650 70.9675 ;
        RECT 4.3110 70.2130 4.3290 70.7810 ;
        RECT 5.2380 71.1120 5.2560 72.0475 ;
        RECT 5.2020 71.1120 5.2200 72.0475 ;
        RECT 5.1660 71.6890 5.1840 72.0115 ;
        RECT 5.0490 71.8860 5.0670 71.9955 ;
        RECT 5.0400 71.1445 5.0580 71.3840 ;
        RECT 5.0040 71.7255 5.0220 71.8790 ;
        RECT 4.9230 71.7510 4.9410 72.0090 ;
        RECT 4.3830 71.1120 4.4010 72.0475 ;
        RECT 4.3470 71.1120 4.3650 72.0475 ;
        RECT 4.3110 71.2930 4.3290 71.8610 ;
        RECT 5.2380 72.1920 5.2560 73.1275 ;
        RECT 5.2020 72.1920 5.2200 73.1275 ;
        RECT 5.1660 72.7690 5.1840 73.0915 ;
        RECT 5.0490 72.9660 5.0670 73.0755 ;
        RECT 5.0400 72.2245 5.0580 72.4640 ;
        RECT 5.0040 72.8055 5.0220 72.9590 ;
        RECT 4.9230 72.8310 4.9410 73.0890 ;
        RECT 4.3830 72.1920 4.4010 73.1275 ;
        RECT 4.3470 72.1920 4.3650 73.1275 ;
        RECT 4.3110 72.3730 4.3290 72.9410 ;
        RECT 5.2380 73.2720 5.2560 74.2075 ;
        RECT 5.2020 73.2720 5.2200 74.2075 ;
        RECT 5.1660 73.8490 5.1840 74.1715 ;
        RECT 5.0490 74.0460 5.0670 74.1555 ;
        RECT 5.0400 73.3045 5.0580 73.5440 ;
        RECT 5.0040 73.8855 5.0220 74.0390 ;
        RECT 4.9230 73.9110 4.9410 74.1690 ;
        RECT 4.3830 73.2720 4.4010 74.2075 ;
        RECT 4.3470 73.2720 4.3650 74.2075 ;
        RECT 4.3110 73.4530 4.3290 74.0210 ;
        RECT 5.2380 74.3520 5.2560 75.2875 ;
        RECT 5.2020 74.3520 5.2200 75.2875 ;
        RECT 5.1660 74.9290 5.1840 75.2515 ;
        RECT 5.0490 75.1260 5.0670 75.2355 ;
        RECT 5.0400 74.3845 5.0580 74.6240 ;
        RECT 5.0040 74.9655 5.0220 75.1190 ;
        RECT 4.9230 74.9910 4.9410 75.2490 ;
        RECT 4.3830 74.3520 4.4010 75.2875 ;
        RECT 4.3470 74.3520 4.3650 75.2875 ;
        RECT 4.3110 74.5330 4.3290 75.1010 ;
        RECT 5.2380 75.4320 5.2560 76.3675 ;
        RECT 5.2020 75.4320 5.2200 76.3675 ;
        RECT 5.1660 76.0090 5.1840 76.3315 ;
        RECT 5.0490 76.2060 5.0670 76.3155 ;
        RECT 5.0400 75.4645 5.0580 75.7040 ;
        RECT 5.0040 76.0455 5.0220 76.1990 ;
        RECT 4.9230 76.0710 4.9410 76.3290 ;
        RECT 4.3830 75.4320 4.4010 76.3675 ;
        RECT 4.3470 75.4320 4.3650 76.3675 ;
        RECT 4.3110 75.6130 4.3290 76.1810 ;
        RECT 5.2380 76.5120 5.2560 77.4475 ;
        RECT 5.2020 76.5120 5.2200 77.4475 ;
        RECT 5.1660 77.0890 5.1840 77.4115 ;
        RECT 5.0490 77.2860 5.0670 77.3955 ;
        RECT 5.0400 76.5445 5.0580 76.7840 ;
        RECT 5.0040 77.1255 5.0220 77.2790 ;
        RECT 4.9230 77.1510 4.9410 77.4090 ;
        RECT 4.3830 76.5120 4.4010 77.4475 ;
        RECT 4.3470 76.5120 4.3650 77.4475 ;
        RECT 4.3110 76.6930 4.3290 77.2610 ;
        RECT 5.2380 77.5920 5.2560 78.5275 ;
        RECT 5.2020 77.5920 5.2200 78.5275 ;
        RECT 5.1660 78.1690 5.1840 78.4915 ;
        RECT 5.0490 78.3660 5.0670 78.4755 ;
        RECT 5.0400 77.6245 5.0580 77.8640 ;
        RECT 5.0040 78.2055 5.0220 78.3590 ;
        RECT 4.9230 78.2310 4.9410 78.4890 ;
        RECT 4.3830 77.5920 4.4010 78.5275 ;
        RECT 4.3470 77.5920 4.3650 78.5275 ;
        RECT 4.3110 77.7730 4.3290 78.3410 ;
        RECT 5.2380 78.6720 5.2560 79.6075 ;
        RECT 5.2020 78.6720 5.2200 79.6075 ;
        RECT 5.1660 79.2490 5.1840 79.5715 ;
        RECT 5.0490 79.4460 5.0670 79.5555 ;
        RECT 5.0400 78.7045 5.0580 78.9440 ;
        RECT 5.0040 79.2855 5.0220 79.4390 ;
        RECT 4.9230 79.3110 4.9410 79.5690 ;
        RECT 4.3830 78.6720 4.4010 79.6075 ;
        RECT 4.3470 78.6720 4.3650 79.6075 ;
        RECT 4.3110 78.8530 4.3290 79.4210 ;
        RECT 5.2380 79.7520 5.2560 80.6875 ;
        RECT 5.2020 79.7520 5.2200 80.6875 ;
        RECT 5.1660 80.3290 5.1840 80.6515 ;
        RECT 5.0490 80.5260 5.0670 80.6355 ;
        RECT 5.0400 79.7845 5.0580 80.0240 ;
        RECT 5.0040 80.3655 5.0220 80.5190 ;
        RECT 4.9230 80.3910 4.9410 80.6490 ;
        RECT 4.3830 79.7520 4.4010 80.6875 ;
        RECT 4.3470 79.7520 4.3650 80.6875 ;
        RECT 4.3110 79.9330 4.3290 80.5010 ;
        RECT 5.2380 80.8320 5.2560 81.7675 ;
        RECT 5.2020 80.8320 5.2200 81.7675 ;
        RECT 5.1660 81.4090 5.1840 81.7315 ;
        RECT 5.0490 81.6060 5.0670 81.7155 ;
        RECT 5.0400 80.8645 5.0580 81.1040 ;
        RECT 5.0040 81.4455 5.0220 81.5990 ;
        RECT 4.9230 81.4710 4.9410 81.7290 ;
        RECT 4.3830 80.8320 4.4010 81.7675 ;
        RECT 4.3470 80.8320 4.3650 81.7675 ;
        RECT 4.3110 81.0130 4.3290 81.5810 ;
        RECT 5.2380 81.9120 5.2560 82.8475 ;
        RECT 5.2020 81.9120 5.2200 82.8475 ;
        RECT 5.1660 82.4890 5.1840 82.8115 ;
        RECT 5.0490 82.6860 5.0670 82.7955 ;
        RECT 5.0400 81.9445 5.0580 82.1840 ;
        RECT 5.0040 82.5255 5.0220 82.6790 ;
        RECT 4.9230 82.5510 4.9410 82.8090 ;
        RECT 4.3830 81.9120 4.4010 82.8475 ;
        RECT 4.3470 81.9120 4.3650 82.8475 ;
        RECT 4.3110 82.0930 4.3290 82.6610 ;
        RECT 5.2380 82.9920 5.2560 83.9275 ;
        RECT 5.2020 82.9920 5.2200 83.9275 ;
        RECT 5.1660 83.5690 5.1840 83.8915 ;
        RECT 5.0490 83.7660 5.0670 83.8755 ;
        RECT 5.0400 83.0245 5.0580 83.2640 ;
        RECT 5.0040 83.6055 5.0220 83.7590 ;
        RECT 4.9230 83.6310 4.9410 83.8890 ;
        RECT 4.3830 82.9920 4.4010 83.9275 ;
        RECT 4.3470 82.9920 4.3650 83.9275 ;
        RECT 4.3110 83.1730 4.3290 83.7410 ;
        RECT 5.2380 84.0720 5.2560 85.0075 ;
        RECT 5.2020 84.0720 5.2200 85.0075 ;
        RECT 5.1660 84.6490 5.1840 84.9715 ;
        RECT 5.0490 84.8460 5.0670 84.9555 ;
        RECT 5.0400 84.1045 5.0580 84.3440 ;
        RECT 5.0040 84.6855 5.0220 84.8390 ;
        RECT 4.9230 84.7110 4.9410 84.9690 ;
        RECT 4.3830 84.0720 4.4010 85.0075 ;
        RECT 4.3470 84.0720 4.3650 85.0075 ;
        RECT 4.3110 84.2530 4.3290 84.8210 ;
        RECT 5.2380 85.1520 5.2560 86.0875 ;
        RECT 5.2020 85.1520 5.2200 86.0875 ;
        RECT 5.1660 85.7290 5.1840 86.0515 ;
        RECT 5.0490 85.9260 5.0670 86.0355 ;
        RECT 5.0400 85.1845 5.0580 85.4240 ;
        RECT 5.0040 85.7655 5.0220 85.9190 ;
        RECT 4.9230 85.7910 4.9410 86.0490 ;
        RECT 4.3830 85.1520 4.4010 86.0875 ;
        RECT 4.3470 85.1520 4.3650 86.0875 ;
        RECT 4.3110 85.3330 4.3290 85.9010 ;
        RECT 5.2380 86.2320 5.2560 87.1675 ;
        RECT 5.2020 86.2320 5.2200 87.1675 ;
        RECT 5.1660 86.8090 5.1840 87.1315 ;
        RECT 5.0490 87.0060 5.0670 87.1155 ;
        RECT 5.0400 86.2645 5.0580 86.5040 ;
        RECT 5.0040 86.8455 5.0220 86.9990 ;
        RECT 4.9230 86.8710 4.9410 87.1290 ;
        RECT 4.3830 86.2320 4.4010 87.1675 ;
        RECT 4.3470 86.2320 4.3650 87.1675 ;
        RECT 4.3110 86.4130 4.3290 86.9810 ;
        RECT 5.2380 87.3120 5.2560 88.2475 ;
        RECT 5.2020 87.3120 5.2200 88.2475 ;
        RECT 5.1660 87.8890 5.1840 88.2115 ;
        RECT 5.0490 88.0860 5.0670 88.1955 ;
        RECT 5.0400 87.3445 5.0580 87.5840 ;
        RECT 5.0040 87.9255 5.0220 88.0790 ;
        RECT 4.9230 87.9510 4.9410 88.2090 ;
        RECT 4.3830 87.3120 4.4010 88.2475 ;
        RECT 4.3470 87.3120 4.3650 88.2475 ;
        RECT 4.3110 87.4930 4.3290 88.0610 ;
        RECT 5.2380 88.3920 5.2560 89.3275 ;
        RECT 5.2020 88.3920 5.2200 89.3275 ;
        RECT 5.1660 88.9690 5.1840 89.2915 ;
        RECT 5.0490 89.1660 5.0670 89.2755 ;
        RECT 5.0400 88.4245 5.0580 88.6640 ;
        RECT 5.0040 89.0055 5.0220 89.1590 ;
        RECT 4.9230 89.0310 4.9410 89.2890 ;
        RECT 4.3830 88.3920 4.4010 89.3275 ;
        RECT 4.3470 88.3920 4.3650 89.3275 ;
        RECT 4.3110 88.5730 4.3290 89.1410 ;
        RECT 5.2380 89.4720 5.2560 90.4075 ;
        RECT 5.2020 89.4720 5.2200 90.4075 ;
        RECT 5.1660 90.0490 5.1840 90.3715 ;
        RECT 5.0490 90.2460 5.0670 90.3555 ;
        RECT 5.0400 89.5045 5.0580 89.7440 ;
        RECT 5.0040 90.0855 5.0220 90.2390 ;
        RECT 4.9230 90.1110 4.9410 90.3690 ;
        RECT 4.3830 89.4720 4.4010 90.4075 ;
        RECT 4.3470 89.4720 4.3650 90.4075 ;
        RECT 4.3110 89.6530 4.3290 90.2210 ;
        RECT 5.2380 90.5520 5.2560 91.4875 ;
        RECT 5.2020 90.5520 5.2200 91.4875 ;
        RECT 5.1660 91.1290 5.1840 91.4515 ;
        RECT 5.0490 91.3260 5.0670 91.4355 ;
        RECT 5.0400 90.5845 5.0580 90.8240 ;
        RECT 5.0040 91.1655 5.0220 91.3190 ;
        RECT 4.9230 91.1910 4.9410 91.4490 ;
        RECT 4.3830 90.5520 4.4010 91.4875 ;
        RECT 4.3470 90.5520 4.3650 91.4875 ;
        RECT 4.3110 90.7330 4.3290 91.3010 ;
        RECT 5.2380 91.6320 5.2560 92.5675 ;
        RECT 5.2020 91.6320 5.2200 92.5675 ;
        RECT 5.1660 92.2090 5.1840 92.5315 ;
        RECT 5.0490 92.4060 5.0670 92.5155 ;
        RECT 5.0400 91.6645 5.0580 91.9040 ;
        RECT 5.0040 92.2455 5.0220 92.3990 ;
        RECT 4.9230 92.2710 4.9410 92.5290 ;
        RECT 4.3830 91.6320 4.4010 92.5675 ;
        RECT 4.3470 91.6320 4.3650 92.5675 ;
        RECT 4.3110 91.8130 4.3290 92.3810 ;
        RECT 5.2380 92.7120 5.2560 93.6475 ;
        RECT 5.2020 92.7120 5.2200 93.6475 ;
        RECT 5.1660 93.2890 5.1840 93.6115 ;
        RECT 5.0490 93.4860 5.0670 93.5955 ;
        RECT 5.0400 92.7445 5.0580 92.9840 ;
        RECT 5.0040 93.3255 5.0220 93.4790 ;
        RECT 4.9230 93.3510 4.9410 93.6090 ;
        RECT 4.3830 92.7120 4.4010 93.6475 ;
        RECT 4.3470 92.7120 4.3650 93.6475 ;
        RECT 4.3110 92.8930 4.3290 93.4610 ;
        RECT 5.2380 93.7920 5.2560 94.7275 ;
        RECT 5.2020 93.7920 5.2200 94.7275 ;
        RECT 5.1660 94.3690 5.1840 94.6915 ;
        RECT 5.0490 94.5660 5.0670 94.6755 ;
        RECT 5.0400 93.8245 5.0580 94.0640 ;
        RECT 5.0040 94.4055 5.0220 94.5590 ;
        RECT 4.9230 94.4310 4.9410 94.6890 ;
        RECT 4.3830 93.7920 4.4010 94.7275 ;
        RECT 4.3470 93.7920 4.3650 94.7275 ;
        RECT 4.3110 93.9730 4.3290 94.5410 ;
  LAYER M3 SPACING 0.018  ;
      RECT 5.1800 0.2565 5.3080 1.3500 ;
      RECT 5.1660 0.9220 5.3080 1.2445 ;
      RECT 5.0180 0.6490 5.0800 1.3500 ;
      RECT 5.0040 0.9585 5.0800 1.1120 ;
      RECT 5.0180 0.2565 5.0440 1.3500 ;
      RECT 5.0180 0.3775 5.0580 0.6170 ;
      RECT 5.0180 0.2565 5.0800 0.3455 ;
      RECT 4.7210 0.7070 4.9270 1.3500 ;
      RECT 4.9010 0.2565 4.9270 1.3500 ;
      RECT 4.7210 0.9840 4.9410 1.2420 ;
      RECT 4.7210 0.2565 4.8190 1.3500 ;
      RECT 4.3040 0.2565 4.3870 1.3500 ;
      RECT 4.3040 0.3450 4.4010 1.2805 ;
      RECT 9.5270 0.2565 9.6120 1.3500 ;
      RECT 9.3830 0.2565 9.4090 1.3500 ;
      RECT 9.2750 0.2565 9.3010 1.3500 ;
      RECT 9.1670 0.2565 9.1930 1.3500 ;
      RECT 9.0590 0.2565 9.0850 1.3500 ;
      RECT 8.9510 0.2565 8.9770 1.3500 ;
      RECT 8.8430 0.2565 8.8690 1.3500 ;
      RECT 8.7350 0.2565 8.7610 1.3500 ;
      RECT 8.6270 0.2565 8.6530 1.3500 ;
      RECT 8.5190 0.2565 8.5450 1.3500 ;
      RECT 8.4110 0.2565 8.4370 1.3500 ;
      RECT 8.3030 0.2565 8.3290 1.3500 ;
      RECT 8.1950 0.2565 8.2210 1.3500 ;
      RECT 8.0870 0.2565 8.1130 1.3500 ;
      RECT 7.9790 0.2565 8.0050 1.3500 ;
      RECT 7.8710 0.2565 7.8970 1.3500 ;
      RECT 7.7630 0.2565 7.7890 1.3500 ;
      RECT 7.6550 0.2565 7.6810 1.3500 ;
      RECT 7.5470 0.2565 7.5730 1.3500 ;
      RECT 7.4390 0.2565 7.4650 1.3500 ;
      RECT 7.3310 0.2565 7.3570 1.3500 ;
      RECT 7.2230 0.2565 7.2490 1.3500 ;
      RECT 7.1150 0.2565 7.1410 1.3500 ;
      RECT 7.0070 0.2565 7.0330 1.3500 ;
      RECT 6.8990 0.2565 6.9250 1.3500 ;
      RECT 6.7910 0.2565 6.8170 1.3500 ;
      RECT 6.6830 0.2565 6.7090 1.3500 ;
      RECT 6.5750 0.2565 6.6010 1.3500 ;
      RECT 6.4670 0.2565 6.4930 1.3500 ;
      RECT 6.3590 0.2565 6.3850 1.3500 ;
      RECT 6.2510 0.2565 6.2770 1.3500 ;
      RECT 6.1430 0.2565 6.1690 1.3500 ;
      RECT 6.0350 0.2565 6.0610 1.3500 ;
      RECT 5.9270 0.2565 5.9530 1.3500 ;
      RECT 5.7140 0.2565 5.7910 1.3500 ;
      RECT 3.8210 0.2565 3.8980 1.3500 ;
      RECT 3.6590 0.2565 3.6850 1.3500 ;
      RECT 3.5510 0.2565 3.5770 1.3500 ;
      RECT 3.4430 0.2565 3.4690 1.3500 ;
      RECT 3.3350 0.2565 3.3610 1.3500 ;
      RECT 3.2270 0.2565 3.2530 1.3500 ;
      RECT 3.1190 0.2565 3.1450 1.3500 ;
      RECT 3.0110 0.2565 3.0370 1.3500 ;
      RECT 2.9030 0.2565 2.9290 1.3500 ;
      RECT 2.7950 0.2565 2.8210 1.3500 ;
      RECT 2.6870 0.2565 2.7130 1.3500 ;
      RECT 2.5790 0.2565 2.6050 1.3500 ;
      RECT 2.4710 0.2565 2.4970 1.3500 ;
      RECT 2.3630 0.2565 2.3890 1.3500 ;
      RECT 2.2550 0.2565 2.2810 1.3500 ;
      RECT 2.1470 0.2565 2.1730 1.3500 ;
      RECT 2.0390 0.2565 2.0650 1.3500 ;
      RECT 1.9310 0.2565 1.9570 1.3500 ;
      RECT 1.8230 0.2565 1.8490 1.3500 ;
      RECT 1.7150 0.2565 1.7410 1.3500 ;
      RECT 1.6070 0.2565 1.6330 1.3500 ;
      RECT 1.4990 0.2565 1.5250 1.3500 ;
      RECT 1.3910 0.2565 1.4170 1.3500 ;
      RECT 1.2830 0.2565 1.3090 1.3500 ;
      RECT 1.1750 0.2565 1.2010 1.3500 ;
      RECT 1.0670 0.2565 1.0930 1.3500 ;
      RECT 0.9590 0.2565 0.9850 1.3500 ;
      RECT 0.8510 0.2565 0.8770 1.3500 ;
      RECT 0.7430 0.2565 0.7690 1.3500 ;
      RECT 0.6350 0.2565 0.6610 1.3500 ;
      RECT 0.5270 0.2565 0.5530 1.3500 ;
      RECT 0.4190 0.2565 0.4450 1.3500 ;
      RECT 0.3110 0.2565 0.3370 1.3500 ;
      RECT 0.2030 0.2565 0.2290 1.3500 ;
      RECT 0.0000 0.2565 0.0850 1.3500 ;
      RECT 5.1800 1.3365 5.3080 2.4300 ;
      RECT 5.1660 2.0020 5.3080 2.3245 ;
      RECT 5.0180 1.7290 5.0800 2.4300 ;
      RECT 5.0040 2.0385 5.0800 2.1920 ;
      RECT 5.0180 1.3365 5.0440 2.4300 ;
      RECT 5.0180 1.4575 5.0580 1.6970 ;
      RECT 5.0180 1.3365 5.0800 1.4255 ;
      RECT 4.7210 1.7870 4.9270 2.4300 ;
      RECT 4.9010 1.3365 4.9270 2.4300 ;
      RECT 4.7210 2.0640 4.9410 2.3220 ;
      RECT 4.7210 1.3365 4.8190 2.4300 ;
      RECT 4.3040 1.3365 4.3870 2.4300 ;
      RECT 4.3040 1.4250 4.4010 2.3605 ;
      RECT 9.5270 1.3365 9.6120 2.4300 ;
      RECT 9.3830 1.3365 9.4090 2.4300 ;
      RECT 9.2750 1.3365 9.3010 2.4300 ;
      RECT 9.1670 1.3365 9.1930 2.4300 ;
      RECT 9.0590 1.3365 9.0850 2.4300 ;
      RECT 8.9510 1.3365 8.9770 2.4300 ;
      RECT 8.8430 1.3365 8.8690 2.4300 ;
      RECT 8.7350 1.3365 8.7610 2.4300 ;
      RECT 8.6270 1.3365 8.6530 2.4300 ;
      RECT 8.5190 1.3365 8.5450 2.4300 ;
      RECT 8.4110 1.3365 8.4370 2.4300 ;
      RECT 8.3030 1.3365 8.3290 2.4300 ;
      RECT 8.1950 1.3365 8.2210 2.4300 ;
      RECT 8.0870 1.3365 8.1130 2.4300 ;
      RECT 7.9790 1.3365 8.0050 2.4300 ;
      RECT 7.8710 1.3365 7.8970 2.4300 ;
      RECT 7.7630 1.3365 7.7890 2.4300 ;
      RECT 7.6550 1.3365 7.6810 2.4300 ;
      RECT 7.5470 1.3365 7.5730 2.4300 ;
      RECT 7.4390 1.3365 7.4650 2.4300 ;
      RECT 7.3310 1.3365 7.3570 2.4300 ;
      RECT 7.2230 1.3365 7.2490 2.4300 ;
      RECT 7.1150 1.3365 7.1410 2.4300 ;
      RECT 7.0070 1.3365 7.0330 2.4300 ;
      RECT 6.8990 1.3365 6.9250 2.4300 ;
      RECT 6.7910 1.3365 6.8170 2.4300 ;
      RECT 6.6830 1.3365 6.7090 2.4300 ;
      RECT 6.5750 1.3365 6.6010 2.4300 ;
      RECT 6.4670 1.3365 6.4930 2.4300 ;
      RECT 6.3590 1.3365 6.3850 2.4300 ;
      RECT 6.2510 1.3365 6.2770 2.4300 ;
      RECT 6.1430 1.3365 6.1690 2.4300 ;
      RECT 6.0350 1.3365 6.0610 2.4300 ;
      RECT 5.9270 1.3365 5.9530 2.4300 ;
      RECT 5.7140 1.3365 5.7910 2.4300 ;
      RECT 3.8210 1.3365 3.8980 2.4300 ;
      RECT 3.6590 1.3365 3.6850 2.4300 ;
      RECT 3.5510 1.3365 3.5770 2.4300 ;
      RECT 3.4430 1.3365 3.4690 2.4300 ;
      RECT 3.3350 1.3365 3.3610 2.4300 ;
      RECT 3.2270 1.3365 3.2530 2.4300 ;
      RECT 3.1190 1.3365 3.1450 2.4300 ;
      RECT 3.0110 1.3365 3.0370 2.4300 ;
      RECT 2.9030 1.3365 2.9290 2.4300 ;
      RECT 2.7950 1.3365 2.8210 2.4300 ;
      RECT 2.6870 1.3365 2.7130 2.4300 ;
      RECT 2.5790 1.3365 2.6050 2.4300 ;
      RECT 2.4710 1.3365 2.4970 2.4300 ;
      RECT 2.3630 1.3365 2.3890 2.4300 ;
      RECT 2.2550 1.3365 2.2810 2.4300 ;
      RECT 2.1470 1.3365 2.1730 2.4300 ;
      RECT 2.0390 1.3365 2.0650 2.4300 ;
      RECT 1.9310 1.3365 1.9570 2.4300 ;
      RECT 1.8230 1.3365 1.8490 2.4300 ;
      RECT 1.7150 1.3365 1.7410 2.4300 ;
      RECT 1.6070 1.3365 1.6330 2.4300 ;
      RECT 1.4990 1.3365 1.5250 2.4300 ;
      RECT 1.3910 1.3365 1.4170 2.4300 ;
      RECT 1.2830 1.3365 1.3090 2.4300 ;
      RECT 1.1750 1.3365 1.2010 2.4300 ;
      RECT 1.0670 1.3365 1.0930 2.4300 ;
      RECT 0.9590 1.3365 0.9850 2.4300 ;
      RECT 0.8510 1.3365 0.8770 2.4300 ;
      RECT 0.7430 1.3365 0.7690 2.4300 ;
      RECT 0.6350 1.3365 0.6610 2.4300 ;
      RECT 0.5270 1.3365 0.5530 2.4300 ;
      RECT 0.4190 1.3365 0.4450 2.4300 ;
      RECT 0.3110 1.3365 0.3370 2.4300 ;
      RECT 0.2030 1.3365 0.2290 2.4300 ;
      RECT 0.0000 1.3365 0.0850 2.4300 ;
      RECT 5.1800 2.4165 5.3080 3.5100 ;
      RECT 5.1660 3.0820 5.3080 3.4045 ;
      RECT 5.0180 2.8090 5.0800 3.5100 ;
      RECT 5.0040 3.1185 5.0800 3.2720 ;
      RECT 5.0180 2.4165 5.0440 3.5100 ;
      RECT 5.0180 2.5375 5.0580 2.7770 ;
      RECT 5.0180 2.4165 5.0800 2.5055 ;
      RECT 4.7210 2.8670 4.9270 3.5100 ;
      RECT 4.9010 2.4165 4.9270 3.5100 ;
      RECT 4.7210 3.1440 4.9410 3.4020 ;
      RECT 4.7210 2.4165 4.8190 3.5100 ;
      RECT 4.3040 2.4165 4.3870 3.5100 ;
      RECT 4.3040 2.5050 4.4010 3.4405 ;
      RECT 9.5270 2.4165 9.6120 3.5100 ;
      RECT 9.3830 2.4165 9.4090 3.5100 ;
      RECT 9.2750 2.4165 9.3010 3.5100 ;
      RECT 9.1670 2.4165 9.1930 3.5100 ;
      RECT 9.0590 2.4165 9.0850 3.5100 ;
      RECT 8.9510 2.4165 8.9770 3.5100 ;
      RECT 8.8430 2.4165 8.8690 3.5100 ;
      RECT 8.7350 2.4165 8.7610 3.5100 ;
      RECT 8.6270 2.4165 8.6530 3.5100 ;
      RECT 8.5190 2.4165 8.5450 3.5100 ;
      RECT 8.4110 2.4165 8.4370 3.5100 ;
      RECT 8.3030 2.4165 8.3290 3.5100 ;
      RECT 8.1950 2.4165 8.2210 3.5100 ;
      RECT 8.0870 2.4165 8.1130 3.5100 ;
      RECT 7.9790 2.4165 8.0050 3.5100 ;
      RECT 7.8710 2.4165 7.8970 3.5100 ;
      RECT 7.7630 2.4165 7.7890 3.5100 ;
      RECT 7.6550 2.4165 7.6810 3.5100 ;
      RECT 7.5470 2.4165 7.5730 3.5100 ;
      RECT 7.4390 2.4165 7.4650 3.5100 ;
      RECT 7.3310 2.4165 7.3570 3.5100 ;
      RECT 7.2230 2.4165 7.2490 3.5100 ;
      RECT 7.1150 2.4165 7.1410 3.5100 ;
      RECT 7.0070 2.4165 7.0330 3.5100 ;
      RECT 6.8990 2.4165 6.9250 3.5100 ;
      RECT 6.7910 2.4165 6.8170 3.5100 ;
      RECT 6.6830 2.4165 6.7090 3.5100 ;
      RECT 6.5750 2.4165 6.6010 3.5100 ;
      RECT 6.4670 2.4165 6.4930 3.5100 ;
      RECT 6.3590 2.4165 6.3850 3.5100 ;
      RECT 6.2510 2.4165 6.2770 3.5100 ;
      RECT 6.1430 2.4165 6.1690 3.5100 ;
      RECT 6.0350 2.4165 6.0610 3.5100 ;
      RECT 5.9270 2.4165 5.9530 3.5100 ;
      RECT 5.7140 2.4165 5.7910 3.5100 ;
      RECT 3.8210 2.4165 3.8980 3.5100 ;
      RECT 3.6590 2.4165 3.6850 3.5100 ;
      RECT 3.5510 2.4165 3.5770 3.5100 ;
      RECT 3.4430 2.4165 3.4690 3.5100 ;
      RECT 3.3350 2.4165 3.3610 3.5100 ;
      RECT 3.2270 2.4165 3.2530 3.5100 ;
      RECT 3.1190 2.4165 3.1450 3.5100 ;
      RECT 3.0110 2.4165 3.0370 3.5100 ;
      RECT 2.9030 2.4165 2.9290 3.5100 ;
      RECT 2.7950 2.4165 2.8210 3.5100 ;
      RECT 2.6870 2.4165 2.7130 3.5100 ;
      RECT 2.5790 2.4165 2.6050 3.5100 ;
      RECT 2.4710 2.4165 2.4970 3.5100 ;
      RECT 2.3630 2.4165 2.3890 3.5100 ;
      RECT 2.2550 2.4165 2.2810 3.5100 ;
      RECT 2.1470 2.4165 2.1730 3.5100 ;
      RECT 2.0390 2.4165 2.0650 3.5100 ;
      RECT 1.9310 2.4165 1.9570 3.5100 ;
      RECT 1.8230 2.4165 1.8490 3.5100 ;
      RECT 1.7150 2.4165 1.7410 3.5100 ;
      RECT 1.6070 2.4165 1.6330 3.5100 ;
      RECT 1.4990 2.4165 1.5250 3.5100 ;
      RECT 1.3910 2.4165 1.4170 3.5100 ;
      RECT 1.2830 2.4165 1.3090 3.5100 ;
      RECT 1.1750 2.4165 1.2010 3.5100 ;
      RECT 1.0670 2.4165 1.0930 3.5100 ;
      RECT 0.9590 2.4165 0.9850 3.5100 ;
      RECT 0.8510 2.4165 0.8770 3.5100 ;
      RECT 0.7430 2.4165 0.7690 3.5100 ;
      RECT 0.6350 2.4165 0.6610 3.5100 ;
      RECT 0.5270 2.4165 0.5530 3.5100 ;
      RECT 0.4190 2.4165 0.4450 3.5100 ;
      RECT 0.3110 2.4165 0.3370 3.5100 ;
      RECT 0.2030 2.4165 0.2290 3.5100 ;
      RECT 0.0000 2.4165 0.0850 3.5100 ;
      RECT 5.1800 3.4965 5.3080 4.5900 ;
      RECT 5.1660 4.1620 5.3080 4.4845 ;
      RECT 5.0180 3.8890 5.0800 4.5900 ;
      RECT 5.0040 4.1985 5.0800 4.3520 ;
      RECT 5.0180 3.4965 5.0440 4.5900 ;
      RECT 5.0180 3.6175 5.0580 3.8570 ;
      RECT 5.0180 3.4965 5.0800 3.5855 ;
      RECT 4.7210 3.9470 4.9270 4.5900 ;
      RECT 4.9010 3.4965 4.9270 4.5900 ;
      RECT 4.7210 4.2240 4.9410 4.4820 ;
      RECT 4.7210 3.4965 4.8190 4.5900 ;
      RECT 4.3040 3.4965 4.3870 4.5900 ;
      RECT 4.3040 3.5850 4.4010 4.5205 ;
      RECT 9.5270 3.4965 9.6120 4.5900 ;
      RECT 9.3830 3.4965 9.4090 4.5900 ;
      RECT 9.2750 3.4965 9.3010 4.5900 ;
      RECT 9.1670 3.4965 9.1930 4.5900 ;
      RECT 9.0590 3.4965 9.0850 4.5900 ;
      RECT 8.9510 3.4965 8.9770 4.5900 ;
      RECT 8.8430 3.4965 8.8690 4.5900 ;
      RECT 8.7350 3.4965 8.7610 4.5900 ;
      RECT 8.6270 3.4965 8.6530 4.5900 ;
      RECT 8.5190 3.4965 8.5450 4.5900 ;
      RECT 8.4110 3.4965 8.4370 4.5900 ;
      RECT 8.3030 3.4965 8.3290 4.5900 ;
      RECT 8.1950 3.4965 8.2210 4.5900 ;
      RECT 8.0870 3.4965 8.1130 4.5900 ;
      RECT 7.9790 3.4965 8.0050 4.5900 ;
      RECT 7.8710 3.4965 7.8970 4.5900 ;
      RECT 7.7630 3.4965 7.7890 4.5900 ;
      RECT 7.6550 3.4965 7.6810 4.5900 ;
      RECT 7.5470 3.4965 7.5730 4.5900 ;
      RECT 7.4390 3.4965 7.4650 4.5900 ;
      RECT 7.3310 3.4965 7.3570 4.5900 ;
      RECT 7.2230 3.4965 7.2490 4.5900 ;
      RECT 7.1150 3.4965 7.1410 4.5900 ;
      RECT 7.0070 3.4965 7.0330 4.5900 ;
      RECT 6.8990 3.4965 6.9250 4.5900 ;
      RECT 6.7910 3.4965 6.8170 4.5900 ;
      RECT 6.6830 3.4965 6.7090 4.5900 ;
      RECT 6.5750 3.4965 6.6010 4.5900 ;
      RECT 6.4670 3.4965 6.4930 4.5900 ;
      RECT 6.3590 3.4965 6.3850 4.5900 ;
      RECT 6.2510 3.4965 6.2770 4.5900 ;
      RECT 6.1430 3.4965 6.1690 4.5900 ;
      RECT 6.0350 3.4965 6.0610 4.5900 ;
      RECT 5.9270 3.4965 5.9530 4.5900 ;
      RECT 5.7140 3.4965 5.7910 4.5900 ;
      RECT 3.8210 3.4965 3.8980 4.5900 ;
      RECT 3.6590 3.4965 3.6850 4.5900 ;
      RECT 3.5510 3.4965 3.5770 4.5900 ;
      RECT 3.4430 3.4965 3.4690 4.5900 ;
      RECT 3.3350 3.4965 3.3610 4.5900 ;
      RECT 3.2270 3.4965 3.2530 4.5900 ;
      RECT 3.1190 3.4965 3.1450 4.5900 ;
      RECT 3.0110 3.4965 3.0370 4.5900 ;
      RECT 2.9030 3.4965 2.9290 4.5900 ;
      RECT 2.7950 3.4965 2.8210 4.5900 ;
      RECT 2.6870 3.4965 2.7130 4.5900 ;
      RECT 2.5790 3.4965 2.6050 4.5900 ;
      RECT 2.4710 3.4965 2.4970 4.5900 ;
      RECT 2.3630 3.4965 2.3890 4.5900 ;
      RECT 2.2550 3.4965 2.2810 4.5900 ;
      RECT 2.1470 3.4965 2.1730 4.5900 ;
      RECT 2.0390 3.4965 2.0650 4.5900 ;
      RECT 1.9310 3.4965 1.9570 4.5900 ;
      RECT 1.8230 3.4965 1.8490 4.5900 ;
      RECT 1.7150 3.4965 1.7410 4.5900 ;
      RECT 1.6070 3.4965 1.6330 4.5900 ;
      RECT 1.4990 3.4965 1.5250 4.5900 ;
      RECT 1.3910 3.4965 1.4170 4.5900 ;
      RECT 1.2830 3.4965 1.3090 4.5900 ;
      RECT 1.1750 3.4965 1.2010 4.5900 ;
      RECT 1.0670 3.4965 1.0930 4.5900 ;
      RECT 0.9590 3.4965 0.9850 4.5900 ;
      RECT 0.8510 3.4965 0.8770 4.5900 ;
      RECT 0.7430 3.4965 0.7690 4.5900 ;
      RECT 0.6350 3.4965 0.6610 4.5900 ;
      RECT 0.5270 3.4965 0.5530 4.5900 ;
      RECT 0.4190 3.4965 0.4450 4.5900 ;
      RECT 0.3110 3.4965 0.3370 4.5900 ;
      RECT 0.2030 3.4965 0.2290 4.5900 ;
      RECT 0.0000 3.4965 0.0850 4.5900 ;
      RECT 5.1800 4.5765 5.3080 5.6700 ;
      RECT 5.1660 5.2420 5.3080 5.5645 ;
      RECT 5.0180 4.9690 5.0800 5.6700 ;
      RECT 5.0040 5.2785 5.0800 5.4320 ;
      RECT 5.0180 4.5765 5.0440 5.6700 ;
      RECT 5.0180 4.6975 5.0580 4.9370 ;
      RECT 5.0180 4.5765 5.0800 4.6655 ;
      RECT 4.7210 5.0270 4.9270 5.6700 ;
      RECT 4.9010 4.5765 4.9270 5.6700 ;
      RECT 4.7210 5.3040 4.9410 5.5620 ;
      RECT 4.7210 4.5765 4.8190 5.6700 ;
      RECT 4.3040 4.5765 4.3870 5.6700 ;
      RECT 4.3040 4.6650 4.4010 5.6005 ;
      RECT 9.5270 4.5765 9.6120 5.6700 ;
      RECT 9.3830 4.5765 9.4090 5.6700 ;
      RECT 9.2750 4.5765 9.3010 5.6700 ;
      RECT 9.1670 4.5765 9.1930 5.6700 ;
      RECT 9.0590 4.5765 9.0850 5.6700 ;
      RECT 8.9510 4.5765 8.9770 5.6700 ;
      RECT 8.8430 4.5765 8.8690 5.6700 ;
      RECT 8.7350 4.5765 8.7610 5.6700 ;
      RECT 8.6270 4.5765 8.6530 5.6700 ;
      RECT 8.5190 4.5765 8.5450 5.6700 ;
      RECT 8.4110 4.5765 8.4370 5.6700 ;
      RECT 8.3030 4.5765 8.3290 5.6700 ;
      RECT 8.1950 4.5765 8.2210 5.6700 ;
      RECT 8.0870 4.5765 8.1130 5.6700 ;
      RECT 7.9790 4.5765 8.0050 5.6700 ;
      RECT 7.8710 4.5765 7.8970 5.6700 ;
      RECT 7.7630 4.5765 7.7890 5.6700 ;
      RECT 7.6550 4.5765 7.6810 5.6700 ;
      RECT 7.5470 4.5765 7.5730 5.6700 ;
      RECT 7.4390 4.5765 7.4650 5.6700 ;
      RECT 7.3310 4.5765 7.3570 5.6700 ;
      RECT 7.2230 4.5765 7.2490 5.6700 ;
      RECT 7.1150 4.5765 7.1410 5.6700 ;
      RECT 7.0070 4.5765 7.0330 5.6700 ;
      RECT 6.8990 4.5765 6.9250 5.6700 ;
      RECT 6.7910 4.5765 6.8170 5.6700 ;
      RECT 6.6830 4.5765 6.7090 5.6700 ;
      RECT 6.5750 4.5765 6.6010 5.6700 ;
      RECT 6.4670 4.5765 6.4930 5.6700 ;
      RECT 6.3590 4.5765 6.3850 5.6700 ;
      RECT 6.2510 4.5765 6.2770 5.6700 ;
      RECT 6.1430 4.5765 6.1690 5.6700 ;
      RECT 6.0350 4.5765 6.0610 5.6700 ;
      RECT 5.9270 4.5765 5.9530 5.6700 ;
      RECT 5.7140 4.5765 5.7910 5.6700 ;
      RECT 3.8210 4.5765 3.8980 5.6700 ;
      RECT 3.6590 4.5765 3.6850 5.6700 ;
      RECT 3.5510 4.5765 3.5770 5.6700 ;
      RECT 3.4430 4.5765 3.4690 5.6700 ;
      RECT 3.3350 4.5765 3.3610 5.6700 ;
      RECT 3.2270 4.5765 3.2530 5.6700 ;
      RECT 3.1190 4.5765 3.1450 5.6700 ;
      RECT 3.0110 4.5765 3.0370 5.6700 ;
      RECT 2.9030 4.5765 2.9290 5.6700 ;
      RECT 2.7950 4.5765 2.8210 5.6700 ;
      RECT 2.6870 4.5765 2.7130 5.6700 ;
      RECT 2.5790 4.5765 2.6050 5.6700 ;
      RECT 2.4710 4.5765 2.4970 5.6700 ;
      RECT 2.3630 4.5765 2.3890 5.6700 ;
      RECT 2.2550 4.5765 2.2810 5.6700 ;
      RECT 2.1470 4.5765 2.1730 5.6700 ;
      RECT 2.0390 4.5765 2.0650 5.6700 ;
      RECT 1.9310 4.5765 1.9570 5.6700 ;
      RECT 1.8230 4.5765 1.8490 5.6700 ;
      RECT 1.7150 4.5765 1.7410 5.6700 ;
      RECT 1.6070 4.5765 1.6330 5.6700 ;
      RECT 1.4990 4.5765 1.5250 5.6700 ;
      RECT 1.3910 4.5765 1.4170 5.6700 ;
      RECT 1.2830 4.5765 1.3090 5.6700 ;
      RECT 1.1750 4.5765 1.2010 5.6700 ;
      RECT 1.0670 4.5765 1.0930 5.6700 ;
      RECT 0.9590 4.5765 0.9850 5.6700 ;
      RECT 0.8510 4.5765 0.8770 5.6700 ;
      RECT 0.7430 4.5765 0.7690 5.6700 ;
      RECT 0.6350 4.5765 0.6610 5.6700 ;
      RECT 0.5270 4.5765 0.5530 5.6700 ;
      RECT 0.4190 4.5765 0.4450 5.6700 ;
      RECT 0.3110 4.5765 0.3370 5.6700 ;
      RECT 0.2030 4.5765 0.2290 5.6700 ;
      RECT 0.0000 4.5765 0.0850 5.6700 ;
      RECT 5.1800 5.6565 5.3080 6.7500 ;
      RECT 5.1660 6.3220 5.3080 6.6445 ;
      RECT 5.0180 6.0490 5.0800 6.7500 ;
      RECT 5.0040 6.3585 5.0800 6.5120 ;
      RECT 5.0180 5.6565 5.0440 6.7500 ;
      RECT 5.0180 5.7775 5.0580 6.0170 ;
      RECT 5.0180 5.6565 5.0800 5.7455 ;
      RECT 4.7210 6.1070 4.9270 6.7500 ;
      RECT 4.9010 5.6565 4.9270 6.7500 ;
      RECT 4.7210 6.3840 4.9410 6.6420 ;
      RECT 4.7210 5.6565 4.8190 6.7500 ;
      RECT 4.3040 5.6565 4.3870 6.7500 ;
      RECT 4.3040 5.7450 4.4010 6.6805 ;
      RECT 9.5270 5.6565 9.6120 6.7500 ;
      RECT 9.3830 5.6565 9.4090 6.7500 ;
      RECT 9.2750 5.6565 9.3010 6.7500 ;
      RECT 9.1670 5.6565 9.1930 6.7500 ;
      RECT 9.0590 5.6565 9.0850 6.7500 ;
      RECT 8.9510 5.6565 8.9770 6.7500 ;
      RECT 8.8430 5.6565 8.8690 6.7500 ;
      RECT 8.7350 5.6565 8.7610 6.7500 ;
      RECT 8.6270 5.6565 8.6530 6.7500 ;
      RECT 8.5190 5.6565 8.5450 6.7500 ;
      RECT 8.4110 5.6565 8.4370 6.7500 ;
      RECT 8.3030 5.6565 8.3290 6.7500 ;
      RECT 8.1950 5.6565 8.2210 6.7500 ;
      RECT 8.0870 5.6565 8.1130 6.7500 ;
      RECT 7.9790 5.6565 8.0050 6.7500 ;
      RECT 7.8710 5.6565 7.8970 6.7500 ;
      RECT 7.7630 5.6565 7.7890 6.7500 ;
      RECT 7.6550 5.6565 7.6810 6.7500 ;
      RECT 7.5470 5.6565 7.5730 6.7500 ;
      RECT 7.4390 5.6565 7.4650 6.7500 ;
      RECT 7.3310 5.6565 7.3570 6.7500 ;
      RECT 7.2230 5.6565 7.2490 6.7500 ;
      RECT 7.1150 5.6565 7.1410 6.7500 ;
      RECT 7.0070 5.6565 7.0330 6.7500 ;
      RECT 6.8990 5.6565 6.9250 6.7500 ;
      RECT 6.7910 5.6565 6.8170 6.7500 ;
      RECT 6.6830 5.6565 6.7090 6.7500 ;
      RECT 6.5750 5.6565 6.6010 6.7500 ;
      RECT 6.4670 5.6565 6.4930 6.7500 ;
      RECT 6.3590 5.6565 6.3850 6.7500 ;
      RECT 6.2510 5.6565 6.2770 6.7500 ;
      RECT 6.1430 5.6565 6.1690 6.7500 ;
      RECT 6.0350 5.6565 6.0610 6.7500 ;
      RECT 5.9270 5.6565 5.9530 6.7500 ;
      RECT 5.7140 5.6565 5.7910 6.7500 ;
      RECT 3.8210 5.6565 3.8980 6.7500 ;
      RECT 3.6590 5.6565 3.6850 6.7500 ;
      RECT 3.5510 5.6565 3.5770 6.7500 ;
      RECT 3.4430 5.6565 3.4690 6.7500 ;
      RECT 3.3350 5.6565 3.3610 6.7500 ;
      RECT 3.2270 5.6565 3.2530 6.7500 ;
      RECT 3.1190 5.6565 3.1450 6.7500 ;
      RECT 3.0110 5.6565 3.0370 6.7500 ;
      RECT 2.9030 5.6565 2.9290 6.7500 ;
      RECT 2.7950 5.6565 2.8210 6.7500 ;
      RECT 2.6870 5.6565 2.7130 6.7500 ;
      RECT 2.5790 5.6565 2.6050 6.7500 ;
      RECT 2.4710 5.6565 2.4970 6.7500 ;
      RECT 2.3630 5.6565 2.3890 6.7500 ;
      RECT 2.2550 5.6565 2.2810 6.7500 ;
      RECT 2.1470 5.6565 2.1730 6.7500 ;
      RECT 2.0390 5.6565 2.0650 6.7500 ;
      RECT 1.9310 5.6565 1.9570 6.7500 ;
      RECT 1.8230 5.6565 1.8490 6.7500 ;
      RECT 1.7150 5.6565 1.7410 6.7500 ;
      RECT 1.6070 5.6565 1.6330 6.7500 ;
      RECT 1.4990 5.6565 1.5250 6.7500 ;
      RECT 1.3910 5.6565 1.4170 6.7500 ;
      RECT 1.2830 5.6565 1.3090 6.7500 ;
      RECT 1.1750 5.6565 1.2010 6.7500 ;
      RECT 1.0670 5.6565 1.0930 6.7500 ;
      RECT 0.9590 5.6565 0.9850 6.7500 ;
      RECT 0.8510 5.6565 0.8770 6.7500 ;
      RECT 0.7430 5.6565 0.7690 6.7500 ;
      RECT 0.6350 5.6565 0.6610 6.7500 ;
      RECT 0.5270 5.6565 0.5530 6.7500 ;
      RECT 0.4190 5.6565 0.4450 6.7500 ;
      RECT 0.3110 5.6565 0.3370 6.7500 ;
      RECT 0.2030 5.6565 0.2290 6.7500 ;
      RECT 0.0000 5.6565 0.0850 6.7500 ;
      RECT 5.1800 6.7365 5.3080 7.8300 ;
      RECT 5.1660 7.4020 5.3080 7.7245 ;
      RECT 5.0180 7.1290 5.0800 7.8300 ;
      RECT 5.0040 7.4385 5.0800 7.5920 ;
      RECT 5.0180 6.7365 5.0440 7.8300 ;
      RECT 5.0180 6.8575 5.0580 7.0970 ;
      RECT 5.0180 6.7365 5.0800 6.8255 ;
      RECT 4.7210 7.1870 4.9270 7.8300 ;
      RECT 4.9010 6.7365 4.9270 7.8300 ;
      RECT 4.7210 7.4640 4.9410 7.7220 ;
      RECT 4.7210 6.7365 4.8190 7.8300 ;
      RECT 4.3040 6.7365 4.3870 7.8300 ;
      RECT 4.3040 6.8250 4.4010 7.7605 ;
      RECT 9.5270 6.7365 9.6120 7.8300 ;
      RECT 9.3830 6.7365 9.4090 7.8300 ;
      RECT 9.2750 6.7365 9.3010 7.8300 ;
      RECT 9.1670 6.7365 9.1930 7.8300 ;
      RECT 9.0590 6.7365 9.0850 7.8300 ;
      RECT 8.9510 6.7365 8.9770 7.8300 ;
      RECT 8.8430 6.7365 8.8690 7.8300 ;
      RECT 8.7350 6.7365 8.7610 7.8300 ;
      RECT 8.6270 6.7365 8.6530 7.8300 ;
      RECT 8.5190 6.7365 8.5450 7.8300 ;
      RECT 8.4110 6.7365 8.4370 7.8300 ;
      RECT 8.3030 6.7365 8.3290 7.8300 ;
      RECT 8.1950 6.7365 8.2210 7.8300 ;
      RECT 8.0870 6.7365 8.1130 7.8300 ;
      RECT 7.9790 6.7365 8.0050 7.8300 ;
      RECT 7.8710 6.7365 7.8970 7.8300 ;
      RECT 7.7630 6.7365 7.7890 7.8300 ;
      RECT 7.6550 6.7365 7.6810 7.8300 ;
      RECT 7.5470 6.7365 7.5730 7.8300 ;
      RECT 7.4390 6.7365 7.4650 7.8300 ;
      RECT 7.3310 6.7365 7.3570 7.8300 ;
      RECT 7.2230 6.7365 7.2490 7.8300 ;
      RECT 7.1150 6.7365 7.1410 7.8300 ;
      RECT 7.0070 6.7365 7.0330 7.8300 ;
      RECT 6.8990 6.7365 6.9250 7.8300 ;
      RECT 6.7910 6.7365 6.8170 7.8300 ;
      RECT 6.6830 6.7365 6.7090 7.8300 ;
      RECT 6.5750 6.7365 6.6010 7.8300 ;
      RECT 6.4670 6.7365 6.4930 7.8300 ;
      RECT 6.3590 6.7365 6.3850 7.8300 ;
      RECT 6.2510 6.7365 6.2770 7.8300 ;
      RECT 6.1430 6.7365 6.1690 7.8300 ;
      RECT 6.0350 6.7365 6.0610 7.8300 ;
      RECT 5.9270 6.7365 5.9530 7.8300 ;
      RECT 5.7140 6.7365 5.7910 7.8300 ;
      RECT 3.8210 6.7365 3.8980 7.8300 ;
      RECT 3.6590 6.7365 3.6850 7.8300 ;
      RECT 3.5510 6.7365 3.5770 7.8300 ;
      RECT 3.4430 6.7365 3.4690 7.8300 ;
      RECT 3.3350 6.7365 3.3610 7.8300 ;
      RECT 3.2270 6.7365 3.2530 7.8300 ;
      RECT 3.1190 6.7365 3.1450 7.8300 ;
      RECT 3.0110 6.7365 3.0370 7.8300 ;
      RECT 2.9030 6.7365 2.9290 7.8300 ;
      RECT 2.7950 6.7365 2.8210 7.8300 ;
      RECT 2.6870 6.7365 2.7130 7.8300 ;
      RECT 2.5790 6.7365 2.6050 7.8300 ;
      RECT 2.4710 6.7365 2.4970 7.8300 ;
      RECT 2.3630 6.7365 2.3890 7.8300 ;
      RECT 2.2550 6.7365 2.2810 7.8300 ;
      RECT 2.1470 6.7365 2.1730 7.8300 ;
      RECT 2.0390 6.7365 2.0650 7.8300 ;
      RECT 1.9310 6.7365 1.9570 7.8300 ;
      RECT 1.8230 6.7365 1.8490 7.8300 ;
      RECT 1.7150 6.7365 1.7410 7.8300 ;
      RECT 1.6070 6.7365 1.6330 7.8300 ;
      RECT 1.4990 6.7365 1.5250 7.8300 ;
      RECT 1.3910 6.7365 1.4170 7.8300 ;
      RECT 1.2830 6.7365 1.3090 7.8300 ;
      RECT 1.1750 6.7365 1.2010 7.8300 ;
      RECT 1.0670 6.7365 1.0930 7.8300 ;
      RECT 0.9590 6.7365 0.9850 7.8300 ;
      RECT 0.8510 6.7365 0.8770 7.8300 ;
      RECT 0.7430 6.7365 0.7690 7.8300 ;
      RECT 0.6350 6.7365 0.6610 7.8300 ;
      RECT 0.5270 6.7365 0.5530 7.8300 ;
      RECT 0.4190 6.7365 0.4450 7.8300 ;
      RECT 0.3110 6.7365 0.3370 7.8300 ;
      RECT 0.2030 6.7365 0.2290 7.8300 ;
      RECT 0.0000 6.7365 0.0850 7.8300 ;
      RECT 5.1800 7.8165 5.3080 8.9100 ;
      RECT 5.1660 8.4820 5.3080 8.8045 ;
      RECT 5.0180 8.2090 5.0800 8.9100 ;
      RECT 5.0040 8.5185 5.0800 8.6720 ;
      RECT 5.0180 7.8165 5.0440 8.9100 ;
      RECT 5.0180 7.9375 5.0580 8.1770 ;
      RECT 5.0180 7.8165 5.0800 7.9055 ;
      RECT 4.7210 8.2670 4.9270 8.9100 ;
      RECT 4.9010 7.8165 4.9270 8.9100 ;
      RECT 4.7210 8.5440 4.9410 8.8020 ;
      RECT 4.7210 7.8165 4.8190 8.9100 ;
      RECT 4.3040 7.8165 4.3870 8.9100 ;
      RECT 4.3040 7.9050 4.4010 8.8405 ;
      RECT 9.5270 7.8165 9.6120 8.9100 ;
      RECT 9.3830 7.8165 9.4090 8.9100 ;
      RECT 9.2750 7.8165 9.3010 8.9100 ;
      RECT 9.1670 7.8165 9.1930 8.9100 ;
      RECT 9.0590 7.8165 9.0850 8.9100 ;
      RECT 8.9510 7.8165 8.9770 8.9100 ;
      RECT 8.8430 7.8165 8.8690 8.9100 ;
      RECT 8.7350 7.8165 8.7610 8.9100 ;
      RECT 8.6270 7.8165 8.6530 8.9100 ;
      RECT 8.5190 7.8165 8.5450 8.9100 ;
      RECT 8.4110 7.8165 8.4370 8.9100 ;
      RECT 8.3030 7.8165 8.3290 8.9100 ;
      RECT 8.1950 7.8165 8.2210 8.9100 ;
      RECT 8.0870 7.8165 8.1130 8.9100 ;
      RECT 7.9790 7.8165 8.0050 8.9100 ;
      RECT 7.8710 7.8165 7.8970 8.9100 ;
      RECT 7.7630 7.8165 7.7890 8.9100 ;
      RECT 7.6550 7.8165 7.6810 8.9100 ;
      RECT 7.5470 7.8165 7.5730 8.9100 ;
      RECT 7.4390 7.8165 7.4650 8.9100 ;
      RECT 7.3310 7.8165 7.3570 8.9100 ;
      RECT 7.2230 7.8165 7.2490 8.9100 ;
      RECT 7.1150 7.8165 7.1410 8.9100 ;
      RECT 7.0070 7.8165 7.0330 8.9100 ;
      RECT 6.8990 7.8165 6.9250 8.9100 ;
      RECT 6.7910 7.8165 6.8170 8.9100 ;
      RECT 6.6830 7.8165 6.7090 8.9100 ;
      RECT 6.5750 7.8165 6.6010 8.9100 ;
      RECT 6.4670 7.8165 6.4930 8.9100 ;
      RECT 6.3590 7.8165 6.3850 8.9100 ;
      RECT 6.2510 7.8165 6.2770 8.9100 ;
      RECT 6.1430 7.8165 6.1690 8.9100 ;
      RECT 6.0350 7.8165 6.0610 8.9100 ;
      RECT 5.9270 7.8165 5.9530 8.9100 ;
      RECT 5.7140 7.8165 5.7910 8.9100 ;
      RECT 3.8210 7.8165 3.8980 8.9100 ;
      RECT 3.6590 7.8165 3.6850 8.9100 ;
      RECT 3.5510 7.8165 3.5770 8.9100 ;
      RECT 3.4430 7.8165 3.4690 8.9100 ;
      RECT 3.3350 7.8165 3.3610 8.9100 ;
      RECT 3.2270 7.8165 3.2530 8.9100 ;
      RECT 3.1190 7.8165 3.1450 8.9100 ;
      RECT 3.0110 7.8165 3.0370 8.9100 ;
      RECT 2.9030 7.8165 2.9290 8.9100 ;
      RECT 2.7950 7.8165 2.8210 8.9100 ;
      RECT 2.6870 7.8165 2.7130 8.9100 ;
      RECT 2.5790 7.8165 2.6050 8.9100 ;
      RECT 2.4710 7.8165 2.4970 8.9100 ;
      RECT 2.3630 7.8165 2.3890 8.9100 ;
      RECT 2.2550 7.8165 2.2810 8.9100 ;
      RECT 2.1470 7.8165 2.1730 8.9100 ;
      RECT 2.0390 7.8165 2.0650 8.9100 ;
      RECT 1.9310 7.8165 1.9570 8.9100 ;
      RECT 1.8230 7.8165 1.8490 8.9100 ;
      RECT 1.7150 7.8165 1.7410 8.9100 ;
      RECT 1.6070 7.8165 1.6330 8.9100 ;
      RECT 1.4990 7.8165 1.5250 8.9100 ;
      RECT 1.3910 7.8165 1.4170 8.9100 ;
      RECT 1.2830 7.8165 1.3090 8.9100 ;
      RECT 1.1750 7.8165 1.2010 8.9100 ;
      RECT 1.0670 7.8165 1.0930 8.9100 ;
      RECT 0.9590 7.8165 0.9850 8.9100 ;
      RECT 0.8510 7.8165 0.8770 8.9100 ;
      RECT 0.7430 7.8165 0.7690 8.9100 ;
      RECT 0.6350 7.8165 0.6610 8.9100 ;
      RECT 0.5270 7.8165 0.5530 8.9100 ;
      RECT 0.4190 7.8165 0.4450 8.9100 ;
      RECT 0.3110 7.8165 0.3370 8.9100 ;
      RECT 0.2030 7.8165 0.2290 8.9100 ;
      RECT 0.0000 7.8165 0.0850 8.9100 ;
      RECT 5.1800 8.8965 5.3080 9.9900 ;
      RECT 5.1660 9.5620 5.3080 9.8845 ;
      RECT 5.0180 9.2890 5.0800 9.9900 ;
      RECT 5.0040 9.5985 5.0800 9.7520 ;
      RECT 5.0180 8.8965 5.0440 9.9900 ;
      RECT 5.0180 9.0175 5.0580 9.2570 ;
      RECT 5.0180 8.8965 5.0800 8.9855 ;
      RECT 4.7210 9.3470 4.9270 9.9900 ;
      RECT 4.9010 8.8965 4.9270 9.9900 ;
      RECT 4.7210 9.6240 4.9410 9.8820 ;
      RECT 4.7210 8.8965 4.8190 9.9900 ;
      RECT 4.3040 8.8965 4.3870 9.9900 ;
      RECT 4.3040 8.9850 4.4010 9.9205 ;
      RECT 9.5270 8.8965 9.6120 9.9900 ;
      RECT 9.3830 8.8965 9.4090 9.9900 ;
      RECT 9.2750 8.8965 9.3010 9.9900 ;
      RECT 9.1670 8.8965 9.1930 9.9900 ;
      RECT 9.0590 8.8965 9.0850 9.9900 ;
      RECT 8.9510 8.8965 8.9770 9.9900 ;
      RECT 8.8430 8.8965 8.8690 9.9900 ;
      RECT 8.7350 8.8965 8.7610 9.9900 ;
      RECT 8.6270 8.8965 8.6530 9.9900 ;
      RECT 8.5190 8.8965 8.5450 9.9900 ;
      RECT 8.4110 8.8965 8.4370 9.9900 ;
      RECT 8.3030 8.8965 8.3290 9.9900 ;
      RECT 8.1950 8.8965 8.2210 9.9900 ;
      RECT 8.0870 8.8965 8.1130 9.9900 ;
      RECT 7.9790 8.8965 8.0050 9.9900 ;
      RECT 7.8710 8.8965 7.8970 9.9900 ;
      RECT 7.7630 8.8965 7.7890 9.9900 ;
      RECT 7.6550 8.8965 7.6810 9.9900 ;
      RECT 7.5470 8.8965 7.5730 9.9900 ;
      RECT 7.4390 8.8965 7.4650 9.9900 ;
      RECT 7.3310 8.8965 7.3570 9.9900 ;
      RECT 7.2230 8.8965 7.2490 9.9900 ;
      RECT 7.1150 8.8965 7.1410 9.9900 ;
      RECT 7.0070 8.8965 7.0330 9.9900 ;
      RECT 6.8990 8.8965 6.9250 9.9900 ;
      RECT 6.7910 8.8965 6.8170 9.9900 ;
      RECT 6.6830 8.8965 6.7090 9.9900 ;
      RECT 6.5750 8.8965 6.6010 9.9900 ;
      RECT 6.4670 8.8965 6.4930 9.9900 ;
      RECT 6.3590 8.8965 6.3850 9.9900 ;
      RECT 6.2510 8.8965 6.2770 9.9900 ;
      RECT 6.1430 8.8965 6.1690 9.9900 ;
      RECT 6.0350 8.8965 6.0610 9.9900 ;
      RECT 5.9270 8.8965 5.9530 9.9900 ;
      RECT 5.7140 8.8965 5.7910 9.9900 ;
      RECT 3.8210 8.8965 3.8980 9.9900 ;
      RECT 3.6590 8.8965 3.6850 9.9900 ;
      RECT 3.5510 8.8965 3.5770 9.9900 ;
      RECT 3.4430 8.8965 3.4690 9.9900 ;
      RECT 3.3350 8.8965 3.3610 9.9900 ;
      RECT 3.2270 8.8965 3.2530 9.9900 ;
      RECT 3.1190 8.8965 3.1450 9.9900 ;
      RECT 3.0110 8.8965 3.0370 9.9900 ;
      RECT 2.9030 8.8965 2.9290 9.9900 ;
      RECT 2.7950 8.8965 2.8210 9.9900 ;
      RECT 2.6870 8.8965 2.7130 9.9900 ;
      RECT 2.5790 8.8965 2.6050 9.9900 ;
      RECT 2.4710 8.8965 2.4970 9.9900 ;
      RECT 2.3630 8.8965 2.3890 9.9900 ;
      RECT 2.2550 8.8965 2.2810 9.9900 ;
      RECT 2.1470 8.8965 2.1730 9.9900 ;
      RECT 2.0390 8.8965 2.0650 9.9900 ;
      RECT 1.9310 8.8965 1.9570 9.9900 ;
      RECT 1.8230 8.8965 1.8490 9.9900 ;
      RECT 1.7150 8.8965 1.7410 9.9900 ;
      RECT 1.6070 8.8965 1.6330 9.9900 ;
      RECT 1.4990 8.8965 1.5250 9.9900 ;
      RECT 1.3910 8.8965 1.4170 9.9900 ;
      RECT 1.2830 8.8965 1.3090 9.9900 ;
      RECT 1.1750 8.8965 1.2010 9.9900 ;
      RECT 1.0670 8.8965 1.0930 9.9900 ;
      RECT 0.9590 8.8965 0.9850 9.9900 ;
      RECT 0.8510 8.8965 0.8770 9.9900 ;
      RECT 0.7430 8.8965 0.7690 9.9900 ;
      RECT 0.6350 8.8965 0.6610 9.9900 ;
      RECT 0.5270 8.8965 0.5530 9.9900 ;
      RECT 0.4190 8.8965 0.4450 9.9900 ;
      RECT 0.3110 8.8965 0.3370 9.9900 ;
      RECT 0.2030 8.8965 0.2290 9.9900 ;
      RECT 0.0000 8.8965 0.0850 9.9900 ;
      RECT 5.1800 9.9765 5.3080 11.0700 ;
      RECT 5.1660 10.6420 5.3080 10.9645 ;
      RECT 5.0180 10.3690 5.0800 11.0700 ;
      RECT 5.0040 10.6785 5.0800 10.8320 ;
      RECT 5.0180 9.9765 5.0440 11.0700 ;
      RECT 5.0180 10.0975 5.0580 10.3370 ;
      RECT 5.0180 9.9765 5.0800 10.0655 ;
      RECT 4.7210 10.4270 4.9270 11.0700 ;
      RECT 4.9010 9.9765 4.9270 11.0700 ;
      RECT 4.7210 10.7040 4.9410 10.9620 ;
      RECT 4.7210 9.9765 4.8190 11.0700 ;
      RECT 4.3040 9.9765 4.3870 11.0700 ;
      RECT 4.3040 10.0650 4.4010 11.0005 ;
      RECT 9.5270 9.9765 9.6120 11.0700 ;
      RECT 9.3830 9.9765 9.4090 11.0700 ;
      RECT 9.2750 9.9765 9.3010 11.0700 ;
      RECT 9.1670 9.9765 9.1930 11.0700 ;
      RECT 9.0590 9.9765 9.0850 11.0700 ;
      RECT 8.9510 9.9765 8.9770 11.0700 ;
      RECT 8.8430 9.9765 8.8690 11.0700 ;
      RECT 8.7350 9.9765 8.7610 11.0700 ;
      RECT 8.6270 9.9765 8.6530 11.0700 ;
      RECT 8.5190 9.9765 8.5450 11.0700 ;
      RECT 8.4110 9.9765 8.4370 11.0700 ;
      RECT 8.3030 9.9765 8.3290 11.0700 ;
      RECT 8.1950 9.9765 8.2210 11.0700 ;
      RECT 8.0870 9.9765 8.1130 11.0700 ;
      RECT 7.9790 9.9765 8.0050 11.0700 ;
      RECT 7.8710 9.9765 7.8970 11.0700 ;
      RECT 7.7630 9.9765 7.7890 11.0700 ;
      RECT 7.6550 9.9765 7.6810 11.0700 ;
      RECT 7.5470 9.9765 7.5730 11.0700 ;
      RECT 7.4390 9.9765 7.4650 11.0700 ;
      RECT 7.3310 9.9765 7.3570 11.0700 ;
      RECT 7.2230 9.9765 7.2490 11.0700 ;
      RECT 7.1150 9.9765 7.1410 11.0700 ;
      RECT 7.0070 9.9765 7.0330 11.0700 ;
      RECT 6.8990 9.9765 6.9250 11.0700 ;
      RECT 6.7910 9.9765 6.8170 11.0700 ;
      RECT 6.6830 9.9765 6.7090 11.0700 ;
      RECT 6.5750 9.9765 6.6010 11.0700 ;
      RECT 6.4670 9.9765 6.4930 11.0700 ;
      RECT 6.3590 9.9765 6.3850 11.0700 ;
      RECT 6.2510 9.9765 6.2770 11.0700 ;
      RECT 6.1430 9.9765 6.1690 11.0700 ;
      RECT 6.0350 9.9765 6.0610 11.0700 ;
      RECT 5.9270 9.9765 5.9530 11.0700 ;
      RECT 5.7140 9.9765 5.7910 11.0700 ;
      RECT 3.8210 9.9765 3.8980 11.0700 ;
      RECT 3.6590 9.9765 3.6850 11.0700 ;
      RECT 3.5510 9.9765 3.5770 11.0700 ;
      RECT 3.4430 9.9765 3.4690 11.0700 ;
      RECT 3.3350 9.9765 3.3610 11.0700 ;
      RECT 3.2270 9.9765 3.2530 11.0700 ;
      RECT 3.1190 9.9765 3.1450 11.0700 ;
      RECT 3.0110 9.9765 3.0370 11.0700 ;
      RECT 2.9030 9.9765 2.9290 11.0700 ;
      RECT 2.7950 9.9765 2.8210 11.0700 ;
      RECT 2.6870 9.9765 2.7130 11.0700 ;
      RECT 2.5790 9.9765 2.6050 11.0700 ;
      RECT 2.4710 9.9765 2.4970 11.0700 ;
      RECT 2.3630 9.9765 2.3890 11.0700 ;
      RECT 2.2550 9.9765 2.2810 11.0700 ;
      RECT 2.1470 9.9765 2.1730 11.0700 ;
      RECT 2.0390 9.9765 2.0650 11.0700 ;
      RECT 1.9310 9.9765 1.9570 11.0700 ;
      RECT 1.8230 9.9765 1.8490 11.0700 ;
      RECT 1.7150 9.9765 1.7410 11.0700 ;
      RECT 1.6070 9.9765 1.6330 11.0700 ;
      RECT 1.4990 9.9765 1.5250 11.0700 ;
      RECT 1.3910 9.9765 1.4170 11.0700 ;
      RECT 1.2830 9.9765 1.3090 11.0700 ;
      RECT 1.1750 9.9765 1.2010 11.0700 ;
      RECT 1.0670 9.9765 1.0930 11.0700 ;
      RECT 0.9590 9.9765 0.9850 11.0700 ;
      RECT 0.8510 9.9765 0.8770 11.0700 ;
      RECT 0.7430 9.9765 0.7690 11.0700 ;
      RECT 0.6350 9.9765 0.6610 11.0700 ;
      RECT 0.5270 9.9765 0.5530 11.0700 ;
      RECT 0.4190 9.9765 0.4450 11.0700 ;
      RECT 0.3110 9.9765 0.3370 11.0700 ;
      RECT 0.2030 9.9765 0.2290 11.0700 ;
      RECT 0.0000 9.9765 0.0850 11.0700 ;
      RECT 5.1800 11.0565 5.3080 12.1500 ;
      RECT 5.1660 11.7220 5.3080 12.0445 ;
      RECT 5.0180 11.4490 5.0800 12.1500 ;
      RECT 5.0040 11.7585 5.0800 11.9120 ;
      RECT 5.0180 11.0565 5.0440 12.1500 ;
      RECT 5.0180 11.1775 5.0580 11.4170 ;
      RECT 5.0180 11.0565 5.0800 11.1455 ;
      RECT 4.7210 11.5070 4.9270 12.1500 ;
      RECT 4.9010 11.0565 4.9270 12.1500 ;
      RECT 4.7210 11.7840 4.9410 12.0420 ;
      RECT 4.7210 11.0565 4.8190 12.1500 ;
      RECT 4.3040 11.0565 4.3870 12.1500 ;
      RECT 4.3040 11.1450 4.4010 12.0805 ;
      RECT 9.5270 11.0565 9.6120 12.1500 ;
      RECT 9.3830 11.0565 9.4090 12.1500 ;
      RECT 9.2750 11.0565 9.3010 12.1500 ;
      RECT 9.1670 11.0565 9.1930 12.1500 ;
      RECT 9.0590 11.0565 9.0850 12.1500 ;
      RECT 8.9510 11.0565 8.9770 12.1500 ;
      RECT 8.8430 11.0565 8.8690 12.1500 ;
      RECT 8.7350 11.0565 8.7610 12.1500 ;
      RECT 8.6270 11.0565 8.6530 12.1500 ;
      RECT 8.5190 11.0565 8.5450 12.1500 ;
      RECT 8.4110 11.0565 8.4370 12.1500 ;
      RECT 8.3030 11.0565 8.3290 12.1500 ;
      RECT 8.1950 11.0565 8.2210 12.1500 ;
      RECT 8.0870 11.0565 8.1130 12.1500 ;
      RECT 7.9790 11.0565 8.0050 12.1500 ;
      RECT 7.8710 11.0565 7.8970 12.1500 ;
      RECT 7.7630 11.0565 7.7890 12.1500 ;
      RECT 7.6550 11.0565 7.6810 12.1500 ;
      RECT 7.5470 11.0565 7.5730 12.1500 ;
      RECT 7.4390 11.0565 7.4650 12.1500 ;
      RECT 7.3310 11.0565 7.3570 12.1500 ;
      RECT 7.2230 11.0565 7.2490 12.1500 ;
      RECT 7.1150 11.0565 7.1410 12.1500 ;
      RECT 7.0070 11.0565 7.0330 12.1500 ;
      RECT 6.8990 11.0565 6.9250 12.1500 ;
      RECT 6.7910 11.0565 6.8170 12.1500 ;
      RECT 6.6830 11.0565 6.7090 12.1500 ;
      RECT 6.5750 11.0565 6.6010 12.1500 ;
      RECT 6.4670 11.0565 6.4930 12.1500 ;
      RECT 6.3590 11.0565 6.3850 12.1500 ;
      RECT 6.2510 11.0565 6.2770 12.1500 ;
      RECT 6.1430 11.0565 6.1690 12.1500 ;
      RECT 6.0350 11.0565 6.0610 12.1500 ;
      RECT 5.9270 11.0565 5.9530 12.1500 ;
      RECT 5.7140 11.0565 5.7910 12.1500 ;
      RECT 3.8210 11.0565 3.8980 12.1500 ;
      RECT 3.6590 11.0565 3.6850 12.1500 ;
      RECT 3.5510 11.0565 3.5770 12.1500 ;
      RECT 3.4430 11.0565 3.4690 12.1500 ;
      RECT 3.3350 11.0565 3.3610 12.1500 ;
      RECT 3.2270 11.0565 3.2530 12.1500 ;
      RECT 3.1190 11.0565 3.1450 12.1500 ;
      RECT 3.0110 11.0565 3.0370 12.1500 ;
      RECT 2.9030 11.0565 2.9290 12.1500 ;
      RECT 2.7950 11.0565 2.8210 12.1500 ;
      RECT 2.6870 11.0565 2.7130 12.1500 ;
      RECT 2.5790 11.0565 2.6050 12.1500 ;
      RECT 2.4710 11.0565 2.4970 12.1500 ;
      RECT 2.3630 11.0565 2.3890 12.1500 ;
      RECT 2.2550 11.0565 2.2810 12.1500 ;
      RECT 2.1470 11.0565 2.1730 12.1500 ;
      RECT 2.0390 11.0565 2.0650 12.1500 ;
      RECT 1.9310 11.0565 1.9570 12.1500 ;
      RECT 1.8230 11.0565 1.8490 12.1500 ;
      RECT 1.7150 11.0565 1.7410 12.1500 ;
      RECT 1.6070 11.0565 1.6330 12.1500 ;
      RECT 1.4990 11.0565 1.5250 12.1500 ;
      RECT 1.3910 11.0565 1.4170 12.1500 ;
      RECT 1.2830 11.0565 1.3090 12.1500 ;
      RECT 1.1750 11.0565 1.2010 12.1500 ;
      RECT 1.0670 11.0565 1.0930 12.1500 ;
      RECT 0.9590 11.0565 0.9850 12.1500 ;
      RECT 0.8510 11.0565 0.8770 12.1500 ;
      RECT 0.7430 11.0565 0.7690 12.1500 ;
      RECT 0.6350 11.0565 0.6610 12.1500 ;
      RECT 0.5270 11.0565 0.5530 12.1500 ;
      RECT 0.4190 11.0565 0.4450 12.1500 ;
      RECT 0.3110 11.0565 0.3370 12.1500 ;
      RECT 0.2030 11.0565 0.2290 12.1500 ;
      RECT 0.0000 11.0565 0.0850 12.1500 ;
      RECT 5.1800 12.1365 5.3080 13.2300 ;
      RECT 5.1660 12.8020 5.3080 13.1245 ;
      RECT 5.0180 12.5290 5.0800 13.2300 ;
      RECT 5.0040 12.8385 5.0800 12.9920 ;
      RECT 5.0180 12.1365 5.0440 13.2300 ;
      RECT 5.0180 12.2575 5.0580 12.4970 ;
      RECT 5.0180 12.1365 5.0800 12.2255 ;
      RECT 4.7210 12.5870 4.9270 13.2300 ;
      RECT 4.9010 12.1365 4.9270 13.2300 ;
      RECT 4.7210 12.8640 4.9410 13.1220 ;
      RECT 4.7210 12.1365 4.8190 13.2300 ;
      RECT 4.3040 12.1365 4.3870 13.2300 ;
      RECT 4.3040 12.2250 4.4010 13.1605 ;
      RECT 9.5270 12.1365 9.6120 13.2300 ;
      RECT 9.3830 12.1365 9.4090 13.2300 ;
      RECT 9.2750 12.1365 9.3010 13.2300 ;
      RECT 9.1670 12.1365 9.1930 13.2300 ;
      RECT 9.0590 12.1365 9.0850 13.2300 ;
      RECT 8.9510 12.1365 8.9770 13.2300 ;
      RECT 8.8430 12.1365 8.8690 13.2300 ;
      RECT 8.7350 12.1365 8.7610 13.2300 ;
      RECT 8.6270 12.1365 8.6530 13.2300 ;
      RECT 8.5190 12.1365 8.5450 13.2300 ;
      RECT 8.4110 12.1365 8.4370 13.2300 ;
      RECT 8.3030 12.1365 8.3290 13.2300 ;
      RECT 8.1950 12.1365 8.2210 13.2300 ;
      RECT 8.0870 12.1365 8.1130 13.2300 ;
      RECT 7.9790 12.1365 8.0050 13.2300 ;
      RECT 7.8710 12.1365 7.8970 13.2300 ;
      RECT 7.7630 12.1365 7.7890 13.2300 ;
      RECT 7.6550 12.1365 7.6810 13.2300 ;
      RECT 7.5470 12.1365 7.5730 13.2300 ;
      RECT 7.4390 12.1365 7.4650 13.2300 ;
      RECT 7.3310 12.1365 7.3570 13.2300 ;
      RECT 7.2230 12.1365 7.2490 13.2300 ;
      RECT 7.1150 12.1365 7.1410 13.2300 ;
      RECT 7.0070 12.1365 7.0330 13.2300 ;
      RECT 6.8990 12.1365 6.9250 13.2300 ;
      RECT 6.7910 12.1365 6.8170 13.2300 ;
      RECT 6.6830 12.1365 6.7090 13.2300 ;
      RECT 6.5750 12.1365 6.6010 13.2300 ;
      RECT 6.4670 12.1365 6.4930 13.2300 ;
      RECT 6.3590 12.1365 6.3850 13.2300 ;
      RECT 6.2510 12.1365 6.2770 13.2300 ;
      RECT 6.1430 12.1365 6.1690 13.2300 ;
      RECT 6.0350 12.1365 6.0610 13.2300 ;
      RECT 5.9270 12.1365 5.9530 13.2300 ;
      RECT 5.7140 12.1365 5.7910 13.2300 ;
      RECT 3.8210 12.1365 3.8980 13.2300 ;
      RECT 3.6590 12.1365 3.6850 13.2300 ;
      RECT 3.5510 12.1365 3.5770 13.2300 ;
      RECT 3.4430 12.1365 3.4690 13.2300 ;
      RECT 3.3350 12.1365 3.3610 13.2300 ;
      RECT 3.2270 12.1365 3.2530 13.2300 ;
      RECT 3.1190 12.1365 3.1450 13.2300 ;
      RECT 3.0110 12.1365 3.0370 13.2300 ;
      RECT 2.9030 12.1365 2.9290 13.2300 ;
      RECT 2.7950 12.1365 2.8210 13.2300 ;
      RECT 2.6870 12.1365 2.7130 13.2300 ;
      RECT 2.5790 12.1365 2.6050 13.2300 ;
      RECT 2.4710 12.1365 2.4970 13.2300 ;
      RECT 2.3630 12.1365 2.3890 13.2300 ;
      RECT 2.2550 12.1365 2.2810 13.2300 ;
      RECT 2.1470 12.1365 2.1730 13.2300 ;
      RECT 2.0390 12.1365 2.0650 13.2300 ;
      RECT 1.9310 12.1365 1.9570 13.2300 ;
      RECT 1.8230 12.1365 1.8490 13.2300 ;
      RECT 1.7150 12.1365 1.7410 13.2300 ;
      RECT 1.6070 12.1365 1.6330 13.2300 ;
      RECT 1.4990 12.1365 1.5250 13.2300 ;
      RECT 1.3910 12.1365 1.4170 13.2300 ;
      RECT 1.2830 12.1365 1.3090 13.2300 ;
      RECT 1.1750 12.1365 1.2010 13.2300 ;
      RECT 1.0670 12.1365 1.0930 13.2300 ;
      RECT 0.9590 12.1365 0.9850 13.2300 ;
      RECT 0.8510 12.1365 0.8770 13.2300 ;
      RECT 0.7430 12.1365 0.7690 13.2300 ;
      RECT 0.6350 12.1365 0.6610 13.2300 ;
      RECT 0.5270 12.1365 0.5530 13.2300 ;
      RECT 0.4190 12.1365 0.4450 13.2300 ;
      RECT 0.3110 12.1365 0.3370 13.2300 ;
      RECT 0.2030 12.1365 0.2290 13.2300 ;
      RECT 0.0000 12.1365 0.0850 13.2300 ;
      RECT 5.1800 13.2165 5.3080 14.3100 ;
      RECT 5.1660 13.8820 5.3080 14.2045 ;
      RECT 5.0180 13.6090 5.0800 14.3100 ;
      RECT 5.0040 13.9185 5.0800 14.0720 ;
      RECT 5.0180 13.2165 5.0440 14.3100 ;
      RECT 5.0180 13.3375 5.0580 13.5770 ;
      RECT 5.0180 13.2165 5.0800 13.3055 ;
      RECT 4.7210 13.6670 4.9270 14.3100 ;
      RECT 4.9010 13.2165 4.9270 14.3100 ;
      RECT 4.7210 13.9440 4.9410 14.2020 ;
      RECT 4.7210 13.2165 4.8190 14.3100 ;
      RECT 4.3040 13.2165 4.3870 14.3100 ;
      RECT 4.3040 13.3050 4.4010 14.2405 ;
      RECT 9.5270 13.2165 9.6120 14.3100 ;
      RECT 9.3830 13.2165 9.4090 14.3100 ;
      RECT 9.2750 13.2165 9.3010 14.3100 ;
      RECT 9.1670 13.2165 9.1930 14.3100 ;
      RECT 9.0590 13.2165 9.0850 14.3100 ;
      RECT 8.9510 13.2165 8.9770 14.3100 ;
      RECT 8.8430 13.2165 8.8690 14.3100 ;
      RECT 8.7350 13.2165 8.7610 14.3100 ;
      RECT 8.6270 13.2165 8.6530 14.3100 ;
      RECT 8.5190 13.2165 8.5450 14.3100 ;
      RECT 8.4110 13.2165 8.4370 14.3100 ;
      RECT 8.3030 13.2165 8.3290 14.3100 ;
      RECT 8.1950 13.2165 8.2210 14.3100 ;
      RECT 8.0870 13.2165 8.1130 14.3100 ;
      RECT 7.9790 13.2165 8.0050 14.3100 ;
      RECT 7.8710 13.2165 7.8970 14.3100 ;
      RECT 7.7630 13.2165 7.7890 14.3100 ;
      RECT 7.6550 13.2165 7.6810 14.3100 ;
      RECT 7.5470 13.2165 7.5730 14.3100 ;
      RECT 7.4390 13.2165 7.4650 14.3100 ;
      RECT 7.3310 13.2165 7.3570 14.3100 ;
      RECT 7.2230 13.2165 7.2490 14.3100 ;
      RECT 7.1150 13.2165 7.1410 14.3100 ;
      RECT 7.0070 13.2165 7.0330 14.3100 ;
      RECT 6.8990 13.2165 6.9250 14.3100 ;
      RECT 6.7910 13.2165 6.8170 14.3100 ;
      RECT 6.6830 13.2165 6.7090 14.3100 ;
      RECT 6.5750 13.2165 6.6010 14.3100 ;
      RECT 6.4670 13.2165 6.4930 14.3100 ;
      RECT 6.3590 13.2165 6.3850 14.3100 ;
      RECT 6.2510 13.2165 6.2770 14.3100 ;
      RECT 6.1430 13.2165 6.1690 14.3100 ;
      RECT 6.0350 13.2165 6.0610 14.3100 ;
      RECT 5.9270 13.2165 5.9530 14.3100 ;
      RECT 5.7140 13.2165 5.7910 14.3100 ;
      RECT 3.8210 13.2165 3.8980 14.3100 ;
      RECT 3.6590 13.2165 3.6850 14.3100 ;
      RECT 3.5510 13.2165 3.5770 14.3100 ;
      RECT 3.4430 13.2165 3.4690 14.3100 ;
      RECT 3.3350 13.2165 3.3610 14.3100 ;
      RECT 3.2270 13.2165 3.2530 14.3100 ;
      RECT 3.1190 13.2165 3.1450 14.3100 ;
      RECT 3.0110 13.2165 3.0370 14.3100 ;
      RECT 2.9030 13.2165 2.9290 14.3100 ;
      RECT 2.7950 13.2165 2.8210 14.3100 ;
      RECT 2.6870 13.2165 2.7130 14.3100 ;
      RECT 2.5790 13.2165 2.6050 14.3100 ;
      RECT 2.4710 13.2165 2.4970 14.3100 ;
      RECT 2.3630 13.2165 2.3890 14.3100 ;
      RECT 2.2550 13.2165 2.2810 14.3100 ;
      RECT 2.1470 13.2165 2.1730 14.3100 ;
      RECT 2.0390 13.2165 2.0650 14.3100 ;
      RECT 1.9310 13.2165 1.9570 14.3100 ;
      RECT 1.8230 13.2165 1.8490 14.3100 ;
      RECT 1.7150 13.2165 1.7410 14.3100 ;
      RECT 1.6070 13.2165 1.6330 14.3100 ;
      RECT 1.4990 13.2165 1.5250 14.3100 ;
      RECT 1.3910 13.2165 1.4170 14.3100 ;
      RECT 1.2830 13.2165 1.3090 14.3100 ;
      RECT 1.1750 13.2165 1.2010 14.3100 ;
      RECT 1.0670 13.2165 1.0930 14.3100 ;
      RECT 0.9590 13.2165 0.9850 14.3100 ;
      RECT 0.8510 13.2165 0.8770 14.3100 ;
      RECT 0.7430 13.2165 0.7690 14.3100 ;
      RECT 0.6350 13.2165 0.6610 14.3100 ;
      RECT 0.5270 13.2165 0.5530 14.3100 ;
      RECT 0.4190 13.2165 0.4450 14.3100 ;
      RECT 0.3110 13.2165 0.3370 14.3100 ;
      RECT 0.2030 13.2165 0.2290 14.3100 ;
      RECT 0.0000 13.2165 0.0850 14.3100 ;
      RECT 5.1800 14.2965 5.3080 15.3900 ;
      RECT 5.1660 14.9620 5.3080 15.2845 ;
      RECT 5.0180 14.6890 5.0800 15.3900 ;
      RECT 5.0040 14.9985 5.0800 15.1520 ;
      RECT 5.0180 14.2965 5.0440 15.3900 ;
      RECT 5.0180 14.4175 5.0580 14.6570 ;
      RECT 5.0180 14.2965 5.0800 14.3855 ;
      RECT 4.7210 14.7470 4.9270 15.3900 ;
      RECT 4.9010 14.2965 4.9270 15.3900 ;
      RECT 4.7210 15.0240 4.9410 15.2820 ;
      RECT 4.7210 14.2965 4.8190 15.3900 ;
      RECT 4.3040 14.2965 4.3870 15.3900 ;
      RECT 4.3040 14.3850 4.4010 15.3205 ;
      RECT 9.5270 14.2965 9.6120 15.3900 ;
      RECT 9.3830 14.2965 9.4090 15.3900 ;
      RECT 9.2750 14.2965 9.3010 15.3900 ;
      RECT 9.1670 14.2965 9.1930 15.3900 ;
      RECT 9.0590 14.2965 9.0850 15.3900 ;
      RECT 8.9510 14.2965 8.9770 15.3900 ;
      RECT 8.8430 14.2965 8.8690 15.3900 ;
      RECT 8.7350 14.2965 8.7610 15.3900 ;
      RECT 8.6270 14.2965 8.6530 15.3900 ;
      RECT 8.5190 14.2965 8.5450 15.3900 ;
      RECT 8.4110 14.2965 8.4370 15.3900 ;
      RECT 8.3030 14.2965 8.3290 15.3900 ;
      RECT 8.1950 14.2965 8.2210 15.3900 ;
      RECT 8.0870 14.2965 8.1130 15.3900 ;
      RECT 7.9790 14.2965 8.0050 15.3900 ;
      RECT 7.8710 14.2965 7.8970 15.3900 ;
      RECT 7.7630 14.2965 7.7890 15.3900 ;
      RECT 7.6550 14.2965 7.6810 15.3900 ;
      RECT 7.5470 14.2965 7.5730 15.3900 ;
      RECT 7.4390 14.2965 7.4650 15.3900 ;
      RECT 7.3310 14.2965 7.3570 15.3900 ;
      RECT 7.2230 14.2965 7.2490 15.3900 ;
      RECT 7.1150 14.2965 7.1410 15.3900 ;
      RECT 7.0070 14.2965 7.0330 15.3900 ;
      RECT 6.8990 14.2965 6.9250 15.3900 ;
      RECT 6.7910 14.2965 6.8170 15.3900 ;
      RECT 6.6830 14.2965 6.7090 15.3900 ;
      RECT 6.5750 14.2965 6.6010 15.3900 ;
      RECT 6.4670 14.2965 6.4930 15.3900 ;
      RECT 6.3590 14.2965 6.3850 15.3900 ;
      RECT 6.2510 14.2965 6.2770 15.3900 ;
      RECT 6.1430 14.2965 6.1690 15.3900 ;
      RECT 6.0350 14.2965 6.0610 15.3900 ;
      RECT 5.9270 14.2965 5.9530 15.3900 ;
      RECT 5.7140 14.2965 5.7910 15.3900 ;
      RECT 3.8210 14.2965 3.8980 15.3900 ;
      RECT 3.6590 14.2965 3.6850 15.3900 ;
      RECT 3.5510 14.2965 3.5770 15.3900 ;
      RECT 3.4430 14.2965 3.4690 15.3900 ;
      RECT 3.3350 14.2965 3.3610 15.3900 ;
      RECT 3.2270 14.2965 3.2530 15.3900 ;
      RECT 3.1190 14.2965 3.1450 15.3900 ;
      RECT 3.0110 14.2965 3.0370 15.3900 ;
      RECT 2.9030 14.2965 2.9290 15.3900 ;
      RECT 2.7950 14.2965 2.8210 15.3900 ;
      RECT 2.6870 14.2965 2.7130 15.3900 ;
      RECT 2.5790 14.2965 2.6050 15.3900 ;
      RECT 2.4710 14.2965 2.4970 15.3900 ;
      RECT 2.3630 14.2965 2.3890 15.3900 ;
      RECT 2.2550 14.2965 2.2810 15.3900 ;
      RECT 2.1470 14.2965 2.1730 15.3900 ;
      RECT 2.0390 14.2965 2.0650 15.3900 ;
      RECT 1.9310 14.2965 1.9570 15.3900 ;
      RECT 1.8230 14.2965 1.8490 15.3900 ;
      RECT 1.7150 14.2965 1.7410 15.3900 ;
      RECT 1.6070 14.2965 1.6330 15.3900 ;
      RECT 1.4990 14.2965 1.5250 15.3900 ;
      RECT 1.3910 14.2965 1.4170 15.3900 ;
      RECT 1.2830 14.2965 1.3090 15.3900 ;
      RECT 1.1750 14.2965 1.2010 15.3900 ;
      RECT 1.0670 14.2965 1.0930 15.3900 ;
      RECT 0.9590 14.2965 0.9850 15.3900 ;
      RECT 0.8510 14.2965 0.8770 15.3900 ;
      RECT 0.7430 14.2965 0.7690 15.3900 ;
      RECT 0.6350 14.2965 0.6610 15.3900 ;
      RECT 0.5270 14.2965 0.5530 15.3900 ;
      RECT 0.4190 14.2965 0.4450 15.3900 ;
      RECT 0.3110 14.2965 0.3370 15.3900 ;
      RECT 0.2030 14.2965 0.2290 15.3900 ;
      RECT 0.0000 14.2965 0.0850 15.3900 ;
      RECT 5.1800 15.3765 5.3080 16.4700 ;
      RECT 5.1660 16.0420 5.3080 16.3645 ;
      RECT 5.0180 15.7690 5.0800 16.4700 ;
      RECT 5.0040 16.0785 5.0800 16.2320 ;
      RECT 5.0180 15.3765 5.0440 16.4700 ;
      RECT 5.0180 15.4975 5.0580 15.7370 ;
      RECT 5.0180 15.3765 5.0800 15.4655 ;
      RECT 4.7210 15.8270 4.9270 16.4700 ;
      RECT 4.9010 15.3765 4.9270 16.4700 ;
      RECT 4.7210 16.1040 4.9410 16.3620 ;
      RECT 4.7210 15.3765 4.8190 16.4700 ;
      RECT 4.3040 15.3765 4.3870 16.4700 ;
      RECT 4.3040 15.4650 4.4010 16.4005 ;
      RECT 9.5270 15.3765 9.6120 16.4700 ;
      RECT 9.3830 15.3765 9.4090 16.4700 ;
      RECT 9.2750 15.3765 9.3010 16.4700 ;
      RECT 9.1670 15.3765 9.1930 16.4700 ;
      RECT 9.0590 15.3765 9.0850 16.4700 ;
      RECT 8.9510 15.3765 8.9770 16.4700 ;
      RECT 8.8430 15.3765 8.8690 16.4700 ;
      RECT 8.7350 15.3765 8.7610 16.4700 ;
      RECT 8.6270 15.3765 8.6530 16.4700 ;
      RECT 8.5190 15.3765 8.5450 16.4700 ;
      RECT 8.4110 15.3765 8.4370 16.4700 ;
      RECT 8.3030 15.3765 8.3290 16.4700 ;
      RECT 8.1950 15.3765 8.2210 16.4700 ;
      RECT 8.0870 15.3765 8.1130 16.4700 ;
      RECT 7.9790 15.3765 8.0050 16.4700 ;
      RECT 7.8710 15.3765 7.8970 16.4700 ;
      RECT 7.7630 15.3765 7.7890 16.4700 ;
      RECT 7.6550 15.3765 7.6810 16.4700 ;
      RECT 7.5470 15.3765 7.5730 16.4700 ;
      RECT 7.4390 15.3765 7.4650 16.4700 ;
      RECT 7.3310 15.3765 7.3570 16.4700 ;
      RECT 7.2230 15.3765 7.2490 16.4700 ;
      RECT 7.1150 15.3765 7.1410 16.4700 ;
      RECT 7.0070 15.3765 7.0330 16.4700 ;
      RECT 6.8990 15.3765 6.9250 16.4700 ;
      RECT 6.7910 15.3765 6.8170 16.4700 ;
      RECT 6.6830 15.3765 6.7090 16.4700 ;
      RECT 6.5750 15.3765 6.6010 16.4700 ;
      RECT 6.4670 15.3765 6.4930 16.4700 ;
      RECT 6.3590 15.3765 6.3850 16.4700 ;
      RECT 6.2510 15.3765 6.2770 16.4700 ;
      RECT 6.1430 15.3765 6.1690 16.4700 ;
      RECT 6.0350 15.3765 6.0610 16.4700 ;
      RECT 5.9270 15.3765 5.9530 16.4700 ;
      RECT 5.7140 15.3765 5.7910 16.4700 ;
      RECT 3.8210 15.3765 3.8980 16.4700 ;
      RECT 3.6590 15.3765 3.6850 16.4700 ;
      RECT 3.5510 15.3765 3.5770 16.4700 ;
      RECT 3.4430 15.3765 3.4690 16.4700 ;
      RECT 3.3350 15.3765 3.3610 16.4700 ;
      RECT 3.2270 15.3765 3.2530 16.4700 ;
      RECT 3.1190 15.3765 3.1450 16.4700 ;
      RECT 3.0110 15.3765 3.0370 16.4700 ;
      RECT 2.9030 15.3765 2.9290 16.4700 ;
      RECT 2.7950 15.3765 2.8210 16.4700 ;
      RECT 2.6870 15.3765 2.7130 16.4700 ;
      RECT 2.5790 15.3765 2.6050 16.4700 ;
      RECT 2.4710 15.3765 2.4970 16.4700 ;
      RECT 2.3630 15.3765 2.3890 16.4700 ;
      RECT 2.2550 15.3765 2.2810 16.4700 ;
      RECT 2.1470 15.3765 2.1730 16.4700 ;
      RECT 2.0390 15.3765 2.0650 16.4700 ;
      RECT 1.9310 15.3765 1.9570 16.4700 ;
      RECT 1.8230 15.3765 1.8490 16.4700 ;
      RECT 1.7150 15.3765 1.7410 16.4700 ;
      RECT 1.6070 15.3765 1.6330 16.4700 ;
      RECT 1.4990 15.3765 1.5250 16.4700 ;
      RECT 1.3910 15.3765 1.4170 16.4700 ;
      RECT 1.2830 15.3765 1.3090 16.4700 ;
      RECT 1.1750 15.3765 1.2010 16.4700 ;
      RECT 1.0670 15.3765 1.0930 16.4700 ;
      RECT 0.9590 15.3765 0.9850 16.4700 ;
      RECT 0.8510 15.3765 0.8770 16.4700 ;
      RECT 0.7430 15.3765 0.7690 16.4700 ;
      RECT 0.6350 15.3765 0.6610 16.4700 ;
      RECT 0.5270 15.3765 0.5530 16.4700 ;
      RECT 0.4190 15.3765 0.4450 16.4700 ;
      RECT 0.3110 15.3765 0.3370 16.4700 ;
      RECT 0.2030 15.3765 0.2290 16.4700 ;
      RECT 0.0000 15.3765 0.0850 16.4700 ;
      RECT 5.1800 16.4565 5.3080 17.5500 ;
      RECT 5.1660 17.1220 5.3080 17.4445 ;
      RECT 5.0180 16.8490 5.0800 17.5500 ;
      RECT 5.0040 17.1585 5.0800 17.3120 ;
      RECT 5.0180 16.4565 5.0440 17.5500 ;
      RECT 5.0180 16.5775 5.0580 16.8170 ;
      RECT 5.0180 16.4565 5.0800 16.5455 ;
      RECT 4.7210 16.9070 4.9270 17.5500 ;
      RECT 4.9010 16.4565 4.9270 17.5500 ;
      RECT 4.7210 17.1840 4.9410 17.4420 ;
      RECT 4.7210 16.4565 4.8190 17.5500 ;
      RECT 4.3040 16.4565 4.3870 17.5500 ;
      RECT 4.3040 16.5450 4.4010 17.4805 ;
      RECT 9.5270 16.4565 9.6120 17.5500 ;
      RECT 9.3830 16.4565 9.4090 17.5500 ;
      RECT 9.2750 16.4565 9.3010 17.5500 ;
      RECT 9.1670 16.4565 9.1930 17.5500 ;
      RECT 9.0590 16.4565 9.0850 17.5500 ;
      RECT 8.9510 16.4565 8.9770 17.5500 ;
      RECT 8.8430 16.4565 8.8690 17.5500 ;
      RECT 8.7350 16.4565 8.7610 17.5500 ;
      RECT 8.6270 16.4565 8.6530 17.5500 ;
      RECT 8.5190 16.4565 8.5450 17.5500 ;
      RECT 8.4110 16.4565 8.4370 17.5500 ;
      RECT 8.3030 16.4565 8.3290 17.5500 ;
      RECT 8.1950 16.4565 8.2210 17.5500 ;
      RECT 8.0870 16.4565 8.1130 17.5500 ;
      RECT 7.9790 16.4565 8.0050 17.5500 ;
      RECT 7.8710 16.4565 7.8970 17.5500 ;
      RECT 7.7630 16.4565 7.7890 17.5500 ;
      RECT 7.6550 16.4565 7.6810 17.5500 ;
      RECT 7.5470 16.4565 7.5730 17.5500 ;
      RECT 7.4390 16.4565 7.4650 17.5500 ;
      RECT 7.3310 16.4565 7.3570 17.5500 ;
      RECT 7.2230 16.4565 7.2490 17.5500 ;
      RECT 7.1150 16.4565 7.1410 17.5500 ;
      RECT 7.0070 16.4565 7.0330 17.5500 ;
      RECT 6.8990 16.4565 6.9250 17.5500 ;
      RECT 6.7910 16.4565 6.8170 17.5500 ;
      RECT 6.6830 16.4565 6.7090 17.5500 ;
      RECT 6.5750 16.4565 6.6010 17.5500 ;
      RECT 6.4670 16.4565 6.4930 17.5500 ;
      RECT 6.3590 16.4565 6.3850 17.5500 ;
      RECT 6.2510 16.4565 6.2770 17.5500 ;
      RECT 6.1430 16.4565 6.1690 17.5500 ;
      RECT 6.0350 16.4565 6.0610 17.5500 ;
      RECT 5.9270 16.4565 5.9530 17.5500 ;
      RECT 5.7140 16.4565 5.7910 17.5500 ;
      RECT 3.8210 16.4565 3.8980 17.5500 ;
      RECT 3.6590 16.4565 3.6850 17.5500 ;
      RECT 3.5510 16.4565 3.5770 17.5500 ;
      RECT 3.4430 16.4565 3.4690 17.5500 ;
      RECT 3.3350 16.4565 3.3610 17.5500 ;
      RECT 3.2270 16.4565 3.2530 17.5500 ;
      RECT 3.1190 16.4565 3.1450 17.5500 ;
      RECT 3.0110 16.4565 3.0370 17.5500 ;
      RECT 2.9030 16.4565 2.9290 17.5500 ;
      RECT 2.7950 16.4565 2.8210 17.5500 ;
      RECT 2.6870 16.4565 2.7130 17.5500 ;
      RECT 2.5790 16.4565 2.6050 17.5500 ;
      RECT 2.4710 16.4565 2.4970 17.5500 ;
      RECT 2.3630 16.4565 2.3890 17.5500 ;
      RECT 2.2550 16.4565 2.2810 17.5500 ;
      RECT 2.1470 16.4565 2.1730 17.5500 ;
      RECT 2.0390 16.4565 2.0650 17.5500 ;
      RECT 1.9310 16.4565 1.9570 17.5500 ;
      RECT 1.8230 16.4565 1.8490 17.5500 ;
      RECT 1.7150 16.4565 1.7410 17.5500 ;
      RECT 1.6070 16.4565 1.6330 17.5500 ;
      RECT 1.4990 16.4565 1.5250 17.5500 ;
      RECT 1.3910 16.4565 1.4170 17.5500 ;
      RECT 1.2830 16.4565 1.3090 17.5500 ;
      RECT 1.1750 16.4565 1.2010 17.5500 ;
      RECT 1.0670 16.4565 1.0930 17.5500 ;
      RECT 0.9590 16.4565 0.9850 17.5500 ;
      RECT 0.8510 16.4565 0.8770 17.5500 ;
      RECT 0.7430 16.4565 0.7690 17.5500 ;
      RECT 0.6350 16.4565 0.6610 17.5500 ;
      RECT 0.5270 16.4565 0.5530 17.5500 ;
      RECT 0.4190 16.4565 0.4450 17.5500 ;
      RECT 0.3110 16.4565 0.3370 17.5500 ;
      RECT 0.2030 16.4565 0.2290 17.5500 ;
      RECT 0.0000 16.4565 0.0850 17.5500 ;
      RECT 5.1800 17.5365 5.3080 18.6300 ;
      RECT 5.1660 18.2020 5.3080 18.5245 ;
      RECT 5.0180 17.9290 5.0800 18.6300 ;
      RECT 5.0040 18.2385 5.0800 18.3920 ;
      RECT 5.0180 17.5365 5.0440 18.6300 ;
      RECT 5.0180 17.6575 5.0580 17.8970 ;
      RECT 5.0180 17.5365 5.0800 17.6255 ;
      RECT 4.7210 17.9870 4.9270 18.6300 ;
      RECT 4.9010 17.5365 4.9270 18.6300 ;
      RECT 4.7210 18.2640 4.9410 18.5220 ;
      RECT 4.7210 17.5365 4.8190 18.6300 ;
      RECT 4.3040 17.5365 4.3870 18.6300 ;
      RECT 4.3040 17.6250 4.4010 18.5605 ;
      RECT 9.5270 17.5365 9.6120 18.6300 ;
      RECT 9.3830 17.5365 9.4090 18.6300 ;
      RECT 9.2750 17.5365 9.3010 18.6300 ;
      RECT 9.1670 17.5365 9.1930 18.6300 ;
      RECT 9.0590 17.5365 9.0850 18.6300 ;
      RECT 8.9510 17.5365 8.9770 18.6300 ;
      RECT 8.8430 17.5365 8.8690 18.6300 ;
      RECT 8.7350 17.5365 8.7610 18.6300 ;
      RECT 8.6270 17.5365 8.6530 18.6300 ;
      RECT 8.5190 17.5365 8.5450 18.6300 ;
      RECT 8.4110 17.5365 8.4370 18.6300 ;
      RECT 8.3030 17.5365 8.3290 18.6300 ;
      RECT 8.1950 17.5365 8.2210 18.6300 ;
      RECT 8.0870 17.5365 8.1130 18.6300 ;
      RECT 7.9790 17.5365 8.0050 18.6300 ;
      RECT 7.8710 17.5365 7.8970 18.6300 ;
      RECT 7.7630 17.5365 7.7890 18.6300 ;
      RECT 7.6550 17.5365 7.6810 18.6300 ;
      RECT 7.5470 17.5365 7.5730 18.6300 ;
      RECT 7.4390 17.5365 7.4650 18.6300 ;
      RECT 7.3310 17.5365 7.3570 18.6300 ;
      RECT 7.2230 17.5365 7.2490 18.6300 ;
      RECT 7.1150 17.5365 7.1410 18.6300 ;
      RECT 7.0070 17.5365 7.0330 18.6300 ;
      RECT 6.8990 17.5365 6.9250 18.6300 ;
      RECT 6.7910 17.5365 6.8170 18.6300 ;
      RECT 6.6830 17.5365 6.7090 18.6300 ;
      RECT 6.5750 17.5365 6.6010 18.6300 ;
      RECT 6.4670 17.5365 6.4930 18.6300 ;
      RECT 6.3590 17.5365 6.3850 18.6300 ;
      RECT 6.2510 17.5365 6.2770 18.6300 ;
      RECT 6.1430 17.5365 6.1690 18.6300 ;
      RECT 6.0350 17.5365 6.0610 18.6300 ;
      RECT 5.9270 17.5365 5.9530 18.6300 ;
      RECT 5.7140 17.5365 5.7910 18.6300 ;
      RECT 3.8210 17.5365 3.8980 18.6300 ;
      RECT 3.6590 17.5365 3.6850 18.6300 ;
      RECT 3.5510 17.5365 3.5770 18.6300 ;
      RECT 3.4430 17.5365 3.4690 18.6300 ;
      RECT 3.3350 17.5365 3.3610 18.6300 ;
      RECT 3.2270 17.5365 3.2530 18.6300 ;
      RECT 3.1190 17.5365 3.1450 18.6300 ;
      RECT 3.0110 17.5365 3.0370 18.6300 ;
      RECT 2.9030 17.5365 2.9290 18.6300 ;
      RECT 2.7950 17.5365 2.8210 18.6300 ;
      RECT 2.6870 17.5365 2.7130 18.6300 ;
      RECT 2.5790 17.5365 2.6050 18.6300 ;
      RECT 2.4710 17.5365 2.4970 18.6300 ;
      RECT 2.3630 17.5365 2.3890 18.6300 ;
      RECT 2.2550 17.5365 2.2810 18.6300 ;
      RECT 2.1470 17.5365 2.1730 18.6300 ;
      RECT 2.0390 17.5365 2.0650 18.6300 ;
      RECT 1.9310 17.5365 1.9570 18.6300 ;
      RECT 1.8230 17.5365 1.8490 18.6300 ;
      RECT 1.7150 17.5365 1.7410 18.6300 ;
      RECT 1.6070 17.5365 1.6330 18.6300 ;
      RECT 1.4990 17.5365 1.5250 18.6300 ;
      RECT 1.3910 17.5365 1.4170 18.6300 ;
      RECT 1.2830 17.5365 1.3090 18.6300 ;
      RECT 1.1750 17.5365 1.2010 18.6300 ;
      RECT 1.0670 17.5365 1.0930 18.6300 ;
      RECT 0.9590 17.5365 0.9850 18.6300 ;
      RECT 0.8510 17.5365 0.8770 18.6300 ;
      RECT 0.7430 17.5365 0.7690 18.6300 ;
      RECT 0.6350 17.5365 0.6610 18.6300 ;
      RECT 0.5270 17.5365 0.5530 18.6300 ;
      RECT 0.4190 17.5365 0.4450 18.6300 ;
      RECT 0.3110 17.5365 0.3370 18.6300 ;
      RECT 0.2030 17.5365 0.2290 18.6300 ;
      RECT 0.0000 17.5365 0.0850 18.6300 ;
      RECT 5.1800 18.6165 5.3080 19.7100 ;
      RECT 5.1660 19.2820 5.3080 19.6045 ;
      RECT 5.0180 19.0090 5.0800 19.7100 ;
      RECT 5.0040 19.3185 5.0800 19.4720 ;
      RECT 5.0180 18.6165 5.0440 19.7100 ;
      RECT 5.0180 18.7375 5.0580 18.9770 ;
      RECT 5.0180 18.6165 5.0800 18.7055 ;
      RECT 4.7210 19.0670 4.9270 19.7100 ;
      RECT 4.9010 18.6165 4.9270 19.7100 ;
      RECT 4.7210 19.3440 4.9410 19.6020 ;
      RECT 4.7210 18.6165 4.8190 19.7100 ;
      RECT 4.3040 18.6165 4.3870 19.7100 ;
      RECT 4.3040 18.7050 4.4010 19.6405 ;
      RECT 9.5270 18.6165 9.6120 19.7100 ;
      RECT 9.3830 18.6165 9.4090 19.7100 ;
      RECT 9.2750 18.6165 9.3010 19.7100 ;
      RECT 9.1670 18.6165 9.1930 19.7100 ;
      RECT 9.0590 18.6165 9.0850 19.7100 ;
      RECT 8.9510 18.6165 8.9770 19.7100 ;
      RECT 8.8430 18.6165 8.8690 19.7100 ;
      RECT 8.7350 18.6165 8.7610 19.7100 ;
      RECT 8.6270 18.6165 8.6530 19.7100 ;
      RECT 8.5190 18.6165 8.5450 19.7100 ;
      RECT 8.4110 18.6165 8.4370 19.7100 ;
      RECT 8.3030 18.6165 8.3290 19.7100 ;
      RECT 8.1950 18.6165 8.2210 19.7100 ;
      RECT 8.0870 18.6165 8.1130 19.7100 ;
      RECT 7.9790 18.6165 8.0050 19.7100 ;
      RECT 7.8710 18.6165 7.8970 19.7100 ;
      RECT 7.7630 18.6165 7.7890 19.7100 ;
      RECT 7.6550 18.6165 7.6810 19.7100 ;
      RECT 7.5470 18.6165 7.5730 19.7100 ;
      RECT 7.4390 18.6165 7.4650 19.7100 ;
      RECT 7.3310 18.6165 7.3570 19.7100 ;
      RECT 7.2230 18.6165 7.2490 19.7100 ;
      RECT 7.1150 18.6165 7.1410 19.7100 ;
      RECT 7.0070 18.6165 7.0330 19.7100 ;
      RECT 6.8990 18.6165 6.9250 19.7100 ;
      RECT 6.7910 18.6165 6.8170 19.7100 ;
      RECT 6.6830 18.6165 6.7090 19.7100 ;
      RECT 6.5750 18.6165 6.6010 19.7100 ;
      RECT 6.4670 18.6165 6.4930 19.7100 ;
      RECT 6.3590 18.6165 6.3850 19.7100 ;
      RECT 6.2510 18.6165 6.2770 19.7100 ;
      RECT 6.1430 18.6165 6.1690 19.7100 ;
      RECT 6.0350 18.6165 6.0610 19.7100 ;
      RECT 5.9270 18.6165 5.9530 19.7100 ;
      RECT 5.7140 18.6165 5.7910 19.7100 ;
      RECT 3.8210 18.6165 3.8980 19.7100 ;
      RECT 3.6590 18.6165 3.6850 19.7100 ;
      RECT 3.5510 18.6165 3.5770 19.7100 ;
      RECT 3.4430 18.6165 3.4690 19.7100 ;
      RECT 3.3350 18.6165 3.3610 19.7100 ;
      RECT 3.2270 18.6165 3.2530 19.7100 ;
      RECT 3.1190 18.6165 3.1450 19.7100 ;
      RECT 3.0110 18.6165 3.0370 19.7100 ;
      RECT 2.9030 18.6165 2.9290 19.7100 ;
      RECT 2.7950 18.6165 2.8210 19.7100 ;
      RECT 2.6870 18.6165 2.7130 19.7100 ;
      RECT 2.5790 18.6165 2.6050 19.7100 ;
      RECT 2.4710 18.6165 2.4970 19.7100 ;
      RECT 2.3630 18.6165 2.3890 19.7100 ;
      RECT 2.2550 18.6165 2.2810 19.7100 ;
      RECT 2.1470 18.6165 2.1730 19.7100 ;
      RECT 2.0390 18.6165 2.0650 19.7100 ;
      RECT 1.9310 18.6165 1.9570 19.7100 ;
      RECT 1.8230 18.6165 1.8490 19.7100 ;
      RECT 1.7150 18.6165 1.7410 19.7100 ;
      RECT 1.6070 18.6165 1.6330 19.7100 ;
      RECT 1.4990 18.6165 1.5250 19.7100 ;
      RECT 1.3910 18.6165 1.4170 19.7100 ;
      RECT 1.2830 18.6165 1.3090 19.7100 ;
      RECT 1.1750 18.6165 1.2010 19.7100 ;
      RECT 1.0670 18.6165 1.0930 19.7100 ;
      RECT 0.9590 18.6165 0.9850 19.7100 ;
      RECT 0.8510 18.6165 0.8770 19.7100 ;
      RECT 0.7430 18.6165 0.7690 19.7100 ;
      RECT 0.6350 18.6165 0.6610 19.7100 ;
      RECT 0.5270 18.6165 0.5530 19.7100 ;
      RECT 0.4190 18.6165 0.4450 19.7100 ;
      RECT 0.3110 18.6165 0.3370 19.7100 ;
      RECT 0.2030 18.6165 0.2290 19.7100 ;
      RECT 0.0000 18.6165 0.0850 19.7100 ;
      RECT 5.1800 19.6965 5.3080 20.7900 ;
      RECT 5.1660 20.3620 5.3080 20.6845 ;
      RECT 5.0180 20.0890 5.0800 20.7900 ;
      RECT 5.0040 20.3985 5.0800 20.5520 ;
      RECT 5.0180 19.6965 5.0440 20.7900 ;
      RECT 5.0180 19.8175 5.0580 20.0570 ;
      RECT 5.0180 19.6965 5.0800 19.7855 ;
      RECT 4.7210 20.1470 4.9270 20.7900 ;
      RECT 4.9010 19.6965 4.9270 20.7900 ;
      RECT 4.7210 20.4240 4.9410 20.6820 ;
      RECT 4.7210 19.6965 4.8190 20.7900 ;
      RECT 4.3040 19.6965 4.3870 20.7900 ;
      RECT 4.3040 19.7850 4.4010 20.7205 ;
      RECT 9.5270 19.6965 9.6120 20.7900 ;
      RECT 9.3830 19.6965 9.4090 20.7900 ;
      RECT 9.2750 19.6965 9.3010 20.7900 ;
      RECT 9.1670 19.6965 9.1930 20.7900 ;
      RECT 9.0590 19.6965 9.0850 20.7900 ;
      RECT 8.9510 19.6965 8.9770 20.7900 ;
      RECT 8.8430 19.6965 8.8690 20.7900 ;
      RECT 8.7350 19.6965 8.7610 20.7900 ;
      RECT 8.6270 19.6965 8.6530 20.7900 ;
      RECT 8.5190 19.6965 8.5450 20.7900 ;
      RECT 8.4110 19.6965 8.4370 20.7900 ;
      RECT 8.3030 19.6965 8.3290 20.7900 ;
      RECT 8.1950 19.6965 8.2210 20.7900 ;
      RECT 8.0870 19.6965 8.1130 20.7900 ;
      RECT 7.9790 19.6965 8.0050 20.7900 ;
      RECT 7.8710 19.6965 7.8970 20.7900 ;
      RECT 7.7630 19.6965 7.7890 20.7900 ;
      RECT 7.6550 19.6965 7.6810 20.7900 ;
      RECT 7.5470 19.6965 7.5730 20.7900 ;
      RECT 7.4390 19.6965 7.4650 20.7900 ;
      RECT 7.3310 19.6965 7.3570 20.7900 ;
      RECT 7.2230 19.6965 7.2490 20.7900 ;
      RECT 7.1150 19.6965 7.1410 20.7900 ;
      RECT 7.0070 19.6965 7.0330 20.7900 ;
      RECT 6.8990 19.6965 6.9250 20.7900 ;
      RECT 6.7910 19.6965 6.8170 20.7900 ;
      RECT 6.6830 19.6965 6.7090 20.7900 ;
      RECT 6.5750 19.6965 6.6010 20.7900 ;
      RECT 6.4670 19.6965 6.4930 20.7900 ;
      RECT 6.3590 19.6965 6.3850 20.7900 ;
      RECT 6.2510 19.6965 6.2770 20.7900 ;
      RECT 6.1430 19.6965 6.1690 20.7900 ;
      RECT 6.0350 19.6965 6.0610 20.7900 ;
      RECT 5.9270 19.6965 5.9530 20.7900 ;
      RECT 5.7140 19.6965 5.7910 20.7900 ;
      RECT 3.8210 19.6965 3.8980 20.7900 ;
      RECT 3.6590 19.6965 3.6850 20.7900 ;
      RECT 3.5510 19.6965 3.5770 20.7900 ;
      RECT 3.4430 19.6965 3.4690 20.7900 ;
      RECT 3.3350 19.6965 3.3610 20.7900 ;
      RECT 3.2270 19.6965 3.2530 20.7900 ;
      RECT 3.1190 19.6965 3.1450 20.7900 ;
      RECT 3.0110 19.6965 3.0370 20.7900 ;
      RECT 2.9030 19.6965 2.9290 20.7900 ;
      RECT 2.7950 19.6965 2.8210 20.7900 ;
      RECT 2.6870 19.6965 2.7130 20.7900 ;
      RECT 2.5790 19.6965 2.6050 20.7900 ;
      RECT 2.4710 19.6965 2.4970 20.7900 ;
      RECT 2.3630 19.6965 2.3890 20.7900 ;
      RECT 2.2550 19.6965 2.2810 20.7900 ;
      RECT 2.1470 19.6965 2.1730 20.7900 ;
      RECT 2.0390 19.6965 2.0650 20.7900 ;
      RECT 1.9310 19.6965 1.9570 20.7900 ;
      RECT 1.8230 19.6965 1.8490 20.7900 ;
      RECT 1.7150 19.6965 1.7410 20.7900 ;
      RECT 1.6070 19.6965 1.6330 20.7900 ;
      RECT 1.4990 19.6965 1.5250 20.7900 ;
      RECT 1.3910 19.6965 1.4170 20.7900 ;
      RECT 1.2830 19.6965 1.3090 20.7900 ;
      RECT 1.1750 19.6965 1.2010 20.7900 ;
      RECT 1.0670 19.6965 1.0930 20.7900 ;
      RECT 0.9590 19.6965 0.9850 20.7900 ;
      RECT 0.8510 19.6965 0.8770 20.7900 ;
      RECT 0.7430 19.6965 0.7690 20.7900 ;
      RECT 0.6350 19.6965 0.6610 20.7900 ;
      RECT 0.5270 19.6965 0.5530 20.7900 ;
      RECT 0.4190 19.6965 0.4450 20.7900 ;
      RECT 0.3110 19.6965 0.3370 20.7900 ;
      RECT 0.2030 19.6965 0.2290 20.7900 ;
      RECT 0.0000 19.6965 0.0850 20.7900 ;
      RECT 5.1800 20.7765 5.3080 21.8700 ;
      RECT 5.1660 21.4420 5.3080 21.7645 ;
      RECT 5.0180 21.1690 5.0800 21.8700 ;
      RECT 5.0040 21.4785 5.0800 21.6320 ;
      RECT 5.0180 20.7765 5.0440 21.8700 ;
      RECT 5.0180 20.8975 5.0580 21.1370 ;
      RECT 5.0180 20.7765 5.0800 20.8655 ;
      RECT 4.7210 21.2270 4.9270 21.8700 ;
      RECT 4.9010 20.7765 4.9270 21.8700 ;
      RECT 4.7210 21.5040 4.9410 21.7620 ;
      RECT 4.7210 20.7765 4.8190 21.8700 ;
      RECT 4.3040 20.7765 4.3870 21.8700 ;
      RECT 4.3040 20.8650 4.4010 21.8005 ;
      RECT 9.5270 20.7765 9.6120 21.8700 ;
      RECT 9.3830 20.7765 9.4090 21.8700 ;
      RECT 9.2750 20.7765 9.3010 21.8700 ;
      RECT 9.1670 20.7765 9.1930 21.8700 ;
      RECT 9.0590 20.7765 9.0850 21.8700 ;
      RECT 8.9510 20.7765 8.9770 21.8700 ;
      RECT 8.8430 20.7765 8.8690 21.8700 ;
      RECT 8.7350 20.7765 8.7610 21.8700 ;
      RECT 8.6270 20.7765 8.6530 21.8700 ;
      RECT 8.5190 20.7765 8.5450 21.8700 ;
      RECT 8.4110 20.7765 8.4370 21.8700 ;
      RECT 8.3030 20.7765 8.3290 21.8700 ;
      RECT 8.1950 20.7765 8.2210 21.8700 ;
      RECT 8.0870 20.7765 8.1130 21.8700 ;
      RECT 7.9790 20.7765 8.0050 21.8700 ;
      RECT 7.8710 20.7765 7.8970 21.8700 ;
      RECT 7.7630 20.7765 7.7890 21.8700 ;
      RECT 7.6550 20.7765 7.6810 21.8700 ;
      RECT 7.5470 20.7765 7.5730 21.8700 ;
      RECT 7.4390 20.7765 7.4650 21.8700 ;
      RECT 7.3310 20.7765 7.3570 21.8700 ;
      RECT 7.2230 20.7765 7.2490 21.8700 ;
      RECT 7.1150 20.7765 7.1410 21.8700 ;
      RECT 7.0070 20.7765 7.0330 21.8700 ;
      RECT 6.8990 20.7765 6.9250 21.8700 ;
      RECT 6.7910 20.7765 6.8170 21.8700 ;
      RECT 6.6830 20.7765 6.7090 21.8700 ;
      RECT 6.5750 20.7765 6.6010 21.8700 ;
      RECT 6.4670 20.7765 6.4930 21.8700 ;
      RECT 6.3590 20.7765 6.3850 21.8700 ;
      RECT 6.2510 20.7765 6.2770 21.8700 ;
      RECT 6.1430 20.7765 6.1690 21.8700 ;
      RECT 6.0350 20.7765 6.0610 21.8700 ;
      RECT 5.9270 20.7765 5.9530 21.8700 ;
      RECT 5.7140 20.7765 5.7910 21.8700 ;
      RECT 3.8210 20.7765 3.8980 21.8700 ;
      RECT 3.6590 20.7765 3.6850 21.8700 ;
      RECT 3.5510 20.7765 3.5770 21.8700 ;
      RECT 3.4430 20.7765 3.4690 21.8700 ;
      RECT 3.3350 20.7765 3.3610 21.8700 ;
      RECT 3.2270 20.7765 3.2530 21.8700 ;
      RECT 3.1190 20.7765 3.1450 21.8700 ;
      RECT 3.0110 20.7765 3.0370 21.8700 ;
      RECT 2.9030 20.7765 2.9290 21.8700 ;
      RECT 2.7950 20.7765 2.8210 21.8700 ;
      RECT 2.6870 20.7765 2.7130 21.8700 ;
      RECT 2.5790 20.7765 2.6050 21.8700 ;
      RECT 2.4710 20.7765 2.4970 21.8700 ;
      RECT 2.3630 20.7765 2.3890 21.8700 ;
      RECT 2.2550 20.7765 2.2810 21.8700 ;
      RECT 2.1470 20.7765 2.1730 21.8700 ;
      RECT 2.0390 20.7765 2.0650 21.8700 ;
      RECT 1.9310 20.7765 1.9570 21.8700 ;
      RECT 1.8230 20.7765 1.8490 21.8700 ;
      RECT 1.7150 20.7765 1.7410 21.8700 ;
      RECT 1.6070 20.7765 1.6330 21.8700 ;
      RECT 1.4990 20.7765 1.5250 21.8700 ;
      RECT 1.3910 20.7765 1.4170 21.8700 ;
      RECT 1.2830 20.7765 1.3090 21.8700 ;
      RECT 1.1750 20.7765 1.2010 21.8700 ;
      RECT 1.0670 20.7765 1.0930 21.8700 ;
      RECT 0.9590 20.7765 0.9850 21.8700 ;
      RECT 0.8510 20.7765 0.8770 21.8700 ;
      RECT 0.7430 20.7765 0.7690 21.8700 ;
      RECT 0.6350 20.7765 0.6610 21.8700 ;
      RECT 0.5270 20.7765 0.5530 21.8700 ;
      RECT 0.4190 20.7765 0.4450 21.8700 ;
      RECT 0.3110 20.7765 0.3370 21.8700 ;
      RECT 0.2030 20.7765 0.2290 21.8700 ;
      RECT 0.0000 20.7765 0.0850 21.8700 ;
      RECT 5.1800 21.8565 5.3080 22.9500 ;
      RECT 5.1660 22.5220 5.3080 22.8445 ;
      RECT 5.0180 22.2490 5.0800 22.9500 ;
      RECT 5.0040 22.5585 5.0800 22.7120 ;
      RECT 5.0180 21.8565 5.0440 22.9500 ;
      RECT 5.0180 21.9775 5.0580 22.2170 ;
      RECT 5.0180 21.8565 5.0800 21.9455 ;
      RECT 4.7210 22.3070 4.9270 22.9500 ;
      RECT 4.9010 21.8565 4.9270 22.9500 ;
      RECT 4.7210 22.5840 4.9410 22.8420 ;
      RECT 4.7210 21.8565 4.8190 22.9500 ;
      RECT 4.3040 21.8565 4.3870 22.9500 ;
      RECT 4.3040 21.9450 4.4010 22.8805 ;
      RECT 9.5270 21.8565 9.6120 22.9500 ;
      RECT 9.3830 21.8565 9.4090 22.9500 ;
      RECT 9.2750 21.8565 9.3010 22.9500 ;
      RECT 9.1670 21.8565 9.1930 22.9500 ;
      RECT 9.0590 21.8565 9.0850 22.9500 ;
      RECT 8.9510 21.8565 8.9770 22.9500 ;
      RECT 8.8430 21.8565 8.8690 22.9500 ;
      RECT 8.7350 21.8565 8.7610 22.9500 ;
      RECT 8.6270 21.8565 8.6530 22.9500 ;
      RECT 8.5190 21.8565 8.5450 22.9500 ;
      RECT 8.4110 21.8565 8.4370 22.9500 ;
      RECT 8.3030 21.8565 8.3290 22.9500 ;
      RECT 8.1950 21.8565 8.2210 22.9500 ;
      RECT 8.0870 21.8565 8.1130 22.9500 ;
      RECT 7.9790 21.8565 8.0050 22.9500 ;
      RECT 7.8710 21.8565 7.8970 22.9500 ;
      RECT 7.7630 21.8565 7.7890 22.9500 ;
      RECT 7.6550 21.8565 7.6810 22.9500 ;
      RECT 7.5470 21.8565 7.5730 22.9500 ;
      RECT 7.4390 21.8565 7.4650 22.9500 ;
      RECT 7.3310 21.8565 7.3570 22.9500 ;
      RECT 7.2230 21.8565 7.2490 22.9500 ;
      RECT 7.1150 21.8565 7.1410 22.9500 ;
      RECT 7.0070 21.8565 7.0330 22.9500 ;
      RECT 6.8990 21.8565 6.9250 22.9500 ;
      RECT 6.7910 21.8565 6.8170 22.9500 ;
      RECT 6.6830 21.8565 6.7090 22.9500 ;
      RECT 6.5750 21.8565 6.6010 22.9500 ;
      RECT 6.4670 21.8565 6.4930 22.9500 ;
      RECT 6.3590 21.8565 6.3850 22.9500 ;
      RECT 6.2510 21.8565 6.2770 22.9500 ;
      RECT 6.1430 21.8565 6.1690 22.9500 ;
      RECT 6.0350 21.8565 6.0610 22.9500 ;
      RECT 5.9270 21.8565 5.9530 22.9500 ;
      RECT 5.7140 21.8565 5.7910 22.9500 ;
      RECT 3.8210 21.8565 3.8980 22.9500 ;
      RECT 3.6590 21.8565 3.6850 22.9500 ;
      RECT 3.5510 21.8565 3.5770 22.9500 ;
      RECT 3.4430 21.8565 3.4690 22.9500 ;
      RECT 3.3350 21.8565 3.3610 22.9500 ;
      RECT 3.2270 21.8565 3.2530 22.9500 ;
      RECT 3.1190 21.8565 3.1450 22.9500 ;
      RECT 3.0110 21.8565 3.0370 22.9500 ;
      RECT 2.9030 21.8565 2.9290 22.9500 ;
      RECT 2.7950 21.8565 2.8210 22.9500 ;
      RECT 2.6870 21.8565 2.7130 22.9500 ;
      RECT 2.5790 21.8565 2.6050 22.9500 ;
      RECT 2.4710 21.8565 2.4970 22.9500 ;
      RECT 2.3630 21.8565 2.3890 22.9500 ;
      RECT 2.2550 21.8565 2.2810 22.9500 ;
      RECT 2.1470 21.8565 2.1730 22.9500 ;
      RECT 2.0390 21.8565 2.0650 22.9500 ;
      RECT 1.9310 21.8565 1.9570 22.9500 ;
      RECT 1.8230 21.8565 1.8490 22.9500 ;
      RECT 1.7150 21.8565 1.7410 22.9500 ;
      RECT 1.6070 21.8565 1.6330 22.9500 ;
      RECT 1.4990 21.8565 1.5250 22.9500 ;
      RECT 1.3910 21.8565 1.4170 22.9500 ;
      RECT 1.2830 21.8565 1.3090 22.9500 ;
      RECT 1.1750 21.8565 1.2010 22.9500 ;
      RECT 1.0670 21.8565 1.0930 22.9500 ;
      RECT 0.9590 21.8565 0.9850 22.9500 ;
      RECT 0.8510 21.8565 0.8770 22.9500 ;
      RECT 0.7430 21.8565 0.7690 22.9500 ;
      RECT 0.6350 21.8565 0.6610 22.9500 ;
      RECT 0.5270 21.8565 0.5530 22.9500 ;
      RECT 0.4190 21.8565 0.4450 22.9500 ;
      RECT 0.3110 21.8565 0.3370 22.9500 ;
      RECT 0.2030 21.8565 0.2290 22.9500 ;
      RECT 0.0000 21.8565 0.0850 22.9500 ;
      RECT 5.1800 22.9365 5.3080 24.0300 ;
      RECT 5.1660 23.6020 5.3080 23.9245 ;
      RECT 5.0180 23.3290 5.0800 24.0300 ;
      RECT 5.0040 23.6385 5.0800 23.7920 ;
      RECT 5.0180 22.9365 5.0440 24.0300 ;
      RECT 5.0180 23.0575 5.0580 23.2970 ;
      RECT 5.0180 22.9365 5.0800 23.0255 ;
      RECT 4.7210 23.3870 4.9270 24.0300 ;
      RECT 4.9010 22.9365 4.9270 24.0300 ;
      RECT 4.7210 23.6640 4.9410 23.9220 ;
      RECT 4.7210 22.9365 4.8190 24.0300 ;
      RECT 4.3040 22.9365 4.3870 24.0300 ;
      RECT 4.3040 23.0250 4.4010 23.9605 ;
      RECT 9.5270 22.9365 9.6120 24.0300 ;
      RECT 9.3830 22.9365 9.4090 24.0300 ;
      RECT 9.2750 22.9365 9.3010 24.0300 ;
      RECT 9.1670 22.9365 9.1930 24.0300 ;
      RECT 9.0590 22.9365 9.0850 24.0300 ;
      RECT 8.9510 22.9365 8.9770 24.0300 ;
      RECT 8.8430 22.9365 8.8690 24.0300 ;
      RECT 8.7350 22.9365 8.7610 24.0300 ;
      RECT 8.6270 22.9365 8.6530 24.0300 ;
      RECT 8.5190 22.9365 8.5450 24.0300 ;
      RECT 8.4110 22.9365 8.4370 24.0300 ;
      RECT 8.3030 22.9365 8.3290 24.0300 ;
      RECT 8.1950 22.9365 8.2210 24.0300 ;
      RECT 8.0870 22.9365 8.1130 24.0300 ;
      RECT 7.9790 22.9365 8.0050 24.0300 ;
      RECT 7.8710 22.9365 7.8970 24.0300 ;
      RECT 7.7630 22.9365 7.7890 24.0300 ;
      RECT 7.6550 22.9365 7.6810 24.0300 ;
      RECT 7.5470 22.9365 7.5730 24.0300 ;
      RECT 7.4390 22.9365 7.4650 24.0300 ;
      RECT 7.3310 22.9365 7.3570 24.0300 ;
      RECT 7.2230 22.9365 7.2490 24.0300 ;
      RECT 7.1150 22.9365 7.1410 24.0300 ;
      RECT 7.0070 22.9365 7.0330 24.0300 ;
      RECT 6.8990 22.9365 6.9250 24.0300 ;
      RECT 6.7910 22.9365 6.8170 24.0300 ;
      RECT 6.6830 22.9365 6.7090 24.0300 ;
      RECT 6.5750 22.9365 6.6010 24.0300 ;
      RECT 6.4670 22.9365 6.4930 24.0300 ;
      RECT 6.3590 22.9365 6.3850 24.0300 ;
      RECT 6.2510 22.9365 6.2770 24.0300 ;
      RECT 6.1430 22.9365 6.1690 24.0300 ;
      RECT 6.0350 22.9365 6.0610 24.0300 ;
      RECT 5.9270 22.9365 5.9530 24.0300 ;
      RECT 5.7140 22.9365 5.7910 24.0300 ;
      RECT 3.8210 22.9365 3.8980 24.0300 ;
      RECT 3.6590 22.9365 3.6850 24.0300 ;
      RECT 3.5510 22.9365 3.5770 24.0300 ;
      RECT 3.4430 22.9365 3.4690 24.0300 ;
      RECT 3.3350 22.9365 3.3610 24.0300 ;
      RECT 3.2270 22.9365 3.2530 24.0300 ;
      RECT 3.1190 22.9365 3.1450 24.0300 ;
      RECT 3.0110 22.9365 3.0370 24.0300 ;
      RECT 2.9030 22.9365 2.9290 24.0300 ;
      RECT 2.7950 22.9365 2.8210 24.0300 ;
      RECT 2.6870 22.9365 2.7130 24.0300 ;
      RECT 2.5790 22.9365 2.6050 24.0300 ;
      RECT 2.4710 22.9365 2.4970 24.0300 ;
      RECT 2.3630 22.9365 2.3890 24.0300 ;
      RECT 2.2550 22.9365 2.2810 24.0300 ;
      RECT 2.1470 22.9365 2.1730 24.0300 ;
      RECT 2.0390 22.9365 2.0650 24.0300 ;
      RECT 1.9310 22.9365 1.9570 24.0300 ;
      RECT 1.8230 22.9365 1.8490 24.0300 ;
      RECT 1.7150 22.9365 1.7410 24.0300 ;
      RECT 1.6070 22.9365 1.6330 24.0300 ;
      RECT 1.4990 22.9365 1.5250 24.0300 ;
      RECT 1.3910 22.9365 1.4170 24.0300 ;
      RECT 1.2830 22.9365 1.3090 24.0300 ;
      RECT 1.1750 22.9365 1.2010 24.0300 ;
      RECT 1.0670 22.9365 1.0930 24.0300 ;
      RECT 0.9590 22.9365 0.9850 24.0300 ;
      RECT 0.8510 22.9365 0.8770 24.0300 ;
      RECT 0.7430 22.9365 0.7690 24.0300 ;
      RECT 0.6350 22.9365 0.6610 24.0300 ;
      RECT 0.5270 22.9365 0.5530 24.0300 ;
      RECT 0.4190 22.9365 0.4450 24.0300 ;
      RECT 0.3110 22.9365 0.3370 24.0300 ;
      RECT 0.2030 22.9365 0.2290 24.0300 ;
      RECT 0.0000 22.9365 0.0850 24.0300 ;
      RECT 5.1800 24.0165 5.3080 25.1100 ;
      RECT 5.1660 24.6820 5.3080 25.0045 ;
      RECT 5.0180 24.4090 5.0800 25.1100 ;
      RECT 5.0040 24.7185 5.0800 24.8720 ;
      RECT 5.0180 24.0165 5.0440 25.1100 ;
      RECT 5.0180 24.1375 5.0580 24.3770 ;
      RECT 5.0180 24.0165 5.0800 24.1055 ;
      RECT 4.7210 24.4670 4.9270 25.1100 ;
      RECT 4.9010 24.0165 4.9270 25.1100 ;
      RECT 4.7210 24.7440 4.9410 25.0020 ;
      RECT 4.7210 24.0165 4.8190 25.1100 ;
      RECT 4.3040 24.0165 4.3870 25.1100 ;
      RECT 4.3040 24.1050 4.4010 25.0405 ;
      RECT 9.5270 24.0165 9.6120 25.1100 ;
      RECT 9.3830 24.0165 9.4090 25.1100 ;
      RECT 9.2750 24.0165 9.3010 25.1100 ;
      RECT 9.1670 24.0165 9.1930 25.1100 ;
      RECT 9.0590 24.0165 9.0850 25.1100 ;
      RECT 8.9510 24.0165 8.9770 25.1100 ;
      RECT 8.8430 24.0165 8.8690 25.1100 ;
      RECT 8.7350 24.0165 8.7610 25.1100 ;
      RECT 8.6270 24.0165 8.6530 25.1100 ;
      RECT 8.5190 24.0165 8.5450 25.1100 ;
      RECT 8.4110 24.0165 8.4370 25.1100 ;
      RECT 8.3030 24.0165 8.3290 25.1100 ;
      RECT 8.1950 24.0165 8.2210 25.1100 ;
      RECT 8.0870 24.0165 8.1130 25.1100 ;
      RECT 7.9790 24.0165 8.0050 25.1100 ;
      RECT 7.8710 24.0165 7.8970 25.1100 ;
      RECT 7.7630 24.0165 7.7890 25.1100 ;
      RECT 7.6550 24.0165 7.6810 25.1100 ;
      RECT 7.5470 24.0165 7.5730 25.1100 ;
      RECT 7.4390 24.0165 7.4650 25.1100 ;
      RECT 7.3310 24.0165 7.3570 25.1100 ;
      RECT 7.2230 24.0165 7.2490 25.1100 ;
      RECT 7.1150 24.0165 7.1410 25.1100 ;
      RECT 7.0070 24.0165 7.0330 25.1100 ;
      RECT 6.8990 24.0165 6.9250 25.1100 ;
      RECT 6.7910 24.0165 6.8170 25.1100 ;
      RECT 6.6830 24.0165 6.7090 25.1100 ;
      RECT 6.5750 24.0165 6.6010 25.1100 ;
      RECT 6.4670 24.0165 6.4930 25.1100 ;
      RECT 6.3590 24.0165 6.3850 25.1100 ;
      RECT 6.2510 24.0165 6.2770 25.1100 ;
      RECT 6.1430 24.0165 6.1690 25.1100 ;
      RECT 6.0350 24.0165 6.0610 25.1100 ;
      RECT 5.9270 24.0165 5.9530 25.1100 ;
      RECT 5.7140 24.0165 5.7910 25.1100 ;
      RECT 3.8210 24.0165 3.8980 25.1100 ;
      RECT 3.6590 24.0165 3.6850 25.1100 ;
      RECT 3.5510 24.0165 3.5770 25.1100 ;
      RECT 3.4430 24.0165 3.4690 25.1100 ;
      RECT 3.3350 24.0165 3.3610 25.1100 ;
      RECT 3.2270 24.0165 3.2530 25.1100 ;
      RECT 3.1190 24.0165 3.1450 25.1100 ;
      RECT 3.0110 24.0165 3.0370 25.1100 ;
      RECT 2.9030 24.0165 2.9290 25.1100 ;
      RECT 2.7950 24.0165 2.8210 25.1100 ;
      RECT 2.6870 24.0165 2.7130 25.1100 ;
      RECT 2.5790 24.0165 2.6050 25.1100 ;
      RECT 2.4710 24.0165 2.4970 25.1100 ;
      RECT 2.3630 24.0165 2.3890 25.1100 ;
      RECT 2.2550 24.0165 2.2810 25.1100 ;
      RECT 2.1470 24.0165 2.1730 25.1100 ;
      RECT 2.0390 24.0165 2.0650 25.1100 ;
      RECT 1.9310 24.0165 1.9570 25.1100 ;
      RECT 1.8230 24.0165 1.8490 25.1100 ;
      RECT 1.7150 24.0165 1.7410 25.1100 ;
      RECT 1.6070 24.0165 1.6330 25.1100 ;
      RECT 1.4990 24.0165 1.5250 25.1100 ;
      RECT 1.3910 24.0165 1.4170 25.1100 ;
      RECT 1.2830 24.0165 1.3090 25.1100 ;
      RECT 1.1750 24.0165 1.2010 25.1100 ;
      RECT 1.0670 24.0165 1.0930 25.1100 ;
      RECT 0.9590 24.0165 0.9850 25.1100 ;
      RECT 0.8510 24.0165 0.8770 25.1100 ;
      RECT 0.7430 24.0165 0.7690 25.1100 ;
      RECT 0.6350 24.0165 0.6610 25.1100 ;
      RECT 0.5270 24.0165 0.5530 25.1100 ;
      RECT 0.4190 24.0165 0.4450 25.1100 ;
      RECT 0.3110 24.0165 0.3370 25.1100 ;
      RECT 0.2030 24.0165 0.2290 25.1100 ;
      RECT 0.0000 24.0165 0.0850 25.1100 ;
      RECT 5.1800 25.0965 5.3080 26.1900 ;
      RECT 5.1660 25.7620 5.3080 26.0845 ;
      RECT 5.0180 25.4890 5.0800 26.1900 ;
      RECT 5.0040 25.7985 5.0800 25.9520 ;
      RECT 5.0180 25.0965 5.0440 26.1900 ;
      RECT 5.0180 25.2175 5.0580 25.4570 ;
      RECT 5.0180 25.0965 5.0800 25.1855 ;
      RECT 4.7210 25.5470 4.9270 26.1900 ;
      RECT 4.9010 25.0965 4.9270 26.1900 ;
      RECT 4.7210 25.8240 4.9410 26.0820 ;
      RECT 4.7210 25.0965 4.8190 26.1900 ;
      RECT 4.3040 25.0965 4.3870 26.1900 ;
      RECT 4.3040 25.1850 4.4010 26.1205 ;
      RECT 9.5270 25.0965 9.6120 26.1900 ;
      RECT 9.3830 25.0965 9.4090 26.1900 ;
      RECT 9.2750 25.0965 9.3010 26.1900 ;
      RECT 9.1670 25.0965 9.1930 26.1900 ;
      RECT 9.0590 25.0965 9.0850 26.1900 ;
      RECT 8.9510 25.0965 8.9770 26.1900 ;
      RECT 8.8430 25.0965 8.8690 26.1900 ;
      RECT 8.7350 25.0965 8.7610 26.1900 ;
      RECT 8.6270 25.0965 8.6530 26.1900 ;
      RECT 8.5190 25.0965 8.5450 26.1900 ;
      RECT 8.4110 25.0965 8.4370 26.1900 ;
      RECT 8.3030 25.0965 8.3290 26.1900 ;
      RECT 8.1950 25.0965 8.2210 26.1900 ;
      RECT 8.0870 25.0965 8.1130 26.1900 ;
      RECT 7.9790 25.0965 8.0050 26.1900 ;
      RECT 7.8710 25.0965 7.8970 26.1900 ;
      RECT 7.7630 25.0965 7.7890 26.1900 ;
      RECT 7.6550 25.0965 7.6810 26.1900 ;
      RECT 7.5470 25.0965 7.5730 26.1900 ;
      RECT 7.4390 25.0965 7.4650 26.1900 ;
      RECT 7.3310 25.0965 7.3570 26.1900 ;
      RECT 7.2230 25.0965 7.2490 26.1900 ;
      RECT 7.1150 25.0965 7.1410 26.1900 ;
      RECT 7.0070 25.0965 7.0330 26.1900 ;
      RECT 6.8990 25.0965 6.9250 26.1900 ;
      RECT 6.7910 25.0965 6.8170 26.1900 ;
      RECT 6.6830 25.0965 6.7090 26.1900 ;
      RECT 6.5750 25.0965 6.6010 26.1900 ;
      RECT 6.4670 25.0965 6.4930 26.1900 ;
      RECT 6.3590 25.0965 6.3850 26.1900 ;
      RECT 6.2510 25.0965 6.2770 26.1900 ;
      RECT 6.1430 25.0965 6.1690 26.1900 ;
      RECT 6.0350 25.0965 6.0610 26.1900 ;
      RECT 5.9270 25.0965 5.9530 26.1900 ;
      RECT 5.7140 25.0965 5.7910 26.1900 ;
      RECT 3.8210 25.0965 3.8980 26.1900 ;
      RECT 3.6590 25.0965 3.6850 26.1900 ;
      RECT 3.5510 25.0965 3.5770 26.1900 ;
      RECT 3.4430 25.0965 3.4690 26.1900 ;
      RECT 3.3350 25.0965 3.3610 26.1900 ;
      RECT 3.2270 25.0965 3.2530 26.1900 ;
      RECT 3.1190 25.0965 3.1450 26.1900 ;
      RECT 3.0110 25.0965 3.0370 26.1900 ;
      RECT 2.9030 25.0965 2.9290 26.1900 ;
      RECT 2.7950 25.0965 2.8210 26.1900 ;
      RECT 2.6870 25.0965 2.7130 26.1900 ;
      RECT 2.5790 25.0965 2.6050 26.1900 ;
      RECT 2.4710 25.0965 2.4970 26.1900 ;
      RECT 2.3630 25.0965 2.3890 26.1900 ;
      RECT 2.2550 25.0965 2.2810 26.1900 ;
      RECT 2.1470 25.0965 2.1730 26.1900 ;
      RECT 2.0390 25.0965 2.0650 26.1900 ;
      RECT 1.9310 25.0965 1.9570 26.1900 ;
      RECT 1.8230 25.0965 1.8490 26.1900 ;
      RECT 1.7150 25.0965 1.7410 26.1900 ;
      RECT 1.6070 25.0965 1.6330 26.1900 ;
      RECT 1.4990 25.0965 1.5250 26.1900 ;
      RECT 1.3910 25.0965 1.4170 26.1900 ;
      RECT 1.2830 25.0965 1.3090 26.1900 ;
      RECT 1.1750 25.0965 1.2010 26.1900 ;
      RECT 1.0670 25.0965 1.0930 26.1900 ;
      RECT 0.9590 25.0965 0.9850 26.1900 ;
      RECT 0.8510 25.0965 0.8770 26.1900 ;
      RECT 0.7430 25.0965 0.7690 26.1900 ;
      RECT 0.6350 25.0965 0.6610 26.1900 ;
      RECT 0.5270 25.0965 0.5530 26.1900 ;
      RECT 0.4190 25.0965 0.4450 26.1900 ;
      RECT 0.3110 25.0965 0.3370 26.1900 ;
      RECT 0.2030 25.0965 0.2290 26.1900 ;
      RECT 0.0000 25.0965 0.0850 26.1900 ;
      RECT 5.1800 26.1765 5.3080 27.2700 ;
      RECT 5.1660 26.8420 5.3080 27.1645 ;
      RECT 5.0180 26.5690 5.0800 27.2700 ;
      RECT 5.0040 26.8785 5.0800 27.0320 ;
      RECT 5.0180 26.1765 5.0440 27.2700 ;
      RECT 5.0180 26.2975 5.0580 26.5370 ;
      RECT 5.0180 26.1765 5.0800 26.2655 ;
      RECT 4.7210 26.6270 4.9270 27.2700 ;
      RECT 4.9010 26.1765 4.9270 27.2700 ;
      RECT 4.7210 26.9040 4.9410 27.1620 ;
      RECT 4.7210 26.1765 4.8190 27.2700 ;
      RECT 4.3040 26.1765 4.3870 27.2700 ;
      RECT 4.3040 26.2650 4.4010 27.2005 ;
      RECT 9.5270 26.1765 9.6120 27.2700 ;
      RECT 9.3830 26.1765 9.4090 27.2700 ;
      RECT 9.2750 26.1765 9.3010 27.2700 ;
      RECT 9.1670 26.1765 9.1930 27.2700 ;
      RECT 9.0590 26.1765 9.0850 27.2700 ;
      RECT 8.9510 26.1765 8.9770 27.2700 ;
      RECT 8.8430 26.1765 8.8690 27.2700 ;
      RECT 8.7350 26.1765 8.7610 27.2700 ;
      RECT 8.6270 26.1765 8.6530 27.2700 ;
      RECT 8.5190 26.1765 8.5450 27.2700 ;
      RECT 8.4110 26.1765 8.4370 27.2700 ;
      RECT 8.3030 26.1765 8.3290 27.2700 ;
      RECT 8.1950 26.1765 8.2210 27.2700 ;
      RECT 8.0870 26.1765 8.1130 27.2700 ;
      RECT 7.9790 26.1765 8.0050 27.2700 ;
      RECT 7.8710 26.1765 7.8970 27.2700 ;
      RECT 7.7630 26.1765 7.7890 27.2700 ;
      RECT 7.6550 26.1765 7.6810 27.2700 ;
      RECT 7.5470 26.1765 7.5730 27.2700 ;
      RECT 7.4390 26.1765 7.4650 27.2700 ;
      RECT 7.3310 26.1765 7.3570 27.2700 ;
      RECT 7.2230 26.1765 7.2490 27.2700 ;
      RECT 7.1150 26.1765 7.1410 27.2700 ;
      RECT 7.0070 26.1765 7.0330 27.2700 ;
      RECT 6.8990 26.1765 6.9250 27.2700 ;
      RECT 6.7910 26.1765 6.8170 27.2700 ;
      RECT 6.6830 26.1765 6.7090 27.2700 ;
      RECT 6.5750 26.1765 6.6010 27.2700 ;
      RECT 6.4670 26.1765 6.4930 27.2700 ;
      RECT 6.3590 26.1765 6.3850 27.2700 ;
      RECT 6.2510 26.1765 6.2770 27.2700 ;
      RECT 6.1430 26.1765 6.1690 27.2700 ;
      RECT 6.0350 26.1765 6.0610 27.2700 ;
      RECT 5.9270 26.1765 5.9530 27.2700 ;
      RECT 5.7140 26.1765 5.7910 27.2700 ;
      RECT 3.8210 26.1765 3.8980 27.2700 ;
      RECT 3.6590 26.1765 3.6850 27.2700 ;
      RECT 3.5510 26.1765 3.5770 27.2700 ;
      RECT 3.4430 26.1765 3.4690 27.2700 ;
      RECT 3.3350 26.1765 3.3610 27.2700 ;
      RECT 3.2270 26.1765 3.2530 27.2700 ;
      RECT 3.1190 26.1765 3.1450 27.2700 ;
      RECT 3.0110 26.1765 3.0370 27.2700 ;
      RECT 2.9030 26.1765 2.9290 27.2700 ;
      RECT 2.7950 26.1765 2.8210 27.2700 ;
      RECT 2.6870 26.1765 2.7130 27.2700 ;
      RECT 2.5790 26.1765 2.6050 27.2700 ;
      RECT 2.4710 26.1765 2.4970 27.2700 ;
      RECT 2.3630 26.1765 2.3890 27.2700 ;
      RECT 2.2550 26.1765 2.2810 27.2700 ;
      RECT 2.1470 26.1765 2.1730 27.2700 ;
      RECT 2.0390 26.1765 2.0650 27.2700 ;
      RECT 1.9310 26.1765 1.9570 27.2700 ;
      RECT 1.8230 26.1765 1.8490 27.2700 ;
      RECT 1.7150 26.1765 1.7410 27.2700 ;
      RECT 1.6070 26.1765 1.6330 27.2700 ;
      RECT 1.4990 26.1765 1.5250 27.2700 ;
      RECT 1.3910 26.1765 1.4170 27.2700 ;
      RECT 1.2830 26.1765 1.3090 27.2700 ;
      RECT 1.1750 26.1765 1.2010 27.2700 ;
      RECT 1.0670 26.1765 1.0930 27.2700 ;
      RECT 0.9590 26.1765 0.9850 27.2700 ;
      RECT 0.8510 26.1765 0.8770 27.2700 ;
      RECT 0.7430 26.1765 0.7690 27.2700 ;
      RECT 0.6350 26.1765 0.6610 27.2700 ;
      RECT 0.5270 26.1765 0.5530 27.2700 ;
      RECT 0.4190 26.1765 0.4450 27.2700 ;
      RECT 0.3110 26.1765 0.3370 27.2700 ;
      RECT 0.2030 26.1765 0.2290 27.2700 ;
      RECT 0.0000 26.1765 0.0850 27.2700 ;
      RECT 5.1800 27.2565 5.3080 28.3500 ;
      RECT 5.1660 27.9220 5.3080 28.2445 ;
      RECT 5.0180 27.6490 5.0800 28.3500 ;
      RECT 5.0040 27.9585 5.0800 28.1120 ;
      RECT 5.0180 27.2565 5.0440 28.3500 ;
      RECT 5.0180 27.3775 5.0580 27.6170 ;
      RECT 5.0180 27.2565 5.0800 27.3455 ;
      RECT 4.7210 27.7070 4.9270 28.3500 ;
      RECT 4.9010 27.2565 4.9270 28.3500 ;
      RECT 4.7210 27.9840 4.9410 28.2420 ;
      RECT 4.7210 27.2565 4.8190 28.3500 ;
      RECT 4.3040 27.2565 4.3870 28.3500 ;
      RECT 4.3040 27.3450 4.4010 28.2805 ;
      RECT 9.5270 27.2565 9.6120 28.3500 ;
      RECT 9.3830 27.2565 9.4090 28.3500 ;
      RECT 9.2750 27.2565 9.3010 28.3500 ;
      RECT 9.1670 27.2565 9.1930 28.3500 ;
      RECT 9.0590 27.2565 9.0850 28.3500 ;
      RECT 8.9510 27.2565 8.9770 28.3500 ;
      RECT 8.8430 27.2565 8.8690 28.3500 ;
      RECT 8.7350 27.2565 8.7610 28.3500 ;
      RECT 8.6270 27.2565 8.6530 28.3500 ;
      RECT 8.5190 27.2565 8.5450 28.3500 ;
      RECT 8.4110 27.2565 8.4370 28.3500 ;
      RECT 8.3030 27.2565 8.3290 28.3500 ;
      RECT 8.1950 27.2565 8.2210 28.3500 ;
      RECT 8.0870 27.2565 8.1130 28.3500 ;
      RECT 7.9790 27.2565 8.0050 28.3500 ;
      RECT 7.8710 27.2565 7.8970 28.3500 ;
      RECT 7.7630 27.2565 7.7890 28.3500 ;
      RECT 7.6550 27.2565 7.6810 28.3500 ;
      RECT 7.5470 27.2565 7.5730 28.3500 ;
      RECT 7.4390 27.2565 7.4650 28.3500 ;
      RECT 7.3310 27.2565 7.3570 28.3500 ;
      RECT 7.2230 27.2565 7.2490 28.3500 ;
      RECT 7.1150 27.2565 7.1410 28.3500 ;
      RECT 7.0070 27.2565 7.0330 28.3500 ;
      RECT 6.8990 27.2565 6.9250 28.3500 ;
      RECT 6.7910 27.2565 6.8170 28.3500 ;
      RECT 6.6830 27.2565 6.7090 28.3500 ;
      RECT 6.5750 27.2565 6.6010 28.3500 ;
      RECT 6.4670 27.2565 6.4930 28.3500 ;
      RECT 6.3590 27.2565 6.3850 28.3500 ;
      RECT 6.2510 27.2565 6.2770 28.3500 ;
      RECT 6.1430 27.2565 6.1690 28.3500 ;
      RECT 6.0350 27.2565 6.0610 28.3500 ;
      RECT 5.9270 27.2565 5.9530 28.3500 ;
      RECT 5.7140 27.2565 5.7910 28.3500 ;
      RECT 3.8210 27.2565 3.8980 28.3500 ;
      RECT 3.6590 27.2565 3.6850 28.3500 ;
      RECT 3.5510 27.2565 3.5770 28.3500 ;
      RECT 3.4430 27.2565 3.4690 28.3500 ;
      RECT 3.3350 27.2565 3.3610 28.3500 ;
      RECT 3.2270 27.2565 3.2530 28.3500 ;
      RECT 3.1190 27.2565 3.1450 28.3500 ;
      RECT 3.0110 27.2565 3.0370 28.3500 ;
      RECT 2.9030 27.2565 2.9290 28.3500 ;
      RECT 2.7950 27.2565 2.8210 28.3500 ;
      RECT 2.6870 27.2565 2.7130 28.3500 ;
      RECT 2.5790 27.2565 2.6050 28.3500 ;
      RECT 2.4710 27.2565 2.4970 28.3500 ;
      RECT 2.3630 27.2565 2.3890 28.3500 ;
      RECT 2.2550 27.2565 2.2810 28.3500 ;
      RECT 2.1470 27.2565 2.1730 28.3500 ;
      RECT 2.0390 27.2565 2.0650 28.3500 ;
      RECT 1.9310 27.2565 1.9570 28.3500 ;
      RECT 1.8230 27.2565 1.8490 28.3500 ;
      RECT 1.7150 27.2565 1.7410 28.3500 ;
      RECT 1.6070 27.2565 1.6330 28.3500 ;
      RECT 1.4990 27.2565 1.5250 28.3500 ;
      RECT 1.3910 27.2565 1.4170 28.3500 ;
      RECT 1.2830 27.2565 1.3090 28.3500 ;
      RECT 1.1750 27.2565 1.2010 28.3500 ;
      RECT 1.0670 27.2565 1.0930 28.3500 ;
      RECT 0.9590 27.2565 0.9850 28.3500 ;
      RECT 0.8510 27.2565 0.8770 28.3500 ;
      RECT 0.7430 27.2565 0.7690 28.3500 ;
      RECT 0.6350 27.2565 0.6610 28.3500 ;
      RECT 0.5270 27.2565 0.5530 28.3500 ;
      RECT 0.4190 27.2565 0.4450 28.3500 ;
      RECT 0.3110 27.2565 0.3370 28.3500 ;
      RECT 0.2030 27.2565 0.2290 28.3500 ;
      RECT 0.0000 27.2565 0.0850 28.3500 ;
      RECT 5.1800 28.3365 5.3080 29.4300 ;
      RECT 5.1660 29.0020 5.3080 29.3245 ;
      RECT 5.0180 28.7290 5.0800 29.4300 ;
      RECT 5.0040 29.0385 5.0800 29.1920 ;
      RECT 5.0180 28.3365 5.0440 29.4300 ;
      RECT 5.0180 28.4575 5.0580 28.6970 ;
      RECT 5.0180 28.3365 5.0800 28.4255 ;
      RECT 4.7210 28.7870 4.9270 29.4300 ;
      RECT 4.9010 28.3365 4.9270 29.4300 ;
      RECT 4.7210 29.0640 4.9410 29.3220 ;
      RECT 4.7210 28.3365 4.8190 29.4300 ;
      RECT 4.3040 28.3365 4.3870 29.4300 ;
      RECT 4.3040 28.4250 4.4010 29.3605 ;
      RECT 9.5270 28.3365 9.6120 29.4300 ;
      RECT 9.3830 28.3365 9.4090 29.4300 ;
      RECT 9.2750 28.3365 9.3010 29.4300 ;
      RECT 9.1670 28.3365 9.1930 29.4300 ;
      RECT 9.0590 28.3365 9.0850 29.4300 ;
      RECT 8.9510 28.3365 8.9770 29.4300 ;
      RECT 8.8430 28.3365 8.8690 29.4300 ;
      RECT 8.7350 28.3365 8.7610 29.4300 ;
      RECT 8.6270 28.3365 8.6530 29.4300 ;
      RECT 8.5190 28.3365 8.5450 29.4300 ;
      RECT 8.4110 28.3365 8.4370 29.4300 ;
      RECT 8.3030 28.3365 8.3290 29.4300 ;
      RECT 8.1950 28.3365 8.2210 29.4300 ;
      RECT 8.0870 28.3365 8.1130 29.4300 ;
      RECT 7.9790 28.3365 8.0050 29.4300 ;
      RECT 7.8710 28.3365 7.8970 29.4300 ;
      RECT 7.7630 28.3365 7.7890 29.4300 ;
      RECT 7.6550 28.3365 7.6810 29.4300 ;
      RECT 7.5470 28.3365 7.5730 29.4300 ;
      RECT 7.4390 28.3365 7.4650 29.4300 ;
      RECT 7.3310 28.3365 7.3570 29.4300 ;
      RECT 7.2230 28.3365 7.2490 29.4300 ;
      RECT 7.1150 28.3365 7.1410 29.4300 ;
      RECT 7.0070 28.3365 7.0330 29.4300 ;
      RECT 6.8990 28.3365 6.9250 29.4300 ;
      RECT 6.7910 28.3365 6.8170 29.4300 ;
      RECT 6.6830 28.3365 6.7090 29.4300 ;
      RECT 6.5750 28.3365 6.6010 29.4300 ;
      RECT 6.4670 28.3365 6.4930 29.4300 ;
      RECT 6.3590 28.3365 6.3850 29.4300 ;
      RECT 6.2510 28.3365 6.2770 29.4300 ;
      RECT 6.1430 28.3365 6.1690 29.4300 ;
      RECT 6.0350 28.3365 6.0610 29.4300 ;
      RECT 5.9270 28.3365 5.9530 29.4300 ;
      RECT 5.7140 28.3365 5.7910 29.4300 ;
      RECT 3.8210 28.3365 3.8980 29.4300 ;
      RECT 3.6590 28.3365 3.6850 29.4300 ;
      RECT 3.5510 28.3365 3.5770 29.4300 ;
      RECT 3.4430 28.3365 3.4690 29.4300 ;
      RECT 3.3350 28.3365 3.3610 29.4300 ;
      RECT 3.2270 28.3365 3.2530 29.4300 ;
      RECT 3.1190 28.3365 3.1450 29.4300 ;
      RECT 3.0110 28.3365 3.0370 29.4300 ;
      RECT 2.9030 28.3365 2.9290 29.4300 ;
      RECT 2.7950 28.3365 2.8210 29.4300 ;
      RECT 2.6870 28.3365 2.7130 29.4300 ;
      RECT 2.5790 28.3365 2.6050 29.4300 ;
      RECT 2.4710 28.3365 2.4970 29.4300 ;
      RECT 2.3630 28.3365 2.3890 29.4300 ;
      RECT 2.2550 28.3365 2.2810 29.4300 ;
      RECT 2.1470 28.3365 2.1730 29.4300 ;
      RECT 2.0390 28.3365 2.0650 29.4300 ;
      RECT 1.9310 28.3365 1.9570 29.4300 ;
      RECT 1.8230 28.3365 1.8490 29.4300 ;
      RECT 1.7150 28.3365 1.7410 29.4300 ;
      RECT 1.6070 28.3365 1.6330 29.4300 ;
      RECT 1.4990 28.3365 1.5250 29.4300 ;
      RECT 1.3910 28.3365 1.4170 29.4300 ;
      RECT 1.2830 28.3365 1.3090 29.4300 ;
      RECT 1.1750 28.3365 1.2010 29.4300 ;
      RECT 1.0670 28.3365 1.0930 29.4300 ;
      RECT 0.9590 28.3365 0.9850 29.4300 ;
      RECT 0.8510 28.3365 0.8770 29.4300 ;
      RECT 0.7430 28.3365 0.7690 29.4300 ;
      RECT 0.6350 28.3365 0.6610 29.4300 ;
      RECT 0.5270 28.3365 0.5530 29.4300 ;
      RECT 0.4190 28.3365 0.4450 29.4300 ;
      RECT 0.3110 28.3365 0.3370 29.4300 ;
      RECT 0.2030 28.3365 0.2290 29.4300 ;
      RECT 0.0000 28.3365 0.0850 29.4300 ;
      RECT 5.1800 29.4165 5.3080 30.5100 ;
      RECT 5.1660 30.0820 5.3080 30.4045 ;
      RECT 5.0180 29.8090 5.0800 30.5100 ;
      RECT 5.0040 30.1185 5.0800 30.2720 ;
      RECT 5.0180 29.4165 5.0440 30.5100 ;
      RECT 5.0180 29.5375 5.0580 29.7770 ;
      RECT 5.0180 29.4165 5.0800 29.5055 ;
      RECT 4.7210 29.8670 4.9270 30.5100 ;
      RECT 4.9010 29.4165 4.9270 30.5100 ;
      RECT 4.7210 30.1440 4.9410 30.4020 ;
      RECT 4.7210 29.4165 4.8190 30.5100 ;
      RECT 4.3040 29.4165 4.3870 30.5100 ;
      RECT 4.3040 29.5050 4.4010 30.4405 ;
      RECT 9.5270 29.4165 9.6120 30.5100 ;
      RECT 9.3830 29.4165 9.4090 30.5100 ;
      RECT 9.2750 29.4165 9.3010 30.5100 ;
      RECT 9.1670 29.4165 9.1930 30.5100 ;
      RECT 9.0590 29.4165 9.0850 30.5100 ;
      RECT 8.9510 29.4165 8.9770 30.5100 ;
      RECT 8.8430 29.4165 8.8690 30.5100 ;
      RECT 8.7350 29.4165 8.7610 30.5100 ;
      RECT 8.6270 29.4165 8.6530 30.5100 ;
      RECT 8.5190 29.4165 8.5450 30.5100 ;
      RECT 8.4110 29.4165 8.4370 30.5100 ;
      RECT 8.3030 29.4165 8.3290 30.5100 ;
      RECT 8.1950 29.4165 8.2210 30.5100 ;
      RECT 8.0870 29.4165 8.1130 30.5100 ;
      RECT 7.9790 29.4165 8.0050 30.5100 ;
      RECT 7.8710 29.4165 7.8970 30.5100 ;
      RECT 7.7630 29.4165 7.7890 30.5100 ;
      RECT 7.6550 29.4165 7.6810 30.5100 ;
      RECT 7.5470 29.4165 7.5730 30.5100 ;
      RECT 7.4390 29.4165 7.4650 30.5100 ;
      RECT 7.3310 29.4165 7.3570 30.5100 ;
      RECT 7.2230 29.4165 7.2490 30.5100 ;
      RECT 7.1150 29.4165 7.1410 30.5100 ;
      RECT 7.0070 29.4165 7.0330 30.5100 ;
      RECT 6.8990 29.4165 6.9250 30.5100 ;
      RECT 6.7910 29.4165 6.8170 30.5100 ;
      RECT 6.6830 29.4165 6.7090 30.5100 ;
      RECT 6.5750 29.4165 6.6010 30.5100 ;
      RECT 6.4670 29.4165 6.4930 30.5100 ;
      RECT 6.3590 29.4165 6.3850 30.5100 ;
      RECT 6.2510 29.4165 6.2770 30.5100 ;
      RECT 6.1430 29.4165 6.1690 30.5100 ;
      RECT 6.0350 29.4165 6.0610 30.5100 ;
      RECT 5.9270 29.4165 5.9530 30.5100 ;
      RECT 5.7140 29.4165 5.7910 30.5100 ;
      RECT 3.8210 29.4165 3.8980 30.5100 ;
      RECT 3.6590 29.4165 3.6850 30.5100 ;
      RECT 3.5510 29.4165 3.5770 30.5100 ;
      RECT 3.4430 29.4165 3.4690 30.5100 ;
      RECT 3.3350 29.4165 3.3610 30.5100 ;
      RECT 3.2270 29.4165 3.2530 30.5100 ;
      RECT 3.1190 29.4165 3.1450 30.5100 ;
      RECT 3.0110 29.4165 3.0370 30.5100 ;
      RECT 2.9030 29.4165 2.9290 30.5100 ;
      RECT 2.7950 29.4165 2.8210 30.5100 ;
      RECT 2.6870 29.4165 2.7130 30.5100 ;
      RECT 2.5790 29.4165 2.6050 30.5100 ;
      RECT 2.4710 29.4165 2.4970 30.5100 ;
      RECT 2.3630 29.4165 2.3890 30.5100 ;
      RECT 2.2550 29.4165 2.2810 30.5100 ;
      RECT 2.1470 29.4165 2.1730 30.5100 ;
      RECT 2.0390 29.4165 2.0650 30.5100 ;
      RECT 1.9310 29.4165 1.9570 30.5100 ;
      RECT 1.8230 29.4165 1.8490 30.5100 ;
      RECT 1.7150 29.4165 1.7410 30.5100 ;
      RECT 1.6070 29.4165 1.6330 30.5100 ;
      RECT 1.4990 29.4165 1.5250 30.5100 ;
      RECT 1.3910 29.4165 1.4170 30.5100 ;
      RECT 1.2830 29.4165 1.3090 30.5100 ;
      RECT 1.1750 29.4165 1.2010 30.5100 ;
      RECT 1.0670 29.4165 1.0930 30.5100 ;
      RECT 0.9590 29.4165 0.9850 30.5100 ;
      RECT 0.8510 29.4165 0.8770 30.5100 ;
      RECT 0.7430 29.4165 0.7690 30.5100 ;
      RECT 0.6350 29.4165 0.6610 30.5100 ;
      RECT 0.5270 29.4165 0.5530 30.5100 ;
      RECT 0.4190 29.4165 0.4450 30.5100 ;
      RECT 0.3110 29.4165 0.3370 30.5100 ;
      RECT 0.2030 29.4165 0.2290 30.5100 ;
      RECT 0.0000 29.4165 0.0850 30.5100 ;
      RECT 5.1800 30.4965 5.3080 31.5900 ;
      RECT 5.1660 31.1620 5.3080 31.4845 ;
      RECT 5.0180 30.8890 5.0800 31.5900 ;
      RECT 5.0040 31.1985 5.0800 31.3520 ;
      RECT 5.0180 30.4965 5.0440 31.5900 ;
      RECT 5.0180 30.6175 5.0580 30.8570 ;
      RECT 5.0180 30.4965 5.0800 30.5855 ;
      RECT 4.7210 30.9470 4.9270 31.5900 ;
      RECT 4.9010 30.4965 4.9270 31.5900 ;
      RECT 4.7210 31.2240 4.9410 31.4820 ;
      RECT 4.7210 30.4965 4.8190 31.5900 ;
      RECT 4.3040 30.4965 4.3870 31.5900 ;
      RECT 4.3040 30.5850 4.4010 31.5205 ;
      RECT 9.5270 30.4965 9.6120 31.5900 ;
      RECT 9.3830 30.4965 9.4090 31.5900 ;
      RECT 9.2750 30.4965 9.3010 31.5900 ;
      RECT 9.1670 30.4965 9.1930 31.5900 ;
      RECT 9.0590 30.4965 9.0850 31.5900 ;
      RECT 8.9510 30.4965 8.9770 31.5900 ;
      RECT 8.8430 30.4965 8.8690 31.5900 ;
      RECT 8.7350 30.4965 8.7610 31.5900 ;
      RECT 8.6270 30.4965 8.6530 31.5900 ;
      RECT 8.5190 30.4965 8.5450 31.5900 ;
      RECT 8.4110 30.4965 8.4370 31.5900 ;
      RECT 8.3030 30.4965 8.3290 31.5900 ;
      RECT 8.1950 30.4965 8.2210 31.5900 ;
      RECT 8.0870 30.4965 8.1130 31.5900 ;
      RECT 7.9790 30.4965 8.0050 31.5900 ;
      RECT 7.8710 30.4965 7.8970 31.5900 ;
      RECT 7.7630 30.4965 7.7890 31.5900 ;
      RECT 7.6550 30.4965 7.6810 31.5900 ;
      RECT 7.5470 30.4965 7.5730 31.5900 ;
      RECT 7.4390 30.4965 7.4650 31.5900 ;
      RECT 7.3310 30.4965 7.3570 31.5900 ;
      RECT 7.2230 30.4965 7.2490 31.5900 ;
      RECT 7.1150 30.4965 7.1410 31.5900 ;
      RECT 7.0070 30.4965 7.0330 31.5900 ;
      RECT 6.8990 30.4965 6.9250 31.5900 ;
      RECT 6.7910 30.4965 6.8170 31.5900 ;
      RECT 6.6830 30.4965 6.7090 31.5900 ;
      RECT 6.5750 30.4965 6.6010 31.5900 ;
      RECT 6.4670 30.4965 6.4930 31.5900 ;
      RECT 6.3590 30.4965 6.3850 31.5900 ;
      RECT 6.2510 30.4965 6.2770 31.5900 ;
      RECT 6.1430 30.4965 6.1690 31.5900 ;
      RECT 6.0350 30.4965 6.0610 31.5900 ;
      RECT 5.9270 30.4965 5.9530 31.5900 ;
      RECT 5.7140 30.4965 5.7910 31.5900 ;
      RECT 3.8210 30.4965 3.8980 31.5900 ;
      RECT 3.6590 30.4965 3.6850 31.5900 ;
      RECT 3.5510 30.4965 3.5770 31.5900 ;
      RECT 3.4430 30.4965 3.4690 31.5900 ;
      RECT 3.3350 30.4965 3.3610 31.5900 ;
      RECT 3.2270 30.4965 3.2530 31.5900 ;
      RECT 3.1190 30.4965 3.1450 31.5900 ;
      RECT 3.0110 30.4965 3.0370 31.5900 ;
      RECT 2.9030 30.4965 2.9290 31.5900 ;
      RECT 2.7950 30.4965 2.8210 31.5900 ;
      RECT 2.6870 30.4965 2.7130 31.5900 ;
      RECT 2.5790 30.4965 2.6050 31.5900 ;
      RECT 2.4710 30.4965 2.4970 31.5900 ;
      RECT 2.3630 30.4965 2.3890 31.5900 ;
      RECT 2.2550 30.4965 2.2810 31.5900 ;
      RECT 2.1470 30.4965 2.1730 31.5900 ;
      RECT 2.0390 30.4965 2.0650 31.5900 ;
      RECT 1.9310 30.4965 1.9570 31.5900 ;
      RECT 1.8230 30.4965 1.8490 31.5900 ;
      RECT 1.7150 30.4965 1.7410 31.5900 ;
      RECT 1.6070 30.4965 1.6330 31.5900 ;
      RECT 1.4990 30.4965 1.5250 31.5900 ;
      RECT 1.3910 30.4965 1.4170 31.5900 ;
      RECT 1.2830 30.4965 1.3090 31.5900 ;
      RECT 1.1750 30.4965 1.2010 31.5900 ;
      RECT 1.0670 30.4965 1.0930 31.5900 ;
      RECT 0.9590 30.4965 0.9850 31.5900 ;
      RECT 0.8510 30.4965 0.8770 31.5900 ;
      RECT 0.7430 30.4965 0.7690 31.5900 ;
      RECT 0.6350 30.4965 0.6610 31.5900 ;
      RECT 0.5270 30.4965 0.5530 31.5900 ;
      RECT 0.4190 30.4965 0.4450 31.5900 ;
      RECT 0.3110 30.4965 0.3370 31.5900 ;
      RECT 0.2030 30.4965 0.2290 31.5900 ;
      RECT 0.0000 30.4965 0.0850 31.5900 ;
      RECT 5.1800 31.5765 5.3080 32.6700 ;
      RECT 5.1660 32.2420 5.3080 32.5645 ;
      RECT 5.0180 31.9690 5.0800 32.6700 ;
      RECT 5.0040 32.2785 5.0800 32.4320 ;
      RECT 5.0180 31.5765 5.0440 32.6700 ;
      RECT 5.0180 31.6975 5.0580 31.9370 ;
      RECT 5.0180 31.5765 5.0800 31.6655 ;
      RECT 4.7210 32.0270 4.9270 32.6700 ;
      RECT 4.9010 31.5765 4.9270 32.6700 ;
      RECT 4.7210 32.3040 4.9410 32.5620 ;
      RECT 4.7210 31.5765 4.8190 32.6700 ;
      RECT 4.3040 31.5765 4.3870 32.6700 ;
      RECT 4.3040 31.6650 4.4010 32.6005 ;
      RECT 9.5270 31.5765 9.6120 32.6700 ;
      RECT 9.3830 31.5765 9.4090 32.6700 ;
      RECT 9.2750 31.5765 9.3010 32.6700 ;
      RECT 9.1670 31.5765 9.1930 32.6700 ;
      RECT 9.0590 31.5765 9.0850 32.6700 ;
      RECT 8.9510 31.5765 8.9770 32.6700 ;
      RECT 8.8430 31.5765 8.8690 32.6700 ;
      RECT 8.7350 31.5765 8.7610 32.6700 ;
      RECT 8.6270 31.5765 8.6530 32.6700 ;
      RECT 8.5190 31.5765 8.5450 32.6700 ;
      RECT 8.4110 31.5765 8.4370 32.6700 ;
      RECT 8.3030 31.5765 8.3290 32.6700 ;
      RECT 8.1950 31.5765 8.2210 32.6700 ;
      RECT 8.0870 31.5765 8.1130 32.6700 ;
      RECT 7.9790 31.5765 8.0050 32.6700 ;
      RECT 7.8710 31.5765 7.8970 32.6700 ;
      RECT 7.7630 31.5765 7.7890 32.6700 ;
      RECT 7.6550 31.5765 7.6810 32.6700 ;
      RECT 7.5470 31.5765 7.5730 32.6700 ;
      RECT 7.4390 31.5765 7.4650 32.6700 ;
      RECT 7.3310 31.5765 7.3570 32.6700 ;
      RECT 7.2230 31.5765 7.2490 32.6700 ;
      RECT 7.1150 31.5765 7.1410 32.6700 ;
      RECT 7.0070 31.5765 7.0330 32.6700 ;
      RECT 6.8990 31.5765 6.9250 32.6700 ;
      RECT 6.7910 31.5765 6.8170 32.6700 ;
      RECT 6.6830 31.5765 6.7090 32.6700 ;
      RECT 6.5750 31.5765 6.6010 32.6700 ;
      RECT 6.4670 31.5765 6.4930 32.6700 ;
      RECT 6.3590 31.5765 6.3850 32.6700 ;
      RECT 6.2510 31.5765 6.2770 32.6700 ;
      RECT 6.1430 31.5765 6.1690 32.6700 ;
      RECT 6.0350 31.5765 6.0610 32.6700 ;
      RECT 5.9270 31.5765 5.9530 32.6700 ;
      RECT 5.7140 31.5765 5.7910 32.6700 ;
      RECT 3.8210 31.5765 3.8980 32.6700 ;
      RECT 3.6590 31.5765 3.6850 32.6700 ;
      RECT 3.5510 31.5765 3.5770 32.6700 ;
      RECT 3.4430 31.5765 3.4690 32.6700 ;
      RECT 3.3350 31.5765 3.3610 32.6700 ;
      RECT 3.2270 31.5765 3.2530 32.6700 ;
      RECT 3.1190 31.5765 3.1450 32.6700 ;
      RECT 3.0110 31.5765 3.0370 32.6700 ;
      RECT 2.9030 31.5765 2.9290 32.6700 ;
      RECT 2.7950 31.5765 2.8210 32.6700 ;
      RECT 2.6870 31.5765 2.7130 32.6700 ;
      RECT 2.5790 31.5765 2.6050 32.6700 ;
      RECT 2.4710 31.5765 2.4970 32.6700 ;
      RECT 2.3630 31.5765 2.3890 32.6700 ;
      RECT 2.2550 31.5765 2.2810 32.6700 ;
      RECT 2.1470 31.5765 2.1730 32.6700 ;
      RECT 2.0390 31.5765 2.0650 32.6700 ;
      RECT 1.9310 31.5765 1.9570 32.6700 ;
      RECT 1.8230 31.5765 1.8490 32.6700 ;
      RECT 1.7150 31.5765 1.7410 32.6700 ;
      RECT 1.6070 31.5765 1.6330 32.6700 ;
      RECT 1.4990 31.5765 1.5250 32.6700 ;
      RECT 1.3910 31.5765 1.4170 32.6700 ;
      RECT 1.2830 31.5765 1.3090 32.6700 ;
      RECT 1.1750 31.5765 1.2010 32.6700 ;
      RECT 1.0670 31.5765 1.0930 32.6700 ;
      RECT 0.9590 31.5765 0.9850 32.6700 ;
      RECT 0.8510 31.5765 0.8770 32.6700 ;
      RECT 0.7430 31.5765 0.7690 32.6700 ;
      RECT 0.6350 31.5765 0.6610 32.6700 ;
      RECT 0.5270 31.5765 0.5530 32.6700 ;
      RECT 0.4190 31.5765 0.4450 32.6700 ;
      RECT 0.3110 31.5765 0.3370 32.6700 ;
      RECT 0.2030 31.5765 0.2290 32.6700 ;
      RECT 0.0000 31.5765 0.0850 32.6700 ;
      RECT 5.1800 32.6565 5.3080 33.7500 ;
      RECT 5.1660 33.3220 5.3080 33.6445 ;
      RECT 5.0180 33.0490 5.0800 33.7500 ;
      RECT 5.0040 33.3585 5.0800 33.5120 ;
      RECT 5.0180 32.6565 5.0440 33.7500 ;
      RECT 5.0180 32.7775 5.0580 33.0170 ;
      RECT 5.0180 32.6565 5.0800 32.7455 ;
      RECT 4.7210 33.1070 4.9270 33.7500 ;
      RECT 4.9010 32.6565 4.9270 33.7500 ;
      RECT 4.7210 33.3840 4.9410 33.6420 ;
      RECT 4.7210 32.6565 4.8190 33.7500 ;
      RECT 4.3040 32.6565 4.3870 33.7500 ;
      RECT 4.3040 32.7450 4.4010 33.6805 ;
      RECT 9.5270 32.6565 9.6120 33.7500 ;
      RECT 9.3830 32.6565 9.4090 33.7500 ;
      RECT 9.2750 32.6565 9.3010 33.7500 ;
      RECT 9.1670 32.6565 9.1930 33.7500 ;
      RECT 9.0590 32.6565 9.0850 33.7500 ;
      RECT 8.9510 32.6565 8.9770 33.7500 ;
      RECT 8.8430 32.6565 8.8690 33.7500 ;
      RECT 8.7350 32.6565 8.7610 33.7500 ;
      RECT 8.6270 32.6565 8.6530 33.7500 ;
      RECT 8.5190 32.6565 8.5450 33.7500 ;
      RECT 8.4110 32.6565 8.4370 33.7500 ;
      RECT 8.3030 32.6565 8.3290 33.7500 ;
      RECT 8.1950 32.6565 8.2210 33.7500 ;
      RECT 8.0870 32.6565 8.1130 33.7500 ;
      RECT 7.9790 32.6565 8.0050 33.7500 ;
      RECT 7.8710 32.6565 7.8970 33.7500 ;
      RECT 7.7630 32.6565 7.7890 33.7500 ;
      RECT 7.6550 32.6565 7.6810 33.7500 ;
      RECT 7.5470 32.6565 7.5730 33.7500 ;
      RECT 7.4390 32.6565 7.4650 33.7500 ;
      RECT 7.3310 32.6565 7.3570 33.7500 ;
      RECT 7.2230 32.6565 7.2490 33.7500 ;
      RECT 7.1150 32.6565 7.1410 33.7500 ;
      RECT 7.0070 32.6565 7.0330 33.7500 ;
      RECT 6.8990 32.6565 6.9250 33.7500 ;
      RECT 6.7910 32.6565 6.8170 33.7500 ;
      RECT 6.6830 32.6565 6.7090 33.7500 ;
      RECT 6.5750 32.6565 6.6010 33.7500 ;
      RECT 6.4670 32.6565 6.4930 33.7500 ;
      RECT 6.3590 32.6565 6.3850 33.7500 ;
      RECT 6.2510 32.6565 6.2770 33.7500 ;
      RECT 6.1430 32.6565 6.1690 33.7500 ;
      RECT 6.0350 32.6565 6.0610 33.7500 ;
      RECT 5.9270 32.6565 5.9530 33.7500 ;
      RECT 5.7140 32.6565 5.7910 33.7500 ;
      RECT 3.8210 32.6565 3.8980 33.7500 ;
      RECT 3.6590 32.6565 3.6850 33.7500 ;
      RECT 3.5510 32.6565 3.5770 33.7500 ;
      RECT 3.4430 32.6565 3.4690 33.7500 ;
      RECT 3.3350 32.6565 3.3610 33.7500 ;
      RECT 3.2270 32.6565 3.2530 33.7500 ;
      RECT 3.1190 32.6565 3.1450 33.7500 ;
      RECT 3.0110 32.6565 3.0370 33.7500 ;
      RECT 2.9030 32.6565 2.9290 33.7500 ;
      RECT 2.7950 32.6565 2.8210 33.7500 ;
      RECT 2.6870 32.6565 2.7130 33.7500 ;
      RECT 2.5790 32.6565 2.6050 33.7500 ;
      RECT 2.4710 32.6565 2.4970 33.7500 ;
      RECT 2.3630 32.6565 2.3890 33.7500 ;
      RECT 2.2550 32.6565 2.2810 33.7500 ;
      RECT 2.1470 32.6565 2.1730 33.7500 ;
      RECT 2.0390 32.6565 2.0650 33.7500 ;
      RECT 1.9310 32.6565 1.9570 33.7500 ;
      RECT 1.8230 32.6565 1.8490 33.7500 ;
      RECT 1.7150 32.6565 1.7410 33.7500 ;
      RECT 1.6070 32.6565 1.6330 33.7500 ;
      RECT 1.4990 32.6565 1.5250 33.7500 ;
      RECT 1.3910 32.6565 1.4170 33.7500 ;
      RECT 1.2830 32.6565 1.3090 33.7500 ;
      RECT 1.1750 32.6565 1.2010 33.7500 ;
      RECT 1.0670 32.6565 1.0930 33.7500 ;
      RECT 0.9590 32.6565 0.9850 33.7500 ;
      RECT 0.8510 32.6565 0.8770 33.7500 ;
      RECT 0.7430 32.6565 0.7690 33.7500 ;
      RECT 0.6350 32.6565 0.6610 33.7500 ;
      RECT 0.5270 32.6565 0.5530 33.7500 ;
      RECT 0.4190 32.6565 0.4450 33.7500 ;
      RECT 0.3110 32.6565 0.3370 33.7500 ;
      RECT 0.2030 32.6565 0.2290 33.7500 ;
      RECT 0.0000 32.6565 0.0850 33.7500 ;
      RECT 5.1800 33.7365 5.3080 34.8300 ;
      RECT 5.1660 34.4020 5.3080 34.7245 ;
      RECT 5.0180 34.1290 5.0800 34.8300 ;
      RECT 5.0040 34.4385 5.0800 34.5920 ;
      RECT 5.0180 33.7365 5.0440 34.8300 ;
      RECT 5.0180 33.8575 5.0580 34.0970 ;
      RECT 5.0180 33.7365 5.0800 33.8255 ;
      RECT 4.7210 34.1870 4.9270 34.8300 ;
      RECT 4.9010 33.7365 4.9270 34.8300 ;
      RECT 4.7210 34.4640 4.9410 34.7220 ;
      RECT 4.7210 33.7365 4.8190 34.8300 ;
      RECT 4.3040 33.7365 4.3870 34.8300 ;
      RECT 4.3040 33.8250 4.4010 34.7605 ;
      RECT 9.5270 33.7365 9.6120 34.8300 ;
      RECT 9.3830 33.7365 9.4090 34.8300 ;
      RECT 9.2750 33.7365 9.3010 34.8300 ;
      RECT 9.1670 33.7365 9.1930 34.8300 ;
      RECT 9.0590 33.7365 9.0850 34.8300 ;
      RECT 8.9510 33.7365 8.9770 34.8300 ;
      RECT 8.8430 33.7365 8.8690 34.8300 ;
      RECT 8.7350 33.7365 8.7610 34.8300 ;
      RECT 8.6270 33.7365 8.6530 34.8300 ;
      RECT 8.5190 33.7365 8.5450 34.8300 ;
      RECT 8.4110 33.7365 8.4370 34.8300 ;
      RECT 8.3030 33.7365 8.3290 34.8300 ;
      RECT 8.1950 33.7365 8.2210 34.8300 ;
      RECT 8.0870 33.7365 8.1130 34.8300 ;
      RECT 7.9790 33.7365 8.0050 34.8300 ;
      RECT 7.8710 33.7365 7.8970 34.8300 ;
      RECT 7.7630 33.7365 7.7890 34.8300 ;
      RECT 7.6550 33.7365 7.6810 34.8300 ;
      RECT 7.5470 33.7365 7.5730 34.8300 ;
      RECT 7.4390 33.7365 7.4650 34.8300 ;
      RECT 7.3310 33.7365 7.3570 34.8300 ;
      RECT 7.2230 33.7365 7.2490 34.8300 ;
      RECT 7.1150 33.7365 7.1410 34.8300 ;
      RECT 7.0070 33.7365 7.0330 34.8300 ;
      RECT 6.8990 33.7365 6.9250 34.8300 ;
      RECT 6.7910 33.7365 6.8170 34.8300 ;
      RECT 6.6830 33.7365 6.7090 34.8300 ;
      RECT 6.5750 33.7365 6.6010 34.8300 ;
      RECT 6.4670 33.7365 6.4930 34.8300 ;
      RECT 6.3590 33.7365 6.3850 34.8300 ;
      RECT 6.2510 33.7365 6.2770 34.8300 ;
      RECT 6.1430 33.7365 6.1690 34.8300 ;
      RECT 6.0350 33.7365 6.0610 34.8300 ;
      RECT 5.9270 33.7365 5.9530 34.8300 ;
      RECT 5.7140 33.7365 5.7910 34.8300 ;
      RECT 3.8210 33.7365 3.8980 34.8300 ;
      RECT 3.6590 33.7365 3.6850 34.8300 ;
      RECT 3.5510 33.7365 3.5770 34.8300 ;
      RECT 3.4430 33.7365 3.4690 34.8300 ;
      RECT 3.3350 33.7365 3.3610 34.8300 ;
      RECT 3.2270 33.7365 3.2530 34.8300 ;
      RECT 3.1190 33.7365 3.1450 34.8300 ;
      RECT 3.0110 33.7365 3.0370 34.8300 ;
      RECT 2.9030 33.7365 2.9290 34.8300 ;
      RECT 2.7950 33.7365 2.8210 34.8300 ;
      RECT 2.6870 33.7365 2.7130 34.8300 ;
      RECT 2.5790 33.7365 2.6050 34.8300 ;
      RECT 2.4710 33.7365 2.4970 34.8300 ;
      RECT 2.3630 33.7365 2.3890 34.8300 ;
      RECT 2.2550 33.7365 2.2810 34.8300 ;
      RECT 2.1470 33.7365 2.1730 34.8300 ;
      RECT 2.0390 33.7365 2.0650 34.8300 ;
      RECT 1.9310 33.7365 1.9570 34.8300 ;
      RECT 1.8230 33.7365 1.8490 34.8300 ;
      RECT 1.7150 33.7365 1.7410 34.8300 ;
      RECT 1.6070 33.7365 1.6330 34.8300 ;
      RECT 1.4990 33.7365 1.5250 34.8300 ;
      RECT 1.3910 33.7365 1.4170 34.8300 ;
      RECT 1.2830 33.7365 1.3090 34.8300 ;
      RECT 1.1750 33.7365 1.2010 34.8300 ;
      RECT 1.0670 33.7365 1.0930 34.8300 ;
      RECT 0.9590 33.7365 0.9850 34.8300 ;
      RECT 0.8510 33.7365 0.8770 34.8300 ;
      RECT 0.7430 33.7365 0.7690 34.8300 ;
      RECT 0.6350 33.7365 0.6610 34.8300 ;
      RECT 0.5270 33.7365 0.5530 34.8300 ;
      RECT 0.4190 33.7365 0.4450 34.8300 ;
      RECT 0.3110 33.7365 0.3370 34.8300 ;
      RECT 0.2030 33.7365 0.2290 34.8300 ;
      RECT 0.0000 33.7365 0.0850 34.8300 ;
      RECT 5.1800 34.8165 5.3080 35.9100 ;
      RECT 5.1660 35.4820 5.3080 35.8045 ;
      RECT 5.0180 35.2090 5.0800 35.9100 ;
      RECT 5.0040 35.5185 5.0800 35.6720 ;
      RECT 5.0180 34.8165 5.0440 35.9100 ;
      RECT 5.0180 34.9375 5.0580 35.1770 ;
      RECT 5.0180 34.8165 5.0800 34.9055 ;
      RECT 4.7210 35.2670 4.9270 35.9100 ;
      RECT 4.9010 34.8165 4.9270 35.9100 ;
      RECT 4.7210 35.5440 4.9410 35.8020 ;
      RECT 4.7210 34.8165 4.8190 35.9100 ;
      RECT 4.3040 34.8165 4.3870 35.9100 ;
      RECT 4.3040 34.9050 4.4010 35.8405 ;
      RECT 9.5270 34.8165 9.6120 35.9100 ;
      RECT 9.3830 34.8165 9.4090 35.9100 ;
      RECT 9.2750 34.8165 9.3010 35.9100 ;
      RECT 9.1670 34.8165 9.1930 35.9100 ;
      RECT 9.0590 34.8165 9.0850 35.9100 ;
      RECT 8.9510 34.8165 8.9770 35.9100 ;
      RECT 8.8430 34.8165 8.8690 35.9100 ;
      RECT 8.7350 34.8165 8.7610 35.9100 ;
      RECT 8.6270 34.8165 8.6530 35.9100 ;
      RECT 8.5190 34.8165 8.5450 35.9100 ;
      RECT 8.4110 34.8165 8.4370 35.9100 ;
      RECT 8.3030 34.8165 8.3290 35.9100 ;
      RECT 8.1950 34.8165 8.2210 35.9100 ;
      RECT 8.0870 34.8165 8.1130 35.9100 ;
      RECT 7.9790 34.8165 8.0050 35.9100 ;
      RECT 7.8710 34.8165 7.8970 35.9100 ;
      RECT 7.7630 34.8165 7.7890 35.9100 ;
      RECT 7.6550 34.8165 7.6810 35.9100 ;
      RECT 7.5470 34.8165 7.5730 35.9100 ;
      RECT 7.4390 34.8165 7.4650 35.9100 ;
      RECT 7.3310 34.8165 7.3570 35.9100 ;
      RECT 7.2230 34.8165 7.2490 35.9100 ;
      RECT 7.1150 34.8165 7.1410 35.9100 ;
      RECT 7.0070 34.8165 7.0330 35.9100 ;
      RECT 6.8990 34.8165 6.9250 35.9100 ;
      RECT 6.7910 34.8165 6.8170 35.9100 ;
      RECT 6.6830 34.8165 6.7090 35.9100 ;
      RECT 6.5750 34.8165 6.6010 35.9100 ;
      RECT 6.4670 34.8165 6.4930 35.9100 ;
      RECT 6.3590 34.8165 6.3850 35.9100 ;
      RECT 6.2510 34.8165 6.2770 35.9100 ;
      RECT 6.1430 34.8165 6.1690 35.9100 ;
      RECT 6.0350 34.8165 6.0610 35.9100 ;
      RECT 5.9270 34.8165 5.9530 35.9100 ;
      RECT 5.7140 34.8165 5.7910 35.9100 ;
      RECT 3.8210 34.8165 3.8980 35.9100 ;
      RECT 3.6590 34.8165 3.6850 35.9100 ;
      RECT 3.5510 34.8165 3.5770 35.9100 ;
      RECT 3.4430 34.8165 3.4690 35.9100 ;
      RECT 3.3350 34.8165 3.3610 35.9100 ;
      RECT 3.2270 34.8165 3.2530 35.9100 ;
      RECT 3.1190 34.8165 3.1450 35.9100 ;
      RECT 3.0110 34.8165 3.0370 35.9100 ;
      RECT 2.9030 34.8165 2.9290 35.9100 ;
      RECT 2.7950 34.8165 2.8210 35.9100 ;
      RECT 2.6870 34.8165 2.7130 35.9100 ;
      RECT 2.5790 34.8165 2.6050 35.9100 ;
      RECT 2.4710 34.8165 2.4970 35.9100 ;
      RECT 2.3630 34.8165 2.3890 35.9100 ;
      RECT 2.2550 34.8165 2.2810 35.9100 ;
      RECT 2.1470 34.8165 2.1730 35.9100 ;
      RECT 2.0390 34.8165 2.0650 35.9100 ;
      RECT 1.9310 34.8165 1.9570 35.9100 ;
      RECT 1.8230 34.8165 1.8490 35.9100 ;
      RECT 1.7150 34.8165 1.7410 35.9100 ;
      RECT 1.6070 34.8165 1.6330 35.9100 ;
      RECT 1.4990 34.8165 1.5250 35.9100 ;
      RECT 1.3910 34.8165 1.4170 35.9100 ;
      RECT 1.2830 34.8165 1.3090 35.9100 ;
      RECT 1.1750 34.8165 1.2010 35.9100 ;
      RECT 1.0670 34.8165 1.0930 35.9100 ;
      RECT 0.9590 34.8165 0.9850 35.9100 ;
      RECT 0.8510 34.8165 0.8770 35.9100 ;
      RECT 0.7430 34.8165 0.7690 35.9100 ;
      RECT 0.6350 34.8165 0.6610 35.9100 ;
      RECT 0.5270 34.8165 0.5530 35.9100 ;
      RECT 0.4190 34.8165 0.4450 35.9100 ;
      RECT 0.3110 34.8165 0.3370 35.9100 ;
      RECT 0.2030 34.8165 0.2290 35.9100 ;
      RECT 0.0000 34.8165 0.0850 35.9100 ;
      RECT 5.1800 35.8965 5.3080 36.9900 ;
      RECT 5.1660 36.5620 5.3080 36.8845 ;
      RECT 5.0180 36.2890 5.0800 36.9900 ;
      RECT 5.0040 36.5985 5.0800 36.7520 ;
      RECT 5.0180 35.8965 5.0440 36.9900 ;
      RECT 5.0180 36.0175 5.0580 36.2570 ;
      RECT 5.0180 35.8965 5.0800 35.9855 ;
      RECT 4.7210 36.3470 4.9270 36.9900 ;
      RECT 4.9010 35.8965 4.9270 36.9900 ;
      RECT 4.7210 36.6240 4.9410 36.8820 ;
      RECT 4.7210 35.8965 4.8190 36.9900 ;
      RECT 4.3040 35.8965 4.3870 36.9900 ;
      RECT 4.3040 35.9850 4.4010 36.9205 ;
      RECT 9.5270 35.8965 9.6120 36.9900 ;
      RECT 9.3830 35.8965 9.4090 36.9900 ;
      RECT 9.2750 35.8965 9.3010 36.9900 ;
      RECT 9.1670 35.8965 9.1930 36.9900 ;
      RECT 9.0590 35.8965 9.0850 36.9900 ;
      RECT 8.9510 35.8965 8.9770 36.9900 ;
      RECT 8.8430 35.8965 8.8690 36.9900 ;
      RECT 8.7350 35.8965 8.7610 36.9900 ;
      RECT 8.6270 35.8965 8.6530 36.9900 ;
      RECT 8.5190 35.8965 8.5450 36.9900 ;
      RECT 8.4110 35.8965 8.4370 36.9900 ;
      RECT 8.3030 35.8965 8.3290 36.9900 ;
      RECT 8.1950 35.8965 8.2210 36.9900 ;
      RECT 8.0870 35.8965 8.1130 36.9900 ;
      RECT 7.9790 35.8965 8.0050 36.9900 ;
      RECT 7.8710 35.8965 7.8970 36.9900 ;
      RECT 7.7630 35.8965 7.7890 36.9900 ;
      RECT 7.6550 35.8965 7.6810 36.9900 ;
      RECT 7.5470 35.8965 7.5730 36.9900 ;
      RECT 7.4390 35.8965 7.4650 36.9900 ;
      RECT 7.3310 35.8965 7.3570 36.9900 ;
      RECT 7.2230 35.8965 7.2490 36.9900 ;
      RECT 7.1150 35.8965 7.1410 36.9900 ;
      RECT 7.0070 35.8965 7.0330 36.9900 ;
      RECT 6.8990 35.8965 6.9250 36.9900 ;
      RECT 6.7910 35.8965 6.8170 36.9900 ;
      RECT 6.6830 35.8965 6.7090 36.9900 ;
      RECT 6.5750 35.8965 6.6010 36.9900 ;
      RECT 6.4670 35.8965 6.4930 36.9900 ;
      RECT 6.3590 35.8965 6.3850 36.9900 ;
      RECT 6.2510 35.8965 6.2770 36.9900 ;
      RECT 6.1430 35.8965 6.1690 36.9900 ;
      RECT 6.0350 35.8965 6.0610 36.9900 ;
      RECT 5.9270 35.8965 5.9530 36.9900 ;
      RECT 5.7140 35.8965 5.7910 36.9900 ;
      RECT 3.8210 35.8965 3.8980 36.9900 ;
      RECT 3.6590 35.8965 3.6850 36.9900 ;
      RECT 3.5510 35.8965 3.5770 36.9900 ;
      RECT 3.4430 35.8965 3.4690 36.9900 ;
      RECT 3.3350 35.8965 3.3610 36.9900 ;
      RECT 3.2270 35.8965 3.2530 36.9900 ;
      RECT 3.1190 35.8965 3.1450 36.9900 ;
      RECT 3.0110 35.8965 3.0370 36.9900 ;
      RECT 2.9030 35.8965 2.9290 36.9900 ;
      RECT 2.7950 35.8965 2.8210 36.9900 ;
      RECT 2.6870 35.8965 2.7130 36.9900 ;
      RECT 2.5790 35.8965 2.6050 36.9900 ;
      RECT 2.4710 35.8965 2.4970 36.9900 ;
      RECT 2.3630 35.8965 2.3890 36.9900 ;
      RECT 2.2550 35.8965 2.2810 36.9900 ;
      RECT 2.1470 35.8965 2.1730 36.9900 ;
      RECT 2.0390 35.8965 2.0650 36.9900 ;
      RECT 1.9310 35.8965 1.9570 36.9900 ;
      RECT 1.8230 35.8965 1.8490 36.9900 ;
      RECT 1.7150 35.8965 1.7410 36.9900 ;
      RECT 1.6070 35.8965 1.6330 36.9900 ;
      RECT 1.4990 35.8965 1.5250 36.9900 ;
      RECT 1.3910 35.8965 1.4170 36.9900 ;
      RECT 1.2830 35.8965 1.3090 36.9900 ;
      RECT 1.1750 35.8965 1.2010 36.9900 ;
      RECT 1.0670 35.8965 1.0930 36.9900 ;
      RECT 0.9590 35.8965 0.9850 36.9900 ;
      RECT 0.8510 35.8965 0.8770 36.9900 ;
      RECT 0.7430 35.8965 0.7690 36.9900 ;
      RECT 0.6350 35.8965 0.6610 36.9900 ;
      RECT 0.5270 35.8965 0.5530 36.9900 ;
      RECT 0.4190 35.8965 0.4450 36.9900 ;
      RECT 0.3110 35.8965 0.3370 36.9900 ;
      RECT 0.2030 35.8965 0.2290 36.9900 ;
      RECT 0.0000 35.8965 0.0850 36.9900 ;
      RECT 5.1800 36.9765 5.3080 38.0700 ;
      RECT 5.1660 37.6420 5.3080 37.9645 ;
      RECT 5.0180 37.3690 5.0800 38.0700 ;
      RECT 5.0040 37.6785 5.0800 37.8320 ;
      RECT 5.0180 36.9765 5.0440 38.0700 ;
      RECT 5.0180 37.0975 5.0580 37.3370 ;
      RECT 5.0180 36.9765 5.0800 37.0655 ;
      RECT 4.7210 37.4270 4.9270 38.0700 ;
      RECT 4.9010 36.9765 4.9270 38.0700 ;
      RECT 4.7210 37.7040 4.9410 37.9620 ;
      RECT 4.7210 36.9765 4.8190 38.0700 ;
      RECT 4.3040 36.9765 4.3870 38.0700 ;
      RECT 4.3040 37.0650 4.4010 38.0005 ;
      RECT 9.5270 36.9765 9.6120 38.0700 ;
      RECT 9.3830 36.9765 9.4090 38.0700 ;
      RECT 9.2750 36.9765 9.3010 38.0700 ;
      RECT 9.1670 36.9765 9.1930 38.0700 ;
      RECT 9.0590 36.9765 9.0850 38.0700 ;
      RECT 8.9510 36.9765 8.9770 38.0700 ;
      RECT 8.8430 36.9765 8.8690 38.0700 ;
      RECT 8.7350 36.9765 8.7610 38.0700 ;
      RECT 8.6270 36.9765 8.6530 38.0700 ;
      RECT 8.5190 36.9765 8.5450 38.0700 ;
      RECT 8.4110 36.9765 8.4370 38.0700 ;
      RECT 8.3030 36.9765 8.3290 38.0700 ;
      RECT 8.1950 36.9765 8.2210 38.0700 ;
      RECT 8.0870 36.9765 8.1130 38.0700 ;
      RECT 7.9790 36.9765 8.0050 38.0700 ;
      RECT 7.8710 36.9765 7.8970 38.0700 ;
      RECT 7.7630 36.9765 7.7890 38.0700 ;
      RECT 7.6550 36.9765 7.6810 38.0700 ;
      RECT 7.5470 36.9765 7.5730 38.0700 ;
      RECT 7.4390 36.9765 7.4650 38.0700 ;
      RECT 7.3310 36.9765 7.3570 38.0700 ;
      RECT 7.2230 36.9765 7.2490 38.0700 ;
      RECT 7.1150 36.9765 7.1410 38.0700 ;
      RECT 7.0070 36.9765 7.0330 38.0700 ;
      RECT 6.8990 36.9765 6.9250 38.0700 ;
      RECT 6.7910 36.9765 6.8170 38.0700 ;
      RECT 6.6830 36.9765 6.7090 38.0700 ;
      RECT 6.5750 36.9765 6.6010 38.0700 ;
      RECT 6.4670 36.9765 6.4930 38.0700 ;
      RECT 6.3590 36.9765 6.3850 38.0700 ;
      RECT 6.2510 36.9765 6.2770 38.0700 ;
      RECT 6.1430 36.9765 6.1690 38.0700 ;
      RECT 6.0350 36.9765 6.0610 38.0700 ;
      RECT 5.9270 36.9765 5.9530 38.0700 ;
      RECT 5.7140 36.9765 5.7910 38.0700 ;
      RECT 3.8210 36.9765 3.8980 38.0700 ;
      RECT 3.6590 36.9765 3.6850 38.0700 ;
      RECT 3.5510 36.9765 3.5770 38.0700 ;
      RECT 3.4430 36.9765 3.4690 38.0700 ;
      RECT 3.3350 36.9765 3.3610 38.0700 ;
      RECT 3.2270 36.9765 3.2530 38.0700 ;
      RECT 3.1190 36.9765 3.1450 38.0700 ;
      RECT 3.0110 36.9765 3.0370 38.0700 ;
      RECT 2.9030 36.9765 2.9290 38.0700 ;
      RECT 2.7950 36.9765 2.8210 38.0700 ;
      RECT 2.6870 36.9765 2.7130 38.0700 ;
      RECT 2.5790 36.9765 2.6050 38.0700 ;
      RECT 2.4710 36.9765 2.4970 38.0700 ;
      RECT 2.3630 36.9765 2.3890 38.0700 ;
      RECT 2.2550 36.9765 2.2810 38.0700 ;
      RECT 2.1470 36.9765 2.1730 38.0700 ;
      RECT 2.0390 36.9765 2.0650 38.0700 ;
      RECT 1.9310 36.9765 1.9570 38.0700 ;
      RECT 1.8230 36.9765 1.8490 38.0700 ;
      RECT 1.7150 36.9765 1.7410 38.0700 ;
      RECT 1.6070 36.9765 1.6330 38.0700 ;
      RECT 1.4990 36.9765 1.5250 38.0700 ;
      RECT 1.3910 36.9765 1.4170 38.0700 ;
      RECT 1.2830 36.9765 1.3090 38.0700 ;
      RECT 1.1750 36.9765 1.2010 38.0700 ;
      RECT 1.0670 36.9765 1.0930 38.0700 ;
      RECT 0.9590 36.9765 0.9850 38.0700 ;
      RECT 0.8510 36.9765 0.8770 38.0700 ;
      RECT 0.7430 36.9765 0.7690 38.0700 ;
      RECT 0.6350 36.9765 0.6610 38.0700 ;
      RECT 0.5270 36.9765 0.5530 38.0700 ;
      RECT 0.4190 36.9765 0.4450 38.0700 ;
      RECT 0.3110 36.9765 0.3370 38.0700 ;
      RECT 0.2030 36.9765 0.2290 38.0700 ;
      RECT 0.0000 36.9765 0.0850 38.0700 ;
      RECT 5.1800 38.0565 5.3080 39.1500 ;
      RECT 5.1660 38.7220 5.3080 39.0445 ;
      RECT 5.0180 38.4490 5.0800 39.1500 ;
      RECT 5.0040 38.7585 5.0800 38.9120 ;
      RECT 5.0180 38.0565 5.0440 39.1500 ;
      RECT 5.0180 38.1775 5.0580 38.4170 ;
      RECT 5.0180 38.0565 5.0800 38.1455 ;
      RECT 4.7210 38.5070 4.9270 39.1500 ;
      RECT 4.9010 38.0565 4.9270 39.1500 ;
      RECT 4.7210 38.7840 4.9410 39.0420 ;
      RECT 4.7210 38.0565 4.8190 39.1500 ;
      RECT 4.3040 38.0565 4.3870 39.1500 ;
      RECT 4.3040 38.1450 4.4010 39.0805 ;
      RECT 9.5270 38.0565 9.6120 39.1500 ;
      RECT 9.3830 38.0565 9.4090 39.1500 ;
      RECT 9.2750 38.0565 9.3010 39.1500 ;
      RECT 9.1670 38.0565 9.1930 39.1500 ;
      RECT 9.0590 38.0565 9.0850 39.1500 ;
      RECT 8.9510 38.0565 8.9770 39.1500 ;
      RECT 8.8430 38.0565 8.8690 39.1500 ;
      RECT 8.7350 38.0565 8.7610 39.1500 ;
      RECT 8.6270 38.0565 8.6530 39.1500 ;
      RECT 8.5190 38.0565 8.5450 39.1500 ;
      RECT 8.4110 38.0565 8.4370 39.1500 ;
      RECT 8.3030 38.0565 8.3290 39.1500 ;
      RECT 8.1950 38.0565 8.2210 39.1500 ;
      RECT 8.0870 38.0565 8.1130 39.1500 ;
      RECT 7.9790 38.0565 8.0050 39.1500 ;
      RECT 7.8710 38.0565 7.8970 39.1500 ;
      RECT 7.7630 38.0565 7.7890 39.1500 ;
      RECT 7.6550 38.0565 7.6810 39.1500 ;
      RECT 7.5470 38.0565 7.5730 39.1500 ;
      RECT 7.4390 38.0565 7.4650 39.1500 ;
      RECT 7.3310 38.0565 7.3570 39.1500 ;
      RECT 7.2230 38.0565 7.2490 39.1500 ;
      RECT 7.1150 38.0565 7.1410 39.1500 ;
      RECT 7.0070 38.0565 7.0330 39.1500 ;
      RECT 6.8990 38.0565 6.9250 39.1500 ;
      RECT 6.7910 38.0565 6.8170 39.1500 ;
      RECT 6.6830 38.0565 6.7090 39.1500 ;
      RECT 6.5750 38.0565 6.6010 39.1500 ;
      RECT 6.4670 38.0565 6.4930 39.1500 ;
      RECT 6.3590 38.0565 6.3850 39.1500 ;
      RECT 6.2510 38.0565 6.2770 39.1500 ;
      RECT 6.1430 38.0565 6.1690 39.1500 ;
      RECT 6.0350 38.0565 6.0610 39.1500 ;
      RECT 5.9270 38.0565 5.9530 39.1500 ;
      RECT 5.7140 38.0565 5.7910 39.1500 ;
      RECT 3.8210 38.0565 3.8980 39.1500 ;
      RECT 3.6590 38.0565 3.6850 39.1500 ;
      RECT 3.5510 38.0565 3.5770 39.1500 ;
      RECT 3.4430 38.0565 3.4690 39.1500 ;
      RECT 3.3350 38.0565 3.3610 39.1500 ;
      RECT 3.2270 38.0565 3.2530 39.1500 ;
      RECT 3.1190 38.0565 3.1450 39.1500 ;
      RECT 3.0110 38.0565 3.0370 39.1500 ;
      RECT 2.9030 38.0565 2.9290 39.1500 ;
      RECT 2.7950 38.0565 2.8210 39.1500 ;
      RECT 2.6870 38.0565 2.7130 39.1500 ;
      RECT 2.5790 38.0565 2.6050 39.1500 ;
      RECT 2.4710 38.0565 2.4970 39.1500 ;
      RECT 2.3630 38.0565 2.3890 39.1500 ;
      RECT 2.2550 38.0565 2.2810 39.1500 ;
      RECT 2.1470 38.0565 2.1730 39.1500 ;
      RECT 2.0390 38.0565 2.0650 39.1500 ;
      RECT 1.9310 38.0565 1.9570 39.1500 ;
      RECT 1.8230 38.0565 1.8490 39.1500 ;
      RECT 1.7150 38.0565 1.7410 39.1500 ;
      RECT 1.6070 38.0565 1.6330 39.1500 ;
      RECT 1.4990 38.0565 1.5250 39.1500 ;
      RECT 1.3910 38.0565 1.4170 39.1500 ;
      RECT 1.2830 38.0565 1.3090 39.1500 ;
      RECT 1.1750 38.0565 1.2010 39.1500 ;
      RECT 1.0670 38.0565 1.0930 39.1500 ;
      RECT 0.9590 38.0565 0.9850 39.1500 ;
      RECT 0.8510 38.0565 0.8770 39.1500 ;
      RECT 0.7430 38.0565 0.7690 39.1500 ;
      RECT 0.6350 38.0565 0.6610 39.1500 ;
      RECT 0.5270 38.0565 0.5530 39.1500 ;
      RECT 0.4190 38.0565 0.4450 39.1500 ;
      RECT 0.3110 38.0565 0.3370 39.1500 ;
      RECT 0.2030 38.0565 0.2290 39.1500 ;
      RECT 0.0000 38.0565 0.0850 39.1500 ;
      RECT 5.1800 39.1365 5.3080 40.2300 ;
      RECT 5.1660 39.8020 5.3080 40.1245 ;
      RECT 5.0180 39.5290 5.0800 40.2300 ;
      RECT 5.0040 39.8385 5.0800 39.9920 ;
      RECT 5.0180 39.1365 5.0440 40.2300 ;
      RECT 5.0180 39.2575 5.0580 39.4970 ;
      RECT 5.0180 39.1365 5.0800 39.2255 ;
      RECT 4.7210 39.5870 4.9270 40.2300 ;
      RECT 4.9010 39.1365 4.9270 40.2300 ;
      RECT 4.7210 39.8640 4.9410 40.1220 ;
      RECT 4.7210 39.1365 4.8190 40.2300 ;
      RECT 4.3040 39.1365 4.3870 40.2300 ;
      RECT 4.3040 39.2250 4.4010 40.1605 ;
      RECT 9.5270 39.1365 9.6120 40.2300 ;
      RECT 9.3830 39.1365 9.4090 40.2300 ;
      RECT 9.2750 39.1365 9.3010 40.2300 ;
      RECT 9.1670 39.1365 9.1930 40.2300 ;
      RECT 9.0590 39.1365 9.0850 40.2300 ;
      RECT 8.9510 39.1365 8.9770 40.2300 ;
      RECT 8.8430 39.1365 8.8690 40.2300 ;
      RECT 8.7350 39.1365 8.7610 40.2300 ;
      RECT 8.6270 39.1365 8.6530 40.2300 ;
      RECT 8.5190 39.1365 8.5450 40.2300 ;
      RECT 8.4110 39.1365 8.4370 40.2300 ;
      RECT 8.3030 39.1365 8.3290 40.2300 ;
      RECT 8.1950 39.1365 8.2210 40.2300 ;
      RECT 8.0870 39.1365 8.1130 40.2300 ;
      RECT 7.9790 39.1365 8.0050 40.2300 ;
      RECT 7.8710 39.1365 7.8970 40.2300 ;
      RECT 7.7630 39.1365 7.7890 40.2300 ;
      RECT 7.6550 39.1365 7.6810 40.2300 ;
      RECT 7.5470 39.1365 7.5730 40.2300 ;
      RECT 7.4390 39.1365 7.4650 40.2300 ;
      RECT 7.3310 39.1365 7.3570 40.2300 ;
      RECT 7.2230 39.1365 7.2490 40.2300 ;
      RECT 7.1150 39.1365 7.1410 40.2300 ;
      RECT 7.0070 39.1365 7.0330 40.2300 ;
      RECT 6.8990 39.1365 6.9250 40.2300 ;
      RECT 6.7910 39.1365 6.8170 40.2300 ;
      RECT 6.6830 39.1365 6.7090 40.2300 ;
      RECT 6.5750 39.1365 6.6010 40.2300 ;
      RECT 6.4670 39.1365 6.4930 40.2300 ;
      RECT 6.3590 39.1365 6.3850 40.2300 ;
      RECT 6.2510 39.1365 6.2770 40.2300 ;
      RECT 6.1430 39.1365 6.1690 40.2300 ;
      RECT 6.0350 39.1365 6.0610 40.2300 ;
      RECT 5.9270 39.1365 5.9530 40.2300 ;
      RECT 5.7140 39.1365 5.7910 40.2300 ;
      RECT 3.8210 39.1365 3.8980 40.2300 ;
      RECT 3.6590 39.1365 3.6850 40.2300 ;
      RECT 3.5510 39.1365 3.5770 40.2300 ;
      RECT 3.4430 39.1365 3.4690 40.2300 ;
      RECT 3.3350 39.1365 3.3610 40.2300 ;
      RECT 3.2270 39.1365 3.2530 40.2300 ;
      RECT 3.1190 39.1365 3.1450 40.2300 ;
      RECT 3.0110 39.1365 3.0370 40.2300 ;
      RECT 2.9030 39.1365 2.9290 40.2300 ;
      RECT 2.7950 39.1365 2.8210 40.2300 ;
      RECT 2.6870 39.1365 2.7130 40.2300 ;
      RECT 2.5790 39.1365 2.6050 40.2300 ;
      RECT 2.4710 39.1365 2.4970 40.2300 ;
      RECT 2.3630 39.1365 2.3890 40.2300 ;
      RECT 2.2550 39.1365 2.2810 40.2300 ;
      RECT 2.1470 39.1365 2.1730 40.2300 ;
      RECT 2.0390 39.1365 2.0650 40.2300 ;
      RECT 1.9310 39.1365 1.9570 40.2300 ;
      RECT 1.8230 39.1365 1.8490 40.2300 ;
      RECT 1.7150 39.1365 1.7410 40.2300 ;
      RECT 1.6070 39.1365 1.6330 40.2300 ;
      RECT 1.4990 39.1365 1.5250 40.2300 ;
      RECT 1.3910 39.1365 1.4170 40.2300 ;
      RECT 1.2830 39.1365 1.3090 40.2300 ;
      RECT 1.1750 39.1365 1.2010 40.2300 ;
      RECT 1.0670 39.1365 1.0930 40.2300 ;
      RECT 0.9590 39.1365 0.9850 40.2300 ;
      RECT 0.8510 39.1365 0.8770 40.2300 ;
      RECT 0.7430 39.1365 0.7690 40.2300 ;
      RECT 0.6350 39.1365 0.6610 40.2300 ;
      RECT 0.5270 39.1365 0.5530 40.2300 ;
      RECT 0.4190 39.1365 0.4450 40.2300 ;
      RECT 0.3110 39.1365 0.3370 40.2300 ;
      RECT 0.2030 39.1365 0.2290 40.2300 ;
      RECT 0.0000 39.1365 0.0850 40.2300 ;
      RECT 5.1800 40.2165 5.3080 41.3100 ;
      RECT 5.1660 40.8820 5.3080 41.2045 ;
      RECT 5.0180 40.6090 5.0800 41.3100 ;
      RECT 5.0040 40.9185 5.0800 41.0720 ;
      RECT 5.0180 40.2165 5.0440 41.3100 ;
      RECT 5.0180 40.3375 5.0580 40.5770 ;
      RECT 5.0180 40.2165 5.0800 40.3055 ;
      RECT 4.7210 40.6670 4.9270 41.3100 ;
      RECT 4.9010 40.2165 4.9270 41.3100 ;
      RECT 4.7210 40.9440 4.9410 41.2020 ;
      RECT 4.7210 40.2165 4.8190 41.3100 ;
      RECT 4.3040 40.2165 4.3870 41.3100 ;
      RECT 4.3040 40.3050 4.4010 41.2405 ;
      RECT 9.5270 40.2165 9.6120 41.3100 ;
      RECT 9.3830 40.2165 9.4090 41.3100 ;
      RECT 9.2750 40.2165 9.3010 41.3100 ;
      RECT 9.1670 40.2165 9.1930 41.3100 ;
      RECT 9.0590 40.2165 9.0850 41.3100 ;
      RECT 8.9510 40.2165 8.9770 41.3100 ;
      RECT 8.8430 40.2165 8.8690 41.3100 ;
      RECT 8.7350 40.2165 8.7610 41.3100 ;
      RECT 8.6270 40.2165 8.6530 41.3100 ;
      RECT 8.5190 40.2165 8.5450 41.3100 ;
      RECT 8.4110 40.2165 8.4370 41.3100 ;
      RECT 8.3030 40.2165 8.3290 41.3100 ;
      RECT 8.1950 40.2165 8.2210 41.3100 ;
      RECT 8.0870 40.2165 8.1130 41.3100 ;
      RECT 7.9790 40.2165 8.0050 41.3100 ;
      RECT 7.8710 40.2165 7.8970 41.3100 ;
      RECT 7.7630 40.2165 7.7890 41.3100 ;
      RECT 7.6550 40.2165 7.6810 41.3100 ;
      RECT 7.5470 40.2165 7.5730 41.3100 ;
      RECT 7.4390 40.2165 7.4650 41.3100 ;
      RECT 7.3310 40.2165 7.3570 41.3100 ;
      RECT 7.2230 40.2165 7.2490 41.3100 ;
      RECT 7.1150 40.2165 7.1410 41.3100 ;
      RECT 7.0070 40.2165 7.0330 41.3100 ;
      RECT 6.8990 40.2165 6.9250 41.3100 ;
      RECT 6.7910 40.2165 6.8170 41.3100 ;
      RECT 6.6830 40.2165 6.7090 41.3100 ;
      RECT 6.5750 40.2165 6.6010 41.3100 ;
      RECT 6.4670 40.2165 6.4930 41.3100 ;
      RECT 6.3590 40.2165 6.3850 41.3100 ;
      RECT 6.2510 40.2165 6.2770 41.3100 ;
      RECT 6.1430 40.2165 6.1690 41.3100 ;
      RECT 6.0350 40.2165 6.0610 41.3100 ;
      RECT 5.9270 40.2165 5.9530 41.3100 ;
      RECT 5.7140 40.2165 5.7910 41.3100 ;
      RECT 3.8210 40.2165 3.8980 41.3100 ;
      RECT 3.6590 40.2165 3.6850 41.3100 ;
      RECT 3.5510 40.2165 3.5770 41.3100 ;
      RECT 3.4430 40.2165 3.4690 41.3100 ;
      RECT 3.3350 40.2165 3.3610 41.3100 ;
      RECT 3.2270 40.2165 3.2530 41.3100 ;
      RECT 3.1190 40.2165 3.1450 41.3100 ;
      RECT 3.0110 40.2165 3.0370 41.3100 ;
      RECT 2.9030 40.2165 2.9290 41.3100 ;
      RECT 2.7950 40.2165 2.8210 41.3100 ;
      RECT 2.6870 40.2165 2.7130 41.3100 ;
      RECT 2.5790 40.2165 2.6050 41.3100 ;
      RECT 2.4710 40.2165 2.4970 41.3100 ;
      RECT 2.3630 40.2165 2.3890 41.3100 ;
      RECT 2.2550 40.2165 2.2810 41.3100 ;
      RECT 2.1470 40.2165 2.1730 41.3100 ;
      RECT 2.0390 40.2165 2.0650 41.3100 ;
      RECT 1.9310 40.2165 1.9570 41.3100 ;
      RECT 1.8230 40.2165 1.8490 41.3100 ;
      RECT 1.7150 40.2165 1.7410 41.3100 ;
      RECT 1.6070 40.2165 1.6330 41.3100 ;
      RECT 1.4990 40.2165 1.5250 41.3100 ;
      RECT 1.3910 40.2165 1.4170 41.3100 ;
      RECT 1.2830 40.2165 1.3090 41.3100 ;
      RECT 1.1750 40.2165 1.2010 41.3100 ;
      RECT 1.0670 40.2165 1.0930 41.3100 ;
      RECT 0.9590 40.2165 0.9850 41.3100 ;
      RECT 0.8510 40.2165 0.8770 41.3100 ;
      RECT 0.7430 40.2165 0.7690 41.3100 ;
      RECT 0.6350 40.2165 0.6610 41.3100 ;
      RECT 0.5270 40.2165 0.5530 41.3100 ;
      RECT 0.4190 40.2165 0.4450 41.3100 ;
      RECT 0.3110 40.2165 0.3370 41.3100 ;
      RECT 0.2030 40.2165 0.2290 41.3100 ;
      RECT 0.0000 40.2165 0.0850 41.3100 ;
      RECT 5.1800 41.2965 5.3080 42.3900 ;
      RECT 5.1660 41.9620 5.3080 42.2845 ;
      RECT 5.0180 41.6890 5.0800 42.3900 ;
      RECT 5.0040 41.9985 5.0800 42.1520 ;
      RECT 5.0180 41.2965 5.0440 42.3900 ;
      RECT 5.0180 41.4175 5.0580 41.6570 ;
      RECT 5.0180 41.2965 5.0800 41.3855 ;
      RECT 4.7210 41.7470 4.9270 42.3900 ;
      RECT 4.9010 41.2965 4.9270 42.3900 ;
      RECT 4.7210 42.0240 4.9410 42.2820 ;
      RECT 4.7210 41.2965 4.8190 42.3900 ;
      RECT 4.3040 41.2965 4.3870 42.3900 ;
      RECT 4.3040 41.3850 4.4010 42.3205 ;
      RECT 9.5270 41.2965 9.6120 42.3900 ;
      RECT 9.3830 41.2965 9.4090 42.3900 ;
      RECT 9.2750 41.2965 9.3010 42.3900 ;
      RECT 9.1670 41.2965 9.1930 42.3900 ;
      RECT 9.0590 41.2965 9.0850 42.3900 ;
      RECT 8.9510 41.2965 8.9770 42.3900 ;
      RECT 8.8430 41.2965 8.8690 42.3900 ;
      RECT 8.7350 41.2965 8.7610 42.3900 ;
      RECT 8.6270 41.2965 8.6530 42.3900 ;
      RECT 8.5190 41.2965 8.5450 42.3900 ;
      RECT 8.4110 41.2965 8.4370 42.3900 ;
      RECT 8.3030 41.2965 8.3290 42.3900 ;
      RECT 8.1950 41.2965 8.2210 42.3900 ;
      RECT 8.0870 41.2965 8.1130 42.3900 ;
      RECT 7.9790 41.2965 8.0050 42.3900 ;
      RECT 7.8710 41.2965 7.8970 42.3900 ;
      RECT 7.7630 41.2965 7.7890 42.3900 ;
      RECT 7.6550 41.2965 7.6810 42.3900 ;
      RECT 7.5470 41.2965 7.5730 42.3900 ;
      RECT 7.4390 41.2965 7.4650 42.3900 ;
      RECT 7.3310 41.2965 7.3570 42.3900 ;
      RECT 7.2230 41.2965 7.2490 42.3900 ;
      RECT 7.1150 41.2965 7.1410 42.3900 ;
      RECT 7.0070 41.2965 7.0330 42.3900 ;
      RECT 6.8990 41.2965 6.9250 42.3900 ;
      RECT 6.7910 41.2965 6.8170 42.3900 ;
      RECT 6.6830 41.2965 6.7090 42.3900 ;
      RECT 6.5750 41.2965 6.6010 42.3900 ;
      RECT 6.4670 41.2965 6.4930 42.3900 ;
      RECT 6.3590 41.2965 6.3850 42.3900 ;
      RECT 6.2510 41.2965 6.2770 42.3900 ;
      RECT 6.1430 41.2965 6.1690 42.3900 ;
      RECT 6.0350 41.2965 6.0610 42.3900 ;
      RECT 5.9270 41.2965 5.9530 42.3900 ;
      RECT 5.7140 41.2965 5.7910 42.3900 ;
      RECT 3.8210 41.2965 3.8980 42.3900 ;
      RECT 3.6590 41.2965 3.6850 42.3900 ;
      RECT 3.5510 41.2965 3.5770 42.3900 ;
      RECT 3.4430 41.2965 3.4690 42.3900 ;
      RECT 3.3350 41.2965 3.3610 42.3900 ;
      RECT 3.2270 41.2965 3.2530 42.3900 ;
      RECT 3.1190 41.2965 3.1450 42.3900 ;
      RECT 3.0110 41.2965 3.0370 42.3900 ;
      RECT 2.9030 41.2965 2.9290 42.3900 ;
      RECT 2.7950 41.2965 2.8210 42.3900 ;
      RECT 2.6870 41.2965 2.7130 42.3900 ;
      RECT 2.5790 41.2965 2.6050 42.3900 ;
      RECT 2.4710 41.2965 2.4970 42.3900 ;
      RECT 2.3630 41.2965 2.3890 42.3900 ;
      RECT 2.2550 41.2965 2.2810 42.3900 ;
      RECT 2.1470 41.2965 2.1730 42.3900 ;
      RECT 2.0390 41.2965 2.0650 42.3900 ;
      RECT 1.9310 41.2965 1.9570 42.3900 ;
      RECT 1.8230 41.2965 1.8490 42.3900 ;
      RECT 1.7150 41.2965 1.7410 42.3900 ;
      RECT 1.6070 41.2965 1.6330 42.3900 ;
      RECT 1.4990 41.2965 1.5250 42.3900 ;
      RECT 1.3910 41.2965 1.4170 42.3900 ;
      RECT 1.2830 41.2965 1.3090 42.3900 ;
      RECT 1.1750 41.2965 1.2010 42.3900 ;
      RECT 1.0670 41.2965 1.0930 42.3900 ;
      RECT 0.9590 41.2965 0.9850 42.3900 ;
      RECT 0.8510 41.2965 0.8770 42.3900 ;
      RECT 0.7430 41.2965 0.7690 42.3900 ;
      RECT 0.6350 41.2965 0.6610 42.3900 ;
      RECT 0.5270 41.2965 0.5530 42.3900 ;
      RECT 0.4190 41.2965 0.4450 42.3900 ;
      RECT 0.3110 41.2965 0.3370 42.3900 ;
      RECT 0.2030 41.2965 0.2290 42.3900 ;
      RECT 0.0000 41.2965 0.0850 42.3900 ;
      RECT 5.1800 42.3765 5.3080 43.4700 ;
      RECT 5.1660 43.0420 5.3080 43.3645 ;
      RECT 5.0180 42.7690 5.0800 43.4700 ;
      RECT 5.0040 43.0785 5.0800 43.2320 ;
      RECT 5.0180 42.3765 5.0440 43.4700 ;
      RECT 5.0180 42.4975 5.0580 42.7370 ;
      RECT 5.0180 42.3765 5.0800 42.4655 ;
      RECT 4.7210 42.8270 4.9270 43.4700 ;
      RECT 4.9010 42.3765 4.9270 43.4700 ;
      RECT 4.7210 43.1040 4.9410 43.3620 ;
      RECT 4.7210 42.3765 4.8190 43.4700 ;
      RECT 4.3040 42.3765 4.3870 43.4700 ;
      RECT 4.3040 42.4650 4.4010 43.4005 ;
      RECT 9.5270 42.3765 9.6120 43.4700 ;
      RECT 9.3830 42.3765 9.4090 43.4700 ;
      RECT 9.2750 42.3765 9.3010 43.4700 ;
      RECT 9.1670 42.3765 9.1930 43.4700 ;
      RECT 9.0590 42.3765 9.0850 43.4700 ;
      RECT 8.9510 42.3765 8.9770 43.4700 ;
      RECT 8.8430 42.3765 8.8690 43.4700 ;
      RECT 8.7350 42.3765 8.7610 43.4700 ;
      RECT 8.6270 42.3765 8.6530 43.4700 ;
      RECT 8.5190 42.3765 8.5450 43.4700 ;
      RECT 8.4110 42.3765 8.4370 43.4700 ;
      RECT 8.3030 42.3765 8.3290 43.4700 ;
      RECT 8.1950 42.3765 8.2210 43.4700 ;
      RECT 8.0870 42.3765 8.1130 43.4700 ;
      RECT 7.9790 42.3765 8.0050 43.4700 ;
      RECT 7.8710 42.3765 7.8970 43.4700 ;
      RECT 7.7630 42.3765 7.7890 43.4700 ;
      RECT 7.6550 42.3765 7.6810 43.4700 ;
      RECT 7.5470 42.3765 7.5730 43.4700 ;
      RECT 7.4390 42.3765 7.4650 43.4700 ;
      RECT 7.3310 42.3765 7.3570 43.4700 ;
      RECT 7.2230 42.3765 7.2490 43.4700 ;
      RECT 7.1150 42.3765 7.1410 43.4700 ;
      RECT 7.0070 42.3765 7.0330 43.4700 ;
      RECT 6.8990 42.3765 6.9250 43.4700 ;
      RECT 6.7910 42.3765 6.8170 43.4700 ;
      RECT 6.6830 42.3765 6.7090 43.4700 ;
      RECT 6.5750 42.3765 6.6010 43.4700 ;
      RECT 6.4670 42.3765 6.4930 43.4700 ;
      RECT 6.3590 42.3765 6.3850 43.4700 ;
      RECT 6.2510 42.3765 6.2770 43.4700 ;
      RECT 6.1430 42.3765 6.1690 43.4700 ;
      RECT 6.0350 42.3765 6.0610 43.4700 ;
      RECT 5.9270 42.3765 5.9530 43.4700 ;
      RECT 5.7140 42.3765 5.7910 43.4700 ;
      RECT 3.8210 42.3765 3.8980 43.4700 ;
      RECT 3.6590 42.3765 3.6850 43.4700 ;
      RECT 3.5510 42.3765 3.5770 43.4700 ;
      RECT 3.4430 42.3765 3.4690 43.4700 ;
      RECT 3.3350 42.3765 3.3610 43.4700 ;
      RECT 3.2270 42.3765 3.2530 43.4700 ;
      RECT 3.1190 42.3765 3.1450 43.4700 ;
      RECT 3.0110 42.3765 3.0370 43.4700 ;
      RECT 2.9030 42.3765 2.9290 43.4700 ;
      RECT 2.7950 42.3765 2.8210 43.4700 ;
      RECT 2.6870 42.3765 2.7130 43.4700 ;
      RECT 2.5790 42.3765 2.6050 43.4700 ;
      RECT 2.4710 42.3765 2.4970 43.4700 ;
      RECT 2.3630 42.3765 2.3890 43.4700 ;
      RECT 2.2550 42.3765 2.2810 43.4700 ;
      RECT 2.1470 42.3765 2.1730 43.4700 ;
      RECT 2.0390 42.3765 2.0650 43.4700 ;
      RECT 1.9310 42.3765 1.9570 43.4700 ;
      RECT 1.8230 42.3765 1.8490 43.4700 ;
      RECT 1.7150 42.3765 1.7410 43.4700 ;
      RECT 1.6070 42.3765 1.6330 43.4700 ;
      RECT 1.4990 42.3765 1.5250 43.4700 ;
      RECT 1.3910 42.3765 1.4170 43.4700 ;
      RECT 1.2830 42.3765 1.3090 43.4700 ;
      RECT 1.1750 42.3765 1.2010 43.4700 ;
      RECT 1.0670 42.3765 1.0930 43.4700 ;
      RECT 0.9590 42.3765 0.9850 43.4700 ;
      RECT 0.8510 42.3765 0.8770 43.4700 ;
      RECT 0.7430 42.3765 0.7690 43.4700 ;
      RECT 0.6350 42.3765 0.6610 43.4700 ;
      RECT 0.5270 42.3765 0.5530 43.4700 ;
      RECT 0.4190 42.3765 0.4450 43.4700 ;
      RECT 0.3110 42.3765 0.3370 43.4700 ;
      RECT 0.2030 42.3765 0.2290 43.4700 ;
      RECT 0.0000 42.3765 0.0850 43.4700 ;
      RECT 0.0000 51.8040 9.6120 52.0965 ;
      RECT 9.5270 43.4430 9.6120 52.0965 ;
      RECT 4.5410 51.6555 9.6120 52.0965 ;
      RECT 0.0000 51.6555 4.3870 52.0965 ;
      RECT 5.9270 44.9470 9.4090 52.0965 ;
      RECT 7.3850 43.4430 9.4090 52.0965 ;
      RECT 4.5410 51.6290 5.8450 52.0965 ;
      RECT 5.1800 51.6280 5.8450 52.0965 ;
      RECT 3.7670 45.0550 4.3870 52.0965 ;
      RECT 3.8210 44.2090 4.3870 52.0965 ;
      RECT 0.2030 44.7520 3.6850 52.0965 ;
      RECT 3.3890 43.4430 3.6850 52.0965 ;
      RECT 0.0000 43.4430 0.0850 52.0965 ;
      RECT 4.5410 51.6260 5.0800 52.0965 ;
      RECT 5.0180 51.3550 5.0800 52.0965 ;
      RECT 5.1800 51.3550 5.7910 52.0965 ;
      RECT 4.5410 51.3550 4.9270 52.0965 ;
      RECT 5.9130 47.2360 9.4090 51.5960 ;
      RECT 0.2030 47.2360 3.6990 51.5960 ;
      RECT 5.9130 47.2360 9.4230 51.5915 ;
      RECT 0.1890 47.2360 3.6990 51.5915 ;
      RECT 5.1890 44.2090 5.7910 52.0965 ;
      RECT 4.7210 44.1280 4.8910 52.0965 ;
      RECT 4.8290 43.4430 4.8910 52.0965 ;
      RECT 4.0370 44.0270 4.4230 51.2050 ;
      RECT 3.7670 51.1630 4.4370 51.2000 ;
      RECT 5.1750 50.0890 5.7910 51.1970 ;
      RECT 4.7070 50.8990 4.8910 51.1250 ;
      RECT 4.7210 50.3230 4.9050 50.5850 ;
      RECT 3.7670 50.1250 4.4370 50.5850 ;
      RECT 4.7070 49.5850 4.8910 50.0450 ;
      RECT 5.1750 47.5510 5.7910 49.8830 ;
      RECT 3.7670 48.1990 4.4370 49.3430 ;
      RECT 4.7210 47.9290 4.9050 49.2350 ;
      RECT 4.7070 48.5050 4.9050 48.9650 ;
      RECT 4.7070 45.2650 4.8910 48.4250 ;
      RECT 4.7070 45.2650 4.9050 47.8850 ;
      RECT 3.7670 47.6590 4.4370 47.8850 ;
      RECT 5.2250 43.6195 5.8450 47.2040 ;
      RECT 5.1750 44.7250 5.8450 46.5110 ;
      RECT 3.7670 45.6970 4.4370 46.0670 ;
      RECT 4.7210 44.9950 4.9050 45.1850 ;
      RECT 3.8210 44.9590 4.4370 45.1490 ;
      RECT 4.7070 44.8510 4.8910 44.9870 ;
      RECT 4.7210 44.7250 4.9050 44.9510 ;
      RECT 6.0890 44.7550 9.4090 52.0965 ;
      RECT 7.1690 44.7520 9.4090 52.0965 ;
      RECT 5.9270 43.4430 6.0070 52.0965 ;
      RECT 3.7670 44.1280 3.9550 44.9420 ;
      RECT 5.9270 43.4430 6.2230 44.8460 ;
      RECT 5.9270 44.5600 7.0870 44.8460 ;
      RECT 7.1690 43.4430 7.3030 52.0965 ;
      RECT 2.5250 44.3710 3.3070 52.0965 ;
      RECT 0.2030 43.4430 2.4430 52.0965 ;
      RECT 5.9270 44.5600 7.3030 44.6540 ;
      RECT 6.9530 43.4430 9.4090 44.6510 ;
      RECT 3.1730 43.4430 3.6850 44.6510 ;
      RECT 4.7070 44.5810 4.9050 44.6450 ;
      RECT 4.7070 44.4550 4.8910 44.6450 ;
      RECT 6.7370 44.1760 9.4090 44.6510 ;
      RECT 5.9270 44.2090 6.6550 44.8460 ;
      RECT 4.7210 44.1850 4.9050 44.4470 ;
      RECT 0.2030 44.1760 3.0910 44.6510 ;
      RECT 2.9570 43.4430 3.0910 52.0965 ;
      RECT 6.5210 43.4430 6.8710 44.3150 ;
      RECT 5.9270 44.1280 6.4390 44.8460 ;
      RECT 6.3050 43.4430 6.4390 52.0965 ;
      RECT 2.7410 44.1280 3.0910 52.0965 ;
      RECT 0.2030 43.4430 2.6590 44.6510 ;
      RECT 4.7210 43.4430 4.7470 52.0965 ;
      RECT 3.8570 43.4430 3.9550 52.0965 ;
      RECT 2.7410 43.4430 2.8750 52.0965 ;
      RECT 6.3050 43.4430 6.8710 44.0780 ;
      RECT 5.1890 43.4430 5.7910 44.0780 ;
      RECT 3.8570 43.4430 4.3870 44.0780 ;
      RECT 2.9570 43.4430 3.6850 44.0780 ;
      RECT 6.3050 43.4430 9.4090 44.0750 ;
      RECT 0.2030 43.4430 2.8750 44.0750 ;
      RECT 5.1750 43.9150 5.8450 44.0690 ;
      RECT 3.8570 43.9150 4.4010 44.0780 ;
      RECT 5.9270 43.4430 9.4090 43.8110 ;
      RECT 4.7210 43.4430 4.8910 43.8110 ;
      RECT 3.7670 43.4430 4.3870 43.8110 ;
      RECT 0.2030 43.4430 3.6850 43.8110 ;
      RECT 4.5410 43.4430 4.8910 43.7080 ;
      RECT 5.1800 43.4430 5.7910 43.6080 ;
      RECT 4.5410 43.4430 4.9270 43.6080 ;
      RECT 5.1800 43.4430 5.8450 43.4640 ;
      RECT 6.3090 43.4165 6.3270 52.0965 ;
      RECT 6.2010 43.4165 6.2190 52.0965 ;
      RECT 2.9610 43.4165 2.9790 52.0965 ;
      RECT 2.8530 43.4165 2.8710 52.0965 ;
      RECT 5.0180 43.4430 5.0800 43.6080 ;
        RECT 5.1800 51.5835 5.3080 52.6770 ;
        RECT 5.1660 52.2490 5.3080 52.5715 ;
        RECT 5.0180 51.9760 5.0800 52.6770 ;
        RECT 5.0040 52.2855 5.0800 52.4390 ;
        RECT 5.0180 51.5835 5.0440 52.6770 ;
        RECT 5.0180 51.7045 5.0580 51.9440 ;
        RECT 5.0180 51.5835 5.0800 51.6725 ;
        RECT 4.7210 52.0340 4.9270 52.6770 ;
        RECT 4.9010 51.5835 4.9270 52.6770 ;
        RECT 4.7210 52.3110 4.9410 52.5690 ;
        RECT 4.7210 51.5835 4.8190 52.6770 ;
        RECT 4.3040 51.5835 4.3870 52.6770 ;
        RECT 4.3040 51.6720 4.4010 52.6075 ;
        RECT 9.5270 51.5835 9.6120 52.6770 ;
        RECT 9.3830 51.5835 9.4090 52.6770 ;
        RECT 9.2750 51.5835 9.3010 52.6770 ;
        RECT 9.1670 51.5835 9.1930 52.6770 ;
        RECT 9.0590 51.5835 9.0850 52.6770 ;
        RECT 8.9510 51.5835 8.9770 52.6770 ;
        RECT 8.8430 51.5835 8.8690 52.6770 ;
        RECT 8.7350 51.5835 8.7610 52.6770 ;
        RECT 8.6270 51.5835 8.6530 52.6770 ;
        RECT 8.5190 51.5835 8.5450 52.6770 ;
        RECT 8.4110 51.5835 8.4370 52.6770 ;
        RECT 8.3030 51.5835 8.3290 52.6770 ;
        RECT 8.1950 51.5835 8.2210 52.6770 ;
        RECT 8.0870 51.5835 8.1130 52.6770 ;
        RECT 7.9790 51.5835 8.0050 52.6770 ;
        RECT 7.8710 51.5835 7.8970 52.6770 ;
        RECT 7.7630 51.5835 7.7890 52.6770 ;
        RECT 7.6550 51.5835 7.6810 52.6770 ;
        RECT 7.5470 51.5835 7.5730 52.6770 ;
        RECT 7.4390 51.5835 7.4650 52.6770 ;
        RECT 7.3310 51.5835 7.3570 52.6770 ;
        RECT 7.2230 51.5835 7.2490 52.6770 ;
        RECT 7.1150 51.5835 7.1410 52.6770 ;
        RECT 7.0070 51.5835 7.0330 52.6770 ;
        RECT 6.8990 51.5835 6.9250 52.6770 ;
        RECT 6.7910 51.5835 6.8170 52.6770 ;
        RECT 6.6830 51.5835 6.7090 52.6770 ;
        RECT 6.5750 51.5835 6.6010 52.6770 ;
        RECT 6.4670 51.5835 6.4930 52.6770 ;
        RECT 6.3590 51.5835 6.3850 52.6770 ;
        RECT 6.2510 51.5835 6.2770 52.6770 ;
        RECT 6.1430 51.5835 6.1690 52.6770 ;
        RECT 6.0350 51.5835 6.0610 52.6770 ;
        RECT 5.9270 51.5835 5.9530 52.6770 ;
        RECT 5.7140 51.5835 5.7910 52.6770 ;
        RECT 3.8210 51.5835 3.8980 52.6770 ;
        RECT 3.6590 51.5835 3.6850 52.6770 ;
        RECT 3.5510 51.5835 3.5770 52.6770 ;
        RECT 3.4430 51.5835 3.4690 52.6770 ;
        RECT 3.3350 51.5835 3.3610 52.6770 ;
        RECT 3.2270 51.5835 3.2530 52.6770 ;
        RECT 3.1190 51.5835 3.1450 52.6770 ;
        RECT 3.0110 51.5835 3.0370 52.6770 ;
        RECT 2.9030 51.5835 2.9290 52.6770 ;
        RECT 2.7950 51.5835 2.8210 52.6770 ;
        RECT 2.6870 51.5835 2.7130 52.6770 ;
        RECT 2.5790 51.5835 2.6050 52.6770 ;
        RECT 2.4710 51.5835 2.4970 52.6770 ;
        RECT 2.3630 51.5835 2.3890 52.6770 ;
        RECT 2.2550 51.5835 2.2810 52.6770 ;
        RECT 2.1470 51.5835 2.1730 52.6770 ;
        RECT 2.0390 51.5835 2.0650 52.6770 ;
        RECT 1.9310 51.5835 1.9570 52.6770 ;
        RECT 1.8230 51.5835 1.8490 52.6770 ;
        RECT 1.7150 51.5835 1.7410 52.6770 ;
        RECT 1.6070 51.5835 1.6330 52.6770 ;
        RECT 1.4990 51.5835 1.5250 52.6770 ;
        RECT 1.3910 51.5835 1.4170 52.6770 ;
        RECT 1.2830 51.5835 1.3090 52.6770 ;
        RECT 1.1750 51.5835 1.2010 52.6770 ;
        RECT 1.0670 51.5835 1.0930 52.6770 ;
        RECT 0.9590 51.5835 0.9850 52.6770 ;
        RECT 0.8510 51.5835 0.8770 52.6770 ;
        RECT 0.7430 51.5835 0.7690 52.6770 ;
        RECT 0.6350 51.5835 0.6610 52.6770 ;
        RECT 0.5270 51.5835 0.5530 52.6770 ;
        RECT 0.4190 51.5835 0.4450 52.6770 ;
        RECT 0.3110 51.5835 0.3370 52.6770 ;
        RECT 0.2030 51.5835 0.2290 52.6770 ;
        RECT 0.0000 51.5835 0.0850 52.6770 ;
        RECT 5.1800 52.6635 5.3080 53.7570 ;
        RECT 5.1660 53.3290 5.3080 53.6515 ;
        RECT 5.0180 53.0560 5.0800 53.7570 ;
        RECT 5.0040 53.3655 5.0800 53.5190 ;
        RECT 5.0180 52.6635 5.0440 53.7570 ;
        RECT 5.0180 52.7845 5.0580 53.0240 ;
        RECT 5.0180 52.6635 5.0800 52.7525 ;
        RECT 4.7210 53.1140 4.9270 53.7570 ;
        RECT 4.9010 52.6635 4.9270 53.7570 ;
        RECT 4.7210 53.3910 4.9410 53.6490 ;
        RECT 4.7210 52.6635 4.8190 53.7570 ;
        RECT 4.3040 52.6635 4.3870 53.7570 ;
        RECT 4.3040 52.7520 4.4010 53.6875 ;
        RECT 9.5270 52.6635 9.6120 53.7570 ;
        RECT 9.3830 52.6635 9.4090 53.7570 ;
        RECT 9.2750 52.6635 9.3010 53.7570 ;
        RECT 9.1670 52.6635 9.1930 53.7570 ;
        RECT 9.0590 52.6635 9.0850 53.7570 ;
        RECT 8.9510 52.6635 8.9770 53.7570 ;
        RECT 8.8430 52.6635 8.8690 53.7570 ;
        RECT 8.7350 52.6635 8.7610 53.7570 ;
        RECT 8.6270 52.6635 8.6530 53.7570 ;
        RECT 8.5190 52.6635 8.5450 53.7570 ;
        RECT 8.4110 52.6635 8.4370 53.7570 ;
        RECT 8.3030 52.6635 8.3290 53.7570 ;
        RECT 8.1950 52.6635 8.2210 53.7570 ;
        RECT 8.0870 52.6635 8.1130 53.7570 ;
        RECT 7.9790 52.6635 8.0050 53.7570 ;
        RECT 7.8710 52.6635 7.8970 53.7570 ;
        RECT 7.7630 52.6635 7.7890 53.7570 ;
        RECT 7.6550 52.6635 7.6810 53.7570 ;
        RECT 7.5470 52.6635 7.5730 53.7570 ;
        RECT 7.4390 52.6635 7.4650 53.7570 ;
        RECT 7.3310 52.6635 7.3570 53.7570 ;
        RECT 7.2230 52.6635 7.2490 53.7570 ;
        RECT 7.1150 52.6635 7.1410 53.7570 ;
        RECT 7.0070 52.6635 7.0330 53.7570 ;
        RECT 6.8990 52.6635 6.9250 53.7570 ;
        RECT 6.7910 52.6635 6.8170 53.7570 ;
        RECT 6.6830 52.6635 6.7090 53.7570 ;
        RECT 6.5750 52.6635 6.6010 53.7570 ;
        RECT 6.4670 52.6635 6.4930 53.7570 ;
        RECT 6.3590 52.6635 6.3850 53.7570 ;
        RECT 6.2510 52.6635 6.2770 53.7570 ;
        RECT 6.1430 52.6635 6.1690 53.7570 ;
        RECT 6.0350 52.6635 6.0610 53.7570 ;
        RECT 5.9270 52.6635 5.9530 53.7570 ;
        RECT 5.7140 52.6635 5.7910 53.7570 ;
        RECT 3.8210 52.6635 3.8980 53.7570 ;
        RECT 3.6590 52.6635 3.6850 53.7570 ;
        RECT 3.5510 52.6635 3.5770 53.7570 ;
        RECT 3.4430 52.6635 3.4690 53.7570 ;
        RECT 3.3350 52.6635 3.3610 53.7570 ;
        RECT 3.2270 52.6635 3.2530 53.7570 ;
        RECT 3.1190 52.6635 3.1450 53.7570 ;
        RECT 3.0110 52.6635 3.0370 53.7570 ;
        RECT 2.9030 52.6635 2.9290 53.7570 ;
        RECT 2.7950 52.6635 2.8210 53.7570 ;
        RECT 2.6870 52.6635 2.7130 53.7570 ;
        RECT 2.5790 52.6635 2.6050 53.7570 ;
        RECT 2.4710 52.6635 2.4970 53.7570 ;
        RECT 2.3630 52.6635 2.3890 53.7570 ;
        RECT 2.2550 52.6635 2.2810 53.7570 ;
        RECT 2.1470 52.6635 2.1730 53.7570 ;
        RECT 2.0390 52.6635 2.0650 53.7570 ;
        RECT 1.9310 52.6635 1.9570 53.7570 ;
        RECT 1.8230 52.6635 1.8490 53.7570 ;
        RECT 1.7150 52.6635 1.7410 53.7570 ;
        RECT 1.6070 52.6635 1.6330 53.7570 ;
        RECT 1.4990 52.6635 1.5250 53.7570 ;
        RECT 1.3910 52.6635 1.4170 53.7570 ;
        RECT 1.2830 52.6635 1.3090 53.7570 ;
        RECT 1.1750 52.6635 1.2010 53.7570 ;
        RECT 1.0670 52.6635 1.0930 53.7570 ;
        RECT 0.9590 52.6635 0.9850 53.7570 ;
        RECT 0.8510 52.6635 0.8770 53.7570 ;
        RECT 0.7430 52.6635 0.7690 53.7570 ;
        RECT 0.6350 52.6635 0.6610 53.7570 ;
        RECT 0.5270 52.6635 0.5530 53.7570 ;
        RECT 0.4190 52.6635 0.4450 53.7570 ;
        RECT 0.3110 52.6635 0.3370 53.7570 ;
        RECT 0.2030 52.6635 0.2290 53.7570 ;
        RECT 0.0000 52.6635 0.0850 53.7570 ;
        RECT 5.1800 53.7435 5.3080 54.8370 ;
        RECT 5.1660 54.4090 5.3080 54.7315 ;
        RECT 5.0180 54.1360 5.0800 54.8370 ;
        RECT 5.0040 54.4455 5.0800 54.5990 ;
        RECT 5.0180 53.7435 5.0440 54.8370 ;
        RECT 5.0180 53.8645 5.0580 54.1040 ;
        RECT 5.0180 53.7435 5.0800 53.8325 ;
        RECT 4.7210 54.1940 4.9270 54.8370 ;
        RECT 4.9010 53.7435 4.9270 54.8370 ;
        RECT 4.7210 54.4710 4.9410 54.7290 ;
        RECT 4.7210 53.7435 4.8190 54.8370 ;
        RECT 4.3040 53.7435 4.3870 54.8370 ;
        RECT 4.3040 53.8320 4.4010 54.7675 ;
        RECT 9.5270 53.7435 9.6120 54.8370 ;
        RECT 9.3830 53.7435 9.4090 54.8370 ;
        RECT 9.2750 53.7435 9.3010 54.8370 ;
        RECT 9.1670 53.7435 9.1930 54.8370 ;
        RECT 9.0590 53.7435 9.0850 54.8370 ;
        RECT 8.9510 53.7435 8.9770 54.8370 ;
        RECT 8.8430 53.7435 8.8690 54.8370 ;
        RECT 8.7350 53.7435 8.7610 54.8370 ;
        RECT 8.6270 53.7435 8.6530 54.8370 ;
        RECT 8.5190 53.7435 8.5450 54.8370 ;
        RECT 8.4110 53.7435 8.4370 54.8370 ;
        RECT 8.3030 53.7435 8.3290 54.8370 ;
        RECT 8.1950 53.7435 8.2210 54.8370 ;
        RECT 8.0870 53.7435 8.1130 54.8370 ;
        RECT 7.9790 53.7435 8.0050 54.8370 ;
        RECT 7.8710 53.7435 7.8970 54.8370 ;
        RECT 7.7630 53.7435 7.7890 54.8370 ;
        RECT 7.6550 53.7435 7.6810 54.8370 ;
        RECT 7.5470 53.7435 7.5730 54.8370 ;
        RECT 7.4390 53.7435 7.4650 54.8370 ;
        RECT 7.3310 53.7435 7.3570 54.8370 ;
        RECT 7.2230 53.7435 7.2490 54.8370 ;
        RECT 7.1150 53.7435 7.1410 54.8370 ;
        RECT 7.0070 53.7435 7.0330 54.8370 ;
        RECT 6.8990 53.7435 6.9250 54.8370 ;
        RECT 6.7910 53.7435 6.8170 54.8370 ;
        RECT 6.6830 53.7435 6.7090 54.8370 ;
        RECT 6.5750 53.7435 6.6010 54.8370 ;
        RECT 6.4670 53.7435 6.4930 54.8370 ;
        RECT 6.3590 53.7435 6.3850 54.8370 ;
        RECT 6.2510 53.7435 6.2770 54.8370 ;
        RECT 6.1430 53.7435 6.1690 54.8370 ;
        RECT 6.0350 53.7435 6.0610 54.8370 ;
        RECT 5.9270 53.7435 5.9530 54.8370 ;
        RECT 5.7140 53.7435 5.7910 54.8370 ;
        RECT 3.8210 53.7435 3.8980 54.8370 ;
        RECT 3.6590 53.7435 3.6850 54.8370 ;
        RECT 3.5510 53.7435 3.5770 54.8370 ;
        RECT 3.4430 53.7435 3.4690 54.8370 ;
        RECT 3.3350 53.7435 3.3610 54.8370 ;
        RECT 3.2270 53.7435 3.2530 54.8370 ;
        RECT 3.1190 53.7435 3.1450 54.8370 ;
        RECT 3.0110 53.7435 3.0370 54.8370 ;
        RECT 2.9030 53.7435 2.9290 54.8370 ;
        RECT 2.7950 53.7435 2.8210 54.8370 ;
        RECT 2.6870 53.7435 2.7130 54.8370 ;
        RECT 2.5790 53.7435 2.6050 54.8370 ;
        RECT 2.4710 53.7435 2.4970 54.8370 ;
        RECT 2.3630 53.7435 2.3890 54.8370 ;
        RECT 2.2550 53.7435 2.2810 54.8370 ;
        RECT 2.1470 53.7435 2.1730 54.8370 ;
        RECT 2.0390 53.7435 2.0650 54.8370 ;
        RECT 1.9310 53.7435 1.9570 54.8370 ;
        RECT 1.8230 53.7435 1.8490 54.8370 ;
        RECT 1.7150 53.7435 1.7410 54.8370 ;
        RECT 1.6070 53.7435 1.6330 54.8370 ;
        RECT 1.4990 53.7435 1.5250 54.8370 ;
        RECT 1.3910 53.7435 1.4170 54.8370 ;
        RECT 1.2830 53.7435 1.3090 54.8370 ;
        RECT 1.1750 53.7435 1.2010 54.8370 ;
        RECT 1.0670 53.7435 1.0930 54.8370 ;
        RECT 0.9590 53.7435 0.9850 54.8370 ;
        RECT 0.8510 53.7435 0.8770 54.8370 ;
        RECT 0.7430 53.7435 0.7690 54.8370 ;
        RECT 0.6350 53.7435 0.6610 54.8370 ;
        RECT 0.5270 53.7435 0.5530 54.8370 ;
        RECT 0.4190 53.7435 0.4450 54.8370 ;
        RECT 0.3110 53.7435 0.3370 54.8370 ;
        RECT 0.2030 53.7435 0.2290 54.8370 ;
        RECT 0.0000 53.7435 0.0850 54.8370 ;
        RECT 5.1800 54.8235 5.3080 55.9170 ;
        RECT 5.1660 55.4890 5.3080 55.8115 ;
        RECT 5.0180 55.2160 5.0800 55.9170 ;
        RECT 5.0040 55.5255 5.0800 55.6790 ;
        RECT 5.0180 54.8235 5.0440 55.9170 ;
        RECT 5.0180 54.9445 5.0580 55.1840 ;
        RECT 5.0180 54.8235 5.0800 54.9125 ;
        RECT 4.7210 55.2740 4.9270 55.9170 ;
        RECT 4.9010 54.8235 4.9270 55.9170 ;
        RECT 4.7210 55.5510 4.9410 55.8090 ;
        RECT 4.7210 54.8235 4.8190 55.9170 ;
        RECT 4.3040 54.8235 4.3870 55.9170 ;
        RECT 4.3040 54.9120 4.4010 55.8475 ;
        RECT 9.5270 54.8235 9.6120 55.9170 ;
        RECT 9.3830 54.8235 9.4090 55.9170 ;
        RECT 9.2750 54.8235 9.3010 55.9170 ;
        RECT 9.1670 54.8235 9.1930 55.9170 ;
        RECT 9.0590 54.8235 9.0850 55.9170 ;
        RECT 8.9510 54.8235 8.9770 55.9170 ;
        RECT 8.8430 54.8235 8.8690 55.9170 ;
        RECT 8.7350 54.8235 8.7610 55.9170 ;
        RECT 8.6270 54.8235 8.6530 55.9170 ;
        RECT 8.5190 54.8235 8.5450 55.9170 ;
        RECT 8.4110 54.8235 8.4370 55.9170 ;
        RECT 8.3030 54.8235 8.3290 55.9170 ;
        RECT 8.1950 54.8235 8.2210 55.9170 ;
        RECT 8.0870 54.8235 8.1130 55.9170 ;
        RECT 7.9790 54.8235 8.0050 55.9170 ;
        RECT 7.8710 54.8235 7.8970 55.9170 ;
        RECT 7.7630 54.8235 7.7890 55.9170 ;
        RECT 7.6550 54.8235 7.6810 55.9170 ;
        RECT 7.5470 54.8235 7.5730 55.9170 ;
        RECT 7.4390 54.8235 7.4650 55.9170 ;
        RECT 7.3310 54.8235 7.3570 55.9170 ;
        RECT 7.2230 54.8235 7.2490 55.9170 ;
        RECT 7.1150 54.8235 7.1410 55.9170 ;
        RECT 7.0070 54.8235 7.0330 55.9170 ;
        RECT 6.8990 54.8235 6.9250 55.9170 ;
        RECT 6.7910 54.8235 6.8170 55.9170 ;
        RECT 6.6830 54.8235 6.7090 55.9170 ;
        RECT 6.5750 54.8235 6.6010 55.9170 ;
        RECT 6.4670 54.8235 6.4930 55.9170 ;
        RECT 6.3590 54.8235 6.3850 55.9170 ;
        RECT 6.2510 54.8235 6.2770 55.9170 ;
        RECT 6.1430 54.8235 6.1690 55.9170 ;
        RECT 6.0350 54.8235 6.0610 55.9170 ;
        RECT 5.9270 54.8235 5.9530 55.9170 ;
        RECT 5.7140 54.8235 5.7910 55.9170 ;
        RECT 3.8210 54.8235 3.8980 55.9170 ;
        RECT 3.6590 54.8235 3.6850 55.9170 ;
        RECT 3.5510 54.8235 3.5770 55.9170 ;
        RECT 3.4430 54.8235 3.4690 55.9170 ;
        RECT 3.3350 54.8235 3.3610 55.9170 ;
        RECT 3.2270 54.8235 3.2530 55.9170 ;
        RECT 3.1190 54.8235 3.1450 55.9170 ;
        RECT 3.0110 54.8235 3.0370 55.9170 ;
        RECT 2.9030 54.8235 2.9290 55.9170 ;
        RECT 2.7950 54.8235 2.8210 55.9170 ;
        RECT 2.6870 54.8235 2.7130 55.9170 ;
        RECT 2.5790 54.8235 2.6050 55.9170 ;
        RECT 2.4710 54.8235 2.4970 55.9170 ;
        RECT 2.3630 54.8235 2.3890 55.9170 ;
        RECT 2.2550 54.8235 2.2810 55.9170 ;
        RECT 2.1470 54.8235 2.1730 55.9170 ;
        RECT 2.0390 54.8235 2.0650 55.9170 ;
        RECT 1.9310 54.8235 1.9570 55.9170 ;
        RECT 1.8230 54.8235 1.8490 55.9170 ;
        RECT 1.7150 54.8235 1.7410 55.9170 ;
        RECT 1.6070 54.8235 1.6330 55.9170 ;
        RECT 1.4990 54.8235 1.5250 55.9170 ;
        RECT 1.3910 54.8235 1.4170 55.9170 ;
        RECT 1.2830 54.8235 1.3090 55.9170 ;
        RECT 1.1750 54.8235 1.2010 55.9170 ;
        RECT 1.0670 54.8235 1.0930 55.9170 ;
        RECT 0.9590 54.8235 0.9850 55.9170 ;
        RECT 0.8510 54.8235 0.8770 55.9170 ;
        RECT 0.7430 54.8235 0.7690 55.9170 ;
        RECT 0.6350 54.8235 0.6610 55.9170 ;
        RECT 0.5270 54.8235 0.5530 55.9170 ;
        RECT 0.4190 54.8235 0.4450 55.9170 ;
        RECT 0.3110 54.8235 0.3370 55.9170 ;
        RECT 0.2030 54.8235 0.2290 55.9170 ;
        RECT 0.0000 54.8235 0.0850 55.9170 ;
        RECT 5.1800 55.9035 5.3080 56.9970 ;
        RECT 5.1660 56.5690 5.3080 56.8915 ;
        RECT 5.0180 56.2960 5.0800 56.9970 ;
        RECT 5.0040 56.6055 5.0800 56.7590 ;
        RECT 5.0180 55.9035 5.0440 56.9970 ;
        RECT 5.0180 56.0245 5.0580 56.2640 ;
        RECT 5.0180 55.9035 5.0800 55.9925 ;
        RECT 4.7210 56.3540 4.9270 56.9970 ;
        RECT 4.9010 55.9035 4.9270 56.9970 ;
        RECT 4.7210 56.6310 4.9410 56.8890 ;
        RECT 4.7210 55.9035 4.8190 56.9970 ;
        RECT 4.3040 55.9035 4.3870 56.9970 ;
        RECT 4.3040 55.9920 4.4010 56.9275 ;
        RECT 9.5270 55.9035 9.6120 56.9970 ;
        RECT 9.3830 55.9035 9.4090 56.9970 ;
        RECT 9.2750 55.9035 9.3010 56.9970 ;
        RECT 9.1670 55.9035 9.1930 56.9970 ;
        RECT 9.0590 55.9035 9.0850 56.9970 ;
        RECT 8.9510 55.9035 8.9770 56.9970 ;
        RECT 8.8430 55.9035 8.8690 56.9970 ;
        RECT 8.7350 55.9035 8.7610 56.9970 ;
        RECT 8.6270 55.9035 8.6530 56.9970 ;
        RECT 8.5190 55.9035 8.5450 56.9970 ;
        RECT 8.4110 55.9035 8.4370 56.9970 ;
        RECT 8.3030 55.9035 8.3290 56.9970 ;
        RECT 8.1950 55.9035 8.2210 56.9970 ;
        RECT 8.0870 55.9035 8.1130 56.9970 ;
        RECT 7.9790 55.9035 8.0050 56.9970 ;
        RECT 7.8710 55.9035 7.8970 56.9970 ;
        RECT 7.7630 55.9035 7.7890 56.9970 ;
        RECT 7.6550 55.9035 7.6810 56.9970 ;
        RECT 7.5470 55.9035 7.5730 56.9970 ;
        RECT 7.4390 55.9035 7.4650 56.9970 ;
        RECT 7.3310 55.9035 7.3570 56.9970 ;
        RECT 7.2230 55.9035 7.2490 56.9970 ;
        RECT 7.1150 55.9035 7.1410 56.9970 ;
        RECT 7.0070 55.9035 7.0330 56.9970 ;
        RECT 6.8990 55.9035 6.9250 56.9970 ;
        RECT 6.7910 55.9035 6.8170 56.9970 ;
        RECT 6.6830 55.9035 6.7090 56.9970 ;
        RECT 6.5750 55.9035 6.6010 56.9970 ;
        RECT 6.4670 55.9035 6.4930 56.9970 ;
        RECT 6.3590 55.9035 6.3850 56.9970 ;
        RECT 6.2510 55.9035 6.2770 56.9970 ;
        RECT 6.1430 55.9035 6.1690 56.9970 ;
        RECT 6.0350 55.9035 6.0610 56.9970 ;
        RECT 5.9270 55.9035 5.9530 56.9970 ;
        RECT 5.7140 55.9035 5.7910 56.9970 ;
        RECT 3.8210 55.9035 3.8980 56.9970 ;
        RECT 3.6590 55.9035 3.6850 56.9970 ;
        RECT 3.5510 55.9035 3.5770 56.9970 ;
        RECT 3.4430 55.9035 3.4690 56.9970 ;
        RECT 3.3350 55.9035 3.3610 56.9970 ;
        RECT 3.2270 55.9035 3.2530 56.9970 ;
        RECT 3.1190 55.9035 3.1450 56.9970 ;
        RECT 3.0110 55.9035 3.0370 56.9970 ;
        RECT 2.9030 55.9035 2.9290 56.9970 ;
        RECT 2.7950 55.9035 2.8210 56.9970 ;
        RECT 2.6870 55.9035 2.7130 56.9970 ;
        RECT 2.5790 55.9035 2.6050 56.9970 ;
        RECT 2.4710 55.9035 2.4970 56.9970 ;
        RECT 2.3630 55.9035 2.3890 56.9970 ;
        RECT 2.2550 55.9035 2.2810 56.9970 ;
        RECT 2.1470 55.9035 2.1730 56.9970 ;
        RECT 2.0390 55.9035 2.0650 56.9970 ;
        RECT 1.9310 55.9035 1.9570 56.9970 ;
        RECT 1.8230 55.9035 1.8490 56.9970 ;
        RECT 1.7150 55.9035 1.7410 56.9970 ;
        RECT 1.6070 55.9035 1.6330 56.9970 ;
        RECT 1.4990 55.9035 1.5250 56.9970 ;
        RECT 1.3910 55.9035 1.4170 56.9970 ;
        RECT 1.2830 55.9035 1.3090 56.9970 ;
        RECT 1.1750 55.9035 1.2010 56.9970 ;
        RECT 1.0670 55.9035 1.0930 56.9970 ;
        RECT 0.9590 55.9035 0.9850 56.9970 ;
        RECT 0.8510 55.9035 0.8770 56.9970 ;
        RECT 0.7430 55.9035 0.7690 56.9970 ;
        RECT 0.6350 55.9035 0.6610 56.9970 ;
        RECT 0.5270 55.9035 0.5530 56.9970 ;
        RECT 0.4190 55.9035 0.4450 56.9970 ;
        RECT 0.3110 55.9035 0.3370 56.9970 ;
        RECT 0.2030 55.9035 0.2290 56.9970 ;
        RECT 0.0000 55.9035 0.0850 56.9970 ;
        RECT 5.1800 56.9835 5.3080 58.0770 ;
        RECT 5.1660 57.6490 5.3080 57.9715 ;
        RECT 5.0180 57.3760 5.0800 58.0770 ;
        RECT 5.0040 57.6855 5.0800 57.8390 ;
        RECT 5.0180 56.9835 5.0440 58.0770 ;
        RECT 5.0180 57.1045 5.0580 57.3440 ;
        RECT 5.0180 56.9835 5.0800 57.0725 ;
        RECT 4.7210 57.4340 4.9270 58.0770 ;
        RECT 4.9010 56.9835 4.9270 58.0770 ;
        RECT 4.7210 57.7110 4.9410 57.9690 ;
        RECT 4.7210 56.9835 4.8190 58.0770 ;
        RECT 4.3040 56.9835 4.3870 58.0770 ;
        RECT 4.3040 57.0720 4.4010 58.0075 ;
        RECT 9.5270 56.9835 9.6120 58.0770 ;
        RECT 9.3830 56.9835 9.4090 58.0770 ;
        RECT 9.2750 56.9835 9.3010 58.0770 ;
        RECT 9.1670 56.9835 9.1930 58.0770 ;
        RECT 9.0590 56.9835 9.0850 58.0770 ;
        RECT 8.9510 56.9835 8.9770 58.0770 ;
        RECT 8.8430 56.9835 8.8690 58.0770 ;
        RECT 8.7350 56.9835 8.7610 58.0770 ;
        RECT 8.6270 56.9835 8.6530 58.0770 ;
        RECT 8.5190 56.9835 8.5450 58.0770 ;
        RECT 8.4110 56.9835 8.4370 58.0770 ;
        RECT 8.3030 56.9835 8.3290 58.0770 ;
        RECT 8.1950 56.9835 8.2210 58.0770 ;
        RECT 8.0870 56.9835 8.1130 58.0770 ;
        RECT 7.9790 56.9835 8.0050 58.0770 ;
        RECT 7.8710 56.9835 7.8970 58.0770 ;
        RECT 7.7630 56.9835 7.7890 58.0770 ;
        RECT 7.6550 56.9835 7.6810 58.0770 ;
        RECT 7.5470 56.9835 7.5730 58.0770 ;
        RECT 7.4390 56.9835 7.4650 58.0770 ;
        RECT 7.3310 56.9835 7.3570 58.0770 ;
        RECT 7.2230 56.9835 7.2490 58.0770 ;
        RECT 7.1150 56.9835 7.1410 58.0770 ;
        RECT 7.0070 56.9835 7.0330 58.0770 ;
        RECT 6.8990 56.9835 6.9250 58.0770 ;
        RECT 6.7910 56.9835 6.8170 58.0770 ;
        RECT 6.6830 56.9835 6.7090 58.0770 ;
        RECT 6.5750 56.9835 6.6010 58.0770 ;
        RECT 6.4670 56.9835 6.4930 58.0770 ;
        RECT 6.3590 56.9835 6.3850 58.0770 ;
        RECT 6.2510 56.9835 6.2770 58.0770 ;
        RECT 6.1430 56.9835 6.1690 58.0770 ;
        RECT 6.0350 56.9835 6.0610 58.0770 ;
        RECT 5.9270 56.9835 5.9530 58.0770 ;
        RECT 5.7140 56.9835 5.7910 58.0770 ;
        RECT 3.8210 56.9835 3.8980 58.0770 ;
        RECT 3.6590 56.9835 3.6850 58.0770 ;
        RECT 3.5510 56.9835 3.5770 58.0770 ;
        RECT 3.4430 56.9835 3.4690 58.0770 ;
        RECT 3.3350 56.9835 3.3610 58.0770 ;
        RECT 3.2270 56.9835 3.2530 58.0770 ;
        RECT 3.1190 56.9835 3.1450 58.0770 ;
        RECT 3.0110 56.9835 3.0370 58.0770 ;
        RECT 2.9030 56.9835 2.9290 58.0770 ;
        RECT 2.7950 56.9835 2.8210 58.0770 ;
        RECT 2.6870 56.9835 2.7130 58.0770 ;
        RECT 2.5790 56.9835 2.6050 58.0770 ;
        RECT 2.4710 56.9835 2.4970 58.0770 ;
        RECT 2.3630 56.9835 2.3890 58.0770 ;
        RECT 2.2550 56.9835 2.2810 58.0770 ;
        RECT 2.1470 56.9835 2.1730 58.0770 ;
        RECT 2.0390 56.9835 2.0650 58.0770 ;
        RECT 1.9310 56.9835 1.9570 58.0770 ;
        RECT 1.8230 56.9835 1.8490 58.0770 ;
        RECT 1.7150 56.9835 1.7410 58.0770 ;
        RECT 1.6070 56.9835 1.6330 58.0770 ;
        RECT 1.4990 56.9835 1.5250 58.0770 ;
        RECT 1.3910 56.9835 1.4170 58.0770 ;
        RECT 1.2830 56.9835 1.3090 58.0770 ;
        RECT 1.1750 56.9835 1.2010 58.0770 ;
        RECT 1.0670 56.9835 1.0930 58.0770 ;
        RECT 0.9590 56.9835 0.9850 58.0770 ;
        RECT 0.8510 56.9835 0.8770 58.0770 ;
        RECT 0.7430 56.9835 0.7690 58.0770 ;
        RECT 0.6350 56.9835 0.6610 58.0770 ;
        RECT 0.5270 56.9835 0.5530 58.0770 ;
        RECT 0.4190 56.9835 0.4450 58.0770 ;
        RECT 0.3110 56.9835 0.3370 58.0770 ;
        RECT 0.2030 56.9835 0.2290 58.0770 ;
        RECT 0.0000 56.9835 0.0850 58.0770 ;
        RECT 5.1800 58.0635 5.3080 59.1570 ;
        RECT 5.1660 58.7290 5.3080 59.0515 ;
        RECT 5.0180 58.4560 5.0800 59.1570 ;
        RECT 5.0040 58.7655 5.0800 58.9190 ;
        RECT 5.0180 58.0635 5.0440 59.1570 ;
        RECT 5.0180 58.1845 5.0580 58.4240 ;
        RECT 5.0180 58.0635 5.0800 58.1525 ;
        RECT 4.7210 58.5140 4.9270 59.1570 ;
        RECT 4.9010 58.0635 4.9270 59.1570 ;
        RECT 4.7210 58.7910 4.9410 59.0490 ;
        RECT 4.7210 58.0635 4.8190 59.1570 ;
        RECT 4.3040 58.0635 4.3870 59.1570 ;
        RECT 4.3040 58.1520 4.4010 59.0875 ;
        RECT 9.5270 58.0635 9.6120 59.1570 ;
        RECT 9.3830 58.0635 9.4090 59.1570 ;
        RECT 9.2750 58.0635 9.3010 59.1570 ;
        RECT 9.1670 58.0635 9.1930 59.1570 ;
        RECT 9.0590 58.0635 9.0850 59.1570 ;
        RECT 8.9510 58.0635 8.9770 59.1570 ;
        RECT 8.8430 58.0635 8.8690 59.1570 ;
        RECT 8.7350 58.0635 8.7610 59.1570 ;
        RECT 8.6270 58.0635 8.6530 59.1570 ;
        RECT 8.5190 58.0635 8.5450 59.1570 ;
        RECT 8.4110 58.0635 8.4370 59.1570 ;
        RECT 8.3030 58.0635 8.3290 59.1570 ;
        RECT 8.1950 58.0635 8.2210 59.1570 ;
        RECT 8.0870 58.0635 8.1130 59.1570 ;
        RECT 7.9790 58.0635 8.0050 59.1570 ;
        RECT 7.8710 58.0635 7.8970 59.1570 ;
        RECT 7.7630 58.0635 7.7890 59.1570 ;
        RECT 7.6550 58.0635 7.6810 59.1570 ;
        RECT 7.5470 58.0635 7.5730 59.1570 ;
        RECT 7.4390 58.0635 7.4650 59.1570 ;
        RECT 7.3310 58.0635 7.3570 59.1570 ;
        RECT 7.2230 58.0635 7.2490 59.1570 ;
        RECT 7.1150 58.0635 7.1410 59.1570 ;
        RECT 7.0070 58.0635 7.0330 59.1570 ;
        RECT 6.8990 58.0635 6.9250 59.1570 ;
        RECT 6.7910 58.0635 6.8170 59.1570 ;
        RECT 6.6830 58.0635 6.7090 59.1570 ;
        RECT 6.5750 58.0635 6.6010 59.1570 ;
        RECT 6.4670 58.0635 6.4930 59.1570 ;
        RECT 6.3590 58.0635 6.3850 59.1570 ;
        RECT 6.2510 58.0635 6.2770 59.1570 ;
        RECT 6.1430 58.0635 6.1690 59.1570 ;
        RECT 6.0350 58.0635 6.0610 59.1570 ;
        RECT 5.9270 58.0635 5.9530 59.1570 ;
        RECT 5.7140 58.0635 5.7910 59.1570 ;
        RECT 3.8210 58.0635 3.8980 59.1570 ;
        RECT 3.6590 58.0635 3.6850 59.1570 ;
        RECT 3.5510 58.0635 3.5770 59.1570 ;
        RECT 3.4430 58.0635 3.4690 59.1570 ;
        RECT 3.3350 58.0635 3.3610 59.1570 ;
        RECT 3.2270 58.0635 3.2530 59.1570 ;
        RECT 3.1190 58.0635 3.1450 59.1570 ;
        RECT 3.0110 58.0635 3.0370 59.1570 ;
        RECT 2.9030 58.0635 2.9290 59.1570 ;
        RECT 2.7950 58.0635 2.8210 59.1570 ;
        RECT 2.6870 58.0635 2.7130 59.1570 ;
        RECT 2.5790 58.0635 2.6050 59.1570 ;
        RECT 2.4710 58.0635 2.4970 59.1570 ;
        RECT 2.3630 58.0635 2.3890 59.1570 ;
        RECT 2.2550 58.0635 2.2810 59.1570 ;
        RECT 2.1470 58.0635 2.1730 59.1570 ;
        RECT 2.0390 58.0635 2.0650 59.1570 ;
        RECT 1.9310 58.0635 1.9570 59.1570 ;
        RECT 1.8230 58.0635 1.8490 59.1570 ;
        RECT 1.7150 58.0635 1.7410 59.1570 ;
        RECT 1.6070 58.0635 1.6330 59.1570 ;
        RECT 1.4990 58.0635 1.5250 59.1570 ;
        RECT 1.3910 58.0635 1.4170 59.1570 ;
        RECT 1.2830 58.0635 1.3090 59.1570 ;
        RECT 1.1750 58.0635 1.2010 59.1570 ;
        RECT 1.0670 58.0635 1.0930 59.1570 ;
        RECT 0.9590 58.0635 0.9850 59.1570 ;
        RECT 0.8510 58.0635 0.8770 59.1570 ;
        RECT 0.7430 58.0635 0.7690 59.1570 ;
        RECT 0.6350 58.0635 0.6610 59.1570 ;
        RECT 0.5270 58.0635 0.5530 59.1570 ;
        RECT 0.4190 58.0635 0.4450 59.1570 ;
        RECT 0.3110 58.0635 0.3370 59.1570 ;
        RECT 0.2030 58.0635 0.2290 59.1570 ;
        RECT 0.0000 58.0635 0.0850 59.1570 ;
        RECT 5.1800 59.1435 5.3080 60.2370 ;
        RECT 5.1660 59.8090 5.3080 60.1315 ;
        RECT 5.0180 59.5360 5.0800 60.2370 ;
        RECT 5.0040 59.8455 5.0800 59.9990 ;
        RECT 5.0180 59.1435 5.0440 60.2370 ;
        RECT 5.0180 59.2645 5.0580 59.5040 ;
        RECT 5.0180 59.1435 5.0800 59.2325 ;
        RECT 4.7210 59.5940 4.9270 60.2370 ;
        RECT 4.9010 59.1435 4.9270 60.2370 ;
        RECT 4.7210 59.8710 4.9410 60.1290 ;
        RECT 4.7210 59.1435 4.8190 60.2370 ;
        RECT 4.3040 59.1435 4.3870 60.2370 ;
        RECT 4.3040 59.2320 4.4010 60.1675 ;
        RECT 9.5270 59.1435 9.6120 60.2370 ;
        RECT 9.3830 59.1435 9.4090 60.2370 ;
        RECT 9.2750 59.1435 9.3010 60.2370 ;
        RECT 9.1670 59.1435 9.1930 60.2370 ;
        RECT 9.0590 59.1435 9.0850 60.2370 ;
        RECT 8.9510 59.1435 8.9770 60.2370 ;
        RECT 8.8430 59.1435 8.8690 60.2370 ;
        RECT 8.7350 59.1435 8.7610 60.2370 ;
        RECT 8.6270 59.1435 8.6530 60.2370 ;
        RECT 8.5190 59.1435 8.5450 60.2370 ;
        RECT 8.4110 59.1435 8.4370 60.2370 ;
        RECT 8.3030 59.1435 8.3290 60.2370 ;
        RECT 8.1950 59.1435 8.2210 60.2370 ;
        RECT 8.0870 59.1435 8.1130 60.2370 ;
        RECT 7.9790 59.1435 8.0050 60.2370 ;
        RECT 7.8710 59.1435 7.8970 60.2370 ;
        RECT 7.7630 59.1435 7.7890 60.2370 ;
        RECT 7.6550 59.1435 7.6810 60.2370 ;
        RECT 7.5470 59.1435 7.5730 60.2370 ;
        RECT 7.4390 59.1435 7.4650 60.2370 ;
        RECT 7.3310 59.1435 7.3570 60.2370 ;
        RECT 7.2230 59.1435 7.2490 60.2370 ;
        RECT 7.1150 59.1435 7.1410 60.2370 ;
        RECT 7.0070 59.1435 7.0330 60.2370 ;
        RECT 6.8990 59.1435 6.9250 60.2370 ;
        RECT 6.7910 59.1435 6.8170 60.2370 ;
        RECT 6.6830 59.1435 6.7090 60.2370 ;
        RECT 6.5750 59.1435 6.6010 60.2370 ;
        RECT 6.4670 59.1435 6.4930 60.2370 ;
        RECT 6.3590 59.1435 6.3850 60.2370 ;
        RECT 6.2510 59.1435 6.2770 60.2370 ;
        RECT 6.1430 59.1435 6.1690 60.2370 ;
        RECT 6.0350 59.1435 6.0610 60.2370 ;
        RECT 5.9270 59.1435 5.9530 60.2370 ;
        RECT 5.7140 59.1435 5.7910 60.2370 ;
        RECT 3.8210 59.1435 3.8980 60.2370 ;
        RECT 3.6590 59.1435 3.6850 60.2370 ;
        RECT 3.5510 59.1435 3.5770 60.2370 ;
        RECT 3.4430 59.1435 3.4690 60.2370 ;
        RECT 3.3350 59.1435 3.3610 60.2370 ;
        RECT 3.2270 59.1435 3.2530 60.2370 ;
        RECT 3.1190 59.1435 3.1450 60.2370 ;
        RECT 3.0110 59.1435 3.0370 60.2370 ;
        RECT 2.9030 59.1435 2.9290 60.2370 ;
        RECT 2.7950 59.1435 2.8210 60.2370 ;
        RECT 2.6870 59.1435 2.7130 60.2370 ;
        RECT 2.5790 59.1435 2.6050 60.2370 ;
        RECT 2.4710 59.1435 2.4970 60.2370 ;
        RECT 2.3630 59.1435 2.3890 60.2370 ;
        RECT 2.2550 59.1435 2.2810 60.2370 ;
        RECT 2.1470 59.1435 2.1730 60.2370 ;
        RECT 2.0390 59.1435 2.0650 60.2370 ;
        RECT 1.9310 59.1435 1.9570 60.2370 ;
        RECT 1.8230 59.1435 1.8490 60.2370 ;
        RECT 1.7150 59.1435 1.7410 60.2370 ;
        RECT 1.6070 59.1435 1.6330 60.2370 ;
        RECT 1.4990 59.1435 1.5250 60.2370 ;
        RECT 1.3910 59.1435 1.4170 60.2370 ;
        RECT 1.2830 59.1435 1.3090 60.2370 ;
        RECT 1.1750 59.1435 1.2010 60.2370 ;
        RECT 1.0670 59.1435 1.0930 60.2370 ;
        RECT 0.9590 59.1435 0.9850 60.2370 ;
        RECT 0.8510 59.1435 0.8770 60.2370 ;
        RECT 0.7430 59.1435 0.7690 60.2370 ;
        RECT 0.6350 59.1435 0.6610 60.2370 ;
        RECT 0.5270 59.1435 0.5530 60.2370 ;
        RECT 0.4190 59.1435 0.4450 60.2370 ;
        RECT 0.3110 59.1435 0.3370 60.2370 ;
        RECT 0.2030 59.1435 0.2290 60.2370 ;
        RECT 0.0000 59.1435 0.0850 60.2370 ;
        RECT 5.1800 60.2235 5.3080 61.3170 ;
        RECT 5.1660 60.8890 5.3080 61.2115 ;
        RECT 5.0180 60.6160 5.0800 61.3170 ;
        RECT 5.0040 60.9255 5.0800 61.0790 ;
        RECT 5.0180 60.2235 5.0440 61.3170 ;
        RECT 5.0180 60.3445 5.0580 60.5840 ;
        RECT 5.0180 60.2235 5.0800 60.3125 ;
        RECT 4.7210 60.6740 4.9270 61.3170 ;
        RECT 4.9010 60.2235 4.9270 61.3170 ;
        RECT 4.7210 60.9510 4.9410 61.2090 ;
        RECT 4.7210 60.2235 4.8190 61.3170 ;
        RECT 4.3040 60.2235 4.3870 61.3170 ;
        RECT 4.3040 60.3120 4.4010 61.2475 ;
        RECT 9.5270 60.2235 9.6120 61.3170 ;
        RECT 9.3830 60.2235 9.4090 61.3170 ;
        RECT 9.2750 60.2235 9.3010 61.3170 ;
        RECT 9.1670 60.2235 9.1930 61.3170 ;
        RECT 9.0590 60.2235 9.0850 61.3170 ;
        RECT 8.9510 60.2235 8.9770 61.3170 ;
        RECT 8.8430 60.2235 8.8690 61.3170 ;
        RECT 8.7350 60.2235 8.7610 61.3170 ;
        RECT 8.6270 60.2235 8.6530 61.3170 ;
        RECT 8.5190 60.2235 8.5450 61.3170 ;
        RECT 8.4110 60.2235 8.4370 61.3170 ;
        RECT 8.3030 60.2235 8.3290 61.3170 ;
        RECT 8.1950 60.2235 8.2210 61.3170 ;
        RECT 8.0870 60.2235 8.1130 61.3170 ;
        RECT 7.9790 60.2235 8.0050 61.3170 ;
        RECT 7.8710 60.2235 7.8970 61.3170 ;
        RECT 7.7630 60.2235 7.7890 61.3170 ;
        RECT 7.6550 60.2235 7.6810 61.3170 ;
        RECT 7.5470 60.2235 7.5730 61.3170 ;
        RECT 7.4390 60.2235 7.4650 61.3170 ;
        RECT 7.3310 60.2235 7.3570 61.3170 ;
        RECT 7.2230 60.2235 7.2490 61.3170 ;
        RECT 7.1150 60.2235 7.1410 61.3170 ;
        RECT 7.0070 60.2235 7.0330 61.3170 ;
        RECT 6.8990 60.2235 6.9250 61.3170 ;
        RECT 6.7910 60.2235 6.8170 61.3170 ;
        RECT 6.6830 60.2235 6.7090 61.3170 ;
        RECT 6.5750 60.2235 6.6010 61.3170 ;
        RECT 6.4670 60.2235 6.4930 61.3170 ;
        RECT 6.3590 60.2235 6.3850 61.3170 ;
        RECT 6.2510 60.2235 6.2770 61.3170 ;
        RECT 6.1430 60.2235 6.1690 61.3170 ;
        RECT 6.0350 60.2235 6.0610 61.3170 ;
        RECT 5.9270 60.2235 5.9530 61.3170 ;
        RECT 5.7140 60.2235 5.7910 61.3170 ;
        RECT 3.8210 60.2235 3.8980 61.3170 ;
        RECT 3.6590 60.2235 3.6850 61.3170 ;
        RECT 3.5510 60.2235 3.5770 61.3170 ;
        RECT 3.4430 60.2235 3.4690 61.3170 ;
        RECT 3.3350 60.2235 3.3610 61.3170 ;
        RECT 3.2270 60.2235 3.2530 61.3170 ;
        RECT 3.1190 60.2235 3.1450 61.3170 ;
        RECT 3.0110 60.2235 3.0370 61.3170 ;
        RECT 2.9030 60.2235 2.9290 61.3170 ;
        RECT 2.7950 60.2235 2.8210 61.3170 ;
        RECT 2.6870 60.2235 2.7130 61.3170 ;
        RECT 2.5790 60.2235 2.6050 61.3170 ;
        RECT 2.4710 60.2235 2.4970 61.3170 ;
        RECT 2.3630 60.2235 2.3890 61.3170 ;
        RECT 2.2550 60.2235 2.2810 61.3170 ;
        RECT 2.1470 60.2235 2.1730 61.3170 ;
        RECT 2.0390 60.2235 2.0650 61.3170 ;
        RECT 1.9310 60.2235 1.9570 61.3170 ;
        RECT 1.8230 60.2235 1.8490 61.3170 ;
        RECT 1.7150 60.2235 1.7410 61.3170 ;
        RECT 1.6070 60.2235 1.6330 61.3170 ;
        RECT 1.4990 60.2235 1.5250 61.3170 ;
        RECT 1.3910 60.2235 1.4170 61.3170 ;
        RECT 1.2830 60.2235 1.3090 61.3170 ;
        RECT 1.1750 60.2235 1.2010 61.3170 ;
        RECT 1.0670 60.2235 1.0930 61.3170 ;
        RECT 0.9590 60.2235 0.9850 61.3170 ;
        RECT 0.8510 60.2235 0.8770 61.3170 ;
        RECT 0.7430 60.2235 0.7690 61.3170 ;
        RECT 0.6350 60.2235 0.6610 61.3170 ;
        RECT 0.5270 60.2235 0.5530 61.3170 ;
        RECT 0.4190 60.2235 0.4450 61.3170 ;
        RECT 0.3110 60.2235 0.3370 61.3170 ;
        RECT 0.2030 60.2235 0.2290 61.3170 ;
        RECT 0.0000 60.2235 0.0850 61.3170 ;
        RECT 5.1800 61.3035 5.3080 62.3970 ;
        RECT 5.1660 61.9690 5.3080 62.2915 ;
        RECT 5.0180 61.6960 5.0800 62.3970 ;
        RECT 5.0040 62.0055 5.0800 62.1590 ;
        RECT 5.0180 61.3035 5.0440 62.3970 ;
        RECT 5.0180 61.4245 5.0580 61.6640 ;
        RECT 5.0180 61.3035 5.0800 61.3925 ;
        RECT 4.7210 61.7540 4.9270 62.3970 ;
        RECT 4.9010 61.3035 4.9270 62.3970 ;
        RECT 4.7210 62.0310 4.9410 62.2890 ;
        RECT 4.7210 61.3035 4.8190 62.3970 ;
        RECT 4.3040 61.3035 4.3870 62.3970 ;
        RECT 4.3040 61.3920 4.4010 62.3275 ;
        RECT 9.5270 61.3035 9.6120 62.3970 ;
        RECT 9.3830 61.3035 9.4090 62.3970 ;
        RECT 9.2750 61.3035 9.3010 62.3970 ;
        RECT 9.1670 61.3035 9.1930 62.3970 ;
        RECT 9.0590 61.3035 9.0850 62.3970 ;
        RECT 8.9510 61.3035 8.9770 62.3970 ;
        RECT 8.8430 61.3035 8.8690 62.3970 ;
        RECT 8.7350 61.3035 8.7610 62.3970 ;
        RECT 8.6270 61.3035 8.6530 62.3970 ;
        RECT 8.5190 61.3035 8.5450 62.3970 ;
        RECT 8.4110 61.3035 8.4370 62.3970 ;
        RECT 8.3030 61.3035 8.3290 62.3970 ;
        RECT 8.1950 61.3035 8.2210 62.3970 ;
        RECT 8.0870 61.3035 8.1130 62.3970 ;
        RECT 7.9790 61.3035 8.0050 62.3970 ;
        RECT 7.8710 61.3035 7.8970 62.3970 ;
        RECT 7.7630 61.3035 7.7890 62.3970 ;
        RECT 7.6550 61.3035 7.6810 62.3970 ;
        RECT 7.5470 61.3035 7.5730 62.3970 ;
        RECT 7.4390 61.3035 7.4650 62.3970 ;
        RECT 7.3310 61.3035 7.3570 62.3970 ;
        RECT 7.2230 61.3035 7.2490 62.3970 ;
        RECT 7.1150 61.3035 7.1410 62.3970 ;
        RECT 7.0070 61.3035 7.0330 62.3970 ;
        RECT 6.8990 61.3035 6.9250 62.3970 ;
        RECT 6.7910 61.3035 6.8170 62.3970 ;
        RECT 6.6830 61.3035 6.7090 62.3970 ;
        RECT 6.5750 61.3035 6.6010 62.3970 ;
        RECT 6.4670 61.3035 6.4930 62.3970 ;
        RECT 6.3590 61.3035 6.3850 62.3970 ;
        RECT 6.2510 61.3035 6.2770 62.3970 ;
        RECT 6.1430 61.3035 6.1690 62.3970 ;
        RECT 6.0350 61.3035 6.0610 62.3970 ;
        RECT 5.9270 61.3035 5.9530 62.3970 ;
        RECT 5.7140 61.3035 5.7910 62.3970 ;
        RECT 3.8210 61.3035 3.8980 62.3970 ;
        RECT 3.6590 61.3035 3.6850 62.3970 ;
        RECT 3.5510 61.3035 3.5770 62.3970 ;
        RECT 3.4430 61.3035 3.4690 62.3970 ;
        RECT 3.3350 61.3035 3.3610 62.3970 ;
        RECT 3.2270 61.3035 3.2530 62.3970 ;
        RECT 3.1190 61.3035 3.1450 62.3970 ;
        RECT 3.0110 61.3035 3.0370 62.3970 ;
        RECT 2.9030 61.3035 2.9290 62.3970 ;
        RECT 2.7950 61.3035 2.8210 62.3970 ;
        RECT 2.6870 61.3035 2.7130 62.3970 ;
        RECT 2.5790 61.3035 2.6050 62.3970 ;
        RECT 2.4710 61.3035 2.4970 62.3970 ;
        RECT 2.3630 61.3035 2.3890 62.3970 ;
        RECT 2.2550 61.3035 2.2810 62.3970 ;
        RECT 2.1470 61.3035 2.1730 62.3970 ;
        RECT 2.0390 61.3035 2.0650 62.3970 ;
        RECT 1.9310 61.3035 1.9570 62.3970 ;
        RECT 1.8230 61.3035 1.8490 62.3970 ;
        RECT 1.7150 61.3035 1.7410 62.3970 ;
        RECT 1.6070 61.3035 1.6330 62.3970 ;
        RECT 1.4990 61.3035 1.5250 62.3970 ;
        RECT 1.3910 61.3035 1.4170 62.3970 ;
        RECT 1.2830 61.3035 1.3090 62.3970 ;
        RECT 1.1750 61.3035 1.2010 62.3970 ;
        RECT 1.0670 61.3035 1.0930 62.3970 ;
        RECT 0.9590 61.3035 0.9850 62.3970 ;
        RECT 0.8510 61.3035 0.8770 62.3970 ;
        RECT 0.7430 61.3035 0.7690 62.3970 ;
        RECT 0.6350 61.3035 0.6610 62.3970 ;
        RECT 0.5270 61.3035 0.5530 62.3970 ;
        RECT 0.4190 61.3035 0.4450 62.3970 ;
        RECT 0.3110 61.3035 0.3370 62.3970 ;
        RECT 0.2030 61.3035 0.2290 62.3970 ;
        RECT 0.0000 61.3035 0.0850 62.3970 ;
        RECT 5.1800 62.3835 5.3080 63.4770 ;
        RECT 5.1660 63.0490 5.3080 63.3715 ;
        RECT 5.0180 62.7760 5.0800 63.4770 ;
        RECT 5.0040 63.0855 5.0800 63.2390 ;
        RECT 5.0180 62.3835 5.0440 63.4770 ;
        RECT 5.0180 62.5045 5.0580 62.7440 ;
        RECT 5.0180 62.3835 5.0800 62.4725 ;
        RECT 4.7210 62.8340 4.9270 63.4770 ;
        RECT 4.9010 62.3835 4.9270 63.4770 ;
        RECT 4.7210 63.1110 4.9410 63.3690 ;
        RECT 4.7210 62.3835 4.8190 63.4770 ;
        RECT 4.3040 62.3835 4.3870 63.4770 ;
        RECT 4.3040 62.4720 4.4010 63.4075 ;
        RECT 9.5270 62.3835 9.6120 63.4770 ;
        RECT 9.3830 62.3835 9.4090 63.4770 ;
        RECT 9.2750 62.3835 9.3010 63.4770 ;
        RECT 9.1670 62.3835 9.1930 63.4770 ;
        RECT 9.0590 62.3835 9.0850 63.4770 ;
        RECT 8.9510 62.3835 8.9770 63.4770 ;
        RECT 8.8430 62.3835 8.8690 63.4770 ;
        RECT 8.7350 62.3835 8.7610 63.4770 ;
        RECT 8.6270 62.3835 8.6530 63.4770 ;
        RECT 8.5190 62.3835 8.5450 63.4770 ;
        RECT 8.4110 62.3835 8.4370 63.4770 ;
        RECT 8.3030 62.3835 8.3290 63.4770 ;
        RECT 8.1950 62.3835 8.2210 63.4770 ;
        RECT 8.0870 62.3835 8.1130 63.4770 ;
        RECT 7.9790 62.3835 8.0050 63.4770 ;
        RECT 7.8710 62.3835 7.8970 63.4770 ;
        RECT 7.7630 62.3835 7.7890 63.4770 ;
        RECT 7.6550 62.3835 7.6810 63.4770 ;
        RECT 7.5470 62.3835 7.5730 63.4770 ;
        RECT 7.4390 62.3835 7.4650 63.4770 ;
        RECT 7.3310 62.3835 7.3570 63.4770 ;
        RECT 7.2230 62.3835 7.2490 63.4770 ;
        RECT 7.1150 62.3835 7.1410 63.4770 ;
        RECT 7.0070 62.3835 7.0330 63.4770 ;
        RECT 6.8990 62.3835 6.9250 63.4770 ;
        RECT 6.7910 62.3835 6.8170 63.4770 ;
        RECT 6.6830 62.3835 6.7090 63.4770 ;
        RECT 6.5750 62.3835 6.6010 63.4770 ;
        RECT 6.4670 62.3835 6.4930 63.4770 ;
        RECT 6.3590 62.3835 6.3850 63.4770 ;
        RECT 6.2510 62.3835 6.2770 63.4770 ;
        RECT 6.1430 62.3835 6.1690 63.4770 ;
        RECT 6.0350 62.3835 6.0610 63.4770 ;
        RECT 5.9270 62.3835 5.9530 63.4770 ;
        RECT 5.7140 62.3835 5.7910 63.4770 ;
        RECT 3.8210 62.3835 3.8980 63.4770 ;
        RECT 3.6590 62.3835 3.6850 63.4770 ;
        RECT 3.5510 62.3835 3.5770 63.4770 ;
        RECT 3.4430 62.3835 3.4690 63.4770 ;
        RECT 3.3350 62.3835 3.3610 63.4770 ;
        RECT 3.2270 62.3835 3.2530 63.4770 ;
        RECT 3.1190 62.3835 3.1450 63.4770 ;
        RECT 3.0110 62.3835 3.0370 63.4770 ;
        RECT 2.9030 62.3835 2.9290 63.4770 ;
        RECT 2.7950 62.3835 2.8210 63.4770 ;
        RECT 2.6870 62.3835 2.7130 63.4770 ;
        RECT 2.5790 62.3835 2.6050 63.4770 ;
        RECT 2.4710 62.3835 2.4970 63.4770 ;
        RECT 2.3630 62.3835 2.3890 63.4770 ;
        RECT 2.2550 62.3835 2.2810 63.4770 ;
        RECT 2.1470 62.3835 2.1730 63.4770 ;
        RECT 2.0390 62.3835 2.0650 63.4770 ;
        RECT 1.9310 62.3835 1.9570 63.4770 ;
        RECT 1.8230 62.3835 1.8490 63.4770 ;
        RECT 1.7150 62.3835 1.7410 63.4770 ;
        RECT 1.6070 62.3835 1.6330 63.4770 ;
        RECT 1.4990 62.3835 1.5250 63.4770 ;
        RECT 1.3910 62.3835 1.4170 63.4770 ;
        RECT 1.2830 62.3835 1.3090 63.4770 ;
        RECT 1.1750 62.3835 1.2010 63.4770 ;
        RECT 1.0670 62.3835 1.0930 63.4770 ;
        RECT 0.9590 62.3835 0.9850 63.4770 ;
        RECT 0.8510 62.3835 0.8770 63.4770 ;
        RECT 0.7430 62.3835 0.7690 63.4770 ;
        RECT 0.6350 62.3835 0.6610 63.4770 ;
        RECT 0.5270 62.3835 0.5530 63.4770 ;
        RECT 0.4190 62.3835 0.4450 63.4770 ;
        RECT 0.3110 62.3835 0.3370 63.4770 ;
        RECT 0.2030 62.3835 0.2290 63.4770 ;
        RECT 0.0000 62.3835 0.0850 63.4770 ;
        RECT 5.1800 63.4635 5.3080 64.5570 ;
        RECT 5.1660 64.1290 5.3080 64.4515 ;
        RECT 5.0180 63.8560 5.0800 64.5570 ;
        RECT 5.0040 64.1655 5.0800 64.3190 ;
        RECT 5.0180 63.4635 5.0440 64.5570 ;
        RECT 5.0180 63.5845 5.0580 63.8240 ;
        RECT 5.0180 63.4635 5.0800 63.5525 ;
        RECT 4.7210 63.9140 4.9270 64.5570 ;
        RECT 4.9010 63.4635 4.9270 64.5570 ;
        RECT 4.7210 64.1910 4.9410 64.4490 ;
        RECT 4.7210 63.4635 4.8190 64.5570 ;
        RECT 4.3040 63.4635 4.3870 64.5570 ;
        RECT 4.3040 63.5520 4.4010 64.4875 ;
        RECT 9.5270 63.4635 9.6120 64.5570 ;
        RECT 9.3830 63.4635 9.4090 64.5570 ;
        RECT 9.2750 63.4635 9.3010 64.5570 ;
        RECT 9.1670 63.4635 9.1930 64.5570 ;
        RECT 9.0590 63.4635 9.0850 64.5570 ;
        RECT 8.9510 63.4635 8.9770 64.5570 ;
        RECT 8.8430 63.4635 8.8690 64.5570 ;
        RECT 8.7350 63.4635 8.7610 64.5570 ;
        RECT 8.6270 63.4635 8.6530 64.5570 ;
        RECT 8.5190 63.4635 8.5450 64.5570 ;
        RECT 8.4110 63.4635 8.4370 64.5570 ;
        RECT 8.3030 63.4635 8.3290 64.5570 ;
        RECT 8.1950 63.4635 8.2210 64.5570 ;
        RECT 8.0870 63.4635 8.1130 64.5570 ;
        RECT 7.9790 63.4635 8.0050 64.5570 ;
        RECT 7.8710 63.4635 7.8970 64.5570 ;
        RECT 7.7630 63.4635 7.7890 64.5570 ;
        RECT 7.6550 63.4635 7.6810 64.5570 ;
        RECT 7.5470 63.4635 7.5730 64.5570 ;
        RECT 7.4390 63.4635 7.4650 64.5570 ;
        RECT 7.3310 63.4635 7.3570 64.5570 ;
        RECT 7.2230 63.4635 7.2490 64.5570 ;
        RECT 7.1150 63.4635 7.1410 64.5570 ;
        RECT 7.0070 63.4635 7.0330 64.5570 ;
        RECT 6.8990 63.4635 6.9250 64.5570 ;
        RECT 6.7910 63.4635 6.8170 64.5570 ;
        RECT 6.6830 63.4635 6.7090 64.5570 ;
        RECT 6.5750 63.4635 6.6010 64.5570 ;
        RECT 6.4670 63.4635 6.4930 64.5570 ;
        RECT 6.3590 63.4635 6.3850 64.5570 ;
        RECT 6.2510 63.4635 6.2770 64.5570 ;
        RECT 6.1430 63.4635 6.1690 64.5570 ;
        RECT 6.0350 63.4635 6.0610 64.5570 ;
        RECT 5.9270 63.4635 5.9530 64.5570 ;
        RECT 5.7140 63.4635 5.7910 64.5570 ;
        RECT 3.8210 63.4635 3.8980 64.5570 ;
        RECT 3.6590 63.4635 3.6850 64.5570 ;
        RECT 3.5510 63.4635 3.5770 64.5570 ;
        RECT 3.4430 63.4635 3.4690 64.5570 ;
        RECT 3.3350 63.4635 3.3610 64.5570 ;
        RECT 3.2270 63.4635 3.2530 64.5570 ;
        RECT 3.1190 63.4635 3.1450 64.5570 ;
        RECT 3.0110 63.4635 3.0370 64.5570 ;
        RECT 2.9030 63.4635 2.9290 64.5570 ;
        RECT 2.7950 63.4635 2.8210 64.5570 ;
        RECT 2.6870 63.4635 2.7130 64.5570 ;
        RECT 2.5790 63.4635 2.6050 64.5570 ;
        RECT 2.4710 63.4635 2.4970 64.5570 ;
        RECT 2.3630 63.4635 2.3890 64.5570 ;
        RECT 2.2550 63.4635 2.2810 64.5570 ;
        RECT 2.1470 63.4635 2.1730 64.5570 ;
        RECT 2.0390 63.4635 2.0650 64.5570 ;
        RECT 1.9310 63.4635 1.9570 64.5570 ;
        RECT 1.8230 63.4635 1.8490 64.5570 ;
        RECT 1.7150 63.4635 1.7410 64.5570 ;
        RECT 1.6070 63.4635 1.6330 64.5570 ;
        RECT 1.4990 63.4635 1.5250 64.5570 ;
        RECT 1.3910 63.4635 1.4170 64.5570 ;
        RECT 1.2830 63.4635 1.3090 64.5570 ;
        RECT 1.1750 63.4635 1.2010 64.5570 ;
        RECT 1.0670 63.4635 1.0930 64.5570 ;
        RECT 0.9590 63.4635 0.9850 64.5570 ;
        RECT 0.8510 63.4635 0.8770 64.5570 ;
        RECT 0.7430 63.4635 0.7690 64.5570 ;
        RECT 0.6350 63.4635 0.6610 64.5570 ;
        RECT 0.5270 63.4635 0.5530 64.5570 ;
        RECT 0.4190 63.4635 0.4450 64.5570 ;
        RECT 0.3110 63.4635 0.3370 64.5570 ;
        RECT 0.2030 63.4635 0.2290 64.5570 ;
        RECT 0.0000 63.4635 0.0850 64.5570 ;
        RECT 5.1800 64.5435 5.3080 65.6370 ;
        RECT 5.1660 65.2090 5.3080 65.5315 ;
        RECT 5.0180 64.9360 5.0800 65.6370 ;
        RECT 5.0040 65.2455 5.0800 65.3990 ;
        RECT 5.0180 64.5435 5.0440 65.6370 ;
        RECT 5.0180 64.6645 5.0580 64.9040 ;
        RECT 5.0180 64.5435 5.0800 64.6325 ;
        RECT 4.7210 64.9940 4.9270 65.6370 ;
        RECT 4.9010 64.5435 4.9270 65.6370 ;
        RECT 4.7210 65.2710 4.9410 65.5290 ;
        RECT 4.7210 64.5435 4.8190 65.6370 ;
        RECT 4.3040 64.5435 4.3870 65.6370 ;
        RECT 4.3040 64.6320 4.4010 65.5675 ;
        RECT 9.5270 64.5435 9.6120 65.6370 ;
        RECT 9.3830 64.5435 9.4090 65.6370 ;
        RECT 9.2750 64.5435 9.3010 65.6370 ;
        RECT 9.1670 64.5435 9.1930 65.6370 ;
        RECT 9.0590 64.5435 9.0850 65.6370 ;
        RECT 8.9510 64.5435 8.9770 65.6370 ;
        RECT 8.8430 64.5435 8.8690 65.6370 ;
        RECT 8.7350 64.5435 8.7610 65.6370 ;
        RECT 8.6270 64.5435 8.6530 65.6370 ;
        RECT 8.5190 64.5435 8.5450 65.6370 ;
        RECT 8.4110 64.5435 8.4370 65.6370 ;
        RECT 8.3030 64.5435 8.3290 65.6370 ;
        RECT 8.1950 64.5435 8.2210 65.6370 ;
        RECT 8.0870 64.5435 8.1130 65.6370 ;
        RECT 7.9790 64.5435 8.0050 65.6370 ;
        RECT 7.8710 64.5435 7.8970 65.6370 ;
        RECT 7.7630 64.5435 7.7890 65.6370 ;
        RECT 7.6550 64.5435 7.6810 65.6370 ;
        RECT 7.5470 64.5435 7.5730 65.6370 ;
        RECT 7.4390 64.5435 7.4650 65.6370 ;
        RECT 7.3310 64.5435 7.3570 65.6370 ;
        RECT 7.2230 64.5435 7.2490 65.6370 ;
        RECT 7.1150 64.5435 7.1410 65.6370 ;
        RECT 7.0070 64.5435 7.0330 65.6370 ;
        RECT 6.8990 64.5435 6.9250 65.6370 ;
        RECT 6.7910 64.5435 6.8170 65.6370 ;
        RECT 6.6830 64.5435 6.7090 65.6370 ;
        RECT 6.5750 64.5435 6.6010 65.6370 ;
        RECT 6.4670 64.5435 6.4930 65.6370 ;
        RECT 6.3590 64.5435 6.3850 65.6370 ;
        RECT 6.2510 64.5435 6.2770 65.6370 ;
        RECT 6.1430 64.5435 6.1690 65.6370 ;
        RECT 6.0350 64.5435 6.0610 65.6370 ;
        RECT 5.9270 64.5435 5.9530 65.6370 ;
        RECT 5.7140 64.5435 5.7910 65.6370 ;
        RECT 3.8210 64.5435 3.8980 65.6370 ;
        RECT 3.6590 64.5435 3.6850 65.6370 ;
        RECT 3.5510 64.5435 3.5770 65.6370 ;
        RECT 3.4430 64.5435 3.4690 65.6370 ;
        RECT 3.3350 64.5435 3.3610 65.6370 ;
        RECT 3.2270 64.5435 3.2530 65.6370 ;
        RECT 3.1190 64.5435 3.1450 65.6370 ;
        RECT 3.0110 64.5435 3.0370 65.6370 ;
        RECT 2.9030 64.5435 2.9290 65.6370 ;
        RECT 2.7950 64.5435 2.8210 65.6370 ;
        RECT 2.6870 64.5435 2.7130 65.6370 ;
        RECT 2.5790 64.5435 2.6050 65.6370 ;
        RECT 2.4710 64.5435 2.4970 65.6370 ;
        RECT 2.3630 64.5435 2.3890 65.6370 ;
        RECT 2.2550 64.5435 2.2810 65.6370 ;
        RECT 2.1470 64.5435 2.1730 65.6370 ;
        RECT 2.0390 64.5435 2.0650 65.6370 ;
        RECT 1.9310 64.5435 1.9570 65.6370 ;
        RECT 1.8230 64.5435 1.8490 65.6370 ;
        RECT 1.7150 64.5435 1.7410 65.6370 ;
        RECT 1.6070 64.5435 1.6330 65.6370 ;
        RECT 1.4990 64.5435 1.5250 65.6370 ;
        RECT 1.3910 64.5435 1.4170 65.6370 ;
        RECT 1.2830 64.5435 1.3090 65.6370 ;
        RECT 1.1750 64.5435 1.2010 65.6370 ;
        RECT 1.0670 64.5435 1.0930 65.6370 ;
        RECT 0.9590 64.5435 0.9850 65.6370 ;
        RECT 0.8510 64.5435 0.8770 65.6370 ;
        RECT 0.7430 64.5435 0.7690 65.6370 ;
        RECT 0.6350 64.5435 0.6610 65.6370 ;
        RECT 0.5270 64.5435 0.5530 65.6370 ;
        RECT 0.4190 64.5435 0.4450 65.6370 ;
        RECT 0.3110 64.5435 0.3370 65.6370 ;
        RECT 0.2030 64.5435 0.2290 65.6370 ;
        RECT 0.0000 64.5435 0.0850 65.6370 ;
        RECT 5.1800 65.6235 5.3080 66.7170 ;
        RECT 5.1660 66.2890 5.3080 66.6115 ;
        RECT 5.0180 66.0160 5.0800 66.7170 ;
        RECT 5.0040 66.3255 5.0800 66.4790 ;
        RECT 5.0180 65.6235 5.0440 66.7170 ;
        RECT 5.0180 65.7445 5.0580 65.9840 ;
        RECT 5.0180 65.6235 5.0800 65.7125 ;
        RECT 4.7210 66.0740 4.9270 66.7170 ;
        RECT 4.9010 65.6235 4.9270 66.7170 ;
        RECT 4.7210 66.3510 4.9410 66.6090 ;
        RECT 4.7210 65.6235 4.8190 66.7170 ;
        RECT 4.3040 65.6235 4.3870 66.7170 ;
        RECT 4.3040 65.7120 4.4010 66.6475 ;
        RECT 9.5270 65.6235 9.6120 66.7170 ;
        RECT 9.3830 65.6235 9.4090 66.7170 ;
        RECT 9.2750 65.6235 9.3010 66.7170 ;
        RECT 9.1670 65.6235 9.1930 66.7170 ;
        RECT 9.0590 65.6235 9.0850 66.7170 ;
        RECT 8.9510 65.6235 8.9770 66.7170 ;
        RECT 8.8430 65.6235 8.8690 66.7170 ;
        RECT 8.7350 65.6235 8.7610 66.7170 ;
        RECT 8.6270 65.6235 8.6530 66.7170 ;
        RECT 8.5190 65.6235 8.5450 66.7170 ;
        RECT 8.4110 65.6235 8.4370 66.7170 ;
        RECT 8.3030 65.6235 8.3290 66.7170 ;
        RECT 8.1950 65.6235 8.2210 66.7170 ;
        RECT 8.0870 65.6235 8.1130 66.7170 ;
        RECT 7.9790 65.6235 8.0050 66.7170 ;
        RECT 7.8710 65.6235 7.8970 66.7170 ;
        RECT 7.7630 65.6235 7.7890 66.7170 ;
        RECT 7.6550 65.6235 7.6810 66.7170 ;
        RECT 7.5470 65.6235 7.5730 66.7170 ;
        RECT 7.4390 65.6235 7.4650 66.7170 ;
        RECT 7.3310 65.6235 7.3570 66.7170 ;
        RECT 7.2230 65.6235 7.2490 66.7170 ;
        RECT 7.1150 65.6235 7.1410 66.7170 ;
        RECT 7.0070 65.6235 7.0330 66.7170 ;
        RECT 6.8990 65.6235 6.9250 66.7170 ;
        RECT 6.7910 65.6235 6.8170 66.7170 ;
        RECT 6.6830 65.6235 6.7090 66.7170 ;
        RECT 6.5750 65.6235 6.6010 66.7170 ;
        RECT 6.4670 65.6235 6.4930 66.7170 ;
        RECT 6.3590 65.6235 6.3850 66.7170 ;
        RECT 6.2510 65.6235 6.2770 66.7170 ;
        RECT 6.1430 65.6235 6.1690 66.7170 ;
        RECT 6.0350 65.6235 6.0610 66.7170 ;
        RECT 5.9270 65.6235 5.9530 66.7170 ;
        RECT 5.7140 65.6235 5.7910 66.7170 ;
        RECT 3.8210 65.6235 3.8980 66.7170 ;
        RECT 3.6590 65.6235 3.6850 66.7170 ;
        RECT 3.5510 65.6235 3.5770 66.7170 ;
        RECT 3.4430 65.6235 3.4690 66.7170 ;
        RECT 3.3350 65.6235 3.3610 66.7170 ;
        RECT 3.2270 65.6235 3.2530 66.7170 ;
        RECT 3.1190 65.6235 3.1450 66.7170 ;
        RECT 3.0110 65.6235 3.0370 66.7170 ;
        RECT 2.9030 65.6235 2.9290 66.7170 ;
        RECT 2.7950 65.6235 2.8210 66.7170 ;
        RECT 2.6870 65.6235 2.7130 66.7170 ;
        RECT 2.5790 65.6235 2.6050 66.7170 ;
        RECT 2.4710 65.6235 2.4970 66.7170 ;
        RECT 2.3630 65.6235 2.3890 66.7170 ;
        RECT 2.2550 65.6235 2.2810 66.7170 ;
        RECT 2.1470 65.6235 2.1730 66.7170 ;
        RECT 2.0390 65.6235 2.0650 66.7170 ;
        RECT 1.9310 65.6235 1.9570 66.7170 ;
        RECT 1.8230 65.6235 1.8490 66.7170 ;
        RECT 1.7150 65.6235 1.7410 66.7170 ;
        RECT 1.6070 65.6235 1.6330 66.7170 ;
        RECT 1.4990 65.6235 1.5250 66.7170 ;
        RECT 1.3910 65.6235 1.4170 66.7170 ;
        RECT 1.2830 65.6235 1.3090 66.7170 ;
        RECT 1.1750 65.6235 1.2010 66.7170 ;
        RECT 1.0670 65.6235 1.0930 66.7170 ;
        RECT 0.9590 65.6235 0.9850 66.7170 ;
        RECT 0.8510 65.6235 0.8770 66.7170 ;
        RECT 0.7430 65.6235 0.7690 66.7170 ;
        RECT 0.6350 65.6235 0.6610 66.7170 ;
        RECT 0.5270 65.6235 0.5530 66.7170 ;
        RECT 0.4190 65.6235 0.4450 66.7170 ;
        RECT 0.3110 65.6235 0.3370 66.7170 ;
        RECT 0.2030 65.6235 0.2290 66.7170 ;
        RECT 0.0000 65.6235 0.0850 66.7170 ;
        RECT 5.1800 66.7035 5.3080 67.7970 ;
        RECT 5.1660 67.3690 5.3080 67.6915 ;
        RECT 5.0180 67.0960 5.0800 67.7970 ;
        RECT 5.0040 67.4055 5.0800 67.5590 ;
        RECT 5.0180 66.7035 5.0440 67.7970 ;
        RECT 5.0180 66.8245 5.0580 67.0640 ;
        RECT 5.0180 66.7035 5.0800 66.7925 ;
        RECT 4.7210 67.1540 4.9270 67.7970 ;
        RECT 4.9010 66.7035 4.9270 67.7970 ;
        RECT 4.7210 67.4310 4.9410 67.6890 ;
        RECT 4.7210 66.7035 4.8190 67.7970 ;
        RECT 4.3040 66.7035 4.3870 67.7970 ;
        RECT 4.3040 66.7920 4.4010 67.7275 ;
        RECT 9.5270 66.7035 9.6120 67.7970 ;
        RECT 9.3830 66.7035 9.4090 67.7970 ;
        RECT 9.2750 66.7035 9.3010 67.7970 ;
        RECT 9.1670 66.7035 9.1930 67.7970 ;
        RECT 9.0590 66.7035 9.0850 67.7970 ;
        RECT 8.9510 66.7035 8.9770 67.7970 ;
        RECT 8.8430 66.7035 8.8690 67.7970 ;
        RECT 8.7350 66.7035 8.7610 67.7970 ;
        RECT 8.6270 66.7035 8.6530 67.7970 ;
        RECT 8.5190 66.7035 8.5450 67.7970 ;
        RECT 8.4110 66.7035 8.4370 67.7970 ;
        RECT 8.3030 66.7035 8.3290 67.7970 ;
        RECT 8.1950 66.7035 8.2210 67.7970 ;
        RECT 8.0870 66.7035 8.1130 67.7970 ;
        RECT 7.9790 66.7035 8.0050 67.7970 ;
        RECT 7.8710 66.7035 7.8970 67.7970 ;
        RECT 7.7630 66.7035 7.7890 67.7970 ;
        RECT 7.6550 66.7035 7.6810 67.7970 ;
        RECT 7.5470 66.7035 7.5730 67.7970 ;
        RECT 7.4390 66.7035 7.4650 67.7970 ;
        RECT 7.3310 66.7035 7.3570 67.7970 ;
        RECT 7.2230 66.7035 7.2490 67.7970 ;
        RECT 7.1150 66.7035 7.1410 67.7970 ;
        RECT 7.0070 66.7035 7.0330 67.7970 ;
        RECT 6.8990 66.7035 6.9250 67.7970 ;
        RECT 6.7910 66.7035 6.8170 67.7970 ;
        RECT 6.6830 66.7035 6.7090 67.7970 ;
        RECT 6.5750 66.7035 6.6010 67.7970 ;
        RECT 6.4670 66.7035 6.4930 67.7970 ;
        RECT 6.3590 66.7035 6.3850 67.7970 ;
        RECT 6.2510 66.7035 6.2770 67.7970 ;
        RECT 6.1430 66.7035 6.1690 67.7970 ;
        RECT 6.0350 66.7035 6.0610 67.7970 ;
        RECT 5.9270 66.7035 5.9530 67.7970 ;
        RECT 5.7140 66.7035 5.7910 67.7970 ;
        RECT 3.8210 66.7035 3.8980 67.7970 ;
        RECT 3.6590 66.7035 3.6850 67.7970 ;
        RECT 3.5510 66.7035 3.5770 67.7970 ;
        RECT 3.4430 66.7035 3.4690 67.7970 ;
        RECT 3.3350 66.7035 3.3610 67.7970 ;
        RECT 3.2270 66.7035 3.2530 67.7970 ;
        RECT 3.1190 66.7035 3.1450 67.7970 ;
        RECT 3.0110 66.7035 3.0370 67.7970 ;
        RECT 2.9030 66.7035 2.9290 67.7970 ;
        RECT 2.7950 66.7035 2.8210 67.7970 ;
        RECT 2.6870 66.7035 2.7130 67.7970 ;
        RECT 2.5790 66.7035 2.6050 67.7970 ;
        RECT 2.4710 66.7035 2.4970 67.7970 ;
        RECT 2.3630 66.7035 2.3890 67.7970 ;
        RECT 2.2550 66.7035 2.2810 67.7970 ;
        RECT 2.1470 66.7035 2.1730 67.7970 ;
        RECT 2.0390 66.7035 2.0650 67.7970 ;
        RECT 1.9310 66.7035 1.9570 67.7970 ;
        RECT 1.8230 66.7035 1.8490 67.7970 ;
        RECT 1.7150 66.7035 1.7410 67.7970 ;
        RECT 1.6070 66.7035 1.6330 67.7970 ;
        RECT 1.4990 66.7035 1.5250 67.7970 ;
        RECT 1.3910 66.7035 1.4170 67.7970 ;
        RECT 1.2830 66.7035 1.3090 67.7970 ;
        RECT 1.1750 66.7035 1.2010 67.7970 ;
        RECT 1.0670 66.7035 1.0930 67.7970 ;
        RECT 0.9590 66.7035 0.9850 67.7970 ;
        RECT 0.8510 66.7035 0.8770 67.7970 ;
        RECT 0.7430 66.7035 0.7690 67.7970 ;
        RECT 0.6350 66.7035 0.6610 67.7970 ;
        RECT 0.5270 66.7035 0.5530 67.7970 ;
        RECT 0.4190 66.7035 0.4450 67.7970 ;
        RECT 0.3110 66.7035 0.3370 67.7970 ;
        RECT 0.2030 66.7035 0.2290 67.7970 ;
        RECT 0.0000 66.7035 0.0850 67.7970 ;
        RECT 5.1800 67.7835 5.3080 68.8770 ;
        RECT 5.1660 68.4490 5.3080 68.7715 ;
        RECT 5.0180 68.1760 5.0800 68.8770 ;
        RECT 5.0040 68.4855 5.0800 68.6390 ;
        RECT 5.0180 67.7835 5.0440 68.8770 ;
        RECT 5.0180 67.9045 5.0580 68.1440 ;
        RECT 5.0180 67.7835 5.0800 67.8725 ;
        RECT 4.7210 68.2340 4.9270 68.8770 ;
        RECT 4.9010 67.7835 4.9270 68.8770 ;
        RECT 4.7210 68.5110 4.9410 68.7690 ;
        RECT 4.7210 67.7835 4.8190 68.8770 ;
        RECT 4.3040 67.7835 4.3870 68.8770 ;
        RECT 4.3040 67.8720 4.4010 68.8075 ;
        RECT 9.5270 67.7835 9.6120 68.8770 ;
        RECT 9.3830 67.7835 9.4090 68.8770 ;
        RECT 9.2750 67.7835 9.3010 68.8770 ;
        RECT 9.1670 67.7835 9.1930 68.8770 ;
        RECT 9.0590 67.7835 9.0850 68.8770 ;
        RECT 8.9510 67.7835 8.9770 68.8770 ;
        RECT 8.8430 67.7835 8.8690 68.8770 ;
        RECT 8.7350 67.7835 8.7610 68.8770 ;
        RECT 8.6270 67.7835 8.6530 68.8770 ;
        RECT 8.5190 67.7835 8.5450 68.8770 ;
        RECT 8.4110 67.7835 8.4370 68.8770 ;
        RECT 8.3030 67.7835 8.3290 68.8770 ;
        RECT 8.1950 67.7835 8.2210 68.8770 ;
        RECT 8.0870 67.7835 8.1130 68.8770 ;
        RECT 7.9790 67.7835 8.0050 68.8770 ;
        RECT 7.8710 67.7835 7.8970 68.8770 ;
        RECT 7.7630 67.7835 7.7890 68.8770 ;
        RECT 7.6550 67.7835 7.6810 68.8770 ;
        RECT 7.5470 67.7835 7.5730 68.8770 ;
        RECT 7.4390 67.7835 7.4650 68.8770 ;
        RECT 7.3310 67.7835 7.3570 68.8770 ;
        RECT 7.2230 67.7835 7.2490 68.8770 ;
        RECT 7.1150 67.7835 7.1410 68.8770 ;
        RECT 7.0070 67.7835 7.0330 68.8770 ;
        RECT 6.8990 67.7835 6.9250 68.8770 ;
        RECT 6.7910 67.7835 6.8170 68.8770 ;
        RECT 6.6830 67.7835 6.7090 68.8770 ;
        RECT 6.5750 67.7835 6.6010 68.8770 ;
        RECT 6.4670 67.7835 6.4930 68.8770 ;
        RECT 6.3590 67.7835 6.3850 68.8770 ;
        RECT 6.2510 67.7835 6.2770 68.8770 ;
        RECT 6.1430 67.7835 6.1690 68.8770 ;
        RECT 6.0350 67.7835 6.0610 68.8770 ;
        RECT 5.9270 67.7835 5.9530 68.8770 ;
        RECT 5.7140 67.7835 5.7910 68.8770 ;
        RECT 3.8210 67.7835 3.8980 68.8770 ;
        RECT 3.6590 67.7835 3.6850 68.8770 ;
        RECT 3.5510 67.7835 3.5770 68.8770 ;
        RECT 3.4430 67.7835 3.4690 68.8770 ;
        RECT 3.3350 67.7835 3.3610 68.8770 ;
        RECT 3.2270 67.7835 3.2530 68.8770 ;
        RECT 3.1190 67.7835 3.1450 68.8770 ;
        RECT 3.0110 67.7835 3.0370 68.8770 ;
        RECT 2.9030 67.7835 2.9290 68.8770 ;
        RECT 2.7950 67.7835 2.8210 68.8770 ;
        RECT 2.6870 67.7835 2.7130 68.8770 ;
        RECT 2.5790 67.7835 2.6050 68.8770 ;
        RECT 2.4710 67.7835 2.4970 68.8770 ;
        RECT 2.3630 67.7835 2.3890 68.8770 ;
        RECT 2.2550 67.7835 2.2810 68.8770 ;
        RECT 2.1470 67.7835 2.1730 68.8770 ;
        RECT 2.0390 67.7835 2.0650 68.8770 ;
        RECT 1.9310 67.7835 1.9570 68.8770 ;
        RECT 1.8230 67.7835 1.8490 68.8770 ;
        RECT 1.7150 67.7835 1.7410 68.8770 ;
        RECT 1.6070 67.7835 1.6330 68.8770 ;
        RECT 1.4990 67.7835 1.5250 68.8770 ;
        RECT 1.3910 67.7835 1.4170 68.8770 ;
        RECT 1.2830 67.7835 1.3090 68.8770 ;
        RECT 1.1750 67.7835 1.2010 68.8770 ;
        RECT 1.0670 67.7835 1.0930 68.8770 ;
        RECT 0.9590 67.7835 0.9850 68.8770 ;
        RECT 0.8510 67.7835 0.8770 68.8770 ;
        RECT 0.7430 67.7835 0.7690 68.8770 ;
        RECT 0.6350 67.7835 0.6610 68.8770 ;
        RECT 0.5270 67.7835 0.5530 68.8770 ;
        RECT 0.4190 67.7835 0.4450 68.8770 ;
        RECT 0.3110 67.7835 0.3370 68.8770 ;
        RECT 0.2030 67.7835 0.2290 68.8770 ;
        RECT 0.0000 67.7835 0.0850 68.8770 ;
        RECT 5.1800 68.8635 5.3080 69.9570 ;
        RECT 5.1660 69.5290 5.3080 69.8515 ;
        RECT 5.0180 69.2560 5.0800 69.9570 ;
        RECT 5.0040 69.5655 5.0800 69.7190 ;
        RECT 5.0180 68.8635 5.0440 69.9570 ;
        RECT 5.0180 68.9845 5.0580 69.2240 ;
        RECT 5.0180 68.8635 5.0800 68.9525 ;
        RECT 4.7210 69.3140 4.9270 69.9570 ;
        RECT 4.9010 68.8635 4.9270 69.9570 ;
        RECT 4.7210 69.5910 4.9410 69.8490 ;
        RECT 4.7210 68.8635 4.8190 69.9570 ;
        RECT 4.3040 68.8635 4.3870 69.9570 ;
        RECT 4.3040 68.9520 4.4010 69.8875 ;
        RECT 9.5270 68.8635 9.6120 69.9570 ;
        RECT 9.3830 68.8635 9.4090 69.9570 ;
        RECT 9.2750 68.8635 9.3010 69.9570 ;
        RECT 9.1670 68.8635 9.1930 69.9570 ;
        RECT 9.0590 68.8635 9.0850 69.9570 ;
        RECT 8.9510 68.8635 8.9770 69.9570 ;
        RECT 8.8430 68.8635 8.8690 69.9570 ;
        RECT 8.7350 68.8635 8.7610 69.9570 ;
        RECT 8.6270 68.8635 8.6530 69.9570 ;
        RECT 8.5190 68.8635 8.5450 69.9570 ;
        RECT 8.4110 68.8635 8.4370 69.9570 ;
        RECT 8.3030 68.8635 8.3290 69.9570 ;
        RECT 8.1950 68.8635 8.2210 69.9570 ;
        RECT 8.0870 68.8635 8.1130 69.9570 ;
        RECT 7.9790 68.8635 8.0050 69.9570 ;
        RECT 7.8710 68.8635 7.8970 69.9570 ;
        RECT 7.7630 68.8635 7.7890 69.9570 ;
        RECT 7.6550 68.8635 7.6810 69.9570 ;
        RECT 7.5470 68.8635 7.5730 69.9570 ;
        RECT 7.4390 68.8635 7.4650 69.9570 ;
        RECT 7.3310 68.8635 7.3570 69.9570 ;
        RECT 7.2230 68.8635 7.2490 69.9570 ;
        RECT 7.1150 68.8635 7.1410 69.9570 ;
        RECT 7.0070 68.8635 7.0330 69.9570 ;
        RECT 6.8990 68.8635 6.9250 69.9570 ;
        RECT 6.7910 68.8635 6.8170 69.9570 ;
        RECT 6.6830 68.8635 6.7090 69.9570 ;
        RECT 6.5750 68.8635 6.6010 69.9570 ;
        RECT 6.4670 68.8635 6.4930 69.9570 ;
        RECT 6.3590 68.8635 6.3850 69.9570 ;
        RECT 6.2510 68.8635 6.2770 69.9570 ;
        RECT 6.1430 68.8635 6.1690 69.9570 ;
        RECT 6.0350 68.8635 6.0610 69.9570 ;
        RECT 5.9270 68.8635 5.9530 69.9570 ;
        RECT 5.7140 68.8635 5.7910 69.9570 ;
        RECT 3.8210 68.8635 3.8980 69.9570 ;
        RECT 3.6590 68.8635 3.6850 69.9570 ;
        RECT 3.5510 68.8635 3.5770 69.9570 ;
        RECT 3.4430 68.8635 3.4690 69.9570 ;
        RECT 3.3350 68.8635 3.3610 69.9570 ;
        RECT 3.2270 68.8635 3.2530 69.9570 ;
        RECT 3.1190 68.8635 3.1450 69.9570 ;
        RECT 3.0110 68.8635 3.0370 69.9570 ;
        RECT 2.9030 68.8635 2.9290 69.9570 ;
        RECT 2.7950 68.8635 2.8210 69.9570 ;
        RECT 2.6870 68.8635 2.7130 69.9570 ;
        RECT 2.5790 68.8635 2.6050 69.9570 ;
        RECT 2.4710 68.8635 2.4970 69.9570 ;
        RECT 2.3630 68.8635 2.3890 69.9570 ;
        RECT 2.2550 68.8635 2.2810 69.9570 ;
        RECT 2.1470 68.8635 2.1730 69.9570 ;
        RECT 2.0390 68.8635 2.0650 69.9570 ;
        RECT 1.9310 68.8635 1.9570 69.9570 ;
        RECT 1.8230 68.8635 1.8490 69.9570 ;
        RECT 1.7150 68.8635 1.7410 69.9570 ;
        RECT 1.6070 68.8635 1.6330 69.9570 ;
        RECT 1.4990 68.8635 1.5250 69.9570 ;
        RECT 1.3910 68.8635 1.4170 69.9570 ;
        RECT 1.2830 68.8635 1.3090 69.9570 ;
        RECT 1.1750 68.8635 1.2010 69.9570 ;
        RECT 1.0670 68.8635 1.0930 69.9570 ;
        RECT 0.9590 68.8635 0.9850 69.9570 ;
        RECT 0.8510 68.8635 0.8770 69.9570 ;
        RECT 0.7430 68.8635 0.7690 69.9570 ;
        RECT 0.6350 68.8635 0.6610 69.9570 ;
        RECT 0.5270 68.8635 0.5530 69.9570 ;
        RECT 0.4190 68.8635 0.4450 69.9570 ;
        RECT 0.3110 68.8635 0.3370 69.9570 ;
        RECT 0.2030 68.8635 0.2290 69.9570 ;
        RECT 0.0000 68.8635 0.0850 69.9570 ;
        RECT 5.1800 69.9435 5.3080 71.0370 ;
        RECT 5.1660 70.6090 5.3080 70.9315 ;
        RECT 5.0180 70.3360 5.0800 71.0370 ;
        RECT 5.0040 70.6455 5.0800 70.7990 ;
        RECT 5.0180 69.9435 5.0440 71.0370 ;
        RECT 5.0180 70.0645 5.0580 70.3040 ;
        RECT 5.0180 69.9435 5.0800 70.0325 ;
        RECT 4.7210 70.3940 4.9270 71.0370 ;
        RECT 4.9010 69.9435 4.9270 71.0370 ;
        RECT 4.7210 70.6710 4.9410 70.9290 ;
        RECT 4.7210 69.9435 4.8190 71.0370 ;
        RECT 4.3040 69.9435 4.3870 71.0370 ;
        RECT 4.3040 70.0320 4.4010 70.9675 ;
        RECT 9.5270 69.9435 9.6120 71.0370 ;
        RECT 9.3830 69.9435 9.4090 71.0370 ;
        RECT 9.2750 69.9435 9.3010 71.0370 ;
        RECT 9.1670 69.9435 9.1930 71.0370 ;
        RECT 9.0590 69.9435 9.0850 71.0370 ;
        RECT 8.9510 69.9435 8.9770 71.0370 ;
        RECT 8.8430 69.9435 8.8690 71.0370 ;
        RECT 8.7350 69.9435 8.7610 71.0370 ;
        RECT 8.6270 69.9435 8.6530 71.0370 ;
        RECT 8.5190 69.9435 8.5450 71.0370 ;
        RECT 8.4110 69.9435 8.4370 71.0370 ;
        RECT 8.3030 69.9435 8.3290 71.0370 ;
        RECT 8.1950 69.9435 8.2210 71.0370 ;
        RECT 8.0870 69.9435 8.1130 71.0370 ;
        RECT 7.9790 69.9435 8.0050 71.0370 ;
        RECT 7.8710 69.9435 7.8970 71.0370 ;
        RECT 7.7630 69.9435 7.7890 71.0370 ;
        RECT 7.6550 69.9435 7.6810 71.0370 ;
        RECT 7.5470 69.9435 7.5730 71.0370 ;
        RECT 7.4390 69.9435 7.4650 71.0370 ;
        RECT 7.3310 69.9435 7.3570 71.0370 ;
        RECT 7.2230 69.9435 7.2490 71.0370 ;
        RECT 7.1150 69.9435 7.1410 71.0370 ;
        RECT 7.0070 69.9435 7.0330 71.0370 ;
        RECT 6.8990 69.9435 6.9250 71.0370 ;
        RECT 6.7910 69.9435 6.8170 71.0370 ;
        RECT 6.6830 69.9435 6.7090 71.0370 ;
        RECT 6.5750 69.9435 6.6010 71.0370 ;
        RECT 6.4670 69.9435 6.4930 71.0370 ;
        RECT 6.3590 69.9435 6.3850 71.0370 ;
        RECT 6.2510 69.9435 6.2770 71.0370 ;
        RECT 6.1430 69.9435 6.1690 71.0370 ;
        RECT 6.0350 69.9435 6.0610 71.0370 ;
        RECT 5.9270 69.9435 5.9530 71.0370 ;
        RECT 5.7140 69.9435 5.7910 71.0370 ;
        RECT 3.8210 69.9435 3.8980 71.0370 ;
        RECT 3.6590 69.9435 3.6850 71.0370 ;
        RECT 3.5510 69.9435 3.5770 71.0370 ;
        RECT 3.4430 69.9435 3.4690 71.0370 ;
        RECT 3.3350 69.9435 3.3610 71.0370 ;
        RECT 3.2270 69.9435 3.2530 71.0370 ;
        RECT 3.1190 69.9435 3.1450 71.0370 ;
        RECT 3.0110 69.9435 3.0370 71.0370 ;
        RECT 2.9030 69.9435 2.9290 71.0370 ;
        RECT 2.7950 69.9435 2.8210 71.0370 ;
        RECT 2.6870 69.9435 2.7130 71.0370 ;
        RECT 2.5790 69.9435 2.6050 71.0370 ;
        RECT 2.4710 69.9435 2.4970 71.0370 ;
        RECT 2.3630 69.9435 2.3890 71.0370 ;
        RECT 2.2550 69.9435 2.2810 71.0370 ;
        RECT 2.1470 69.9435 2.1730 71.0370 ;
        RECT 2.0390 69.9435 2.0650 71.0370 ;
        RECT 1.9310 69.9435 1.9570 71.0370 ;
        RECT 1.8230 69.9435 1.8490 71.0370 ;
        RECT 1.7150 69.9435 1.7410 71.0370 ;
        RECT 1.6070 69.9435 1.6330 71.0370 ;
        RECT 1.4990 69.9435 1.5250 71.0370 ;
        RECT 1.3910 69.9435 1.4170 71.0370 ;
        RECT 1.2830 69.9435 1.3090 71.0370 ;
        RECT 1.1750 69.9435 1.2010 71.0370 ;
        RECT 1.0670 69.9435 1.0930 71.0370 ;
        RECT 0.9590 69.9435 0.9850 71.0370 ;
        RECT 0.8510 69.9435 0.8770 71.0370 ;
        RECT 0.7430 69.9435 0.7690 71.0370 ;
        RECT 0.6350 69.9435 0.6610 71.0370 ;
        RECT 0.5270 69.9435 0.5530 71.0370 ;
        RECT 0.4190 69.9435 0.4450 71.0370 ;
        RECT 0.3110 69.9435 0.3370 71.0370 ;
        RECT 0.2030 69.9435 0.2290 71.0370 ;
        RECT 0.0000 69.9435 0.0850 71.0370 ;
        RECT 5.1800 71.0235 5.3080 72.1170 ;
        RECT 5.1660 71.6890 5.3080 72.0115 ;
        RECT 5.0180 71.4160 5.0800 72.1170 ;
        RECT 5.0040 71.7255 5.0800 71.8790 ;
        RECT 5.0180 71.0235 5.0440 72.1170 ;
        RECT 5.0180 71.1445 5.0580 71.3840 ;
        RECT 5.0180 71.0235 5.0800 71.1125 ;
        RECT 4.7210 71.4740 4.9270 72.1170 ;
        RECT 4.9010 71.0235 4.9270 72.1170 ;
        RECT 4.7210 71.7510 4.9410 72.0090 ;
        RECT 4.7210 71.0235 4.8190 72.1170 ;
        RECT 4.3040 71.0235 4.3870 72.1170 ;
        RECT 4.3040 71.1120 4.4010 72.0475 ;
        RECT 9.5270 71.0235 9.6120 72.1170 ;
        RECT 9.3830 71.0235 9.4090 72.1170 ;
        RECT 9.2750 71.0235 9.3010 72.1170 ;
        RECT 9.1670 71.0235 9.1930 72.1170 ;
        RECT 9.0590 71.0235 9.0850 72.1170 ;
        RECT 8.9510 71.0235 8.9770 72.1170 ;
        RECT 8.8430 71.0235 8.8690 72.1170 ;
        RECT 8.7350 71.0235 8.7610 72.1170 ;
        RECT 8.6270 71.0235 8.6530 72.1170 ;
        RECT 8.5190 71.0235 8.5450 72.1170 ;
        RECT 8.4110 71.0235 8.4370 72.1170 ;
        RECT 8.3030 71.0235 8.3290 72.1170 ;
        RECT 8.1950 71.0235 8.2210 72.1170 ;
        RECT 8.0870 71.0235 8.1130 72.1170 ;
        RECT 7.9790 71.0235 8.0050 72.1170 ;
        RECT 7.8710 71.0235 7.8970 72.1170 ;
        RECT 7.7630 71.0235 7.7890 72.1170 ;
        RECT 7.6550 71.0235 7.6810 72.1170 ;
        RECT 7.5470 71.0235 7.5730 72.1170 ;
        RECT 7.4390 71.0235 7.4650 72.1170 ;
        RECT 7.3310 71.0235 7.3570 72.1170 ;
        RECT 7.2230 71.0235 7.2490 72.1170 ;
        RECT 7.1150 71.0235 7.1410 72.1170 ;
        RECT 7.0070 71.0235 7.0330 72.1170 ;
        RECT 6.8990 71.0235 6.9250 72.1170 ;
        RECT 6.7910 71.0235 6.8170 72.1170 ;
        RECT 6.6830 71.0235 6.7090 72.1170 ;
        RECT 6.5750 71.0235 6.6010 72.1170 ;
        RECT 6.4670 71.0235 6.4930 72.1170 ;
        RECT 6.3590 71.0235 6.3850 72.1170 ;
        RECT 6.2510 71.0235 6.2770 72.1170 ;
        RECT 6.1430 71.0235 6.1690 72.1170 ;
        RECT 6.0350 71.0235 6.0610 72.1170 ;
        RECT 5.9270 71.0235 5.9530 72.1170 ;
        RECT 5.7140 71.0235 5.7910 72.1170 ;
        RECT 3.8210 71.0235 3.8980 72.1170 ;
        RECT 3.6590 71.0235 3.6850 72.1170 ;
        RECT 3.5510 71.0235 3.5770 72.1170 ;
        RECT 3.4430 71.0235 3.4690 72.1170 ;
        RECT 3.3350 71.0235 3.3610 72.1170 ;
        RECT 3.2270 71.0235 3.2530 72.1170 ;
        RECT 3.1190 71.0235 3.1450 72.1170 ;
        RECT 3.0110 71.0235 3.0370 72.1170 ;
        RECT 2.9030 71.0235 2.9290 72.1170 ;
        RECT 2.7950 71.0235 2.8210 72.1170 ;
        RECT 2.6870 71.0235 2.7130 72.1170 ;
        RECT 2.5790 71.0235 2.6050 72.1170 ;
        RECT 2.4710 71.0235 2.4970 72.1170 ;
        RECT 2.3630 71.0235 2.3890 72.1170 ;
        RECT 2.2550 71.0235 2.2810 72.1170 ;
        RECT 2.1470 71.0235 2.1730 72.1170 ;
        RECT 2.0390 71.0235 2.0650 72.1170 ;
        RECT 1.9310 71.0235 1.9570 72.1170 ;
        RECT 1.8230 71.0235 1.8490 72.1170 ;
        RECT 1.7150 71.0235 1.7410 72.1170 ;
        RECT 1.6070 71.0235 1.6330 72.1170 ;
        RECT 1.4990 71.0235 1.5250 72.1170 ;
        RECT 1.3910 71.0235 1.4170 72.1170 ;
        RECT 1.2830 71.0235 1.3090 72.1170 ;
        RECT 1.1750 71.0235 1.2010 72.1170 ;
        RECT 1.0670 71.0235 1.0930 72.1170 ;
        RECT 0.9590 71.0235 0.9850 72.1170 ;
        RECT 0.8510 71.0235 0.8770 72.1170 ;
        RECT 0.7430 71.0235 0.7690 72.1170 ;
        RECT 0.6350 71.0235 0.6610 72.1170 ;
        RECT 0.5270 71.0235 0.5530 72.1170 ;
        RECT 0.4190 71.0235 0.4450 72.1170 ;
        RECT 0.3110 71.0235 0.3370 72.1170 ;
        RECT 0.2030 71.0235 0.2290 72.1170 ;
        RECT 0.0000 71.0235 0.0850 72.1170 ;
        RECT 5.1800 72.1035 5.3080 73.1970 ;
        RECT 5.1660 72.7690 5.3080 73.0915 ;
        RECT 5.0180 72.4960 5.0800 73.1970 ;
        RECT 5.0040 72.8055 5.0800 72.9590 ;
        RECT 5.0180 72.1035 5.0440 73.1970 ;
        RECT 5.0180 72.2245 5.0580 72.4640 ;
        RECT 5.0180 72.1035 5.0800 72.1925 ;
        RECT 4.7210 72.5540 4.9270 73.1970 ;
        RECT 4.9010 72.1035 4.9270 73.1970 ;
        RECT 4.7210 72.8310 4.9410 73.0890 ;
        RECT 4.7210 72.1035 4.8190 73.1970 ;
        RECT 4.3040 72.1035 4.3870 73.1970 ;
        RECT 4.3040 72.1920 4.4010 73.1275 ;
        RECT 9.5270 72.1035 9.6120 73.1970 ;
        RECT 9.3830 72.1035 9.4090 73.1970 ;
        RECT 9.2750 72.1035 9.3010 73.1970 ;
        RECT 9.1670 72.1035 9.1930 73.1970 ;
        RECT 9.0590 72.1035 9.0850 73.1970 ;
        RECT 8.9510 72.1035 8.9770 73.1970 ;
        RECT 8.8430 72.1035 8.8690 73.1970 ;
        RECT 8.7350 72.1035 8.7610 73.1970 ;
        RECT 8.6270 72.1035 8.6530 73.1970 ;
        RECT 8.5190 72.1035 8.5450 73.1970 ;
        RECT 8.4110 72.1035 8.4370 73.1970 ;
        RECT 8.3030 72.1035 8.3290 73.1970 ;
        RECT 8.1950 72.1035 8.2210 73.1970 ;
        RECT 8.0870 72.1035 8.1130 73.1970 ;
        RECT 7.9790 72.1035 8.0050 73.1970 ;
        RECT 7.8710 72.1035 7.8970 73.1970 ;
        RECT 7.7630 72.1035 7.7890 73.1970 ;
        RECT 7.6550 72.1035 7.6810 73.1970 ;
        RECT 7.5470 72.1035 7.5730 73.1970 ;
        RECT 7.4390 72.1035 7.4650 73.1970 ;
        RECT 7.3310 72.1035 7.3570 73.1970 ;
        RECT 7.2230 72.1035 7.2490 73.1970 ;
        RECT 7.1150 72.1035 7.1410 73.1970 ;
        RECT 7.0070 72.1035 7.0330 73.1970 ;
        RECT 6.8990 72.1035 6.9250 73.1970 ;
        RECT 6.7910 72.1035 6.8170 73.1970 ;
        RECT 6.6830 72.1035 6.7090 73.1970 ;
        RECT 6.5750 72.1035 6.6010 73.1970 ;
        RECT 6.4670 72.1035 6.4930 73.1970 ;
        RECT 6.3590 72.1035 6.3850 73.1970 ;
        RECT 6.2510 72.1035 6.2770 73.1970 ;
        RECT 6.1430 72.1035 6.1690 73.1970 ;
        RECT 6.0350 72.1035 6.0610 73.1970 ;
        RECT 5.9270 72.1035 5.9530 73.1970 ;
        RECT 5.7140 72.1035 5.7910 73.1970 ;
        RECT 3.8210 72.1035 3.8980 73.1970 ;
        RECT 3.6590 72.1035 3.6850 73.1970 ;
        RECT 3.5510 72.1035 3.5770 73.1970 ;
        RECT 3.4430 72.1035 3.4690 73.1970 ;
        RECT 3.3350 72.1035 3.3610 73.1970 ;
        RECT 3.2270 72.1035 3.2530 73.1970 ;
        RECT 3.1190 72.1035 3.1450 73.1970 ;
        RECT 3.0110 72.1035 3.0370 73.1970 ;
        RECT 2.9030 72.1035 2.9290 73.1970 ;
        RECT 2.7950 72.1035 2.8210 73.1970 ;
        RECT 2.6870 72.1035 2.7130 73.1970 ;
        RECT 2.5790 72.1035 2.6050 73.1970 ;
        RECT 2.4710 72.1035 2.4970 73.1970 ;
        RECT 2.3630 72.1035 2.3890 73.1970 ;
        RECT 2.2550 72.1035 2.2810 73.1970 ;
        RECT 2.1470 72.1035 2.1730 73.1970 ;
        RECT 2.0390 72.1035 2.0650 73.1970 ;
        RECT 1.9310 72.1035 1.9570 73.1970 ;
        RECT 1.8230 72.1035 1.8490 73.1970 ;
        RECT 1.7150 72.1035 1.7410 73.1970 ;
        RECT 1.6070 72.1035 1.6330 73.1970 ;
        RECT 1.4990 72.1035 1.5250 73.1970 ;
        RECT 1.3910 72.1035 1.4170 73.1970 ;
        RECT 1.2830 72.1035 1.3090 73.1970 ;
        RECT 1.1750 72.1035 1.2010 73.1970 ;
        RECT 1.0670 72.1035 1.0930 73.1970 ;
        RECT 0.9590 72.1035 0.9850 73.1970 ;
        RECT 0.8510 72.1035 0.8770 73.1970 ;
        RECT 0.7430 72.1035 0.7690 73.1970 ;
        RECT 0.6350 72.1035 0.6610 73.1970 ;
        RECT 0.5270 72.1035 0.5530 73.1970 ;
        RECT 0.4190 72.1035 0.4450 73.1970 ;
        RECT 0.3110 72.1035 0.3370 73.1970 ;
        RECT 0.2030 72.1035 0.2290 73.1970 ;
        RECT 0.0000 72.1035 0.0850 73.1970 ;
        RECT 5.1800 73.1835 5.3080 74.2770 ;
        RECT 5.1660 73.8490 5.3080 74.1715 ;
        RECT 5.0180 73.5760 5.0800 74.2770 ;
        RECT 5.0040 73.8855 5.0800 74.0390 ;
        RECT 5.0180 73.1835 5.0440 74.2770 ;
        RECT 5.0180 73.3045 5.0580 73.5440 ;
        RECT 5.0180 73.1835 5.0800 73.2725 ;
        RECT 4.7210 73.6340 4.9270 74.2770 ;
        RECT 4.9010 73.1835 4.9270 74.2770 ;
        RECT 4.7210 73.9110 4.9410 74.1690 ;
        RECT 4.7210 73.1835 4.8190 74.2770 ;
        RECT 4.3040 73.1835 4.3870 74.2770 ;
        RECT 4.3040 73.2720 4.4010 74.2075 ;
        RECT 9.5270 73.1835 9.6120 74.2770 ;
        RECT 9.3830 73.1835 9.4090 74.2770 ;
        RECT 9.2750 73.1835 9.3010 74.2770 ;
        RECT 9.1670 73.1835 9.1930 74.2770 ;
        RECT 9.0590 73.1835 9.0850 74.2770 ;
        RECT 8.9510 73.1835 8.9770 74.2770 ;
        RECT 8.8430 73.1835 8.8690 74.2770 ;
        RECT 8.7350 73.1835 8.7610 74.2770 ;
        RECT 8.6270 73.1835 8.6530 74.2770 ;
        RECT 8.5190 73.1835 8.5450 74.2770 ;
        RECT 8.4110 73.1835 8.4370 74.2770 ;
        RECT 8.3030 73.1835 8.3290 74.2770 ;
        RECT 8.1950 73.1835 8.2210 74.2770 ;
        RECT 8.0870 73.1835 8.1130 74.2770 ;
        RECT 7.9790 73.1835 8.0050 74.2770 ;
        RECT 7.8710 73.1835 7.8970 74.2770 ;
        RECT 7.7630 73.1835 7.7890 74.2770 ;
        RECT 7.6550 73.1835 7.6810 74.2770 ;
        RECT 7.5470 73.1835 7.5730 74.2770 ;
        RECT 7.4390 73.1835 7.4650 74.2770 ;
        RECT 7.3310 73.1835 7.3570 74.2770 ;
        RECT 7.2230 73.1835 7.2490 74.2770 ;
        RECT 7.1150 73.1835 7.1410 74.2770 ;
        RECT 7.0070 73.1835 7.0330 74.2770 ;
        RECT 6.8990 73.1835 6.9250 74.2770 ;
        RECT 6.7910 73.1835 6.8170 74.2770 ;
        RECT 6.6830 73.1835 6.7090 74.2770 ;
        RECT 6.5750 73.1835 6.6010 74.2770 ;
        RECT 6.4670 73.1835 6.4930 74.2770 ;
        RECT 6.3590 73.1835 6.3850 74.2770 ;
        RECT 6.2510 73.1835 6.2770 74.2770 ;
        RECT 6.1430 73.1835 6.1690 74.2770 ;
        RECT 6.0350 73.1835 6.0610 74.2770 ;
        RECT 5.9270 73.1835 5.9530 74.2770 ;
        RECT 5.7140 73.1835 5.7910 74.2770 ;
        RECT 3.8210 73.1835 3.8980 74.2770 ;
        RECT 3.6590 73.1835 3.6850 74.2770 ;
        RECT 3.5510 73.1835 3.5770 74.2770 ;
        RECT 3.4430 73.1835 3.4690 74.2770 ;
        RECT 3.3350 73.1835 3.3610 74.2770 ;
        RECT 3.2270 73.1835 3.2530 74.2770 ;
        RECT 3.1190 73.1835 3.1450 74.2770 ;
        RECT 3.0110 73.1835 3.0370 74.2770 ;
        RECT 2.9030 73.1835 2.9290 74.2770 ;
        RECT 2.7950 73.1835 2.8210 74.2770 ;
        RECT 2.6870 73.1835 2.7130 74.2770 ;
        RECT 2.5790 73.1835 2.6050 74.2770 ;
        RECT 2.4710 73.1835 2.4970 74.2770 ;
        RECT 2.3630 73.1835 2.3890 74.2770 ;
        RECT 2.2550 73.1835 2.2810 74.2770 ;
        RECT 2.1470 73.1835 2.1730 74.2770 ;
        RECT 2.0390 73.1835 2.0650 74.2770 ;
        RECT 1.9310 73.1835 1.9570 74.2770 ;
        RECT 1.8230 73.1835 1.8490 74.2770 ;
        RECT 1.7150 73.1835 1.7410 74.2770 ;
        RECT 1.6070 73.1835 1.6330 74.2770 ;
        RECT 1.4990 73.1835 1.5250 74.2770 ;
        RECT 1.3910 73.1835 1.4170 74.2770 ;
        RECT 1.2830 73.1835 1.3090 74.2770 ;
        RECT 1.1750 73.1835 1.2010 74.2770 ;
        RECT 1.0670 73.1835 1.0930 74.2770 ;
        RECT 0.9590 73.1835 0.9850 74.2770 ;
        RECT 0.8510 73.1835 0.8770 74.2770 ;
        RECT 0.7430 73.1835 0.7690 74.2770 ;
        RECT 0.6350 73.1835 0.6610 74.2770 ;
        RECT 0.5270 73.1835 0.5530 74.2770 ;
        RECT 0.4190 73.1835 0.4450 74.2770 ;
        RECT 0.3110 73.1835 0.3370 74.2770 ;
        RECT 0.2030 73.1835 0.2290 74.2770 ;
        RECT 0.0000 73.1835 0.0850 74.2770 ;
        RECT 5.1800 74.2635 5.3080 75.3570 ;
        RECT 5.1660 74.9290 5.3080 75.2515 ;
        RECT 5.0180 74.6560 5.0800 75.3570 ;
        RECT 5.0040 74.9655 5.0800 75.1190 ;
        RECT 5.0180 74.2635 5.0440 75.3570 ;
        RECT 5.0180 74.3845 5.0580 74.6240 ;
        RECT 5.0180 74.2635 5.0800 74.3525 ;
        RECT 4.7210 74.7140 4.9270 75.3570 ;
        RECT 4.9010 74.2635 4.9270 75.3570 ;
        RECT 4.7210 74.9910 4.9410 75.2490 ;
        RECT 4.7210 74.2635 4.8190 75.3570 ;
        RECT 4.3040 74.2635 4.3870 75.3570 ;
        RECT 4.3040 74.3520 4.4010 75.2875 ;
        RECT 9.5270 74.2635 9.6120 75.3570 ;
        RECT 9.3830 74.2635 9.4090 75.3570 ;
        RECT 9.2750 74.2635 9.3010 75.3570 ;
        RECT 9.1670 74.2635 9.1930 75.3570 ;
        RECT 9.0590 74.2635 9.0850 75.3570 ;
        RECT 8.9510 74.2635 8.9770 75.3570 ;
        RECT 8.8430 74.2635 8.8690 75.3570 ;
        RECT 8.7350 74.2635 8.7610 75.3570 ;
        RECT 8.6270 74.2635 8.6530 75.3570 ;
        RECT 8.5190 74.2635 8.5450 75.3570 ;
        RECT 8.4110 74.2635 8.4370 75.3570 ;
        RECT 8.3030 74.2635 8.3290 75.3570 ;
        RECT 8.1950 74.2635 8.2210 75.3570 ;
        RECT 8.0870 74.2635 8.1130 75.3570 ;
        RECT 7.9790 74.2635 8.0050 75.3570 ;
        RECT 7.8710 74.2635 7.8970 75.3570 ;
        RECT 7.7630 74.2635 7.7890 75.3570 ;
        RECT 7.6550 74.2635 7.6810 75.3570 ;
        RECT 7.5470 74.2635 7.5730 75.3570 ;
        RECT 7.4390 74.2635 7.4650 75.3570 ;
        RECT 7.3310 74.2635 7.3570 75.3570 ;
        RECT 7.2230 74.2635 7.2490 75.3570 ;
        RECT 7.1150 74.2635 7.1410 75.3570 ;
        RECT 7.0070 74.2635 7.0330 75.3570 ;
        RECT 6.8990 74.2635 6.9250 75.3570 ;
        RECT 6.7910 74.2635 6.8170 75.3570 ;
        RECT 6.6830 74.2635 6.7090 75.3570 ;
        RECT 6.5750 74.2635 6.6010 75.3570 ;
        RECT 6.4670 74.2635 6.4930 75.3570 ;
        RECT 6.3590 74.2635 6.3850 75.3570 ;
        RECT 6.2510 74.2635 6.2770 75.3570 ;
        RECT 6.1430 74.2635 6.1690 75.3570 ;
        RECT 6.0350 74.2635 6.0610 75.3570 ;
        RECT 5.9270 74.2635 5.9530 75.3570 ;
        RECT 5.7140 74.2635 5.7910 75.3570 ;
        RECT 3.8210 74.2635 3.8980 75.3570 ;
        RECT 3.6590 74.2635 3.6850 75.3570 ;
        RECT 3.5510 74.2635 3.5770 75.3570 ;
        RECT 3.4430 74.2635 3.4690 75.3570 ;
        RECT 3.3350 74.2635 3.3610 75.3570 ;
        RECT 3.2270 74.2635 3.2530 75.3570 ;
        RECT 3.1190 74.2635 3.1450 75.3570 ;
        RECT 3.0110 74.2635 3.0370 75.3570 ;
        RECT 2.9030 74.2635 2.9290 75.3570 ;
        RECT 2.7950 74.2635 2.8210 75.3570 ;
        RECT 2.6870 74.2635 2.7130 75.3570 ;
        RECT 2.5790 74.2635 2.6050 75.3570 ;
        RECT 2.4710 74.2635 2.4970 75.3570 ;
        RECT 2.3630 74.2635 2.3890 75.3570 ;
        RECT 2.2550 74.2635 2.2810 75.3570 ;
        RECT 2.1470 74.2635 2.1730 75.3570 ;
        RECT 2.0390 74.2635 2.0650 75.3570 ;
        RECT 1.9310 74.2635 1.9570 75.3570 ;
        RECT 1.8230 74.2635 1.8490 75.3570 ;
        RECT 1.7150 74.2635 1.7410 75.3570 ;
        RECT 1.6070 74.2635 1.6330 75.3570 ;
        RECT 1.4990 74.2635 1.5250 75.3570 ;
        RECT 1.3910 74.2635 1.4170 75.3570 ;
        RECT 1.2830 74.2635 1.3090 75.3570 ;
        RECT 1.1750 74.2635 1.2010 75.3570 ;
        RECT 1.0670 74.2635 1.0930 75.3570 ;
        RECT 0.9590 74.2635 0.9850 75.3570 ;
        RECT 0.8510 74.2635 0.8770 75.3570 ;
        RECT 0.7430 74.2635 0.7690 75.3570 ;
        RECT 0.6350 74.2635 0.6610 75.3570 ;
        RECT 0.5270 74.2635 0.5530 75.3570 ;
        RECT 0.4190 74.2635 0.4450 75.3570 ;
        RECT 0.3110 74.2635 0.3370 75.3570 ;
        RECT 0.2030 74.2635 0.2290 75.3570 ;
        RECT 0.0000 74.2635 0.0850 75.3570 ;
        RECT 5.1800 75.3435 5.3080 76.4370 ;
        RECT 5.1660 76.0090 5.3080 76.3315 ;
        RECT 5.0180 75.7360 5.0800 76.4370 ;
        RECT 5.0040 76.0455 5.0800 76.1990 ;
        RECT 5.0180 75.3435 5.0440 76.4370 ;
        RECT 5.0180 75.4645 5.0580 75.7040 ;
        RECT 5.0180 75.3435 5.0800 75.4325 ;
        RECT 4.7210 75.7940 4.9270 76.4370 ;
        RECT 4.9010 75.3435 4.9270 76.4370 ;
        RECT 4.7210 76.0710 4.9410 76.3290 ;
        RECT 4.7210 75.3435 4.8190 76.4370 ;
        RECT 4.3040 75.3435 4.3870 76.4370 ;
        RECT 4.3040 75.4320 4.4010 76.3675 ;
        RECT 9.5270 75.3435 9.6120 76.4370 ;
        RECT 9.3830 75.3435 9.4090 76.4370 ;
        RECT 9.2750 75.3435 9.3010 76.4370 ;
        RECT 9.1670 75.3435 9.1930 76.4370 ;
        RECT 9.0590 75.3435 9.0850 76.4370 ;
        RECT 8.9510 75.3435 8.9770 76.4370 ;
        RECT 8.8430 75.3435 8.8690 76.4370 ;
        RECT 8.7350 75.3435 8.7610 76.4370 ;
        RECT 8.6270 75.3435 8.6530 76.4370 ;
        RECT 8.5190 75.3435 8.5450 76.4370 ;
        RECT 8.4110 75.3435 8.4370 76.4370 ;
        RECT 8.3030 75.3435 8.3290 76.4370 ;
        RECT 8.1950 75.3435 8.2210 76.4370 ;
        RECT 8.0870 75.3435 8.1130 76.4370 ;
        RECT 7.9790 75.3435 8.0050 76.4370 ;
        RECT 7.8710 75.3435 7.8970 76.4370 ;
        RECT 7.7630 75.3435 7.7890 76.4370 ;
        RECT 7.6550 75.3435 7.6810 76.4370 ;
        RECT 7.5470 75.3435 7.5730 76.4370 ;
        RECT 7.4390 75.3435 7.4650 76.4370 ;
        RECT 7.3310 75.3435 7.3570 76.4370 ;
        RECT 7.2230 75.3435 7.2490 76.4370 ;
        RECT 7.1150 75.3435 7.1410 76.4370 ;
        RECT 7.0070 75.3435 7.0330 76.4370 ;
        RECT 6.8990 75.3435 6.9250 76.4370 ;
        RECT 6.7910 75.3435 6.8170 76.4370 ;
        RECT 6.6830 75.3435 6.7090 76.4370 ;
        RECT 6.5750 75.3435 6.6010 76.4370 ;
        RECT 6.4670 75.3435 6.4930 76.4370 ;
        RECT 6.3590 75.3435 6.3850 76.4370 ;
        RECT 6.2510 75.3435 6.2770 76.4370 ;
        RECT 6.1430 75.3435 6.1690 76.4370 ;
        RECT 6.0350 75.3435 6.0610 76.4370 ;
        RECT 5.9270 75.3435 5.9530 76.4370 ;
        RECT 5.7140 75.3435 5.7910 76.4370 ;
        RECT 3.8210 75.3435 3.8980 76.4370 ;
        RECT 3.6590 75.3435 3.6850 76.4370 ;
        RECT 3.5510 75.3435 3.5770 76.4370 ;
        RECT 3.4430 75.3435 3.4690 76.4370 ;
        RECT 3.3350 75.3435 3.3610 76.4370 ;
        RECT 3.2270 75.3435 3.2530 76.4370 ;
        RECT 3.1190 75.3435 3.1450 76.4370 ;
        RECT 3.0110 75.3435 3.0370 76.4370 ;
        RECT 2.9030 75.3435 2.9290 76.4370 ;
        RECT 2.7950 75.3435 2.8210 76.4370 ;
        RECT 2.6870 75.3435 2.7130 76.4370 ;
        RECT 2.5790 75.3435 2.6050 76.4370 ;
        RECT 2.4710 75.3435 2.4970 76.4370 ;
        RECT 2.3630 75.3435 2.3890 76.4370 ;
        RECT 2.2550 75.3435 2.2810 76.4370 ;
        RECT 2.1470 75.3435 2.1730 76.4370 ;
        RECT 2.0390 75.3435 2.0650 76.4370 ;
        RECT 1.9310 75.3435 1.9570 76.4370 ;
        RECT 1.8230 75.3435 1.8490 76.4370 ;
        RECT 1.7150 75.3435 1.7410 76.4370 ;
        RECT 1.6070 75.3435 1.6330 76.4370 ;
        RECT 1.4990 75.3435 1.5250 76.4370 ;
        RECT 1.3910 75.3435 1.4170 76.4370 ;
        RECT 1.2830 75.3435 1.3090 76.4370 ;
        RECT 1.1750 75.3435 1.2010 76.4370 ;
        RECT 1.0670 75.3435 1.0930 76.4370 ;
        RECT 0.9590 75.3435 0.9850 76.4370 ;
        RECT 0.8510 75.3435 0.8770 76.4370 ;
        RECT 0.7430 75.3435 0.7690 76.4370 ;
        RECT 0.6350 75.3435 0.6610 76.4370 ;
        RECT 0.5270 75.3435 0.5530 76.4370 ;
        RECT 0.4190 75.3435 0.4450 76.4370 ;
        RECT 0.3110 75.3435 0.3370 76.4370 ;
        RECT 0.2030 75.3435 0.2290 76.4370 ;
        RECT 0.0000 75.3435 0.0850 76.4370 ;
        RECT 5.1800 76.4235 5.3080 77.5170 ;
        RECT 5.1660 77.0890 5.3080 77.4115 ;
        RECT 5.0180 76.8160 5.0800 77.5170 ;
        RECT 5.0040 77.1255 5.0800 77.2790 ;
        RECT 5.0180 76.4235 5.0440 77.5170 ;
        RECT 5.0180 76.5445 5.0580 76.7840 ;
        RECT 5.0180 76.4235 5.0800 76.5125 ;
        RECT 4.7210 76.8740 4.9270 77.5170 ;
        RECT 4.9010 76.4235 4.9270 77.5170 ;
        RECT 4.7210 77.1510 4.9410 77.4090 ;
        RECT 4.7210 76.4235 4.8190 77.5170 ;
        RECT 4.3040 76.4235 4.3870 77.5170 ;
        RECT 4.3040 76.5120 4.4010 77.4475 ;
        RECT 9.5270 76.4235 9.6120 77.5170 ;
        RECT 9.3830 76.4235 9.4090 77.5170 ;
        RECT 9.2750 76.4235 9.3010 77.5170 ;
        RECT 9.1670 76.4235 9.1930 77.5170 ;
        RECT 9.0590 76.4235 9.0850 77.5170 ;
        RECT 8.9510 76.4235 8.9770 77.5170 ;
        RECT 8.8430 76.4235 8.8690 77.5170 ;
        RECT 8.7350 76.4235 8.7610 77.5170 ;
        RECT 8.6270 76.4235 8.6530 77.5170 ;
        RECT 8.5190 76.4235 8.5450 77.5170 ;
        RECT 8.4110 76.4235 8.4370 77.5170 ;
        RECT 8.3030 76.4235 8.3290 77.5170 ;
        RECT 8.1950 76.4235 8.2210 77.5170 ;
        RECT 8.0870 76.4235 8.1130 77.5170 ;
        RECT 7.9790 76.4235 8.0050 77.5170 ;
        RECT 7.8710 76.4235 7.8970 77.5170 ;
        RECT 7.7630 76.4235 7.7890 77.5170 ;
        RECT 7.6550 76.4235 7.6810 77.5170 ;
        RECT 7.5470 76.4235 7.5730 77.5170 ;
        RECT 7.4390 76.4235 7.4650 77.5170 ;
        RECT 7.3310 76.4235 7.3570 77.5170 ;
        RECT 7.2230 76.4235 7.2490 77.5170 ;
        RECT 7.1150 76.4235 7.1410 77.5170 ;
        RECT 7.0070 76.4235 7.0330 77.5170 ;
        RECT 6.8990 76.4235 6.9250 77.5170 ;
        RECT 6.7910 76.4235 6.8170 77.5170 ;
        RECT 6.6830 76.4235 6.7090 77.5170 ;
        RECT 6.5750 76.4235 6.6010 77.5170 ;
        RECT 6.4670 76.4235 6.4930 77.5170 ;
        RECT 6.3590 76.4235 6.3850 77.5170 ;
        RECT 6.2510 76.4235 6.2770 77.5170 ;
        RECT 6.1430 76.4235 6.1690 77.5170 ;
        RECT 6.0350 76.4235 6.0610 77.5170 ;
        RECT 5.9270 76.4235 5.9530 77.5170 ;
        RECT 5.7140 76.4235 5.7910 77.5170 ;
        RECT 3.8210 76.4235 3.8980 77.5170 ;
        RECT 3.6590 76.4235 3.6850 77.5170 ;
        RECT 3.5510 76.4235 3.5770 77.5170 ;
        RECT 3.4430 76.4235 3.4690 77.5170 ;
        RECT 3.3350 76.4235 3.3610 77.5170 ;
        RECT 3.2270 76.4235 3.2530 77.5170 ;
        RECT 3.1190 76.4235 3.1450 77.5170 ;
        RECT 3.0110 76.4235 3.0370 77.5170 ;
        RECT 2.9030 76.4235 2.9290 77.5170 ;
        RECT 2.7950 76.4235 2.8210 77.5170 ;
        RECT 2.6870 76.4235 2.7130 77.5170 ;
        RECT 2.5790 76.4235 2.6050 77.5170 ;
        RECT 2.4710 76.4235 2.4970 77.5170 ;
        RECT 2.3630 76.4235 2.3890 77.5170 ;
        RECT 2.2550 76.4235 2.2810 77.5170 ;
        RECT 2.1470 76.4235 2.1730 77.5170 ;
        RECT 2.0390 76.4235 2.0650 77.5170 ;
        RECT 1.9310 76.4235 1.9570 77.5170 ;
        RECT 1.8230 76.4235 1.8490 77.5170 ;
        RECT 1.7150 76.4235 1.7410 77.5170 ;
        RECT 1.6070 76.4235 1.6330 77.5170 ;
        RECT 1.4990 76.4235 1.5250 77.5170 ;
        RECT 1.3910 76.4235 1.4170 77.5170 ;
        RECT 1.2830 76.4235 1.3090 77.5170 ;
        RECT 1.1750 76.4235 1.2010 77.5170 ;
        RECT 1.0670 76.4235 1.0930 77.5170 ;
        RECT 0.9590 76.4235 0.9850 77.5170 ;
        RECT 0.8510 76.4235 0.8770 77.5170 ;
        RECT 0.7430 76.4235 0.7690 77.5170 ;
        RECT 0.6350 76.4235 0.6610 77.5170 ;
        RECT 0.5270 76.4235 0.5530 77.5170 ;
        RECT 0.4190 76.4235 0.4450 77.5170 ;
        RECT 0.3110 76.4235 0.3370 77.5170 ;
        RECT 0.2030 76.4235 0.2290 77.5170 ;
        RECT 0.0000 76.4235 0.0850 77.5170 ;
        RECT 5.1800 77.5035 5.3080 78.5970 ;
        RECT 5.1660 78.1690 5.3080 78.4915 ;
        RECT 5.0180 77.8960 5.0800 78.5970 ;
        RECT 5.0040 78.2055 5.0800 78.3590 ;
        RECT 5.0180 77.5035 5.0440 78.5970 ;
        RECT 5.0180 77.6245 5.0580 77.8640 ;
        RECT 5.0180 77.5035 5.0800 77.5925 ;
        RECT 4.7210 77.9540 4.9270 78.5970 ;
        RECT 4.9010 77.5035 4.9270 78.5970 ;
        RECT 4.7210 78.2310 4.9410 78.4890 ;
        RECT 4.7210 77.5035 4.8190 78.5970 ;
        RECT 4.3040 77.5035 4.3870 78.5970 ;
        RECT 4.3040 77.5920 4.4010 78.5275 ;
        RECT 9.5270 77.5035 9.6120 78.5970 ;
        RECT 9.3830 77.5035 9.4090 78.5970 ;
        RECT 9.2750 77.5035 9.3010 78.5970 ;
        RECT 9.1670 77.5035 9.1930 78.5970 ;
        RECT 9.0590 77.5035 9.0850 78.5970 ;
        RECT 8.9510 77.5035 8.9770 78.5970 ;
        RECT 8.8430 77.5035 8.8690 78.5970 ;
        RECT 8.7350 77.5035 8.7610 78.5970 ;
        RECT 8.6270 77.5035 8.6530 78.5970 ;
        RECT 8.5190 77.5035 8.5450 78.5970 ;
        RECT 8.4110 77.5035 8.4370 78.5970 ;
        RECT 8.3030 77.5035 8.3290 78.5970 ;
        RECT 8.1950 77.5035 8.2210 78.5970 ;
        RECT 8.0870 77.5035 8.1130 78.5970 ;
        RECT 7.9790 77.5035 8.0050 78.5970 ;
        RECT 7.8710 77.5035 7.8970 78.5970 ;
        RECT 7.7630 77.5035 7.7890 78.5970 ;
        RECT 7.6550 77.5035 7.6810 78.5970 ;
        RECT 7.5470 77.5035 7.5730 78.5970 ;
        RECT 7.4390 77.5035 7.4650 78.5970 ;
        RECT 7.3310 77.5035 7.3570 78.5970 ;
        RECT 7.2230 77.5035 7.2490 78.5970 ;
        RECT 7.1150 77.5035 7.1410 78.5970 ;
        RECT 7.0070 77.5035 7.0330 78.5970 ;
        RECT 6.8990 77.5035 6.9250 78.5970 ;
        RECT 6.7910 77.5035 6.8170 78.5970 ;
        RECT 6.6830 77.5035 6.7090 78.5970 ;
        RECT 6.5750 77.5035 6.6010 78.5970 ;
        RECT 6.4670 77.5035 6.4930 78.5970 ;
        RECT 6.3590 77.5035 6.3850 78.5970 ;
        RECT 6.2510 77.5035 6.2770 78.5970 ;
        RECT 6.1430 77.5035 6.1690 78.5970 ;
        RECT 6.0350 77.5035 6.0610 78.5970 ;
        RECT 5.9270 77.5035 5.9530 78.5970 ;
        RECT 5.7140 77.5035 5.7910 78.5970 ;
        RECT 3.8210 77.5035 3.8980 78.5970 ;
        RECT 3.6590 77.5035 3.6850 78.5970 ;
        RECT 3.5510 77.5035 3.5770 78.5970 ;
        RECT 3.4430 77.5035 3.4690 78.5970 ;
        RECT 3.3350 77.5035 3.3610 78.5970 ;
        RECT 3.2270 77.5035 3.2530 78.5970 ;
        RECT 3.1190 77.5035 3.1450 78.5970 ;
        RECT 3.0110 77.5035 3.0370 78.5970 ;
        RECT 2.9030 77.5035 2.9290 78.5970 ;
        RECT 2.7950 77.5035 2.8210 78.5970 ;
        RECT 2.6870 77.5035 2.7130 78.5970 ;
        RECT 2.5790 77.5035 2.6050 78.5970 ;
        RECT 2.4710 77.5035 2.4970 78.5970 ;
        RECT 2.3630 77.5035 2.3890 78.5970 ;
        RECT 2.2550 77.5035 2.2810 78.5970 ;
        RECT 2.1470 77.5035 2.1730 78.5970 ;
        RECT 2.0390 77.5035 2.0650 78.5970 ;
        RECT 1.9310 77.5035 1.9570 78.5970 ;
        RECT 1.8230 77.5035 1.8490 78.5970 ;
        RECT 1.7150 77.5035 1.7410 78.5970 ;
        RECT 1.6070 77.5035 1.6330 78.5970 ;
        RECT 1.4990 77.5035 1.5250 78.5970 ;
        RECT 1.3910 77.5035 1.4170 78.5970 ;
        RECT 1.2830 77.5035 1.3090 78.5970 ;
        RECT 1.1750 77.5035 1.2010 78.5970 ;
        RECT 1.0670 77.5035 1.0930 78.5970 ;
        RECT 0.9590 77.5035 0.9850 78.5970 ;
        RECT 0.8510 77.5035 0.8770 78.5970 ;
        RECT 0.7430 77.5035 0.7690 78.5970 ;
        RECT 0.6350 77.5035 0.6610 78.5970 ;
        RECT 0.5270 77.5035 0.5530 78.5970 ;
        RECT 0.4190 77.5035 0.4450 78.5970 ;
        RECT 0.3110 77.5035 0.3370 78.5970 ;
        RECT 0.2030 77.5035 0.2290 78.5970 ;
        RECT 0.0000 77.5035 0.0850 78.5970 ;
        RECT 5.1800 78.5835 5.3080 79.6770 ;
        RECT 5.1660 79.2490 5.3080 79.5715 ;
        RECT 5.0180 78.9760 5.0800 79.6770 ;
        RECT 5.0040 79.2855 5.0800 79.4390 ;
        RECT 5.0180 78.5835 5.0440 79.6770 ;
        RECT 5.0180 78.7045 5.0580 78.9440 ;
        RECT 5.0180 78.5835 5.0800 78.6725 ;
        RECT 4.7210 79.0340 4.9270 79.6770 ;
        RECT 4.9010 78.5835 4.9270 79.6770 ;
        RECT 4.7210 79.3110 4.9410 79.5690 ;
        RECT 4.7210 78.5835 4.8190 79.6770 ;
        RECT 4.3040 78.5835 4.3870 79.6770 ;
        RECT 4.3040 78.6720 4.4010 79.6075 ;
        RECT 9.5270 78.5835 9.6120 79.6770 ;
        RECT 9.3830 78.5835 9.4090 79.6770 ;
        RECT 9.2750 78.5835 9.3010 79.6770 ;
        RECT 9.1670 78.5835 9.1930 79.6770 ;
        RECT 9.0590 78.5835 9.0850 79.6770 ;
        RECT 8.9510 78.5835 8.9770 79.6770 ;
        RECT 8.8430 78.5835 8.8690 79.6770 ;
        RECT 8.7350 78.5835 8.7610 79.6770 ;
        RECT 8.6270 78.5835 8.6530 79.6770 ;
        RECT 8.5190 78.5835 8.5450 79.6770 ;
        RECT 8.4110 78.5835 8.4370 79.6770 ;
        RECT 8.3030 78.5835 8.3290 79.6770 ;
        RECT 8.1950 78.5835 8.2210 79.6770 ;
        RECT 8.0870 78.5835 8.1130 79.6770 ;
        RECT 7.9790 78.5835 8.0050 79.6770 ;
        RECT 7.8710 78.5835 7.8970 79.6770 ;
        RECT 7.7630 78.5835 7.7890 79.6770 ;
        RECT 7.6550 78.5835 7.6810 79.6770 ;
        RECT 7.5470 78.5835 7.5730 79.6770 ;
        RECT 7.4390 78.5835 7.4650 79.6770 ;
        RECT 7.3310 78.5835 7.3570 79.6770 ;
        RECT 7.2230 78.5835 7.2490 79.6770 ;
        RECT 7.1150 78.5835 7.1410 79.6770 ;
        RECT 7.0070 78.5835 7.0330 79.6770 ;
        RECT 6.8990 78.5835 6.9250 79.6770 ;
        RECT 6.7910 78.5835 6.8170 79.6770 ;
        RECT 6.6830 78.5835 6.7090 79.6770 ;
        RECT 6.5750 78.5835 6.6010 79.6770 ;
        RECT 6.4670 78.5835 6.4930 79.6770 ;
        RECT 6.3590 78.5835 6.3850 79.6770 ;
        RECT 6.2510 78.5835 6.2770 79.6770 ;
        RECT 6.1430 78.5835 6.1690 79.6770 ;
        RECT 6.0350 78.5835 6.0610 79.6770 ;
        RECT 5.9270 78.5835 5.9530 79.6770 ;
        RECT 5.7140 78.5835 5.7910 79.6770 ;
        RECT 3.8210 78.5835 3.8980 79.6770 ;
        RECT 3.6590 78.5835 3.6850 79.6770 ;
        RECT 3.5510 78.5835 3.5770 79.6770 ;
        RECT 3.4430 78.5835 3.4690 79.6770 ;
        RECT 3.3350 78.5835 3.3610 79.6770 ;
        RECT 3.2270 78.5835 3.2530 79.6770 ;
        RECT 3.1190 78.5835 3.1450 79.6770 ;
        RECT 3.0110 78.5835 3.0370 79.6770 ;
        RECT 2.9030 78.5835 2.9290 79.6770 ;
        RECT 2.7950 78.5835 2.8210 79.6770 ;
        RECT 2.6870 78.5835 2.7130 79.6770 ;
        RECT 2.5790 78.5835 2.6050 79.6770 ;
        RECT 2.4710 78.5835 2.4970 79.6770 ;
        RECT 2.3630 78.5835 2.3890 79.6770 ;
        RECT 2.2550 78.5835 2.2810 79.6770 ;
        RECT 2.1470 78.5835 2.1730 79.6770 ;
        RECT 2.0390 78.5835 2.0650 79.6770 ;
        RECT 1.9310 78.5835 1.9570 79.6770 ;
        RECT 1.8230 78.5835 1.8490 79.6770 ;
        RECT 1.7150 78.5835 1.7410 79.6770 ;
        RECT 1.6070 78.5835 1.6330 79.6770 ;
        RECT 1.4990 78.5835 1.5250 79.6770 ;
        RECT 1.3910 78.5835 1.4170 79.6770 ;
        RECT 1.2830 78.5835 1.3090 79.6770 ;
        RECT 1.1750 78.5835 1.2010 79.6770 ;
        RECT 1.0670 78.5835 1.0930 79.6770 ;
        RECT 0.9590 78.5835 0.9850 79.6770 ;
        RECT 0.8510 78.5835 0.8770 79.6770 ;
        RECT 0.7430 78.5835 0.7690 79.6770 ;
        RECT 0.6350 78.5835 0.6610 79.6770 ;
        RECT 0.5270 78.5835 0.5530 79.6770 ;
        RECT 0.4190 78.5835 0.4450 79.6770 ;
        RECT 0.3110 78.5835 0.3370 79.6770 ;
        RECT 0.2030 78.5835 0.2290 79.6770 ;
        RECT 0.0000 78.5835 0.0850 79.6770 ;
        RECT 5.1800 79.6635 5.3080 80.7570 ;
        RECT 5.1660 80.3290 5.3080 80.6515 ;
        RECT 5.0180 80.0560 5.0800 80.7570 ;
        RECT 5.0040 80.3655 5.0800 80.5190 ;
        RECT 5.0180 79.6635 5.0440 80.7570 ;
        RECT 5.0180 79.7845 5.0580 80.0240 ;
        RECT 5.0180 79.6635 5.0800 79.7525 ;
        RECT 4.7210 80.1140 4.9270 80.7570 ;
        RECT 4.9010 79.6635 4.9270 80.7570 ;
        RECT 4.7210 80.3910 4.9410 80.6490 ;
        RECT 4.7210 79.6635 4.8190 80.7570 ;
        RECT 4.3040 79.6635 4.3870 80.7570 ;
        RECT 4.3040 79.7520 4.4010 80.6875 ;
        RECT 9.5270 79.6635 9.6120 80.7570 ;
        RECT 9.3830 79.6635 9.4090 80.7570 ;
        RECT 9.2750 79.6635 9.3010 80.7570 ;
        RECT 9.1670 79.6635 9.1930 80.7570 ;
        RECT 9.0590 79.6635 9.0850 80.7570 ;
        RECT 8.9510 79.6635 8.9770 80.7570 ;
        RECT 8.8430 79.6635 8.8690 80.7570 ;
        RECT 8.7350 79.6635 8.7610 80.7570 ;
        RECT 8.6270 79.6635 8.6530 80.7570 ;
        RECT 8.5190 79.6635 8.5450 80.7570 ;
        RECT 8.4110 79.6635 8.4370 80.7570 ;
        RECT 8.3030 79.6635 8.3290 80.7570 ;
        RECT 8.1950 79.6635 8.2210 80.7570 ;
        RECT 8.0870 79.6635 8.1130 80.7570 ;
        RECT 7.9790 79.6635 8.0050 80.7570 ;
        RECT 7.8710 79.6635 7.8970 80.7570 ;
        RECT 7.7630 79.6635 7.7890 80.7570 ;
        RECT 7.6550 79.6635 7.6810 80.7570 ;
        RECT 7.5470 79.6635 7.5730 80.7570 ;
        RECT 7.4390 79.6635 7.4650 80.7570 ;
        RECT 7.3310 79.6635 7.3570 80.7570 ;
        RECT 7.2230 79.6635 7.2490 80.7570 ;
        RECT 7.1150 79.6635 7.1410 80.7570 ;
        RECT 7.0070 79.6635 7.0330 80.7570 ;
        RECT 6.8990 79.6635 6.9250 80.7570 ;
        RECT 6.7910 79.6635 6.8170 80.7570 ;
        RECT 6.6830 79.6635 6.7090 80.7570 ;
        RECT 6.5750 79.6635 6.6010 80.7570 ;
        RECT 6.4670 79.6635 6.4930 80.7570 ;
        RECT 6.3590 79.6635 6.3850 80.7570 ;
        RECT 6.2510 79.6635 6.2770 80.7570 ;
        RECT 6.1430 79.6635 6.1690 80.7570 ;
        RECT 6.0350 79.6635 6.0610 80.7570 ;
        RECT 5.9270 79.6635 5.9530 80.7570 ;
        RECT 5.7140 79.6635 5.7910 80.7570 ;
        RECT 3.8210 79.6635 3.8980 80.7570 ;
        RECT 3.6590 79.6635 3.6850 80.7570 ;
        RECT 3.5510 79.6635 3.5770 80.7570 ;
        RECT 3.4430 79.6635 3.4690 80.7570 ;
        RECT 3.3350 79.6635 3.3610 80.7570 ;
        RECT 3.2270 79.6635 3.2530 80.7570 ;
        RECT 3.1190 79.6635 3.1450 80.7570 ;
        RECT 3.0110 79.6635 3.0370 80.7570 ;
        RECT 2.9030 79.6635 2.9290 80.7570 ;
        RECT 2.7950 79.6635 2.8210 80.7570 ;
        RECT 2.6870 79.6635 2.7130 80.7570 ;
        RECT 2.5790 79.6635 2.6050 80.7570 ;
        RECT 2.4710 79.6635 2.4970 80.7570 ;
        RECT 2.3630 79.6635 2.3890 80.7570 ;
        RECT 2.2550 79.6635 2.2810 80.7570 ;
        RECT 2.1470 79.6635 2.1730 80.7570 ;
        RECT 2.0390 79.6635 2.0650 80.7570 ;
        RECT 1.9310 79.6635 1.9570 80.7570 ;
        RECT 1.8230 79.6635 1.8490 80.7570 ;
        RECT 1.7150 79.6635 1.7410 80.7570 ;
        RECT 1.6070 79.6635 1.6330 80.7570 ;
        RECT 1.4990 79.6635 1.5250 80.7570 ;
        RECT 1.3910 79.6635 1.4170 80.7570 ;
        RECT 1.2830 79.6635 1.3090 80.7570 ;
        RECT 1.1750 79.6635 1.2010 80.7570 ;
        RECT 1.0670 79.6635 1.0930 80.7570 ;
        RECT 0.9590 79.6635 0.9850 80.7570 ;
        RECT 0.8510 79.6635 0.8770 80.7570 ;
        RECT 0.7430 79.6635 0.7690 80.7570 ;
        RECT 0.6350 79.6635 0.6610 80.7570 ;
        RECT 0.5270 79.6635 0.5530 80.7570 ;
        RECT 0.4190 79.6635 0.4450 80.7570 ;
        RECT 0.3110 79.6635 0.3370 80.7570 ;
        RECT 0.2030 79.6635 0.2290 80.7570 ;
        RECT 0.0000 79.6635 0.0850 80.7570 ;
        RECT 5.1800 80.7435 5.3080 81.8370 ;
        RECT 5.1660 81.4090 5.3080 81.7315 ;
        RECT 5.0180 81.1360 5.0800 81.8370 ;
        RECT 5.0040 81.4455 5.0800 81.5990 ;
        RECT 5.0180 80.7435 5.0440 81.8370 ;
        RECT 5.0180 80.8645 5.0580 81.1040 ;
        RECT 5.0180 80.7435 5.0800 80.8325 ;
        RECT 4.7210 81.1940 4.9270 81.8370 ;
        RECT 4.9010 80.7435 4.9270 81.8370 ;
        RECT 4.7210 81.4710 4.9410 81.7290 ;
        RECT 4.7210 80.7435 4.8190 81.8370 ;
        RECT 4.3040 80.7435 4.3870 81.8370 ;
        RECT 4.3040 80.8320 4.4010 81.7675 ;
        RECT 9.5270 80.7435 9.6120 81.8370 ;
        RECT 9.3830 80.7435 9.4090 81.8370 ;
        RECT 9.2750 80.7435 9.3010 81.8370 ;
        RECT 9.1670 80.7435 9.1930 81.8370 ;
        RECT 9.0590 80.7435 9.0850 81.8370 ;
        RECT 8.9510 80.7435 8.9770 81.8370 ;
        RECT 8.8430 80.7435 8.8690 81.8370 ;
        RECT 8.7350 80.7435 8.7610 81.8370 ;
        RECT 8.6270 80.7435 8.6530 81.8370 ;
        RECT 8.5190 80.7435 8.5450 81.8370 ;
        RECT 8.4110 80.7435 8.4370 81.8370 ;
        RECT 8.3030 80.7435 8.3290 81.8370 ;
        RECT 8.1950 80.7435 8.2210 81.8370 ;
        RECT 8.0870 80.7435 8.1130 81.8370 ;
        RECT 7.9790 80.7435 8.0050 81.8370 ;
        RECT 7.8710 80.7435 7.8970 81.8370 ;
        RECT 7.7630 80.7435 7.7890 81.8370 ;
        RECT 7.6550 80.7435 7.6810 81.8370 ;
        RECT 7.5470 80.7435 7.5730 81.8370 ;
        RECT 7.4390 80.7435 7.4650 81.8370 ;
        RECT 7.3310 80.7435 7.3570 81.8370 ;
        RECT 7.2230 80.7435 7.2490 81.8370 ;
        RECT 7.1150 80.7435 7.1410 81.8370 ;
        RECT 7.0070 80.7435 7.0330 81.8370 ;
        RECT 6.8990 80.7435 6.9250 81.8370 ;
        RECT 6.7910 80.7435 6.8170 81.8370 ;
        RECT 6.6830 80.7435 6.7090 81.8370 ;
        RECT 6.5750 80.7435 6.6010 81.8370 ;
        RECT 6.4670 80.7435 6.4930 81.8370 ;
        RECT 6.3590 80.7435 6.3850 81.8370 ;
        RECT 6.2510 80.7435 6.2770 81.8370 ;
        RECT 6.1430 80.7435 6.1690 81.8370 ;
        RECT 6.0350 80.7435 6.0610 81.8370 ;
        RECT 5.9270 80.7435 5.9530 81.8370 ;
        RECT 5.7140 80.7435 5.7910 81.8370 ;
        RECT 3.8210 80.7435 3.8980 81.8370 ;
        RECT 3.6590 80.7435 3.6850 81.8370 ;
        RECT 3.5510 80.7435 3.5770 81.8370 ;
        RECT 3.4430 80.7435 3.4690 81.8370 ;
        RECT 3.3350 80.7435 3.3610 81.8370 ;
        RECT 3.2270 80.7435 3.2530 81.8370 ;
        RECT 3.1190 80.7435 3.1450 81.8370 ;
        RECT 3.0110 80.7435 3.0370 81.8370 ;
        RECT 2.9030 80.7435 2.9290 81.8370 ;
        RECT 2.7950 80.7435 2.8210 81.8370 ;
        RECT 2.6870 80.7435 2.7130 81.8370 ;
        RECT 2.5790 80.7435 2.6050 81.8370 ;
        RECT 2.4710 80.7435 2.4970 81.8370 ;
        RECT 2.3630 80.7435 2.3890 81.8370 ;
        RECT 2.2550 80.7435 2.2810 81.8370 ;
        RECT 2.1470 80.7435 2.1730 81.8370 ;
        RECT 2.0390 80.7435 2.0650 81.8370 ;
        RECT 1.9310 80.7435 1.9570 81.8370 ;
        RECT 1.8230 80.7435 1.8490 81.8370 ;
        RECT 1.7150 80.7435 1.7410 81.8370 ;
        RECT 1.6070 80.7435 1.6330 81.8370 ;
        RECT 1.4990 80.7435 1.5250 81.8370 ;
        RECT 1.3910 80.7435 1.4170 81.8370 ;
        RECT 1.2830 80.7435 1.3090 81.8370 ;
        RECT 1.1750 80.7435 1.2010 81.8370 ;
        RECT 1.0670 80.7435 1.0930 81.8370 ;
        RECT 0.9590 80.7435 0.9850 81.8370 ;
        RECT 0.8510 80.7435 0.8770 81.8370 ;
        RECT 0.7430 80.7435 0.7690 81.8370 ;
        RECT 0.6350 80.7435 0.6610 81.8370 ;
        RECT 0.5270 80.7435 0.5530 81.8370 ;
        RECT 0.4190 80.7435 0.4450 81.8370 ;
        RECT 0.3110 80.7435 0.3370 81.8370 ;
        RECT 0.2030 80.7435 0.2290 81.8370 ;
        RECT 0.0000 80.7435 0.0850 81.8370 ;
        RECT 5.1800 81.8235 5.3080 82.9170 ;
        RECT 5.1660 82.4890 5.3080 82.8115 ;
        RECT 5.0180 82.2160 5.0800 82.9170 ;
        RECT 5.0040 82.5255 5.0800 82.6790 ;
        RECT 5.0180 81.8235 5.0440 82.9170 ;
        RECT 5.0180 81.9445 5.0580 82.1840 ;
        RECT 5.0180 81.8235 5.0800 81.9125 ;
        RECT 4.7210 82.2740 4.9270 82.9170 ;
        RECT 4.9010 81.8235 4.9270 82.9170 ;
        RECT 4.7210 82.5510 4.9410 82.8090 ;
        RECT 4.7210 81.8235 4.8190 82.9170 ;
        RECT 4.3040 81.8235 4.3870 82.9170 ;
        RECT 4.3040 81.9120 4.4010 82.8475 ;
        RECT 9.5270 81.8235 9.6120 82.9170 ;
        RECT 9.3830 81.8235 9.4090 82.9170 ;
        RECT 9.2750 81.8235 9.3010 82.9170 ;
        RECT 9.1670 81.8235 9.1930 82.9170 ;
        RECT 9.0590 81.8235 9.0850 82.9170 ;
        RECT 8.9510 81.8235 8.9770 82.9170 ;
        RECT 8.8430 81.8235 8.8690 82.9170 ;
        RECT 8.7350 81.8235 8.7610 82.9170 ;
        RECT 8.6270 81.8235 8.6530 82.9170 ;
        RECT 8.5190 81.8235 8.5450 82.9170 ;
        RECT 8.4110 81.8235 8.4370 82.9170 ;
        RECT 8.3030 81.8235 8.3290 82.9170 ;
        RECT 8.1950 81.8235 8.2210 82.9170 ;
        RECT 8.0870 81.8235 8.1130 82.9170 ;
        RECT 7.9790 81.8235 8.0050 82.9170 ;
        RECT 7.8710 81.8235 7.8970 82.9170 ;
        RECT 7.7630 81.8235 7.7890 82.9170 ;
        RECT 7.6550 81.8235 7.6810 82.9170 ;
        RECT 7.5470 81.8235 7.5730 82.9170 ;
        RECT 7.4390 81.8235 7.4650 82.9170 ;
        RECT 7.3310 81.8235 7.3570 82.9170 ;
        RECT 7.2230 81.8235 7.2490 82.9170 ;
        RECT 7.1150 81.8235 7.1410 82.9170 ;
        RECT 7.0070 81.8235 7.0330 82.9170 ;
        RECT 6.8990 81.8235 6.9250 82.9170 ;
        RECT 6.7910 81.8235 6.8170 82.9170 ;
        RECT 6.6830 81.8235 6.7090 82.9170 ;
        RECT 6.5750 81.8235 6.6010 82.9170 ;
        RECT 6.4670 81.8235 6.4930 82.9170 ;
        RECT 6.3590 81.8235 6.3850 82.9170 ;
        RECT 6.2510 81.8235 6.2770 82.9170 ;
        RECT 6.1430 81.8235 6.1690 82.9170 ;
        RECT 6.0350 81.8235 6.0610 82.9170 ;
        RECT 5.9270 81.8235 5.9530 82.9170 ;
        RECT 5.7140 81.8235 5.7910 82.9170 ;
        RECT 3.8210 81.8235 3.8980 82.9170 ;
        RECT 3.6590 81.8235 3.6850 82.9170 ;
        RECT 3.5510 81.8235 3.5770 82.9170 ;
        RECT 3.4430 81.8235 3.4690 82.9170 ;
        RECT 3.3350 81.8235 3.3610 82.9170 ;
        RECT 3.2270 81.8235 3.2530 82.9170 ;
        RECT 3.1190 81.8235 3.1450 82.9170 ;
        RECT 3.0110 81.8235 3.0370 82.9170 ;
        RECT 2.9030 81.8235 2.9290 82.9170 ;
        RECT 2.7950 81.8235 2.8210 82.9170 ;
        RECT 2.6870 81.8235 2.7130 82.9170 ;
        RECT 2.5790 81.8235 2.6050 82.9170 ;
        RECT 2.4710 81.8235 2.4970 82.9170 ;
        RECT 2.3630 81.8235 2.3890 82.9170 ;
        RECT 2.2550 81.8235 2.2810 82.9170 ;
        RECT 2.1470 81.8235 2.1730 82.9170 ;
        RECT 2.0390 81.8235 2.0650 82.9170 ;
        RECT 1.9310 81.8235 1.9570 82.9170 ;
        RECT 1.8230 81.8235 1.8490 82.9170 ;
        RECT 1.7150 81.8235 1.7410 82.9170 ;
        RECT 1.6070 81.8235 1.6330 82.9170 ;
        RECT 1.4990 81.8235 1.5250 82.9170 ;
        RECT 1.3910 81.8235 1.4170 82.9170 ;
        RECT 1.2830 81.8235 1.3090 82.9170 ;
        RECT 1.1750 81.8235 1.2010 82.9170 ;
        RECT 1.0670 81.8235 1.0930 82.9170 ;
        RECT 0.9590 81.8235 0.9850 82.9170 ;
        RECT 0.8510 81.8235 0.8770 82.9170 ;
        RECT 0.7430 81.8235 0.7690 82.9170 ;
        RECT 0.6350 81.8235 0.6610 82.9170 ;
        RECT 0.5270 81.8235 0.5530 82.9170 ;
        RECT 0.4190 81.8235 0.4450 82.9170 ;
        RECT 0.3110 81.8235 0.3370 82.9170 ;
        RECT 0.2030 81.8235 0.2290 82.9170 ;
        RECT 0.0000 81.8235 0.0850 82.9170 ;
        RECT 5.1800 82.9035 5.3080 83.9970 ;
        RECT 5.1660 83.5690 5.3080 83.8915 ;
        RECT 5.0180 83.2960 5.0800 83.9970 ;
        RECT 5.0040 83.6055 5.0800 83.7590 ;
        RECT 5.0180 82.9035 5.0440 83.9970 ;
        RECT 5.0180 83.0245 5.0580 83.2640 ;
        RECT 5.0180 82.9035 5.0800 82.9925 ;
        RECT 4.7210 83.3540 4.9270 83.9970 ;
        RECT 4.9010 82.9035 4.9270 83.9970 ;
        RECT 4.7210 83.6310 4.9410 83.8890 ;
        RECT 4.7210 82.9035 4.8190 83.9970 ;
        RECT 4.3040 82.9035 4.3870 83.9970 ;
        RECT 4.3040 82.9920 4.4010 83.9275 ;
        RECT 9.5270 82.9035 9.6120 83.9970 ;
        RECT 9.3830 82.9035 9.4090 83.9970 ;
        RECT 9.2750 82.9035 9.3010 83.9970 ;
        RECT 9.1670 82.9035 9.1930 83.9970 ;
        RECT 9.0590 82.9035 9.0850 83.9970 ;
        RECT 8.9510 82.9035 8.9770 83.9970 ;
        RECT 8.8430 82.9035 8.8690 83.9970 ;
        RECT 8.7350 82.9035 8.7610 83.9970 ;
        RECT 8.6270 82.9035 8.6530 83.9970 ;
        RECT 8.5190 82.9035 8.5450 83.9970 ;
        RECT 8.4110 82.9035 8.4370 83.9970 ;
        RECT 8.3030 82.9035 8.3290 83.9970 ;
        RECT 8.1950 82.9035 8.2210 83.9970 ;
        RECT 8.0870 82.9035 8.1130 83.9970 ;
        RECT 7.9790 82.9035 8.0050 83.9970 ;
        RECT 7.8710 82.9035 7.8970 83.9970 ;
        RECT 7.7630 82.9035 7.7890 83.9970 ;
        RECT 7.6550 82.9035 7.6810 83.9970 ;
        RECT 7.5470 82.9035 7.5730 83.9970 ;
        RECT 7.4390 82.9035 7.4650 83.9970 ;
        RECT 7.3310 82.9035 7.3570 83.9970 ;
        RECT 7.2230 82.9035 7.2490 83.9970 ;
        RECT 7.1150 82.9035 7.1410 83.9970 ;
        RECT 7.0070 82.9035 7.0330 83.9970 ;
        RECT 6.8990 82.9035 6.9250 83.9970 ;
        RECT 6.7910 82.9035 6.8170 83.9970 ;
        RECT 6.6830 82.9035 6.7090 83.9970 ;
        RECT 6.5750 82.9035 6.6010 83.9970 ;
        RECT 6.4670 82.9035 6.4930 83.9970 ;
        RECT 6.3590 82.9035 6.3850 83.9970 ;
        RECT 6.2510 82.9035 6.2770 83.9970 ;
        RECT 6.1430 82.9035 6.1690 83.9970 ;
        RECT 6.0350 82.9035 6.0610 83.9970 ;
        RECT 5.9270 82.9035 5.9530 83.9970 ;
        RECT 5.7140 82.9035 5.7910 83.9970 ;
        RECT 3.8210 82.9035 3.8980 83.9970 ;
        RECT 3.6590 82.9035 3.6850 83.9970 ;
        RECT 3.5510 82.9035 3.5770 83.9970 ;
        RECT 3.4430 82.9035 3.4690 83.9970 ;
        RECT 3.3350 82.9035 3.3610 83.9970 ;
        RECT 3.2270 82.9035 3.2530 83.9970 ;
        RECT 3.1190 82.9035 3.1450 83.9970 ;
        RECT 3.0110 82.9035 3.0370 83.9970 ;
        RECT 2.9030 82.9035 2.9290 83.9970 ;
        RECT 2.7950 82.9035 2.8210 83.9970 ;
        RECT 2.6870 82.9035 2.7130 83.9970 ;
        RECT 2.5790 82.9035 2.6050 83.9970 ;
        RECT 2.4710 82.9035 2.4970 83.9970 ;
        RECT 2.3630 82.9035 2.3890 83.9970 ;
        RECT 2.2550 82.9035 2.2810 83.9970 ;
        RECT 2.1470 82.9035 2.1730 83.9970 ;
        RECT 2.0390 82.9035 2.0650 83.9970 ;
        RECT 1.9310 82.9035 1.9570 83.9970 ;
        RECT 1.8230 82.9035 1.8490 83.9970 ;
        RECT 1.7150 82.9035 1.7410 83.9970 ;
        RECT 1.6070 82.9035 1.6330 83.9970 ;
        RECT 1.4990 82.9035 1.5250 83.9970 ;
        RECT 1.3910 82.9035 1.4170 83.9970 ;
        RECT 1.2830 82.9035 1.3090 83.9970 ;
        RECT 1.1750 82.9035 1.2010 83.9970 ;
        RECT 1.0670 82.9035 1.0930 83.9970 ;
        RECT 0.9590 82.9035 0.9850 83.9970 ;
        RECT 0.8510 82.9035 0.8770 83.9970 ;
        RECT 0.7430 82.9035 0.7690 83.9970 ;
        RECT 0.6350 82.9035 0.6610 83.9970 ;
        RECT 0.5270 82.9035 0.5530 83.9970 ;
        RECT 0.4190 82.9035 0.4450 83.9970 ;
        RECT 0.3110 82.9035 0.3370 83.9970 ;
        RECT 0.2030 82.9035 0.2290 83.9970 ;
        RECT 0.0000 82.9035 0.0850 83.9970 ;
        RECT 5.1800 83.9835 5.3080 85.0770 ;
        RECT 5.1660 84.6490 5.3080 84.9715 ;
        RECT 5.0180 84.3760 5.0800 85.0770 ;
        RECT 5.0040 84.6855 5.0800 84.8390 ;
        RECT 5.0180 83.9835 5.0440 85.0770 ;
        RECT 5.0180 84.1045 5.0580 84.3440 ;
        RECT 5.0180 83.9835 5.0800 84.0725 ;
        RECT 4.7210 84.4340 4.9270 85.0770 ;
        RECT 4.9010 83.9835 4.9270 85.0770 ;
        RECT 4.7210 84.7110 4.9410 84.9690 ;
        RECT 4.7210 83.9835 4.8190 85.0770 ;
        RECT 4.3040 83.9835 4.3870 85.0770 ;
        RECT 4.3040 84.0720 4.4010 85.0075 ;
        RECT 9.5270 83.9835 9.6120 85.0770 ;
        RECT 9.3830 83.9835 9.4090 85.0770 ;
        RECT 9.2750 83.9835 9.3010 85.0770 ;
        RECT 9.1670 83.9835 9.1930 85.0770 ;
        RECT 9.0590 83.9835 9.0850 85.0770 ;
        RECT 8.9510 83.9835 8.9770 85.0770 ;
        RECT 8.8430 83.9835 8.8690 85.0770 ;
        RECT 8.7350 83.9835 8.7610 85.0770 ;
        RECT 8.6270 83.9835 8.6530 85.0770 ;
        RECT 8.5190 83.9835 8.5450 85.0770 ;
        RECT 8.4110 83.9835 8.4370 85.0770 ;
        RECT 8.3030 83.9835 8.3290 85.0770 ;
        RECT 8.1950 83.9835 8.2210 85.0770 ;
        RECT 8.0870 83.9835 8.1130 85.0770 ;
        RECT 7.9790 83.9835 8.0050 85.0770 ;
        RECT 7.8710 83.9835 7.8970 85.0770 ;
        RECT 7.7630 83.9835 7.7890 85.0770 ;
        RECT 7.6550 83.9835 7.6810 85.0770 ;
        RECT 7.5470 83.9835 7.5730 85.0770 ;
        RECT 7.4390 83.9835 7.4650 85.0770 ;
        RECT 7.3310 83.9835 7.3570 85.0770 ;
        RECT 7.2230 83.9835 7.2490 85.0770 ;
        RECT 7.1150 83.9835 7.1410 85.0770 ;
        RECT 7.0070 83.9835 7.0330 85.0770 ;
        RECT 6.8990 83.9835 6.9250 85.0770 ;
        RECT 6.7910 83.9835 6.8170 85.0770 ;
        RECT 6.6830 83.9835 6.7090 85.0770 ;
        RECT 6.5750 83.9835 6.6010 85.0770 ;
        RECT 6.4670 83.9835 6.4930 85.0770 ;
        RECT 6.3590 83.9835 6.3850 85.0770 ;
        RECT 6.2510 83.9835 6.2770 85.0770 ;
        RECT 6.1430 83.9835 6.1690 85.0770 ;
        RECT 6.0350 83.9835 6.0610 85.0770 ;
        RECT 5.9270 83.9835 5.9530 85.0770 ;
        RECT 5.7140 83.9835 5.7910 85.0770 ;
        RECT 3.8210 83.9835 3.8980 85.0770 ;
        RECT 3.6590 83.9835 3.6850 85.0770 ;
        RECT 3.5510 83.9835 3.5770 85.0770 ;
        RECT 3.4430 83.9835 3.4690 85.0770 ;
        RECT 3.3350 83.9835 3.3610 85.0770 ;
        RECT 3.2270 83.9835 3.2530 85.0770 ;
        RECT 3.1190 83.9835 3.1450 85.0770 ;
        RECT 3.0110 83.9835 3.0370 85.0770 ;
        RECT 2.9030 83.9835 2.9290 85.0770 ;
        RECT 2.7950 83.9835 2.8210 85.0770 ;
        RECT 2.6870 83.9835 2.7130 85.0770 ;
        RECT 2.5790 83.9835 2.6050 85.0770 ;
        RECT 2.4710 83.9835 2.4970 85.0770 ;
        RECT 2.3630 83.9835 2.3890 85.0770 ;
        RECT 2.2550 83.9835 2.2810 85.0770 ;
        RECT 2.1470 83.9835 2.1730 85.0770 ;
        RECT 2.0390 83.9835 2.0650 85.0770 ;
        RECT 1.9310 83.9835 1.9570 85.0770 ;
        RECT 1.8230 83.9835 1.8490 85.0770 ;
        RECT 1.7150 83.9835 1.7410 85.0770 ;
        RECT 1.6070 83.9835 1.6330 85.0770 ;
        RECT 1.4990 83.9835 1.5250 85.0770 ;
        RECT 1.3910 83.9835 1.4170 85.0770 ;
        RECT 1.2830 83.9835 1.3090 85.0770 ;
        RECT 1.1750 83.9835 1.2010 85.0770 ;
        RECT 1.0670 83.9835 1.0930 85.0770 ;
        RECT 0.9590 83.9835 0.9850 85.0770 ;
        RECT 0.8510 83.9835 0.8770 85.0770 ;
        RECT 0.7430 83.9835 0.7690 85.0770 ;
        RECT 0.6350 83.9835 0.6610 85.0770 ;
        RECT 0.5270 83.9835 0.5530 85.0770 ;
        RECT 0.4190 83.9835 0.4450 85.0770 ;
        RECT 0.3110 83.9835 0.3370 85.0770 ;
        RECT 0.2030 83.9835 0.2290 85.0770 ;
        RECT 0.0000 83.9835 0.0850 85.0770 ;
        RECT 5.1800 85.0635 5.3080 86.1570 ;
        RECT 5.1660 85.7290 5.3080 86.0515 ;
        RECT 5.0180 85.4560 5.0800 86.1570 ;
        RECT 5.0040 85.7655 5.0800 85.9190 ;
        RECT 5.0180 85.0635 5.0440 86.1570 ;
        RECT 5.0180 85.1845 5.0580 85.4240 ;
        RECT 5.0180 85.0635 5.0800 85.1525 ;
        RECT 4.7210 85.5140 4.9270 86.1570 ;
        RECT 4.9010 85.0635 4.9270 86.1570 ;
        RECT 4.7210 85.7910 4.9410 86.0490 ;
        RECT 4.7210 85.0635 4.8190 86.1570 ;
        RECT 4.3040 85.0635 4.3870 86.1570 ;
        RECT 4.3040 85.1520 4.4010 86.0875 ;
        RECT 9.5270 85.0635 9.6120 86.1570 ;
        RECT 9.3830 85.0635 9.4090 86.1570 ;
        RECT 9.2750 85.0635 9.3010 86.1570 ;
        RECT 9.1670 85.0635 9.1930 86.1570 ;
        RECT 9.0590 85.0635 9.0850 86.1570 ;
        RECT 8.9510 85.0635 8.9770 86.1570 ;
        RECT 8.8430 85.0635 8.8690 86.1570 ;
        RECT 8.7350 85.0635 8.7610 86.1570 ;
        RECT 8.6270 85.0635 8.6530 86.1570 ;
        RECT 8.5190 85.0635 8.5450 86.1570 ;
        RECT 8.4110 85.0635 8.4370 86.1570 ;
        RECT 8.3030 85.0635 8.3290 86.1570 ;
        RECT 8.1950 85.0635 8.2210 86.1570 ;
        RECT 8.0870 85.0635 8.1130 86.1570 ;
        RECT 7.9790 85.0635 8.0050 86.1570 ;
        RECT 7.8710 85.0635 7.8970 86.1570 ;
        RECT 7.7630 85.0635 7.7890 86.1570 ;
        RECT 7.6550 85.0635 7.6810 86.1570 ;
        RECT 7.5470 85.0635 7.5730 86.1570 ;
        RECT 7.4390 85.0635 7.4650 86.1570 ;
        RECT 7.3310 85.0635 7.3570 86.1570 ;
        RECT 7.2230 85.0635 7.2490 86.1570 ;
        RECT 7.1150 85.0635 7.1410 86.1570 ;
        RECT 7.0070 85.0635 7.0330 86.1570 ;
        RECT 6.8990 85.0635 6.9250 86.1570 ;
        RECT 6.7910 85.0635 6.8170 86.1570 ;
        RECT 6.6830 85.0635 6.7090 86.1570 ;
        RECT 6.5750 85.0635 6.6010 86.1570 ;
        RECT 6.4670 85.0635 6.4930 86.1570 ;
        RECT 6.3590 85.0635 6.3850 86.1570 ;
        RECT 6.2510 85.0635 6.2770 86.1570 ;
        RECT 6.1430 85.0635 6.1690 86.1570 ;
        RECT 6.0350 85.0635 6.0610 86.1570 ;
        RECT 5.9270 85.0635 5.9530 86.1570 ;
        RECT 5.7140 85.0635 5.7910 86.1570 ;
        RECT 3.8210 85.0635 3.8980 86.1570 ;
        RECT 3.6590 85.0635 3.6850 86.1570 ;
        RECT 3.5510 85.0635 3.5770 86.1570 ;
        RECT 3.4430 85.0635 3.4690 86.1570 ;
        RECT 3.3350 85.0635 3.3610 86.1570 ;
        RECT 3.2270 85.0635 3.2530 86.1570 ;
        RECT 3.1190 85.0635 3.1450 86.1570 ;
        RECT 3.0110 85.0635 3.0370 86.1570 ;
        RECT 2.9030 85.0635 2.9290 86.1570 ;
        RECT 2.7950 85.0635 2.8210 86.1570 ;
        RECT 2.6870 85.0635 2.7130 86.1570 ;
        RECT 2.5790 85.0635 2.6050 86.1570 ;
        RECT 2.4710 85.0635 2.4970 86.1570 ;
        RECT 2.3630 85.0635 2.3890 86.1570 ;
        RECT 2.2550 85.0635 2.2810 86.1570 ;
        RECT 2.1470 85.0635 2.1730 86.1570 ;
        RECT 2.0390 85.0635 2.0650 86.1570 ;
        RECT 1.9310 85.0635 1.9570 86.1570 ;
        RECT 1.8230 85.0635 1.8490 86.1570 ;
        RECT 1.7150 85.0635 1.7410 86.1570 ;
        RECT 1.6070 85.0635 1.6330 86.1570 ;
        RECT 1.4990 85.0635 1.5250 86.1570 ;
        RECT 1.3910 85.0635 1.4170 86.1570 ;
        RECT 1.2830 85.0635 1.3090 86.1570 ;
        RECT 1.1750 85.0635 1.2010 86.1570 ;
        RECT 1.0670 85.0635 1.0930 86.1570 ;
        RECT 0.9590 85.0635 0.9850 86.1570 ;
        RECT 0.8510 85.0635 0.8770 86.1570 ;
        RECT 0.7430 85.0635 0.7690 86.1570 ;
        RECT 0.6350 85.0635 0.6610 86.1570 ;
        RECT 0.5270 85.0635 0.5530 86.1570 ;
        RECT 0.4190 85.0635 0.4450 86.1570 ;
        RECT 0.3110 85.0635 0.3370 86.1570 ;
        RECT 0.2030 85.0635 0.2290 86.1570 ;
        RECT 0.0000 85.0635 0.0850 86.1570 ;
        RECT 5.1800 86.1435 5.3080 87.2370 ;
        RECT 5.1660 86.8090 5.3080 87.1315 ;
        RECT 5.0180 86.5360 5.0800 87.2370 ;
        RECT 5.0040 86.8455 5.0800 86.9990 ;
        RECT 5.0180 86.1435 5.0440 87.2370 ;
        RECT 5.0180 86.2645 5.0580 86.5040 ;
        RECT 5.0180 86.1435 5.0800 86.2325 ;
        RECT 4.7210 86.5940 4.9270 87.2370 ;
        RECT 4.9010 86.1435 4.9270 87.2370 ;
        RECT 4.7210 86.8710 4.9410 87.1290 ;
        RECT 4.7210 86.1435 4.8190 87.2370 ;
        RECT 4.3040 86.1435 4.3870 87.2370 ;
        RECT 4.3040 86.2320 4.4010 87.1675 ;
        RECT 9.5270 86.1435 9.6120 87.2370 ;
        RECT 9.3830 86.1435 9.4090 87.2370 ;
        RECT 9.2750 86.1435 9.3010 87.2370 ;
        RECT 9.1670 86.1435 9.1930 87.2370 ;
        RECT 9.0590 86.1435 9.0850 87.2370 ;
        RECT 8.9510 86.1435 8.9770 87.2370 ;
        RECT 8.8430 86.1435 8.8690 87.2370 ;
        RECT 8.7350 86.1435 8.7610 87.2370 ;
        RECT 8.6270 86.1435 8.6530 87.2370 ;
        RECT 8.5190 86.1435 8.5450 87.2370 ;
        RECT 8.4110 86.1435 8.4370 87.2370 ;
        RECT 8.3030 86.1435 8.3290 87.2370 ;
        RECT 8.1950 86.1435 8.2210 87.2370 ;
        RECT 8.0870 86.1435 8.1130 87.2370 ;
        RECT 7.9790 86.1435 8.0050 87.2370 ;
        RECT 7.8710 86.1435 7.8970 87.2370 ;
        RECT 7.7630 86.1435 7.7890 87.2370 ;
        RECT 7.6550 86.1435 7.6810 87.2370 ;
        RECT 7.5470 86.1435 7.5730 87.2370 ;
        RECT 7.4390 86.1435 7.4650 87.2370 ;
        RECT 7.3310 86.1435 7.3570 87.2370 ;
        RECT 7.2230 86.1435 7.2490 87.2370 ;
        RECT 7.1150 86.1435 7.1410 87.2370 ;
        RECT 7.0070 86.1435 7.0330 87.2370 ;
        RECT 6.8990 86.1435 6.9250 87.2370 ;
        RECT 6.7910 86.1435 6.8170 87.2370 ;
        RECT 6.6830 86.1435 6.7090 87.2370 ;
        RECT 6.5750 86.1435 6.6010 87.2370 ;
        RECT 6.4670 86.1435 6.4930 87.2370 ;
        RECT 6.3590 86.1435 6.3850 87.2370 ;
        RECT 6.2510 86.1435 6.2770 87.2370 ;
        RECT 6.1430 86.1435 6.1690 87.2370 ;
        RECT 6.0350 86.1435 6.0610 87.2370 ;
        RECT 5.9270 86.1435 5.9530 87.2370 ;
        RECT 5.7140 86.1435 5.7910 87.2370 ;
        RECT 3.8210 86.1435 3.8980 87.2370 ;
        RECT 3.6590 86.1435 3.6850 87.2370 ;
        RECT 3.5510 86.1435 3.5770 87.2370 ;
        RECT 3.4430 86.1435 3.4690 87.2370 ;
        RECT 3.3350 86.1435 3.3610 87.2370 ;
        RECT 3.2270 86.1435 3.2530 87.2370 ;
        RECT 3.1190 86.1435 3.1450 87.2370 ;
        RECT 3.0110 86.1435 3.0370 87.2370 ;
        RECT 2.9030 86.1435 2.9290 87.2370 ;
        RECT 2.7950 86.1435 2.8210 87.2370 ;
        RECT 2.6870 86.1435 2.7130 87.2370 ;
        RECT 2.5790 86.1435 2.6050 87.2370 ;
        RECT 2.4710 86.1435 2.4970 87.2370 ;
        RECT 2.3630 86.1435 2.3890 87.2370 ;
        RECT 2.2550 86.1435 2.2810 87.2370 ;
        RECT 2.1470 86.1435 2.1730 87.2370 ;
        RECT 2.0390 86.1435 2.0650 87.2370 ;
        RECT 1.9310 86.1435 1.9570 87.2370 ;
        RECT 1.8230 86.1435 1.8490 87.2370 ;
        RECT 1.7150 86.1435 1.7410 87.2370 ;
        RECT 1.6070 86.1435 1.6330 87.2370 ;
        RECT 1.4990 86.1435 1.5250 87.2370 ;
        RECT 1.3910 86.1435 1.4170 87.2370 ;
        RECT 1.2830 86.1435 1.3090 87.2370 ;
        RECT 1.1750 86.1435 1.2010 87.2370 ;
        RECT 1.0670 86.1435 1.0930 87.2370 ;
        RECT 0.9590 86.1435 0.9850 87.2370 ;
        RECT 0.8510 86.1435 0.8770 87.2370 ;
        RECT 0.7430 86.1435 0.7690 87.2370 ;
        RECT 0.6350 86.1435 0.6610 87.2370 ;
        RECT 0.5270 86.1435 0.5530 87.2370 ;
        RECT 0.4190 86.1435 0.4450 87.2370 ;
        RECT 0.3110 86.1435 0.3370 87.2370 ;
        RECT 0.2030 86.1435 0.2290 87.2370 ;
        RECT 0.0000 86.1435 0.0850 87.2370 ;
        RECT 5.1800 87.2235 5.3080 88.3170 ;
        RECT 5.1660 87.8890 5.3080 88.2115 ;
        RECT 5.0180 87.6160 5.0800 88.3170 ;
        RECT 5.0040 87.9255 5.0800 88.0790 ;
        RECT 5.0180 87.2235 5.0440 88.3170 ;
        RECT 5.0180 87.3445 5.0580 87.5840 ;
        RECT 5.0180 87.2235 5.0800 87.3125 ;
        RECT 4.7210 87.6740 4.9270 88.3170 ;
        RECT 4.9010 87.2235 4.9270 88.3170 ;
        RECT 4.7210 87.9510 4.9410 88.2090 ;
        RECT 4.7210 87.2235 4.8190 88.3170 ;
        RECT 4.3040 87.2235 4.3870 88.3170 ;
        RECT 4.3040 87.3120 4.4010 88.2475 ;
        RECT 9.5270 87.2235 9.6120 88.3170 ;
        RECT 9.3830 87.2235 9.4090 88.3170 ;
        RECT 9.2750 87.2235 9.3010 88.3170 ;
        RECT 9.1670 87.2235 9.1930 88.3170 ;
        RECT 9.0590 87.2235 9.0850 88.3170 ;
        RECT 8.9510 87.2235 8.9770 88.3170 ;
        RECT 8.8430 87.2235 8.8690 88.3170 ;
        RECT 8.7350 87.2235 8.7610 88.3170 ;
        RECT 8.6270 87.2235 8.6530 88.3170 ;
        RECT 8.5190 87.2235 8.5450 88.3170 ;
        RECT 8.4110 87.2235 8.4370 88.3170 ;
        RECT 8.3030 87.2235 8.3290 88.3170 ;
        RECT 8.1950 87.2235 8.2210 88.3170 ;
        RECT 8.0870 87.2235 8.1130 88.3170 ;
        RECT 7.9790 87.2235 8.0050 88.3170 ;
        RECT 7.8710 87.2235 7.8970 88.3170 ;
        RECT 7.7630 87.2235 7.7890 88.3170 ;
        RECT 7.6550 87.2235 7.6810 88.3170 ;
        RECT 7.5470 87.2235 7.5730 88.3170 ;
        RECT 7.4390 87.2235 7.4650 88.3170 ;
        RECT 7.3310 87.2235 7.3570 88.3170 ;
        RECT 7.2230 87.2235 7.2490 88.3170 ;
        RECT 7.1150 87.2235 7.1410 88.3170 ;
        RECT 7.0070 87.2235 7.0330 88.3170 ;
        RECT 6.8990 87.2235 6.9250 88.3170 ;
        RECT 6.7910 87.2235 6.8170 88.3170 ;
        RECT 6.6830 87.2235 6.7090 88.3170 ;
        RECT 6.5750 87.2235 6.6010 88.3170 ;
        RECT 6.4670 87.2235 6.4930 88.3170 ;
        RECT 6.3590 87.2235 6.3850 88.3170 ;
        RECT 6.2510 87.2235 6.2770 88.3170 ;
        RECT 6.1430 87.2235 6.1690 88.3170 ;
        RECT 6.0350 87.2235 6.0610 88.3170 ;
        RECT 5.9270 87.2235 5.9530 88.3170 ;
        RECT 5.7140 87.2235 5.7910 88.3170 ;
        RECT 3.8210 87.2235 3.8980 88.3170 ;
        RECT 3.6590 87.2235 3.6850 88.3170 ;
        RECT 3.5510 87.2235 3.5770 88.3170 ;
        RECT 3.4430 87.2235 3.4690 88.3170 ;
        RECT 3.3350 87.2235 3.3610 88.3170 ;
        RECT 3.2270 87.2235 3.2530 88.3170 ;
        RECT 3.1190 87.2235 3.1450 88.3170 ;
        RECT 3.0110 87.2235 3.0370 88.3170 ;
        RECT 2.9030 87.2235 2.9290 88.3170 ;
        RECT 2.7950 87.2235 2.8210 88.3170 ;
        RECT 2.6870 87.2235 2.7130 88.3170 ;
        RECT 2.5790 87.2235 2.6050 88.3170 ;
        RECT 2.4710 87.2235 2.4970 88.3170 ;
        RECT 2.3630 87.2235 2.3890 88.3170 ;
        RECT 2.2550 87.2235 2.2810 88.3170 ;
        RECT 2.1470 87.2235 2.1730 88.3170 ;
        RECT 2.0390 87.2235 2.0650 88.3170 ;
        RECT 1.9310 87.2235 1.9570 88.3170 ;
        RECT 1.8230 87.2235 1.8490 88.3170 ;
        RECT 1.7150 87.2235 1.7410 88.3170 ;
        RECT 1.6070 87.2235 1.6330 88.3170 ;
        RECT 1.4990 87.2235 1.5250 88.3170 ;
        RECT 1.3910 87.2235 1.4170 88.3170 ;
        RECT 1.2830 87.2235 1.3090 88.3170 ;
        RECT 1.1750 87.2235 1.2010 88.3170 ;
        RECT 1.0670 87.2235 1.0930 88.3170 ;
        RECT 0.9590 87.2235 0.9850 88.3170 ;
        RECT 0.8510 87.2235 0.8770 88.3170 ;
        RECT 0.7430 87.2235 0.7690 88.3170 ;
        RECT 0.6350 87.2235 0.6610 88.3170 ;
        RECT 0.5270 87.2235 0.5530 88.3170 ;
        RECT 0.4190 87.2235 0.4450 88.3170 ;
        RECT 0.3110 87.2235 0.3370 88.3170 ;
        RECT 0.2030 87.2235 0.2290 88.3170 ;
        RECT 0.0000 87.2235 0.0850 88.3170 ;
        RECT 5.1800 88.3035 5.3080 89.3970 ;
        RECT 5.1660 88.9690 5.3080 89.2915 ;
        RECT 5.0180 88.6960 5.0800 89.3970 ;
        RECT 5.0040 89.0055 5.0800 89.1590 ;
        RECT 5.0180 88.3035 5.0440 89.3970 ;
        RECT 5.0180 88.4245 5.0580 88.6640 ;
        RECT 5.0180 88.3035 5.0800 88.3925 ;
        RECT 4.7210 88.7540 4.9270 89.3970 ;
        RECT 4.9010 88.3035 4.9270 89.3970 ;
        RECT 4.7210 89.0310 4.9410 89.2890 ;
        RECT 4.7210 88.3035 4.8190 89.3970 ;
        RECT 4.3040 88.3035 4.3870 89.3970 ;
        RECT 4.3040 88.3920 4.4010 89.3275 ;
        RECT 9.5270 88.3035 9.6120 89.3970 ;
        RECT 9.3830 88.3035 9.4090 89.3970 ;
        RECT 9.2750 88.3035 9.3010 89.3970 ;
        RECT 9.1670 88.3035 9.1930 89.3970 ;
        RECT 9.0590 88.3035 9.0850 89.3970 ;
        RECT 8.9510 88.3035 8.9770 89.3970 ;
        RECT 8.8430 88.3035 8.8690 89.3970 ;
        RECT 8.7350 88.3035 8.7610 89.3970 ;
        RECT 8.6270 88.3035 8.6530 89.3970 ;
        RECT 8.5190 88.3035 8.5450 89.3970 ;
        RECT 8.4110 88.3035 8.4370 89.3970 ;
        RECT 8.3030 88.3035 8.3290 89.3970 ;
        RECT 8.1950 88.3035 8.2210 89.3970 ;
        RECT 8.0870 88.3035 8.1130 89.3970 ;
        RECT 7.9790 88.3035 8.0050 89.3970 ;
        RECT 7.8710 88.3035 7.8970 89.3970 ;
        RECT 7.7630 88.3035 7.7890 89.3970 ;
        RECT 7.6550 88.3035 7.6810 89.3970 ;
        RECT 7.5470 88.3035 7.5730 89.3970 ;
        RECT 7.4390 88.3035 7.4650 89.3970 ;
        RECT 7.3310 88.3035 7.3570 89.3970 ;
        RECT 7.2230 88.3035 7.2490 89.3970 ;
        RECT 7.1150 88.3035 7.1410 89.3970 ;
        RECT 7.0070 88.3035 7.0330 89.3970 ;
        RECT 6.8990 88.3035 6.9250 89.3970 ;
        RECT 6.7910 88.3035 6.8170 89.3970 ;
        RECT 6.6830 88.3035 6.7090 89.3970 ;
        RECT 6.5750 88.3035 6.6010 89.3970 ;
        RECT 6.4670 88.3035 6.4930 89.3970 ;
        RECT 6.3590 88.3035 6.3850 89.3970 ;
        RECT 6.2510 88.3035 6.2770 89.3970 ;
        RECT 6.1430 88.3035 6.1690 89.3970 ;
        RECT 6.0350 88.3035 6.0610 89.3970 ;
        RECT 5.9270 88.3035 5.9530 89.3970 ;
        RECT 5.7140 88.3035 5.7910 89.3970 ;
        RECT 3.8210 88.3035 3.8980 89.3970 ;
        RECT 3.6590 88.3035 3.6850 89.3970 ;
        RECT 3.5510 88.3035 3.5770 89.3970 ;
        RECT 3.4430 88.3035 3.4690 89.3970 ;
        RECT 3.3350 88.3035 3.3610 89.3970 ;
        RECT 3.2270 88.3035 3.2530 89.3970 ;
        RECT 3.1190 88.3035 3.1450 89.3970 ;
        RECT 3.0110 88.3035 3.0370 89.3970 ;
        RECT 2.9030 88.3035 2.9290 89.3970 ;
        RECT 2.7950 88.3035 2.8210 89.3970 ;
        RECT 2.6870 88.3035 2.7130 89.3970 ;
        RECT 2.5790 88.3035 2.6050 89.3970 ;
        RECT 2.4710 88.3035 2.4970 89.3970 ;
        RECT 2.3630 88.3035 2.3890 89.3970 ;
        RECT 2.2550 88.3035 2.2810 89.3970 ;
        RECT 2.1470 88.3035 2.1730 89.3970 ;
        RECT 2.0390 88.3035 2.0650 89.3970 ;
        RECT 1.9310 88.3035 1.9570 89.3970 ;
        RECT 1.8230 88.3035 1.8490 89.3970 ;
        RECT 1.7150 88.3035 1.7410 89.3970 ;
        RECT 1.6070 88.3035 1.6330 89.3970 ;
        RECT 1.4990 88.3035 1.5250 89.3970 ;
        RECT 1.3910 88.3035 1.4170 89.3970 ;
        RECT 1.2830 88.3035 1.3090 89.3970 ;
        RECT 1.1750 88.3035 1.2010 89.3970 ;
        RECT 1.0670 88.3035 1.0930 89.3970 ;
        RECT 0.9590 88.3035 0.9850 89.3970 ;
        RECT 0.8510 88.3035 0.8770 89.3970 ;
        RECT 0.7430 88.3035 0.7690 89.3970 ;
        RECT 0.6350 88.3035 0.6610 89.3970 ;
        RECT 0.5270 88.3035 0.5530 89.3970 ;
        RECT 0.4190 88.3035 0.4450 89.3970 ;
        RECT 0.3110 88.3035 0.3370 89.3970 ;
        RECT 0.2030 88.3035 0.2290 89.3970 ;
        RECT 0.0000 88.3035 0.0850 89.3970 ;
        RECT 5.1800 89.3835 5.3080 90.4770 ;
        RECT 5.1660 90.0490 5.3080 90.3715 ;
        RECT 5.0180 89.7760 5.0800 90.4770 ;
        RECT 5.0040 90.0855 5.0800 90.2390 ;
        RECT 5.0180 89.3835 5.0440 90.4770 ;
        RECT 5.0180 89.5045 5.0580 89.7440 ;
        RECT 5.0180 89.3835 5.0800 89.4725 ;
        RECT 4.7210 89.8340 4.9270 90.4770 ;
        RECT 4.9010 89.3835 4.9270 90.4770 ;
        RECT 4.7210 90.1110 4.9410 90.3690 ;
        RECT 4.7210 89.3835 4.8190 90.4770 ;
        RECT 4.3040 89.3835 4.3870 90.4770 ;
        RECT 4.3040 89.4720 4.4010 90.4075 ;
        RECT 9.5270 89.3835 9.6120 90.4770 ;
        RECT 9.3830 89.3835 9.4090 90.4770 ;
        RECT 9.2750 89.3835 9.3010 90.4770 ;
        RECT 9.1670 89.3835 9.1930 90.4770 ;
        RECT 9.0590 89.3835 9.0850 90.4770 ;
        RECT 8.9510 89.3835 8.9770 90.4770 ;
        RECT 8.8430 89.3835 8.8690 90.4770 ;
        RECT 8.7350 89.3835 8.7610 90.4770 ;
        RECT 8.6270 89.3835 8.6530 90.4770 ;
        RECT 8.5190 89.3835 8.5450 90.4770 ;
        RECT 8.4110 89.3835 8.4370 90.4770 ;
        RECT 8.3030 89.3835 8.3290 90.4770 ;
        RECT 8.1950 89.3835 8.2210 90.4770 ;
        RECT 8.0870 89.3835 8.1130 90.4770 ;
        RECT 7.9790 89.3835 8.0050 90.4770 ;
        RECT 7.8710 89.3835 7.8970 90.4770 ;
        RECT 7.7630 89.3835 7.7890 90.4770 ;
        RECT 7.6550 89.3835 7.6810 90.4770 ;
        RECT 7.5470 89.3835 7.5730 90.4770 ;
        RECT 7.4390 89.3835 7.4650 90.4770 ;
        RECT 7.3310 89.3835 7.3570 90.4770 ;
        RECT 7.2230 89.3835 7.2490 90.4770 ;
        RECT 7.1150 89.3835 7.1410 90.4770 ;
        RECT 7.0070 89.3835 7.0330 90.4770 ;
        RECT 6.8990 89.3835 6.9250 90.4770 ;
        RECT 6.7910 89.3835 6.8170 90.4770 ;
        RECT 6.6830 89.3835 6.7090 90.4770 ;
        RECT 6.5750 89.3835 6.6010 90.4770 ;
        RECT 6.4670 89.3835 6.4930 90.4770 ;
        RECT 6.3590 89.3835 6.3850 90.4770 ;
        RECT 6.2510 89.3835 6.2770 90.4770 ;
        RECT 6.1430 89.3835 6.1690 90.4770 ;
        RECT 6.0350 89.3835 6.0610 90.4770 ;
        RECT 5.9270 89.3835 5.9530 90.4770 ;
        RECT 5.7140 89.3835 5.7910 90.4770 ;
        RECT 3.8210 89.3835 3.8980 90.4770 ;
        RECT 3.6590 89.3835 3.6850 90.4770 ;
        RECT 3.5510 89.3835 3.5770 90.4770 ;
        RECT 3.4430 89.3835 3.4690 90.4770 ;
        RECT 3.3350 89.3835 3.3610 90.4770 ;
        RECT 3.2270 89.3835 3.2530 90.4770 ;
        RECT 3.1190 89.3835 3.1450 90.4770 ;
        RECT 3.0110 89.3835 3.0370 90.4770 ;
        RECT 2.9030 89.3835 2.9290 90.4770 ;
        RECT 2.7950 89.3835 2.8210 90.4770 ;
        RECT 2.6870 89.3835 2.7130 90.4770 ;
        RECT 2.5790 89.3835 2.6050 90.4770 ;
        RECT 2.4710 89.3835 2.4970 90.4770 ;
        RECT 2.3630 89.3835 2.3890 90.4770 ;
        RECT 2.2550 89.3835 2.2810 90.4770 ;
        RECT 2.1470 89.3835 2.1730 90.4770 ;
        RECT 2.0390 89.3835 2.0650 90.4770 ;
        RECT 1.9310 89.3835 1.9570 90.4770 ;
        RECT 1.8230 89.3835 1.8490 90.4770 ;
        RECT 1.7150 89.3835 1.7410 90.4770 ;
        RECT 1.6070 89.3835 1.6330 90.4770 ;
        RECT 1.4990 89.3835 1.5250 90.4770 ;
        RECT 1.3910 89.3835 1.4170 90.4770 ;
        RECT 1.2830 89.3835 1.3090 90.4770 ;
        RECT 1.1750 89.3835 1.2010 90.4770 ;
        RECT 1.0670 89.3835 1.0930 90.4770 ;
        RECT 0.9590 89.3835 0.9850 90.4770 ;
        RECT 0.8510 89.3835 0.8770 90.4770 ;
        RECT 0.7430 89.3835 0.7690 90.4770 ;
        RECT 0.6350 89.3835 0.6610 90.4770 ;
        RECT 0.5270 89.3835 0.5530 90.4770 ;
        RECT 0.4190 89.3835 0.4450 90.4770 ;
        RECT 0.3110 89.3835 0.3370 90.4770 ;
        RECT 0.2030 89.3835 0.2290 90.4770 ;
        RECT 0.0000 89.3835 0.0850 90.4770 ;
        RECT 5.1800 90.4635 5.3080 91.5570 ;
        RECT 5.1660 91.1290 5.3080 91.4515 ;
        RECT 5.0180 90.8560 5.0800 91.5570 ;
        RECT 5.0040 91.1655 5.0800 91.3190 ;
        RECT 5.0180 90.4635 5.0440 91.5570 ;
        RECT 5.0180 90.5845 5.0580 90.8240 ;
        RECT 5.0180 90.4635 5.0800 90.5525 ;
        RECT 4.7210 90.9140 4.9270 91.5570 ;
        RECT 4.9010 90.4635 4.9270 91.5570 ;
        RECT 4.7210 91.1910 4.9410 91.4490 ;
        RECT 4.7210 90.4635 4.8190 91.5570 ;
        RECT 4.3040 90.4635 4.3870 91.5570 ;
        RECT 4.3040 90.5520 4.4010 91.4875 ;
        RECT 9.5270 90.4635 9.6120 91.5570 ;
        RECT 9.3830 90.4635 9.4090 91.5570 ;
        RECT 9.2750 90.4635 9.3010 91.5570 ;
        RECT 9.1670 90.4635 9.1930 91.5570 ;
        RECT 9.0590 90.4635 9.0850 91.5570 ;
        RECT 8.9510 90.4635 8.9770 91.5570 ;
        RECT 8.8430 90.4635 8.8690 91.5570 ;
        RECT 8.7350 90.4635 8.7610 91.5570 ;
        RECT 8.6270 90.4635 8.6530 91.5570 ;
        RECT 8.5190 90.4635 8.5450 91.5570 ;
        RECT 8.4110 90.4635 8.4370 91.5570 ;
        RECT 8.3030 90.4635 8.3290 91.5570 ;
        RECT 8.1950 90.4635 8.2210 91.5570 ;
        RECT 8.0870 90.4635 8.1130 91.5570 ;
        RECT 7.9790 90.4635 8.0050 91.5570 ;
        RECT 7.8710 90.4635 7.8970 91.5570 ;
        RECT 7.7630 90.4635 7.7890 91.5570 ;
        RECT 7.6550 90.4635 7.6810 91.5570 ;
        RECT 7.5470 90.4635 7.5730 91.5570 ;
        RECT 7.4390 90.4635 7.4650 91.5570 ;
        RECT 7.3310 90.4635 7.3570 91.5570 ;
        RECT 7.2230 90.4635 7.2490 91.5570 ;
        RECT 7.1150 90.4635 7.1410 91.5570 ;
        RECT 7.0070 90.4635 7.0330 91.5570 ;
        RECT 6.8990 90.4635 6.9250 91.5570 ;
        RECT 6.7910 90.4635 6.8170 91.5570 ;
        RECT 6.6830 90.4635 6.7090 91.5570 ;
        RECT 6.5750 90.4635 6.6010 91.5570 ;
        RECT 6.4670 90.4635 6.4930 91.5570 ;
        RECT 6.3590 90.4635 6.3850 91.5570 ;
        RECT 6.2510 90.4635 6.2770 91.5570 ;
        RECT 6.1430 90.4635 6.1690 91.5570 ;
        RECT 6.0350 90.4635 6.0610 91.5570 ;
        RECT 5.9270 90.4635 5.9530 91.5570 ;
        RECT 5.7140 90.4635 5.7910 91.5570 ;
        RECT 3.8210 90.4635 3.8980 91.5570 ;
        RECT 3.6590 90.4635 3.6850 91.5570 ;
        RECT 3.5510 90.4635 3.5770 91.5570 ;
        RECT 3.4430 90.4635 3.4690 91.5570 ;
        RECT 3.3350 90.4635 3.3610 91.5570 ;
        RECT 3.2270 90.4635 3.2530 91.5570 ;
        RECT 3.1190 90.4635 3.1450 91.5570 ;
        RECT 3.0110 90.4635 3.0370 91.5570 ;
        RECT 2.9030 90.4635 2.9290 91.5570 ;
        RECT 2.7950 90.4635 2.8210 91.5570 ;
        RECT 2.6870 90.4635 2.7130 91.5570 ;
        RECT 2.5790 90.4635 2.6050 91.5570 ;
        RECT 2.4710 90.4635 2.4970 91.5570 ;
        RECT 2.3630 90.4635 2.3890 91.5570 ;
        RECT 2.2550 90.4635 2.2810 91.5570 ;
        RECT 2.1470 90.4635 2.1730 91.5570 ;
        RECT 2.0390 90.4635 2.0650 91.5570 ;
        RECT 1.9310 90.4635 1.9570 91.5570 ;
        RECT 1.8230 90.4635 1.8490 91.5570 ;
        RECT 1.7150 90.4635 1.7410 91.5570 ;
        RECT 1.6070 90.4635 1.6330 91.5570 ;
        RECT 1.4990 90.4635 1.5250 91.5570 ;
        RECT 1.3910 90.4635 1.4170 91.5570 ;
        RECT 1.2830 90.4635 1.3090 91.5570 ;
        RECT 1.1750 90.4635 1.2010 91.5570 ;
        RECT 1.0670 90.4635 1.0930 91.5570 ;
        RECT 0.9590 90.4635 0.9850 91.5570 ;
        RECT 0.8510 90.4635 0.8770 91.5570 ;
        RECT 0.7430 90.4635 0.7690 91.5570 ;
        RECT 0.6350 90.4635 0.6610 91.5570 ;
        RECT 0.5270 90.4635 0.5530 91.5570 ;
        RECT 0.4190 90.4635 0.4450 91.5570 ;
        RECT 0.3110 90.4635 0.3370 91.5570 ;
        RECT 0.2030 90.4635 0.2290 91.5570 ;
        RECT 0.0000 90.4635 0.0850 91.5570 ;
        RECT 5.1800 91.5435 5.3080 92.6370 ;
        RECT 5.1660 92.2090 5.3080 92.5315 ;
        RECT 5.0180 91.9360 5.0800 92.6370 ;
        RECT 5.0040 92.2455 5.0800 92.3990 ;
        RECT 5.0180 91.5435 5.0440 92.6370 ;
        RECT 5.0180 91.6645 5.0580 91.9040 ;
        RECT 5.0180 91.5435 5.0800 91.6325 ;
        RECT 4.7210 91.9940 4.9270 92.6370 ;
        RECT 4.9010 91.5435 4.9270 92.6370 ;
        RECT 4.7210 92.2710 4.9410 92.5290 ;
        RECT 4.7210 91.5435 4.8190 92.6370 ;
        RECT 4.3040 91.5435 4.3870 92.6370 ;
        RECT 4.3040 91.6320 4.4010 92.5675 ;
        RECT 9.5270 91.5435 9.6120 92.6370 ;
        RECT 9.3830 91.5435 9.4090 92.6370 ;
        RECT 9.2750 91.5435 9.3010 92.6370 ;
        RECT 9.1670 91.5435 9.1930 92.6370 ;
        RECT 9.0590 91.5435 9.0850 92.6370 ;
        RECT 8.9510 91.5435 8.9770 92.6370 ;
        RECT 8.8430 91.5435 8.8690 92.6370 ;
        RECT 8.7350 91.5435 8.7610 92.6370 ;
        RECT 8.6270 91.5435 8.6530 92.6370 ;
        RECT 8.5190 91.5435 8.5450 92.6370 ;
        RECT 8.4110 91.5435 8.4370 92.6370 ;
        RECT 8.3030 91.5435 8.3290 92.6370 ;
        RECT 8.1950 91.5435 8.2210 92.6370 ;
        RECT 8.0870 91.5435 8.1130 92.6370 ;
        RECT 7.9790 91.5435 8.0050 92.6370 ;
        RECT 7.8710 91.5435 7.8970 92.6370 ;
        RECT 7.7630 91.5435 7.7890 92.6370 ;
        RECT 7.6550 91.5435 7.6810 92.6370 ;
        RECT 7.5470 91.5435 7.5730 92.6370 ;
        RECT 7.4390 91.5435 7.4650 92.6370 ;
        RECT 7.3310 91.5435 7.3570 92.6370 ;
        RECT 7.2230 91.5435 7.2490 92.6370 ;
        RECT 7.1150 91.5435 7.1410 92.6370 ;
        RECT 7.0070 91.5435 7.0330 92.6370 ;
        RECT 6.8990 91.5435 6.9250 92.6370 ;
        RECT 6.7910 91.5435 6.8170 92.6370 ;
        RECT 6.6830 91.5435 6.7090 92.6370 ;
        RECT 6.5750 91.5435 6.6010 92.6370 ;
        RECT 6.4670 91.5435 6.4930 92.6370 ;
        RECT 6.3590 91.5435 6.3850 92.6370 ;
        RECT 6.2510 91.5435 6.2770 92.6370 ;
        RECT 6.1430 91.5435 6.1690 92.6370 ;
        RECT 6.0350 91.5435 6.0610 92.6370 ;
        RECT 5.9270 91.5435 5.9530 92.6370 ;
        RECT 5.7140 91.5435 5.7910 92.6370 ;
        RECT 3.8210 91.5435 3.8980 92.6370 ;
        RECT 3.6590 91.5435 3.6850 92.6370 ;
        RECT 3.5510 91.5435 3.5770 92.6370 ;
        RECT 3.4430 91.5435 3.4690 92.6370 ;
        RECT 3.3350 91.5435 3.3610 92.6370 ;
        RECT 3.2270 91.5435 3.2530 92.6370 ;
        RECT 3.1190 91.5435 3.1450 92.6370 ;
        RECT 3.0110 91.5435 3.0370 92.6370 ;
        RECT 2.9030 91.5435 2.9290 92.6370 ;
        RECT 2.7950 91.5435 2.8210 92.6370 ;
        RECT 2.6870 91.5435 2.7130 92.6370 ;
        RECT 2.5790 91.5435 2.6050 92.6370 ;
        RECT 2.4710 91.5435 2.4970 92.6370 ;
        RECT 2.3630 91.5435 2.3890 92.6370 ;
        RECT 2.2550 91.5435 2.2810 92.6370 ;
        RECT 2.1470 91.5435 2.1730 92.6370 ;
        RECT 2.0390 91.5435 2.0650 92.6370 ;
        RECT 1.9310 91.5435 1.9570 92.6370 ;
        RECT 1.8230 91.5435 1.8490 92.6370 ;
        RECT 1.7150 91.5435 1.7410 92.6370 ;
        RECT 1.6070 91.5435 1.6330 92.6370 ;
        RECT 1.4990 91.5435 1.5250 92.6370 ;
        RECT 1.3910 91.5435 1.4170 92.6370 ;
        RECT 1.2830 91.5435 1.3090 92.6370 ;
        RECT 1.1750 91.5435 1.2010 92.6370 ;
        RECT 1.0670 91.5435 1.0930 92.6370 ;
        RECT 0.9590 91.5435 0.9850 92.6370 ;
        RECT 0.8510 91.5435 0.8770 92.6370 ;
        RECT 0.7430 91.5435 0.7690 92.6370 ;
        RECT 0.6350 91.5435 0.6610 92.6370 ;
        RECT 0.5270 91.5435 0.5530 92.6370 ;
        RECT 0.4190 91.5435 0.4450 92.6370 ;
        RECT 0.3110 91.5435 0.3370 92.6370 ;
        RECT 0.2030 91.5435 0.2290 92.6370 ;
        RECT 0.0000 91.5435 0.0850 92.6370 ;
        RECT 5.1800 92.6235 5.3080 93.7170 ;
        RECT 5.1660 93.2890 5.3080 93.6115 ;
        RECT 5.0180 93.0160 5.0800 93.7170 ;
        RECT 5.0040 93.3255 5.0800 93.4790 ;
        RECT 5.0180 92.6235 5.0440 93.7170 ;
        RECT 5.0180 92.7445 5.0580 92.9840 ;
        RECT 5.0180 92.6235 5.0800 92.7125 ;
        RECT 4.7210 93.0740 4.9270 93.7170 ;
        RECT 4.9010 92.6235 4.9270 93.7170 ;
        RECT 4.7210 93.3510 4.9410 93.6090 ;
        RECT 4.7210 92.6235 4.8190 93.7170 ;
        RECT 4.3040 92.6235 4.3870 93.7170 ;
        RECT 4.3040 92.7120 4.4010 93.6475 ;
        RECT 9.5270 92.6235 9.6120 93.7170 ;
        RECT 9.3830 92.6235 9.4090 93.7170 ;
        RECT 9.2750 92.6235 9.3010 93.7170 ;
        RECT 9.1670 92.6235 9.1930 93.7170 ;
        RECT 9.0590 92.6235 9.0850 93.7170 ;
        RECT 8.9510 92.6235 8.9770 93.7170 ;
        RECT 8.8430 92.6235 8.8690 93.7170 ;
        RECT 8.7350 92.6235 8.7610 93.7170 ;
        RECT 8.6270 92.6235 8.6530 93.7170 ;
        RECT 8.5190 92.6235 8.5450 93.7170 ;
        RECT 8.4110 92.6235 8.4370 93.7170 ;
        RECT 8.3030 92.6235 8.3290 93.7170 ;
        RECT 8.1950 92.6235 8.2210 93.7170 ;
        RECT 8.0870 92.6235 8.1130 93.7170 ;
        RECT 7.9790 92.6235 8.0050 93.7170 ;
        RECT 7.8710 92.6235 7.8970 93.7170 ;
        RECT 7.7630 92.6235 7.7890 93.7170 ;
        RECT 7.6550 92.6235 7.6810 93.7170 ;
        RECT 7.5470 92.6235 7.5730 93.7170 ;
        RECT 7.4390 92.6235 7.4650 93.7170 ;
        RECT 7.3310 92.6235 7.3570 93.7170 ;
        RECT 7.2230 92.6235 7.2490 93.7170 ;
        RECT 7.1150 92.6235 7.1410 93.7170 ;
        RECT 7.0070 92.6235 7.0330 93.7170 ;
        RECT 6.8990 92.6235 6.9250 93.7170 ;
        RECT 6.7910 92.6235 6.8170 93.7170 ;
        RECT 6.6830 92.6235 6.7090 93.7170 ;
        RECT 6.5750 92.6235 6.6010 93.7170 ;
        RECT 6.4670 92.6235 6.4930 93.7170 ;
        RECT 6.3590 92.6235 6.3850 93.7170 ;
        RECT 6.2510 92.6235 6.2770 93.7170 ;
        RECT 6.1430 92.6235 6.1690 93.7170 ;
        RECT 6.0350 92.6235 6.0610 93.7170 ;
        RECT 5.9270 92.6235 5.9530 93.7170 ;
        RECT 5.7140 92.6235 5.7910 93.7170 ;
        RECT 3.8210 92.6235 3.8980 93.7170 ;
        RECT 3.6590 92.6235 3.6850 93.7170 ;
        RECT 3.5510 92.6235 3.5770 93.7170 ;
        RECT 3.4430 92.6235 3.4690 93.7170 ;
        RECT 3.3350 92.6235 3.3610 93.7170 ;
        RECT 3.2270 92.6235 3.2530 93.7170 ;
        RECT 3.1190 92.6235 3.1450 93.7170 ;
        RECT 3.0110 92.6235 3.0370 93.7170 ;
        RECT 2.9030 92.6235 2.9290 93.7170 ;
        RECT 2.7950 92.6235 2.8210 93.7170 ;
        RECT 2.6870 92.6235 2.7130 93.7170 ;
        RECT 2.5790 92.6235 2.6050 93.7170 ;
        RECT 2.4710 92.6235 2.4970 93.7170 ;
        RECT 2.3630 92.6235 2.3890 93.7170 ;
        RECT 2.2550 92.6235 2.2810 93.7170 ;
        RECT 2.1470 92.6235 2.1730 93.7170 ;
        RECT 2.0390 92.6235 2.0650 93.7170 ;
        RECT 1.9310 92.6235 1.9570 93.7170 ;
        RECT 1.8230 92.6235 1.8490 93.7170 ;
        RECT 1.7150 92.6235 1.7410 93.7170 ;
        RECT 1.6070 92.6235 1.6330 93.7170 ;
        RECT 1.4990 92.6235 1.5250 93.7170 ;
        RECT 1.3910 92.6235 1.4170 93.7170 ;
        RECT 1.2830 92.6235 1.3090 93.7170 ;
        RECT 1.1750 92.6235 1.2010 93.7170 ;
        RECT 1.0670 92.6235 1.0930 93.7170 ;
        RECT 0.9590 92.6235 0.9850 93.7170 ;
        RECT 0.8510 92.6235 0.8770 93.7170 ;
        RECT 0.7430 92.6235 0.7690 93.7170 ;
        RECT 0.6350 92.6235 0.6610 93.7170 ;
        RECT 0.5270 92.6235 0.5530 93.7170 ;
        RECT 0.4190 92.6235 0.4450 93.7170 ;
        RECT 0.3110 92.6235 0.3370 93.7170 ;
        RECT 0.2030 92.6235 0.2290 93.7170 ;
        RECT 0.0000 92.6235 0.0850 93.7170 ;
        RECT 5.1800 93.7035 5.3080 94.7970 ;
        RECT 5.1660 94.3690 5.3080 94.6915 ;
        RECT 5.0180 94.0960 5.0800 94.7970 ;
        RECT 5.0040 94.4055 5.0800 94.5590 ;
        RECT 5.0180 93.7035 5.0440 94.7970 ;
        RECT 5.0180 93.8245 5.0580 94.0640 ;
        RECT 5.0180 93.7035 5.0800 93.7925 ;
        RECT 4.7210 94.1540 4.9270 94.7970 ;
        RECT 4.9010 93.7035 4.9270 94.7970 ;
        RECT 4.7210 94.4310 4.9410 94.6890 ;
        RECT 4.7210 93.7035 4.8190 94.7970 ;
        RECT 4.3040 93.7035 4.3870 94.7970 ;
        RECT 4.3040 93.7920 4.4010 94.7275 ;
        RECT 9.5270 93.7035 9.6120 94.7970 ;
        RECT 9.3830 93.7035 9.4090 94.7970 ;
        RECT 9.2750 93.7035 9.3010 94.7970 ;
        RECT 9.1670 93.7035 9.1930 94.7970 ;
        RECT 9.0590 93.7035 9.0850 94.7970 ;
        RECT 8.9510 93.7035 8.9770 94.7970 ;
        RECT 8.8430 93.7035 8.8690 94.7970 ;
        RECT 8.7350 93.7035 8.7610 94.7970 ;
        RECT 8.6270 93.7035 8.6530 94.7970 ;
        RECT 8.5190 93.7035 8.5450 94.7970 ;
        RECT 8.4110 93.7035 8.4370 94.7970 ;
        RECT 8.3030 93.7035 8.3290 94.7970 ;
        RECT 8.1950 93.7035 8.2210 94.7970 ;
        RECT 8.0870 93.7035 8.1130 94.7970 ;
        RECT 7.9790 93.7035 8.0050 94.7970 ;
        RECT 7.8710 93.7035 7.8970 94.7970 ;
        RECT 7.7630 93.7035 7.7890 94.7970 ;
        RECT 7.6550 93.7035 7.6810 94.7970 ;
        RECT 7.5470 93.7035 7.5730 94.7970 ;
        RECT 7.4390 93.7035 7.4650 94.7970 ;
        RECT 7.3310 93.7035 7.3570 94.7970 ;
        RECT 7.2230 93.7035 7.2490 94.7970 ;
        RECT 7.1150 93.7035 7.1410 94.7970 ;
        RECT 7.0070 93.7035 7.0330 94.7970 ;
        RECT 6.8990 93.7035 6.9250 94.7970 ;
        RECT 6.7910 93.7035 6.8170 94.7970 ;
        RECT 6.6830 93.7035 6.7090 94.7970 ;
        RECT 6.5750 93.7035 6.6010 94.7970 ;
        RECT 6.4670 93.7035 6.4930 94.7970 ;
        RECT 6.3590 93.7035 6.3850 94.7970 ;
        RECT 6.2510 93.7035 6.2770 94.7970 ;
        RECT 6.1430 93.7035 6.1690 94.7970 ;
        RECT 6.0350 93.7035 6.0610 94.7970 ;
        RECT 5.9270 93.7035 5.9530 94.7970 ;
        RECT 5.7140 93.7035 5.7910 94.7970 ;
        RECT 3.8210 93.7035 3.8980 94.7970 ;
        RECT 3.6590 93.7035 3.6850 94.7970 ;
        RECT 3.5510 93.7035 3.5770 94.7970 ;
        RECT 3.4430 93.7035 3.4690 94.7970 ;
        RECT 3.3350 93.7035 3.3610 94.7970 ;
        RECT 3.2270 93.7035 3.2530 94.7970 ;
        RECT 3.1190 93.7035 3.1450 94.7970 ;
        RECT 3.0110 93.7035 3.0370 94.7970 ;
        RECT 2.9030 93.7035 2.9290 94.7970 ;
        RECT 2.7950 93.7035 2.8210 94.7970 ;
        RECT 2.6870 93.7035 2.7130 94.7970 ;
        RECT 2.5790 93.7035 2.6050 94.7970 ;
        RECT 2.4710 93.7035 2.4970 94.7970 ;
        RECT 2.3630 93.7035 2.3890 94.7970 ;
        RECT 2.2550 93.7035 2.2810 94.7970 ;
        RECT 2.1470 93.7035 2.1730 94.7970 ;
        RECT 2.0390 93.7035 2.0650 94.7970 ;
        RECT 1.9310 93.7035 1.9570 94.7970 ;
        RECT 1.8230 93.7035 1.8490 94.7970 ;
        RECT 1.7150 93.7035 1.7410 94.7970 ;
        RECT 1.6070 93.7035 1.6330 94.7970 ;
        RECT 1.4990 93.7035 1.5250 94.7970 ;
        RECT 1.3910 93.7035 1.4170 94.7970 ;
        RECT 1.2830 93.7035 1.3090 94.7970 ;
        RECT 1.1750 93.7035 1.2010 94.7970 ;
        RECT 1.0670 93.7035 1.0930 94.7970 ;
        RECT 0.9590 93.7035 0.9850 94.7970 ;
        RECT 0.8510 93.7035 0.8770 94.7970 ;
        RECT 0.7430 93.7035 0.7690 94.7970 ;
        RECT 0.6350 93.7035 0.6610 94.7970 ;
        RECT 0.5270 93.7035 0.5530 94.7970 ;
        RECT 0.4190 93.7035 0.4450 94.7970 ;
        RECT 0.3110 93.7035 0.3370 94.7970 ;
        RECT 0.2030 93.7035 0.2290 94.7970 ;
        RECT 0.0000 93.7035 0.0850 94.7970 ;
  LAYER V3  ;
      RECT 0.0000 1.2200 9.6120 1.3500 ;
      RECT 9.4950 0.2565 9.6120 1.3500 ;
      RECT 5.8410 1.1240 9.4770 1.3500 ;
      RECT 4.5090 1.1240 5.8230 1.3500 ;
      RECT 3.7890 0.2565 4.4190 1.3500 ;
      RECT 0.1350 1.1240 3.7710 1.3500 ;
      RECT 0.0000 0.2565 0.1170 1.3500 ;
      RECT 9.4590 0.2565 9.6120 1.1720 ;
      RECT 5.8950 0.2565 9.4410 1.3500 ;
      RECT 5.1480 0.2565 5.8770 1.1720 ;
      RECT 4.9860 0.4520 5.1120 1.3500 ;
      RECT 3.7350 0.3560 4.9590 1.1720 ;
      RECT 0.1710 0.2565 3.7170 1.3500 ;
      RECT 0.0000 0.2565 0.1530 1.1720 ;
      RECT 5.0940 0.2565 9.6120 1.0760 ;
      RECT 0.0000 0.3560 5.0760 1.0760 ;
      RECT 4.8690 0.2565 9.6120 0.4280 ;
      RECT 0.0000 0.2565 4.8510 1.0760 ;
      RECT 0.0000 0.2565 9.6120 0.3320 ;
      RECT 0.0000 2.3000 9.6120 2.4300 ;
      RECT 9.4950 1.3365 9.6120 2.4300 ;
      RECT 5.8410 2.2040 9.4770 2.4300 ;
      RECT 4.5090 2.2040 5.8230 2.4300 ;
      RECT 3.7890 1.3365 4.4190 2.4300 ;
      RECT 0.1350 2.2040 3.7710 2.4300 ;
      RECT 0.0000 1.3365 0.1170 2.4300 ;
      RECT 9.4590 1.3365 9.6120 2.2520 ;
      RECT 5.8950 1.3365 9.4410 2.4300 ;
      RECT 5.1480 1.3365 5.8770 2.2520 ;
      RECT 4.9860 1.5320 5.1120 2.4300 ;
      RECT 3.7350 1.4360 4.9590 2.2520 ;
      RECT 0.1710 1.3365 3.7170 2.4300 ;
      RECT 0.0000 1.3365 0.1530 2.2520 ;
      RECT 5.0940 1.3365 9.6120 2.1560 ;
      RECT 0.0000 1.4360 5.0760 2.1560 ;
      RECT 4.8690 1.3365 9.6120 1.5080 ;
      RECT 0.0000 1.3365 4.8510 2.1560 ;
      RECT 0.0000 1.3365 9.6120 1.4120 ;
      RECT 0.0000 3.3800 9.6120 3.5100 ;
      RECT 9.4950 2.4165 9.6120 3.5100 ;
      RECT 5.8410 3.2840 9.4770 3.5100 ;
      RECT 4.5090 3.2840 5.8230 3.5100 ;
      RECT 3.7890 2.4165 4.4190 3.5100 ;
      RECT 0.1350 3.2840 3.7710 3.5100 ;
      RECT 0.0000 2.4165 0.1170 3.5100 ;
      RECT 9.4590 2.4165 9.6120 3.3320 ;
      RECT 5.8950 2.4165 9.4410 3.5100 ;
      RECT 5.1480 2.4165 5.8770 3.3320 ;
      RECT 4.9860 2.6120 5.1120 3.5100 ;
      RECT 3.7350 2.5160 4.9590 3.3320 ;
      RECT 0.1710 2.4165 3.7170 3.5100 ;
      RECT 0.0000 2.4165 0.1530 3.3320 ;
      RECT 5.0940 2.4165 9.6120 3.2360 ;
      RECT 0.0000 2.5160 5.0760 3.2360 ;
      RECT 4.8690 2.4165 9.6120 2.5880 ;
      RECT 0.0000 2.4165 4.8510 3.2360 ;
      RECT 0.0000 2.4165 9.6120 2.4920 ;
      RECT 0.0000 4.4600 9.6120 4.5900 ;
      RECT 9.4950 3.4965 9.6120 4.5900 ;
      RECT 5.8410 4.3640 9.4770 4.5900 ;
      RECT 4.5090 4.3640 5.8230 4.5900 ;
      RECT 3.7890 3.4965 4.4190 4.5900 ;
      RECT 0.1350 4.3640 3.7710 4.5900 ;
      RECT 0.0000 3.4965 0.1170 4.5900 ;
      RECT 9.4590 3.4965 9.6120 4.4120 ;
      RECT 5.8950 3.4965 9.4410 4.5900 ;
      RECT 5.1480 3.4965 5.8770 4.4120 ;
      RECT 4.9860 3.6920 5.1120 4.5900 ;
      RECT 3.7350 3.5960 4.9590 4.4120 ;
      RECT 0.1710 3.4965 3.7170 4.5900 ;
      RECT 0.0000 3.4965 0.1530 4.4120 ;
      RECT 5.0940 3.4965 9.6120 4.3160 ;
      RECT 0.0000 3.5960 5.0760 4.3160 ;
      RECT 4.8690 3.4965 9.6120 3.6680 ;
      RECT 0.0000 3.4965 4.8510 4.3160 ;
      RECT 0.0000 3.4965 9.6120 3.5720 ;
      RECT 0.0000 5.5400 9.6120 5.6700 ;
      RECT 9.4950 4.5765 9.6120 5.6700 ;
      RECT 5.8410 5.4440 9.4770 5.6700 ;
      RECT 4.5090 5.4440 5.8230 5.6700 ;
      RECT 3.7890 4.5765 4.4190 5.6700 ;
      RECT 0.1350 5.4440 3.7710 5.6700 ;
      RECT 0.0000 4.5765 0.1170 5.6700 ;
      RECT 9.4590 4.5765 9.6120 5.4920 ;
      RECT 5.8950 4.5765 9.4410 5.6700 ;
      RECT 5.1480 4.5765 5.8770 5.4920 ;
      RECT 4.9860 4.7720 5.1120 5.6700 ;
      RECT 3.7350 4.6760 4.9590 5.4920 ;
      RECT 0.1710 4.5765 3.7170 5.6700 ;
      RECT 0.0000 4.5765 0.1530 5.4920 ;
      RECT 5.0940 4.5765 9.6120 5.3960 ;
      RECT 0.0000 4.6760 5.0760 5.3960 ;
      RECT 4.8690 4.5765 9.6120 4.7480 ;
      RECT 0.0000 4.5765 4.8510 5.3960 ;
      RECT 0.0000 4.5765 9.6120 4.6520 ;
      RECT 0.0000 6.6200 9.6120 6.7500 ;
      RECT 9.4950 5.6565 9.6120 6.7500 ;
      RECT 5.8410 6.5240 9.4770 6.7500 ;
      RECT 4.5090 6.5240 5.8230 6.7500 ;
      RECT 3.7890 5.6565 4.4190 6.7500 ;
      RECT 0.1350 6.5240 3.7710 6.7500 ;
      RECT 0.0000 5.6565 0.1170 6.7500 ;
      RECT 9.4590 5.6565 9.6120 6.5720 ;
      RECT 5.8950 5.6565 9.4410 6.7500 ;
      RECT 5.1480 5.6565 5.8770 6.5720 ;
      RECT 4.9860 5.8520 5.1120 6.7500 ;
      RECT 3.7350 5.7560 4.9590 6.5720 ;
      RECT 0.1710 5.6565 3.7170 6.7500 ;
      RECT 0.0000 5.6565 0.1530 6.5720 ;
      RECT 5.0940 5.6565 9.6120 6.4760 ;
      RECT 0.0000 5.7560 5.0760 6.4760 ;
      RECT 4.8690 5.6565 9.6120 5.8280 ;
      RECT 0.0000 5.6565 4.8510 6.4760 ;
      RECT 0.0000 5.6565 9.6120 5.7320 ;
      RECT 0.0000 7.7000 9.6120 7.8300 ;
      RECT 9.4950 6.7365 9.6120 7.8300 ;
      RECT 5.8410 7.6040 9.4770 7.8300 ;
      RECT 4.5090 7.6040 5.8230 7.8300 ;
      RECT 3.7890 6.7365 4.4190 7.8300 ;
      RECT 0.1350 7.6040 3.7710 7.8300 ;
      RECT 0.0000 6.7365 0.1170 7.8300 ;
      RECT 9.4590 6.7365 9.6120 7.6520 ;
      RECT 5.8950 6.7365 9.4410 7.8300 ;
      RECT 5.1480 6.7365 5.8770 7.6520 ;
      RECT 4.9860 6.9320 5.1120 7.8300 ;
      RECT 3.7350 6.8360 4.9590 7.6520 ;
      RECT 0.1710 6.7365 3.7170 7.8300 ;
      RECT 0.0000 6.7365 0.1530 7.6520 ;
      RECT 5.0940 6.7365 9.6120 7.5560 ;
      RECT 0.0000 6.8360 5.0760 7.5560 ;
      RECT 4.8690 6.7365 9.6120 6.9080 ;
      RECT 0.0000 6.7365 4.8510 7.5560 ;
      RECT 0.0000 6.7365 9.6120 6.8120 ;
      RECT 0.0000 8.7800 9.6120 8.9100 ;
      RECT 9.4950 7.8165 9.6120 8.9100 ;
      RECT 5.8410 8.6840 9.4770 8.9100 ;
      RECT 4.5090 8.6840 5.8230 8.9100 ;
      RECT 3.7890 7.8165 4.4190 8.9100 ;
      RECT 0.1350 8.6840 3.7710 8.9100 ;
      RECT 0.0000 7.8165 0.1170 8.9100 ;
      RECT 9.4590 7.8165 9.6120 8.7320 ;
      RECT 5.8950 7.8165 9.4410 8.9100 ;
      RECT 5.1480 7.8165 5.8770 8.7320 ;
      RECT 4.9860 8.0120 5.1120 8.9100 ;
      RECT 3.7350 7.9160 4.9590 8.7320 ;
      RECT 0.1710 7.8165 3.7170 8.9100 ;
      RECT 0.0000 7.8165 0.1530 8.7320 ;
      RECT 5.0940 7.8165 9.6120 8.6360 ;
      RECT 0.0000 7.9160 5.0760 8.6360 ;
      RECT 4.8690 7.8165 9.6120 7.9880 ;
      RECT 0.0000 7.8165 4.8510 8.6360 ;
      RECT 0.0000 7.8165 9.6120 7.8920 ;
      RECT 0.0000 9.8600 9.6120 9.9900 ;
      RECT 9.4950 8.8965 9.6120 9.9900 ;
      RECT 5.8410 9.7640 9.4770 9.9900 ;
      RECT 4.5090 9.7640 5.8230 9.9900 ;
      RECT 3.7890 8.8965 4.4190 9.9900 ;
      RECT 0.1350 9.7640 3.7710 9.9900 ;
      RECT 0.0000 8.8965 0.1170 9.9900 ;
      RECT 9.4590 8.8965 9.6120 9.8120 ;
      RECT 5.8950 8.8965 9.4410 9.9900 ;
      RECT 5.1480 8.8965 5.8770 9.8120 ;
      RECT 4.9860 9.0920 5.1120 9.9900 ;
      RECT 3.7350 8.9960 4.9590 9.8120 ;
      RECT 0.1710 8.8965 3.7170 9.9900 ;
      RECT 0.0000 8.8965 0.1530 9.8120 ;
      RECT 5.0940 8.8965 9.6120 9.7160 ;
      RECT 0.0000 8.9960 5.0760 9.7160 ;
      RECT 4.8690 8.8965 9.6120 9.0680 ;
      RECT 0.0000 8.8965 4.8510 9.7160 ;
      RECT 0.0000 8.8965 9.6120 8.9720 ;
      RECT 0.0000 10.9400 9.6120 11.0700 ;
      RECT 9.4950 9.9765 9.6120 11.0700 ;
      RECT 5.8410 10.8440 9.4770 11.0700 ;
      RECT 4.5090 10.8440 5.8230 11.0700 ;
      RECT 3.7890 9.9765 4.4190 11.0700 ;
      RECT 0.1350 10.8440 3.7710 11.0700 ;
      RECT 0.0000 9.9765 0.1170 11.0700 ;
      RECT 9.4590 9.9765 9.6120 10.8920 ;
      RECT 5.8950 9.9765 9.4410 11.0700 ;
      RECT 5.1480 9.9765 5.8770 10.8920 ;
      RECT 4.9860 10.1720 5.1120 11.0700 ;
      RECT 3.7350 10.0760 4.9590 10.8920 ;
      RECT 0.1710 9.9765 3.7170 11.0700 ;
      RECT 0.0000 9.9765 0.1530 10.8920 ;
      RECT 5.0940 9.9765 9.6120 10.7960 ;
      RECT 0.0000 10.0760 5.0760 10.7960 ;
      RECT 4.8690 9.9765 9.6120 10.1480 ;
      RECT 0.0000 9.9765 4.8510 10.7960 ;
      RECT 0.0000 9.9765 9.6120 10.0520 ;
      RECT 0.0000 12.0200 9.6120 12.1500 ;
      RECT 9.4950 11.0565 9.6120 12.1500 ;
      RECT 5.8410 11.9240 9.4770 12.1500 ;
      RECT 4.5090 11.9240 5.8230 12.1500 ;
      RECT 3.7890 11.0565 4.4190 12.1500 ;
      RECT 0.1350 11.9240 3.7710 12.1500 ;
      RECT 0.0000 11.0565 0.1170 12.1500 ;
      RECT 9.4590 11.0565 9.6120 11.9720 ;
      RECT 5.8950 11.0565 9.4410 12.1500 ;
      RECT 5.1480 11.0565 5.8770 11.9720 ;
      RECT 4.9860 11.2520 5.1120 12.1500 ;
      RECT 3.7350 11.1560 4.9590 11.9720 ;
      RECT 0.1710 11.0565 3.7170 12.1500 ;
      RECT 0.0000 11.0565 0.1530 11.9720 ;
      RECT 5.0940 11.0565 9.6120 11.8760 ;
      RECT 0.0000 11.1560 5.0760 11.8760 ;
      RECT 4.8690 11.0565 9.6120 11.2280 ;
      RECT 0.0000 11.0565 4.8510 11.8760 ;
      RECT 0.0000 11.0565 9.6120 11.1320 ;
      RECT 0.0000 13.1000 9.6120 13.2300 ;
      RECT 9.4950 12.1365 9.6120 13.2300 ;
      RECT 5.8410 13.0040 9.4770 13.2300 ;
      RECT 4.5090 13.0040 5.8230 13.2300 ;
      RECT 3.7890 12.1365 4.4190 13.2300 ;
      RECT 0.1350 13.0040 3.7710 13.2300 ;
      RECT 0.0000 12.1365 0.1170 13.2300 ;
      RECT 9.4590 12.1365 9.6120 13.0520 ;
      RECT 5.8950 12.1365 9.4410 13.2300 ;
      RECT 5.1480 12.1365 5.8770 13.0520 ;
      RECT 4.9860 12.3320 5.1120 13.2300 ;
      RECT 3.7350 12.2360 4.9590 13.0520 ;
      RECT 0.1710 12.1365 3.7170 13.2300 ;
      RECT 0.0000 12.1365 0.1530 13.0520 ;
      RECT 5.0940 12.1365 9.6120 12.9560 ;
      RECT 0.0000 12.2360 5.0760 12.9560 ;
      RECT 4.8690 12.1365 9.6120 12.3080 ;
      RECT 0.0000 12.1365 4.8510 12.9560 ;
      RECT 0.0000 12.1365 9.6120 12.2120 ;
      RECT 0.0000 14.1800 9.6120 14.3100 ;
      RECT 9.4950 13.2165 9.6120 14.3100 ;
      RECT 5.8410 14.0840 9.4770 14.3100 ;
      RECT 4.5090 14.0840 5.8230 14.3100 ;
      RECT 3.7890 13.2165 4.4190 14.3100 ;
      RECT 0.1350 14.0840 3.7710 14.3100 ;
      RECT 0.0000 13.2165 0.1170 14.3100 ;
      RECT 9.4590 13.2165 9.6120 14.1320 ;
      RECT 5.8950 13.2165 9.4410 14.3100 ;
      RECT 5.1480 13.2165 5.8770 14.1320 ;
      RECT 4.9860 13.4120 5.1120 14.3100 ;
      RECT 3.7350 13.3160 4.9590 14.1320 ;
      RECT 0.1710 13.2165 3.7170 14.3100 ;
      RECT 0.0000 13.2165 0.1530 14.1320 ;
      RECT 5.0940 13.2165 9.6120 14.0360 ;
      RECT 0.0000 13.3160 5.0760 14.0360 ;
      RECT 4.8690 13.2165 9.6120 13.3880 ;
      RECT 0.0000 13.2165 4.8510 14.0360 ;
      RECT 0.0000 13.2165 9.6120 13.2920 ;
      RECT 0.0000 15.2600 9.6120 15.3900 ;
      RECT 9.4950 14.2965 9.6120 15.3900 ;
      RECT 5.8410 15.1640 9.4770 15.3900 ;
      RECT 4.5090 15.1640 5.8230 15.3900 ;
      RECT 3.7890 14.2965 4.4190 15.3900 ;
      RECT 0.1350 15.1640 3.7710 15.3900 ;
      RECT 0.0000 14.2965 0.1170 15.3900 ;
      RECT 9.4590 14.2965 9.6120 15.2120 ;
      RECT 5.8950 14.2965 9.4410 15.3900 ;
      RECT 5.1480 14.2965 5.8770 15.2120 ;
      RECT 4.9860 14.4920 5.1120 15.3900 ;
      RECT 3.7350 14.3960 4.9590 15.2120 ;
      RECT 0.1710 14.2965 3.7170 15.3900 ;
      RECT 0.0000 14.2965 0.1530 15.2120 ;
      RECT 5.0940 14.2965 9.6120 15.1160 ;
      RECT 0.0000 14.3960 5.0760 15.1160 ;
      RECT 4.8690 14.2965 9.6120 14.4680 ;
      RECT 0.0000 14.2965 4.8510 15.1160 ;
      RECT 0.0000 14.2965 9.6120 14.3720 ;
      RECT 0.0000 16.3400 9.6120 16.4700 ;
      RECT 9.4950 15.3765 9.6120 16.4700 ;
      RECT 5.8410 16.2440 9.4770 16.4700 ;
      RECT 4.5090 16.2440 5.8230 16.4700 ;
      RECT 3.7890 15.3765 4.4190 16.4700 ;
      RECT 0.1350 16.2440 3.7710 16.4700 ;
      RECT 0.0000 15.3765 0.1170 16.4700 ;
      RECT 9.4590 15.3765 9.6120 16.2920 ;
      RECT 5.8950 15.3765 9.4410 16.4700 ;
      RECT 5.1480 15.3765 5.8770 16.2920 ;
      RECT 4.9860 15.5720 5.1120 16.4700 ;
      RECT 3.7350 15.4760 4.9590 16.2920 ;
      RECT 0.1710 15.3765 3.7170 16.4700 ;
      RECT 0.0000 15.3765 0.1530 16.2920 ;
      RECT 5.0940 15.3765 9.6120 16.1960 ;
      RECT 0.0000 15.4760 5.0760 16.1960 ;
      RECT 4.8690 15.3765 9.6120 15.5480 ;
      RECT 0.0000 15.3765 4.8510 16.1960 ;
      RECT 0.0000 15.3765 9.6120 15.4520 ;
      RECT 0.0000 17.4200 9.6120 17.5500 ;
      RECT 9.4950 16.4565 9.6120 17.5500 ;
      RECT 5.8410 17.3240 9.4770 17.5500 ;
      RECT 4.5090 17.3240 5.8230 17.5500 ;
      RECT 3.7890 16.4565 4.4190 17.5500 ;
      RECT 0.1350 17.3240 3.7710 17.5500 ;
      RECT 0.0000 16.4565 0.1170 17.5500 ;
      RECT 9.4590 16.4565 9.6120 17.3720 ;
      RECT 5.8950 16.4565 9.4410 17.5500 ;
      RECT 5.1480 16.4565 5.8770 17.3720 ;
      RECT 4.9860 16.6520 5.1120 17.5500 ;
      RECT 3.7350 16.5560 4.9590 17.3720 ;
      RECT 0.1710 16.4565 3.7170 17.5500 ;
      RECT 0.0000 16.4565 0.1530 17.3720 ;
      RECT 5.0940 16.4565 9.6120 17.2760 ;
      RECT 0.0000 16.5560 5.0760 17.2760 ;
      RECT 4.8690 16.4565 9.6120 16.6280 ;
      RECT 0.0000 16.4565 4.8510 17.2760 ;
      RECT 0.0000 16.4565 9.6120 16.5320 ;
      RECT 0.0000 18.5000 9.6120 18.6300 ;
      RECT 9.4950 17.5365 9.6120 18.6300 ;
      RECT 5.8410 18.4040 9.4770 18.6300 ;
      RECT 4.5090 18.4040 5.8230 18.6300 ;
      RECT 3.7890 17.5365 4.4190 18.6300 ;
      RECT 0.1350 18.4040 3.7710 18.6300 ;
      RECT 0.0000 17.5365 0.1170 18.6300 ;
      RECT 9.4590 17.5365 9.6120 18.4520 ;
      RECT 5.8950 17.5365 9.4410 18.6300 ;
      RECT 5.1480 17.5365 5.8770 18.4520 ;
      RECT 4.9860 17.7320 5.1120 18.6300 ;
      RECT 3.7350 17.6360 4.9590 18.4520 ;
      RECT 0.1710 17.5365 3.7170 18.6300 ;
      RECT 0.0000 17.5365 0.1530 18.4520 ;
      RECT 5.0940 17.5365 9.6120 18.3560 ;
      RECT 0.0000 17.6360 5.0760 18.3560 ;
      RECT 4.8690 17.5365 9.6120 17.7080 ;
      RECT 0.0000 17.5365 4.8510 18.3560 ;
      RECT 0.0000 17.5365 9.6120 17.6120 ;
      RECT 0.0000 19.5800 9.6120 19.7100 ;
      RECT 9.4950 18.6165 9.6120 19.7100 ;
      RECT 5.8410 19.4840 9.4770 19.7100 ;
      RECT 4.5090 19.4840 5.8230 19.7100 ;
      RECT 3.7890 18.6165 4.4190 19.7100 ;
      RECT 0.1350 19.4840 3.7710 19.7100 ;
      RECT 0.0000 18.6165 0.1170 19.7100 ;
      RECT 9.4590 18.6165 9.6120 19.5320 ;
      RECT 5.8950 18.6165 9.4410 19.7100 ;
      RECT 5.1480 18.6165 5.8770 19.5320 ;
      RECT 4.9860 18.8120 5.1120 19.7100 ;
      RECT 3.7350 18.7160 4.9590 19.5320 ;
      RECT 0.1710 18.6165 3.7170 19.7100 ;
      RECT 0.0000 18.6165 0.1530 19.5320 ;
      RECT 5.0940 18.6165 9.6120 19.4360 ;
      RECT 0.0000 18.7160 5.0760 19.4360 ;
      RECT 4.8690 18.6165 9.6120 18.7880 ;
      RECT 0.0000 18.6165 4.8510 19.4360 ;
      RECT 0.0000 18.6165 9.6120 18.6920 ;
      RECT 0.0000 20.6600 9.6120 20.7900 ;
      RECT 9.4950 19.6965 9.6120 20.7900 ;
      RECT 5.8410 20.5640 9.4770 20.7900 ;
      RECT 4.5090 20.5640 5.8230 20.7900 ;
      RECT 3.7890 19.6965 4.4190 20.7900 ;
      RECT 0.1350 20.5640 3.7710 20.7900 ;
      RECT 0.0000 19.6965 0.1170 20.7900 ;
      RECT 9.4590 19.6965 9.6120 20.6120 ;
      RECT 5.8950 19.6965 9.4410 20.7900 ;
      RECT 5.1480 19.6965 5.8770 20.6120 ;
      RECT 4.9860 19.8920 5.1120 20.7900 ;
      RECT 3.7350 19.7960 4.9590 20.6120 ;
      RECT 0.1710 19.6965 3.7170 20.7900 ;
      RECT 0.0000 19.6965 0.1530 20.6120 ;
      RECT 5.0940 19.6965 9.6120 20.5160 ;
      RECT 0.0000 19.7960 5.0760 20.5160 ;
      RECT 4.8690 19.6965 9.6120 19.8680 ;
      RECT 0.0000 19.6965 4.8510 20.5160 ;
      RECT 0.0000 19.6965 9.6120 19.7720 ;
      RECT 0.0000 21.7400 9.6120 21.8700 ;
      RECT 9.4950 20.7765 9.6120 21.8700 ;
      RECT 5.8410 21.6440 9.4770 21.8700 ;
      RECT 4.5090 21.6440 5.8230 21.8700 ;
      RECT 3.7890 20.7765 4.4190 21.8700 ;
      RECT 0.1350 21.6440 3.7710 21.8700 ;
      RECT 0.0000 20.7765 0.1170 21.8700 ;
      RECT 9.4590 20.7765 9.6120 21.6920 ;
      RECT 5.8950 20.7765 9.4410 21.8700 ;
      RECT 5.1480 20.7765 5.8770 21.6920 ;
      RECT 4.9860 20.9720 5.1120 21.8700 ;
      RECT 3.7350 20.8760 4.9590 21.6920 ;
      RECT 0.1710 20.7765 3.7170 21.8700 ;
      RECT 0.0000 20.7765 0.1530 21.6920 ;
      RECT 5.0940 20.7765 9.6120 21.5960 ;
      RECT 0.0000 20.8760 5.0760 21.5960 ;
      RECT 4.8690 20.7765 9.6120 20.9480 ;
      RECT 0.0000 20.7765 4.8510 21.5960 ;
      RECT 0.0000 20.7765 9.6120 20.8520 ;
      RECT 0.0000 22.8200 9.6120 22.9500 ;
      RECT 9.4950 21.8565 9.6120 22.9500 ;
      RECT 5.8410 22.7240 9.4770 22.9500 ;
      RECT 4.5090 22.7240 5.8230 22.9500 ;
      RECT 3.7890 21.8565 4.4190 22.9500 ;
      RECT 0.1350 22.7240 3.7710 22.9500 ;
      RECT 0.0000 21.8565 0.1170 22.9500 ;
      RECT 9.4590 21.8565 9.6120 22.7720 ;
      RECT 5.8950 21.8565 9.4410 22.9500 ;
      RECT 5.1480 21.8565 5.8770 22.7720 ;
      RECT 4.9860 22.0520 5.1120 22.9500 ;
      RECT 3.7350 21.9560 4.9590 22.7720 ;
      RECT 0.1710 21.8565 3.7170 22.9500 ;
      RECT 0.0000 21.8565 0.1530 22.7720 ;
      RECT 5.0940 21.8565 9.6120 22.6760 ;
      RECT 0.0000 21.9560 5.0760 22.6760 ;
      RECT 4.8690 21.8565 9.6120 22.0280 ;
      RECT 0.0000 21.8565 4.8510 22.6760 ;
      RECT 0.0000 21.8565 9.6120 21.9320 ;
      RECT 0.0000 23.9000 9.6120 24.0300 ;
      RECT 9.4950 22.9365 9.6120 24.0300 ;
      RECT 5.8410 23.8040 9.4770 24.0300 ;
      RECT 4.5090 23.8040 5.8230 24.0300 ;
      RECT 3.7890 22.9365 4.4190 24.0300 ;
      RECT 0.1350 23.8040 3.7710 24.0300 ;
      RECT 0.0000 22.9365 0.1170 24.0300 ;
      RECT 9.4590 22.9365 9.6120 23.8520 ;
      RECT 5.8950 22.9365 9.4410 24.0300 ;
      RECT 5.1480 22.9365 5.8770 23.8520 ;
      RECT 4.9860 23.1320 5.1120 24.0300 ;
      RECT 3.7350 23.0360 4.9590 23.8520 ;
      RECT 0.1710 22.9365 3.7170 24.0300 ;
      RECT 0.0000 22.9365 0.1530 23.8520 ;
      RECT 5.0940 22.9365 9.6120 23.7560 ;
      RECT 0.0000 23.0360 5.0760 23.7560 ;
      RECT 4.8690 22.9365 9.6120 23.1080 ;
      RECT 0.0000 22.9365 4.8510 23.7560 ;
      RECT 0.0000 22.9365 9.6120 23.0120 ;
      RECT 0.0000 24.9800 9.6120 25.1100 ;
      RECT 9.4950 24.0165 9.6120 25.1100 ;
      RECT 5.8410 24.8840 9.4770 25.1100 ;
      RECT 4.5090 24.8840 5.8230 25.1100 ;
      RECT 3.7890 24.0165 4.4190 25.1100 ;
      RECT 0.1350 24.8840 3.7710 25.1100 ;
      RECT 0.0000 24.0165 0.1170 25.1100 ;
      RECT 9.4590 24.0165 9.6120 24.9320 ;
      RECT 5.8950 24.0165 9.4410 25.1100 ;
      RECT 5.1480 24.0165 5.8770 24.9320 ;
      RECT 4.9860 24.2120 5.1120 25.1100 ;
      RECT 3.7350 24.1160 4.9590 24.9320 ;
      RECT 0.1710 24.0165 3.7170 25.1100 ;
      RECT 0.0000 24.0165 0.1530 24.9320 ;
      RECT 5.0940 24.0165 9.6120 24.8360 ;
      RECT 0.0000 24.1160 5.0760 24.8360 ;
      RECT 4.8690 24.0165 9.6120 24.1880 ;
      RECT 0.0000 24.0165 4.8510 24.8360 ;
      RECT 0.0000 24.0165 9.6120 24.0920 ;
      RECT 0.0000 26.0600 9.6120 26.1900 ;
      RECT 9.4950 25.0965 9.6120 26.1900 ;
      RECT 5.8410 25.9640 9.4770 26.1900 ;
      RECT 4.5090 25.9640 5.8230 26.1900 ;
      RECT 3.7890 25.0965 4.4190 26.1900 ;
      RECT 0.1350 25.9640 3.7710 26.1900 ;
      RECT 0.0000 25.0965 0.1170 26.1900 ;
      RECT 9.4590 25.0965 9.6120 26.0120 ;
      RECT 5.8950 25.0965 9.4410 26.1900 ;
      RECT 5.1480 25.0965 5.8770 26.0120 ;
      RECT 4.9860 25.2920 5.1120 26.1900 ;
      RECT 3.7350 25.1960 4.9590 26.0120 ;
      RECT 0.1710 25.0965 3.7170 26.1900 ;
      RECT 0.0000 25.0965 0.1530 26.0120 ;
      RECT 5.0940 25.0965 9.6120 25.9160 ;
      RECT 0.0000 25.1960 5.0760 25.9160 ;
      RECT 4.8690 25.0965 9.6120 25.2680 ;
      RECT 0.0000 25.0965 4.8510 25.9160 ;
      RECT 0.0000 25.0965 9.6120 25.1720 ;
      RECT 0.0000 27.1400 9.6120 27.2700 ;
      RECT 9.4950 26.1765 9.6120 27.2700 ;
      RECT 5.8410 27.0440 9.4770 27.2700 ;
      RECT 4.5090 27.0440 5.8230 27.2700 ;
      RECT 3.7890 26.1765 4.4190 27.2700 ;
      RECT 0.1350 27.0440 3.7710 27.2700 ;
      RECT 0.0000 26.1765 0.1170 27.2700 ;
      RECT 9.4590 26.1765 9.6120 27.0920 ;
      RECT 5.8950 26.1765 9.4410 27.2700 ;
      RECT 5.1480 26.1765 5.8770 27.0920 ;
      RECT 4.9860 26.3720 5.1120 27.2700 ;
      RECT 3.7350 26.2760 4.9590 27.0920 ;
      RECT 0.1710 26.1765 3.7170 27.2700 ;
      RECT 0.0000 26.1765 0.1530 27.0920 ;
      RECT 5.0940 26.1765 9.6120 26.9960 ;
      RECT 0.0000 26.2760 5.0760 26.9960 ;
      RECT 4.8690 26.1765 9.6120 26.3480 ;
      RECT 0.0000 26.1765 4.8510 26.9960 ;
      RECT 0.0000 26.1765 9.6120 26.2520 ;
      RECT 0.0000 28.2200 9.6120 28.3500 ;
      RECT 9.4950 27.2565 9.6120 28.3500 ;
      RECT 5.8410 28.1240 9.4770 28.3500 ;
      RECT 4.5090 28.1240 5.8230 28.3500 ;
      RECT 3.7890 27.2565 4.4190 28.3500 ;
      RECT 0.1350 28.1240 3.7710 28.3500 ;
      RECT 0.0000 27.2565 0.1170 28.3500 ;
      RECT 9.4590 27.2565 9.6120 28.1720 ;
      RECT 5.8950 27.2565 9.4410 28.3500 ;
      RECT 5.1480 27.2565 5.8770 28.1720 ;
      RECT 4.9860 27.4520 5.1120 28.3500 ;
      RECT 3.7350 27.3560 4.9590 28.1720 ;
      RECT 0.1710 27.2565 3.7170 28.3500 ;
      RECT 0.0000 27.2565 0.1530 28.1720 ;
      RECT 5.0940 27.2565 9.6120 28.0760 ;
      RECT 0.0000 27.3560 5.0760 28.0760 ;
      RECT 4.8690 27.2565 9.6120 27.4280 ;
      RECT 0.0000 27.2565 4.8510 28.0760 ;
      RECT 0.0000 27.2565 9.6120 27.3320 ;
      RECT 0.0000 29.3000 9.6120 29.4300 ;
      RECT 9.4950 28.3365 9.6120 29.4300 ;
      RECT 5.8410 29.2040 9.4770 29.4300 ;
      RECT 4.5090 29.2040 5.8230 29.4300 ;
      RECT 3.7890 28.3365 4.4190 29.4300 ;
      RECT 0.1350 29.2040 3.7710 29.4300 ;
      RECT 0.0000 28.3365 0.1170 29.4300 ;
      RECT 9.4590 28.3365 9.6120 29.2520 ;
      RECT 5.8950 28.3365 9.4410 29.4300 ;
      RECT 5.1480 28.3365 5.8770 29.2520 ;
      RECT 4.9860 28.5320 5.1120 29.4300 ;
      RECT 3.7350 28.4360 4.9590 29.2520 ;
      RECT 0.1710 28.3365 3.7170 29.4300 ;
      RECT 0.0000 28.3365 0.1530 29.2520 ;
      RECT 5.0940 28.3365 9.6120 29.1560 ;
      RECT 0.0000 28.4360 5.0760 29.1560 ;
      RECT 4.8690 28.3365 9.6120 28.5080 ;
      RECT 0.0000 28.3365 4.8510 29.1560 ;
      RECT 0.0000 28.3365 9.6120 28.4120 ;
      RECT 0.0000 30.3800 9.6120 30.5100 ;
      RECT 9.4950 29.4165 9.6120 30.5100 ;
      RECT 5.8410 30.2840 9.4770 30.5100 ;
      RECT 4.5090 30.2840 5.8230 30.5100 ;
      RECT 3.7890 29.4165 4.4190 30.5100 ;
      RECT 0.1350 30.2840 3.7710 30.5100 ;
      RECT 0.0000 29.4165 0.1170 30.5100 ;
      RECT 9.4590 29.4165 9.6120 30.3320 ;
      RECT 5.8950 29.4165 9.4410 30.5100 ;
      RECT 5.1480 29.4165 5.8770 30.3320 ;
      RECT 4.9860 29.6120 5.1120 30.5100 ;
      RECT 3.7350 29.5160 4.9590 30.3320 ;
      RECT 0.1710 29.4165 3.7170 30.5100 ;
      RECT 0.0000 29.4165 0.1530 30.3320 ;
      RECT 5.0940 29.4165 9.6120 30.2360 ;
      RECT 0.0000 29.5160 5.0760 30.2360 ;
      RECT 4.8690 29.4165 9.6120 29.5880 ;
      RECT 0.0000 29.4165 4.8510 30.2360 ;
      RECT 0.0000 29.4165 9.6120 29.4920 ;
      RECT 0.0000 31.4600 9.6120 31.5900 ;
      RECT 9.4950 30.4965 9.6120 31.5900 ;
      RECT 5.8410 31.3640 9.4770 31.5900 ;
      RECT 4.5090 31.3640 5.8230 31.5900 ;
      RECT 3.7890 30.4965 4.4190 31.5900 ;
      RECT 0.1350 31.3640 3.7710 31.5900 ;
      RECT 0.0000 30.4965 0.1170 31.5900 ;
      RECT 9.4590 30.4965 9.6120 31.4120 ;
      RECT 5.8950 30.4965 9.4410 31.5900 ;
      RECT 5.1480 30.4965 5.8770 31.4120 ;
      RECT 4.9860 30.6920 5.1120 31.5900 ;
      RECT 3.7350 30.5960 4.9590 31.4120 ;
      RECT 0.1710 30.4965 3.7170 31.5900 ;
      RECT 0.0000 30.4965 0.1530 31.4120 ;
      RECT 5.0940 30.4965 9.6120 31.3160 ;
      RECT 0.0000 30.5960 5.0760 31.3160 ;
      RECT 4.8690 30.4965 9.6120 30.6680 ;
      RECT 0.0000 30.4965 4.8510 31.3160 ;
      RECT 0.0000 30.4965 9.6120 30.5720 ;
      RECT 0.0000 32.5400 9.6120 32.6700 ;
      RECT 9.4950 31.5765 9.6120 32.6700 ;
      RECT 5.8410 32.4440 9.4770 32.6700 ;
      RECT 4.5090 32.4440 5.8230 32.6700 ;
      RECT 3.7890 31.5765 4.4190 32.6700 ;
      RECT 0.1350 32.4440 3.7710 32.6700 ;
      RECT 0.0000 31.5765 0.1170 32.6700 ;
      RECT 9.4590 31.5765 9.6120 32.4920 ;
      RECT 5.8950 31.5765 9.4410 32.6700 ;
      RECT 5.1480 31.5765 5.8770 32.4920 ;
      RECT 4.9860 31.7720 5.1120 32.6700 ;
      RECT 3.7350 31.6760 4.9590 32.4920 ;
      RECT 0.1710 31.5765 3.7170 32.6700 ;
      RECT 0.0000 31.5765 0.1530 32.4920 ;
      RECT 5.0940 31.5765 9.6120 32.3960 ;
      RECT 0.0000 31.6760 5.0760 32.3960 ;
      RECT 4.8690 31.5765 9.6120 31.7480 ;
      RECT 0.0000 31.5765 4.8510 32.3960 ;
      RECT 0.0000 31.5765 9.6120 31.6520 ;
      RECT 0.0000 33.6200 9.6120 33.7500 ;
      RECT 9.4950 32.6565 9.6120 33.7500 ;
      RECT 5.8410 33.5240 9.4770 33.7500 ;
      RECT 4.5090 33.5240 5.8230 33.7500 ;
      RECT 3.7890 32.6565 4.4190 33.7500 ;
      RECT 0.1350 33.5240 3.7710 33.7500 ;
      RECT 0.0000 32.6565 0.1170 33.7500 ;
      RECT 9.4590 32.6565 9.6120 33.5720 ;
      RECT 5.8950 32.6565 9.4410 33.7500 ;
      RECT 5.1480 32.6565 5.8770 33.5720 ;
      RECT 4.9860 32.8520 5.1120 33.7500 ;
      RECT 3.7350 32.7560 4.9590 33.5720 ;
      RECT 0.1710 32.6565 3.7170 33.7500 ;
      RECT 0.0000 32.6565 0.1530 33.5720 ;
      RECT 5.0940 32.6565 9.6120 33.4760 ;
      RECT 0.0000 32.7560 5.0760 33.4760 ;
      RECT 4.8690 32.6565 9.6120 32.8280 ;
      RECT 0.0000 32.6565 4.8510 33.4760 ;
      RECT 0.0000 32.6565 9.6120 32.7320 ;
      RECT 0.0000 34.7000 9.6120 34.8300 ;
      RECT 9.4950 33.7365 9.6120 34.8300 ;
      RECT 5.8410 34.6040 9.4770 34.8300 ;
      RECT 4.5090 34.6040 5.8230 34.8300 ;
      RECT 3.7890 33.7365 4.4190 34.8300 ;
      RECT 0.1350 34.6040 3.7710 34.8300 ;
      RECT 0.0000 33.7365 0.1170 34.8300 ;
      RECT 9.4590 33.7365 9.6120 34.6520 ;
      RECT 5.8950 33.7365 9.4410 34.8300 ;
      RECT 5.1480 33.7365 5.8770 34.6520 ;
      RECT 4.9860 33.9320 5.1120 34.8300 ;
      RECT 3.7350 33.8360 4.9590 34.6520 ;
      RECT 0.1710 33.7365 3.7170 34.8300 ;
      RECT 0.0000 33.7365 0.1530 34.6520 ;
      RECT 5.0940 33.7365 9.6120 34.5560 ;
      RECT 0.0000 33.8360 5.0760 34.5560 ;
      RECT 4.8690 33.7365 9.6120 33.9080 ;
      RECT 0.0000 33.7365 4.8510 34.5560 ;
      RECT 0.0000 33.7365 9.6120 33.8120 ;
      RECT 0.0000 35.7800 9.6120 35.9100 ;
      RECT 9.4950 34.8165 9.6120 35.9100 ;
      RECT 5.8410 35.6840 9.4770 35.9100 ;
      RECT 4.5090 35.6840 5.8230 35.9100 ;
      RECT 3.7890 34.8165 4.4190 35.9100 ;
      RECT 0.1350 35.6840 3.7710 35.9100 ;
      RECT 0.0000 34.8165 0.1170 35.9100 ;
      RECT 9.4590 34.8165 9.6120 35.7320 ;
      RECT 5.8950 34.8165 9.4410 35.9100 ;
      RECT 5.1480 34.8165 5.8770 35.7320 ;
      RECT 4.9860 35.0120 5.1120 35.9100 ;
      RECT 3.7350 34.9160 4.9590 35.7320 ;
      RECT 0.1710 34.8165 3.7170 35.9100 ;
      RECT 0.0000 34.8165 0.1530 35.7320 ;
      RECT 5.0940 34.8165 9.6120 35.6360 ;
      RECT 0.0000 34.9160 5.0760 35.6360 ;
      RECT 4.8690 34.8165 9.6120 34.9880 ;
      RECT 0.0000 34.8165 4.8510 35.6360 ;
      RECT 0.0000 34.8165 9.6120 34.8920 ;
      RECT 0.0000 36.8600 9.6120 36.9900 ;
      RECT 9.4950 35.8965 9.6120 36.9900 ;
      RECT 5.8410 36.7640 9.4770 36.9900 ;
      RECT 4.5090 36.7640 5.8230 36.9900 ;
      RECT 3.7890 35.8965 4.4190 36.9900 ;
      RECT 0.1350 36.7640 3.7710 36.9900 ;
      RECT 0.0000 35.8965 0.1170 36.9900 ;
      RECT 9.4590 35.8965 9.6120 36.8120 ;
      RECT 5.8950 35.8965 9.4410 36.9900 ;
      RECT 5.1480 35.8965 5.8770 36.8120 ;
      RECT 4.9860 36.0920 5.1120 36.9900 ;
      RECT 3.7350 35.9960 4.9590 36.8120 ;
      RECT 0.1710 35.8965 3.7170 36.9900 ;
      RECT 0.0000 35.8965 0.1530 36.8120 ;
      RECT 5.0940 35.8965 9.6120 36.7160 ;
      RECT 0.0000 35.9960 5.0760 36.7160 ;
      RECT 4.8690 35.8965 9.6120 36.0680 ;
      RECT 0.0000 35.8965 4.8510 36.7160 ;
      RECT 0.0000 35.8965 9.6120 35.9720 ;
      RECT 0.0000 37.9400 9.6120 38.0700 ;
      RECT 9.4950 36.9765 9.6120 38.0700 ;
      RECT 5.8410 37.8440 9.4770 38.0700 ;
      RECT 4.5090 37.8440 5.8230 38.0700 ;
      RECT 3.7890 36.9765 4.4190 38.0700 ;
      RECT 0.1350 37.8440 3.7710 38.0700 ;
      RECT 0.0000 36.9765 0.1170 38.0700 ;
      RECT 9.4590 36.9765 9.6120 37.8920 ;
      RECT 5.8950 36.9765 9.4410 38.0700 ;
      RECT 5.1480 36.9765 5.8770 37.8920 ;
      RECT 4.9860 37.1720 5.1120 38.0700 ;
      RECT 3.7350 37.0760 4.9590 37.8920 ;
      RECT 0.1710 36.9765 3.7170 38.0700 ;
      RECT 0.0000 36.9765 0.1530 37.8920 ;
      RECT 5.0940 36.9765 9.6120 37.7960 ;
      RECT 0.0000 37.0760 5.0760 37.7960 ;
      RECT 4.8690 36.9765 9.6120 37.1480 ;
      RECT 0.0000 36.9765 4.8510 37.7960 ;
      RECT 0.0000 36.9765 9.6120 37.0520 ;
      RECT 0.0000 39.0200 9.6120 39.1500 ;
      RECT 9.4950 38.0565 9.6120 39.1500 ;
      RECT 5.8410 38.9240 9.4770 39.1500 ;
      RECT 4.5090 38.9240 5.8230 39.1500 ;
      RECT 3.7890 38.0565 4.4190 39.1500 ;
      RECT 0.1350 38.9240 3.7710 39.1500 ;
      RECT 0.0000 38.0565 0.1170 39.1500 ;
      RECT 9.4590 38.0565 9.6120 38.9720 ;
      RECT 5.8950 38.0565 9.4410 39.1500 ;
      RECT 5.1480 38.0565 5.8770 38.9720 ;
      RECT 4.9860 38.2520 5.1120 39.1500 ;
      RECT 3.7350 38.1560 4.9590 38.9720 ;
      RECT 0.1710 38.0565 3.7170 39.1500 ;
      RECT 0.0000 38.0565 0.1530 38.9720 ;
      RECT 5.0940 38.0565 9.6120 38.8760 ;
      RECT 0.0000 38.1560 5.0760 38.8760 ;
      RECT 4.8690 38.0565 9.6120 38.2280 ;
      RECT 0.0000 38.0565 4.8510 38.8760 ;
      RECT 0.0000 38.0565 9.6120 38.1320 ;
      RECT 0.0000 40.1000 9.6120 40.2300 ;
      RECT 9.4950 39.1365 9.6120 40.2300 ;
      RECT 5.8410 40.0040 9.4770 40.2300 ;
      RECT 4.5090 40.0040 5.8230 40.2300 ;
      RECT 3.7890 39.1365 4.4190 40.2300 ;
      RECT 0.1350 40.0040 3.7710 40.2300 ;
      RECT 0.0000 39.1365 0.1170 40.2300 ;
      RECT 9.4590 39.1365 9.6120 40.0520 ;
      RECT 5.8950 39.1365 9.4410 40.2300 ;
      RECT 5.1480 39.1365 5.8770 40.0520 ;
      RECT 4.9860 39.3320 5.1120 40.2300 ;
      RECT 3.7350 39.2360 4.9590 40.0520 ;
      RECT 0.1710 39.1365 3.7170 40.2300 ;
      RECT 0.0000 39.1365 0.1530 40.0520 ;
      RECT 5.0940 39.1365 9.6120 39.9560 ;
      RECT 0.0000 39.2360 5.0760 39.9560 ;
      RECT 4.8690 39.1365 9.6120 39.3080 ;
      RECT 0.0000 39.1365 4.8510 39.9560 ;
      RECT 0.0000 39.1365 9.6120 39.2120 ;
      RECT 0.0000 41.1800 9.6120 41.3100 ;
      RECT 9.4950 40.2165 9.6120 41.3100 ;
      RECT 5.8410 41.0840 9.4770 41.3100 ;
      RECT 4.5090 41.0840 5.8230 41.3100 ;
      RECT 3.7890 40.2165 4.4190 41.3100 ;
      RECT 0.1350 41.0840 3.7710 41.3100 ;
      RECT 0.0000 40.2165 0.1170 41.3100 ;
      RECT 9.4590 40.2165 9.6120 41.1320 ;
      RECT 5.8950 40.2165 9.4410 41.3100 ;
      RECT 5.1480 40.2165 5.8770 41.1320 ;
      RECT 4.9860 40.4120 5.1120 41.3100 ;
      RECT 3.7350 40.3160 4.9590 41.1320 ;
      RECT 0.1710 40.2165 3.7170 41.3100 ;
      RECT 0.0000 40.2165 0.1530 41.1320 ;
      RECT 5.0940 40.2165 9.6120 41.0360 ;
      RECT 0.0000 40.3160 5.0760 41.0360 ;
      RECT 4.8690 40.2165 9.6120 40.3880 ;
      RECT 0.0000 40.2165 4.8510 41.0360 ;
      RECT 0.0000 40.2165 9.6120 40.2920 ;
      RECT 0.0000 42.2600 9.6120 42.3900 ;
      RECT 9.4950 41.2965 9.6120 42.3900 ;
      RECT 5.8410 42.1640 9.4770 42.3900 ;
      RECT 4.5090 42.1640 5.8230 42.3900 ;
      RECT 3.7890 41.2965 4.4190 42.3900 ;
      RECT 0.1350 42.1640 3.7710 42.3900 ;
      RECT 0.0000 41.2965 0.1170 42.3900 ;
      RECT 9.4590 41.2965 9.6120 42.2120 ;
      RECT 5.8950 41.2965 9.4410 42.3900 ;
      RECT 5.1480 41.2965 5.8770 42.2120 ;
      RECT 4.9860 41.4920 5.1120 42.3900 ;
      RECT 3.7350 41.3960 4.9590 42.2120 ;
      RECT 0.1710 41.2965 3.7170 42.3900 ;
      RECT 0.0000 41.2965 0.1530 42.2120 ;
      RECT 5.0940 41.2965 9.6120 42.1160 ;
      RECT 0.0000 41.3960 5.0760 42.1160 ;
      RECT 4.8690 41.2965 9.6120 41.4680 ;
      RECT 0.0000 41.2965 4.8510 42.1160 ;
      RECT 0.0000 41.2965 9.6120 41.3720 ;
      RECT 0.0000 43.3400 9.6120 43.4700 ;
      RECT 9.4950 42.3765 9.6120 43.4700 ;
      RECT 5.8410 43.2440 9.4770 43.4700 ;
      RECT 4.5090 43.2440 5.8230 43.4700 ;
      RECT 3.7890 42.3765 4.4190 43.4700 ;
      RECT 0.1350 43.2440 3.7710 43.4700 ;
      RECT 0.0000 42.3765 0.1170 43.4700 ;
      RECT 9.4590 42.3765 9.6120 43.2920 ;
      RECT 5.8950 42.3765 9.4410 43.4700 ;
      RECT 5.1480 42.3765 5.8770 43.2920 ;
      RECT 4.9860 42.5720 5.1120 43.4700 ;
      RECT 3.7350 42.4760 4.9590 43.2920 ;
      RECT 0.1710 42.3765 3.7170 43.4700 ;
      RECT 0.0000 42.3765 0.1530 43.2920 ;
      RECT 5.0940 42.3765 9.6120 43.1960 ;
      RECT 0.0000 42.4760 5.0760 43.1960 ;
      RECT 4.8690 42.3765 9.6120 42.5480 ;
      RECT 0.0000 42.3765 4.8510 43.1960 ;
      RECT 0.0000 42.3765 9.6120 42.4520 ;
      RECT 0.0000 50.7630 9.6120 52.0965 ;
      RECT 7.3530 43.4430 9.6120 52.0965 ;
      RECT 5.1530 47.3070 9.6120 52.0965 ;
      RECT 6.0570 44.7150 9.6120 52.0965 ;
      RECT 5.1010 43.4430 5.1350 52.0965 ;
      RECT 5.0490 43.4430 5.0830 52.0965 ;
      RECT 4.9970 43.4430 5.0310 52.0965 ;
      RECT 4.9450 43.4430 4.9790 52.0965 ;
      RECT 0.0000 50.3310 4.9270 52.0965 ;
      RECT 4.6850 47.5950 9.6120 50.5470 ;
      RECT 4.6330 43.4430 4.6670 52.0965 ;
      RECT 4.5810 43.4430 4.6150 52.0965 ;
      RECT 4.5290 43.4430 4.5630 52.0965 ;
      RECT 4.4770 43.4430 4.5110 52.0965 ;
      RECT 0.0000 45.0030 4.4590 52.0965 ;
      RECT 0.0000 47.1630 4.9270 50.1150 ;
      RECT 4.6850 44.4270 5.8230 47.3790 ;
      RECT 5.8410 44.9070 9.6120 52.0965 ;
      RECT 5.1930 43.5230 6.0390 47.2830 ;
      RECT 4.0050 43.9950 4.7790 46.9470 ;
      RECT 3.7890 44.1390 4.4590 52.0965 ;
      RECT 0.0000 44.7150 3.7710 52.0965 ;
      RECT 3.3570 43.4430 3.8070 44.9790 ;
      RECT 7.1370 43.4430 7.3350 52.0965 ;
      RECT 3.3570 44.5230 7.1190 44.8830 ;
      RECT 2.4930 44.1390 3.3390 52.0965 ;
      RECT 0.0000 44.4270 2.4750 52.0965 ;
      RECT 6.9210 43.4430 9.6120 44.6910 ;
      RECT 6.7050 44.1390 9.6120 44.6910 ;
      RECT 0.0000 44.4270 6.6870 44.6910 ;
      RECT 6.4890 43.4430 6.9030 44.4990 ;
      RECT 5.1530 44.1390 9.6120 44.4990 ;
      RECT 0.1710 44.1390 4.9270 44.6910 ;
      RECT 4.6850 44.0910 4.9270 52.0965 ;
      RECT 0.0000 43.9950 0.1530 52.0965 ;
      RECT 4.7970 43.4430 5.1750 44.2110 ;
      RECT 5.1930 44.0910 6.4710 44.8830 ;
      RECT 3.1410 44.0910 3.9870 44.6910 ;
      RECT 2.7090 44.0910 3.1230 52.0965 ;
      RECT 0.0000 43.9950 2.6910 44.2110 ;
      RECT 6.2730 43.4430 9.6120 44.1150 ;
      RECT 4.7970 43.5230 6.2550 44.1150 ;
      RECT 3.8250 43.9950 4.7790 44.1150 ;
      RECT 2.9250 43.4430 3.8070 44.1150 ;
      RECT 0.0000 43.9950 2.9070 44.1150 ;
      RECT 5.8410 43.4430 9.6120 44.0670 ;
      RECT 4.6850 43.5230 9.6120 44.0670 ;
      RECT 0.1350 43.4430 4.4590 44.0670 ;
      RECT 0.0000 43.4430 0.1170 52.0965 ;
      RECT 0.0000 43.4430 5.8230 43.7790 ;
      RECT 0.0000 43.4430 9.6120 43.4990 ;
        RECT 0.0000 52.5470 9.6120 52.6770 ;
        RECT 9.4950 51.5835 9.6120 52.6770 ;
        RECT 5.8410 52.4510 9.4770 52.6770 ;
        RECT 4.5090 52.4510 5.8230 52.6770 ;
        RECT 3.7890 51.5835 4.4190 52.6770 ;
        RECT 0.1350 52.4510 3.7710 52.6770 ;
        RECT 0.0000 51.5835 0.1170 52.6770 ;
        RECT 9.4590 51.5835 9.6120 52.4990 ;
        RECT 5.8950 51.5835 9.4410 52.6770 ;
        RECT 5.1480 51.5835 5.8770 52.4990 ;
        RECT 4.9860 51.7790 5.1120 52.6770 ;
        RECT 3.7350 51.6830 4.9590 52.4990 ;
        RECT 0.1710 51.5835 3.7170 52.6770 ;
        RECT 0.0000 51.5835 0.1530 52.4990 ;
        RECT 5.0940 51.5835 9.6120 52.4030 ;
        RECT 0.0000 51.6830 5.0760 52.4030 ;
        RECT 4.8690 51.5835 9.6120 51.7550 ;
        RECT 0.0000 51.5835 4.8510 52.4030 ;
        RECT 0.0000 51.5835 9.6120 51.6590 ;
        RECT 0.0000 53.6270 9.6120 53.7570 ;
        RECT 9.4950 52.6635 9.6120 53.7570 ;
        RECT 5.8410 53.5310 9.4770 53.7570 ;
        RECT 4.5090 53.5310 5.8230 53.7570 ;
        RECT 3.7890 52.6635 4.4190 53.7570 ;
        RECT 0.1350 53.5310 3.7710 53.7570 ;
        RECT 0.0000 52.6635 0.1170 53.7570 ;
        RECT 9.4590 52.6635 9.6120 53.5790 ;
        RECT 5.8950 52.6635 9.4410 53.7570 ;
        RECT 5.1480 52.6635 5.8770 53.5790 ;
        RECT 4.9860 52.8590 5.1120 53.7570 ;
        RECT 3.7350 52.7630 4.9590 53.5790 ;
        RECT 0.1710 52.6635 3.7170 53.7570 ;
        RECT 0.0000 52.6635 0.1530 53.5790 ;
        RECT 5.0940 52.6635 9.6120 53.4830 ;
        RECT 0.0000 52.7630 5.0760 53.4830 ;
        RECT 4.8690 52.6635 9.6120 52.8350 ;
        RECT 0.0000 52.6635 4.8510 53.4830 ;
        RECT 0.0000 52.6635 9.6120 52.7390 ;
        RECT 0.0000 54.7070 9.6120 54.8370 ;
        RECT 9.4950 53.7435 9.6120 54.8370 ;
        RECT 5.8410 54.6110 9.4770 54.8370 ;
        RECT 4.5090 54.6110 5.8230 54.8370 ;
        RECT 3.7890 53.7435 4.4190 54.8370 ;
        RECT 0.1350 54.6110 3.7710 54.8370 ;
        RECT 0.0000 53.7435 0.1170 54.8370 ;
        RECT 9.4590 53.7435 9.6120 54.6590 ;
        RECT 5.8950 53.7435 9.4410 54.8370 ;
        RECT 5.1480 53.7435 5.8770 54.6590 ;
        RECT 4.9860 53.9390 5.1120 54.8370 ;
        RECT 3.7350 53.8430 4.9590 54.6590 ;
        RECT 0.1710 53.7435 3.7170 54.8370 ;
        RECT 0.0000 53.7435 0.1530 54.6590 ;
        RECT 5.0940 53.7435 9.6120 54.5630 ;
        RECT 0.0000 53.8430 5.0760 54.5630 ;
        RECT 4.8690 53.7435 9.6120 53.9150 ;
        RECT 0.0000 53.7435 4.8510 54.5630 ;
        RECT 0.0000 53.7435 9.6120 53.8190 ;
        RECT 0.0000 55.7870 9.6120 55.9170 ;
        RECT 9.4950 54.8235 9.6120 55.9170 ;
        RECT 5.8410 55.6910 9.4770 55.9170 ;
        RECT 4.5090 55.6910 5.8230 55.9170 ;
        RECT 3.7890 54.8235 4.4190 55.9170 ;
        RECT 0.1350 55.6910 3.7710 55.9170 ;
        RECT 0.0000 54.8235 0.1170 55.9170 ;
        RECT 9.4590 54.8235 9.6120 55.7390 ;
        RECT 5.8950 54.8235 9.4410 55.9170 ;
        RECT 5.1480 54.8235 5.8770 55.7390 ;
        RECT 4.9860 55.0190 5.1120 55.9170 ;
        RECT 3.7350 54.9230 4.9590 55.7390 ;
        RECT 0.1710 54.8235 3.7170 55.9170 ;
        RECT 0.0000 54.8235 0.1530 55.7390 ;
        RECT 5.0940 54.8235 9.6120 55.6430 ;
        RECT 0.0000 54.9230 5.0760 55.6430 ;
        RECT 4.8690 54.8235 9.6120 54.9950 ;
        RECT 0.0000 54.8235 4.8510 55.6430 ;
        RECT 0.0000 54.8235 9.6120 54.8990 ;
        RECT 0.0000 56.8670 9.6120 56.9970 ;
        RECT 9.4950 55.9035 9.6120 56.9970 ;
        RECT 5.8410 56.7710 9.4770 56.9970 ;
        RECT 4.5090 56.7710 5.8230 56.9970 ;
        RECT 3.7890 55.9035 4.4190 56.9970 ;
        RECT 0.1350 56.7710 3.7710 56.9970 ;
        RECT 0.0000 55.9035 0.1170 56.9970 ;
        RECT 9.4590 55.9035 9.6120 56.8190 ;
        RECT 5.8950 55.9035 9.4410 56.9970 ;
        RECT 5.1480 55.9035 5.8770 56.8190 ;
        RECT 4.9860 56.0990 5.1120 56.9970 ;
        RECT 3.7350 56.0030 4.9590 56.8190 ;
        RECT 0.1710 55.9035 3.7170 56.9970 ;
        RECT 0.0000 55.9035 0.1530 56.8190 ;
        RECT 5.0940 55.9035 9.6120 56.7230 ;
        RECT 0.0000 56.0030 5.0760 56.7230 ;
        RECT 4.8690 55.9035 9.6120 56.0750 ;
        RECT 0.0000 55.9035 4.8510 56.7230 ;
        RECT 0.0000 55.9035 9.6120 55.9790 ;
        RECT 0.0000 57.9470 9.6120 58.0770 ;
        RECT 9.4950 56.9835 9.6120 58.0770 ;
        RECT 5.8410 57.8510 9.4770 58.0770 ;
        RECT 4.5090 57.8510 5.8230 58.0770 ;
        RECT 3.7890 56.9835 4.4190 58.0770 ;
        RECT 0.1350 57.8510 3.7710 58.0770 ;
        RECT 0.0000 56.9835 0.1170 58.0770 ;
        RECT 9.4590 56.9835 9.6120 57.8990 ;
        RECT 5.8950 56.9835 9.4410 58.0770 ;
        RECT 5.1480 56.9835 5.8770 57.8990 ;
        RECT 4.9860 57.1790 5.1120 58.0770 ;
        RECT 3.7350 57.0830 4.9590 57.8990 ;
        RECT 0.1710 56.9835 3.7170 58.0770 ;
        RECT 0.0000 56.9835 0.1530 57.8990 ;
        RECT 5.0940 56.9835 9.6120 57.8030 ;
        RECT 0.0000 57.0830 5.0760 57.8030 ;
        RECT 4.8690 56.9835 9.6120 57.1550 ;
        RECT 0.0000 56.9835 4.8510 57.8030 ;
        RECT 0.0000 56.9835 9.6120 57.0590 ;
        RECT 0.0000 59.0270 9.6120 59.1570 ;
        RECT 9.4950 58.0635 9.6120 59.1570 ;
        RECT 5.8410 58.9310 9.4770 59.1570 ;
        RECT 4.5090 58.9310 5.8230 59.1570 ;
        RECT 3.7890 58.0635 4.4190 59.1570 ;
        RECT 0.1350 58.9310 3.7710 59.1570 ;
        RECT 0.0000 58.0635 0.1170 59.1570 ;
        RECT 9.4590 58.0635 9.6120 58.9790 ;
        RECT 5.8950 58.0635 9.4410 59.1570 ;
        RECT 5.1480 58.0635 5.8770 58.9790 ;
        RECT 4.9860 58.2590 5.1120 59.1570 ;
        RECT 3.7350 58.1630 4.9590 58.9790 ;
        RECT 0.1710 58.0635 3.7170 59.1570 ;
        RECT 0.0000 58.0635 0.1530 58.9790 ;
        RECT 5.0940 58.0635 9.6120 58.8830 ;
        RECT 0.0000 58.1630 5.0760 58.8830 ;
        RECT 4.8690 58.0635 9.6120 58.2350 ;
        RECT 0.0000 58.0635 4.8510 58.8830 ;
        RECT 0.0000 58.0635 9.6120 58.1390 ;
        RECT 0.0000 60.1070 9.6120 60.2370 ;
        RECT 9.4950 59.1435 9.6120 60.2370 ;
        RECT 5.8410 60.0110 9.4770 60.2370 ;
        RECT 4.5090 60.0110 5.8230 60.2370 ;
        RECT 3.7890 59.1435 4.4190 60.2370 ;
        RECT 0.1350 60.0110 3.7710 60.2370 ;
        RECT 0.0000 59.1435 0.1170 60.2370 ;
        RECT 9.4590 59.1435 9.6120 60.0590 ;
        RECT 5.8950 59.1435 9.4410 60.2370 ;
        RECT 5.1480 59.1435 5.8770 60.0590 ;
        RECT 4.9860 59.3390 5.1120 60.2370 ;
        RECT 3.7350 59.2430 4.9590 60.0590 ;
        RECT 0.1710 59.1435 3.7170 60.2370 ;
        RECT 0.0000 59.1435 0.1530 60.0590 ;
        RECT 5.0940 59.1435 9.6120 59.9630 ;
        RECT 0.0000 59.2430 5.0760 59.9630 ;
        RECT 4.8690 59.1435 9.6120 59.3150 ;
        RECT 0.0000 59.1435 4.8510 59.9630 ;
        RECT 0.0000 59.1435 9.6120 59.2190 ;
        RECT 0.0000 61.1870 9.6120 61.3170 ;
        RECT 9.4950 60.2235 9.6120 61.3170 ;
        RECT 5.8410 61.0910 9.4770 61.3170 ;
        RECT 4.5090 61.0910 5.8230 61.3170 ;
        RECT 3.7890 60.2235 4.4190 61.3170 ;
        RECT 0.1350 61.0910 3.7710 61.3170 ;
        RECT 0.0000 60.2235 0.1170 61.3170 ;
        RECT 9.4590 60.2235 9.6120 61.1390 ;
        RECT 5.8950 60.2235 9.4410 61.3170 ;
        RECT 5.1480 60.2235 5.8770 61.1390 ;
        RECT 4.9860 60.4190 5.1120 61.3170 ;
        RECT 3.7350 60.3230 4.9590 61.1390 ;
        RECT 0.1710 60.2235 3.7170 61.3170 ;
        RECT 0.0000 60.2235 0.1530 61.1390 ;
        RECT 5.0940 60.2235 9.6120 61.0430 ;
        RECT 0.0000 60.3230 5.0760 61.0430 ;
        RECT 4.8690 60.2235 9.6120 60.3950 ;
        RECT 0.0000 60.2235 4.8510 61.0430 ;
        RECT 0.0000 60.2235 9.6120 60.2990 ;
        RECT 0.0000 62.2670 9.6120 62.3970 ;
        RECT 9.4950 61.3035 9.6120 62.3970 ;
        RECT 5.8410 62.1710 9.4770 62.3970 ;
        RECT 4.5090 62.1710 5.8230 62.3970 ;
        RECT 3.7890 61.3035 4.4190 62.3970 ;
        RECT 0.1350 62.1710 3.7710 62.3970 ;
        RECT 0.0000 61.3035 0.1170 62.3970 ;
        RECT 9.4590 61.3035 9.6120 62.2190 ;
        RECT 5.8950 61.3035 9.4410 62.3970 ;
        RECT 5.1480 61.3035 5.8770 62.2190 ;
        RECT 4.9860 61.4990 5.1120 62.3970 ;
        RECT 3.7350 61.4030 4.9590 62.2190 ;
        RECT 0.1710 61.3035 3.7170 62.3970 ;
        RECT 0.0000 61.3035 0.1530 62.2190 ;
        RECT 5.0940 61.3035 9.6120 62.1230 ;
        RECT 0.0000 61.4030 5.0760 62.1230 ;
        RECT 4.8690 61.3035 9.6120 61.4750 ;
        RECT 0.0000 61.3035 4.8510 62.1230 ;
        RECT 0.0000 61.3035 9.6120 61.3790 ;
        RECT 0.0000 63.3470 9.6120 63.4770 ;
        RECT 9.4950 62.3835 9.6120 63.4770 ;
        RECT 5.8410 63.2510 9.4770 63.4770 ;
        RECT 4.5090 63.2510 5.8230 63.4770 ;
        RECT 3.7890 62.3835 4.4190 63.4770 ;
        RECT 0.1350 63.2510 3.7710 63.4770 ;
        RECT 0.0000 62.3835 0.1170 63.4770 ;
        RECT 9.4590 62.3835 9.6120 63.2990 ;
        RECT 5.8950 62.3835 9.4410 63.4770 ;
        RECT 5.1480 62.3835 5.8770 63.2990 ;
        RECT 4.9860 62.5790 5.1120 63.4770 ;
        RECT 3.7350 62.4830 4.9590 63.2990 ;
        RECT 0.1710 62.3835 3.7170 63.4770 ;
        RECT 0.0000 62.3835 0.1530 63.2990 ;
        RECT 5.0940 62.3835 9.6120 63.2030 ;
        RECT 0.0000 62.4830 5.0760 63.2030 ;
        RECT 4.8690 62.3835 9.6120 62.5550 ;
        RECT 0.0000 62.3835 4.8510 63.2030 ;
        RECT 0.0000 62.3835 9.6120 62.4590 ;
        RECT 0.0000 64.4270 9.6120 64.5570 ;
        RECT 9.4950 63.4635 9.6120 64.5570 ;
        RECT 5.8410 64.3310 9.4770 64.5570 ;
        RECT 4.5090 64.3310 5.8230 64.5570 ;
        RECT 3.7890 63.4635 4.4190 64.5570 ;
        RECT 0.1350 64.3310 3.7710 64.5570 ;
        RECT 0.0000 63.4635 0.1170 64.5570 ;
        RECT 9.4590 63.4635 9.6120 64.3790 ;
        RECT 5.8950 63.4635 9.4410 64.5570 ;
        RECT 5.1480 63.4635 5.8770 64.3790 ;
        RECT 4.9860 63.6590 5.1120 64.5570 ;
        RECT 3.7350 63.5630 4.9590 64.3790 ;
        RECT 0.1710 63.4635 3.7170 64.5570 ;
        RECT 0.0000 63.4635 0.1530 64.3790 ;
        RECT 5.0940 63.4635 9.6120 64.2830 ;
        RECT 0.0000 63.5630 5.0760 64.2830 ;
        RECT 4.8690 63.4635 9.6120 63.6350 ;
        RECT 0.0000 63.4635 4.8510 64.2830 ;
        RECT 0.0000 63.4635 9.6120 63.5390 ;
        RECT 0.0000 65.5070 9.6120 65.6370 ;
        RECT 9.4950 64.5435 9.6120 65.6370 ;
        RECT 5.8410 65.4110 9.4770 65.6370 ;
        RECT 4.5090 65.4110 5.8230 65.6370 ;
        RECT 3.7890 64.5435 4.4190 65.6370 ;
        RECT 0.1350 65.4110 3.7710 65.6370 ;
        RECT 0.0000 64.5435 0.1170 65.6370 ;
        RECT 9.4590 64.5435 9.6120 65.4590 ;
        RECT 5.8950 64.5435 9.4410 65.6370 ;
        RECT 5.1480 64.5435 5.8770 65.4590 ;
        RECT 4.9860 64.7390 5.1120 65.6370 ;
        RECT 3.7350 64.6430 4.9590 65.4590 ;
        RECT 0.1710 64.5435 3.7170 65.6370 ;
        RECT 0.0000 64.5435 0.1530 65.4590 ;
        RECT 5.0940 64.5435 9.6120 65.3630 ;
        RECT 0.0000 64.6430 5.0760 65.3630 ;
        RECT 4.8690 64.5435 9.6120 64.7150 ;
        RECT 0.0000 64.5435 4.8510 65.3630 ;
        RECT 0.0000 64.5435 9.6120 64.6190 ;
        RECT 0.0000 66.5870 9.6120 66.7170 ;
        RECT 9.4950 65.6235 9.6120 66.7170 ;
        RECT 5.8410 66.4910 9.4770 66.7170 ;
        RECT 4.5090 66.4910 5.8230 66.7170 ;
        RECT 3.7890 65.6235 4.4190 66.7170 ;
        RECT 0.1350 66.4910 3.7710 66.7170 ;
        RECT 0.0000 65.6235 0.1170 66.7170 ;
        RECT 9.4590 65.6235 9.6120 66.5390 ;
        RECT 5.8950 65.6235 9.4410 66.7170 ;
        RECT 5.1480 65.6235 5.8770 66.5390 ;
        RECT 4.9860 65.8190 5.1120 66.7170 ;
        RECT 3.7350 65.7230 4.9590 66.5390 ;
        RECT 0.1710 65.6235 3.7170 66.7170 ;
        RECT 0.0000 65.6235 0.1530 66.5390 ;
        RECT 5.0940 65.6235 9.6120 66.4430 ;
        RECT 0.0000 65.7230 5.0760 66.4430 ;
        RECT 4.8690 65.6235 9.6120 65.7950 ;
        RECT 0.0000 65.6235 4.8510 66.4430 ;
        RECT 0.0000 65.6235 9.6120 65.6990 ;
        RECT 0.0000 67.6670 9.6120 67.7970 ;
        RECT 9.4950 66.7035 9.6120 67.7970 ;
        RECT 5.8410 67.5710 9.4770 67.7970 ;
        RECT 4.5090 67.5710 5.8230 67.7970 ;
        RECT 3.7890 66.7035 4.4190 67.7970 ;
        RECT 0.1350 67.5710 3.7710 67.7970 ;
        RECT 0.0000 66.7035 0.1170 67.7970 ;
        RECT 9.4590 66.7035 9.6120 67.6190 ;
        RECT 5.8950 66.7035 9.4410 67.7970 ;
        RECT 5.1480 66.7035 5.8770 67.6190 ;
        RECT 4.9860 66.8990 5.1120 67.7970 ;
        RECT 3.7350 66.8030 4.9590 67.6190 ;
        RECT 0.1710 66.7035 3.7170 67.7970 ;
        RECT 0.0000 66.7035 0.1530 67.6190 ;
        RECT 5.0940 66.7035 9.6120 67.5230 ;
        RECT 0.0000 66.8030 5.0760 67.5230 ;
        RECT 4.8690 66.7035 9.6120 66.8750 ;
        RECT 0.0000 66.7035 4.8510 67.5230 ;
        RECT 0.0000 66.7035 9.6120 66.7790 ;
        RECT 0.0000 68.7470 9.6120 68.8770 ;
        RECT 9.4950 67.7835 9.6120 68.8770 ;
        RECT 5.8410 68.6510 9.4770 68.8770 ;
        RECT 4.5090 68.6510 5.8230 68.8770 ;
        RECT 3.7890 67.7835 4.4190 68.8770 ;
        RECT 0.1350 68.6510 3.7710 68.8770 ;
        RECT 0.0000 67.7835 0.1170 68.8770 ;
        RECT 9.4590 67.7835 9.6120 68.6990 ;
        RECT 5.8950 67.7835 9.4410 68.8770 ;
        RECT 5.1480 67.7835 5.8770 68.6990 ;
        RECT 4.9860 67.9790 5.1120 68.8770 ;
        RECT 3.7350 67.8830 4.9590 68.6990 ;
        RECT 0.1710 67.7835 3.7170 68.8770 ;
        RECT 0.0000 67.7835 0.1530 68.6990 ;
        RECT 5.0940 67.7835 9.6120 68.6030 ;
        RECT 0.0000 67.8830 5.0760 68.6030 ;
        RECT 4.8690 67.7835 9.6120 67.9550 ;
        RECT 0.0000 67.7835 4.8510 68.6030 ;
        RECT 0.0000 67.7835 9.6120 67.8590 ;
        RECT 0.0000 69.8270 9.6120 69.9570 ;
        RECT 9.4950 68.8635 9.6120 69.9570 ;
        RECT 5.8410 69.7310 9.4770 69.9570 ;
        RECT 4.5090 69.7310 5.8230 69.9570 ;
        RECT 3.7890 68.8635 4.4190 69.9570 ;
        RECT 0.1350 69.7310 3.7710 69.9570 ;
        RECT 0.0000 68.8635 0.1170 69.9570 ;
        RECT 9.4590 68.8635 9.6120 69.7790 ;
        RECT 5.8950 68.8635 9.4410 69.9570 ;
        RECT 5.1480 68.8635 5.8770 69.7790 ;
        RECT 4.9860 69.0590 5.1120 69.9570 ;
        RECT 3.7350 68.9630 4.9590 69.7790 ;
        RECT 0.1710 68.8635 3.7170 69.9570 ;
        RECT 0.0000 68.8635 0.1530 69.7790 ;
        RECT 5.0940 68.8635 9.6120 69.6830 ;
        RECT 0.0000 68.9630 5.0760 69.6830 ;
        RECT 4.8690 68.8635 9.6120 69.0350 ;
        RECT 0.0000 68.8635 4.8510 69.6830 ;
        RECT 0.0000 68.8635 9.6120 68.9390 ;
        RECT 0.0000 70.9070 9.6120 71.0370 ;
        RECT 9.4950 69.9435 9.6120 71.0370 ;
        RECT 5.8410 70.8110 9.4770 71.0370 ;
        RECT 4.5090 70.8110 5.8230 71.0370 ;
        RECT 3.7890 69.9435 4.4190 71.0370 ;
        RECT 0.1350 70.8110 3.7710 71.0370 ;
        RECT 0.0000 69.9435 0.1170 71.0370 ;
        RECT 9.4590 69.9435 9.6120 70.8590 ;
        RECT 5.8950 69.9435 9.4410 71.0370 ;
        RECT 5.1480 69.9435 5.8770 70.8590 ;
        RECT 4.9860 70.1390 5.1120 71.0370 ;
        RECT 3.7350 70.0430 4.9590 70.8590 ;
        RECT 0.1710 69.9435 3.7170 71.0370 ;
        RECT 0.0000 69.9435 0.1530 70.8590 ;
        RECT 5.0940 69.9435 9.6120 70.7630 ;
        RECT 0.0000 70.0430 5.0760 70.7630 ;
        RECT 4.8690 69.9435 9.6120 70.1150 ;
        RECT 0.0000 69.9435 4.8510 70.7630 ;
        RECT 0.0000 69.9435 9.6120 70.0190 ;
        RECT 0.0000 71.9870 9.6120 72.1170 ;
        RECT 9.4950 71.0235 9.6120 72.1170 ;
        RECT 5.8410 71.8910 9.4770 72.1170 ;
        RECT 4.5090 71.8910 5.8230 72.1170 ;
        RECT 3.7890 71.0235 4.4190 72.1170 ;
        RECT 0.1350 71.8910 3.7710 72.1170 ;
        RECT 0.0000 71.0235 0.1170 72.1170 ;
        RECT 9.4590 71.0235 9.6120 71.9390 ;
        RECT 5.8950 71.0235 9.4410 72.1170 ;
        RECT 5.1480 71.0235 5.8770 71.9390 ;
        RECT 4.9860 71.2190 5.1120 72.1170 ;
        RECT 3.7350 71.1230 4.9590 71.9390 ;
        RECT 0.1710 71.0235 3.7170 72.1170 ;
        RECT 0.0000 71.0235 0.1530 71.9390 ;
        RECT 5.0940 71.0235 9.6120 71.8430 ;
        RECT 0.0000 71.1230 5.0760 71.8430 ;
        RECT 4.8690 71.0235 9.6120 71.1950 ;
        RECT 0.0000 71.0235 4.8510 71.8430 ;
        RECT 0.0000 71.0235 9.6120 71.0990 ;
        RECT 0.0000 73.0670 9.6120 73.1970 ;
        RECT 9.4950 72.1035 9.6120 73.1970 ;
        RECT 5.8410 72.9710 9.4770 73.1970 ;
        RECT 4.5090 72.9710 5.8230 73.1970 ;
        RECT 3.7890 72.1035 4.4190 73.1970 ;
        RECT 0.1350 72.9710 3.7710 73.1970 ;
        RECT 0.0000 72.1035 0.1170 73.1970 ;
        RECT 9.4590 72.1035 9.6120 73.0190 ;
        RECT 5.8950 72.1035 9.4410 73.1970 ;
        RECT 5.1480 72.1035 5.8770 73.0190 ;
        RECT 4.9860 72.2990 5.1120 73.1970 ;
        RECT 3.7350 72.2030 4.9590 73.0190 ;
        RECT 0.1710 72.1035 3.7170 73.1970 ;
        RECT 0.0000 72.1035 0.1530 73.0190 ;
        RECT 5.0940 72.1035 9.6120 72.9230 ;
        RECT 0.0000 72.2030 5.0760 72.9230 ;
        RECT 4.8690 72.1035 9.6120 72.2750 ;
        RECT 0.0000 72.1035 4.8510 72.9230 ;
        RECT 0.0000 72.1035 9.6120 72.1790 ;
        RECT 0.0000 74.1470 9.6120 74.2770 ;
        RECT 9.4950 73.1835 9.6120 74.2770 ;
        RECT 5.8410 74.0510 9.4770 74.2770 ;
        RECT 4.5090 74.0510 5.8230 74.2770 ;
        RECT 3.7890 73.1835 4.4190 74.2770 ;
        RECT 0.1350 74.0510 3.7710 74.2770 ;
        RECT 0.0000 73.1835 0.1170 74.2770 ;
        RECT 9.4590 73.1835 9.6120 74.0990 ;
        RECT 5.8950 73.1835 9.4410 74.2770 ;
        RECT 5.1480 73.1835 5.8770 74.0990 ;
        RECT 4.9860 73.3790 5.1120 74.2770 ;
        RECT 3.7350 73.2830 4.9590 74.0990 ;
        RECT 0.1710 73.1835 3.7170 74.2770 ;
        RECT 0.0000 73.1835 0.1530 74.0990 ;
        RECT 5.0940 73.1835 9.6120 74.0030 ;
        RECT 0.0000 73.2830 5.0760 74.0030 ;
        RECT 4.8690 73.1835 9.6120 73.3550 ;
        RECT 0.0000 73.1835 4.8510 74.0030 ;
        RECT 0.0000 73.1835 9.6120 73.2590 ;
        RECT 0.0000 75.2270 9.6120 75.3570 ;
        RECT 9.4950 74.2635 9.6120 75.3570 ;
        RECT 5.8410 75.1310 9.4770 75.3570 ;
        RECT 4.5090 75.1310 5.8230 75.3570 ;
        RECT 3.7890 74.2635 4.4190 75.3570 ;
        RECT 0.1350 75.1310 3.7710 75.3570 ;
        RECT 0.0000 74.2635 0.1170 75.3570 ;
        RECT 9.4590 74.2635 9.6120 75.1790 ;
        RECT 5.8950 74.2635 9.4410 75.3570 ;
        RECT 5.1480 74.2635 5.8770 75.1790 ;
        RECT 4.9860 74.4590 5.1120 75.3570 ;
        RECT 3.7350 74.3630 4.9590 75.1790 ;
        RECT 0.1710 74.2635 3.7170 75.3570 ;
        RECT 0.0000 74.2635 0.1530 75.1790 ;
        RECT 5.0940 74.2635 9.6120 75.0830 ;
        RECT 0.0000 74.3630 5.0760 75.0830 ;
        RECT 4.8690 74.2635 9.6120 74.4350 ;
        RECT 0.0000 74.2635 4.8510 75.0830 ;
        RECT 0.0000 74.2635 9.6120 74.3390 ;
        RECT 0.0000 76.3070 9.6120 76.4370 ;
        RECT 9.4950 75.3435 9.6120 76.4370 ;
        RECT 5.8410 76.2110 9.4770 76.4370 ;
        RECT 4.5090 76.2110 5.8230 76.4370 ;
        RECT 3.7890 75.3435 4.4190 76.4370 ;
        RECT 0.1350 76.2110 3.7710 76.4370 ;
        RECT 0.0000 75.3435 0.1170 76.4370 ;
        RECT 9.4590 75.3435 9.6120 76.2590 ;
        RECT 5.8950 75.3435 9.4410 76.4370 ;
        RECT 5.1480 75.3435 5.8770 76.2590 ;
        RECT 4.9860 75.5390 5.1120 76.4370 ;
        RECT 3.7350 75.4430 4.9590 76.2590 ;
        RECT 0.1710 75.3435 3.7170 76.4370 ;
        RECT 0.0000 75.3435 0.1530 76.2590 ;
        RECT 5.0940 75.3435 9.6120 76.1630 ;
        RECT 0.0000 75.4430 5.0760 76.1630 ;
        RECT 4.8690 75.3435 9.6120 75.5150 ;
        RECT 0.0000 75.3435 4.8510 76.1630 ;
        RECT 0.0000 75.3435 9.6120 75.4190 ;
        RECT 0.0000 77.3870 9.6120 77.5170 ;
        RECT 9.4950 76.4235 9.6120 77.5170 ;
        RECT 5.8410 77.2910 9.4770 77.5170 ;
        RECT 4.5090 77.2910 5.8230 77.5170 ;
        RECT 3.7890 76.4235 4.4190 77.5170 ;
        RECT 0.1350 77.2910 3.7710 77.5170 ;
        RECT 0.0000 76.4235 0.1170 77.5170 ;
        RECT 9.4590 76.4235 9.6120 77.3390 ;
        RECT 5.8950 76.4235 9.4410 77.5170 ;
        RECT 5.1480 76.4235 5.8770 77.3390 ;
        RECT 4.9860 76.6190 5.1120 77.5170 ;
        RECT 3.7350 76.5230 4.9590 77.3390 ;
        RECT 0.1710 76.4235 3.7170 77.5170 ;
        RECT 0.0000 76.4235 0.1530 77.3390 ;
        RECT 5.0940 76.4235 9.6120 77.2430 ;
        RECT 0.0000 76.5230 5.0760 77.2430 ;
        RECT 4.8690 76.4235 9.6120 76.5950 ;
        RECT 0.0000 76.4235 4.8510 77.2430 ;
        RECT 0.0000 76.4235 9.6120 76.4990 ;
        RECT 0.0000 78.4670 9.6120 78.5970 ;
        RECT 9.4950 77.5035 9.6120 78.5970 ;
        RECT 5.8410 78.3710 9.4770 78.5970 ;
        RECT 4.5090 78.3710 5.8230 78.5970 ;
        RECT 3.7890 77.5035 4.4190 78.5970 ;
        RECT 0.1350 78.3710 3.7710 78.5970 ;
        RECT 0.0000 77.5035 0.1170 78.5970 ;
        RECT 9.4590 77.5035 9.6120 78.4190 ;
        RECT 5.8950 77.5035 9.4410 78.5970 ;
        RECT 5.1480 77.5035 5.8770 78.4190 ;
        RECT 4.9860 77.6990 5.1120 78.5970 ;
        RECT 3.7350 77.6030 4.9590 78.4190 ;
        RECT 0.1710 77.5035 3.7170 78.5970 ;
        RECT 0.0000 77.5035 0.1530 78.4190 ;
        RECT 5.0940 77.5035 9.6120 78.3230 ;
        RECT 0.0000 77.6030 5.0760 78.3230 ;
        RECT 4.8690 77.5035 9.6120 77.6750 ;
        RECT 0.0000 77.5035 4.8510 78.3230 ;
        RECT 0.0000 77.5035 9.6120 77.5790 ;
        RECT 0.0000 79.5470 9.6120 79.6770 ;
        RECT 9.4950 78.5835 9.6120 79.6770 ;
        RECT 5.8410 79.4510 9.4770 79.6770 ;
        RECT 4.5090 79.4510 5.8230 79.6770 ;
        RECT 3.7890 78.5835 4.4190 79.6770 ;
        RECT 0.1350 79.4510 3.7710 79.6770 ;
        RECT 0.0000 78.5835 0.1170 79.6770 ;
        RECT 9.4590 78.5835 9.6120 79.4990 ;
        RECT 5.8950 78.5835 9.4410 79.6770 ;
        RECT 5.1480 78.5835 5.8770 79.4990 ;
        RECT 4.9860 78.7790 5.1120 79.6770 ;
        RECT 3.7350 78.6830 4.9590 79.4990 ;
        RECT 0.1710 78.5835 3.7170 79.6770 ;
        RECT 0.0000 78.5835 0.1530 79.4990 ;
        RECT 5.0940 78.5835 9.6120 79.4030 ;
        RECT 0.0000 78.6830 5.0760 79.4030 ;
        RECT 4.8690 78.5835 9.6120 78.7550 ;
        RECT 0.0000 78.5835 4.8510 79.4030 ;
        RECT 0.0000 78.5835 9.6120 78.6590 ;
        RECT 0.0000 80.6270 9.6120 80.7570 ;
        RECT 9.4950 79.6635 9.6120 80.7570 ;
        RECT 5.8410 80.5310 9.4770 80.7570 ;
        RECT 4.5090 80.5310 5.8230 80.7570 ;
        RECT 3.7890 79.6635 4.4190 80.7570 ;
        RECT 0.1350 80.5310 3.7710 80.7570 ;
        RECT 0.0000 79.6635 0.1170 80.7570 ;
        RECT 9.4590 79.6635 9.6120 80.5790 ;
        RECT 5.8950 79.6635 9.4410 80.7570 ;
        RECT 5.1480 79.6635 5.8770 80.5790 ;
        RECT 4.9860 79.8590 5.1120 80.7570 ;
        RECT 3.7350 79.7630 4.9590 80.5790 ;
        RECT 0.1710 79.6635 3.7170 80.7570 ;
        RECT 0.0000 79.6635 0.1530 80.5790 ;
        RECT 5.0940 79.6635 9.6120 80.4830 ;
        RECT 0.0000 79.7630 5.0760 80.4830 ;
        RECT 4.8690 79.6635 9.6120 79.8350 ;
        RECT 0.0000 79.6635 4.8510 80.4830 ;
        RECT 0.0000 79.6635 9.6120 79.7390 ;
        RECT 0.0000 81.7070 9.6120 81.8370 ;
        RECT 9.4950 80.7435 9.6120 81.8370 ;
        RECT 5.8410 81.6110 9.4770 81.8370 ;
        RECT 4.5090 81.6110 5.8230 81.8370 ;
        RECT 3.7890 80.7435 4.4190 81.8370 ;
        RECT 0.1350 81.6110 3.7710 81.8370 ;
        RECT 0.0000 80.7435 0.1170 81.8370 ;
        RECT 9.4590 80.7435 9.6120 81.6590 ;
        RECT 5.8950 80.7435 9.4410 81.8370 ;
        RECT 5.1480 80.7435 5.8770 81.6590 ;
        RECT 4.9860 80.9390 5.1120 81.8370 ;
        RECT 3.7350 80.8430 4.9590 81.6590 ;
        RECT 0.1710 80.7435 3.7170 81.8370 ;
        RECT 0.0000 80.7435 0.1530 81.6590 ;
        RECT 5.0940 80.7435 9.6120 81.5630 ;
        RECT 0.0000 80.8430 5.0760 81.5630 ;
        RECT 4.8690 80.7435 9.6120 80.9150 ;
        RECT 0.0000 80.7435 4.8510 81.5630 ;
        RECT 0.0000 80.7435 9.6120 80.8190 ;
        RECT 0.0000 82.7870 9.6120 82.9170 ;
        RECT 9.4950 81.8235 9.6120 82.9170 ;
        RECT 5.8410 82.6910 9.4770 82.9170 ;
        RECT 4.5090 82.6910 5.8230 82.9170 ;
        RECT 3.7890 81.8235 4.4190 82.9170 ;
        RECT 0.1350 82.6910 3.7710 82.9170 ;
        RECT 0.0000 81.8235 0.1170 82.9170 ;
        RECT 9.4590 81.8235 9.6120 82.7390 ;
        RECT 5.8950 81.8235 9.4410 82.9170 ;
        RECT 5.1480 81.8235 5.8770 82.7390 ;
        RECT 4.9860 82.0190 5.1120 82.9170 ;
        RECT 3.7350 81.9230 4.9590 82.7390 ;
        RECT 0.1710 81.8235 3.7170 82.9170 ;
        RECT 0.0000 81.8235 0.1530 82.7390 ;
        RECT 5.0940 81.8235 9.6120 82.6430 ;
        RECT 0.0000 81.9230 5.0760 82.6430 ;
        RECT 4.8690 81.8235 9.6120 81.9950 ;
        RECT 0.0000 81.8235 4.8510 82.6430 ;
        RECT 0.0000 81.8235 9.6120 81.8990 ;
        RECT 0.0000 83.8670 9.6120 83.9970 ;
        RECT 9.4950 82.9035 9.6120 83.9970 ;
        RECT 5.8410 83.7710 9.4770 83.9970 ;
        RECT 4.5090 83.7710 5.8230 83.9970 ;
        RECT 3.7890 82.9035 4.4190 83.9970 ;
        RECT 0.1350 83.7710 3.7710 83.9970 ;
        RECT 0.0000 82.9035 0.1170 83.9970 ;
        RECT 9.4590 82.9035 9.6120 83.8190 ;
        RECT 5.8950 82.9035 9.4410 83.9970 ;
        RECT 5.1480 82.9035 5.8770 83.8190 ;
        RECT 4.9860 83.0990 5.1120 83.9970 ;
        RECT 3.7350 83.0030 4.9590 83.8190 ;
        RECT 0.1710 82.9035 3.7170 83.9970 ;
        RECT 0.0000 82.9035 0.1530 83.8190 ;
        RECT 5.0940 82.9035 9.6120 83.7230 ;
        RECT 0.0000 83.0030 5.0760 83.7230 ;
        RECT 4.8690 82.9035 9.6120 83.0750 ;
        RECT 0.0000 82.9035 4.8510 83.7230 ;
        RECT 0.0000 82.9035 9.6120 82.9790 ;
        RECT 0.0000 84.9470 9.6120 85.0770 ;
        RECT 9.4950 83.9835 9.6120 85.0770 ;
        RECT 5.8410 84.8510 9.4770 85.0770 ;
        RECT 4.5090 84.8510 5.8230 85.0770 ;
        RECT 3.7890 83.9835 4.4190 85.0770 ;
        RECT 0.1350 84.8510 3.7710 85.0770 ;
        RECT 0.0000 83.9835 0.1170 85.0770 ;
        RECT 9.4590 83.9835 9.6120 84.8990 ;
        RECT 5.8950 83.9835 9.4410 85.0770 ;
        RECT 5.1480 83.9835 5.8770 84.8990 ;
        RECT 4.9860 84.1790 5.1120 85.0770 ;
        RECT 3.7350 84.0830 4.9590 84.8990 ;
        RECT 0.1710 83.9835 3.7170 85.0770 ;
        RECT 0.0000 83.9835 0.1530 84.8990 ;
        RECT 5.0940 83.9835 9.6120 84.8030 ;
        RECT 0.0000 84.0830 5.0760 84.8030 ;
        RECT 4.8690 83.9835 9.6120 84.1550 ;
        RECT 0.0000 83.9835 4.8510 84.8030 ;
        RECT 0.0000 83.9835 9.6120 84.0590 ;
        RECT 0.0000 86.0270 9.6120 86.1570 ;
        RECT 9.4950 85.0635 9.6120 86.1570 ;
        RECT 5.8410 85.9310 9.4770 86.1570 ;
        RECT 4.5090 85.9310 5.8230 86.1570 ;
        RECT 3.7890 85.0635 4.4190 86.1570 ;
        RECT 0.1350 85.9310 3.7710 86.1570 ;
        RECT 0.0000 85.0635 0.1170 86.1570 ;
        RECT 9.4590 85.0635 9.6120 85.9790 ;
        RECT 5.8950 85.0635 9.4410 86.1570 ;
        RECT 5.1480 85.0635 5.8770 85.9790 ;
        RECT 4.9860 85.2590 5.1120 86.1570 ;
        RECT 3.7350 85.1630 4.9590 85.9790 ;
        RECT 0.1710 85.0635 3.7170 86.1570 ;
        RECT 0.0000 85.0635 0.1530 85.9790 ;
        RECT 5.0940 85.0635 9.6120 85.8830 ;
        RECT 0.0000 85.1630 5.0760 85.8830 ;
        RECT 4.8690 85.0635 9.6120 85.2350 ;
        RECT 0.0000 85.0635 4.8510 85.8830 ;
        RECT 0.0000 85.0635 9.6120 85.1390 ;
        RECT 0.0000 87.1070 9.6120 87.2370 ;
        RECT 9.4950 86.1435 9.6120 87.2370 ;
        RECT 5.8410 87.0110 9.4770 87.2370 ;
        RECT 4.5090 87.0110 5.8230 87.2370 ;
        RECT 3.7890 86.1435 4.4190 87.2370 ;
        RECT 0.1350 87.0110 3.7710 87.2370 ;
        RECT 0.0000 86.1435 0.1170 87.2370 ;
        RECT 9.4590 86.1435 9.6120 87.0590 ;
        RECT 5.8950 86.1435 9.4410 87.2370 ;
        RECT 5.1480 86.1435 5.8770 87.0590 ;
        RECT 4.9860 86.3390 5.1120 87.2370 ;
        RECT 3.7350 86.2430 4.9590 87.0590 ;
        RECT 0.1710 86.1435 3.7170 87.2370 ;
        RECT 0.0000 86.1435 0.1530 87.0590 ;
        RECT 5.0940 86.1435 9.6120 86.9630 ;
        RECT 0.0000 86.2430 5.0760 86.9630 ;
        RECT 4.8690 86.1435 9.6120 86.3150 ;
        RECT 0.0000 86.1435 4.8510 86.9630 ;
        RECT 0.0000 86.1435 9.6120 86.2190 ;
        RECT 0.0000 88.1870 9.6120 88.3170 ;
        RECT 9.4950 87.2235 9.6120 88.3170 ;
        RECT 5.8410 88.0910 9.4770 88.3170 ;
        RECT 4.5090 88.0910 5.8230 88.3170 ;
        RECT 3.7890 87.2235 4.4190 88.3170 ;
        RECT 0.1350 88.0910 3.7710 88.3170 ;
        RECT 0.0000 87.2235 0.1170 88.3170 ;
        RECT 9.4590 87.2235 9.6120 88.1390 ;
        RECT 5.8950 87.2235 9.4410 88.3170 ;
        RECT 5.1480 87.2235 5.8770 88.1390 ;
        RECT 4.9860 87.4190 5.1120 88.3170 ;
        RECT 3.7350 87.3230 4.9590 88.1390 ;
        RECT 0.1710 87.2235 3.7170 88.3170 ;
        RECT 0.0000 87.2235 0.1530 88.1390 ;
        RECT 5.0940 87.2235 9.6120 88.0430 ;
        RECT 0.0000 87.3230 5.0760 88.0430 ;
        RECT 4.8690 87.2235 9.6120 87.3950 ;
        RECT 0.0000 87.2235 4.8510 88.0430 ;
        RECT 0.0000 87.2235 9.6120 87.2990 ;
        RECT 0.0000 89.2670 9.6120 89.3970 ;
        RECT 9.4950 88.3035 9.6120 89.3970 ;
        RECT 5.8410 89.1710 9.4770 89.3970 ;
        RECT 4.5090 89.1710 5.8230 89.3970 ;
        RECT 3.7890 88.3035 4.4190 89.3970 ;
        RECT 0.1350 89.1710 3.7710 89.3970 ;
        RECT 0.0000 88.3035 0.1170 89.3970 ;
        RECT 9.4590 88.3035 9.6120 89.2190 ;
        RECT 5.8950 88.3035 9.4410 89.3970 ;
        RECT 5.1480 88.3035 5.8770 89.2190 ;
        RECT 4.9860 88.4990 5.1120 89.3970 ;
        RECT 3.7350 88.4030 4.9590 89.2190 ;
        RECT 0.1710 88.3035 3.7170 89.3970 ;
        RECT 0.0000 88.3035 0.1530 89.2190 ;
        RECT 5.0940 88.3035 9.6120 89.1230 ;
        RECT 0.0000 88.4030 5.0760 89.1230 ;
        RECT 4.8690 88.3035 9.6120 88.4750 ;
        RECT 0.0000 88.3035 4.8510 89.1230 ;
        RECT 0.0000 88.3035 9.6120 88.3790 ;
        RECT 0.0000 90.3470 9.6120 90.4770 ;
        RECT 9.4950 89.3835 9.6120 90.4770 ;
        RECT 5.8410 90.2510 9.4770 90.4770 ;
        RECT 4.5090 90.2510 5.8230 90.4770 ;
        RECT 3.7890 89.3835 4.4190 90.4770 ;
        RECT 0.1350 90.2510 3.7710 90.4770 ;
        RECT 0.0000 89.3835 0.1170 90.4770 ;
        RECT 9.4590 89.3835 9.6120 90.2990 ;
        RECT 5.8950 89.3835 9.4410 90.4770 ;
        RECT 5.1480 89.3835 5.8770 90.2990 ;
        RECT 4.9860 89.5790 5.1120 90.4770 ;
        RECT 3.7350 89.4830 4.9590 90.2990 ;
        RECT 0.1710 89.3835 3.7170 90.4770 ;
        RECT 0.0000 89.3835 0.1530 90.2990 ;
        RECT 5.0940 89.3835 9.6120 90.2030 ;
        RECT 0.0000 89.4830 5.0760 90.2030 ;
        RECT 4.8690 89.3835 9.6120 89.5550 ;
        RECT 0.0000 89.3835 4.8510 90.2030 ;
        RECT 0.0000 89.3835 9.6120 89.4590 ;
        RECT 0.0000 91.4270 9.6120 91.5570 ;
        RECT 9.4950 90.4635 9.6120 91.5570 ;
        RECT 5.8410 91.3310 9.4770 91.5570 ;
        RECT 4.5090 91.3310 5.8230 91.5570 ;
        RECT 3.7890 90.4635 4.4190 91.5570 ;
        RECT 0.1350 91.3310 3.7710 91.5570 ;
        RECT 0.0000 90.4635 0.1170 91.5570 ;
        RECT 9.4590 90.4635 9.6120 91.3790 ;
        RECT 5.8950 90.4635 9.4410 91.5570 ;
        RECT 5.1480 90.4635 5.8770 91.3790 ;
        RECT 4.9860 90.6590 5.1120 91.5570 ;
        RECT 3.7350 90.5630 4.9590 91.3790 ;
        RECT 0.1710 90.4635 3.7170 91.5570 ;
        RECT 0.0000 90.4635 0.1530 91.3790 ;
        RECT 5.0940 90.4635 9.6120 91.2830 ;
        RECT 0.0000 90.5630 5.0760 91.2830 ;
        RECT 4.8690 90.4635 9.6120 90.6350 ;
        RECT 0.0000 90.4635 4.8510 91.2830 ;
        RECT 0.0000 90.4635 9.6120 90.5390 ;
        RECT 0.0000 92.5070 9.6120 92.6370 ;
        RECT 9.4950 91.5435 9.6120 92.6370 ;
        RECT 5.8410 92.4110 9.4770 92.6370 ;
        RECT 4.5090 92.4110 5.8230 92.6370 ;
        RECT 3.7890 91.5435 4.4190 92.6370 ;
        RECT 0.1350 92.4110 3.7710 92.6370 ;
        RECT 0.0000 91.5435 0.1170 92.6370 ;
        RECT 9.4590 91.5435 9.6120 92.4590 ;
        RECT 5.8950 91.5435 9.4410 92.6370 ;
        RECT 5.1480 91.5435 5.8770 92.4590 ;
        RECT 4.9860 91.7390 5.1120 92.6370 ;
        RECT 3.7350 91.6430 4.9590 92.4590 ;
        RECT 0.1710 91.5435 3.7170 92.6370 ;
        RECT 0.0000 91.5435 0.1530 92.4590 ;
        RECT 5.0940 91.5435 9.6120 92.3630 ;
        RECT 0.0000 91.6430 5.0760 92.3630 ;
        RECT 4.8690 91.5435 9.6120 91.7150 ;
        RECT 0.0000 91.5435 4.8510 92.3630 ;
        RECT 0.0000 91.5435 9.6120 91.6190 ;
        RECT 0.0000 93.5870 9.6120 93.7170 ;
        RECT 9.4950 92.6235 9.6120 93.7170 ;
        RECT 5.8410 93.4910 9.4770 93.7170 ;
        RECT 4.5090 93.4910 5.8230 93.7170 ;
        RECT 3.7890 92.6235 4.4190 93.7170 ;
        RECT 0.1350 93.4910 3.7710 93.7170 ;
        RECT 0.0000 92.6235 0.1170 93.7170 ;
        RECT 9.4590 92.6235 9.6120 93.5390 ;
        RECT 5.8950 92.6235 9.4410 93.7170 ;
        RECT 5.1480 92.6235 5.8770 93.5390 ;
        RECT 4.9860 92.8190 5.1120 93.7170 ;
        RECT 3.7350 92.7230 4.9590 93.5390 ;
        RECT 0.1710 92.6235 3.7170 93.7170 ;
        RECT 0.0000 92.6235 0.1530 93.5390 ;
        RECT 5.0940 92.6235 9.6120 93.4430 ;
        RECT 0.0000 92.7230 5.0760 93.4430 ;
        RECT 4.8690 92.6235 9.6120 92.7950 ;
        RECT 0.0000 92.6235 4.8510 93.4430 ;
        RECT 0.0000 92.6235 9.6120 92.6990 ;
        RECT 0.0000 94.6670 9.6120 94.7970 ;
        RECT 9.4950 93.7035 9.6120 94.7970 ;
        RECT 5.8410 94.5710 9.4770 94.7970 ;
        RECT 4.5090 94.5710 5.8230 94.7970 ;
        RECT 3.7890 93.7035 4.4190 94.7970 ;
        RECT 0.1350 94.5710 3.7710 94.7970 ;
        RECT 0.0000 93.7035 0.1170 94.7970 ;
        RECT 9.4590 93.7035 9.6120 94.6190 ;
        RECT 5.8950 93.7035 9.4410 94.7970 ;
        RECT 5.1480 93.7035 5.8770 94.6190 ;
        RECT 4.9860 93.8990 5.1120 94.7970 ;
        RECT 3.7350 93.8030 4.9590 94.6190 ;
        RECT 0.1710 93.7035 3.7170 94.7970 ;
        RECT 0.0000 93.7035 0.1530 94.6190 ;
        RECT 5.0940 93.7035 9.6120 94.5230 ;
        RECT 0.0000 93.8030 5.0760 94.5230 ;
        RECT 4.8690 93.7035 9.6120 93.8750 ;
        RECT 0.0000 93.7035 4.8510 94.5230 ;
        RECT 0.0000 93.7035 9.6120 93.7790 ;
  LAYER M4  ;
      RECT 1.6070 45.1560 8.0025 45.1800 ;
      RECT 1.6070 45.4440 8.0025 45.4680 ;
      RECT 1.6070 45.8280 8.0025 45.8520 ;
      RECT 1.6070 45.9240 8.0025 45.9480 ;
      RECT 1.6070 46.2600 8.0025 46.2840 ;
      RECT 7.4990 44.1150 7.5830 44.1390 ;
      RECT 7.3190 44.5470 7.4360 44.5710 ;
      RECT 7.3190 45.2040 7.4360 45.2280 ;
      RECT 7.3190 45.4920 7.4360 45.5160 ;
      RECT 6.6785 44.5470 7.2480 44.5710 ;
      RECT 6.7430 45.3240 6.8510 45.3480 ;
      RECT 5.4070 45.6990 6.5000 45.7230 ;
      RECT 6.0950 45.2670 6.1790 45.2910 ;
      RECT 5.3110 46.4670 6.1790 46.4910 ;
      RECT 6.0950 46.5630 6.1790 46.5870 ;
      RECT 5.9170 44.7870 6.0010 44.8110 ;
      RECT 5.8790 46.1310 5.9630 46.1550 ;
      RECT 5.7010 44.6910 5.7850 44.7150 ;
      RECT 5.4870 43.4030 5.7500 43.4270 ;
      RECT 5.4870 52.0430 5.7500 52.0670 ;
      RECT 5.5030 46.1790 5.7470 46.2030 ;
      RECT 5.6630 46.3230 5.7470 46.3470 ;
      RECT 4.2070 46.5630 5.7470 46.5870 ;
      RECT 5.6630 46.8510 5.7470 46.8750 ;
      RECT 5.4290 51.9470 5.6920 51.9710 ;
      RECT 5.4280 43.3070 5.6910 43.3310 ;
      RECT 5.3900 43.2110 5.6530 43.2350 ;
      RECT 5.3900 51.7550 5.6530 51.7790 ;
      RECT 5.5550 47.2830 5.6390 47.3070 ;
      RECT 4.7830 47.6670 5.6390 47.6910 ;
      RECT 5.1670 49.9230 5.6390 49.9470 ;
      RECT 5.5550 50.0190 5.6390 50.0430 ;
      RECT 5.3420 43.1150 5.6050 43.1390 ;
      RECT 5.3420 51.6590 5.6050 51.6830 ;
      RECT 5.1190 49.0110 5.5640 49.0350 ;
      RECT 5.2980 43.0190 5.5610 43.0430 ;
      RECT 5.2980 51.9950 5.5610 52.0190 ;
      RECT 5.2490 43.3550 5.5120 43.3790 ;
      RECT 5.2490 51.8990 5.5120 51.9230 ;
      RECT 5.3800 46.3230 5.5010 46.3470 ;
      RECT 5.3590 48.4350 5.4920 48.4590 ;
      RECT 5.2020 43.2590 5.4650 43.2830 ;
      RECT 5.2020 51.8030 5.4650 51.8270 ;
      RECT 5.1670 42.9710 5.4300 42.9950 ;
      RECT 5.1670 51.7070 5.4300 51.7310 ;
      RECT 4.3510 50.0190 5.4200 50.0430 ;
      RECT 5.3360 51.1710 5.4200 51.1950 ;
      RECT 5.1110 42.8270 5.3740 42.8510 ;
      RECT 5.1110 51.6110 5.3740 51.6350 ;
      RECT 5.2630 47.2830 5.3480 47.3070 ;
      RECT 4.1590 47.8590 5.2760 47.8830 ;
      RECT 4.8040 45.6990 5.2610 45.7230 ;
      RECT 4.6310 43.5470 4.8980 43.5710 ;
      RECT 4.6310 51.4670 4.8980 51.4910 ;
      RECT 4.7680 47.2350 4.8770 47.2590 ;
      RECT 4.6080 43.4510 4.8500 43.4750 ;
      RECT 4.6080 52.0910 4.8500 52.1150 ;
      RECT 4.5520 42.9710 4.7940 42.9950 ;
      RECT 4.5810 52.1870 4.7940 52.2110 ;
      RECT 4.6970 46.8510 4.7810 46.8750 ;
      RECT 4.4980 43.0670 4.7460 43.0910 ;
      RECT 4.4980 52.0430 4.7460 52.0670 ;
      RECT 4.2640 49.4430 4.6850 49.4670 ;
      RECT 4.2320 43.4030 4.4990 43.4270 ;
      RECT 4.2320 52.1870 4.4990 52.2110 ;
      RECT 4.3720 48.0030 4.4930 48.0270 ;
      RECT 4.3640 51.1710 4.4480 51.1950 ;
      RECT 4.1980 43.3070 4.4450 43.3310 ;
      RECT 4.1310 51.7550 4.4450 51.7790 ;
      RECT 4.1720 43.2110 4.4020 43.2350 ;
      RECT 4.1600 52.0910 4.4020 52.1150 ;
      RECT 4.1190 43.1150 4.3490 43.1390 ;
      RECT 4.2650 49.5870 4.3490 49.6110 ;
      RECT 4.0690 51.6590 4.3490 51.6830 ;
      RECT 4.0740 43.0190 4.3040 43.0430 ;
      RECT 4.0740 51.9950 4.3040 52.0190 ;
      RECT 3.1120 46.8510 4.3010 46.8750 ;
      RECT 4.0360 43.2590 4.2660 43.2830 ;
      RECT 4.0360 51.8990 4.2660 51.9230 ;
      RECT 4.0180 43.1630 4.2110 43.1870 ;
      RECT 4.0180 51.8030 4.2110 51.8270 ;
      RECT 3.9690 43.0670 4.1620 43.0910 ;
      RECT 3.9690 51.7070 4.1620 51.7310 ;
      RECT 3.9730 47.7630 4.1570 47.7870 ;
      RECT 3.9170 42.9710 4.1100 42.9950 ;
      RECT 3.9170 51.6110 4.1100 51.6350 ;
      RECT 3.4330 45.0750 4.1090 45.0990 ;
      RECT 3.9730 47.8590 4.0570 47.8830 ;
      RECT 3.7040 43.4990 3.9670 43.5230 ;
      RECT 3.7580 47.2830 3.8700 47.3070 ;
      RECT 3.3950 45.2670 3.4790 45.2910 ;
  LAYER V4  ;
      RECT 7.5480 44.1150 7.5720 44.1390 ;
      RECT 7.5480 45.1560 7.5720 45.1800 ;
      RECT 7.3800 44.5470 7.4040 44.5710 ;
      RECT 7.3800 45.2040 7.4040 45.2280 ;
      RECT 7.3800 45.4920 7.4040 45.5160 ;
      RECT 6.7560 44.5470 6.7800 44.5710 ;
      RECT 6.7560 45.3240 6.7800 45.3480 ;
      RECT 6.1440 45.2670 6.1680 45.2910 ;
      RECT 6.1440 45.4440 6.1680 45.4680 ;
      RECT 6.1440 46.4670 6.1680 46.4910 ;
      RECT 6.1440 46.5630 6.1680 46.5870 ;
      RECT 5.9280 44.7870 5.9520 44.8110 ;
      RECT 5.9280 45.8280 5.9520 45.8520 ;
      RECT 5.9280 46.1310 5.9520 46.1550 ;
      RECT 5.9280 46.2600 5.9520 46.2840 ;
      RECT 5.7120 44.6910 5.7360 44.7150 ;
      RECT 5.7120 45.9240 5.7360 45.9480 ;
      RECT 5.7120 46.1790 5.7360 46.2030 ;
      RECT 5.7120 46.3230 5.7360 46.3470 ;
      RECT 5.7120 46.5630 5.7360 46.5870 ;
      RECT 5.7120 46.8510 5.7360 46.8750 ;
      RECT 5.6040 47.2830 5.6280 47.3070 ;
      RECT 5.6040 47.6670 5.6280 47.6910 ;
      RECT 5.6040 49.9230 5.6280 49.9470 ;
      RECT 5.6040 50.0190 5.6280 50.0430 ;
      RECT 5.5140 43.4030 5.5380 43.4270 ;
      RECT 5.5140 46.1790 5.5380 46.2030 ;
      RECT 5.5140 52.0430 5.5380 52.0670 ;
      RECT 5.4660 43.3070 5.4900 43.3310 ;
      RECT 5.4660 46.3230 5.4900 46.3470 ;
      RECT 5.4660 51.9470 5.4900 51.9710 ;
      RECT 5.4180 43.2110 5.4420 43.2350 ;
      RECT 5.4180 45.6990 5.4420 45.7230 ;
      RECT 5.4180 51.7550 5.4420 51.7790 ;
      RECT 5.3700 43.1150 5.3940 43.1390 ;
      RECT 5.3700 48.4350 5.3940 48.4590 ;
      RECT 5.3700 51.1710 5.3940 51.1950 ;
      RECT 5.3700 51.6590 5.3940 51.6830 ;
      RECT 5.3220 43.0190 5.3460 43.0430 ;
      RECT 5.3220 46.4670 5.3460 46.4910 ;
      RECT 5.3220 51.9950 5.3460 52.0190 ;
      RECT 5.2740 43.3550 5.2980 43.3790 ;
      RECT 5.2740 47.2830 5.2980 47.3070 ;
      RECT 5.2740 51.8990 5.2980 51.9230 ;
      RECT 5.2260 43.2590 5.2500 43.2830 ;
      RECT 5.2260 45.6990 5.2500 45.7230 ;
      RECT 5.2260 51.8030 5.2500 51.8270 ;
      RECT 5.1780 42.9710 5.2020 42.9950 ;
      RECT 5.1780 49.9230 5.2020 49.9470 ;
      RECT 5.1780 51.7070 5.2020 51.7310 ;
      RECT 5.1300 42.8270 5.1540 42.8510 ;
      RECT 5.1300 49.0110 5.1540 49.0350 ;
      RECT 5.1300 51.6110 5.1540 51.6350 ;
      RECT 4.8420 43.5470 4.8660 43.5710 ;
      RECT 4.8420 47.2350 4.8660 47.2590 ;
      RECT 4.8420 51.4670 4.8660 51.4910 ;
      RECT 4.7940 43.4510 4.8180 43.4750 ;
      RECT 4.7940 47.6670 4.8180 47.6910 ;
      RECT 4.7940 52.0910 4.8180 52.1150 ;
      RECT 4.7460 42.9710 4.7700 42.9950 ;
      RECT 4.7460 46.8510 4.7700 46.8750 ;
      RECT 4.7460 52.1870 4.7700 52.2110 ;
      RECT 4.6500 43.0670 4.6740 43.0910 ;
      RECT 4.6500 49.4430 4.6740 49.4670 ;
      RECT 4.6500 52.0430 4.6740 52.0670 ;
      RECT 4.4580 43.4030 4.4820 43.4270 ;
      RECT 4.4580 48.0030 4.4820 48.0270 ;
      RECT 4.4580 52.1870 4.4820 52.2110 ;
      RECT 4.4100 43.3070 4.4340 43.3310 ;
      RECT 4.4100 51.1710 4.4340 51.1950 ;
      RECT 4.4100 51.7550 4.4340 51.7790 ;
      RECT 4.3620 43.2110 4.3860 43.2350 ;
      RECT 4.3620 50.0190 4.3860 50.0430 ;
      RECT 4.3620 52.0910 4.3860 52.1150 ;
      RECT 4.3140 43.1150 4.3380 43.1390 ;
      RECT 4.3140 49.5870 4.3380 49.6110 ;
      RECT 4.3140 51.6590 4.3380 51.6830 ;
      RECT 4.2660 43.0190 4.2900 43.0430 ;
      RECT 4.2660 46.8510 4.2900 46.8750 ;
      RECT 4.2660 51.9950 4.2900 52.0190 ;
      RECT 4.2180 43.2590 4.2420 43.2830 ;
      RECT 4.2180 46.5630 4.2420 46.5870 ;
      RECT 4.2180 51.8990 4.2420 51.9230 ;
      RECT 4.1700 43.1630 4.1940 43.1870 ;
      RECT 4.1700 47.8590 4.1940 47.8830 ;
      RECT 4.1700 51.8030 4.1940 51.8270 ;
      RECT 4.1220 43.0670 4.1460 43.0910 ;
      RECT 4.1220 47.7630 4.1460 47.7870 ;
      RECT 4.1220 51.7070 4.1460 51.7310 ;
      RECT 4.0740 42.9710 4.0980 42.9950 ;
      RECT 4.0740 45.0750 4.0980 45.0990 ;
      RECT 4.0740 51.6110 4.0980 51.6350 ;
      RECT 3.9840 47.7630 4.0080 47.7870 ;
      RECT 3.9840 47.8590 4.0080 47.8830 ;
      RECT 3.8170 43.4990 3.8410 43.5230 ;
      RECT 3.8170 47.2830 3.8410 47.3070 ;
      RECT 3.4440 45.0750 3.4680 45.0990 ;
      RECT 3.4440 45.2670 3.4680 45.2910 ;
  LAYER M5  ;
      RECT 7.5480 44.1040 7.5720 45.1910 ;
      RECT 7.3800 44.5335 7.4040 45.5660 ;
      RECT 6.7560 44.5275 6.7800 45.3600 ;
      RECT 6.1440 45.2560 6.1680 45.4790 ;
      RECT 6.1440 46.4560 6.1680 46.5980 ;
      RECT 5.9280 44.7760 5.9520 45.8630 ;
      RECT 5.9280 46.1200 5.9520 46.2950 ;
      RECT 5.7120 44.6800 5.7360 45.9590 ;
      RECT 5.7120 46.1680 5.7360 46.3580 ;
      RECT 5.7120 46.5520 5.7360 46.8860 ;
      RECT 5.6040 47.2720 5.6280 47.7020 ;
      RECT 5.6040 49.9120 5.6280 50.0540 ;
      RECT 5.5140 43.7400 5.5380 51.3230 ;
      RECT 5.4660 43.7400 5.4900 51.3230 ;
      RECT 5.4180 43.7400 5.4420 51.3230 ;
      RECT 5.3700 43.7400 5.3940 51.3230 ;
      RECT 5.3220 43.7400 5.3460 51.3230 ;
      RECT 5.2740 43.7400 5.2980 51.3230 ;
      RECT 5.2260 43.7400 5.2500 51.3230 ;
      RECT 5.1780 43.7400 5.2020 51.3230 ;
      RECT 5.1300 43.7400 5.1540 51.3230 ;
      RECT 4.8420 43.4780 4.8660 51.5110 ;
      RECT 4.7940 42.9570 4.8180 52.2860 ;
      RECT 4.7460 42.9260 4.7700 52.2850 ;
      RECT 4.6500 42.9720 4.6740 52.2860 ;
      RECT 4.4580 42.9710 4.4820 52.2390 ;
      RECT 4.4100 42.9710 4.4340 52.2390 ;
      RECT 4.3620 42.9710 4.3860 52.2390 ;
      RECT 4.3140 42.9710 4.3380 52.2390 ;
      RECT 4.2660 42.9710 4.2900 52.2390 ;
      RECT 4.2180 42.9420 4.2420 52.2390 ;
      RECT 4.1700 42.8980 4.1940 52.2400 ;
      RECT 4.1220 42.8610 4.1460 52.2410 ;
      RECT 4.0740 42.8010 4.0980 52.2410 ;
      RECT 3.9840 47.7520 4.0080 47.8940 ;
      RECT 3.8170 43.4810 3.8410 47.3250 ;
      RECT 3.4440 45.0640 3.4680 45.3020 ;
  LAYER M2  ;
    RECT 0.108 0.036 9.5040 95.0040 ;
  LAYER M1  ;
    RECT 0.108 0.036 9.5040 95.0040 ;
  END
END srambank_64x4x80_6t122 
