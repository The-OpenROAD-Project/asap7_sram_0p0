VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_128x4x48_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_128x4x48_6t122 0 0 ; 
  SIZE 64 BY 241.92 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.688 65.768 4.88 ; 
        RECT 0.376 9.008 65.768 9.2 ; 
        RECT 0.376 13.328 65.768 13.52 ; 
        RECT 0.376 17.648 65.768 17.84 ; 
        RECT 0.376 21.968 65.768 22.16 ; 
        RECT 0.376 26.288 65.768 26.48 ; 
        RECT 0.376 30.608 65.768 30.8 ; 
        RECT 0.376 34.928 65.768 35.12 ; 
        RECT 0.376 39.248 65.768 39.44 ; 
        RECT 0.376 43.568 65.768 43.76 ; 
        RECT 0.376 47.888 65.768 48.08 ; 
        RECT 0.376 52.208 65.768 52.4 ; 
        RECT 0.376 56.528 65.768 56.72 ; 
        RECT 0.376 60.848 65.768 61.04 ; 
        RECT 0.376 65.168 65.768 65.36 ; 
        RECT 0.376 69.488 65.768 69.68 ; 
        RECT 0.376 73.808 65.768 74 ; 
        RECT 0.376 78.128 65.768 78.32 ; 
        RECT 0.376 82.448 65.768 82.64 ; 
        RECT 0.376 86.768 65.768 86.96 ; 
        RECT 0.376 91.088 65.768 91.28 ; 
        RECT 0.376 95.408 65.768 95.6 ; 
        RECT 0.376 99.728 65.768 99.92 ; 
        RECT 0.376 104.048 65.768 104.24 ; 
        RECT 14.256 105.972 51.84 106.836 ; 
        RECT 36.788 119.988 37.352 120.084 ; 
        RECT 36.264 104.852 37.316 104.948 ; 
        RECT 29.592 118.644 36.504 119.508 ; 
        RECT 29.592 131.316 36.504 132.18 ; 
        RECT 0.376 140.876 65.768 141.068 ; 
        RECT 0.376 145.196 65.768 145.388 ; 
        RECT 0.376 149.516 65.768 149.708 ; 
        RECT 0.376 153.836 65.768 154.028 ; 
        RECT 0.376 158.156 65.768 158.348 ; 
        RECT 0.376 162.476 65.768 162.668 ; 
        RECT 0.376 166.796 65.768 166.988 ; 
        RECT 0.376 171.116 65.768 171.308 ; 
        RECT 0.376 175.436 65.768 175.628 ; 
        RECT 0.376 179.756 65.768 179.948 ; 
        RECT 0.376 184.076 65.768 184.268 ; 
        RECT 0.376 188.396 65.768 188.588 ; 
        RECT 0.376 192.716 65.768 192.908 ; 
        RECT 0.376 197.036 65.768 197.228 ; 
        RECT 0.376 201.356 65.768 201.548 ; 
        RECT 0.376 205.676 65.768 205.868 ; 
        RECT 0.376 209.996 65.768 210.188 ; 
        RECT 0.376 214.316 65.768 214.508 ; 
        RECT 0.376 218.636 65.768 218.828 ; 
        RECT 0.376 222.956 65.768 223.148 ; 
        RECT 0.376 227.276 65.768 227.468 ; 
        RECT 0.376 231.596 65.768 231.788 ; 
        RECT 0.376 235.916 65.768 236.108 ; 
        RECT 0.376 240.236 65.768 240.428 ; 
      LAYER M3 ; 
        RECT 65.576 0.866 65.648 5.506 ; 
        RECT 37.136 0.868 37.208 5.504 ; 
        RECT 31.52 1.028 31.88 5.484 ; 
        RECT 28.928 0.868 29 5.504 ; 
        RECT 0.488 0.866 0.56 5.506 ; 
        RECT 65.576 5.186 65.648 9.826 ; 
        RECT 37.136 5.188 37.208 9.824 ; 
        RECT 31.52 5.348 31.88 9.804 ; 
        RECT 28.928 5.188 29 9.824 ; 
        RECT 0.488 5.186 0.56 9.826 ; 
        RECT 65.576 9.506 65.648 14.146 ; 
        RECT 37.136 9.508 37.208 14.144 ; 
        RECT 31.52 9.668 31.88 14.124 ; 
        RECT 28.928 9.508 29 14.144 ; 
        RECT 0.488 9.506 0.56 14.146 ; 
        RECT 65.576 13.826 65.648 18.466 ; 
        RECT 37.136 13.828 37.208 18.464 ; 
        RECT 31.52 13.988 31.88 18.444 ; 
        RECT 28.928 13.828 29 18.464 ; 
        RECT 0.488 13.826 0.56 18.466 ; 
        RECT 65.576 18.146 65.648 22.786 ; 
        RECT 37.136 18.148 37.208 22.784 ; 
        RECT 31.52 18.308 31.88 22.764 ; 
        RECT 28.928 18.148 29 22.784 ; 
        RECT 0.488 18.146 0.56 22.786 ; 
        RECT 65.576 22.466 65.648 27.106 ; 
        RECT 37.136 22.468 37.208 27.104 ; 
        RECT 31.52 22.628 31.88 27.084 ; 
        RECT 28.928 22.468 29 27.104 ; 
        RECT 0.488 22.466 0.56 27.106 ; 
        RECT 65.576 26.786 65.648 31.426 ; 
        RECT 37.136 26.788 37.208 31.424 ; 
        RECT 31.52 26.948 31.88 31.404 ; 
        RECT 28.928 26.788 29 31.424 ; 
        RECT 0.488 26.786 0.56 31.426 ; 
        RECT 65.576 31.106 65.648 35.746 ; 
        RECT 37.136 31.108 37.208 35.744 ; 
        RECT 31.52 31.268 31.88 35.724 ; 
        RECT 28.928 31.108 29 35.744 ; 
        RECT 0.488 31.106 0.56 35.746 ; 
        RECT 65.576 35.426 65.648 40.066 ; 
        RECT 37.136 35.428 37.208 40.064 ; 
        RECT 31.52 35.588 31.88 40.044 ; 
        RECT 28.928 35.428 29 40.064 ; 
        RECT 0.488 35.426 0.56 40.066 ; 
        RECT 65.576 39.746 65.648 44.386 ; 
        RECT 37.136 39.748 37.208 44.384 ; 
        RECT 31.52 39.908 31.88 44.364 ; 
        RECT 28.928 39.748 29 44.384 ; 
        RECT 0.488 39.746 0.56 44.386 ; 
        RECT 65.576 44.066 65.648 48.706 ; 
        RECT 37.136 44.068 37.208 48.704 ; 
        RECT 31.52 44.228 31.88 48.684 ; 
        RECT 28.928 44.068 29 48.704 ; 
        RECT 0.488 44.066 0.56 48.706 ; 
        RECT 65.576 48.386 65.648 53.026 ; 
        RECT 37.136 48.388 37.208 53.024 ; 
        RECT 31.52 48.548 31.88 53.004 ; 
        RECT 28.928 48.388 29 53.024 ; 
        RECT 0.488 48.386 0.56 53.026 ; 
        RECT 65.576 52.706 65.648 57.346 ; 
        RECT 37.136 52.708 37.208 57.344 ; 
        RECT 31.52 52.868 31.88 57.324 ; 
        RECT 28.928 52.708 29 57.344 ; 
        RECT 0.488 52.706 0.56 57.346 ; 
        RECT 65.576 57.026 65.648 61.666 ; 
        RECT 37.136 57.028 37.208 61.664 ; 
        RECT 31.52 57.188 31.88 61.644 ; 
        RECT 28.928 57.028 29 61.664 ; 
        RECT 0.488 57.026 0.56 61.666 ; 
        RECT 65.576 61.346 65.648 65.986 ; 
        RECT 37.136 61.348 37.208 65.984 ; 
        RECT 31.52 61.508 31.88 65.964 ; 
        RECT 28.928 61.348 29 65.984 ; 
        RECT 0.488 61.346 0.56 65.986 ; 
        RECT 65.576 65.666 65.648 70.306 ; 
        RECT 37.136 65.668 37.208 70.304 ; 
        RECT 31.52 65.828 31.88 70.284 ; 
        RECT 28.928 65.668 29 70.304 ; 
        RECT 0.488 65.666 0.56 70.306 ; 
        RECT 65.576 69.986 65.648 74.626 ; 
        RECT 37.136 69.988 37.208 74.624 ; 
        RECT 31.52 70.148 31.88 74.604 ; 
        RECT 28.928 69.988 29 74.624 ; 
        RECT 0.488 69.986 0.56 74.626 ; 
        RECT 65.576 74.306 65.648 78.946 ; 
        RECT 37.136 74.308 37.208 78.944 ; 
        RECT 31.52 74.468 31.88 78.924 ; 
        RECT 28.928 74.308 29 78.944 ; 
        RECT 0.488 74.306 0.56 78.946 ; 
        RECT 65.576 78.626 65.648 83.266 ; 
        RECT 37.136 78.628 37.208 83.264 ; 
        RECT 31.52 78.788 31.88 83.244 ; 
        RECT 28.928 78.628 29 83.264 ; 
        RECT 0.488 78.626 0.56 83.266 ; 
        RECT 65.576 82.946 65.648 87.586 ; 
        RECT 37.136 82.948 37.208 87.584 ; 
        RECT 31.52 83.108 31.88 87.564 ; 
        RECT 28.928 82.948 29 87.584 ; 
        RECT 0.488 82.946 0.56 87.586 ; 
        RECT 65.576 87.266 65.648 91.906 ; 
        RECT 37.136 87.268 37.208 91.904 ; 
        RECT 31.52 87.428 31.88 91.884 ; 
        RECT 28.928 87.268 29 91.904 ; 
        RECT 0.488 87.266 0.56 91.906 ; 
        RECT 65.576 91.586 65.648 96.226 ; 
        RECT 37.136 91.588 37.208 96.224 ; 
        RECT 31.52 91.748 31.88 96.204 ; 
        RECT 28.928 91.588 29 96.224 ; 
        RECT 0.488 91.586 0.56 96.226 ; 
        RECT 65.576 95.906 65.648 100.546 ; 
        RECT 37.136 95.908 37.208 100.544 ; 
        RECT 31.52 96.068 31.88 100.524 ; 
        RECT 28.928 95.908 29 100.544 ; 
        RECT 0.488 95.906 0.56 100.546 ; 
        RECT 65.576 100.226 65.648 104.866 ; 
        RECT 37.136 100.228 37.208 104.864 ; 
        RECT 31.52 100.388 31.88 104.844 ; 
        RECT 28.928 100.228 29 104.864 ; 
        RECT 0.488 100.226 0.56 104.866 ; 
        RECT 65.556 104.522 65.628 137.35 ; 
        RECT 37.188 119.8 37.26 137.194 ; 
        RECT 37.116 104.654 37.188 105.206 ; 
        RECT 31.644 105.816 32.58 136.148 ; 
        RECT 31.5 135.816 31.86 137.32 ; 
        RECT 31.5 104.68 31.86 106.184 ; 
        RECT 0.468 104.522 0.54 137.35 ; 
        RECT 65.576 137.054 65.648 141.694 ; 
        RECT 37.136 137.056 37.208 141.692 ; 
        RECT 31.52 137.216 31.88 141.672 ; 
        RECT 28.928 137.056 29 141.692 ; 
        RECT 0.488 137.054 0.56 141.694 ; 
        RECT 65.576 141.374 65.648 146.014 ; 
        RECT 37.136 141.376 37.208 146.012 ; 
        RECT 31.52 141.536 31.88 145.992 ; 
        RECT 28.928 141.376 29 146.012 ; 
        RECT 0.488 141.374 0.56 146.014 ; 
        RECT 65.576 145.694 65.648 150.334 ; 
        RECT 37.136 145.696 37.208 150.332 ; 
        RECT 31.52 145.856 31.88 150.312 ; 
        RECT 28.928 145.696 29 150.332 ; 
        RECT 0.488 145.694 0.56 150.334 ; 
        RECT 65.576 150.014 65.648 154.654 ; 
        RECT 37.136 150.016 37.208 154.652 ; 
        RECT 31.52 150.176 31.88 154.632 ; 
        RECT 28.928 150.016 29 154.652 ; 
        RECT 0.488 150.014 0.56 154.654 ; 
        RECT 65.576 154.334 65.648 158.974 ; 
        RECT 37.136 154.336 37.208 158.972 ; 
        RECT 31.52 154.496 31.88 158.952 ; 
        RECT 28.928 154.336 29 158.972 ; 
        RECT 0.488 154.334 0.56 158.974 ; 
        RECT 65.576 158.654 65.648 163.294 ; 
        RECT 37.136 158.656 37.208 163.292 ; 
        RECT 31.52 158.816 31.88 163.272 ; 
        RECT 28.928 158.656 29 163.292 ; 
        RECT 0.488 158.654 0.56 163.294 ; 
        RECT 65.576 162.974 65.648 167.614 ; 
        RECT 37.136 162.976 37.208 167.612 ; 
        RECT 31.52 163.136 31.88 167.592 ; 
        RECT 28.928 162.976 29 167.612 ; 
        RECT 0.488 162.974 0.56 167.614 ; 
        RECT 65.576 167.294 65.648 171.934 ; 
        RECT 37.136 167.296 37.208 171.932 ; 
        RECT 31.52 167.456 31.88 171.912 ; 
        RECT 28.928 167.296 29 171.932 ; 
        RECT 0.488 167.294 0.56 171.934 ; 
        RECT 65.576 171.614 65.648 176.254 ; 
        RECT 37.136 171.616 37.208 176.252 ; 
        RECT 31.52 171.776 31.88 176.232 ; 
        RECT 28.928 171.616 29 176.252 ; 
        RECT 0.488 171.614 0.56 176.254 ; 
        RECT 65.576 175.934 65.648 180.574 ; 
        RECT 37.136 175.936 37.208 180.572 ; 
        RECT 31.52 176.096 31.88 180.552 ; 
        RECT 28.928 175.936 29 180.572 ; 
        RECT 0.488 175.934 0.56 180.574 ; 
        RECT 65.576 180.254 65.648 184.894 ; 
        RECT 37.136 180.256 37.208 184.892 ; 
        RECT 31.52 180.416 31.88 184.872 ; 
        RECT 28.928 180.256 29 184.892 ; 
        RECT 0.488 180.254 0.56 184.894 ; 
        RECT 65.576 184.574 65.648 189.214 ; 
        RECT 37.136 184.576 37.208 189.212 ; 
        RECT 31.52 184.736 31.88 189.192 ; 
        RECT 28.928 184.576 29 189.212 ; 
        RECT 0.488 184.574 0.56 189.214 ; 
        RECT 65.576 188.894 65.648 193.534 ; 
        RECT 37.136 188.896 37.208 193.532 ; 
        RECT 31.52 189.056 31.88 193.512 ; 
        RECT 28.928 188.896 29 193.532 ; 
        RECT 0.488 188.894 0.56 193.534 ; 
        RECT 65.576 193.214 65.648 197.854 ; 
        RECT 37.136 193.216 37.208 197.852 ; 
        RECT 31.52 193.376 31.88 197.832 ; 
        RECT 28.928 193.216 29 197.852 ; 
        RECT 0.488 193.214 0.56 197.854 ; 
        RECT 65.576 197.534 65.648 202.174 ; 
        RECT 37.136 197.536 37.208 202.172 ; 
        RECT 31.52 197.696 31.88 202.152 ; 
        RECT 28.928 197.536 29 202.172 ; 
        RECT 0.488 197.534 0.56 202.174 ; 
        RECT 65.576 201.854 65.648 206.494 ; 
        RECT 37.136 201.856 37.208 206.492 ; 
        RECT 31.52 202.016 31.88 206.472 ; 
        RECT 28.928 201.856 29 206.492 ; 
        RECT 0.488 201.854 0.56 206.494 ; 
        RECT 65.576 206.174 65.648 210.814 ; 
        RECT 37.136 206.176 37.208 210.812 ; 
        RECT 31.52 206.336 31.88 210.792 ; 
        RECT 28.928 206.176 29 210.812 ; 
        RECT 0.488 206.174 0.56 210.814 ; 
        RECT 65.576 210.494 65.648 215.134 ; 
        RECT 37.136 210.496 37.208 215.132 ; 
        RECT 31.52 210.656 31.88 215.112 ; 
        RECT 28.928 210.496 29 215.132 ; 
        RECT 0.488 210.494 0.56 215.134 ; 
        RECT 65.576 214.814 65.648 219.454 ; 
        RECT 37.136 214.816 37.208 219.452 ; 
        RECT 31.52 214.976 31.88 219.432 ; 
        RECT 28.928 214.816 29 219.452 ; 
        RECT 0.488 214.814 0.56 219.454 ; 
        RECT 65.576 219.134 65.648 223.774 ; 
        RECT 37.136 219.136 37.208 223.772 ; 
        RECT 31.52 219.296 31.88 223.752 ; 
        RECT 28.928 219.136 29 223.772 ; 
        RECT 0.488 219.134 0.56 223.774 ; 
        RECT 65.576 223.454 65.648 228.094 ; 
        RECT 37.136 223.456 37.208 228.092 ; 
        RECT 31.52 223.616 31.88 228.072 ; 
        RECT 28.928 223.456 29 228.092 ; 
        RECT 0.488 223.454 0.56 228.094 ; 
        RECT 65.576 227.774 65.648 232.414 ; 
        RECT 37.136 227.776 37.208 232.412 ; 
        RECT 31.52 227.936 31.88 232.392 ; 
        RECT 28.928 227.776 29 232.412 ; 
        RECT 0.488 227.774 0.56 232.414 ; 
        RECT 65.576 232.094 65.648 236.734 ; 
        RECT 37.136 232.096 37.208 236.732 ; 
        RECT 31.52 232.256 31.88 236.712 ; 
        RECT 28.928 232.096 29 236.732 ; 
        RECT 0.488 232.094 0.56 236.734 ; 
        RECT 65.576 236.414 65.648 241.054 ; 
        RECT 37.136 236.416 37.208 241.052 ; 
        RECT 31.52 236.576 31.88 241.032 ; 
        RECT 28.928 236.416 29 241.052 ; 
        RECT 0.488 236.414 0.56 241.054 ; 
      LAYER V3 ; 
        RECT 0.488 4.688 0.56 4.88 ; 
        RECT 28.928 4.688 29 4.88 ; 
        RECT 31.52 4.688 31.88 4.88 ; 
        RECT 37.136 4.688 37.208 4.88 ; 
        RECT 65.576 4.688 65.648 4.88 ; 
        RECT 0.488 9.008 0.56 9.2 ; 
        RECT 28.928 9.008 29 9.2 ; 
        RECT 31.52 9.008 31.88 9.2 ; 
        RECT 37.136 9.008 37.208 9.2 ; 
        RECT 65.576 9.008 65.648 9.2 ; 
        RECT 0.488 13.328 0.56 13.52 ; 
        RECT 28.928 13.328 29 13.52 ; 
        RECT 31.52 13.328 31.88 13.52 ; 
        RECT 37.136 13.328 37.208 13.52 ; 
        RECT 65.576 13.328 65.648 13.52 ; 
        RECT 0.488 17.648 0.56 17.84 ; 
        RECT 28.928 17.648 29 17.84 ; 
        RECT 31.52 17.648 31.88 17.84 ; 
        RECT 37.136 17.648 37.208 17.84 ; 
        RECT 65.576 17.648 65.648 17.84 ; 
        RECT 0.488 21.968 0.56 22.16 ; 
        RECT 28.928 21.968 29 22.16 ; 
        RECT 31.52 21.968 31.88 22.16 ; 
        RECT 37.136 21.968 37.208 22.16 ; 
        RECT 65.576 21.968 65.648 22.16 ; 
        RECT 0.488 26.288 0.56 26.48 ; 
        RECT 28.928 26.288 29 26.48 ; 
        RECT 31.52 26.288 31.88 26.48 ; 
        RECT 37.136 26.288 37.208 26.48 ; 
        RECT 65.576 26.288 65.648 26.48 ; 
        RECT 0.488 30.608 0.56 30.8 ; 
        RECT 28.928 30.608 29 30.8 ; 
        RECT 31.52 30.608 31.88 30.8 ; 
        RECT 37.136 30.608 37.208 30.8 ; 
        RECT 65.576 30.608 65.648 30.8 ; 
        RECT 0.488 34.928 0.56 35.12 ; 
        RECT 28.928 34.928 29 35.12 ; 
        RECT 31.52 34.928 31.88 35.12 ; 
        RECT 37.136 34.928 37.208 35.12 ; 
        RECT 65.576 34.928 65.648 35.12 ; 
        RECT 0.488 39.248 0.56 39.44 ; 
        RECT 28.928 39.248 29 39.44 ; 
        RECT 31.52 39.248 31.88 39.44 ; 
        RECT 37.136 39.248 37.208 39.44 ; 
        RECT 65.576 39.248 65.648 39.44 ; 
        RECT 0.488 43.568 0.56 43.76 ; 
        RECT 28.928 43.568 29 43.76 ; 
        RECT 31.52 43.568 31.88 43.76 ; 
        RECT 37.136 43.568 37.208 43.76 ; 
        RECT 65.576 43.568 65.648 43.76 ; 
        RECT 0.488 47.888 0.56 48.08 ; 
        RECT 28.928 47.888 29 48.08 ; 
        RECT 31.52 47.888 31.88 48.08 ; 
        RECT 37.136 47.888 37.208 48.08 ; 
        RECT 65.576 47.888 65.648 48.08 ; 
        RECT 0.488 52.208 0.56 52.4 ; 
        RECT 28.928 52.208 29 52.4 ; 
        RECT 31.52 52.208 31.88 52.4 ; 
        RECT 37.136 52.208 37.208 52.4 ; 
        RECT 65.576 52.208 65.648 52.4 ; 
        RECT 0.488 56.528 0.56 56.72 ; 
        RECT 28.928 56.528 29 56.72 ; 
        RECT 31.52 56.528 31.88 56.72 ; 
        RECT 37.136 56.528 37.208 56.72 ; 
        RECT 65.576 56.528 65.648 56.72 ; 
        RECT 0.488 60.848 0.56 61.04 ; 
        RECT 28.928 60.848 29 61.04 ; 
        RECT 31.52 60.848 31.88 61.04 ; 
        RECT 37.136 60.848 37.208 61.04 ; 
        RECT 65.576 60.848 65.648 61.04 ; 
        RECT 0.488 65.168 0.56 65.36 ; 
        RECT 28.928 65.168 29 65.36 ; 
        RECT 31.52 65.168 31.88 65.36 ; 
        RECT 37.136 65.168 37.208 65.36 ; 
        RECT 65.576 65.168 65.648 65.36 ; 
        RECT 0.488 69.488 0.56 69.68 ; 
        RECT 28.928 69.488 29 69.68 ; 
        RECT 31.52 69.488 31.88 69.68 ; 
        RECT 37.136 69.488 37.208 69.68 ; 
        RECT 65.576 69.488 65.648 69.68 ; 
        RECT 0.488 73.808 0.56 74 ; 
        RECT 28.928 73.808 29 74 ; 
        RECT 31.52 73.808 31.88 74 ; 
        RECT 37.136 73.808 37.208 74 ; 
        RECT 65.576 73.808 65.648 74 ; 
        RECT 0.488 78.128 0.56 78.32 ; 
        RECT 28.928 78.128 29 78.32 ; 
        RECT 31.52 78.128 31.88 78.32 ; 
        RECT 37.136 78.128 37.208 78.32 ; 
        RECT 65.576 78.128 65.648 78.32 ; 
        RECT 0.488 82.448 0.56 82.64 ; 
        RECT 28.928 82.448 29 82.64 ; 
        RECT 31.52 82.448 31.88 82.64 ; 
        RECT 37.136 82.448 37.208 82.64 ; 
        RECT 65.576 82.448 65.648 82.64 ; 
        RECT 0.488 86.768 0.56 86.96 ; 
        RECT 28.928 86.768 29 86.96 ; 
        RECT 31.52 86.768 31.88 86.96 ; 
        RECT 37.136 86.768 37.208 86.96 ; 
        RECT 65.576 86.768 65.648 86.96 ; 
        RECT 0.488 91.088 0.56 91.28 ; 
        RECT 28.928 91.088 29 91.28 ; 
        RECT 31.52 91.088 31.88 91.28 ; 
        RECT 37.136 91.088 37.208 91.28 ; 
        RECT 65.576 91.088 65.648 91.28 ; 
        RECT 0.488 95.408 0.56 95.6 ; 
        RECT 28.928 95.408 29 95.6 ; 
        RECT 31.52 95.408 31.88 95.6 ; 
        RECT 37.136 95.408 37.208 95.6 ; 
        RECT 65.576 95.408 65.648 95.6 ; 
        RECT 0.488 99.728 0.56 99.92 ; 
        RECT 28.928 99.728 29 99.92 ; 
        RECT 31.52 99.728 31.88 99.92 ; 
        RECT 37.136 99.728 37.208 99.92 ; 
        RECT 65.576 99.728 65.648 99.92 ; 
        RECT 0.488 104.048 0.56 104.24 ; 
        RECT 28.928 104.048 29 104.24 ; 
        RECT 31.52 104.048 31.88 104.24 ; 
        RECT 37.136 104.048 37.208 104.24 ; 
        RECT 65.576 104.048 65.648 104.24 ; 
        RECT 31.66 131.316 31.732 132.18 ; 
        RECT 31.66 118.644 31.732 119.508 ; 
        RECT 31.66 105.972 31.732 106.836 ; 
        RECT 31.868 131.316 31.94 132.18 ; 
        RECT 31.868 118.644 31.94 119.508 ; 
        RECT 31.868 105.972 31.94 106.836 ; 
        RECT 32.076 131.316 32.148 132.18 ; 
        RECT 32.076 118.644 32.148 119.508 ; 
        RECT 32.076 105.972 32.148 106.836 ; 
        RECT 32.284 131.316 32.356 132.18 ; 
        RECT 32.284 118.644 32.356 119.508 ; 
        RECT 32.284 105.972 32.356 106.836 ; 
        RECT 32.492 131.316 32.564 132.18 ; 
        RECT 32.492 118.644 32.564 119.508 ; 
        RECT 32.492 105.972 32.564 106.836 ; 
        RECT 37.116 104.852 37.188 104.948 ; 
        RECT 37.188 119.988 37.26 120.084 ; 
        RECT 0.488 140.876 0.56 141.068 ; 
        RECT 28.928 140.876 29 141.068 ; 
        RECT 31.52 140.876 31.88 141.068 ; 
        RECT 37.136 140.876 37.208 141.068 ; 
        RECT 65.576 140.876 65.648 141.068 ; 
        RECT 0.488 145.196 0.56 145.388 ; 
        RECT 28.928 145.196 29 145.388 ; 
        RECT 31.52 145.196 31.88 145.388 ; 
        RECT 37.136 145.196 37.208 145.388 ; 
        RECT 65.576 145.196 65.648 145.388 ; 
        RECT 0.488 149.516 0.56 149.708 ; 
        RECT 28.928 149.516 29 149.708 ; 
        RECT 31.52 149.516 31.88 149.708 ; 
        RECT 37.136 149.516 37.208 149.708 ; 
        RECT 65.576 149.516 65.648 149.708 ; 
        RECT 0.488 153.836 0.56 154.028 ; 
        RECT 28.928 153.836 29 154.028 ; 
        RECT 31.52 153.836 31.88 154.028 ; 
        RECT 37.136 153.836 37.208 154.028 ; 
        RECT 65.576 153.836 65.648 154.028 ; 
        RECT 0.488 158.156 0.56 158.348 ; 
        RECT 28.928 158.156 29 158.348 ; 
        RECT 31.52 158.156 31.88 158.348 ; 
        RECT 37.136 158.156 37.208 158.348 ; 
        RECT 65.576 158.156 65.648 158.348 ; 
        RECT 0.488 162.476 0.56 162.668 ; 
        RECT 28.928 162.476 29 162.668 ; 
        RECT 31.52 162.476 31.88 162.668 ; 
        RECT 37.136 162.476 37.208 162.668 ; 
        RECT 65.576 162.476 65.648 162.668 ; 
        RECT 0.488 166.796 0.56 166.988 ; 
        RECT 28.928 166.796 29 166.988 ; 
        RECT 31.52 166.796 31.88 166.988 ; 
        RECT 37.136 166.796 37.208 166.988 ; 
        RECT 65.576 166.796 65.648 166.988 ; 
        RECT 0.488 171.116 0.56 171.308 ; 
        RECT 28.928 171.116 29 171.308 ; 
        RECT 31.52 171.116 31.88 171.308 ; 
        RECT 37.136 171.116 37.208 171.308 ; 
        RECT 65.576 171.116 65.648 171.308 ; 
        RECT 0.488 175.436 0.56 175.628 ; 
        RECT 28.928 175.436 29 175.628 ; 
        RECT 31.52 175.436 31.88 175.628 ; 
        RECT 37.136 175.436 37.208 175.628 ; 
        RECT 65.576 175.436 65.648 175.628 ; 
        RECT 0.488 179.756 0.56 179.948 ; 
        RECT 28.928 179.756 29 179.948 ; 
        RECT 31.52 179.756 31.88 179.948 ; 
        RECT 37.136 179.756 37.208 179.948 ; 
        RECT 65.576 179.756 65.648 179.948 ; 
        RECT 0.488 184.076 0.56 184.268 ; 
        RECT 28.928 184.076 29 184.268 ; 
        RECT 31.52 184.076 31.88 184.268 ; 
        RECT 37.136 184.076 37.208 184.268 ; 
        RECT 65.576 184.076 65.648 184.268 ; 
        RECT 0.488 188.396 0.56 188.588 ; 
        RECT 28.928 188.396 29 188.588 ; 
        RECT 31.52 188.396 31.88 188.588 ; 
        RECT 37.136 188.396 37.208 188.588 ; 
        RECT 65.576 188.396 65.648 188.588 ; 
        RECT 0.488 192.716 0.56 192.908 ; 
        RECT 28.928 192.716 29 192.908 ; 
        RECT 31.52 192.716 31.88 192.908 ; 
        RECT 37.136 192.716 37.208 192.908 ; 
        RECT 65.576 192.716 65.648 192.908 ; 
        RECT 0.488 197.036 0.56 197.228 ; 
        RECT 28.928 197.036 29 197.228 ; 
        RECT 31.52 197.036 31.88 197.228 ; 
        RECT 37.136 197.036 37.208 197.228 ; 
        RECT 65.576 197.036 65.648 197.228 ; 
        RECT 0.488 201.356 0.56 201.548 ; 
        RECT 28.928 201.356 29 201.548 ; 
        RECT 31.52 201.356 31.88 201.548 ; 
        RECT 37.136 201.356 37.208 201.548 ; 
        RECT 65.576 201.356 65.648 201.548 ; 
        RECT 0.488 205.676 0.56 205.868 ; 
        RECT 28.928 205.676 29 205.868 ; 
        RECT 31.52 205.676 31.88 205.868 ; 
        RECT 37.136 205.676 37.208 205.868 ; 
        RECT 65.576 205.676 65.648 205.868 ; 
        RECT 0.488 209.996 0.56 210.188 ; 
        RECT 28.928 209.996 29 210.188 ; 
        RECT 31.52 209.996 31.88 210.188 ; 
        RECT 37.136 209.996 37.208 210.188 ; 
        RECT 65.576 209.996 65.648 210.188 ; 
        RECT 0.488 214.316 0.56 214.508 ; 
        RECT 28.928 214.316 29 214.508 ; 
        RECT 31.52 214.316 31.88 214.508 ; 
        RECT 37.136 214.316 37.208 214.508 ; 
        RECT 65.576 214.316 65.648 214.508 ; 
        RECT 0.488 218.636 0.56 218.828 ; 
        RECT 28.928 218.636 29 218.828 ; 
        RECT 31.52 218.636 31.88 218.828 ; 
        RECT 37.136 218.636 37.208 218.828 ; 
        RECT 65.576 218.636 65.648 218.828 ; 
        RECT 0.488 222.956 0.56 223.148 ; 
        RECT 28.928 222.956 29 223.148 ; 
        RECT 31.52 222.956 31.88 223.148 ; 
        RECT 37.136 222.956 37.208 223.148 ; 
        RECT 65.576 222.956 65.648 223.148 ; 
        RECT 0.488 227.276 0.56 227.468 ; 
        RECT 28.928 227.276 29 227.468 ; 
        RECT 31.52 227.276 31.88 227.468 ; 
        RECT 37.136 227.276 37.208 227.468 ; 
        RECT 65.576 227.276 65.648 227.468 ; 
        RECT 0.488 231.596 0.56 231.788 ; 
        RECT 28.928 231.596 29 231.788 ; 
        RECT 31.52 231.596 31.88 231.788 ; 
        RECT 37.136 231.596 37.208 231.788 ; 
        RECT 65.576 231.596 65.648 231.788 ; 
        RECT 0.488 235.916 0.56 236.108 ; 
        RECT 28.928 235.916 29 236.108 ; 
        RECT 31.52 235.916 31.88 236.108 ; 
        RECT 37.136 235.916 37.208 236.108 ; 
        RECT 65.576 235.916 65.648 236.108 ; 
        RECT 0.488 240.236 0.56 240.428 ; 
        RECT 28.928 240.236 29 240.428 ; 
        RECT 31.52 240.236 31.88 240.428 ; 
        RECT 37.136 240.236 37.208 240.428 ; 
        RECT 65.576 240.236 65.648 240.428 ; 
      LAYER M5 ; 
        RECT 36.864 104.78 36.96 120.156 ; 
      LAYER V4 ; 
        RECT 36.864 119.988 36.96 120.084 ; 
        RECT 36.864 105.972 36.96 106.836 ; 
        RECT 36.864 104.852 36.96 104.948 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.376 4.304 65.748 4.496 ; 
        RECT 0.376 8.624 65.748 8.816 ; 
        RECT 0.376 12.944 65.748 13.136 ; 
        RECT 0.376 17.264 65.748 17.456 ; 
        RECT 0.376 21.584 65.748 21.776 ; 
        RECT 0.376 25.904 65.748 26.096 ; 
        RECT 0.376 30.224 65.748 30.416 ; 
        RECT 0.376 34.544 65.748 34.736 ; 
        RECT 0.376 38.864 65.748 39.056 ; 
        RECT 0.376 43.184 65.748 43.376 ; 
        RECT 0.376 47.504 65.748 47.696 ; 
        RECT 0.376 51.824 65.748 52.016 ; 
        RECT 0.376 56.144 65.748 56.336 ; 
        RECT 0.376 60.464 65.748 60.656 ; 
        RECT 0.376 64.784 65.748 64.976 ; 
        RECT 0.376 69.104 65.748 69.296 ; 
        RECT 0.376 73.424 65.748 73.616 ; 
        RECT 0.376 77.744 65.748 77.936 ; 
        RECT 0.376 82.064 65.748 82.256 ; 
        RECT 0.376 86.384 65.748 86.576 ; 
        RECT 0.376 90.704 65.748 90.896 ; 
        RECT 0.376 95.024 65.748 95.216 ; 
        RECT 0.376 99.344 65.748 99.536 ; 
        RECT 0.376 103.664 65.748 103.856 ; 
        RECT 14.256 107.7 51.84 108.564 ; 
        RECT 29.592 120.372 36.504 121.236 ; 
        RECT 29.592 133.044 36.504 133.908 ; 
        RECT 0.376 140.492 65.748 140.684 ; 
        RECT 0.376 144.812 65.748 145.004 ; 
        RECT 0.376 149.132 65.748 149.324 ; 
        RECT 0.376 153.452 65.748 153.644 ; 
        RECT 0.376 157.772 65.748 157.964 ; 
        RECT 0.376 162.092 65.748 162.284 ; 
        RECT 0.376 166.412 65.748 166.604 ; 
        RECT 0.376 170.732 65.748 170.924 ; 
        RECT 0.376 175.052 65.748 175.244 ; 
        RECT 0.376 179.372 65.748 179.564 ; 
        RECT 0.376 183.692 65.748 183.884 ; 
        RECT 0.376 188.012 65.748 188.204 ; 
        RECT 0.376 192.332 65.748 192.524 ; 
        RECT 0.376 196.652 65.748 196.844 ; 
        RECT 0.376 200.972 65.748 201.164 ; 
        RECT 0.376 205.292 65.748 205.484 ; 
        RECT 0.376 209.612 65.748 209.804 ; 
        RECT 0.376 213.932 65.748 214.124 ; 
        RECT 0.376 218.252 65.748 218.444 ; 
        RECT 0.376 222.572 65.748 222.764 ; 
        RECT 0.376 226.892 65.748 227.084 ; 
        RECT 0.376 231.212 65.748 231.404 ; 
        RECT 0.376 235.532 65.748 235.724 ; 
        RECT 0.376 239.852 65.748 240.044 ; 
      LAYER M3 ; 
        RECT 65.432 0.866 65.504 5.506 ; 
        RECT 37.352 0.866 37.424 5.506 ; 
        RECT 34.292 1.012 34.436 5.468 ; 
        RECT 33.68 1.012 33.788 5.468 ; 
        RECT 28.712 0.866 28.784 5.506 ; 
        RECT 0.632 0.866 0.704 5.506 ; 
        RECT 65.432 5.186 65.504 9.826 ; 
        RECT 37.352 5.186 37.424 9.826 ; 
        RECT 34.292 5.332 34.436 9.788 ; 
        RECT 33.68 5.332 33.788 9.788 ; 
        RECT 28.712 5.186 28.784 9.826 ; 
        RECT 0.632 5.186 0.704 9.826 ; 
        RECT 65.432 9.506 65.504 14.146 ; 
        RECT 37.352 9.506 37.424 14.146 ; 
        RECT 34.292 9.652 34.436 14.108 ; 
        RECT 33.68 9.652 33.788 14.108 ; 
        RECT 28.712 9.506 28.784 14.146 ; 
        RECT 0.632 9.506 0.704 14.146 ; 
        RECT 65.432 13.826 65.504 18.466 ; 
        RECT 37.352 13.826 37.424 18.466 ; 
        RECT 34.292 13.972 34.436 18.428 ; 
        RECT 33.68 13.972 33.788 18.428 ; 
        RECT 28.712 13.826 28.784 18.466 ; 
        RECT 0.632 13.826 0.704 18.466 ; 
        RECT 65.432 18.146 65.504 22.786 ; 
        RECT 37.352 18.146 37.424 22.786 ; 
        RECT 34.292 18.292 34.436 22.748 ; 
        RECT 33.68 18.292 33.788 22.748 ; 
        RECT 28.712 18.146 28.784 22.786 ; 
        RECT 0.632 18.146 0.704 22.786 ; 
        RECT 65.432 22.466 65.504 27.106 ; 
        RECT 37.352 22.466 37.424 27.106 ; 
        RECT 34.292 22.612 34.436 27.068 ; 
        RECT 33.68 22.612 33.788 27.068 ; 
        RECT 28.712 22.466 28.784 27.106 ; 
        RECT 0.632 22.466 0.704 27.106 ; 
        RECT 65.432 26.786 65.504 31.426 ; 
        RECT 37.352 26.786 37.424 31.426 ; 
        RECT 34.292 26.932 34.436 31.388 ; 
        RECT 33.68 26.932 33.788 31.388 ; 
        RECT 28.712 26.786 28.784 31.426 ; 
        RECT 0.632 26.786 0.704 31.426 ; 
        RECT 65.432 31.106 65.504 35.746 ; 
        RECT 37.352 31.106 37.424 35.746 ; 
        RECT 34.292 31.252 34.436 35.708 ; 
        RECT 33.68 31.252 33.788 35.708 ; 
        RECT 28.712 31.106 28.784 35.746 ; 
        RECT 0.632 31.106 0.704 35.746 ; 
        RECT 65.432 35.426 65.504 40.066 ; 
        RECT 37.352 35.426 37.424 40.066 ; 
        RECT 34.292 35.572 34.436 40.028 ; 
        RECT 33.68 35.572 33.788 40.028 ; 
        RECT 28.712 35.426 28.784 40.066 ; 
        RECT 0.632 35.426 0.704 40.066 ; 
        RECT 65.432 39.746 65.504 44.386 ; 
        RECT 37.352 39.746 37.424 44.386 ; 
        RECT 34.292 39.892 34.436 44.348 ; 
        RECT 33.68 39.892 33.788 44.348 ; 
        RECT 28.712 39.746 28.784 44.386 ; 
        RECT 0.632 39.746 0.704 44.386 ; 
        RECT 65.432 44.066 65.504 48.706 ; 
        RECT 37.352 44.066 37.424 48.706 ; 
        RECT 34.292 44.212 34.436 48.668 ; 
        RECT 33.68 44.212 33.788 48.668 ; 
        RECT 28.712 44.066 28.784 48.706 ; 
        RECT 0.632 44.066 0.704 48.706 ; 
        RECT 65.432 48.386 65.504 53.026 ; 
        RECT 37.352 48.386 37.424 53.026 ; 
        RECT 34.292 48.532 34.436 52.988 ; 
        RECT 33.68 48.532 33.788 52.988 ; 
        RECT 28.712 48.386 28.784 53.026 ; 
        RECT 0.632 48.386 0.704 53.026 ; 
        RECT 65.432 52.706 65.504 57.346 ; 
        RECT 37.352 52.706 37.424 57.346 ; 
        RECT 34.292 52.852 34.436 57.308 ; 
        RECT 33.68 52.852 33.788 57.308 ; 
        RECT 28.712 52.706 28.784 57.346 ; 
        RECT 0.632 52.706 0.704 57.346 ; 
        RECT 65.432 57.026 65.504 61.666 ; 
        RECT 37.352 57.026 37.424 61.666 ; 
        RECT 34.292 57.172 34.436 61.628 ; 
        RECT 33.68 57.172 33.788 61.628 ; 
        RECT 28.712 57.026 28.784 61.666 ; 
        RECT 0.632 57.026 0.704 61.666 ; 
        RECT 65.432 61.346 65.504 65.986 ; 
        RECT 37.352 61.346 37.424 65.986 ; 
        RECT 34.292 61.492 34.436 65.948 ; 
        RECT 33.68 61.492 33.788 65.948 ; 
        RECT 28.712 61.346 28.784 65.986 ; 
        RECT 0.632 61.346 0.704 65.986 ; 
        RECT 65.432 65.666 65.504 70.306 ; 
        RECT 37.352 65.666 37.424 70.306 ; 
        RECT 34.292 65.812 34.436 70.268 ; 
        RECT 33.68 65.812 33.788 70.268 ; 
        RECT 28.712 65.666 28.784 70.306 ; 
        RECT 0.632 65.666 0.704 70.306 ; 
        RECT 65.432 69.986 65.504 74.626 ; 
        RECT 37.352 69.986 37.424 74.626 ; 
        RECT 34.292 70.132 34.436 74.588 ; 
        RECT 33.68 70.132 33.788 74.588 ; 
        RECT 28.712 69.986 28.784 74.626 ; 
        RECT 0.632 69.986 0.704 74.626 ; 
        RECT 65.432 74.306 65.504 78.946 ; 
        RECT 37.352 74.306 37.424 78.946 ; 
        RECT 34.292 74.452 34.436 78.908 ; 
        RECT 33.68 74.452 33.788 78.908 ; 
        RECT 28.712 74.306 28.784 78.946 ; 
        RECT 0.632 74.306 0.704 78.946 ; 
        RECT 65.432 78.626 65.504 83.266 ; 
        RECT 37.352 78.626 37.424 83.266 ; 
        RECT 34.292 78.772 34.436 83.228 ; 
        RECT 33.68 78.772 33.788 83.228 ; 
        RECT 28.712 78.626 28.784 83.266 ; 
        RECT 0.632 78.626 0.704 83.266 ; 
        RECT 65.432 82.946 65.504 87.586 ; 
        RECT 37.352 82.946 37.424 87.586 ; 
        RECT 34.292 83.092 34.436 87.548 ; 
        RECT 33.68 83.092 33.788 87.548 ; 
        RECT 28.712 82.946 28.784 87.586 ; 
        RECT 0.632 82.946 0.704 87.586 ; 
        RECT 65.432 87.266 65.504 91.906 ; 
        RECT 37.352 87.266 37.424 91.906 ; 
        RECT 34.292 87.412 34.436 91.868 ; 
        RECT 33.68 87.412 33.788 91.868 ; 
        RECT 28.712 87.266 28.784 91.906 ; 
        RECT 0.632 87.266 0.704 91.906 ; 
        RECT 65.432 91.586 65.504 96.226 ; 
        RECT 37.352 91.586 37.424 96.226 ; 
        RECT 34.292 91.732 34.436 96.188 ; 
        RECT 33.68 91.732 33.788 96.188 ; 
        RECT 28.712 91.586 28.784 96.226 ; 
        RECT 0.632 91.586 0.704 96.226 ; 
        RECT 65.432 95.906 65.504 100.546 ; 
        RECT 37.352 95.906 37.424 100.546 ; 
        RECT 34.292 96.052 34.436 100.508 ; 
        RECT 33.68 96.052 33.788 100.508 ; 
        RECT 28.712 95.906 28.784 100.546 ; 
        RECT 0.632 95.906 0.704 100.546 ; 
        RECT 65.432 100.226 65.504 104.866 ; 
        RECT 37.352 100.226 37.424 104.866 ; 
        RECT 34.292 100.372 34.436 104.828 ; 
        RECT 33.68 100.372 33.788 104.828 ; 
        RECT 28.712 100.226 28.784 104.866 ; 
        RECT 0.632 100.226 0.704 104.866 ; 
        RECT 65.412 104.522 65.484 137.35 ; 
        RECT 37.332 104.522 37.404 137.35 ; 
        RECT 33.516 105.416 34.452 136.148 ; 
        RECT 34.272 104.698 34.416 137.176 ; 
        RECT 33.66 104.696 33.768 137.176 ; 
        RECT 28.692 104.522 28.764 137.35 ; 
        RECT 0.612 104.522 0.684 137.35 ; 
        RECT 65.432 137.054 65.504 141.694 ; 
        RECT 37.352 137.054 37.424 141.694 ; 
        RECT 34.292 137.2 34.436 141.656 ; 
        RECT 33.68 137.2 33.788 141.656 ; 
        RECT 28.712 137.054 28.784 141.694 ; 
        RECT 0.632 137.054 0.704 141.694 ; 
        RECT 65.432 141.374 65.504 146.014 ; 
        RECT 37.352 141.374 37.424 146.014 ; 
        RECT 34.292 141.52 34.436 145.976 ; 
        RECT 33.68 141.52 33.788 145.976 ; 
        RECT 28.712 141.374 28.784 146.014 ; 
        RECT 0.632 141.374 0.704 146.014 ; 
        RECT 65.432 145.694 65.504 150.334 ; 
        RECT 37.352 145.694 37.424 150.334 ; 
        RECT 34.292 145.84 34.436 150.296 ; 
        RECT 33.68 145.84 33.788 150.296 ; 
        RECT 28.712 145.694 28.784 150.334 ; 
        RECT 0.632 145.694 0.704 150.334 ; 
        RECT 65.432 150.014 65.504 154.654 ; 
        RECT 37.352 150.014 37.424 154.654 ; 
        RECT 34.292 150.16 34.436 154.616 ; 
        RECT 33.68 150.16 33.788 154.616 ; 
        RECT 28.712 150.014 28.784 154.654 ; 
        RECT 0.632 150.014 0.704 154.654 ; 
        RECT 65.432 154.334 65.504 158.974 ; 
        RECT 37.352 154.334 37.424 158.974 ; 
        RECT 34.292 154.48 34.436 158.936 ; 
        RECT 33.68 154.48 33.788 158.936 ; 
        RECT 28.712 154.334 28.784 158.974 ; 
        RECT 0.632 154.334 0.704 158.974 ; 
        RECT 65.432 158.654 65.504 163.294 ; 
        RECT 37.352 158.654 37.424 163.294 ; 
        RECT 34.292 158.8 34.436 163.256 ; 
        RECT 33.68 158.8 33.788 163.256 ; 
        RECT 28.712 158.654 28.784 163.294 ; 
        RECT 0.632 158.654 0.704 163.294 ; 
        RECT 65.432 162.974 65.504 167.614 ; 
        RECT 37.352 162.974 37.424 167.614 ; 
        RECT 34.292 163.12 34.436 167.576 ; 
        RECT 33.68 163.12 33.788 167.576 ; 
        RECT 28.712 162.974 28.784 167.614 ; 
        RECT 0.632 162.974 0.704 167.614 ; 
        RECT 65.432 167.294 65.504 171.934 ; 
        RECT 37.352 167.294 37.424 171.934 ; 
        RECT 34.292 167.44 34.436 171.896 ; 
        RECT 33.68 167.44 33.788 171.896 ; 
        RECT 28.712 167.294 28.784 171.934 ; 
        RECT 0.632 167.294 0.704 171.934 ; 
        RECT 65.432 171.614 65.504 176.254 ; 
        RECT 37.352 171.614 37.424 176.254 ; 
        RECT 34.292 171.76 34.436 176.216 ; 
        RECT 33.68 171.76 33.788 176.216 ; 
        RECT 28.712 171.614 28.784 176.254 ; 
        RECT 0.632 171.614 0.704 176.254 ; 
        RECT 65.432 175.934 65.504 180.574 ; 
        RECT 37.352 175.934 37.424 180.574 ; 
        RECT 34.292 176.08 34.436 180.536 ; 
        RECT 33.68 176.08 33.788 180.536 ; 
        RECT 28.712 175.934 28.784 180.574 ; 
        RECT 0.632 175.934 0.704 180.574 ; 
        RECT 65.432 180.254 65.504 184.894 ; 
        RECT 37.352 180.254 37.424 184.894 ; 
        RECT 34.292 180.4 34.436 184.856 ; 
        RECT 33.68 180.4 33.788 184.856 ; 
        RECT 28.712 180.254 28.784 184.894 ; 
        RECT 0.632 180.254 0.704 184.894 ; 
        RECT 65.432 184.574 65.504 189.214 ; 
        RECT 37.352 184.574 37.424 189.214 ; 
        RECT 34.292 184.72 34.436 189.176 ; 
        RECT 33.68 184.72 33.788 189.176 ; 
        RECT 28.712 184.574 28.784 189.214 ; 
        RECT 0.632 184.574 0.704 189.214 ; 
        RECT 65.432 188.894 65.504 193.534 ; 
        RECT 37.352 188.894 37.424 193.534 ; 
        RECT 34.292 189.04 34.436 193.496 ; 
        RECT 33.68 189.04 33.788 193.496 ; 
        RECT 28.712 188.894 28.784 193.534 ; 
        RECT 0.632 188.894 0.704 193.534 ; 
        RECT 65.432 193.214 65.504 197.854 ; 
        RECT 37.352 193.214 37.424 197.854 ; 
        RECT 34.292 193.36 34.436 197.816 ; 
        RECT 33.68 193.36 33.788 197.816 ; 
        RECT 28.712 193.214 28.784 197.854 ; 
        RECT 0.632 193.214 0.704 197.854 ; 
        RECT 65.432 197.534 65.504 202.174 ; 
        RECT 37.352 197.534 37.424 202.174 ; 
        RECT 34.292 197.68 34.436 202.136 ; 
        RECT 33.68 197.68 33.788 202.136 ; 
        RECT 28.712 197.534 28.784 202.174 ; 
        RECT 0.632 197.534 0.704 202.174 ; 
        RECT 65.432 201.854 65.504 206.494 ; 
        RECT 37.352 201.854 37.424 206.494 ; 
        RECT 34.292 202 34.436 206.456 ; 
        RECT 33.68 202 33.788 206.456 ; 
        RECT 28.712 201.854 28.784 206.494 ; 
        RECT 0.632 201.854 0.704 206.494 ; 
        RECT 65.432 206.174 65.504 210.814 ; 
        RECT 37.352 206.174 37.424 210.814 ; 
        RECT 34.292 206.32 34.436 210.776 ; 
        RECT 33.68 206.32 33.788 210.776 ; 
        RECT 28.712 206.174 28.784 210.814 ; 
        RECT 0.632 206.174 0.704 210.814 ; 
        RECT 65.432 210.494 65.504 215.134 ; 
        RECT 37.352 210.494 37.424 215.134 ; 
        RECT 34.292 210.64 34.436 215.096 ; 
        RECT 33.68 210.64 33.788 215.096 ; 
        RECT 28.712 210.494 28.784 215.134 ; 
        RECT 0.632 210.494 0.704 215.134 ; 
        RECT 65.432 214.814 65.504 219.454 ; 
        RECT 37.352 214.814 37.424 219.454 ; 
        RECT 34.292 214.96 34.436 219.416 ; 
        RECT 33.68 214.96 33.788 219.416 ; 
        RECT 28.712 214.814 28.784 219.454 ; 
        RECT 0.632 214.814 0.704 219.454 ; 
        RECT 65.432 219.134 65.504 223.774 ; 
        RECT 37.352 219.134 37.424 223.774 ; 
        RECT 34.292 219.28 34.436 223.736 ; 
        RECT 33.68 219.28 33.788 223.736 ; 
        RECT 28.712 219.134 28.784 223.774 ; 
        RECT 0.632 219.134 0.704 223.774 ; 
        RECT 65.432 223.454 65.504 228.094 ; 
        RECT 37.352 223.454 37.424 228.094 ; 
        RECT 34.292 223.6 34.436 228.056 ; 
        RECT 33.68 223.6 33.788 228.056 ; 
        RECT 28.712 223.454 28.784 228.094 ; 
        RECT 0.632 223.454 0.704 228.094 ; 
        RECT 65.432 227.774 65.504 232.414 ; 
        RECT 37.352 227.774 37.424 232.414 ; 
        RECT 34.292 227.92 34.436 232.376 ; 
        RECT 33.68 227.92 33.788 232.376 ; 
        RECT 28.712 227.774 28.784 232.414 ; 
        RECT 0.632 227.774 0.704 232.414 ; 
        RECT 65.432 232.094 65.504 236.734 ; 
        RECT 37.352 232.094 37.424 236.734 ; 
        RECT 34.292 232.24 34.436 236.696 ; 
        RECT 33.68 232.24 33.788 236.696 ; 
        RECT 28.712 232.094 28.784 236.734 ; 
        RECT 0.632 232.094 0.704 236.734 ; 
        RECT 65.432 236.414 65.504 241.054 ; 
        RECT 37.352 236.414 37.424 241.054 ; 
        RECT 34.292 236.56 34.436 241.016 ; 
        RECT 33.68 236.56 33.788 241.016 ; 
        RECT 28.712 236.414 28.784 241.054 ; 
        RECT 0.632 236.414 0.704 241.054 ; 
      LAYER V3 ; 
        RECT 0.632 4.304 0.704 4.496 ; 
        RECT 28.712 4.304 28.784 4.496 ; 
        RECT 33.68 4.304 33.788 4.496 ; 
        RECT 34.292 4.304 34.436 4.496 ; 
        RECT 37.352 4.304 37.424 4.496 ; 
        RECT 65.432 4.304 65.504 4.496 ; 
        RECT 0.632 8.624 0.704 8.816 ; 
        RECT 28.712 8.624 28.784 8.816 ; 
        RECT 33.68 8.624 33.788 8.816 ; 
        RECT 34.292 8.624 34.436 8.816 ; 
        RECT 37.352 8.624 37.424 8.816 ; 
        RECT 65.432 8.624 65.504 8.816 ; 
        RECT 0.632 12.944 0.704 13.136 ; 
        RECT 28.712 12.944 28.784 13.136 ; 
        RECT 33.68 12.944 33.788 13.136 ; 
        RECT 34.292 12.944 34.436 13.136 ; 
        RECT 37.352 12.944 37.424 13.136 ; 
        RECT 65.432 12.944 65.504 13.136 ; 
        RECT 0.632 17.264 0.704 17.456 ; 
        RECT 28.712 17.264 28.784 17.456 ; 
        RECT 33.68 17.264 33.788 17.456 ; 
        RECT 34.292 17.264 34.436 17.456 ; 
        RECT 37.352 17.264 37.424 17.456 ; 
        RECT 65.432 17.264 65.504 17.456 ; 
        RECT 0.632 21.584 0.704 21.776 ; 
        RECT 28.712 21.584 28.784 21.776 ; 
        RECT 33.68 21.584 33.788 21.776 ; 
        RECT 34.292 21.584 34.436 21.776 ; 
        RECT 37.352 21.584 37.424 21.776 ; 
        RECT 65.432 21.584 65.504 21.776 ; 
        RECT 0.632 25.904 0.704 26.096 ; 
        RECT 28.712 25.904 28.784 26.096 ; 
        RECT 33.68 25.904 33.788 26.096 ; 
        RECT 34.292 25.904 34.436 26.096 ; 
        RECT 37.352 25.904 37.424 26.096 ; 
        RECT 65.432 25.904 65.504 26.096 ; 
        RECT 0.632 30.224 0.704 30.416 ; 
        RECT 28.712 30.224 28.784 30.416 ; 
        RECT 33.68 30.224 33.788 30.416 ; 
        RECT 34.292 30.224 34.436 30.416 ; 
        RECT 37.352 30.224 37.424 30.416 ; 
        RECT 65.432 30.224 65.504 30.416 ; 
        RECT 0.632 34.544 0.704 34.736 ; 
        RECT 28.712 34.544 28.784 34.736 ; 
        RECT 33.68 34.544 33.788 34.736 ; 
        RECT 34.292 34.544 34.436 34.736 ; 
        RECT 37.352 34.544 37.424 34.736 ; 
        RECT 65.432 34.544 65.504 34.736 ; 
        RECT 0.632 38.864 0.704 39.056 ; 
        RECT 28.712 38.864 28.784 39.056 ; 
        RECT 33.68 38.864 33.788 39.056 ; 
        RECT 34.292 38.864 34.436 39.056 ; 
        RECT 37.352 38.864 37.424 39.056 ; 
        RECT 65.432 38.864 65.504 39.056 ; 
        RECT 0.632 43.184 0.704 43.376 ; 
        RECT 28.712 43.184 28.784 43.376 ; 
        RECT 33.68 43.184 33.788 43.376 ; 
        RECT 34.292 43.184 34.436 43.376 ; 
        RECT 37.352 43.184 37.424 43.376 ; 
        RECT 65.432 43.184 65.504 43.376 ; 
        RECT 0.632 47.504 0.704 47.696 ; 
        RECT 28.712 47.504 28.784 47.696 ; 
        RECT 33.68 47.504 33.788 47.696 ; 
        RECT 34.292 47.504 34.436 47.696 ; 
        RECT 37.352 47.504 37.424 47.696 ; 
        RECT 65.432 47.504 65.504 47.696 ; 
        RECT 0.632 51.824 0.704 52.016 ; 
        RECT 28.712 51.824 28.784 52.016 ; 
        RECT 33.68 51.824 33.788 52.016 ; 
        RECT 34.292 51.824 34.436 52.016 ; 
        RECT 37.352 51.824 37.424 52.016 ; 
        RECT 65.432 51.824 65.504 52.016 ; 
        RECT 0.632 56.144 0.704 56.336 ; 
        RECT 28.712 56.144 28.784 56.336 ; 
        RECT 33.68 56.144 33.788 56.336 ; 
        RECT 34.292 56.144 34.436 56.336 ; 
        RECT 37.352 56.144 37.424 56.336 ; 
        RECT 65.432 56.144 65.504 56.336 ; 
        RECT 0.632 60.464 0.704 60.656 ; 
        RECT 28.712 60.464 28.784 60.656 ; 
        RECT 33.68 60.464 33.788 60.656 ; 
        RECT 34.292 60.464 34.436 60.656 ; 
        RECT 37.352 60.464 37.424 60.656 ; 
        RECT 65.432 60.464 65.504 60.656 ; 
        RECT 0.632 64.784 0.704 64.976 ; 
        RECT 28.712 64.784 28.784 64.976 ; 
        RECT 33.68 64.784 33.788 64.976 ; 
        RECT 34.292 64.784 34.436 64.976 ; 
        RECT 37.352 64.784 37.424 64.976 ; 
        RECT 65.432 64.784 65.504 64.976 ; 
        RECT 0.632 69.104 0.704 69.296 ; 
        RECT 28.712 69.104 28.784 69.296 ; 
        RECT 33.68 69.104 33.788 69.296 ; 
        RECT 34.292 69.104 34.436 69.296 ; 
        RECT 37.352 69.104 37.424 69.296 ; 
        RECT 65.432 69.104 65.504 69.296 ; 
        RECT 0.632 73.424 0.704 73.616 ; 
        RECT 28.712 73.424 28.784 73.616 ; 
        RECT 33.68 73.424 33.788 73.616 ; 
        RECT 34.292 73.424 34.436 73.616 ; 
        RECT 37.352 73.424 37.424 73.616 ; 
        RECT 65.432 73.424 65.504 73.616 ; 
        RECT 0.632 77.744 0.704 77.936 ; 
        RECT 28.712 77.744 28.784 77.936 ; 
        RECT 33.68 77.744 33.788 77.936 ; 
        RECT 34.292 77.744 34.436 77.936 ; 
        RECT 37.352 77.744 37.424 77.936 ; 
        RECT 65.432 77.744 65.504 77.936 ; 
        RECT 0.632 82.064 0.704 82.256 ; 
        RECT 28.712 82.064 28.784 82.256 ; 
        RECT 33.68 82.064 33.788 82.256 ; 
        RECT 34.292 82.064 34.436 82.256 ; 
        RECT 37.352 82.064 37.424 82.256 ; 
        RECT 65.432 82.064 65.504 82.256 ; 
        RECT 0.632 86.384 0.704 86.576 ; 
        RECT 28.712 86.384 28.784 86.576 ; 
        RECT 33.68 86.384 33.788 86.576 ; 
        RECT 34.292 86.384 34.436 86.576 ; 
        RECT 37.352 86.384 37.424 86.576 ; 
        RECT 65.432 86.384 65.504 86.576 ; 
        RECT 0.632 90.704 0.704 90.896 ; 
        RECT 28.712 90.704 28.784 90.896 ; 
        RECT 33.68 90.704 33.788 90.896 ; 
        RECT 34.292 90.704 34.436 90.896 ; 
        RECT 37.352 90.704 37.424 90.896 ; 
        RECT 65.432 90.704 65.504 90.896 ; 
        RECT 0.632 95.024 0.704 95.216 ; 
        RECT 28.712 95.024 28.784 95.216 ; 
        RECT 33.68 95.024 33.788 95.216 ; 
        RECT 34.292 95.024 34.436 95.216 ; 
        RECT 37.352 95.024 37.424 95.216 ; 
        RECT 65.432 95.024 65.504 95.216 ; 
        RECT 0.632 99.344 0.704 99.536 ; 
        RECT 28.712 99.344 28.784 99.536 ; 
        RECT 33.68 99.344 33.788 99.536 ; 
        RECT 34.292 99.344 34.436 99.536 ; 
        RECT 37.352 99.344 37.424 99.536 ; 
        RECT 65.432 99.344 65.504 99.536 ; 
        RECT 0.632 103.664 0.704 103.856 ; 
        RECT 28.712 103.664 28.784 103.856 ; 
        RECT 33.68 103.664 33.788 103.856 ; 
        RECT 34.292 103.664 34.436 103.856 ; 
        RECT 37.352 103.664 37.424 103.856 ; 
        RECT 65.432 103.664 65.504 103.856 ; 
        RECT 33.532 133.044 33.604 133.908 ; 
        RECT 33.532 120.372 33.604 121.236 ; 
        RECT 33.532 107.7 33.604 108.564 ; 
        RECT 33.74 133.044 33.812 133.908 ; 
        RECT 33.74 120.372 33.812 121.236 ; 
        RECT 33.74 107.7 33.812 108.564 ; 
        RECT 33.948 133.044 34.02 133.908 ; 
        RECT 33.948 120.372 34.02 121.236 ; 
        RECT 33.948 107.7 34.02 108.564 ; 
        RECT 34.156 133.044 34.228 133.908 ; 
        RECT 34.156 120.372 34.228 121.236 ; 
        RECT 34.156 107.7 34.228 108.564 ; 
        RECT 34.364 133.044 34.436 133.908 ; 
        RECT 34.364 120.372 34.436 121.236 ; 
        RECT 34.364 107.7 34.436 108.564 ; 
        RECT 37.332 107.702 37.404 108.566 ; 
        RECT 0.632 140.492 0.704 140.684 ; 
        RECT 28.712 140.492 28.784 140.684 ; 
        RECT 33.68 140.492 33.788 140.684 ; 
        RECT 34.292 140.492 34.436 140.684 ; 
        RECT 37.352 140.492 37.424 140.684 ; 
        RECT 65.432 140.492 65.504 140.684 ; 
        RECT 0.632 144.812 0.704 145.004 ; 
        RECT 28.712 144.812 28.784 145.004 ; 
        RECT 33.68 144.812 33.788 145.004 ; 
        RECT 34.292 144.812 34.436 145.004 ; 
        RECT 37.352 144.812 37.424 145.004 ; 
        RECT 65.432 144.812 65.504 145.004 ; 
        RECT 0.632 149.132 0.704 149.324 ; 
        RECT 28.712 149.132 28.784 149.324 ; 
        RECT 33.68 149.132 33.788 149.324 ; 
        RECT 34.292 149.132 34.436 149.324 ; 
        RECT 37.352 149.132 37.424 149.324 ; 
        RECT 65.432 149.132 65.504 149.324 ; 
        RECT 0.632 153.452 0.704 153.644 ; 
        RECT 28.712 153.452 28.784 153.644 ; 
        RECT 33.68 153.452 33.788 153.644 ; 
        RECT 34.292 153.452 34.436 153.644 ; 
        RECT 37.352 153.452 37.424 153.644 ; 
        RECT 65.432 153.452 65.504 153.644 ; 
        RECT 0.632 157.772 0.704 157.964 ; 
        RECT 28.712 157.772 28.784 157.964 ; 
        RECT 33.68 157.772 33.788 157.964 ; 
        RECT 34.292 157.772 34.436 157.964 ; 
        RECT 37.352 157.772 37.424 157.964 ; 
        RECT 65.432 157.772 65.504 157.964 ; 
        RECT 0.632 162.092 0.704 162.284 ; 
        RECT 28.712 162.092 28.784 162.284 ; 
        RECT 33.68 162.092 33.788 162.284 ; 
        RECT 34.292 162.092 34.436 162.284 ; 
        RECT 37.352 162.092 37.424 162.284 ; 
        RECT 65.432 162.092 65.504 162.284 ; 
        RECT 0.632 166.412 0.704 166.604 ; 
        RECT 28.712 166.412 28.784 166.604 ; 
        RECT 33.68 166.412 33.788 166.604 ; 
        RECT 34.292 166.412 34.436 166.604 ; 
        RECT 37.352 166.412 37.424 166.604 ; 
        RECT 65.432 166.412 65.504 166.604 ; 
        RECT 0.632 170.732 0.704 170.924 ; 
        RECT 28.712 170.732 28.784 170.924 ; 
        RECT 33.68 170.732 33.788 170.924 ; 
        RECT 34.292 170.732 34.436 170.924 ; 
        RECT 37.352 170.732 37.424 170.924 ; 
        RECT 65.432 170.732 65.504 170.924 ; 
        RECT 0.632 175.052 0.704 175.244 ; 
        RECT 28.712 175.052 28.784 175.244 ; 
        RECT 33.68 175.052 33.788 175.244 ; 
        RECT 34.292 175.052 34.436 175.244 ; 
        RECT 37.352 175.052 37.424 175.244 ; 
        RECT 65.432 175.052 65.504 175.244 ; 
        RECT 0.632 179.372 0.704 179.564 ; 
        RECT 28.712 179.372 28.784 179.564 ; 
        RECT 33.68 179.372 33.788 179.564 ; 
        RECT 34.292 179.372 34.436 179.564 ; 
        RECT 37.352 179.372 37.424 179.564 ; 
        RECT 65.432 179.372 65.504 179.564 ; 
        RECT 0.632 183.692 0.704 183.884 ; 
        RECT 28.712 183.692 28.784 183.884 ; 
        RECT 33.68 183.692 33.788 183.884 ; 
        RECT 34.292 183.692 34.436 183.884 ; 
        RECT 37.352 183.692 37.424 183.884 ; 
        RECT 65.432 183.692 65.504 183.884 ; 
        RECT 0.632 188.012 0.704 188.204 ; 
        RECT 28.712 188.012 28.784 188.204 ; 
        RECT 33.68 188.012 33.788 188.204 ; 
        RECT 34.292 188.012 34.436 188.204 ; 
        RECT 37.352 188.012 37.424 188.204 ; 
        RECT 65.432 188.012 65.504 188.204 ; 
        RECT 0.632 192.332 0.704 192.524 ; 
        RECT 28.712 192.332 28.784 192.524 ; 
        RECT 33.68 192.332 33.788 192.524 ; 
        RECT 34.292 192.332 34.436 192.524 ; 
        RECT 37.352 192.332 37.424 192.524 ; 
        RECT 65.432 192.332 65.504 192.524 ; 
        RECT 0.632 196.652 0.704 196.844 ; 
        RECT 28.712 196.652 28.784 196.844 ; 
        RECT 33.68 196.652 33.788 196.844 ; 
        RECT 34.292 196.652 34.436 196.844 ; 
        RECT 37.352 196.652 37.424 196.844 ; 
        RECT 65.432 196.652 65.504 196.844 ; 
        RECT 0.632 200.972 0.704 201.164 ; 
        RECT 28.712 200.972 28.784 201.164 ; 
        RECT 33.68 200.972 33.788 201.164 ; 
        RECT 34.292 200.972 34.436 201.164 ; 
        RECT 37.352 200.972 37.424 201.164 ; 
        RECT 65.432 200.972 65.504 201.164 ; 
        RECT 0.632 205.292 0.704 205.484 ; 
        RECT 28.712 205.292 28.784 205.484 ; 
        RECT 33.68 205.292 33.788 205.484 ; 
        RECT 34.292 205.292 34.436 205.484 ; 
        RECT 37.352 205.292 37.424 205.484 ; 
        RECT 65.432 205.292 65.504 205.484 ; 
        RECT 0.632 209.612 0.704 209.804 ; 
        RECT 28.712 209.612 28.784 209.804 ; 
        RECT 33.68 209.612 33.788 209.804 ; 
        RECT 34.292 209.612 34.436 209.804 ; 
        RECT 37.352 209.612 37.424 209.804 ; 
        RECT 65.432 209.612 65.504 209.804 ; 
        RECT 0.632 213.932 0.704 214.124 ; 
        RECT 28.712 213.932 28.784 214.124 ; 
        RECT 33.68 213.932 33.788 214.124 ; 
        RECT 34.292 213.932 34.436 214.124 ; 
        RECT 37.352 213.932 37.424 214.124 ; 
        RECT 65.432 213.932 65.504 214.124 ; 
        RECT 0.632 218.252 0.704 218.444 ; 
        RECT 28.712 218.252 28.784 218.444 ; 
        RECT 33.68 218.252 33.788 218.444 ; 
        RECT 34.292 218.252 34.436 218.444 ; 
        RECT 37.352 218.252 37.424 218.444 ; 
        RECT 65.432 218.252 65.504 218.444 ; 
        RECT 0.632 222.572 0.704 222.764 ; 
        RECT 28.712 222.572 28.784 222.764 ; 
        RECT 33.68 222.572 33.788 222.764 ; 
        RECT 34.292 222.572 34.436 222.764 ; 
        RECT 37.352 222.572 37.424 222.764 ; 
        RECT 65.432 222.572 65.504 222.764 ; 
        RECT 0.632 226.892 0.704 227.084 ; 
        RECT 28.712 226.892 28.784 227.084 ; 
        RECT 33.68 226.892 33.788 227.084 ; 
        RECT 34.292 226.892 34.436 227.084 ; 
        RECT 37.352 226.892 37.424 227.084 ; 
        RECT 65.432 226.892 65.504 227.084 ; 
        RECT 0.632 231.212 0.704 231.404 ; 
        RECT 28.712 231.212 28.784 231.404 ; 
        RECT 33.68 231.212 33.788 231.404 ; 
        RECT 34.292 231.212 34.436 231.404 ; 
        RECT 37.352 231.212 37.424 231.404 ; 
        RECT 65.432 231.212 65.504 231.404 ; 
        RECT 0.632 235.532 0.704 235.724 ; 
        RECT 28.712 235.532 28.784 235.724 ; 
        RECT 33.68 235.532 33.788 235.724 ; 
        RECT 34.292 235.532 34.436 235.724 ; 
        RECT 37.352 235.532 37.424 235.724 ; 
        RECT 65.432 235.532 65.504 235.724 ; 
        RECT 0.632 239.852 0.704 240.044 ; 
        RECT 28.712 239.852 28.784 240.044 ; 
        RECT 33.68 239.852 33.788 240.044 ; 
        RECT 34.292 239.852 34.436 240.044 ; 
        RECT 37.352 239.852 37.424 240.044 ; 
        RECT 65.432 239.852 65.504 240.044 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 43.164 109.588 43.236 109.736 ; 
      LAYER M4 ; 
        RECT 42.956 109.62 43.292 109.716 ; 
      LAYER M5 ; 
        RECT 43.152 105.816 43.248 118.776 ; 
      LAYER V3 ; 
        RECT 43.164 109.62 43.236 109.716 ; 
      LAYER V4 ; 
        RECT 43.152 109.62 43.248 109.716 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 42.3 109.6 42.372 109.748 ; 
      LAYER M4 ; 
        RECT 42.092 109.62 42.428 109.716 ; 
      LAYER M5 ; 
        RECT 42.288 105.816 42.384 118.776 ; 
      LAYER V3 ; 
        RECT 42.3 109.62 42.372 109.716 ; 
      LAYER V4 ; 
        RECT 42.288 109.62 42.384 109.716 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 41.436 107.284 41.508 107.432 ; 
      LAYER M4 ; 
        RECT 41.228 107.316 41.564 107.412 ; 
      LAYER M5 ; 
        RECT 41.424 105.816 41.52 118.776 ; 
      LAYER V3 ; 
        RECT 41.436 107.316 41.508 107.412 ; 
      LAYER V4 ; 
        RECT 41.424 107.316 41.52 107.412 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 40.572 108.244 40.644 108.968 ; 
      LAYER M4 ; 
        RECT 40.364 108.852 40.7 108.948 ; 
      LAYER M5 ; 
        RECT 40.56 105.816 40.656 118.776 ; 
      LAYER V3 ; 
        RECT 40.572 108.852 40.644 108.948 ; 
      LAYER V4 ; 
        RECT 40.56 108.852 40.656 108.948 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 39.708 107.296 39.78 107.564 ; 
      LAYER M4 ; 
        RECT 39.5 107.316 39.836 107.412 ; 
      LAYER M5 ; 
        RECT 39.696 105.816 39.792 118.776 ; 
      LAYER V3 ; 
        RECT 39.708 107.316 39.78 107.412 ; 
      LAYER V4 ; 
        RECT 39.696 107.316 39.792 107.412 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 38.844 106.228 38.916 107.24 ; 
      LAYER M4 ; 
        RECT 38.636 107.124 38.972 107.22 ; 
      LAYER M5 ; 
        RECT 38.832 105.816 38.928 118.776 ; 
      LAYER V3 ; 
        RECT 38.844 107.124 38.916 107.22 ; 
      LAYER V4 ; 
        RECT 38.832 107.124 38.928 107.22 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.98 110.368 38.052 110.516 ; 
      LAYER M4 ; 
        RECT 37.772 110.388 38.108 110.484 ; 
      LAYER M5 ; 
        RECT 37.968 105.816 38.064 118.776 ; 
      LAYER V3 ; 
        RECT 37.98 110.388 38.052 110.484 ; 
      LAYER V4 ; 
        RECT 37.968 110.388 38.064 110.484 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 37.116 109.756 37.188 110.12 ; 
      LAYER M4 ; 
        RECT 36.908 110.004 37.244 110.1 ; 
      LAYER M5 ; 
        RECT 37.104 105.816 37.2 118.776 ; 
      LAYER V3 ; 
        RECT 37.116 110.004 37.188 110.1 ; 
      LAYER V4 ; 
        RECT 37.104 110.004 37.2 110.1 ; 
    END 
  END ADDRESS[7] 
  PIN ADDRESS[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 34.524 107.296 34.596 107.564 ; 
      LAYER M4 ; 
        RECT 33.388 107.316 34.64 107.412 ; 
      LAYER M5 ; 
        RECT 33.432 105.816 33.528 118.776 ; 
      LAYER V3 ; 
        RECT 34.524 107.316 34.596 107.412 ; 
      LAYER V4 ; 
        RECT 33.432 107.316 33.528 107.412 ; 
    END 
  END ADDRESS[8] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 32.94 106.228 33.012 107.24 ; 
      LAYER M4 ; 
        RECT 32.092 107.124 33.056 107.22 ; 
      LAYER M5 ; 
        RECT 32.136 105.816 32.232 118.776 ; 
      LAYER V3 ; 
        RECT 32.94 107.124 33.012 107.22 ; 
      LAYER V4 ; 
        RECT 32.136 107.124 32.232 107.22 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.772 107.296 29.844 107.564 ; 
      LAYER M4 ; 
        RECT 29.564 107.316 29.9 107.412 ; 
      LAYER M5 ; 
        RECT 29.76 105.816 29.856 118.776 ; 
      LAYER V3 ; 
        RECT 29.772 107.316 29.844 107.412 ; 
      LAYER V4 ; 
        RECT 29.76 107.316 29.856 107.412 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.908 110.752 28.98 110.948 ; 
      LAYER M4 ; 
        RECT 28.7 110.772 29.036 110.868 ; 
      LAYER M5 ; 
        RECT 28.896 105.816 28.992 118.776 ; 
      LAYER V3 ; 
        RECT 28.908 110.772 28.98 110.868 ; 
      LAYER V4 ; 
        RECT 28.896 110.772 28.992 110.868 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.052 106.228 29.124 107.24 ; 
      LAYER M4 ; 
        RECT 27.988 107.124 29.168 107.22 ; 
      LAYER M5 ; 
        RECT 28.032 105.816 28.128 118.776 ; 
      LAYER V3 ; 
        RECT 29.052 107.124 29.124 107.22 ; 
      LAYER V4 ; 
        RECT 28.032 107.124 28.128 107.22 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.18 109.588 27.252 109.736 ; 
      LAYER M4 ; 
        RECT 26.972 109.62 27.308 109.716 ; 
      LAYER M5 ; 
        RECT 27.168 105.816 27.264 118.776 ; 
      LAYER V3 ; 
        RECT 27.18 109.62 27.252 109.716 ; 
      LAYER V4 ; 
        RECT 27.168 109.62 27.264 109.716 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.316 107.296 26.388 108.212 ; 
      LAYER M4 ; 
        RECT 26.108 107.316 26.444 107.412 ; 
      LAYER M5 ; 
        RECT 26.304 105.816 26.4 118.776 ; 
      LAYER V3 ; 
        RECT 26.316 107.316 26.388 107.412 ; 
      LAYER V4 ; 
        RECT 26.304 107.316 26.4 107.412 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.452 106.228 25.524 107.24 ; 
      LAYER M4 ; 
        RECT 25.244 107.124 25.58 107.22 ; 
      LAYER M5 ; 
        RECT 25.44 105.816 25.536 118.776 ; 
      LAYER V3 ; 
        RECT 25.452 107.124 25.524 107.22 ; 
      LAYER V4 ; 
        RECT 25.44 107.124 25.536 107.22 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.588 107.284 24.66 107.432 ; 
      LAYER M4 ; 
        RECT 24.38 107.316 24.716 107.412 ; 
      LAYER M5 ; 
        RECT 24.576 105.816 24.672 118.776 ; 
      LAYER V3 ; 
        RECT 24.588 107.316 24.66 107.412 ; 
      LAYER V4 ; 
        RECT 24.576 107.316 24.672 107.412 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 23.724 109.588 23.796 109.736 ; 
      LAYER M4 ; 
        RECT 23.516 109.62 23.852 109.716 ; 
      LAYER M5 ; 
        RECT 23.712 105.816 23.808 118.776 ; 
      LAYER V3 ; 
        RECT 23.724 109.62 23.796 109.716 ; 
      LAYER V4 ; 
        RECT 23.712 109.62 23.808 109.716 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.712 34.388 1.808 ; 
      LAYER M3 ; 
        RECT 34.148 1.51 34.22 2.468 ; 
      LAYER V3 ; 
        RECT 34.148 1.712 34.22 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 1.328 34.66 1.424 ; 
      LAYER M3 ; 
        RECT 33.248 1.08 33.32 2.7 ; 
      LAYER V3 ; 
        RECT 33.248 1.328 33.32 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 6.032 34.388 6.128 ; 
      LAYER M3 ; 
        RECT 34.148 5.83 34.22 6.788 ; 
      LAYER V3 ; 
        RECT 34.148 6.032 34.22 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 5.648 34.66 5.744 ; 
      LAYER M3 ; 
        RECT 33.248 5.4 33.32 7.02 ; 
      LAYER V3 ; 
        RECT 33.248 5.648 33.32 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 10.352 34.388 10.448 ; 
      LAYER M3 ; 
        RECT 34.148 10.15 34.22 11.108 ; 
      LAYER V3 ; 
        RECT 34.148 10.352 34.22 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 9.968 34.66 10.064 ; 
      LAYER M3 ; 
        RECT 33.248 9.72 33.32 11.34 ; 
      LAYER V3 ; 
        RECT 33.248 9.968 33.32 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.672 34.388 14.768 ; 
      LAYER M3 ; 
        RECT 34.148 14.47 34.22 15.428 ; 
      LAYER V3 ; 
        RECT 34.148 14.672 34.22 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 14.288 34.66 14.384 ; 
      LAYER M3 ; 
        RECT 33.248 14.04 33.32 15.66 ; 
      LAYER V3 ; 
        RECT 33.248 14.288 33.32 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.992 34.388 19.088 ; 
      LAYER M3 ; 
        RECT 34.148 18.79 34.22 19.748 ; 
      LAYER V3 ; 
        RECT 34.148 18.992 34.22 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 18.608 34.66 18.704 ; 
      LAYER M3 ; 
        RECT 33.248 18.36 33.32 19.98 ; 
      LAYER V3 ; 
        RECT 33.248 18.608 33.32 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 23.312 34.388 23.408 ; 
      LAYER M3 ; 
        RECT 34.148 23.11 34.22 24.068 ; 
      LAYER V3 ; 
        RECT 34.148 23.312 34.22 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 22.928 34.66 23.024 ; 
      LAYER M3 ; 
        RECT 33.248 22.68 33.32 24.3 ; 
      LAYER V3 ; 
        RECT 33.248 22.928 33.32 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.632 34.388 27.728 ; 
      LAYER M3 ; 
        RECT 34.148 27.43 34.22 28.388 ; 
      LAYER V3 ; 
        RECT 34.148 27.632 34.22 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 27.248 34.66 27.344 ; 
      LAYER M3 ; 
        RECT 33.248 27 33.32 28.62 ; 
      LAYER V3 ; 
        RECT 33.248 27.248 33.32 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.952 34.388 32.048 ; 
      LAYER M3 ; 
        RECT 34.148 31.75 34.22 32.708 ; 
      LAYER V3 ; 
        RECT 34.148 31.952 34.22 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 31.568 34.66 31.664 ; 
      LAYER M3 ; 
        RECT 33.248 31.32 33.32 32.94 ; 
      LAYER V3 ; 
        RECT 33.248 31.568 33.32 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 36.272 34.388 36.368 ; 
      LAYER M3 ; 
        RECT 34.148 36.07 34.22 37.028 ; 
      LAYER V3 ; 
        RECT 34.148 36.272 34.22 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 35.888 34.66 35.984 ; 
      LAYER M3 ; 
        RECT 33.248 35.64 33.32 37.26 ; 
      LAYER V3 ; 
        RECT 33.248 35.888 33.32 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.592 34.388 40.688 ; 
      LAYER M3 ; 
        RECT 34.148 40.39 34.22 41.348 ; 
      LAYER V3 ; 
        RECT 34.148 40.592 34.22 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 40.208 34.66 40.304 ; 
      LAYER M3 ; 
        RECT 33.248 39.96 33.32 41.58 ; 
      LAYER V3 ; 
        RECT 33.248 40.208 33.32 40.304 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 44.912 34.388 45.008 ; 
      LAYER M3 ; 
        RECT 34.148 44.71 34.22 45.668 ; 
      LAYER V3 ; 
        RECT 34.148 44.912 34.22 45.008 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 44.528 34.66 44.624 ; 
      LAYER M3 ; 
        RECT 33.248 44.28 33.32 45.9 ; 
      LAYER V3 ; 
        RECT 33.248 44.528 33.32 44.624 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 49.232 34.388 49.328 ; 
      LAYER M3 ; 
        RECT 34.148 49.03 34.22 49.988 ; 
      LAYER V3 ; 
        RECT 34.148 49.232 34.22 49.328 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 48.848 34.66 48.944 ; 
      LAYER M3 ; 
        RECT 33.248 48.6 33.32 50.22 ; 
      LAYER V3 ; 
        RECT 33.248 48.848 33.32 48.944 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 53.552 34.388 53.648 ; 
      LAYER M3 ; 
        RECT 34.148 53.35 34.22 54.308 ; 
      LAYER V3 ; 
        RECT 34.148 53.552 34.22 53.648 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 53.168 34.66 53.264 ; 
      LAYER M3 ; 
        RECT 33.248 52.92 33.32 54.54 ; 
      LAYER V3 ; 
        RECT 33.248 53.168 33.32 53.264 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 57.872 34.388 57.968 ; 
      LAYER M3 ; 
        RECT 34.148 57.67 34.22 58.628 ; 
      LAYER V3 ; 
        RECT 34.148 57.872 34.22 57.968 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 57.488 34.66 57.584 ; 
      LAYER M3 ; 
        RECT 33.248 57.24 33.32 58.86 ; 
      LAYER V3 ; 
        RECT 33.248 57.488 33.32 57.584 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 62.192 34.388 62.288 ; 
      LAYER M3 ; 
        RECT 34.148 61.99 34.22 62.948 ; 
      LAYER V3 ; 
        RECT 34.148 62.192 34.22 62.288 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 61.808 34.66 61.904 ; 
      LAYER M3 ; 
        RECT 33.248 61.56 33.32 63.18 ; 
      LAYER V3 ; 
        RECT 33.248 61.808 33.32 61.904 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 66.512 34.388 66.608 ; 
      LAYER M3 ; 
        RECT 34.148 66.31 34.22 67.268 ; 
      LAYER V3 ; 
        RECT 34.148 66.512 34.22 66.608 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 66.128 34.66 66.224 ; 
      LAYER M3 ; 
        RECT 33.248 65.88 33.32 67.5 ; 
      LAYER V3 ; 
        RECT 33.248 66.128 33.32 66.224 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 70.832 34.388 70.928 ; 
      LAYER M3 ; 
        RECT 34.148 70.63 34.22 71.588 ; 
      LAYER V3 ; 
        RECT 34.148 70.832 34.22 70.928 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 70.448 34.66 70.544 ; 
      LAYER M3 ; 
        RECT 33.248 70.2 33.32 71.82 ; 
      LAYER V3 ; 
        RECT 33.248 70.448 33.32 70.544 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 75.152 34.388 75.248 ; 
      LAYER M3 ; 
        RECT 34.148 74.95 34.22 75.908 ; 
      LAYER V3 ; 
        RECT 34.148 75.152 34.22 75.248 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 74.768 34.66 74.864 ; 
      LAYER M3 ; 
        RECT 33.248 74.52 33.32 76.14 ; 
      LAYER V3 ; 
        RECT 33.248 74.768 33.32 74.864 ; 
    END 
  END wd[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 79.472 34.388 79.568 ; 
      LAYER M3 ; 
        RECT 34.148 79.27 34.22 80.228 ; 
      LAYER V3 ; 
        RECT 34.148 79.472 34.22 79.568 ; 
    END 
  END dataout[18] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 79.088 34.66 79.184 ; 
      LAYER M3 ; 
        RECT 33.248 78.84 33.32 80.46 ; 
      LAYER V3 ; 
        RECT 33.248 79.088 33.32 79.184 ; 
    END 
  END wd[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 83.792 34.388 83.888 ; 
      LAYER M3 ; 
        RECT 34.148 83.59 34.22 84.548 ; 
      LAYER V3 ; 
        RECT 34.148 83.792 34.22 83.888 ; 
    END 
  END dataout[19] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 83.408 34.66 83.504 ; 
      LAYER M3 ; 
        RECT 33.248 83.16 33.32 84.78 ; 
      LAYER V3 ; 
        RECT 33.248 83.408 33.32 83.504 ; 
    END 
  END wd[19] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 88.112 34.388 88.208 ; 
      LAYER M3 ; 
        RECT 34.148 87.91 34.22 88.868 ; 
      LAYER V3 ; 
        RECT 34.148 88.112 34.22 88.208 ; 
    END 
  END dataout[20] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 87.728 34.66 87.824 ; 
      LAYER M3 ; 
        RECT 33.248 87.48 33.32 89.1 ; 
      LAYER V3 ; 
        RECT 33.248 87.728 33.32 87.824 ; 
    END 
  END wd[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 92.432 34.388 92.528 ; 
      LAYER M3 ; 
        RECT 34.148 92.23 34.22 93.188 ; 
      LAYER V3 ; 
        RECT 34.148 92.432 34.22 92.528 ; 
    END 
  END dataout[21] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 92.048 34.66 92.144 ; 
      LAYER M3 ; 
        RECT 33.248 91.8 33.32 93.42 ; 
      LAYER V3 ; 
        RECT 33.248 92.048 33.32 92.144 ; 
    END 
  END wd[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 96.752 34.388 96.848 ; 
      LAYER M3 ; 
        RECT 34.148 96.55 34.22 97.508 ; 
      LAYER V3 ; 
        RECT 34.148 96.752 34.22 96.848 ; 
    END 
  END dataout[22] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 96.368 34.66 96.464 ; 
      LAYER M3 ; 
        RECT 33.248 96.12 33.32 97.74 ; 
      LAYER V3 ; 
        RECT 33.248 96.368 33.32 96.464 ; 
    END 
  END wd[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 101.072 34.388 101.168 ; 
      LAYER M3 ; 
        RECT 34.148 100.87 34.22 101.828 ; 
      LAYER V3 ; 
        RECT 34.148 101.072 34.22 101.168 ; 
    END 
  END dataout[23] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 100.688 34.66 100.784 ; 
      LAYER M3 ; 
        RECT 33.248 100.44 33.32 102.06 ; 
      LAYER V3 ; 
        RECT 33.248 100.688 33.32 100.784 ; 
    END 
  END wd[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 137.9 34.388 137.996 ; 
      LAYER M3 ; 
        RECT 34.148 137.698 34.22 138.656 ; 
      LAYER V3 ; 
        RECT 34.148 137.9 34.22 137.996 ; 
    END 
  END dataout[24] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 137.516 34.66 137.612 ; 
      LAYER M3 ; 
        RECT 33.248 137.268 33.32 138.888 ; 
      LAYER V3 ; 
        RECT 33.248 137.516 33.32 137.612 ; 
    END 
  END wd[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 142.22 34.388 142.316 ; 
      LAYER M3 ; 
        RECT 34.148 142.018 34.22 142.976 ; 
      LAYER V3 ; 
        RECT 34.148 142.22 34.22 142.316 ; 
    END 
  END dataout[25] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 141.836 34.66 141.932 ; 
      LAYER M3 ; 
        RECT 33.248 141.588 33.32 143.208 ; 
      LAYER V3 ; 
        RECT 33.248 141.836 33.32 141.932 ; 
    END 
  END wd[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 146.54 34.388 146.636 ; 
      LAYER M3 ; 
        RECT 34.148 146.338 34.22 147.296 ; 
      LAYER V3 ; 
        RECT 34.148 146.54 34.22 146.636 ; 
    END 
  END dataout[26] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 146.156 34.66 146.252 ; 
      LAYER M3 ; 
        RECT 33.248 145.908 33.32 147.528 ; 
      LAYER V3 ; 
        RECT 33.248 146.156 33.32 146.252 ; 
    END 
  END wd[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 150.86 34.388 150.956 ; 
      LAYER M3 ; 
        RECT 34.148 150.658 34.22 151.616 ; 
      LAYER V3 ; 
        RECT 34.148 150.86 34.22 150.956 ; 
    END 
  END dataout[27] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 150.476 34.66 150.572 ; 
      LAYER M3 ; 
        RECT 33.248 150.228 33.32 151.848 ; 
      LAYER V3 ; 
        RECT 33.248 150.476 33.32 150.572 ; 
    END 
  END wd[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 155.18 34.388 155.276 ; 
      LAYER M3 ; 
        RECT 34.148 154.978 34.22 155.936 ; 
      LAYER V3 ; 
        RECT 34.148 155.18 34.22 155.276 ; 
    END 
  END dataout[28] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 154.796 34.66 154.892 ; 
      LAYER M3 ; 
        RECT 33.248 154.548 33.32 156.168 ; 
      LAYER V3 ; 
        RECT 33.248 154.796 33.32 154.892 ; 
    END 
  END wd[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 159.5 34.388 159.596 ; 
      LAYER M3 ; 
        RECT 34.148 159.298 34.22 160.256 ; 
      LAYER V3 ; 
        RECT 34.148 159.5 34.22 159.596 ; 
    END 
  END dataout[29] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 159.116 34.66 159.212 ; 
      LAYER M3 ; 
        RECT 33.248 158.868 33.32 160.488 ; 
      LAYER V3 ; 
        RECT 33.248 159.116 33.32 159.212 ; 
    END 
  END wd[29] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 163.82 34.388 163.916 ; 
      LAYER M3 ; 
        RECT 34.148 163.618 34.22 164.576 ; 
      LAYER V3 ; 
        RECT 34.148 163.82 34.22 163.916 ; 
    END 
  END dataout[30] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 163.436 34.66 163.532 ; 
      LAYER M3 ; 
        RECT 33.248 163.188 33.32 164.808 ; 
      LAYER V3 ; 
        RECT 33.248 163.436 33.32 163.532 ; 
    END 
  END wd[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 168.14 34.388 168.236 ; 
      LAYER M3 ; 
        RECT 34.148 167.938 34.22 168.896 ; 
      LAYER V3 ; 
        RECT 34.148 168.14 34.22 168.236 ; 
    END 
  END dataout[31] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 167.756 34.66 167.852 ; 
      LAYER M3 ; 
        RECT 33.248 167.508 33.32 169.128 ; 
      LAYER V3 ; 
        RECT 33.248 167.756 33.32 167.852 ; 
    END 
  END wd[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 172.46 34.388 172.556 ; 
      LAYER M3 ; 
        RECT 34.148 172.258 34.22 173.216 ; 
      LAYER V3 ; 
        RECT 34.148 172.46 34.22 172.556 ; 
    END 
  END dataout[32] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 172.076 34.66 172.172 ; 
      LAYER M3 ; 
        RECT 33.248 171.828 33.32 173.448 ; 
      LAYER V3 ; 
        RECT 33.248 172.076 33.32 172.172 ; 
    END 
  END wd[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 176.78 34.388 176.876 ; 
      LAYER M3 ; 
        RECT 34.148 176.578 34.22 177.536 ; 
      LAYER V3 ; 
        RECT 34.148 176.78 34.22 176.876 ; 
    END 
  END dataout[33] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 176.396 34.66 176.492 ; 
      LAYER M3 ; 
        RECT 33.248 176.148 33.32 177.768 ; 
      LAYER V3 ; 
        RECT 33.248 176.396 33.32 176.492 ; 
    END 
  END wd[33] 
  PIN dataout[34] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 181.1 34.388 181.196 ; 
      LAYER M3 ; 
        RECT 34.148 180.898 34.22 181.856 ; 
      LAYER V3 ; 
        RECT 34.148 181.1 34.22 181.196 ; 
    END 
  END dataout[34] 
  PIN wd[34] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 180.716 34.66 180.812 ; 
      LAYER M3 ; 
        RECT 33.248 180.468 33.32 182.088 ; 
      LAYER V3 ; 
        RECT 33.248 180.716 33.32 180.812 ; 
    END 
  END wd[34] 
  PIN dataout[35] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 185.42 34.388 185.516 ; 
      LAYER M3 ; 
        RECT 34.148 185.218 34.22 186.176 ; 
      LAYER V3 ; 
        RECT 34.148 185.42 34.22 185.516 ; 
    END 
  END dataout[35] 
  PIN wd[35] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 185.036 34.66 185.132 ; 
      LAYER M3 ; 
        RECT 33.248 184.788 33.32 186.408 ; 
      LAYER V3 ; 
        RECT 33.248 185.036 33.32 185.132 ; 
    END 
  END wd[35] 
  PIN dataout[36] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 189.74 34.388 189.836 ; 
      LAYER M3 ; 
        RECT 34.148 189.538 34.22 190.496 ; 
      LAYER V3 ; 
        RECT 34.148 189.74 34.22 189.836 ; 
    END 
  END dataout[36] 
  PIN wd[36] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 189.356 34.66 189.452 ; 
      LAYER M3 ; 
        RECT 33.248 189.108 33.32 190.728 ; 
      LAYER V3 ; 
        RECT 33.248 189.356 33.32 189.452 ; 
    END 
  END wd[36] 
  PIN dataout[37] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 194.06 34.388 194.156 ; 
      LAYER M3 ; 
        RECT 34.148 193.858 34.22 194.816 ; 
      LAYER V3 ; 
        RECT 34.148 194.06 34.22 194.156 ; 
    END 
  END dataout[37] 
  PIN wd[37] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 193.676 34.66 193.772 ; 
      LAYER M3 ; 
        RECT 33.248 193.428 33.32 195.048 ; 
      LAYER V3 ; 
        RECT 33.248 193.676 33.32 193.772 ; 
    END 
  END wd[37] 
  PIN dataout[38] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 198.38 34.388 198.476 ; 
      LAYER M3 ; 
        RECT 34.148 198.178 34.22 199.136 ; 
      LAYER V3 ; 
        RECT 34.148 198.38 34.22 198.476 ; 
    END 
  END dataout[38] 
  PIN wd[38] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 197.996 34.66 198.092 ; 
      LAYER M3 ; 
        RECT 33.248 197.748 33.32 199.368 ; 
      LAYER V3 ; 
        RECT 33.248 197.996 33.32 198.092 ; 
    END 
  END wd[38] 
  PIN dataout[39] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 202.7 34.388 202.796 ; 
      LAYER M3 ; 
        RECT 34.148 202.498 34.22 203.456 ; 
      LAYER V3 ; 
        RECT 34.148 202.7 34.22 202.796 ; 
    END 
  END dataout[39] 
  PIN wd[39] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 202.316 34.66 202.412 ; 
      LAYER M3 ; 
        RECT 33.248 202.068 33.32 203.688 ; 
      LAYER V3 ; 
        RECT 33.248 202.316 33.32 202.412 ; 
    END 
  END wd[39] 
  PIN dataout[40] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 207.02 34.388 207.116 ; 
      LAYER M3 ; 
        RECT 34.148 206.818 34.22 207.776 ; 
      LAYER V3 ; 
        RECT 34.148 207.02 34.22 207.116 ; 
    END 
  END dataout[40] 
  PIN wd[40] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 206.636 34.66 206.732 ; 
      LAYER M3 ; 
        RECT 33.248 206.388 33.32 208.008 ; 
      LAYER V3 ; 
        RECT 33.248 206.636 33.32 206.732 ; 
    END 
  END wd[40] 
  PIN dataout[41] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 211.34 34.388 211.436 ; 
      LAYER M3 ; 
        RECT 34.148 211.138 34.22 212.096 ; 
      LAYER V3 ; 
        RECT 34.148 211.34 34.22 211.436 ; 
    END 
  END dataout[41] 
  PIN wd[41] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 210.956 34.66 211.052 ; 
      LAYER M3 ; 
        RECT 33.248 210.708 33.32 212.328 ; 
      LAYER V3 ; 
        RECT 33.248 210.956 33.32 211.052 ; 
    END 
  END wd[41] 
  PIN dataout[42] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 215.66 34.388 215.756 ; 
      LAYER M3 ; 
        RECT 34.148 215.458 34.22 216.416 ; 
      LAYER V3 ; 
        RECT 34.148 215.66 34.22 215.756 ; 
    END 
  END dataout[42] 
  PIN wd[42] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 215.276 34.66 215.372 ; 
      LAYER M3 ; 
        RECT 33.248 215.028 33.32 216.648 ; 
      LAYER V3 ; 
        RECT 33.248 215.276 33.32 215.372 ; 
    END 
  END wd[42] 
  PIN dataout[43] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 219.98 34.388 220.076 ; 
      LAYER M3 ; 
        RECT 34.148 219.778 34.22 220.736 ; 
      LAYER V3 ; 
        RECT 34.148 219.98 34.22 220.076 ; 
    END 
  END dataout[43] 
  PIN wd[43] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 219.596 34.66 219.692 ; 
      LAYER M3 ; 
        RECT 33.248 219.348 33.32 220.968 ; 
      LAYER V3 ; 
        RECT 33.248 219.596 33.32 219.692 ; 
    END 
  END wd[43] 
  PIN dataout[44] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 224.3 34.388 224.396 ; 
      LAYER M3 ; 
        RECT 34.148 224.098 34.22 225.056 ; 
      LAYER V3 ; 
        RECT 34.148 224.3 34.22 224.396 ; 
    END 
  END dataout[44] 
  PIN wd[44] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 223.916 34.66 224.012 ; 
      LAYER M3 ; 
        RECT 33.248 223.668 33.32 225.288 ; 
      LAYER V3 ; 
        RECT 33.248 223.916 33.32 224.012 ; 
    END 
  END wd[44] 
  PIN dataout[45] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 228.62 34.388 228.716 ; 
      LAYER M3 ; 
        RECT 34.148 228.418 34.22 229.376 ; 
      LAYER V3 ; 
        RECT 34.148 228.62 34.22 228.716 ; 
    END 
  END dataout[45] 
  PIN wd[45] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 228.236 34.66 228.332 ; 
      LAYER M3 ; 
        RECT 33.248 227.988 33.32 229.608 ; 
      LAYER V3 ; 
        RECT 33.248 228.236 33.32 228.332 ; 
    END 
  END wd[45] 
  PIN dataout[46] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 232.94 34.388 233.036 ; 
      LAYER M3 ; 
        RECT 34.148 232.738 34.22 233.696 ; 
      LAYER V3 ; 
        RECT 34.148 232.94 34.22 233.036 ; 
    END 
  END dataout[46] 
  PIN wd[46] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 232.556 34.66 232.652 ; 
      LAYER M3 ; 
        RECT 33.248 232.308 33.32 233.928 ; 
      LAYER V3 ; 
        RECT 33.248 232.556 33.32 232.652 ; 
    END 
  END wd[46] 
  PIN dataout[47] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 237.26 34.388 237.356 ; 
      LAYER M3 ; 
        RECT 34.148 237.058 34.22 238.016 ; 
      LAYER V3 ; 
        RECT 34.148 237.26 34.22 237.356 ; 
    END 
  END dataout[47] 
  PIN wd[47] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 31.796 236.876 34.66 236.972 ; 
      LAYER M3 ; 
        RECT 33.248 236.628 33.32 238.248 ; 
      LAYER V3 ; 
        RECT 33.248 236.876 33.32 236.972 ; 
    END 
  END wd[47] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0 104.628 66.096 139.242 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
        RECT 0.02 180.414 66.116 184.788 ; 
        RECT 0.02 184.734 66.116 189.108 ; 
        RECT 0.02 189.054 66.116 193.428 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0 104.628 66.096 139.242 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
        RECT 0.02 180.414 66.116 184.788 ; 
        RECT 0.02 184.734 66.116 189.108 ; 
        RECT 0.02 189.054 66.116 193.428 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
  LAYER V1 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0 104.628 66.096 139.242 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
        RECT 0.02 180.414 66.116 184.788 ; 
        RECT 0.02 184.734 66.116 189.108 ; 
        RECT 0.02 189.054 66.116 193.428 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
  LAYER V2 SPACING 0.072 ; 
      RECT 0.02 1.026 66.116 5.4 ; 
      RECT 0.02 5.346 66.116 9.72 ; 
      RECT 0.02 9.666 66.116 14.04 ; 
      RECT 0.02 13.986 66.116 18.36 ; 
      RECT 0.02 18.306 66.116 22.68 ; 
      RECT 0.02 22.626 66.116 27 ; 
      RECT 0.02 26.946 66.116 31.32 ; 
      RECT 0.02 31.266 66.116 35.64 ; 
      RECT 0.02 35.586 66.116 39.96 ; 
      RECT 0.02 39.906 66.116 44.28 ; 
      RECT 0.02 44.226 66.116 48.6 ; 
      RECT 0.02 48.546 66.116 52.92 ; 
      RECT 0.02 52.866 66.116 57.24 ; 
      RECT 0.02 57.186 66.116 61.56 ; 
      RECT 0.02 61.506 66.116 65.88 ; 
      RECT 0.02 65.826 66.116 70.2 ; 
      RECT 0.02 70.146 66.116 74.52 ; 
      RECT 0.02 74.466 66.116 78.84 ; 
      RECT 0.02 78.786 66.116 83.16 ; 
      RECT 0.02 83.106 66.116 87.48 ; 
      RECT 0.02 87.426 66.116 91.8 ; 
      RECT 0.02 91.746 66.116 96.12 ; 
      RECT 0.02 96.066 66.116 100.44 ; 
      RECT 0.02 100.386 66.116 104.76 ; 
      RECT 0 104.628 66.096 139.242 ; 
        RECT 0.02 137.214 66.116 141.588 ; 
        RECT 0.02 141.534 66.116 145.908 ; 
        RECT 0.02 145.854 66.116 150.228 ; 
        RECT 0.02 150.174 66.116 154.548 ; 
        RECT 0.02 154.494 66.116 158.868 ; 
        RECT 0.02 158.814 66.116 163.188 ; 
        RECT 0.02 163.134 66.116 167.508 ; 
        RECT 0.02 167.454 66.116 171.828 ; 
        RECT 0.02 171.774 66.116 176.148 ; 
        RECT 0.02 176.094 66.116 180.468 ; 
        RECT 0.02 180.414 66.116 184.788 ; 
        RECT 0.02 184.734 66.116 189.108 ; 
        RECT 0.02 189.054 66.116 193.428 ; 
        RECT 0.02 193.374 66.116 197.748 ; 
        RECT 0.02 197.694 66.116 202.068 ; 
        RECT 0.02 202.014 66.116 206.388 ; 
        RECT 0.02 206.334 66.116 210.708 ; 
        RECT 0.02 210.654 66.116 215.028 ; 
        RECT 0.02 214.974 66.116 219.348 ; 
        RECT 0.02 219.294 66.116 223.668 ; 
        RECT 0.02 223.614 66.116 227.988 ; 
        RECT 0.02 227.934 66.116 232.308 ; 
        RECT 0.02 232.254 66.116 236.628 ; 
        RECT 0.02 236.574 66.116 240.948 ; 
  LAYER M3 ; 
      RECT 34.796 1.38 34.868 5.122 ; 
      RECT 34.652 1.38 34.724 5.122 ; 
      RECT 34.508 3.688 34.58 4.978 ; 
      RECT 34.04 4.476 34.112 4.914 ; 
      RECT 34.004 1.51 34.076 2.468 ; 
      RECT 33.86 3.834 33.932 4.448 ; 
      RECT 33.536 3.936 33.608 4.968 ; 
      RECT 31.376 1.38 31.448 5.122 ; 
      RECT 31.232 1.38 31.304 5.122 ; 
      RECT 31.088 2.104 31.16 4.376 ; 
      RECT 34.796 5.7 34.868 9.442 ; 
      RECT 34.652 5.7 34.724 9.442 ; 
      RECT 34.508 8.008 34.58 9.298 ; 
      RECT 34.04 8.796 34.112 9.234 ; 
      RECT 34.004 5.83 34.076 6.788 ; 
      RECT 33.86 8.154 33.932 8.768 ; 
      RECT 33.536 8.256 33.608 9.288 ; 
      RECT 31.376 5.7 31.448 9.442 ; 
      RECT 31.232 5.7 31.304 9.442 ; 
      RECT 31.088 6.424 31.16 8.696 ; 
      RECT 34.796 10.02 34.868 13.762 ; 
      RECT 34.652 10.02 34.724 13.762 ; 
      RECT 34.508 12.328 34.58 13.618 ; 
      RECT 34.04 13.116 34.112 13.554 ; 
      RECT 34.004 10.15 34.076 11.108 ; 
      RECT 33.86 12.474 33.932 13.088 ; 
      RECT 33.536 12.576 33.608 13.608 ; 
      RECT 31.376 10.02 31.448 13.762 ; 
      RECT 31.232 10.02 31.304 13.762 ; 
      RECT 31.088 10.744 31.16 13.016 ; 
      RECT 34.796 14.34 34.868 18.082 ; 
      RECT 34.652 14.34 34.724 18.082 ; 
      RECT 34.508 16.648 34.58 17.938 ; 
      RECT 34.04 17.436 34.112 17.874 ; 
      RECT 34.004 14.47 34.076 15.428 ; 
      RECT 33.86 16.794 33.932 17.408 ; 
      RECT 33.536 16.896 33.608 17.928 ; 
      RECT 31.376 14.34 31.448 18.082 ; 
      RECT 31.232 14.34 31.304 18.082 ; 
      RECT 31.088 15.064 31.16 17.336 ; 
      RECT 34.796 18.66 34.868 22.402 ; 
      RECT 34.652 18.66 34.724 22.402 ; 
      RECT 34.508 20.968 34.58 22.258 ; 
      RECT 34.04 21.756 34.112 22.194 ; 
      RECT 34.004 18.79 34.076 19.748 ; 
      RECT 33.86 21.114 33.932 21.728 ; 
      RECT 33.536 21.216 33.608 22.248 ; 
      RECT 31.376 18.66 31.448 22.402 ; 
      RECT 31.232 18.66 31.304 22.402 ; 
      RECT 31.088 19.384 31.16 21.656 ; 
      RECT 34.796 22.98 34.868 26.722 ; 
      RECT 34.652 22.98 34.724 26.722 ; 
      RECT 34.508 25.288 34.58 26.578 ; 
      RECT 34.04 26.076 34.112 26.514 ; 
      RECT 34.004 23.11 34.076 24.068 ; 
      RECT 33.86 25.434 33.932 26.048 ; 
      RECT 33.536 25.536 33.608 26.568 ; 
      RECT 31.376 22.98 31.448 26.722 ; 
      RECT 31.232 22.98 31.304 26.722 ; 
      RECT 31.088 23.704 31.16 25.976 ; 
      RECT 34.796 27.3 34.868 31.042 ; 
      RECT 34.652 27.3 34.724 31.042 ; 
      RECT 34.508 29.608 34.58 30.898 ; 
      RECT 34.04 30.396 34.112 30.834 ; 
      RECT 34.004 27.43 34.076 28.388 ; 
      RECT 33.86 29.754 33.932 30.368 ; 
      RECT 33.536 29.856 33.608 30.888 ; 
      RECT 31.376 27.3 31.448 31.042 ; 
      RECT 31.232 27.3 31.304 31.042 ; 
      RECT 31.088 28.024 31.16 30.296 ; 
      RECT 34.796 31.62 34.868 35.362 ; 
      RECT 34.652 31.62 34.724 35.362 ; 
      RECT 34.508 33.928 34.58 35.218 ; 
      RECT 34.04 34.716 34.112 35.154 ; 
      RECT 34.004 31.75 34.076 32.708 ; 
      RECT 33.86 34.074 33.932 34.688 ; 
      RECT 33.536 34.176 33.608 35.208 ; 
      RECT 31.376 31.62 31.448 35.362 ; 
      RECT 31.232 31.62 31.304 35.362 ; 
      RECT 31.088 32.344 31.16 34.616 ; 
      RECT 34.796 35.94 34.868 39.682 ; 
      RECT 34.652 35.94 34.724 39.682 ; 
      RECT 34.508 38.248 34.58 39.538 ; 
      RECT 34.04 39.036 34.112 39.474 ; 
      RECT 34.004 36.07 34.076 37.028 ; 
      RECT 33.86 38.394 33.932 39.008 ; 
      RECT 33.536 38.496 33.608 39.528 ; 
      RECT 31.376 35.94 31.448 39.682 ; 
      RECT 31.232 35.94 31.304 39.682 ; 
      RECT 31.088 36.664 31.16 38.936 ; 
      RECT 34.796 40.26 34.868 44.002 ; 
      RECT 34.652 40.26 34.724 44.002 ; 
      RECT 34.508 42.568 34.58 43.858 ; 
      RECT 34.04 43.356 34.112 43.794 ; 
      RECT 34.004 40.39 34.076 41.348 ; 
      RECT 33.86 42.714 33.932 43.328 ; 
      RECT 33.536 42.816 33.608 43.848 ; 
      RECT 31.376 40.26 31.448 44.002 ; 
      RECT 31.232 40.26 31.304 44.002 ; 
      RECT 31.088 40.984 31.16 43.256 ; 
      RECT 34.796 44.58 34.868 48.322 ; 
      RECT 34.652 44.58 34.724 48.322 ; 
      RECT 34.508 46.888 34.58 48.178 ; 
      RECT 34.04 47.676 34.112 48.114 ; 
      RECT 34.004 44.71 34.076 45.668 ; 
      RECT 33.86 47.034 33.932 47.648 ; 
      RECT 33.536 47.136 33.608 48.168 ; 
      RECT 31.376 44.58 31.448 48.322 ; 
      RECT 31.232 44.58 31.304 48.322 ; 
      RECT 31.088 45.304 31.16 47.576 ; 
      RECT 34.796 48.9 34.868 52.642 ; 
      RECT 34.652 48.9 34.724 52.642 ; 
      RECT 34.508 51.208 34.58 52.498 ; 
      RECT 34.04 51.996 34.112 52.434 ; 
      RECT 34.004 49.03 34.076 49.988 ; 
      RECT 33.86 51.354 33.932 51.968 ; 
      RECT 33.536 51.456 33.608 52.488 ; 
      RECT 31.376 48.9 31.448 52.642 ; 
      RECT 31.232 48.9 31.304 52.642 ; 
      RECT 31.088 49.624 31.16 51.896 ; 
      RECT 34.796 53.22 34.868 56.962 ; 
      RECT 34.652 53.22 34.724 56.962 ; 
      RECT 34.508 55.528 34.58 56.818 ; 
      RECT 34.04 56.316 34.112 56.754 ; 
      RECT 34.004 53.35 34.076 54.308 ; 
      RECT 33.86 55.674 33.932 56.288 ; 
      RECT 33.536 55.776 33.608 56.808 ; 
      RECT 31.376 53.22 31.448 56.962 ; 
      RECT 31.232 53.22 31.304 56.962 ; 
      RECT 31.088 53.944 31.16 56.216 ; 
      RECT 34.796 57.54 34.868 61.282 ; 
      RECT 34.652 57.54 34.724 61.282 ; 
      RECT 34.508 59.848 34.58 61.138 ; 
      RECT 34.04 60.636 34.112 61.074 ; 
      RECT 34.004 57.67 34.076 58.628 ; 
      RECT 33.86 59.994 33.932 60.608 ; 
      RECT 33.536 60.096 33.608 61.128 ; 
      RECT 31.376 57.54 31.448 61.282 ; 
      RECT 31.232 57.54 31.304 61.282 ; 
      RECT 31.088 58.264 31.16 60.536 ; 
      RECT 34.796 61.86 34.868 65.602 ; 
      RECT 34.652 61.86 34.724 65.602 ; 
      RECT 34.508 64.168 34.58 65.458 ; 
      RECT 34.04 64.956 34.112 65.394 ; 
      RECT 34.004 61.99 34.076 62.948 ; 
      RECT 33.86 64.314 33.932 64.928 ; 
      RECT 33.536 64.416 33.608 65.448 ; 
      RECT 31.376 61.86 31.448 65.602 ; 
      RECT 31.232 61.86 31.304 65.602 ; 
      RECT 31.088 62.584 31.16 64.856 ; 
      RECT 34.796 66.18 34.868 69.922 ; 
      RECT 34.652 66.18 34.724 69.922 ; 
      RECT 34.508 68.488 34.58 69.778 ; 
      RECT 34.04 69.276 34.112 69.714 ; 
      RECT 34.004 66.31 34.076 67.268 ; 
      RECT 33.86 68.634 33.932 69.248 ; 
      RECT 33.536 68.736 33.608 69.768 ; 
      RECT 31.376 66.18 31.448 69.922 ; 
      RECT 31.232 66.18 31.304 69.922 ; 
      RECT 31.088 66.904 31.16 69.176 ; 
      RECT 34.796 70.5 34.868 74.242 ; 
      RECT 34.652 70.5 34.724 74.242 ; 
      RECT 34.508 72.808 34.58 74.098 ; 
      RECT 34.04 73.596 34.112 74.034 ; 
      RECT 34.004 70.63 34.076 71.588 ; 
      RECT 33.86 72.954 33.932 73.568 ; 
      RECT 33.536 73.056 33.608 74.088 ; 
      RECT 31.376 70.5 31.448 74.242 ; 
      RECT 31.232 70.5 31.304 74.242 ; 
      RECT 31.088 71.224 31.16 73.496 ; 
      RECT 34.796 74.82 34.868 78.562 ; 
      RECT 34.652 74.82 34.724 78.562 ; 
      RECT 34.508 77.128 34.58 78.418 ; 
      RECT 34.04 77.916 34.112 78.354 ; 
      RECT 34.004 74.95 34.076 75.908 ; 
      RECT 33.86 77.274 33.932 77.888 ; 
      RECT 33.536 77.376 33.608 78.408 ; 
      RECT 31.376 74.82 31.448 78.562 ; 
      RECT 31.232 74.82 31.304 78.562 ; 
      RECT 31.088 75.544 31.16 77.816 ; 
      RECT 34.796 79.14 34.868 82.882 ; 
      RECT 34.652 79.14 34.724 82.882 ; 
      RECT 34.508 81.448 34.58 82.738 ; 
      RECT 34.04 82.236 34.112 82.674 ; 
      RECT 34.004 79.27 34.076 80.228 ; 
      RECT 33.86 81.594 33.932 82.208 ; 
      RECT 33.536 81.696 33.608 82.728 ; 
      RECT 31.376 79.14 31.448 82.882 ; 
      RECT 31.232 79.14 31.304 82.882 ; 
      RECT 31.088 79.864 31.16 82.136 ; 
      RECT 34.796 83.46 34.868 87.202 ; 
      RECT 34.652 83.46 34.724 87.202 ; 
      RECT 34.508 85.768 34.58 87.058 ; 
      RECT 34.04 86.556 34.112 86.994 ; 
      RECT 34.004 83.59 34.076 84.548 ; 
      RECT 33.86 85.914 33.932 86.528 ; 
      RECT 33.536 86.016 33.608 87.048 ; 
      RECT 31.376 83.46 31.448 87.202 ; 
      RECT 31.232 83.46 31.304 87.202 ; 
      RECT 31.088 84.184 31.16 86.456 ; 
      RECT 34.796 87.78 34.868 91.522 ; 
      RECT 34.652 87.78 34.724 91.522 ; 
      RECT 34.508 90.088 34.58 91.378 ; 
      RECT 34.04 90.876 34.112 91.314 ; 
      RECT 34.004 87.91 34.076 88.868 ; 
      RECT 33.86 90.234 33.932 90.848 ; 
      RECT 33.536 90.336 33.608 91.368 ; 
      RECT 31.376 87.78 31.448 91.522 ; 
      RECT 31.232 87.78 31.304 91.522 ; 
      RECT 31.088 88.504 31.16 90.776 ; 
      RECT 34.796 92.1 34.868 95.842 ; 
      RECT 34.652 92.1 34.724 95.842 ; 
      RECT 34.508 94.408 34.58 95.698 ; 
      RECT 34.04 95.196 34.112 95.634 ; 
      RECT 34.004 92.23 34.076 93.188 ; 
      RECT 33.86 94.554 33.932 95.168 ; 
      RECT 33.536 94.656 33.608 95.688 ; 
      RECT 31.376 92.1 31.448 95.842 ; 
      RECT 31.232 92.1 31.304 95.842 ; 
      RECT 31.088 92.824 31.16 95.096 ; 
      RECT 34.796 96.42 34.868 100.162 ; 
      RECT 34.652 96.42 34.724 100.162 ; 
      RECT 34.508 98.728 34.58 100.018 ; 
      RECT 34.04 99.516 34.112 99.954 ; 
      RECT 34.004 96.55 34.076 97.508 ; 
      RECT 33.86 98.874 33.932 99.488 ; 
      RECT 33.536 98.976 33.608 100.008 ; 
      RECT 31.376 96.42 31.448 100.162 ; 
      RECT 31.232 96.42 31.304 100.162 ; 
      RECT 31.088 97.144 31.16 99.416 ; 
      RECT 34.796 100.74 34.868 104.482 ; 
      RECT 34.652 100.74 34.724 104.482 ; 
      RECT 34.508 103.048 34.58 104.338 ; 
      RECT 34.04 103.836 34.112 104.274 ; 
      RECT 34.004 100.87 34.076 101.828 ; 
      RECT 33.86 103.194 33.932 103.808 ; 
      RECT 33.536 103.296 33.608 104.328 ; 
      RECT 31.376 100.74 31.448 104.482 ; 
      RECT 31.232 100.74 31.304 104.482 ; 
      RECT 31.088 101.464 31.16 103.736 ; 
      RECT 65.268 119.8 65.34 137.216 ; 
      RECT 65.124 114.54 65.196 114.816 ; 
      RECT 65.124 121.02 65.196 121.352 ; 
      RECT 64.98 104.522 65.052 137.35 ; 
      RECT 64.836 119.93 64.908 122.69 ; 
      RECT 64.836 122.894 64.908 126.84 ; 
      RECT 64.836 127 64.908 129.468 ; 
      RECT 64.692 119.676 64.764 122.4948 ; 
      RECT 64.692 125.508 64.764 130.188 ; 
      RECT 64.548 104.522 64.62 118.908 ; 
      RECT 64.116 104.522 64.188 118.908 ; 
      RECT 63.684 104.522 63.756 118.908 ; 
      RECT 63.252 104.522 63.324 118.908 ; 
      RECT 62.82 104.522 62.892 118.908 ; 
      RECT 62.388 104.522 62.46 118.908 ; 
      RECT 61.956 104.522 62.028 118.908 ; 
      RECT 61.524 104.522 61.596 118.908 ; 
      RECT 61.092 104.522 61.164 118.908 ; 
      RECT 60.66 104.522 60.732 118.908 ; 
      RECT 60.228 104.522 60.3 118.908 ; 
      RECT 59.796 104.522 59.868 118.908 ; 
      RECT 59.364 104.522 59.436 118.908 ; 
      RECT 58.932 104.522 59.004 118.908 ; 
      RECT 58.5 104.522 58.572 118.908 ; 
      RECT 58.068 104.522 58.14 118.908 ; 
      RECT 57.636 104.522 57.708 118.908 ; 
      RECT 57.204 104.522 57.276 118.908 ; 
      RECT 56.772 104.522 56.844 118.908 ; 
      RECT 56.34 104.522 56.412 118.908 ; 
      RECT 55.908 104.522 55.98 118.908 ; 
      RECT 55.476 104.522 55.548 118.908 ; 
      RECT 55.044 104.522 55.116 118.908 ; 
      RECT 54.612 104.522 54.684 118.908 ; 
      RECT 54.18 104.522 54.252 118.908 ; 
      RECT 53.748 104.522 53.82 118.908 ; 
      RECT 53.316 104.522 53.388 118.908 ; 
      RECT 52.884 104.522 52.956 118.908 ; 
      RECT 52.452 104.522 52.524 118.908 ; 
      RECT 52.02 104.522 52.092 118.908 ; 
      RECT 51.588 104.522 51.66 118.908 ; 
      RECT 51.156 104.522 51.228 118.908 ; 
      RECT 50.724 104.522 50.796 118.908 ; 
      RECT 50.292 104.522 50.364 118.908 ; 
      RECT 49.86 104.522 49.932 118.908 ; 
      RECT 49.428 104.522 49.5 118.908 ; 
      RECT 48.996 104.522 49.068 118.908 ; 
      RECT 48.564 104.522 48.636 118.908 ; 
      RECT 48.132 104.522 48.204 118.908 ; 
      RECT 47.7 104.522 47.772 118.908 ; 
      RECT 47.268 104.522 47.34 118.908 ; 
      RECT 46.836 104.522 46.908 118.908 ; 
      RECT 46.404 104.522 46.476 118.908 ; 
      RECT 45.972 104.522 46.044 118.908 ; 
      RECT 45.54 104.522 45.612 118.908 ; 
      RECT 45.108 104.522 45.18 118.908 ; 
      RECT 44.676 104.522 44.748 118.908 ; 
      RECT 44.244 104.522 44.316 118.908 ; 
      RECT 43.812 104.522 43.884 118.908 ; 
      RECT 43.38 104.522 43.452 118.908 ; 
      RECT 42.948 104.522 43.02 118.908 ; 
      RECT 42.516 104.522 42.588 118.908 ; 
      RECT 42.084 104.522 42.156 118.908 ; 
      RECT 41.652 104.522 41.724 118.908 ; 
      RECT 41.22 104.522 41.292 118.908 ; 
      RECT 40.788 104.522 40.86 118.908 ; 
      RECT 40.356 104.522 40.428 118.908 ; 
      RECT 39.924 104.522 39.996 118.908 ; 
      RECT 39.492 104.522 39.564 118.908 ; 
      RECT 39.06 104.522 39.132 118.908 ; 
      RECT 38.628 104.522 38.7 118.908 ; 
      RECT 38.196 104.522 38.268 118.908 ; 
      RECT 38.052 119.942 38.124 122.51 ; 
      RECT 38.052 125.22 38.124 127.348 ; 
      RECT 37.98 107.164 38.052 109.868 ; 
      RECT 37.98 112.852 38.052 114.044 ; 
      RECT 37.98 117.316 38.052 118.364 ; 
      RECT 37.908 119.6 37.98 122.69 ; 
      RECT 37.908 122.8948 37.98 124.86 ; 
      RECT 37.908 125.04 37.98 126.524 ; 
      RECT 37.908 126.828 37.98 129.468 ; 
      RECT 37.764 104.522 37.836 137.35 ; 
      RECT 37.62 121.772 37.692 123.63 ; 
      RECT 37.548 107.596 37.62 110.12 ; 
      RECT 37.548 111.772 37.62 112.532 ; 
      RECT 37.548 115.3 37.62 115.496 ; 
      RECT 37.548 118.228 37.62 118.376 ; 
      RECT 37.476 119.8 37.548 137.198 ; 
      RECT 37.116 106.084 37.188 109.292 ; 
      RECT 37.116 111.484 37.188 113.756 ; 
      RECT 36.972 111.772 37.044 113.252 ; 
      RECT 36.828 109.18 36.9 109.724 ; 
      RECT 36.828 113.14 36.9 114.044 ; 
      RECT 36.828 118.108 36.9 118.364 ; 
      RECT 36.684 109.588 36.756 109.736 ; 
      RECT 36.684 116.092 36.756 116.264 ; 
      RECT 36.684 118.228 36.756 118.376 ; 
      RECT 36.54 110.836 36.612 112.82 ; 
      RECT 36.54 112.996 36.612 113.756 ; 
      RECT 36.54 116.836 36.612 118.076 ; 
      RECT 36.396 110.404 36.468 115.392 ; 
      RECT 36.396 125.956 36.468 128.876 ; 
      RECT 36.396 130.276 36.468 133.196 ; 
      RECT 35.1 109.324 35.172 110.516 ; 
      RECT 35.1 114.076 35.172 114.332 ; 
      RECT 35.1 115.156 35.172 116.996 ; 
      RECT 35.1 119.956 35.172 120.104 ; 
      RECT 35.1 128.116 35.172 129.308 ; 
      RECT 34.956 109.612 35.028 111.632 ; 
      RECT 34.956 112.708 35.028 115.916 ; 
      RECT 34.956 120.088 35.028 121.172 ; 
      RECT 34.956 121.492 35.028 122.396 ; 
      RECT 34.812 109.324 34.884 112.028 ; 
      RECT 34.812 112.42 34.884 113.756 ; 
      RECT 34.812 114.58 34.884 115.124 ; 
      RECT 34.812 117.316 34.884 120.524 ; 
      RECT 34.812 122.26 34.884 122.408 ; 
      RECT 34.812 130.924 34.884 132.26 ; 
      RECT 34.668 110.26 34.74 110.804 ; 
      RECT 34.668 117.82 34.74 121.748 ; 
      RECT 34.668 123.508 34.74 124.7 ; 
      RECT 34.668 130.276 34.74 131.324 ; 
      RECT 34.524 106.516 34.596 107.132 ; 
      RECT 34.524 109.756 34.596 116.9 ; 
      RECT 34.524 121.06 34.596 130.388 ; 
      RECT 34.524 131.212 34.596 135.644 ; 
      RECT 33.372 107.596 33.444 108.644 ; 
      RECT 33.372 109.18 33.444 109.436 ; 
      RECT 33.372 109.756 33.444 110.66 ; 
      RECT 33.372 110.836 33.444 111.596 ; 
      RECT 33.372 111.916 33.444 122.396 ; 
      RECT 33.372 122.572 33.444 127.796 ; 
      RECT 33.372 132.148 33.444 133.196 ; 
      RECT 33.228 111.592 33.3 112.676 ; 
      RECT 33.228 112.996 33.3 116.348 ; 
      RECT 33.228 117.028 33.3 120.38 ; 
      RECT 33.228 120.556 33.3 125.636 ; 
      RECT 33.228 126.46 33.3 127.148 ; 
      RECT 33.228 129.988 33.3 134.276 ; 
      RECT 33.084 111.916 33.156 113 ; 
      RECT 33.084 113.62 33.156 113.768 ; 
      RECT 33.084 116.74 33.156 120.668 ; 
      RECT 33.084 121.636 33.156 123.476 ; 
      RECT 33.084 124.876 33.156 127.832 ; 
      RECT 32.94 108.388 33.012 112.676 ; 
      RECT 32.94 119.044 33.012 119.912 ; 
      RECT 32.94 124.588 33.012 125.78 ; 
      RECT 32.796 110.98 32.868 112.82 ; 
      RECT 32.796 117.316 32.868 118.076 ; 
      RECT 32.796 118.24 32.868 118.388 ; 
      RECT 32.796 119.332 32.868 120.668 ; 
      RECT 32.796 121.204 32.868 126.572 ; 
      RECT 32.796 127 32.868 131.468 ; 
      RECT 32.652 108.676 32.724 109.436 ; 
      RECT 32.652 110.26 32.724 110.804 ; 
      RECT 32.652 111.916 32.724 124.556 ; 
      RECT 32.652 124.876 32.724 126.716 ; 
      RECT 32.652 129.196 32.724 131.036 ; 
      RECT 32.652 134.452 32.724 135.356 ; 
      RECT 32.508 104.628 32.58 105.244 ; 
      RECT 32.508 136.608 32.58 137.272 ; 
      RECT 32.364 104.628 32.436 104.828 ; 
      RECT 32.076 104.628 32.148 104.914 ; 
      RECT 32.076 136.886 32.148 137.35 ; 
      RECT 31.5 110.692 31.572 111.452 ; 
      RECT 31.5 113.644 31.572 115.124 ; 
      RECT 31.5 121.492 31.572 122.396 ; 
      RECT 31.5 123.652 31.572 128.228 ; 
      RECT 31.5 131.356 31.572 133.196 ; 
      RECT 31.5 135.508 31.572 135.656 ; 
      RECT 31.356 106.516 31.428 108.5 ; 
      RECT 31.356 122.836 31.428 122.984 ; 
      RECT 31.356 127.144 31.428 130.388 ; 
      RECT 31.212 108.388 31.284 109.436 ; 
      RECT 31.212 110.548 31.284 111.884 ; 
      RECT 31.212 112.708 31.284 113.108 ; 
      RECT 31.212 116.236 31.284 127.292 ; 
      RECT 31.212 127.828 31.284 128.732 ; 
      RECT 31.068 107.02 31.14 111.596 ; 
      RECT 31.068 125.956 31.14 126.716 ; 
      RECT 31.068 129.172 31.14 129.32 ; 
      RECT 31.068 130.276 31.14 133.484 ; 
      RECT 30.924 110.836 30.996 114.836 ; 
      RECT 30.924 128.596 30.996 128.744 ; 
      RECT 29.484 109.18 29.556 110.804 ; 
      RECT 29.196 109.324 29.268 111.74 ; 
      RECT 29.052 108.676 29.124 108.932 ; 
      RECT 28.908 104.84 28.98 105.044 ; 
      RECT 28.908 117.316 28.98 118.076 ; 
      RECT 28.836 119.8 28.908 137.194 ; 
      RECT 28.548 119.8 28.62 137.198 ; 
      RECT 28.476 106.516 28.548 107.276 ; 
      RECT 28.476 109.612 28.548 118.652 ; 
      RECT 28.404 121.772 28.476 123.63 ; 
      RECT 28.26 104.522 28.332 137.35 ; 
      RECT 28.116 119.6 28.188 122.69 ; 
      RECT 28.116 122.8948 28.188 124.86 ; 
      RECT 28.116 125.04 28.188 126.524 ; 
      RECT 28.116 126.828 28.188 129.468 ; 
      RECT 28.044 106.516 28.116 108.5 ; 
      RECT 28.044 111.628 28.116 113.9 ; 
      RECT 28.044 115.156 28.116 118.076 ; 
      RECT 27.972 119.942 28.044 122.51 ; 
      RECT 27.972 125.22 28.044 127.348 ; 
      RECT 27.828 104.522 27.9 118.908 ; 
      RECT 27.396 104.522 27.468 118.908 ; 
      RECT 26.964 104.522 27.036 118.908 ; 
      RECT 26.532 104.522 26.604 118.908 ; 
      RECT 26.1 104.522 26.172 118.908 ; 
      RECT 25.668 104.522 25.74 118.908 ; 
      RECT 25.236 104.522 25.308 118.908 ; 
      RECT 24.804 104.522 24.876 118.908 ; 
      RECT 24.372 104.522 24.444 118.908 ; 
      RECT 23.94 104.522 24.012 118.908 ; 
      RECT 23.508 104.522 23.58 118.908 ; 
      RECT 23.076 104.522 23.148 118.908 ; 
      RECT 22.644 104.522 22.716 118.908 ; 
      RECT 22.212 104.522 22.284 118.908 ; 
      RECT 21.78 104.522 21.852 118.908 ; 
      RECT 21.348 104.522 21.42 118.908 ; 
      RECT 20.916 104.522 20.988 118.908 ; 
      RECT 20.484 104.522 20.556 118.908 ; 
      RECT 20.052 104.522 20.124 118.908 ; 
      RECT 19.62 104.522 19.692 118.908 ; 
      RECT 19.188 104.522 19.26 118.908 ; 
      RECT 18.756 104.522 18.828 118.908 ; 
      RECT 18.324 104.522 18.396 118.908 ; 
      RECT 17.892 104.522 17.964 118.908 ; 
      RECT 17.46 104.522 17.532 118.908 ; 
      RECT 17.028 104.522 17.1 118.908 ; 
      RECT 16.596 104.522 16.668 118.908 ; 
      RECT 16.164 104.522 16.236 118.908 ; 
      RECT 15.732 104.522 15.804 118.908 ; 
      RECT 15.3 104.522 15.372 118.908 ; 
      RECT 14.868 104.522 14.94 118.908 ; 
      RECT 14.436 104.522 14.508 118.908 ; 
      RECT 14.004 104.522 14.076 118.908 ; 
      RECT 13.572 104.522 13.644 118.908 ; 
      RECT 13.14 104.522 13.212 118.908 ; 
      RECT 12.708 104.522 12.78 118.908 ; 
      RECT 12.276 104.522 12.348 118.908 ; 
      RECT 11.844 104.522 11.916 118.908 ; 
      RECT 11.412 104.522 11.484 118.908 ; 
      RECT 10.98 104.522 11.052 118.908 ; 
      RECT 10.548 104.522 10.62 118.908 ; 
      RECT 10.116 104.522 10.188 118.908 ; 
      RECT 9.684 104.522 9.756 118.908 ; 
      RECT 9.252 104.522 9.324 118.908 ; 
      RECT 8.82 104.522 8.892 118.908 ; 
      RECT 8.388 104.522 8.46 118.908 ; 
      RECT 7.956 104.522 8.028 118.908 ; 
      RECT 7.524 104.522 7.596 118.908 ; 
      RECT 7.092 104.522 7.164 118.908 ; 
      RECT 6.66 104.522 6.732 118.908 ; 
      RECT 6.228 104.522 6.3 118.908 ; 
      RECT 5.796 104.522 5.868 118.908 ; 
      RECT 5.364 104.522 5.436 118.908 ; 
      RECT 4.932 104.522 5.004 118.908 ; 
      RECT 4.5 104.522 4.572 118.908 ; 
      RECT 4.068 104.522 4.14 118.908 ; 
      RECT 3.636 104.522 3.708 118.908 ; 
      RECT 3.204 104.522 3.276 118.908 ; 
      RECT 2.772 104.522 2.844 118.908 ; 
      RECT 2.34 104.522 2.412 118.908 ; 
      RECT 1.908 104.522 1.98 118.908 ; 
      RECT 1.476 104.522 1.548 118.908 ; 
      RECT 1.332 119.676 1.404 122.4948 ; 
      RECT 1.332 125.508 1.404 130.188 ; 
      RECT 1.188 119.93 1.26 122.69 ; 
      RECT 1.188 122.894 1.26 126.84 ; 
      RECT 1.188 127 1.26 129.468 ; 
      RECT 1.044 104.522 1.116 137.35 ; 
      RECT 0.9 114.54 0.972 114.816 ; 
      RECT 0.9 121.02 0.972 121.352 ; 
      RECT 0.756 119.8 0.828 137.216 ; 
        RECT 34.796 137.568 34.868 141.31 ; 
        RECT 34.652 137.568 34.724 141.31 ; 
        RECT 34.508 139.876 34.58 141.166 ; 
        RECT 34.04 140.664 34.112 141.102 ; 
        RECT 34.004 137.698 34.076 138.656 ; 
        RECT 33.86 140.022 33.932 140.636 ; 
        RECT 33.536 140.124 33.608 141.156 ; 
        RECT 31.376 137.568 31.448 141.31 ; 
        RECT 31.232 137.568 31.304 141.31 ; 
        RECT 31.088 138.292 31.16 140.564 ; 
        RECT 34.796 141.888 34.868 145.63 ; 
        RECT 34.652 141.888 34.724 145.63 ; 
        RECT 34.508 144.196 34.58 145.486 ; 
        RECT 34.04 144.984 34.112 145.422 ; 
        RECT 34.004 142.018 34.076 142.976 ; 
        RECT 33.86 144.342 33.932 144.956 ; 
        RECT 33.536 144.444 33.608 145.476 ; 
        RECT 31.376 141.888 31.448 145.63 ; 
        RECT 31.232 141.888 31.304 145.63 ; 
        RECT 31.088 142.612 31.16 144.884 ; 
        RECT 34.796 146.208 34.868 149.95 ; 
        RECT 34.652 146.208 34.724 149.95 ; 
        RECT 34.508 148.516 34.58 149.806 ; 
        RECT 34.04 149.304 34.112 149.742 ; 
        RECT 34.004 146.338 34.076 147.296 ; 
        RECT 33.86 148.662 33.932 149.276 ; 
        RECT 33.536 148.764 33.608 149.796 ; 
        RECT 31.376 146.208 31.448 149.95 ; 
        RECT 31.232 146.208 31.304 149.95 ; 
        RECT 31.088 146.932 31.16 149.204 ; 
        RECT 34.796 150.528 34.868 154.27 ; 
        RECT 34.652 150.528 34.724 154.27 ; 
        RECT 34.508 152.836 34.58 154.126 ; 
        RECT 34.04 153.624 34.112 154.062 ; 
        RECT 34.004 150.658 34.076 151.616 ; 
        RECT 33.86 152.982 33.932 153.596 ; 
        RECT 33.536 153.084 33.608 154.116 ; 
        RECT 31.376 150.528 31.448 154.27 ; 
        RECT 31.232 150.528 31.304 154.27 ; 
        RECT 31.088 151.252 31.16 153.524 ; 
        RECT 34.796 154.848 34.868 158.59 ; 
        RECT 34.652 154.848 34.724 158.59 ; 
        RECT 34.508 157.156 34.58 158.446 ; 
        RECT 34.04 157.944 34.112 158.382 ; 
        RECT 34.004 154.978 34.076 155.936 ; 
        RECT 33.86 157.302 33.932 157.916 ; 
        RECT 33.536 157.404 33.608 158.436 ; 
        RECT 31.376 154.848 31.448 158.59 ; 
        RECT 31.232 154.848 31.304 158.59 ; 
        RECT 31.088 155.572 31.16 157.844 ; 
        RECT 34.796 159.168 34.868 162.91 ; 
        RECT 34.652 159.168 34.724 162.91 ; 
        RECT 34.508 161.476 34.58 162.766 ; 
        RECT 34.04 162.264 34.112 162.702 ; 
        RECT 34.004 159.298 34.076 160.256 ; 
        RECT 33.86 161.622 33.932 162.236 ; 
        RECT 33.536 161.724 33.608 162.756 ; 
        RECT 31.376 159.168 31.448 162.91 ; 
        RECT 31.232 159.168 31.304 162.91 ; 
        RECT 31.088 159.892 31.16 162.164 ; 
        RECT 34.796 163.488 34.868 167.23 ; 
        RECT 34.652 163.488 34.724 167.23 ; 
        RECT 34.508 165.796 34.58 167.086 ; 
        RECT 34.04 166.584 34.112 167.022 ; 
        RECT 34.004 163.618 34.076 164.576 ; 
        RECT 33.86 165.942 33.932 166.556 ; 
        RECT 33.536 166.044 33.608 167.076 ; 
        RECT 31.376 163.488 31.448 167.23 ; 
        RECT 31.232 163.488 31.304 167.23 ; 
        RECT 31.088 164.212 31.16 166.484 ; 
        RECT 34.796 167.808 34.868 171.55 ; 
        RECT 34.652 167.808 34.724 171.55 ; 
        RECT 34.508 170.116 34.58 171.406 ; 
        RECT 34.04 170.904 34.112 171.342 ; 
        RECT 34.004 167.938 34.076 168.896 ; 
        RECT 33.86 170.262 33.932 170.876 ; 
        RECT 33.536 170.364 33.608 171.396 ; 
        RECT 31.376 167.808 31.448 171.55 ; 
        RECT 31.232 167.808 31.304 171.55 ; 
        RECT 31.088 168.532 31.16 170.804 ; 
        RECT 34.796 172.128 34.868 175.87 ; 
        RECT 34.652 172.128 34.724 175.87 ; 
        RECT 34.508 174.436 34.58 175.726 ; 
        RECT 34.04 175.224 34.112 175.662 ; 
        RECT 34.004 172.258 34.076 173.216 ; 
        RECT 33.86 174.582 33.932 175.196 ; 
        RECT 33.536 174.684 33.608 175.716 ; 
        RECT 31.376 172.128 31.448 175.87 ; 
        RECT 31.232 172.128 31.304 175.87 ; 
        RECT 31.088 172.852 31.16 175.124 ; 
        RECT 34.796 176.448 34.868 180.19 ; 
        RECT 34.652 176.448 34.724 180.19 ; 
        RECT 34.508 178.756 34.58 180.046 ; 
        RECT 34.04 179.544 34.112 179.982 ; 
        RECT 34.004 176.578 34.076 177.536 ; 
        RECT 33.86 178.902 33.932 179.516 ; 
        RECT 33.536 179.004 33.608 180.036 ; 
        RECT 31.376 176.448 31.448 180.19 ; 
        RECT 31.232 176.448 31.304 180.19 ; 
        RECT 31.088 177.172 31.16 179.444 ; 
        RECT 34.796 180.768 34.868 184.51 ; 
        RECT 34.652 180.768 34.724 184.51 ; 
        RECT 34.508 183.076 34.58 184.366 ; 
        RECT 34.04 183.864 34.112 184.302 ; 
        RECT 34.004 180.898 34.076 181.856 ; 
        RECT 33.86 183.222 33.932 183.836 ; 
        RECT 33.536 183.324 33.608 184.356 ; 
        RECT 31.376 180.768 31.448 184.51 ; 
        RECT 31.232 180.768 31.304 184.51 ; 
        RECT 31.088 181.492 31.16 183.764 ; 
        RECT 34.796 185.088 34.868 188.83 ; 
        RECT 34.652 185.088 34.724 188.83 ; 
        RECT 34.508 187.396 34.58 188.686 ; 
        RECT 34.04 188.184 34.112 188.622 ; 
        RECT 34.004 185.218 34.076 186.176 ; 
        RECT 33.86 187.542 33.932 188.156 ; 
        RECT 33.536 187.644 33.608 188.676 ; 
        RECT 31.376 185.088 31.448 188.83 ; 
        RECT 31.232 185.088 31.304 188.83 ; 
        RECT 31.088 185.812 31.16 188.084 ; 
        RECT 34.796 189.408 34.868 193.15 ; 
        RECT 34.652 189.408 34.724 193.15 ; 
        RECT 34.508 191.716 34.58 193.006 ; 
        RECT 34.04 192.504 34.112 192.942 ; 
        RECT 34.004 189.538 34.076 190.496 ; 
        RECT 33.86 191.862 33.932 192.476 ; 
        RECT 33.536 191.964 33.608 192.996 ; 
        RECT 31.376 189.408 31.448 193.15 ; 
        RECT 31.232 189.408 31.304 193.15 ; 
        RECT 31.088 190.132 31.16 192.404 ; 
        RECT 34.796 193.728 34.868 197.47 ; 
        RECT 34.652 193.728 34.724 197.47 ; 
        RECT 34.508 196.036 34.58 197.326 ; 
        RECT 34.04 196.824 34.112 197.262 ; 
        RECT 34.004 193.858 34.076 194.816 ; 
        RECT 33.86 196.182 33.932 196.796 ; 
        RECT 33.536 196.284 33.608 197.316 ; 
        RECT 31.376 193.728 31.448 197.47 ; 
        RECT 31.232 193.728 31.304 197.47 ; 
        RECT 31.088 194.452 31.16 196.724 ; 
        RECT 34.796 198.048 34.868 201.79 ; 
        RECT 34.652 198.048 34.724 201.79 ; 
        RECT 34.508 200.356 34.58 201.646 ; 
        RECT 34.04 201.144 34.112 201.582 ; 
        RECT 34.004 198.178 34.076 199.136 ; 
        RECT 33.86 200.502 33.932 201.116 ; 
        RECT 33.536 200.604 33.608 201.636 ; 
        RECT 31.376 198.048 31.448 201.79 ; 
        RECT 31.232 198.048 31.304 201.79 ; 
        RECT 31.088 198.772 31.16 201.044 ; 
        RECT 34.796 202.368 34.868 206.11 ; 
        RECT 34.652 202.368 34.724 206.11 ; 
        RECT 34.508 204.676 34.58 205.966 ; 
        RECT 34.04 205.464 34.112 205.902 ; 
        RECT 34.004 202.498 34.076 203.456 ; 
        RECT 33.86 204.822 33.932 205.436 ; 
        RECT 33.536 204.924 33.608 205.956 ; 
        RECT 31.376 202.368 31.448 206.11 ; 
        RECT 31.232 202.368 31.304 206.11 ; 
        RECT 31.088 203.092 31.16 205.364 ; 
        RECT 34.796 206.688 34.868 210.43 ; 
        RECT 34.652 206.688 34.724 210.43 ; 
        RECT 34.508 208.996 34.58 210.286 ; 
        RECT 34.04 209.784 34.112 210.222 ; 
        RECT 34.004 206.818 34.076 207.776 ; 
        RECT 33.86 209.142 33.932 209.756 ; 
        RECT 33.536 209.244 33.608 210.276 ; 
        RECT 31.376 206.688 31.448 210.43 ; 
        RECT 31.232 206.688 31.304 210.43 ; 
        RECT 31.088 207.412 31.16 209.684 ; 
        RECT 34.796 211.008 34.868 214.75 ; 
        RECT 34.652 211.008 34.724 214.75 ; 
        RECT 34.508 213.316 34.58 214.606 ; 
        RECT 34.04 214.104 34.112 214.542 ; 
        RECT 34.004 211.138 34.076 212.096 ; 
        RECT 33.86 213.462 33.932 214.076 ; 
        RECT 33.536 213.564 33.608 214.596 ; 
        RECT 31.376 211.008 31.448 214.75 ; 
        RECT 31.232 211.008 31.304 214.75 ; 
        RECT 31.088 211.732 31.16 214.004 ; 
        RECT 34.796 215.328 34.868 219.07 ; 
        RECT 34.652 215.328 34.724 219.07 ; 
        RECT 34.508 217.636 34.58 218.926 ; 
        RECT 34.04 218.424 34.112 218.862 ; 
        RECT 34.004 215.458 34.076 216.416 ; 
        RECT 33.86 217.782 33.932 218.396 ; 
        RECT 33.536 217.884 33.608 218.916 ; 
        RECT 31.376 215.328 31.448 219.07 ; 
        RECT 31.232 215.328 31.304 219.07 ; 
        RECT 31.088 216.052 31.16 218.324 ; 
        RECT 34.796 219.648 34.868 223.39 ; 
        RECT 34.652 219.648 34.724 223.39 ; 
        RECT 34.508 221.956 34.58 223.246 ; 
        RECT 34.04 222.744 34.112 223.182 ; 
        RECT 34.004 219.778 34.076 220.736 ; 
        RECT 33.86 222.102 33.932 222.716 ; 
        RECT 33.536 222.204 33.608 223.236 ; 
        RECT 31.376 219.648 31.448 223.39 ; 
        RECT 31.232 219.648 31.304 223.39 ; 
        RECT 31.088 220.372 31.16 222.644 ; 
        RECT 34.796 223.968 34.868 227.71 ; 
        RECT 34.652 223.968 34.724 227.71 ; 
        RECT 34.508 226.276 34.58 227.566 ; 
        RECT 34.04 227.064 34.112 227.502 ; 
        RECT 34.004 224.098 34.076 225.056 ; 
        RECT 33.86 226.422 33.932 227.036 ; 
        RECT 33.536 226.524 33.608 227.556 ; 
        RECT 31.376 223.968 31.448 227.71 ; 
        RECT 31.232 223.968 31.304 227.71 ; 
        RECT 31.088 224.692 31.16 226.964 ; 
        RECT 34.796 228.288 34.868 232.03 ; 
        RECT 34.652 228.288 34.724 232.03 ; 
        RECT 34.508 230.596 34.58 231.886 ; 
        RECT 34.04 231.384 34.112 231.822 ; 
        RECT 34.004 228.418 34.076 229.376 ; 
        RECT 33.86 230.742 33.932 231.356 ; 
        RECT 33.536 230.844 33.608 231.876 ; 
        RECT 31.376 228.288 31.448 232.03 ; 
        RECT 31.232 228.288 31.304 232.03 ; 
        RECT 31.088 229.012 31.16 231.284 ; 
        RECT 34.796 232.608 34.868 236.35 ; 
        RECT 34.652 232.608 34.724 236.35 ; 
        RECT 34.508 234.916 34.58 236.206 ; 
        RECT 34.04 235.704 34.112 236.142 ; 
        RECT 34.004 232.738 34.076 233.696 ; 
        RECT 33.86 235.062 33.932 235.676 ; 
        RECT 33.536 235.164 33.608 236.196 ; 
        RECT 31.376 232.608 31.448 236.35 ; 
        RECT 31.232 232.608 31.304 236.35 ; 
        RECT 31.088 233.332 31.16 235.604 ; 
        RECT 34.796 236.928 34.868 240.67 ; 
        RECT 34.652 236.928 34.724 240.67 ; 
        RECT 34.508 239.236 34.58 240.526 ; 
        RECT 34.04 240.024 34.112 240.462 ; 
        RECT 34.004 237.058 34.076 238.016 ; 
        RECT 33.86 239.382 33.932 239.996 ; 
        RECT 33.536 239.484 33.608 240.516 ; 
        RECT 31.376 236.928 31.448 240.67 ; 
        RECT 31.232 236.928 31.304 240.67 ; 
        RECT 31.088 237.652 31.16 239.924 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 34.564 1.026 35.076 5.4 ; 
      RECT 34.508 3.688 35.076 4.978 ; 
      RECT 33.916 2.596 34.164 5.4 ; 
      RECT 33.86 3.834 34.164 4.448 ; 
      RECT 33.916 1.026 34.02 5.4 ; 
      RECT 33.916 1.51 34.076 2.468 ; 
      RECT 33.916 1.026 34.164 1.382 ; 
      RECT 32.728 2.828 33.552 5.4 ; 
      RECT 33.448 1.026 33.552 5.4 ; 
      RECT 32.728 3.936 33.608 4.968 ; 
      RECT 32.728 1.026 33.12 5.4 ; 
      RECT 31.06 1.026 31.392 5.4 ; 
      RECT 31.06 1.38 31.448 5.122 ; 
      RECT 65.776 1.026 66.116 5.4 ; 
      RECT 65.2 1.026 65.304 5.4 ; 
      RECT 64.768 1.026 64.872 5.4 ; 
      RECT 64.336 1.026 64.44 5.4 ; 
      RECT 63.904 1.026 64.008 5.4 ; 
      RECT 63.472 1.026 63.576 5.4 ; 
      RECT 63.04 1.026 63.144 5.4 ; 
      RECT 62.608 1.026 62.712 5.4 ; 
      RECT 62.176 1.026 62.28 5.4 ; 
      RECT 61.744 1.026 61.848 5.4 ; 
      RECT 61.312 1.026 61.416 5.4 ; 
      RECT 60.88 1.026 60.984 5.4 ; 
      RECT 60.448 1.026 60.552 5.4 ; 
      RECT 60.016 1.026 60.12 5.4 ; 
      RECT 59.584 1.026 59.688 5.4 ; 
      RECT 59.152 1.026 59.256 5.4 ; 
      RECT 58.72 1.026 58.824 5.4 ; 
      RECT 58.288 1.026 58.392 5.4 ; 
      RECT 57.856 1.026 57.96 5.4 ; 
      RECT 57.424 1.026 57.528 5.4 ; 
      RECT 56.992 1.026 57.096 5.4 ; 
      RECT 56.56 1.026 56.664 5.4 ; 
      RECT 56.128 1.026 56.232 5.4 ; 
      RECT 55.696 1.026 55.8 5.4 ; 
      RECT 55.264 1.026 55.368 5.4 ; 
      RECT 54.832 1.026 54.936 5.4 ; 
      RECT 54.4 1.026 54.504 5.4 ; 
      RECT 53.968 1.026 54.072 5.4 ; 
      RECT 53.536 1.026 53.64 5.4 ; 
      RECT 53.104 1.026 53.208 5.4 ; 
      RECT 52.672 1.026 52.776 5.4 ; 
      RECT 52.24 1.026 52.344 5.4 ; 
      RECT 51.808 1.026 51.912 5.4 ; 
      RECT 51.376 1.026 51.48 5.4 ; 
      RECT 50.944 1.026 51.048 5.4 ; 
      RECT 50.512 1.026 50.616 5.4 ; 
      RECT 50.08 1.026 50.184 5.4 ; 
      RECT 49.648 1.026 49.752 5.4 ; 
      RECT 49.216 1.026 49.32 5.4 ; 
      RECT 48.784 1.026 48.888 5.4 ; 
      RECT 48.352 1.026 48.456 5.4 ; 
      RECT 47.92 1.026 48.024 5.4 ; 
      RECT 47.488 1.026 47.592 5.4 ; 
      RECT 47.056 1.026 47.16 5.4 ; 
      RECT 46.624 1.026 46.728 5.4 ; 
      RECT 46.192 1.026 46.296 5.4 ; 
      RECT 45.76 1.026 45.864 5.4 ; 
      RECT 45.328 1.026 45.432 5.4 ; 
      RECT 44.896 1.026 45 5.4 ; 
      RECT 44.464 1.026 44.568 5.4 ; 
      RECT 44.032 1.026 44.136 5.4 ; 
      RECT 43.6 1.026 43.704 5.4 ; 
      RECT 43.168 1.026 43.272 5.4 ; 
      RECT 42.736 1.026 42.84 5.4 ; 
      RECT 42.304 1.026 42.408 5.4 ; 
      RECT 41.872 1.026 41.976 5.4 ; 
      RECT 41.44 1.026 41.544 5.4 ; 
      RECT 41.008 1.026 41.112 5.4 ; 
      RECT 40.576 1.026 40.68 5.4 ; 
      RECT 40.144 1.026 40.248 5.4 ; 
      RECT 39.712 1.026 39.816 5.4 ; 
      RECT 39.28 1.026 39.384 5.4 ; 
      RECT 38.848 1.026 38.952 5.4 ; 
      RECT 38.416 1.026 38.52 5.4 ; 
      RECT 37.984 1.026 38.088 5.4 ; 
      RECT 37.552 1.026 37.656 5.4 ; 
      RECT 36.7 1.026 37.008 5.4 ; 
      RECT 29.128 1.026 29.436 5.4 ; 
      RECT 28.48 1.026 28.584 5.4 ; 
      RECT 28.048 1.026 28.152 5.4 ; 
      RECT 27.616 1.026 27.72 5.4 ; 
      RECT 27.184 1.026 27.288 5.4 ; 
      RECT 26.752 1.026 26.856 5.4 ; 
      RECT 26.32 1.026 26.424 5.4 ; 
      RECT 25.888 1.026 25.992 5.4 ; 
      RECT 25.456 1.026 25.56 5.4 ; 
      RECT 25.024 1.026 25.128 5.4 ; 
      RECT 24.592 1.026 24.696 5.4 ; 
      RECT 24.16 1.026 24.264 5.4 ; 
      RECT 23.728 1.026 23.832 5.4 ; 
      RECT 23.296 1.026 23.4 5.4 ; 
      RECT 22.864 1.026 22.968 5.4 ; 
      RECT 22.432 1.026 22.536 5.4 ; 
      RECT 22 1.026 22.104 5.4 ; 
      RECT 21.568 1.026 21.672 5.4 ; 
      RECT 21.136 1.026 21.24 5.4 ; 
      RECT 20.704 1.026 20.808 5.4 ; 
      RECT 20.272 1.026 20.376 5.4 ; 
      RECT 19.84 1.026 19.944 5.4 ; 
      RECT 19.408 1.026 19.512 5.4 ; 
      RECT 18.976 1.026 19.08 5.4 ; 
      RECT 18.544 1.026 18.648 5.4 ; 
      RECT 18.112 1.026 18.216 5.4 ; 
      RECT 17.68 1.026 17.784 5.4 ; 
      RECT 17.248 1.026 17.352 5.4 ; 
      RECT 16.816 1.026 16.92 5.4 ; 
      RECT 16.384 1.026 16.488 5.4 ; 
      RECT 15.952 1.026 16.056 5.4 ; 
      RECT 15.52 1.026 15.624 5.4 ; 
      RECT 15.088 1.026 15.192 5.4 ; 
      RECT 14.656 1.026 14.76 5.4 ; 
      RECT 14.224 1.026 14.328 5.4 ; 
      RECT 13.792 1.026 13.896 5.4 ; 
      RECT 13.36 1.026 13.464 5.4 ; 
      RECT 12.928 1.026 13.032 5.4 ; 
      RECT 12.496 1.026 12.6 5.4 ; 
      RECT 12.064 1.026 12.168 5.4 ; 
      RECT 11.632 1.026 11.736 5.4 ; 
      RECT 11.2 1.026 11.304 5.4 ; 
      RECT 10.768 1.026 10.872 5.4 ; 
      RECT 10.336 1.026 10.44 5.4 ; 
      RECT 9.904 1.026 10.008 5.4 ; 
      RECT 9.472 1.026 9.576 5.4 ; 
      RECT 9.04 1.026 9.144 5.4 ; 
      RECT 8.608 1.026 8.712 5.4 ; 
      RECT 8.176 1.026 8.28 5.4 ; 
      RECT 7.744 1.026 7.848 5.4 ; 
      RECT 7.312 1.026 7.416 5.4 ; 
      RECT 6.88 1.026 6.984 5.4 ; 
      RECT 6.448 1.026 6.552 5.4 ; 
      RECT 6.016 1.026 6.12 5.4 ; 
      RECT 5.584 1.026 5.688 5.4 ; 
      RECT 5.152 1.026 5.256 5.4 ; 
      RECT 4.72 1.026 4.824 5.4 ; 
      RECT 4.288 1.026 4.392 5.4 ; 
      RECT 3.856 1.026 3.96 5.4 ; 
      RECT 3.424 1.026 3.528 5.4 ; 
      RECT 2.992 1.026 3.096 5.4 ; 
      RECT 2.56 1.026 2.664 5.4 ; 
      RECT 2.128 1.026 2.232 5.4 ; 
      RECT 1.696 1.026 1.8 5.4 ; 
      RECT 1.264 1.026 1.368 5.4 ; 
      RECT 0.832 1.026 0.936 5.4 ; 
      RECT 0.02 1.026 0.36 5.4 ; 
      RECT 34.564 5.346 35.076 9.72 ; 
      RECT 34.508 8.008 35.076 9.298 ; 
      RECT 33.916 6.916 34.164 9.72 ; 
      RECT 33.86 8.154 34.164 8.768 ; 
      RECT 33.916 5.346 34.02 9.72 ; 
      RECT 33.916 5.83 34.076 6.788 ; 
      RECT 33.916 5.346 34.164 5.702 ; 
      RECT 32.728 7.148 33.552 9.72 ; 
      RECT 33.448 5.346 33.552 9.72 ; 
      RECT 32.728 8.256 33.608 9.288 ; 
      RECT 32.728 5.346 33.12 9.72 ; 
      RECT 31.06 5.346 31.392 9.72 ; 
      RECT 31.06 5.7 31.448 9.442 ; 
      RECT 65.776 5.346 66.116 9.72 ; 
      RECT 65.2 5.346 65.304 9.72 ; 
      RECT 64.768 5.346 64.872 9.72 ; 
      RECT 64.336 5.346 64.44 9.72 ; 
      RECT 63.904 5.346 64.008 9.72 ; 
      RECT 63.472 5.346 63.576 9.72 ; 
      RECT 63.04 5.346 63.144 9.72 ; 
      RECT 62.608 5.346 62.712 9.72 ; 
      RECT 62.176 5.346 62.28 9.72 ; 
      RECT 61.744 5.346 61.848 9.72 ; 
      RECT 61.312 5.346 61.416 9.72 ; 
      RECT 60.88 5.346 60.984 9.72 ; 
      RECT 60.448 5.346 60.552 9.72 ; 
      RECT 60.016 5.346 60.12 9.72 ; 
      RECT 59.584 5.346 59.688 9.72 ; 
      RECT 59.152 5.346 59.256 9.72 ; 
      RECT 58.72 5.346 58.824 9.72 ; 
      RECT 58.288 5.346 58.392 9.72 ; 
      RECT 57.856 5.346 57.96 9.72 ; 
      RECT 57.424 5.346 57.528 9.72 ; 
      RECT 56.992 5.346 57.096 9.72 ; 
      RECT 56.56 5.346 56.664 9.72 ; 
      RECT 56.128 5.346 56.232 9.72 ; 
      RECT 55.696 5.346 55.8 9.72 ; 
      RECT 55.264 5.346 55.368 9.72 ; 
      RECT 54.832 5.346 54.936 9.72 ; 
      RECT 54.4 5.346 54.504 9.72 ; 
      RECT 53.968 5.346 54.072 9.72 ; 
      RECT 53.536 5.346 53.64 9.72 ; 
      RECT 53.104 5.346 53.208 9.72 ; 
      RECT 52.672 5.346 52.776 9.72 ; 
      RECT 52.24 5.346 52.344 9.72 ; 
      RECT 51.808 5.346 51.912 9.72 ; 
      RECT 51.376 5.346 51.48 9.72 ; 
      RECT 50.944 5.346 51.048 9.72 ; 
      RECT 50.512 5.346 50.616 9.72 ; 
      RECT 50.08 5.346 50.184 9.72 ; 
      RECT 49.648 5.346 49.752 9.72 ; 
      RECT 49.216 5.346 49.32 9.72 ; 
      RECT 48.784 5.346 48.888 9.72 ; 
      RECT 48.352 5.346 48.456 9.72 ; 
      RECT 47.92 5.346 48.024 9.72 ; 
      RECT 47.488 5.346 47.592 9.72 ; 
      RECT 47.056 5.346 47.16 9.72 ; 
      RECT 46.624 5.346 46.728 9.72 ; 
      RECT 46.192 5.346 46.296 9.72 ; 
      RECT 45.76 5.346 45.864 9.72 ; 
      RECT 45.328 5.346 45.432 9.72 ; 
      RECT 44.896 5.346 45 9.72 ; 
      RECT 44.464 5.346 44.568 9.72 ; 
      RECT 44.032 5.346 44.136 9.72 ; 
      RECT 43.6 5.346 43.704 9.72 ; 
      RECT 43.168 5.346 43.272 9.72 ; 
      RECT 42.736 5.346 42.84 9.72 ; 
      RECT 42.304 5.346 42.408 9.72 ; 
      RECT 41.872 5.346 41.976 9.72 ; 
      RECT 41.44 5.346 41.544 9.72 ; 
      RECT 41.008 5.346 41.112 9.72 ; 
      RECT 40.576 5.346 40.68 9.72 ; 
      RECT 40.144 5.346 40.248 9.72 ; 
      RECT 39.712 5.346 39.816 9.72 ; 
      RECT 39.28 5.346 39.384 9.72 ; 
      RECT 38.848 5.346 38.952 9.72 ; 
      RECT 38.416 5.346 38.52 9.72 ; 
      RECT 37.984 5.346 38.088 9.72 ; 
      RECT 37.552 5.346 37.656 9.72 ; 
      RECT 36.7 5.346 37.008 9.72 ; 
      RECT 29.128 5.346 29.436 9.72 ; 
      RECT 28.48 5.346 28.584 9.72 ; 
      RECT 28.048 5.346 28.152 9.72 ; 
      RECT 27.616 5.346 27.72 9.72 ; 
      RECT 27.184 5.346 27.288 9.72 ; 
      RECT 26.752 5.346 26.856 9.72 ; 
      RECT 26.32 5.346 26.424 9.72 ; 
      RECT 25.888 5.346 25.992 9.72 ; 
      RECT 25.456 5.346 25.56 9.72 ; 
      RECT 25.024 5.346 25.128 9.72 ; 
      RECT 24.592 5.346 24.696 9.72 ; 
      RECT 24.16 5.346 24.264 9.72 ; 
      RECT 23.728 5.346 23.832 9.72 ; 
      RECT 23.296 5.346 23.4 9.72 ; 
      RECT 22.864 5.346 22.968 9.72 ; 
      RECT 22.432 5.346 22.536 9.72 ; 
      RECT 22 5.346 22.104 9.72 ; 
      RECT 21.568 5.346 21.672 9.72 ; 
      RECT 21.136 5.346 21.24 9.72 ; 
      RECT 20.704 5.346 20.808 9.72 ; 
      RECT 20.272 5.346 20.376 9.72 ; 
      RECT 19.84 5.346 19.944 9.72 ; 
      RECT 19.408 5.346 19.512 9.72 ; 
      RECT 18.976 5.346 19.08 9.72 ; 
      RECT 18.544 5.346 18.648 9.72 ; 
      RECT 18.112 5.346 18.216 9.72 ; 
      RECT 17.68 5.346 17.784 9.72 ; 
      RECT 17.248 5.346 17.352 9.72 ; 
      RECT 16.816 5.346 16.92 9.72 ; 
      RECT 16.384 5.346 16.488 9.72 ; 
      RECT 15.952 5.346 16.056 9.72 ; 
      RECT 15.52 5.346 15.624 9.72 ; 
      RECT 15.088 5.346 15.192 9.72 ; 
      RECT 14.656 5.346 14.76 9.72 ; 
      RECT 14.224 5.346 14.328 9.72 ; 
      RECT 13.792 5.346 13.896 9.72 ; 
      RECT 13.36 5.346 13.464 9.72 ; 
      RECT 12.928 5.346 13.032 9.72 ; 
      RECT 12.496 5.346 12.6 9.72 ; 
      RECT 12.064 5.346 12.168 9.72 ; 
      RECT 11.632 5.346 11.736 9.72 ; 
      RECT 11.2 5.346 11.304 9.72 ; 
      RECT 10.768 5.346 10.872 9.72 ; 
      RECT 10.336 5.346 10.44 9.72 ; 
      RECT 9.904 5.346 10.008 9.72 ; 
      RECT 9.472 5.346 9.576 9.72 ; 
      RECT 9.04 5.346 9.144 9.72 ; 
      RECT 8.608 5.346 8.712 9.72 ; 
      RECT 8.176 5.346 8.28 9.72 ; 
      RECT 7.744 5.346 7.848 9.72 ; 
      RECT 7.312 5.346 7.416 9.72 ; 
      RECT 6.88 5.346 6.984 9.72 ; 
      RECT 6.448 5.346 6.552 9.72 ; 
      RECT 6.016 5.346 6.12 9.72 ; 
      RECT 5.584 5.346 5.688 9.72 ; 
      RECT 5.152 5.346 5.256 9.72 ; 
      RECT 4.72 5.346 4.824 9.72 ; 
      RECT 4.288 5.346 4.392 9.72 ; 
      RECT 3.856 5.346 3.96 9.72 ; 
      RECT 3.424 5.346 3.528 9.72 ; 
      RECT 2.992 5.346 3.096 9.72 ; 
      RECT 2.56 5.346 2.664 9.72 ; 
      RECT 2.128 5.346 2.232 9.72 ; 
      RECT 1.696 5.346 1.8 9.72 ; 
      RECT 1.264 5.346 1.368 9.72 ; 
      RECT 0.832 5.346 0.936 9.72 ; 
      RECT 0.02 5.346 0.36 9.72 ; 
      RECT 34.564 9.666 35.076 14.04 ; 
      RECT 34.508 12.328 35.076 13.618 ; 
      RECT 33.916 11.236 34.164 14.04 ; 
      RECT 33.86 12.474 34.164 13.088 ; 
      RECT 33.916 9.666 34.02 14.04 ; 
      RECT 33.916 10.15 34.076 11.108 ; 
      RECT 33.916 9.666 34.164 10.022 ; 
      RECT 32.728 11.468 33.552 14.04 ; 
      RECT 33.448 9.666 33.552 14.04 ; 
      RECT 32.728 12.576 33.608 13.608 ; 
      RECT 32.728 9.666 33.12 14.04 ; 
      RECT 31.06 9.666 31.392 14.04 ; 
      RECT 31.06 10.02 31.448 13.762 ; 
      RECT 65.776 9.666 66.116 14.04 ; 
      RECT 65.2 9.666 65.304 14.04 ; 
      RECT 64.768 9.666 64.872 14.04 ; 
      RECT 64.336 9.666 64.44 14.04 ; 
      RECT 63.904 9.666 64.008 14.04 ; 
      RECT 63.472 9.666 63.576 14.04 ; 
      RECT 63.04 9.666 63.144 14.04 ; 
      RECT 62.608 9.666 62.712 14.04 ; 
      RECT 62.176 9.666 62.28 14.04 ; 
      RECT 61.744 9.666 61.848 14.04 ; 
      RECT 61.312 9.666 61.416 14.04 ; 
      RECT 60.88 9.666 60.984 14.04 ; 
      RECT 60.448 9.666 60.552 14.04 ; 
      RECT 60.016 9.666 60.12 14.04 ; 
      RECT 59.584 9.666 59.688 14.04 ; 
      RECT 59.152 9.666 59.256 14.04 ; 
      RECT 58.72 9.666 58.824 14.04 ; 
      RECT 58.288 9.666 58.392 14.04 ; 
      RECT 57.856 9.666 57.96 14.04 ; 
      RECT 57.424 9.666 57.528 14.04 ; 
      RECT 56.992 9.666 57.096 14.04 ; 
      RECT 56.56 9.666 56.664 14.04 ; 
      RECT 56.128 9.666 56.232 14.04 ; 
      RECT 55.696 9.666 55.8 14.04 ; 
      RECT 55.264 9.666 55.368 14.04 ; 
      RECT 54.832 9.666 54.936 14.04 ; 
      RECT 54.4 9.666 54.504 14.04 ; 
      RECT 53.968 9.666 54.072 14.04 ; 
      RECT 53.536 9.666 53.64 14.04 ; 
      RECT 53.104 9.666 53.208 14.04 ; 
      RECT 52.672 9.666 52.776 14.04 ; 
      RECT 52.24 9.666 52.344 14.04 ; 
      RECT 51.808 9.666 51.912 14.04 ; 
      RECT 51.376 9.666 51.48 14.04 ; 
      RECT 50.944 9.666 51.048 14.04 ; 
      RECT 50.512 9.666 50.616 14.04 ; 
      RECT 50.08 9.666 50.184 14.04 ; 
      RECT 49.648 9.666 49.752 14.04 ; 
      RECT 49.216 9.666 49.32 14.04 ; 
      RECT 48.784 9.666 48.888 14.04 ; 
      RECT 48.352 9.666 48.456 14.04 ; 
      RECT 47.92 9.666 48.024 14.04 ; 
      RECT 47.488 9.666 47.592 14.04 ; 
      RECT 47.056 9.666 47.16 14.04 ; 
      RECT 46.624 9.666 46.728 14.04 ; 
      RECT 46.192 9.666 46.296 14.04 ; 
      RECT 45.76 9.666 45.864 14.04 ; 
      RECT 45.328 9.666 45.432 14.04 ; 
      RECT 44.896 9.666 45 14.04 ; 
      RECT 44.464 9.666 44.568 14.04 ; 
      RECT 44.032 9.666 44.136 14.04 ; 
      RECT 43.6 9.666 43.704 14.04 ; 
      RECT 43.168 9.666 43.272 14.04 ; 
      RECT 42.736 9.666 42.84 14.04 ; 
      RECT 42.304 9.666 42.408 14.04 ; 
      RECT 41.872 9.666 41.976 14.04 ; 
      RECT 41.44 9.666 41.544 14.04 ; 
      RECT 41.008 9.666 41.112 14.04 ; 
      RECT 40.576 9.666 40.68 14.04 ; 
      RECT 40.144 9.666 40.248 14.04 ; 
      RECT 39.712 9.666 39.816 14.04 ; 
      RECT 39.28 9.666 39.384 14.04 ; 
      RECT 38.848 9.666 38.952 14.04 ; 
      RECT 38.416 9.666 38.52 14.04 ; 
      RECT 37.984 9.666 38.088 14.04 ; 
      RECT 37.552 9.666 37.656 14.04 ; 
      RECT 36.7 9.666 37.008 14.04 ; 
      RECT 29.128 9.666 29.436 14.04 ; 
      RECT 28.48 9.666 28.584 14.04 ; 
      RECT 28.048 9.666 28.152 14.04 ; 
      RECT 27.616 9.666 27.72 14.04 ; 
      RECT 27.184 9.666 27.288 14.04 ; 
      RECT 26.752 9.666 26.856 14.04 ; 
      RECT 26.32 9.666 26.424 14.04 ; 
      RECT 25.888 9.666 25.992 14.04 ; 
      RECT 25.456 9.666 25.56 14.04 ; 
      RECT 25.024 9.666 25.128 14.04 ; 
      RECT 24.592 9.666 24.696 14.04 ; 
      RECT 24.16 9.666 24.264 14.04 ; 
      RECT 23.728 9.666 23.832 14.04 ; 
      RECT 23.296 9.666 23.4 14.04 ; 
      RECT 22.864 9.666 22.968 14.04 ; 
      RECT 22.432 9.666 22.536 14.04 ; 
      RECT 22 9.666 22.104 14.04 ; 
      RECT 21.568 9.666 21.672 14.04 ; 
      RECT 21.136 9.666 21.24 14.04 ; 
      RECT 20.704 9.666 20.808 14.04 ; 
      RECT 20.272 9.666 20.376 14.04 ; 
      RECT 19.84 9.666 19.944 14.04 ; 
      RECT 19.408 9.666 19.512 14.04 ; 
      RECT 18.976 9.666 19.08 14.04 ; 
      RECT 18.544 9.666 18.648 14.04 ; 
      RECT 18.112 9.666 18.216 14.04 ; 
      RECT 17.68 9.666 17.784 14.04 ; 
      RECT 17.248 9.666 17.352 14.04 ; 
      RECT 16.816 9.666 16.92 14.04 ; 
      RECT 16.384 9.666 16.488 14.04 ; 
      RECT 15.952 9.666 16.056 14.04 ; 
      RECT 15.52 9.666 15.624 14.04 ; 
      RECT 15.088 9.666 15.192 14.04 ; 
      RECT 14.656 9.666 14.76 14.04 ; 
      RECT 14.224 9.666 14.328 14.04 ; 
      RECT 13.792 9.666 13.896 14.04 ; 
      RECT 13.36 9.666 13.464 14.04 ; 
      RECT 12.928 9.666 13.032 14.04 ; 
      RECT 12.496 9.666 12.6 14.04 ; 
      RECT 12.064 9.666 12.168 14.04 ; 
      RECT 11.632 9.666 11.736 14.04 ; 
      RECT 11.2 9.666 11.304 14.04 ; 
      RECT 10.768 9.666 10.872 14.04 ; 
      RECT 10.336 9.666 10.44 14.04 ; 
      RECT 9.904 9.666 10.008 14.04 ; 
      RECT 9.472 9.666 9.576 14.04 ; 
      RECT 9.04 9.666 9.144 14.04 ; 
      RECT 8.608 9.666 8.712 14.04 ; 
      RECT 8.176 9.666 8.28 14.04 ; 
      RECT 7.744 9.666 7.848 14.04 ; 
      RECT 7.312 9.666 7.416 14.04 ; 
      RECT 6.88 9.666 6.984 14.04 ; 
      RECT 6.448 9.666 6.552 14.04 ; 
      RECT 6.016 9.666 6.12 14.04 ; 
      RECT 5.584 9.666 5.688 14.04 ; 
      RECT 5.152 9.666 5.256 14.04 ; 
      RECT 4.72 9.666 4.824 14.04 ; 
      RECT 4.288 9.666 4.392 14.04 ; 
      RECT 3.856 9.666 3.96 14.04 ; 
      RECT 3.424 9.666 3.528 14.04 ; 
      RECT 2.992 9.666 3.096 14.04 ; 
      RECT 2.56 9.666 2.664 14.04 ; 
      RECT 2.128 9.666 2.232 14.04 ; 
      RECT 1.696 9.666 1.8 14.04 ; 
      RECT 1.264 9.666 1.368 14.04 ; 
      RECT 0.832 9.666 0.936 14.04 ; 
      RECT 0.02 9.666 0.36 14.04 ; 
      RECT 34.564 13.986 35.076 18.36 ; 
      RECT 34.508 16.648 35.076 17.938 ; 
      RECT 33.916 15.556 34.164 18.36 ; 
      RECT 33.86 16.794 34.164 17.408 ; 
      RECT 33.916 13.986 34.02 18.36 ; 
      RECT 33.916 14.47 34.076 15.428 ; 
      RECT 33.916 13.986 34.164 14.342 ; 
      RECT 32.728 15.788 33.552 18.36 ; 
      RECT 33.448 13.986 33.552 18.36 ; 
      RECT 32.728 16.896 33.608 17.928 ; 
      RECT 32.728 13.986 33.12 18.36 ; 
      RECT 31.06 13.986 31.392 18.36 ; 
      RECT 31.06 14.34 31.448 18.082 ; 
      RECT 65.776 13.986 66.116 18.36 ; 
      RECT 65.2 13.986 65.304 18.36 ; 
      RECT 64.768 13.986 64.872 18.36 ; 
      RECT 64.336 13.986 64.44 18.36 ; 
      RECT 63.904 13.986 64.008 18.36 ; 
      RECT 63.472 13.986 63.576 18.36 ; 
      RECT 63.04 13.986 63.144 18.36 ; 
      RECT 62.608 13.986 62.712 18.36 ; 
      RECT 62.176 13.986 62.28 18.36 ; 
      RECT 61.744 13.986 61.848 18.36 ; 
      RECT 61.312 13.986 61.416 18.36 ; 
      RECT 60.88 13.986 60.984 18.36 ; 
      RECT 60.448 13.986 60.552 18.36 ; 
      RECT 60.016 13.986 60.12 18.36 ; 
      RECT 59.584 13.986 59.688 18.36 ; 
      RECT 59.152 13.986 59.256 18.36 ; 
      RECT 58.72 13.986 58.824 18.36 ; 
      RECT 58.288 13.986 58.392 18.36 ; 
      RECT 57.856 13.986 57.96 18.36 ; 
      RECT 57.424 13.986 57.528 18.36 ; 
      RECT 56.992 13.986 57.096 18.36 ; 
      RECT 56.56 13.986 56.664 18.36 ; 
      RECT 56.128 13.986 56.232 18.36 ; 
      RECT 55.696 13.986 55.8 18.36 ; 
      RECT 55.264 13.986 55.368 18.36 ; 
      RECT 54.832 13.986 54.936 18.36 ; 
      RECT 54.4 13.986 54.504 18.36 ; 
      RECT 53.968 13.986 54.072 18.36 ; 
      RECT 53.536 13.986 53.64 18.36 ; 
      RECT 53.104 13.986 53.208 18.36 ; 
      RECT 52.672 13.986 52.776 18.36 ; 
      RECT 52.24 13.986 52.344 18.36 ; 
      RECT 51.808 13.986 51.912 18.36 ; 
      RECT 51.376 13.986 51.48 18.36 ; 
      RECT 50.944 13.986 51.048 18.36 ; 
      RECT 50.512 13.986 50.616 18.36 ; 
      RECT 50.08 13.986 50.184 18.36 ; 
      RECT 49.648 13.986 49.752 18.36 ; 
      RECT 49.216 13.986 49.32 18.36 ; 
      RECT 48.784 13.986 48.888 18.36 ; 
      RECT 48.352 13.986 48.456 18.36 ; 
      RECT 47.92 13.986 48.024 18.36 ; 
      RECT 47.488 13.986 47.592 18.36 ; 
      RECT 47.056 13.986 47.16 18.36 ; 
      RECT 46.624 13.986 46.728 18.36 ; 
      RECT 46.192 13.986 46.296 18.36 ; 
      RECT 45.76 13.986 45.864 18.36 ; 
      RECT 45.328 13.986 45.432 18.36 ; 
      RECT 44.896 13.986 45 18.36 ; 
      RECT 44.464 13.986 44.568 18.36 ; 
      RECT 44.032 13.986 44.136 18.36 ; 
      RECT 43.6 13.986 43.704 18.36 ; 
      RECT 43.168 13.986 43.272 18.36 ; 
      RECT 42.736 13.986 42.84 18.36 ; 
      RECT 42.304 13.986 42.408 18.36 ; 
      RECT 41.872 13.986 41.976 18.36 ; 
      RECT 41.44 13.986 41.544 18.36 ; 
      RECT 41.008 13.986 41.112 18.36 ; 
      RECT 40.576 13.986 40.68 18.36 ; 
      RECT 40.144 13.986 40.248 18.36 ; 
      RECT 39.712 13.986 39.816 18.36 ; 
      RECT 39.28 13.986 39.384 18.36 ; 
      RECT 38.848 13.986 38.952 18.36 ; 
      RECT 38.416 13.986 38.52 18.36 ; 
      RECT 37.984 13.986 38.088 18.36 ; 
      RECT 37.552 13.986 37.656 18.36 ; 
      RECT 36.7 13.986 37.008 18.36 ; 
      RECT 29.128 13.986 29.436 18.36 ; 
      RECT 28.48 13.986 28.584 18.36 ; 
      RECT 28.048 13.986 28.152 18.36 ; 
      RECT 27.616 13.986 27.72 18.36 ; 
      RECT 27.184 13.986 27.288 18.36 ; 
      RECT 26.752 13.986 26.856 18.36 ; 
      RECT 26.32 13.986 26.424 18.36 ; 
      RECT 25.888 13.986 25.992 18.36 ; 
      RECT 25.456 13.986 25.56 18.36 ; 
      RECT 25.024 13.986 25.128 18.36 ; 
      RECT 24.592 13.986 24.696 18.36 ; 
      RECT 24.16 13.986 24.264 18.36 ; 
      RECT 23.728 13.986 23.832 18.36 ; 
      RECT 23.296 13.986 23.4 18.36 ; 
      RECT 22.864 13.986 22.968 18.36 ; 
      RECT 22.432 13.986 22.536 18.36 ; 
      RECT 22 13.986 22.104 18.36 ; 
      RECT 21.568 13.986 21.672 18.36 ; 
      RECT 21.136 13.986 21.24 18.36 ; 
      RECT 20.704 13.986 20.808 18.36 ; 
      RECT 20.272 13.986 20.376 18.36 ; 
      RECT 19.84 13.986 19.944 18.36 ; 
      RECT 19.408 13.986 19.512 18.36 ; 
      RECT 18.976 13.986 19.08 18.36 ; 
      RECT 18.544 13.986 18.648 18.36 ; 
      RECT 18.112 13.986 18.216 18.36 ; 
      RECT 17.68 13.986 17.784 18.36 ; 
      RECT 17.248 13.986 17.352 18.36 ; 
      RECT 16.816 13.986 16.92 18.36 ; 
      RECT 16.384 13.986 16.488 18.36 ; 
      RECT 15.952 13.986 16.056 18.36 ; 
      RECT 15.52 13.986 15.624 18.36 ; 
      RECT 15.088 13.986 15.192 18.36 ; 
      RECT 14.656 13.986 14.76 18.36 ; 
      RECT 14.224 13.986 14.328 18.36 ; 
      RECT 13.792 13.986 13.896 18.36 ; 
      RECT 13.36 13.986 13.464 18.36 ; 
      RECT 12.928 13.986 13.032 18.36 ; 
      RECT 12.496 13.986 12.6 18.36 ; 
      RECT 12.064 13.986 12.168 18.36 ; 
      RECT 11.632 13.986 11.736 18.36 ; 
      RECT 11.2 13.986 11.304 18.36 ; 
      RECT 10.768 13.986 10.872 18.36 ; 
      RECT 10.336 13.986 10.44 18.36 ; 
      RECT 9.904 13.986 10.008 18.36 ; 
      RECT 9.472 13.986 9.576 18.36 ; 
      RECT 9.04 13.986 9.144 18.36 ; 
      RECT 8.608 13.986 8.712 18.36 ; 
      RECT 8.176 13.986 8.28 18.36 ; 
      RECT 7.744 13.986 7.848 18.36 ; 
      RECT 7.312 13.986 7.416 18.36 ; 
      RECT 6.88 13.986 6.984 18.36 ; 
      RECT 6.448 13.986 6.552 18.36 ; 
      RECT 6.016 13.986 6.12 18.36 ; 
      RECT 5.584 13.986 5.688 18.36 ; 
      RECT 5.152 13.986 5.256 18.36 ; 
      RECT 4.72 13.986 4.824 18.36 ; 
      RECT 4.288 13.986 4.392 18.36 ; 
      RECT 3.856 13.986 3.96 18.36 ; 
      RECT 3.424 13.986 3.528 18.36 ; 
      RECT 2.992 13.986 3.096 18.36 ; 
      RECT 2.56 13.986 2.664 18.36 ; 
      RECT 2.128 13.986 2.232 18.36 ; 
      RECT 1.696 13.986 1.8 18.36 ; 
      RECT 1.264 13.986 1.368 18.36 ; 
      RECT 0.832 13.986 0.936 18.36 ; 
      RECT 0.02 13.986 0.36 18.36 ; 
      RECT 34.564 18.306 35.076 22.68 ; 
      RECT 34.508 20.968 35.076 22.258 ; 
      RECT 33.916 19.876 34.164 22.68 ; 
      RECT 33.86 21.114 34.164 21.728 ; 
      RECT 33.916 18.306 34.02 22.68 ; 
      RECT 33.916 18.79 34.076 19.748 ; 
      RECT 33.916 18.306 34.164 18.662 ; 
      RECT 32.728 20.108 33.552 22.68 ; 
      RECT 33.448 18.306 33.552 22.68 ; 
      RECT 32.728 21.216 33.608 22.248 ; 
      RECT 32.728 18.306 33.12 22.68 ; 
      RECT 31.06 18.306 31.392 22.68 ; 
      RECT 31.06 18.66 31.448 22.402 ; 
      RECT 65.776 18.306 66.116 22.68 ; 
      RECT 65.2 18.306 65.304 22.68 ; 
      RECT 64.768 18.306 64.872 22.68 ; 
      RECT 64.336 18.306 64.44 22.68 ; 
      RECT 63.904 18.306 64.008 22.68 ; 
      RECT 63.472 18.306 63.576 22.68 ; 
      RECT 63.04 18.306 63.144 22.68 ; 
      RECT 62.608 18.306 62.712 22.68 ; 
      RECT 62.176 18.306 62.28 22.68 ; 
      RECT 61.744 18.306 61.848 22.68 ; 
      RECT 61.312 18.306 61.416 22.68 ; 
      RECT 60.88 18.306 60.984 22.68 ; 
      RECT 60.448 18.306 60.552 22.68 ; 
      RECT 60.016 18.306 60.12 22.68 ; 
      RECT 59.584 18.306 59.688 22.68 ; 
      RECT 59.152 18.306 59.256 22.68 ; 
      RECT 58.72 18.306 58.824 22.68 ; 
      RECT 58.288 18.306 58.392 22.68 ; 
      RECT 57.856 18.306 57.96 22.68 ; 
      RECT 57.424 18.306 57.528 22.68 ; 
      RECT 56.992 18.306 57.096 22.68 ; 
      RECT 56.56 18.306 56.664 22.68 ; 
      RECT 56.128 18.306 56.232 22.68 ; 
      RECT 55.696 18.306 55.8 22.68 ; 
      RECT 55.264 18.306 55.368 22.68 ; 
      RECT 54.832 18.306 54.936 22.68 ; 
      RECT 54.4 18.306 54.504 22.68 ; 
      RECT 53.968 18.306 54.072 22.68 ; 
      RECT 53.536 18.306 53.64 22.68 ; 
      RECT 53.104 18.306 53.208 22.68 ; 
      RECT 52.672 18.306 52.776 22.68 ; 
      RECT 52.24 18.306 52.344 22.68 ; 
      RECT 51.808 18.306 51.912 22.68 ; 
      RECT 51.376 18.306 51.48 22.68 ; 
      RECT 50.944 18.306 51.048 22.68 ; 
      RECT 50.512 18.306 50.616 22.68 ; 
      RECT 50.08 18.306 50.184 22.68 ; 
      RECT 49.648 18.306 49.752 22.68 ; 
      RECT 49.216 18.306 49.32 22.68 ; 
      RECT 48.784 18.306 48.888 22.68 ; 
      RECT 48.352 18.306 48.456 22.68 ; 
      RECT 47.92 18.306 48.024 22.68 ; 
      RECT 47.488 18.306 47.592 22.68 ; 
      RECT 47.056 18.306 47.16 22.68 ; 
      RECT 46.624 18.306 46.728 22.68 ; 
      RECT 46.192 18.306 46.296 22.68 ; 
      RECT 45.76 18.306 45.864 22.68 ; 
      RECT 45.328 18.306 45.432 22.68 ; 
      RECT 44.896 18.306 45 22.68 ; 
      RECT 44.464 18.306 44.568 22.68 ; 
      RECT 44.032 18.306 44.136 22.68 ; 
      RECT 43.6 18.306 43.704 22.68 ; 
      RECT 43.168 18.306 43.272 22.68 ; 
      RECT 42.736 18.306 42.84 22.68 ; 
      RECT 42.304 18.306 42.408 22.68 ; 
      RECT 41.872 18.306 41.976 22.68 ; 
      RECT 41.44 18.306 41.544 22.68 ; 
      RECT 41.008 18.306 41.112 22.68 ; 
      RECT 40.576 18.306 40.68 22.68 ; 
      RECT 40.144 18.306 40.248 22.68 ; 
      RECT 39.712 18.306 39.816 22.68 ; 
      RECT 39.28 18.306 39.384 22.68 ; 
      RECT 38.848 18.306 38.952 22.68 ; 
      RECT 38.416 18.306 38.52 22.68 ; 
      RECT 37.984 18.306 38.088 22.68 ; 
      RECT 37.552 18.306 37.656 22.68 ; 
      RECT 36.7 18.306 37.008 22.68 ; 
      RECT 29.128 18.306 29.436 22.68 ; 
      RECT 28.48 18.306 28.584 22.68 ; 
      RECT 28.048 18.306 28.152 22.68 ; 
      RECT 27.616 18.306 27.72 22.68 ; 
      RECT 27.184 18.306 27.288 22.68 ; 
      RECT 26.752 18.306 26.856 22.68 ; 
      RECT 26.32 18.306 26.424 22.68 ; 
      RECT 25.888 18.306 25.992 22.68 ; 
      RECT 25.456 18.306 25.56 22.68 ; 
      RECT 25.024 18.306 25.128 22.68 ; 
      RECT 24.592 18.306 24.696 22.68 ; 
      RECT 24.16 18.306 24.264 22.68 ; 
      RECT 23.728 18.306 23.832 22.68 ; 
      RECT 23.296 18.306 23.4 22.68 ; 
      RECT 22.864 18.306 22.968 22.68 ; 
      RECT 22.432 18.306 22.536 22.68 ; 
      RECT 22 18.306 22.104 22.68 ; 
      RECT 21.568 18.306 21.672 22.68 ; 
      RECT 21.136 18.306 21.24 22.68 ; 
      RECT 20.704 18.306 20.808 22.68 ; 
      RECT 20.272 18.306 20.376 22.68 ; 
      RECT 19.84 18.306 19.944 22.68 ; 
      RECT 19.408 18.306 19.512 22.68 ; 
      RECT 18.976 18.306 19.08 22.68 ; 
      RECT 18.544 18.306 18.648 22.68 ; 
      RECT 18.112 18.306 18.216 22.68 ; 
      RECT 17.68 18.306 17.784 22.68 ; 
      RECT 17.248 18.306 17.352 22.68 ; 
      RECT 16.816 18.306 16.92 22.68 ; 
      RECT 16.384 18.306 16.488 22.68 ; 
      RECT 15.952 18.306 16.056 22.68 ; 
      RECT 15.52 18.306 15.624 22.68 ; 
      RECT 15.088 18.306 15.192 22.68 ; 
      RECT 14.656 18.306 14.76 22.68 ; 
      RECT 14.224 18.306 14.328 22.68 ; 
      RECT 13.792 18.306 13.896 22.68 ; 
      RECT 13.36 18.306 13.464 22.68 ; 
      RECT 12.928 18.306 13.032 22.68 ; 
      RECT 12.496 18.306 12.6 22.68 ; 
      RECT 12.064 18.306 12.168 22.68 ; 
      RECT 11.632 18.306 11.736 22.68 ; 
      RECT 11.2 18.306 11.304 22.68 ; 
      RECT 10.768 18.306 10.872 22.68 ; 
      RECT 10.336 18.306 10.44 22.68 ; 
      RECT 9.904 18.306 10.008 22.68 ; 
      RECT 9.472 18.306 9.576 22.68 ; 
      RECT 9.04 18.306 9.144 22.68 ; 
      RECT 8.608 18.306 8.712 22.68 ; 
      RECT 8.176 18.306 8.28 22.68 ; 
      RECT 7.744 18.306 7.848 22.68 ; 
      RECT 7.312 18.306 7.416 22.68 ; 
      RECT 6.88 18.306 6.984 22.68 ; 
      RECT 6.448 18.306 6.552 22.68 ; 
      RECT 6.016 18.306 6.12 22.68 ; 
      RECT 5.584 18.306 5.688 22.68 ; 
      RECT 5.152 18.306 5.256 22.68 ; 
      RECT 4.72 18.306 4.824 22.68 ; 
      RECT 4.288 18.306 4.392 22.68 ; 
      RECT 3.856 18.306 3.96 22.68 ; 
      RECT 3.424 18.306 3.528 22.68 ; 
      RECT 2.992 18.306 3.096 22.68 ; 
      RECT 2.56 18.306 2.664 22.68 ; 
      RECT 2.128 18.306 2.232 22.68 ; 
      RECT 1.696 18.306 1.8 22.68 ; 
      RECT 1.264 18.306 1.368 22.68 ; 
      RECT 0.832 18.306 0.936 22.68 ; 
      RECT 0.02 18.306 0.36 22.68 ; 
      RECT 34.564 22.626 35.076 27 ; 
      RECT 34.508 25.288 35.076 26.578 ; 
      RECT 33.916 24.196 34.164 27 ; 
      RECT 33.86 25.434 34.164 26.048 ; 
      RECT 33.916 22.626 34.02 27 ; 
      RECT 33.916 23.11 34.076 24.068 ; 
      RECT 33.916 22.626 34.164 22.982 ; 
      RECT 32.728 24.428 33.552 27 ; 
      RECT 33.448 22.626 33.552 27 ; 
      RECT 32.728 25.536 33.608 26.568 ; 
      RECT 32.728 22.626 33.12 27 ; 
      RECT 31.06 22.626 31.392 27 ; 
      RECT 31.06 22.98 31.448 26.722 ; 
      RECT 65.776 22.626 66.116 27 ; 
      RECT 65.2 22.626 65.304 27 ; 
      RECT 64.768 22.626 64.872 27 ; 
      RECT 64.336 22.626 64.44 27 ; 
      RECT 63.904 22.626 64.008 27 ; 
      RECT 63.472 22.626 63.576 27 ; 
      RECT 63.04 22.626 63.144 27 ; 
      RECT 62.608 22.626 62.712 27 ; 
      RECT 62.176 22.626 62.28 27 ; 
      RECT 61.744 22.626 61.848 27 ; 
      RECT 61.312 22.626 61.416 27 ; 
      RECT 60.88 22.626 60.984 27 ; 
      RECT 60.448 22.626 60.552 27 ; 
      RECT 60.016 22.626 60.12 27 ; 
      RECT 59.584 22.626 59.688 27 ; 
      RECT 59.152 22.626 59.256 27 ; 
      RECT 58.72 22.626 58.824 27 ; 
      RECT 58.288 22.626 58.392 27 ; 
      RECT 57.856 22.626 57.96 27 ; 
      RECT 57.424 22.626 57.528 27 ; 
      RECT 56.992 22.626 57.096 27 ; 
      RECT 56.56 22.626 56.664 27 ; 
      RECT 56.128 22.626 56.232 27 ; 
      RECT 55.696 22.626 55.8 27 ; 
      RECT 55.264 22.626 55.368 27 ; 
      RECT 54.832 22.626 54.936 27 ; 
      RECT 54.4 22.626 54.504 27 ; 
      RECT 53.968 22.626 54.072 27 ; 
      RECT 53.536 22.626 53.64 27 ; 
      RECT 53.104 22.626 53.208 27 ; 
      RECT 52.672 22.626 52.776 27 ; 
      RECT 52.24 22.626 52.344 27 ; 
      RECT 51.808 22.626 51.912 27 ; 
      RECT 51.376 22.626 51.48 27 ; 
      RECT 50.944 22.626 51.048 27 ; 
      RECT 50.512 22.626 50.616 27 ; 
      RECT 50.08 22.626 50.184 27 ; 
      RECT 49.648 22.626 49.752 27 ; 
      RECT 49.216 22.626 49.32 27 ; 
      RECT 48.784 22.626 48.888 27 ; 
      RECT 48.352 22.626 48.456 27 ; 
      RECT 47.92 22.626 48.024 27 ; 
      RECT 47.488 22.626 47.592 27 ; 
      RECT 47.056 22.626 47.16 27 ; 
      RECT 46.624 22.626 46.728 27 ; 
      RECT 46.192 22.626 46.296 27 ; 
      RECT 45.76 22.626 45.864 27 ; 
      RECT 45.328 22.626 45.432 27 ; 
      RECT 44.896 22.626 45 27 ; 
      RECT 44.464 22.626 44.568 27 ; 
      RECT 44.032 22.626 44.136 27 ; 
      RECT 43.6 22.626 43.704 27 ; 
      RECT 43.168 22.626 43.272 27 ; 
      RECT 42.736 22.626 42.84 27 ; 
      RECT 42.304 22.626 42.408 27 ; 
      RECT 41.872 22.626 41.976 27 ; 
      RECT 41.44 22.626 41.544 27 ; 
      RECT 41.008 22.626 41.112 27 ; 
      RECT 40.576 22.626 40.68 27 ; 
      RECT 40.144 22.626 40.248 27 ; 
      RECT 39.712 22.626 39.816 27 ; 
      RECT 39.28 22.626 39.384 27 ; 
      RECT 38.848 22.626 38.952 27 ; 
      RECT 38.416 22.626 38.52 27 ; 
      RECT 37.984 22.626 38.088 27 ; 
      RECT 37.552 22.626 37.656 27 ; 
      RECT 36.7 22.626 37.008 27 ; 
      RECT 29.128 22.626 29.436 27 ; 
      RECT 28.48 22.626 28.584 27 ; 
      RECT 28.048 22.626 28.152 27 ; 
      RECT 27.616 22.626 27.72 27 ; 
      RECT 27.184 22.626 27.288 27 ; 
      RECT 26.752 22.626 26.856 27 ; 
      RECT 26.32 22.626 26.424 27 ; 
      RECT 25.888 22.626 25.992 27 ; 
      RECT 25.456 22.626 25.56 27 ; 
      RECT 25.024 22.626 25.128 27 ; 
      RECT 24.592 22.626 24.696 27 ; 
      RECT 24.16 22.626 24.264 27 ; 
      RECT 23.728 22.626 23.832 27 ; 
      RECT 23.296 22.626 23.4 27 ; 
      RECT 22.864 22.626 22.968 27 ; 
      RECT 22.432 22.626 22.536 27 ; 
      RECT 22 22.626 22.104 27 ; 
      RECT 21.568 22.626 21.672 27 ; 
      RECT 21.136 22.626 21.24 27 ; 
      RECT 20.704 22.626 20.808 27 ; 
      RECT 20.272 22.626 20.376 27 ; 
      RECT 19.84 22.626 19.944 27 ; 
      RECT 19.408 22.626 19.512 27 ; 
      RECT 18.976 22.626 19.08 27 ; 
      RECT 18.544 22.626 18.648 27 ; 
      RECT 18.112 22.626 18.216 27 ; 
      RECT 17.68 22.626 17.784 27 ; 
      RECT 17.248 22.626 17.352 27 ; 
      RECT 16.816 22.626 16.92 27 ; 
      RECT 16.384 22.626 16.488 27 ; 
      RECT 15.952 22.626 16.056 27 ; 
      RECT 15.52 22.626 15.624 27 ; 
      RECT 15.088 22.626 15.192 27 ; 
      RECT 14.656 22.626 14.76 27 ; 
      RECT 14.224 22.626 14.328 27 ; 
      RECT 13.792 22.626 13.896 27 ; 
      RECT 13.36 22.626 13.464 27 ; 
      RECT 12.928 22.626 13.032 27 ; 
      RECT 12.496 22.626 12.6 27 ; 
      RECT 12.064 22.626 12.168 27 ; 
      RECT 11.632 22.626 11.736 27 ; 
      RECT 11.2 22.626 11.304 27 ; 
      RECT 10.768 22.626 10.872 27 ; 
      RECT 10.336 22.626 10.44 27 ; 
      RECT 9.904 22.626 10.008 27 ; 
      RECT 9.472 22.626 9.576 27 ; 
      RECT 9.04 22.626 9.144 27 ; 
      RECT 8.608 22.626 8.712 27 ; 
      RECT 8.176 22.626 8.28 27 ; 
      RECT 7.744 22.626 7.848 27 ; 
      RECT 7.312 22.626 7.416 27 ; 
      RECT 6.88 22.626 6.984 27 ; 
      RECT 6.448 22.626 6.552 27 ; 
      RECT 6.016 22.626 6.12 27 ; 
      RECT 5.584 22.626 5.688 27 ; 
      RECT 5.152 22.626 5.256 27 ; 
      RECT 4.72 22.626 4.824 27 ; 
      RECT 4.288 22.626 4.392 27 ; 
      RECT 3.856 22.626 3.96 27 ; 
      RECT 3.424 22.626 3.528 27 ; 
      RECT 2.992 22.626 3.096 27 ; 
      RECT 2.56 22.626 2.664 27 ; 
      RECT 2.128 22.626 2.232 27 ; 
      RECT 1.696 22.626 1.8 27 ; 
      RECT 1.264 22.626 1.368 27 ; 
      RECT 0.832 22.626 0.936 27 ; 
      RECT 0.02 22.626 0.36 27 ; 
      RECT 34.564 26.946 35.076 31.32 ; 
      RECT 34.508 29.608 35.076 30.898 ; 
      RECT 33.916 28.516 34.164 31.32 ; 
      RECT 33.86 29.754 34.164 30.368 ; 
      RECT 33.916 26.946 34.02 31.32 ; 
      RECT 33.916 27.43 34.076 28.388 ; 
      RECT 33.916 26.946 34.164 27.302 ; 
      RECT 32.728 28.748 33.552 31.32 ; 
      RECT 33.448 26.946 33.552 31.32 ; 
      RECT 32.728 29.856 33.608 30.888 ; 
      RECT 32.728 26.946 33.12 31.32 ; 
      RECT 31.06 26.946 31.392 31.32 ; 
      RECT 31.06 27.3 31.448 31.042 ; 
      RECT 65.776 26.946 66.116 31.32 ; 
      RECT 65.2 26.946 65.304 31.32 ; 
      RECT 64.768 26.946 64.872 31.32 ; 
      RECT 64.336 26.946 64.44 31.32 ; 
      RECT 63.904 26.946 64.008 31.32 ; 
      RECT 63.472 26.946 63.576 31.32 ; 
      RECT 63.04 26.946 63.144 31.32 ; 
      RECT 62.608 26.946 62.712 31.32 ; 
      RECT 62.176 26.946 62.28 31.32 ; 
      RECT 61.744 26.946 61.848 31.32 ; 
      RECT 61.312 26.946 61.416 31.32 ; 
      RECT 60.88 26.946 60.984 31.32 ; 
      RECT 60.448 26.946 60.552 31.32 ; 
      RECT 60.016 26.946 60.12 31.32 ; 
      RECT 59.584 26.946 59.688 31.32 ; 
      RECT 59.152 26.946 59.256 31.32 ; 
      RECT 58.72 26.946 58.824 31.32 ; 
      RECT 58.288 26.946 58.392 31.32 ; 
      RECT 57.856 26.946 57.96 31.32 ; 
      RECT 57.424 26.946 57.528 31.32 ; 
      RECT 56.992 26.946 57.096 31.32 ; 
      RECT 56.56 26.946 56.664 31.32 ; 
      RECT 56.128 26.946 56.232 31.32 ; 
      RECT 55.696 26.946 55.8 31.32 ; 
      RECT 55.264 26.946 55.368 31.32 ; 
      RECT 54.832 26.946 54.936 31.32 ; 
      RECT 54.4 26.946 54.504 31.32 ; 
      RECT 53.968 26.946 54.072 31.32 ; 
      RECT 53.536 26.946 53.64 31.32 ; 
      RECT 53.104 26.946 53.208 31.32 ; 
      RECT 52.672 26.946 52.776 31.32 ; 
      RECT 52.24 26.946 52.344 31.32 ; 
      RECT 51.808 26.946 51.912 31.32 ; 
      RECT 51.376 26.946 51.48 31.32 ; 
      RECT 50.944 26.946 51.048 31.32 ; 
      RECT 50.512 26.946 50.616 31.32 ; 
      RECT 50.08 26.946 50.184 31.32 ; 
      RECT 49.648 26.946 49.752 31.32 ; 
      RECT 49.216 26.946 49.32 31.32 ; 
      RECT 48.784 26.946 48.888 31.32 ; 
      RECT 48.352 26.946 48.456 31.32 ; 
      RECT 47.92 26.946 48.024 31.32 ; 
      RECT 47.488 26.946 47.592 31.32 ; 
      RECT 47.056 26.946 47.16 31.32 ; 
      RECT 46.624 26.946 46.728 31.32 ; 
      RECT 46.192 26.946 46.296 31.32 ; 
      RECT 45.76 26.946 45.864 31.32 ; 
      RECT 45.328 26.946 45.432 31.32 ; 
      RECT 44.896 26.946 45 31.32 ; 
      RECT 44.464 26.946 44.568 31.32 ; 
      RECT 44.032 26.946 44.136 31.32 ; 
      RECT 43.6 26.946 43.704 31.32 ; 
      RECT 43.168 26.946 43.272 31.32 ; 
      RECT 42.736 26.946 42.84 31.32 ; 
      RECT 42.304 26.946 42.408 31.32 ; 
      RECT 41.872 26.946 41.976 31.32 ; 
      RECT 41.44 26.946 41.544 31.32 ; 
      RECT 41.008 26.946 41.112 31.32 ; 
      RECT 40.576 26.946 40.68 31.32 ; 
      RECT 40.144 26.946 40.248 31.32 ; 
      RECT 39.712 26.946 39.816 31.32 ; 
      RECT 39.28 26.946 39.384 31.32 ; 
      RECT 38.848 26.946 38.952 31.32 ; 
      RECT 38.416 26.946 38.52 31.32 ; 
      RECT 37.984 26.946 38.088 31.32 ; 
      RECT 37.552 26.946 37.656 31.32 ; 
      RECT 36.7 26.946 37.008 31.32 ; 
      RECT 29.128 26.946 29.436 31.32 ; 
      RECT 28.48 26.946 28.584 31.32 ; 
      RECT 28.048 26.946 28.152 31.32 ; 
      RECT 27.616 26.946 27.72 31.32 ; 
      RECT 27.184 26.946 27.288 31.32 ; 
      RECT 26.752 26.946 26.856 31.32 ; 
      RECT 26.32 26.946 26.424 31.32 ; 
      RECT 25.888 26.946 25.992 31.32 ; 
      RECT 25.456 26.946 25.56 31.32 ; 
      RECT 25.024 26.946 25.128 31.32 ; 
      RECT 24.592 26.946 24.696 31.32 ; 
      RECT 24.16 26.946 24.264 31.32 ; 
      RECT 23.728 26.946 23.832 31.32 ; 
      RECT 23.296 26.946 23.4 31.32 ; 
      RECT 22.864 26.946 22.968 31.32 ; 
      RECT 22.432 26.946 22.536 31.32 ; 
      RECT 22 26.946 22.104 31.32 ; 
      RECT 21.568 26.946 21.672 31.32 ; 
      RECT 21.136 26.946 21.24 31.32 ; 
      RECT 20.704 26.946 20.808 31.32 ; 
      RECT 20.272 26.946 20.376 31.32 ; 
      RECT 19.84 26.946 19.944 31.32 ; 
      RECT 19.408 26.946 19.512 31.32 ; 
      RECT 18.976 26.946 19.08 31.32 ; 
      RECT 18.544 26.946 18.648 31.32 ; 
      RECT 18.112 26.946 18.216 31.32 ; 
      RECT 17.68 26.946 17.784 31.32 ; 
      RECT 17.248 26.946 17.352 31.32 ; 
      RECT 16.816 26.946 16.92 31.32 ; 
      RECT 16.384 26.946 16.488 31.32 ; 
      RECT 15.952 26.946 16.056 31.32 ; 
      RECT 15.52 26.946 15.624 31.32 ; 
      RECT 15.088 26.946 15.192 31.32 ; 
      RECT 14.656 26.946 14.76 31.32 ; 
      RECT 14.224 26.946 14.328 31.32 ; 
      RECT 13.792 26.946 13.896 31.32 ; 
      RECT 13.36 26.946 13.464 31.32 ; 
      RECT 12.928 26.946 13.032 31.32 ; 
      RECT 12.496 26.946 12.6 31.32 ; 
      RECT 12.064 26.946 12.168 31.32 ; 
      RECT 11.632 26.946 11.736 31.32 ; 
      RECT 11.2 26.946 11.304 31.32 ; 
      RECT 10.768 26.946 10.872 31.32 ; 
      RECT 10.336 26.946 10.44 31.32 ; 
      RECT 9.904 26.946 10.008 31.32 ; 
      RECT 9.472 26.946 9.576 31.32 ; 
      RECT 9.04 26.946 9.144 31.32 ; 
      RECT 8.608 26.946 8.712 31.32 ; 
      RECT 8.176 26.946 8.28 31.32 ; 
      RECT 7.744 26.946 7.848 31.32 ; 
      RECT 7.312 26.946 7.416 31.32 ; 
      RECT 6.88 26.946 6.984 31.32 ; 
      RECT 6.448 26.946 6.552 31.32 ; 
      RECT 6.016 26.946 6.12 31.32 ; 
      RECT 5.584 26.946 5.688 31.32 ; 
      RECT 5.152 26.946 5.256 31.32 ; 
      RECT 4.72 26.946 4.824 31.32 ; 
      RECT 4.288 26.946 4.392 31.32 ; 
      RECT 3.856 26.946 3.96 31.32 ; 
      RECT 3.424 26.946 3.528 31.32 ; 
      RECT 2.992 26.946 3.096 31.32 ; 
      RECT 2.56 26.946 2.664 31.32 ; 
      RECT 2.128 26.946 2.232 31.32 ; 
      RECT 1.696 26.946 1.8 31.32 ; 
      RECT 1.264 26.946 1.368 31.32 ; 
      RECT 0.832 26.946 0.936 31.32 ; 
      RECT 0.02 26.946 0.36 31.32 ; 
      RECT 34.564 31.266 35.076 35.64 ; 
      RECT 34.508 33.928 35.076 35.218 ; 
      RECT 33.916 32.836 34.164 35.64 ; 
      RECT 33.86 34.074 34.164 34.688 ; 
      RECT 33.916 31.266 34.02 35.64 ; 
      RECT 33.916 31.75 34.076 32.708 ; 
      RECT 33.916 31.266 34.164 31.622 ; 
      RECT 32.728 33.068 33.552 35.64 ; 
      RECT 33.448 31.266 33.552 35.64 ; 
      RECT 32.728 34.176 33.608 35.208 ; 
      RECT 32.728 31.266 33.12 35.64 ; 
      RECT 31.06 31.266 31.392 35.64 ; 
      RECT 31.06 31.62 31.448 35.362 ; 
      RECT 65.776 31.266 66.116 35.64 ; 
      RECT 65.2 31.266 65.304 35.64 ; 
      RECT 64.768 31.266 64.872 35.64 ; 
      RECT 64.336 31.266 64.44 35.64 ; 
      RECT 63.904 31.266 64.008 35.64 ; 
      RECT 63.472 31.266 63.576 35.64 ; 
      RECT 63.04 31.266 63.144 35.64 ; 
      RECT 62.608 31.266 62.712 35.64 ; 
      RECT 62.176 31.266 62.28 35.64 ; 
      RECT 61.744 31.266 61.848 35.64 ; 
      RECT 61.312 31.266 61.416 35.64 ; 
      RECT 60.88 31.266 60.984 35.64 ; 
      RECT 60.448 31.266 60.552 35.64 ; 
      RECT 60.016 31.266 60.12 35.64 ; 
      RECT 59.584 31.266 59.688 35.64 ; 
      RECT 59.152 31.266 59.256 35.64 ; 
      RECT 58.72 31.266 58.824 35.64 ; 
      RECT 58.288 31.266 58.392 35.64 ; 
      RECT 57.856 31.266 57.96 35.64 ; 
      RECT 57.424 31.266 57.528 35.64 ; 
      RECT 56.992 31.266 57.096 35.64 ; 
      RECT 56.56 31.266 56.664 35.64 ; 
      RECT 56.128 31.266 56.232 35.64 ; 
      RECT 55.696 31.266 55.8 35.64 ; 
      RECT 55.264 31.266 55.368 35.64 ; 
      RECT 54.832 31.266 54.936 35.64 ; 
      RECT 54.4 31.266 54.504 35.64 ; 
      RECT 53.968 31.266 54.072 35.64 ; 
      RECT 53.536 31.266 53.64 35.64 ; 
      RECT 53.104 31.266 53.208 35.64 ; 
      RECT 52.672 31.266 52.776 35.64 ; 
      RECT 52.24 31.266 52.344 35.64 ; 
      RECT 51.808 31.266 51.912 35.64 ; 
      RECT 51.376 31.266 51.48 35.64 ; 
      RECT 50.944 31.266 51.048 35.64 ; 
      RECT 50.512 31.266 50.616 35.64 ; 
      RECT 50.08 31.266 50.184 35.64 ; 
      RECT 49.648 31.266 49.752 35.64 ; 
      RECT 49.216 31.266 49.32 35.64 ; 
      RECT 48.784 31.266 48.888 35.64 ; 
      RECT 48.352 31.266 48.456 35.64 ; 
      RECT 47.92 31.266 48.024 35.64 ; 
      RECT 47.488 31.266 47.592 35.64 ; 
      RECT 47.056 31.266 47.16 35.64 ; 
      RECT 46.624 31.266 46.728 35.64 ; 
      RECT 46.192 31.266 46.296 35.64 ; 
      RECT 45.76 31.266 45.864 35.64 ; 
      RECT 45.328 31.266 45.432 35.64 ; 
      RECT 44.896 31.266 45 35.64 ; 
      RECT 44.464 31.266 44.568 35.64 ; 
      RECT 44.032 31.266 44.136 35.64 ; 
      RECT 43.6 31.266 43.704 35.64 ; 
      RECT 43.168 31.266 43.272 35.64 ; 
      RECT 42.736 31.266 42.84 35.64 ; 
      RECT 42.304 31.266 42.408 35.64 ; 
      RECT 41.872 31.266 41.976 35.64 ; 
      RECT 41.44 31.266 41.544 35.64 ; 
      RECT 41.008 31.266 41.112 35.64 ; 
      RECT 40.576 31.266 40.68 35.64 ; 
      RECT 40.144 31.266 40.248 35.64 ; 
      RECT 39.712 31.266 39.816 35.64 ; 
      RECT 39.28 31.266 39.384 35.64 ; 
      RECT 38.848 31.266 38.952 35.64 ; 
      RECT 38.416 31.266 38.52 35.64 ; 
      RECT 37.984 31.266 38.088 35.64 ; 
      RECT 37.552 31.266 37.656 35.64 ; 
      RECT 36.7 31.266 37.008 35.64 ; 
      RECT 29.128 31.266 29.436 35.64 ; 
      RECT 28.48 31.266 28.584 35.64 ; 
      RECT 28.048 31.266 28.152 35.64 ; 
      RECT 27.616 31.266 27.72 35.64 ; 
      RECT 27.184 31.266 27.288 35.64 ; 
      RECT 26.752 31.266 26.856 35.64 ; 
      RECT 26.32 31.266 26.424 35.64 ; 
      RECT 25.888 31.266 25.992 35.64 ; 
      RECT 25.456 31.266 25.56 35.64 ; 
      RECT 25.024 31.266 25.128 35.64 ; 
      RECT 24.592 31.266 24.696 35.64 ; 
      RECT 24.16 31.266 24.264 35.64 ; 
      RECT 23.728 31.266 23.832 35.64 ; 
      RECT 23.296 31.266 23.4 35.64 ; 
      RECT 22.864 31.266 22.968 35.64 ; 
      RECT 22.432 31.266 22.536 35.64 ; 
      RECT 22 31.266 22.104 35.64 ; 
      RECT 21.568 31.266 21.672 35.64 ; 
      RECT 21.136 31.266 21.24 35.64 ; 
      RECT 20.704 31.266 20.808 35.64 ; 
      RECT 20.272 31.266 20.376 35.64 ; 
      RECT 19.84 31.266 19.944 35.64 ; 
      RECT 19.408 31.266 19.512 35.64 ; 
      RECT 18.976 31.266 19.08 35.64 ; 
      RECT 18.544 31.266 18.648 35.64 ; 
      RECT 18.112 31.266 18.216 35.64 ; 
      RECT 17.68 31.266 17.784 35.64 ; 
      RECT 17.248 31.266 17.352 35.64 ; 
      RECT 16.816 31.266 16.92 35.64 ; 
      RECT 16.384 31.266 16.488 35.64 ; 
      RECT 15.952 31.266 16.056 35.64 ; 
      RECT 15.52 31.266 15.624 35.64 ; 
      RECT 15.088 31.266 15.192 35.64 ; 
      RECT 14.656 31.266 14.76 35.64 ; 
      RECT 14.224 31.266 14.328 35.64 ; 
      RECT 13.792 31.266 13.896 35.64 ; 
      RECT 13.36 31.266 13.464 35.64 ; 
      RECT 12.928 31.266 13.032 35.64 ; 
      RECT 12.496 31.266 12.6 35.64 ; 
      RECT 12.064 31.266 12.168 35.64 ; 
      RECT 11.632 31.266 11.736 35.64 ; 
      RECT 11.2 31.266 11.304 35.64 ; 
      RECT 10.768 31.266 10.872 35.64 ; 
      RECT 10.336 31.266 10.44 35.64 ; 
      RECT 9.904 31.266 10.008 35.64 ; 
      RECT 9.472 31.266 9.576 35.64 ; 
      RECT 9.04 31.266 9.144 35.64 ; 
      RECT 8.608 31.266 8.712 35.64 ; 
      RECT 8.176 31.266 8.28 35.64 ; 
      RECT 7.744 31.266 7.848 35.64 ; 
      RECT 7.312 31.266 7.416 35.64 ; 
      RECT 6.88 31.266 6.984 35.64 ; 
      RECT 6.448 31.266 6.552 35.64 ; 
      RECT 6.016 31.266 6.12 35.64 ; 
      RECT 5.584 31.266 5.688 35.64 ; 
      RECT 5.152 31.266 5.256 35.64 ; 
      RECT 4.72 31.266 4.824 35.64 ; 
      RECT 4.288 31.266 4.392 35.64 ; 
      RECT 3.856 31.266 3.96 35.64 ; 
      RECT 3.424 31.266 3.528 35.64 ; 
      RECT 2.992 31.266 3.096 35.64 ; 
      RECT 2.56 31.266 2.664 35.64 ; 
      RECT 2.128 31.266 2.232 35.64 ; 
      RECT 1.696 31.266 1.8 35.64 ; 
      RECT 1.264 31.266 1.368 35.64 ; 
      RECT 0.832 31.266 0.936 35.64 ; 
      RECT 0.02 31.266 0.36 35.64 ; 
      RECT 34.564 35.586 35.076 39.96 ; 
      RECT 34.508 38.248 35.076 39.538 ; 
      RECT 33.916 37.156 34.164 39.96 ; 
      RECT 33.86 38.394 34.164 39.008 ; 
      RECT 33.916 35.586 34.02 39.96 ; 
      RECT 33.916 36.07 34.076 37.028 ; 
      RECT 33.916 35.586 34.164 35.942 ; 
      RECT 32.728 37.388 33.552 39.96 ; 
      RECT 33.448 35.586 33.552 39.96 ; 
      RECT 32.728 38.496 33.608 39.528 ; 
      RECT 32.728 35.586 33.12 39.96 ; 
      RECT 31.06 35.586 31.392 39.96 ; 
      RECT 31.06 35.94 31.448 39.682 ; 
      RECT 65.776 35.586 66.116 39.96 ; 
      RECT 65.2 35.586 65.304 39.96 ; 
      RECT 64.768 35.586 64.872 39.96 ; 
      RECT 64.336 35.586 64.44 39.96 ; 
      RECT 63.904 35.586 64.008 39.96 ; 
      RECT 63.472 35.586 63.576 39.96 ; 
      RECT 63.04 35.586 63.144 39.96 ; 
      RECT 62.608 35.586 62.712 39.96 ; 
      RECT 62.176 35.586 62.28 39.96 ; 
      RECT 61.744 35.586 61.848 39.96 ; 
      RECT 61.312 35.586 61.416 39.96 ; 
      RECT 60.88 35.586 60.984 39.96 ; 
      RECT 60.448 35.586 60.552 39.96 ; 
      RECT 60.016 35.586 60.12 39.96 ; 
      RECT 59.584 35.586 59.688 39.96 ; 
      RECT 59.152 35.586 59.256 39.96 ; 
      RECT 58.72 35.586 58.824 39.96 ; 
      RECT 58.288 35.586 58.392 39.96 ; 
      RECT 57.856 35.586 57.96 39.96 ; 
      RECT 57.424 35.586 57.528 39.96 ; 
      RECT 56.992 35.586 57.096 39.96 ; 
      RECT 56.56 35.586 56.664 39.96 ; 
      RECT 56.128 35.586 56.232 39.96 ; 
      RECT 55.696 35.586 55.8 39.96 ; 
      RECT 55.264 35.586 55.368 39.96 ; 
      RECT 54.832 35.586 54.936 39.96 ; 
      RECT 54.4 35.586 54.504 39.96 ; 
      RECT 53.968 35.586 54.072 39.96 ; 
      RECT 53.536 35.586 53.64 39.96 ; 
      RECT 53.104 35.586 53.208 39.96 ; 
      RECT 52.672 35.586 52.776 39.96 ; 
      RECT 52.24 35.586 52.344 39.96 ; 
      RECT 51.808 35.586 51.912 39.96 ; 
      RECT 51.376 35.586 51.48 39.96 ; 
      RECT 50.944 35.586 51.048 39.96 ; 
      RECT 50.512 35.586 50.616 39.96 ; 
      RECT 50.08 35.586 50.184 39.96 ; 
      RECT 49.648 35.586 49.752 39.96 ; 
      RECT 49.216 35.586 49.32 39.96 ; 
      RECT 48.784 35.586 48.888 39.96 ; 
      RECT 48.352 35.586 48.456 39.96 ; 
      RECT 47.92 35.586 48.024 39.96 ; 
      RECT 47.488 35.586 47.592 39.96 ; 
      RECT 47.056 35.586 47.16 39.96 ; 
      RECT 46.624 35.586 46.728 39.96 ; 
      RECT 46.192 35.586 46.296 39.96 ; 
      RECT 45.76 35.586 45.864 39.96 ; 
      RECT 45.328 35.586 45.432 39.96 ; 
      RECT 44.896 35.586 45 39.96 ; 
      RECT 44.464 35.586 44.568 39.96 ; 
      RECT 44.032 35.586 44.136 39.96 ; 
      RECT 43.6 35.586 43.704 39.96 ; 
      RECT 43.168 35.586 43.272 39.96 ; 
      RECT 42.736 35.586 42.84 39.96 ; 
      RECT 42.304 35.586 42.408 39.96 ; 
      RECT 41.872 35.586 41.976 39.96 ; 
      RECT 41.44 35.586 41.544 39.96 ; 
      RECT 41.008 35.586 41.112 39.96 ; 
      RECT 40.576 35.586 40.68 39.96 ; 
      RECT 40.144 35.586 40.248 39.96 ; 
      RECT 39.712 35.586 39.816 39.96 ; 
      RECT 39.28 35.586 39.384 39.96 ; 
      RECT 38.848 35.586 38.952 39.96 ; 
      RECT 38.416 35.586 38.52 39.96 ; 
      RECT 37.984 35.586 38.088 39.96 ; 
      RECT 37.552 35.586 37.656 39.96 ; 
      RECT 36.7 35.586 37.008 39.96 ; 
      RECT 29.128 35.586 29.436 39.96 ; 
      RECT 28.48 35.586 28.584 39.96 ; 
      RECT 28.048 35.586 28.152 39.96 ; 
      RECT 27.616 35.586 27.72 39.96 ; 
      RECT 27.184 35.586 27.288 39.96 ; 
      RECT 26.752 35.586 26.856 39.96 ; 
      RECT 26.32 35.586 26.424 39.96 ; 
      RECT 25.888 35.586 25.992 39.96 ; 
      RECT 25.456 35.586 25.56 39.96 ; 
      RECT 25.024 35.586 25.128 39.96 ; 
      RECT 24.592 35.586 24.696 39.96 ; 
      RECT 24.16 35.586 24.264 39.96 ; 
      RECT 23.728 35.586 23.832 39.96 ; 
      RECT 23.296 35.586 23.4 39.96 ; 
      RECT 22.864 35.586 22.968 39.96 ; 
      RECT 22.432 35.586 22.536 39.96 ; 
      RECT 22 35.586 22.104 39.96 ; 
      RECT 21.568 35.586 21.672 39.96 ; 
      RECT 21.136 35.586 21.24 39.96 ; 
      RECT 20.704 35.586 20.808 39.96 ; 
      RECT 20.272 35.586 20.376 39.96 ; 
      RECT 19.84 35.586 19.944 39.96 ; 
      RECT 19.408 35.586 19.512 39.96 ; 
      RECT 18.976 35.586 19.08 39.96 ; 
      RECT 18.544 35.586 18.648 39.96 ; 
      RECT 18.112 35.586 18.216 39.96 ; 
      RECT 17.68 35.586 17.784 39.96 ; 
      RECT 17.248 35.586 17.352 39.96 ; 
      RECT 16.816 35.586 16.92 39.96 ; 
      RECT 16.384 35.586 16.488 39.96 ; 
      RECT 15.952 35.586 16.056 39.96 ; 
      RECT 15.52 35.586 15.624 39.96 ; 
      RECT 15.088 35.586 15.192 39.96 ; 
      RECT 14.656 35.586 14.76 39.96 ; 
      RECT 14.224 35.586 14.328 39.96 ; 
      RECT 13.792 35.586 13.896 39.96 ; 
      RECT 13.36 35.586 13.464 39.96 ; 
      RECT 12.928 35.586 13.032 39.96 ; 
      RECT 12.496 35.586 12.6 39.96 ; 
      RECT 12.064 35.586 12.168 39.96 ; 
      RECT 11.632 35.586 11.736 39.96 ; 
      RECT 11.2 35.586 11.304 39.96 ; 
      RECT 10.768 35.586 10.872 39.96 ; 
      RECT 10.336 35.586 10.44 39.96 ; 
      RECT 9.904 35.586 10.008 39.96 ; 
      RECT 9.472 35.586 9.576 39.96 ; 
      RECT 9.04 35.586 9.144 39.96 ; 
      RECT 8.608 35.586 8.712 39.96 ; 
      RECT 8.176 35.586 8.28 39.96 ; 
      RECT 7.744 35.586 7.848 39.96 ; 
      RECT 7.312 35.586 7.416 39.96 ; 
      RECT 6.88 35.586 6.984 39.96 ; 
      RECT 6.448 35.586 6.552 39.96 ; 
      RECT 6.016 35.586 6.12 39.96 ; 
      RECT 5.584 35.586 5.688 39.96 ; 
      RECT 5.152 35.586 5.256 39.96 ; 
      RECT 4.72 35.586 4.824 39.96 ; 
      RECT 4.288 35.586 4.392 39.96 ; 
      RECT 3.856 35.586 3.96 39.96 ; 
      RECT 3.424 35.586 3.528 39.96 ; 
      RECT 2.992 35.586 3.096 39.96 ; 
      RECT 2.56 35.586 2.664 39.96 ; 
      RECT 2.128 35.586 2.232 39.96 ; 
      RECT 1.696 35.586 1.8 39.96 ; 
      RECT 1.264 35.586 1.368 39.96 ; 
      RECT 0.832 35.586 0.936 39.96 ; 
      RECT 0.02 35.586 0.36 39.96 ; 
      RECT 34.564 39.906 35.076 44.28 ; 
      RECT 34.508 42.568 35.076 43.858 ; 
      RECT 33.916 41.476 34.164 44.28 ; 
      RECT 33.86 42.714 34.164 43.328 ; 
      RECT 33.916 39.906 34.02 44.28 ; 
      RECT 33.916 40.39 34.076 41.348 ; 
      RECT 33.916 39.906 34.164 40.262 ; 
      RECT 32.728 41.708 33.552 44.28 ; 
      RECT 33.448 39.906 33.552 44.28 ; 
      RECT 32.728 42.816 33.608 43.848 ; 
      RECT 32.728 39.906 33.12 44.28 ; 
      RECT 31.06 39.906 31.392 44.28 ; 
      RECT 31.06 40.26 31.448 44.002 ; 
      RECT 65.776 39.906 66.116 44.28 ; 
      RECT 65.2 39.906 65.304 44.28 ; 
      RECT 64.768 39.906 64.872 44.28 ; 
      RECT 64.336 39.906 64.44 44.28 ; 
      RECT 63.904 39.906 64.008 44.28 ; 
      RECT 63.472 39.906 63.576 44.28 ; 
      RECT 63.04 39.906 63.144 44.28 ; 
      RECT 62.608 39.906 62.712 44.28 ; 
      RECT 62.176 39.906 62.28 44.28 ; 
      RECT 61.744 39.906 61.848 44.28 ; 
      RECT 61.312 39.906 61.416 44.28 ; 
      RECT 60.88 39.906 60.984 44.28 ; 
      RECT 60.448 39.906 60.552 44.28 ; 
      RECT 60.016 39.906 60.12 44.28 ; 
      RECT 59.584 39.906 59.688 44.28 ; 
      RECT 59.152 39.906 59.256 44.28 ; 
      RECT 58.72 39.906 58.824 44.28 ; 
      RECT 58.288 39.906 58.392 44.28 ; 
      RECT 57.856 39.906 57.96 44.28 ; 
      RECT 57.424 39.906 57.528 44.28 ; 
      RECT 56.992 39.906 57.096 44.28 ; 
      RECT 56.56 39.906 56.664 44.28 ; 
      RECT 56.128 39.906 56.232 44.28 ; 
      RECT 55.696 39.906 55.8 44.28 ; 
      RECT 55.264 39.906 55.368 44.28 ; 
      RECT 54.832 39.906 54.936 44.28 ; 
      RECT 54.4 39.906 54.504 44.28 ; 
      RECT 53.968 39.906 54.072 44.28 ; 
      RECT 53.536 39.906 53.64 44.28 ; 
      RECT 53.104 39.906 53.208 44.28 ; 
      RECT 52.672 39.906 52.776 44.28 ; 
      RECT 52.24 39.906 52.344 44.28 ; 
      RECT 51.808 39.906 51.912 44.28 ; 
      RECT 51.376 39.906 51.48 44.28 ; 
      RECT 50.944 39.906 51.048 44.28 ; 
      RECT 50.512 39.906 50.616 44.28 ; 
      RECT 50.08 39.906 50.184 44.28 ; 
      RECT 49.648 39.906 49.752 44.28 ; 
      RECT 49.216 39.906 49.32 44.28 ; 
      RECT 48.784 39.906 48.888 44.28 ; 
      RECT 48.352 39.906 48.456 44.28 ; 
      RECT 47.92 39.906 48.024 44.28 ; 
      RECT 47.488 39.906 47.592 44.28 ; 
      RECT 47.056 39.906 47.16 44.28 ; 
      RECT 46.624 39.906 46.728 44.28 ; 
      RECT 46.192 39.906 46.296 44.28 ; 
      RECT 45.76 39.906 45.864 44.28 ; 
      RECT 45.328 39.906 45.432 44.28 ; 
      RECT 44.896 39.906 45 44.28 ; 
      RECT 44.464 39.906 44.568 44.28 ; 
      RECT 44.032 39.906 44.136 44.28 ; 
      RECT 43.6 39.906 43.704 44.28 ; 
      RECT 43.168 39.906 43.272 44.28 ; 
      RECT 42.736 39.906 42.84 44.28 ; 
      RECT 42.304 39.906 42.408 44.28 ; 
      RECT 41.872 39.906 41.976 44.28 ; 
      RECT 41.44 39.906 41.544 44.28 ; 
      RECT 41.008 39.906 41.112 44.28 ; 
      RECT 40.576 39.906 40.68 44.28 ; 
      RECT 40.144 39.906 40.248 44.28 ; 
      RECT 39.712 39.906 39.816 44.28 ; 
      RECT 39.28 39.906 39.384 44.28 ; 
      RECT 38.848 39.906 38.952 44.28 ; 
      RECT 38.416 39.906 38.52 44.28 ; 
      RECT 37.984 39.906 38.088 44.28 ; 
      RECT 37.552 39.906 37.656 44.28 ; 
      RECT 36.7 39.906 37.008 44.28 ; 
      RECT 29.128 39.906 29.436 44.28 ; 
      RECT 28.48 39.906 28.584 44.28 ; 
      RECT 28.048 39.906 28.152 44.28 ; 
      RECT 27.616 39.906 27.72 44.28 ; 
      RECT 27.184 39.906 27.288 44.28 ; 
      RECT 26.752 39.906 26.856 44.28 ; 
      RECT 26.32 39.906 26.424 44.28 ; 
      RECT 25.888 39.906 25.992 44.28 ; 
      RECT 25.456 39.906 25.56 44.28 ; 
      RECT 25.024 39.906 25.128 44.28 ; 
      RECT 24.592 39.906 24.696 44.28 ; 
      RECT 24.16 39.906 24.264 44.28 ; 
      RECT 23.728 39.906 23.832 44.28 ; 
      RECT 23.296 39.906 23.4 44.28 ; 
      RECT 22.864 39.906 22.968 44.28 ; 
      RECT 22.432 39.906 22.536 44.28 ; 
      RECT 22 39.906 22.104 44.28 ; 
      RECT 21.568 39.906 21.672 44.28 ; 
      RECT 21.136 39.906 21.24 44.28 ; 
      RECT 20.704 39.906 20.808 44.28 ; 
      RECT 20.272 39.906 20.376 44.28 ; 
      RECT 19.84 39.906 19.944 44.28 ; 
      RECT 19.408 39.906 19.512 44.28 ; 
      RECT 18.976 39.906 19.08 44.28 ; 
      RECT 18.544 39.906 18.648 44.28 ; 
      RECT 18.112 39.906 18.216 44.28 ; 
      RECT 17.68 39.906 17.784 44.28 ; 
      RECT 17.248 39.906 17.352 44.28 ; 
      RECT 16.816 39.906 16.92 44.28 ; 
      RECT 16.384 39.906 16.488 44.28 ; 
      RECT 15.952 39.906 16.056 44.28 ; 
      RECT 15.52 39.906 15.624 44.28 ; 
      RECT 15.088 39.906 15.192 44.28 ; 
      RECT 14.656 39.906 14.76 44.28 ; 
      RECT 14.224 39.906 14.328 44.28 ; 
      RECT 13.792 39.906 13.896 44.28 ; 
      RECT 13.36 39.906 13.464 44.28 ; 
      RECT 12.928 39.906 13.032 44.28 ; 
      RECT 12.496 39.906 12.6 44.28 ; 
      RECT 12.064 39.906 12.168 44.28 ; 
      RECT 11.632 39.906 11.736 44.28 ; 
      RECT 11.2 39.906 11.304 44.28 ; 
      RECT 10.768 39.906 10.872 44.28 ; 
      RECT 10.336 39.906 10.44 44.28 ; 
      RECT 9.904 39.906 10.008 44.28 ; 
      RECT 9.472 39.906 9.576 44.28 ; 
      RECT 9.04 39.906 9.144 44.28 ; 
      RECT 8.608 39.906 8.712 44.28 ; 
      RECT 8.176 39.906 8.28 44.28 ; 
      RECT 7.744 39.906 7.848 44.28 ; 
      RECT 7.312 39.906 7.416 44.28 ; 
      RECT 6.88 39.906 6.984 44.28 ; 
      RECT 6.448 39.906 6.552 44.28 ; 
      RECT 6.016 39.906 6.12 44.28 ; 
      RECT 5.584 39.906 5.688 44.28 ; 
      RECT 5.152 39.906 5.256 44.28 ; 
      RECT 4.72 39.906 4.824 44.28 ; 
      RECT 4.288 39.906 4.392 44.28 ; 
      RECT 3.856 39.906 3.96 44.28 ; 
      RECT 3.424 39.906 3.528 44.28 ; 
      RECT 2.992 39.906 3.096 44.28 ; 
      RECT 2.56 39.906 2.664 44.28 ; 
      RECT 2.128 39.906 2.232 44.28 ; 
      RECT 1.696 39.906 1.8 44.28 ; 
      RECT 1.264 39.906 1.368 44.28 ; 
      RECT 0.832 39.906 0.936 44.28 ; 
      RECT 0.02 39.906 0.36 44.28 ; 
      RECT 34.564 44.226 35.076 48.6 ; 
      RECT 34.508 46.888 35.076 48.178 ; 
      RECT 33.916 45.796 34.164 48.6 ; 
      RECT 33.86 47.034 34.164 47.648 ; 
      RECT 33.916 44.226 34.02 48.6 ; 
      RECT 33.916 44.71 34.076 45.668 ; 
      RECT 33.916 44.226 34.164 44.582 ; 
      RECT 32.728 46.028 33.552 48.6 ; 
      RECT 33.448 44.226 33.552 48.6 ; 
      RECT 32.728 47.136 33.608 48.168 ; 
      RECT 32.728 44.226 33.12 48.6 ; 
      RECT 31.06 44.226 31.392 48.6 ; 
      RECT 31.06 44.58 31.448 48.322 ; 
      RECT 65.776 44.226 66.116 48.6 ; 
      RECT 65.2 44.226 65.304 48.6 ; 
      RECT 64.768 44.226 64.872 48.6 ; 
      RECT 64.336 44.226 64.44 48.6 ; 
      RECT 63.904 44.226 64.008 48.6 ; 
      RECT 63.472 44.226 63.576 48.6 ; 
      RECT 63.04 44.226 63.144 48.6 ; 
      RECT 62.608 44.226 62.712 48.6 ; 
      RECT 62.176 44.226 62.28 48.6 ; 
      RECT 61.744 44.226 61.848 48.6 ; 
      RECT 61.312 44.226 61.416 48.6 ; 
      RECT 60.88 44.226 60.984 48.6 ; 
      RECT 60.448 44.226 60.552 48.6 ; 
      RECT 60.016 44.226 60.12 48.6 ; 
      RECT 59.584 44.226 59.688 48.6 ; 
      RECT 59.152 44.226 59.256 48.6 ; 
      RECT 58.72 44.226 58.824 48.6 ; 
      RECT 58.288 44.226 58.392 48.6 ; 
      RECT 57.856 44.226 57.96 48.6 ; 
      RECT 57.424 44.226 57.528 48.6 ; 
      RECT 56.992 44.226 57.096 48.6 ; 
      RECT 56.56 44.226 56.664 48.6 ; 
      RECT 56.128 44.226 56.232 48.6 ; 
      RECT 55.696 44.226 55.8 48.6 ; 
      RECT 55.264 44.226 55.368 48.6 ; 
      RECT 54.832 44.226 54.936 48.6 ; 
      RECT 54.4 44.226 54.504 48.6 ; 
      RECT 53.968 44.226 54.072 48.6 ; 
      RECT 53.536 44.226 53.64 48.6 ; 
      RECT 53.104 44.226 53.208 48.6 ; 
      RECT 52.672 44.226 52.776 48.6 ; 
      RECT 52.24 44.226 52.344 48.6 ; 
      RECT 51.808 44.226 51.912 48.6 ; 
      RECT 51.376 44.226 51.48 48.6 ; 
      RECT 50.944 44.226 51.048 48.6 ; 
      RECT 50.512 44.226 50.616 48.6 ; 
      RECT 50.08 44.226 50.184 48.6 ; 
      RECT 49.648 44.226 49.752 48.6 ; 
      RECT 49.216 44.226 49.32 48.6 ; 
      RECT 48.784 44.226 48.888 48.6 ; 
      RECT 48.352 44.226 48.456 48.6 ; 
      RECT 47.92 44.226 48.024 48.6 ; 
      RECT 47.488 44.226 47.592 48.6 ; 
      RECT 47.056 44.226 47.16 48.6 ; 
      RECT 46.624 44.226 46.728 48.6 ; 
      RECT 46.192 44.226 46.296 48.6 ; 
      RECT 45.76 44.226 45.864 48.6 ; 
      RECT 45.328 44.226 45.432 48.6 ; 
      RECT 44.896 44.226 45 48.6 ; 
      RECT 44.464 44.226 44.568 48.6 ; 
      RECT 44.032 44.226 44.136 48.6 ; 
      RECT 43.6 44.226 43.704 48.6 ; 
      RECT 43.168 44.226 43.272 48.6 ; 
      RECT 42.736 44.226 42.84 48.6 ; 
      RECT 42.304 44.226 42.408 48.6 ; 
      RECT 41.872 44.226 41.976 48.6 ; 
      RECT 41.44 44.226 41.544 48.6 ; 
      RECT 41.008 44.226 41.112 48.6 ; 
      RECT 40.576 44.226 40.68 48.6 ; 
      RECT 40.144 44.226 40.248 48.6 ; 
      RECT 39.712 44.226 39.816 48.6 ; 
      RECT 39.28 44.226 39.384 48.6 ; 
      RECT 38.848 44.226 38.952 48.6 ; 
      RECT 38.416 44.226 38.52 48.6 ; 
      RECT 37.984 44.226 38.088 48.6 ; 
      RECT 37.552 44.226 37.656 48.6 ; 
      RECT 36.7 44.226 37.008 48.6 ; 
      RECT 29.128 44.226 29.436 48.6 ; 
      RECT 28.48 44.226 28.584 48.6 ; 
      RECT 28.048 44.226 28.152 48.6 ; 
      RECT 27.616 44.226 27.72 48.6 ; 
      RECT 27.184 44.226 27.288 48.6 ; 
      RECT 26.752 44.226 26.856 48.6 ; 
      RECT 26.32 44.226 26.424 48.6 ; 
      RECT 25.888 44.226 25.992 48.6 ; 
      RECT 25.456 44.226 25.56 48.6 ; 
      RECT 25.024 44.226 25.128 48.6 ; 
      RECT 24.592 44.226 24.696 48.6 ; 
      RECT 24.16 44.226 24.264 48.6 ; 
      RECT 23.728 44.226 23.832 48.6 ; 
      RECT 23.296 44.226 23.4 48.6 ; 
      RECT 22.864 44.226 22.968 48.6 ; 
      RECT 22.432 44.226 22.536 48.6 ; 
      RECT 22 44.226 22.104 48.6 ; 
      RECT 21.568 44.226 21.672 48.6 ; 
      RECT 21.136 44.226 21.24 48.6 ; 
      RECT 20.704 44.226 20.808 48.6 ; 
      RECT 20.272 44.226 20.376 48.6 ; 
      RECT 19.84 44.226 19.944 48.6 ; 
      RECT 19.408 44.226 19.512 48.6 ; 
      RECT 18.976 44.226 19.08 48.6 ; 
      RECT 18.544 44.226 18.648 48.6 ; 
      RECT 18.112 44.226 18.216 48.6 ; 
      RECT 17.68 44.226 17.784 48.6 ; 
      RECT 17.248 44.226 17.352 48.6 ; 
      RECT 16.816 44.226 16.92 48.6 ; 
      RECT 16.384 44.226 16.488 48.6 ; 
      RECT 15.952 44.226 16.056 48.6 ; 
      RECT 15.52 44.226 15.624 48.6 ; 
      RECT 15.088 44.226 15.192 48.6 ; 
      RECT 14.656 44.226 14.76 48.6 ; 
      RECT 14.224 44.226 14.328 48.6 ; 
      RECT 13.792 44.226 13.896 48.6 ; 
      RECT 13.36 44.226 13.464 48.6 ; 
      RECT 12.928 44.226 13.032 48.6 ; 
      RECT 12.496 44.226 12.6 48.6 ; 
      RECT 12.064 44.226 12.168 48.6 ; 
      RECT 11.632 44.226 11.736 48.6 ; 
      RECT 11.2 44.226 11.304 48.6 ; 
      RECT 10.768 44.226 10.872 48.6 ; 
      RECT 10.336 44.226 10.44 48.6 ; 
      RECT 9.904 44.226 10.008 48.6 ; 
      RECT 9.472 44.226 9.576 48.6 ; 
      RECT 9.04 44.226 9.144 48.6 ; 
      RECT 8.608 44.226 8.712 48.6 ; 
      RECT 8.176 44.226 8.28 48.6 ; 
      RECT 7.744 44.226 7.848 48.6 ; 
      RECT 7.312 44.226 7.416 48.6 ; 
      RECT 6.88 44.226 6.984 48.6 ; 
      RECT 6.448 44.226 6.552 48.6 ; 
      RECT 6.016 44.226 6.12 48.6 ; 
      RECT 5.584 44.226 5.688 48.6 ; 
      RECT 5.152 44.226 5.256 48.6 ; 
      RECT 4.72 44.226 4.824 48.6 ; 
      RECT 4.288 44.226 4.392 48.6 ; 
      RECT 3.856 44.226 3.96 48.6 ; 
      RECT 3.424 44.226 3.528 48.6 ; 
      RECT 2.992 44.226 3.096 48.6 ; 
      RECT 2.56 44.226 2.664 48.6 ; 
      RECT 2.128 44.226 2.232 48.6 ; 
      RECT 1.696 44.226 1.8 48.6 ; 
      RECT 1.264 44.226 1.368 48.6 ; 
      RECT 0.832 44.226 0.936 48.6 ; 
      RECT 0.02 44.226 0.36 48.6 ; 
      RECT 34.564 48.546 35.076 52.92 ; 
      RECT 34.508 51.208 35.076 52.498 ; 
      RECT 33.916 50.116 34.164 52.92 ; 
      RECT 33.86 51.354 34.164 51.968 ; 
      RECT 33.916 48.546 34.02 52.92 ; 
      RECT 33.916 49.03 34.076 49.988 ; 
      RECT 33.916 48.546 34.164 48.902 ; 
      RECT 32.728 50.348 33.552 52.92 ; 
      RECT 33.448 48.546 33.552 52.92 ; 
      RECT 32.728 51.456 33.608 52.488 ; 
      RECT 32.728 48.546 33.12 52.92 ; 
      RECT 31.06 48.546 31.392 52.92 ; 
      RECT 31.06 48.9 31.448 52.642 ; 
      RECT 65.776 48.546 66.116 52.92 ; 
      RECT 65.2 48.546 65.304 52.92 ; 
      RECT 64.768 48.546 64.872 52.92 ; 
      RECT 64.336 48.546 64.44 52.92 ; 
      RECT 63.904 48.546 64.008 52.92 ; 
      RECT 63.472 48.546 63.576 52.92 ; 
      RECT 63.04 48.546 63.144 52.92 ; 
      RECT 62.608 48.546 62.712 52.92 ; 
      RECT 62.176 48.546 62.28 52.92 ; 
      RECT 61.744 48.546 61.848 52.92 ; 
      RECT 61.312 48.546 61.416 52.92 ; 
      RECT 60.88 48.546 60.984 52.92 ; 
      RECT 60.448 48.546 60.552 52.92 ; 
      RECT 60.016 48.546 60.12 52.92 ; 
      RECT 59.584 48.546 59.688 52.92 ; 
      RECT 59.152 48.546 59.256 52.92 ; 
      RECT 58.72 48.546 58.824 52.92 ; 
      RECT 58.288 48.546 58.392 52.92 ; 
      RECT 57.856 48.546 57.96 52.92 ; 
      RECT 57.424 48.546 57.528 52.92 ; 
      RECT 56.992 48.546 57.096 52.92 ; 
      RECT 56.56 48.546 56.664 52.92 ; 
      RECT 56.128 48.546 56.232 52.92 ; 
      RECT 55.696 48.546 55.8 52.92 ; 
      RECT 55.264 48.546 55.368 52.92 ; 
      RECT 54.832 48.546 54.936 52.92 ; 
      RECT 54.4 48.546 54.504 52.92 ; 
      RECT 53.968 48.546 54.072 52.92 ; 
      RECT 53.536 48.546 53.64 52.92 ; 
      RECT 53.104 48.546 53.208 52.92 ; 
      RECT 52.672 48.546 52.776 52.92 ; 
      RECT 52.24 48.546 52.344 52.92 ; 
      RECT 51.808 48.546 51.912 52.92 ; 
      RECT 51.376 48.546 51.48 52.92 ; 
      RECT 50.944 48.546 51.048 52.92 ; 
      RECT 50.512 48.546 50.616 52.92 ; 
      RECT 50.08 48.546 50.184 52.92 ; 
      RECT 49.648 48.546 49.752 52.92 ; 
      RECT 49.216 48.546 49.32 52.92 ; 
      RECT 48.784 48.546 48.888 52.92 ; 
      RECT 48.352 48.546 48.456 52.92 ; 
      RECT 47.92 48.546 48.024 52.92 ; 
      RECT 47.488 48.546 47.592 52.92 ; 
      RECT 47.056 48.546 47.16 52.92 ; 
      RECT 46.624 48.546 46.728 52.92 ; 
      RECT 46.192 48.546 46.296 52.92 ; 
      RECT 45.76 48.546 45.864 52.92 ; 
      RECT 45.328 48.546 45.432 52.92 ; 
      RECT 44.896 48.546 45 52.92 ; 
      RECT 44.464 48.546 44.568 52.92 ; 
      RECT 44.032 48.546 44.136 52.92 ; 
      RECT 43.6 48.546 43.704 52.92 ; 
      RECT 43.168 48.546 43.272 52.92 ; 
      RECT 42.736 48.546 42.84 52.92 ; 
      RECT 42.304 48.546 42.408 52.92 ; 
      RECT 41.872 48.546 41.976 52.92 ; 
      RECT 41.44 48.546 41.544 52.92 ; 
      RECT 41.008 48.546 41.112 52.92 ; 
      RECT 40.576 48.546 40.68 52.92 ; 
      RECT 40.144 48.546 40.248 52.92 ; 
      RECT 39.712 48.546 39.816 52.92 ; 
      RECT 39.28 48.546 39.384 52.92 ; 
      RECT 38.848 48.546 38.952 52.92 ; 
      RECT 38.416 48.546 38.52 52.92 ; 
      RECT 37.984 48.546 38.088 52.92 ; 
      RECT 37.552 48.546 37.656 52.92 ; 
      RECT 36.7 48.546 37.008 52.92 ; 
      RECT 29.128 48.546 29.436 52.92 ; 
      RECT 28.48 48.546 28.584 52.92 ; 
      RECT 28.048 48.546 28.152 52.92 ; 
      RECT 27.616 48.546 27.72 52.92 ; 
      RECT 27.184 48.546 27.288 52.92 ; 
      RECT 26.752 48.546 26.856 52.92 ; 
      RECT 26.32 48.546 26.424 52.92 ; 
      RECT 25.888 48.546 25.992 52.92 ; 
      RECT 25.456 48.546 25.56 52.92 ; 
      RECT 25.024 48.546 25.128 52.92 ; 
      RECT 24.592 48.546 24.696 52.92 ; 
      RECT 24.16 48.546 24.264 52.92 ; 
      RECT 23.728 48.546 23.832 52.92 ; 
      RECT 23.296 48.546 23.4 52.92 ; 
      RECT 22.864 48.546 22.968 52.92 ; 
      RECT 22.432 48.546 22.536 52.92 ; 
      RECT 22 48.546 22.104 52.92 ; 
      RECT 21.568 48.546 21.672 52.92 ; 
      RECT 21.136 48.546 21.24 52.92 ; 
      RECT 20.704 48.546 20.808 52.92 ; 
      RECT 20.272 48.546 20.376 52.92 ; 
      RECT 19.84 48.546 19.944 52.92 ; 
      RECT 19.408 48.546 19.512 52.92 ; 
      RECT 18.976 48.546 19.08 52.92 ; 
      RECT 18.544 48.546 18.648 52.92 ; 
      RECT 18.112 48.546 18.216 52.92 ; 
      RECT 17.68 48.546 17.784 52.92 ; 
      RECT 17.248 48.546 17.352 52.92 ; 
      RECT 16.816 48.546 16.92 52.92 ; 
      RECT 16.384 48.546 16.488 52.92 ; 
      RECT 15.952 48.546 16.056 52.92 ; 
      RECT 15.52 48.546 15.624 52.92 ; 
      RECT 15.088 48.546 15.192 52.92 ; 
      RECT 14.656 48.546 14.76 52.92 ; 
      RECT 14.224 48.546 14.328 52.92 ; 
      RECT 13.792 48.546 13.896 52.92 ; 
      RECT 13.36 48.546 13.464 52.92 ; 
      RECT 12.928 48.546 13.032 52.92 ; 
      RECT 12.496 48.546 12.6 52.92 ; 
      RECT 12.064 48.546 12.168 52.92 ; 
      RECT 11.632 48.546 11.736 52.92 ; 
      RECT 11.2 48.546 11.304 52.92 ; 
      RECT 10.768 48.546 10.872 52.92 ; 
      RECT 10.336 48.546 10.44 52.92 ; 
      RECT 9.904 48.546 10.008 52.92 ; 
      RECT 9.472 48.546 9.576 52.92 ; 
      RECT 9.04 48.546 9.144 52.92 ; 
      RECT 8.608 48.546 8.712 52.92 ; 
      RECT 8.176 48.546 8.28 52.92 ; 
      RECT 7.744 48.546 7.848 52.92 ; 
      RECT 7.312 48.546 7.416 52.92 ; 
      RECT 6.88 48.546 6.984 52.92 ; 
      RECT 6.448 48.546 6.552 52.92 ; 
      RECT 6.016 48.546 6.12 52.92 ; 
      RECT 5.584 48.546 5.688 52.92 ; 
      RECT 5.152 48.546 5.256 52.92 ; 
      RECT 4.72 48.546 4.824 52.92 ; 
      RECT 4.288 48.546 4.392 52.92 ; 
      RECT 3.856 48.546 3.96 52.92 ; 
      RECT 3.424 48.546 3.528 52.92 ; 
      RECT 2.992 48.546 3.096 52.92 ; 
      RECT 2.56 48.546 2.664 52.92 ; 
      RECT 2.128 48.546 2.232 52.92 ; 
      RECT 1.696 48.546 1.8 52.92 ; 
      RECT 1.264 48.546 1.368 52.92 ; 
      RECT 0.832 48.546 0.936 52.92 ; 
      RECT 0.02 48.546 0.36 52.92 ; 
      RECT 34.564 52.866 35.076 57.24 ; 
      RECT 34.508 55.528 35.076 56.818 ; 
      RECT 33.916 54.436 34.164 57.24 ; 
      RECT 33.86 55.674 34.164 56.288 ; 
      RECT 33.916 52.866 34.02 57.24 ; 
      RECT 33.916 53.35 34.076 54.308 ; 
      RECT 33.916 52.866 34.164 53.222 ; 
      RECT 32.728 54.668 33.552 57.24 ; 
      RECT 33.448 52.866 33.552 57.24 ; 
      RECT 32.728 55.776 33.608 56.808 ; 
      RECT 32.728 52.866 33.12 57.24 ; 
      RECT 31.06 52.866 31.392 57.24 ; 
      RECT 31.06 53.22 31.448 56.962 ; 
      RECT 65.776 52.866 66.116 57.24 ; 
      RECT 65.2 52.866 65.304 57.24 ; 
      RECT 64.768 52.866 64.872 57.24 ; 
      RECT 64.336 52.866 64.44 57.24 ; 
      RECT 63.904 52.866 64.008 57.24 ; 
      RECT 63.472 52.866 63.576 57.24 ; 
      RECT 63.04 52.866 63.144 57.24 ; 
      RECT 62.608 52.866 62.712 57.24 ; 
      RECT 62.176 52.866 62.28 57.24 ; 
      RECT 61.744 52.866 61.848 57.24 ; 
      RECT 61.312 52.866 61.416 57.24 ; 
      RECT 60.88 52.866 60.984 57.24 ; 
      RECT 60.448 52.866 60.552 57.24 ; 
      RECT 60.016 52.866 60.12 57.24 ; 
      RECT 59.584 52.866 59.688 57.24 ; 
      RECT 59.152 52.866 59.256 57.24 ; 
      RECT 58.72 52.866 58.824 57.24 ; 
      RECT 58.288 52.866 58.392 57.24 ; 
      RECT 57.856 52.866 57.96 57.24 ; 
      RECT 57.424 52.866 57.528 57.24 ; 
      RECT 56.992 52.866 57.096 57.24 ; 
      RECT 56.56 52.866 56.664 57.24 ; 
      RECT 56.128 52.866 56.232 57.24 ; 
      RECT 55.696 52.866 55.8 57.24 ; 
      RECT 55.264 52.866 55.368 57.24 ; 
      RECT 54.832 52.866 54.936 57.24 ; 
      RECT 54.4 52.866 54.504 57.24 ; 
      RECT 53.968 52.866 54.072 57.24 ; 
      RECT 53.536 52.866 53.64 57.24 ; 
      RECT 53.104 52.866 53.208 57.24 ; 
      RECT 52.672 52.866 52.776 57.24 ; 
      RECT 52.24 52.866 52.344 57.24 ; 
      RECT 51.808 52.866 51.912 57.24 ; 
      RECT 51.376 52.866 51.48 57.24 ; 
      RECT 50.944 52.866 51.048 57.24 ; 
      RECT 50.512 52.866 50.616 57.24 ; 
      RECT 50.08 52.866 50.184 57.24 ; 
      RECT 49.648 52.866 49.752 57.24 ; 
      RECT 49.216 52.866 49.32 57.24 ; 
      RECT 48.784 52.866 48.888 57.24 ; 
      RECT 48.352 52.866 48.456 57.24 ; 
      RECT 47.92 52.866 48.024 57.24 ; 
      RECT 47.488 52.866 47.592 57.24 ; 
      RECT 47.056 52.866 47.16 57.24 ; 
      RECT 46.624 52.866 46.728 57.24 ; 
      RECT 46.192 52.866 46.296 57.24 ; 
      RECT 45.76 52.866 45.864 57.24 ; 
      RECT 45.328 52.866 45.432 57.24 ; 
      RECT 44.896 52.866 45 57.24 ; 
      RECT 44.464 52.866 44.568 57.24 ; 
      RECT 44.032 52.866 44.136 57.24 ; 
      RECT 43.6 52.866 43.704 57.24 ; 
      RECT 43.168 52.866 43.272 57.24 ; 
      RECT 42.736 52.866 42.84 57.24 ; 
      RECT 42.304 52.866 42.408 57.24 ; 
      RECT 41.872 52.866 41.976 57.24 ; 
      RECT 41.44 52.866 41.544 57.24 ; 
      RECT 41.008 52.866 41.112 57.24 ; 
      RECT 40.576 52.866 40.68 57.24 ; 
      RECT 40.144 52.866 40.248 57.24 ; 
      RECT 39.712 52.866 39.816 57.24 ; 
      RECT 39.28 52.866 39.384 57.24 ; 
      RECT 38.848 52.866 38.952 57.24 ; 
      RECT 38.416 52.866 38.52 57.24 ; 
      RECT 37.984 52.866 38.088 57.24 ; 
      RECT 37.552 52.866 37.656 57.24 ; 
      RECT 36.7 52.866 37.008 57.24 ; 
      RECT 29.128 52.866 29.436 57.24 ; 
      RECT 28.48 52.866 28.584 57.24 ; 
      RECT 28.048 52.866 28.152 57.24 ; 
      RECT 27.616 52.866 27.72 57.24 ; 
      RECT 27.184 52.866 27.288 57.24 ; 
      RECT 26.752 52.866 26.856 57.24 ; 
      RECT 26.32 52.866 26.424 57.24 ; 
      RECT 25.888 52.866 25.992 57.24 ; 
      RECT 25.456 52.866 25.56 57.24 ; 
      RECT 25.024 52.866 25.128 57.24 ; 
      RECT 24.592 52.866 24.696 57.24 ; 
      RECT 24.16 52.866 24.264 57.24 ; 
      RECT 23.728 52.866 23.832 57.24 ; 
      RECT 23.296 52.866 23.4 57.24 ; 
      RECT 22.864 52.866 22.968 57.24 ; 
      RECT 22.432 52.866 22.536 57.24 ; 
      RECT 22 52.866 22.104 57.24 ; 
      RECT 21.568 52.866 21.672 57.24 ; 
      RECT 21.136 52.866 21.24 57.24 ; 
      RECT 20.704 52.866 20.808 57.24 ; 
      RECT 20.272 52.866 20.376 57.24 ; 
      RECT 19.84 52.866 19.944 57.24 ; 
      RECT 19.408 52.866 19.512 57.24 ; 
      RECT 18.976 52.866 19.08 57.24 ; 
      RECT 18.544 52.866 18.648 57.24 ; 
      RECT 18.112 52.866 18.216 57.24 ; 
      RECT 17.68 52.866 17.784 57.24 ; 
      RECT 17.248 52.866 17.352 57.24 ; 
      RECT 16.816 52.866 16.92 57.24 ; 
      RECT 16.384 52.866 16.488 57.24 ; 
      RECT 15.952 52.866 16.056 57.24 ; 
      RECT 15.52 52.866 15.624 57.24 ; 
      RECT 15.088 52.866 15.192 57.24 ; 
      RECT 14.656 52.866 14.76 57.24 ; 
      RECT 14.224 52.866 14.328 57.24 ; 
      RECT 13.792 52.866 13.896 57.24 ; 
      RECT 13.36 52.866 13.464 57.24 ; 
      RECT 12.928 52.866 13.032 57.24 ; 
      RECT 12.496 52.866 12.6 57.24 ; 
      RECT 12.064 52.866 12.168 57.24 ; 
      RECT 11.632 52.866 11.736 57.24 ; 
      RECT 11.2 52.866 11.304 57.24 ; 
      RECT 10.768 52.866 10.872 57.24 ; 
      RECT 10.336 52.866 10.44 57.24 ; 
      RECT 9.904 52.866 10.008 57.24 ; 
      RECT 9.472 52.866 9.576 57.24 ; 
      RECT 9.04 52.866 9.144 57.24 ; 
      RECT 8.608 52.866 8.712 57.24 ; 
      RECT 8.176 52.866 8.28 57.24 ; 
      RECT 7.744 52.866 7.848 57.24 ; 
      RECT 7.312 52.866 7.416 57.24 ; 
      RECT 6.88 52.866 6.984 57.24 ; 
      RECT 6.448 52.866 6.552 57.24 ; 
      RECT 6.016 52.866 6.12 57.24 ; 
      RECT 5.584 52.866 5.688 57.24 ; 
      RECT 5.152 52.866 5.256 57.24 ; 
      RECT 4.72 52.866 4.824 57.24 ; 
      RECT 4.288 52.866 4.392 57.24 ; 
      RECT 3.856 52.866 3.96 57.24 ; 
      RECT 3.424 52.866 3.528 57.24 ; 
      RECT 2.992 52.866 3.096 57.24 ; 
      RECT 2.56 52.866 2.664 57.24 ; 
      RECT 2.128 52.866 2.232 57.24 ; 
      RECT 1.696 52.866 1.8 57.24 ; 
      RECT 1.264 52.866 1.368 57.24 ; 
      RECT 0.832 52.866 0.936 57.24 ; 
      RECT 0.02 52.866 0.36 57.24 ; 
      RECT 34.564 57.186 35.076 61.56 ; 
      RECT 34.508 59.848 35.076 61.138 ; 
      RECT 33.916 58.756 34.164 61.56 ; 
      RECT 33.86 59.994 34.164 60.608 ; 
      RECT 33.916 57.186 34.02 61.56 ; 
      RECT 33.916 57.67 34.076 58.628 ; 
      RECT 33.916 57.186 34.164 57.542 ; 
      RECT 32.728 58.988 33.552 61.56 ; 
      RECT 33.448 57.186 33.552 61.56 ; 
      RECT 32.728 60.096 33.608 61.128 ; 
      RECT 32.728 57.186 33.12 61.56 ; 
      RECT 31.06 57.186 31.392 61.56 ; 
      RECT 31.06 57.54 31.448 61.282 ; 
      RECT 65.776 57.186 66.116 61.56 ; 
      RECT 65.2 57.186 65.304 61.56 ; 
      RECT 64.768 57.186 64.872 61.56 ; 
      RECT 64.336 57.186 64.44 61.56 ; 
      RECT 63.904 57.186 64.008 61.56 ; 
      RECT 63.472 57.186 63.576 61.56 ; 
      RECT 63.04 57.186 63.144 61.56 ; 
      RECT 62.608 57.186 62.712 61.56 ; 
      RECT 62.176 57.186 62.28 61.56 ; 
      RECT 61.744 57.186 61.848 61.56 ; 
      RECT 61.312 57.186 61.416 61.56 ; 
      RECT 60.88 57.186 60.984 61.56 ; 
      RECT 60.448 57.186 60.552 61.56 ; 
      RECT 60.016 57.186 60.12 61.56 ; 
      RECT 59.584 57.186 59.688 61.56 ; 
      RECT 59.152 57.186 59.256 61.56 ; 
      RECT 58.72 57.186 58.824 61.56 ; 
      RECT 58.288 57.186 58.392 61.56 ; 
      RECT 57.856 57.186 57.96 61.56 ; 
      RECT 57.424 57.186 57.528 61.56 ; 
      RECT 56.992 57.186 57.096 61.56 ; 
      RECT 56.56 57.186 56.664 61.56 ; 
      RECT 56.128 57.186 56.232 61.56 ; 
      RECT 55.696 57.186 55.8 61.56 ; 
      RECT 55.264 57.186 55.368 61.56 ; 
      RECT 54.832 57.186 54.936 61.56 ; 
      RECT 54.4 57.186 54.504 61.56 ; 
      RECT 53.968 57.186 54.072 61.56 ; 
      RECT 53.536 57.186 53.64 61.56 ; 
      RECT 53.104 57.186 53.208 61.56 ; 
      RECT 52.672 57.186 52.776 61.56 ; 
      RECT 52.24 57.186 52.344 61.56 ; 
      RECT 51.808 57.186 51.912 61.56 ; 
      RECT 51.376 57.186 51.48 61.56 ; 
      RECT 50.944 57.186 51.048 61.56 ; 
      RECT 50.512 57.186 50.616 61.56 ; 
      RECT 50.08 57.186 50.184 61.56 ; 
      RECT 49.648 57.186 49.752 61.56 ; 
      RECT 49.216 57.186 49.32 61.56 ; 
      RECT 48.784 57.186 48.888 61.56 ; 
      RECT 48.352 57.186 48.456 61.56 ; 
      RECT 47.92 57.186 48.024 61.56 ; 
      RECT 47.488 57.186 47.592 61.56 ; 
      RECT 47.056 57.186 47.16 61.56 ; 
      RECT 46.624 57.186 46.728 61.56 ; 
      RECT 46.192 57.186 46.296 61.56 ; 
      RECT 45.76 57.186 45.864 61.56 ; 
      RECT 45.328 57.186 45.432 61.56 ; 
      RECT 44.896 57.186 45 61.56 ; 
      RECT 44.464 57.186 44.568 61.56 ; 
      RECT 44.032 57.186 44.136 61.56 ; 
      RECT 43.6 57.186 43.704 61.56 ; 
      RECT 43.168 57.186 43.272 61.56 ; 
      RECT 42.736 57.186 42.84 61.56 ; 
      RECT 42.304 57.186 42.408 61.56 ; 
      RECT 41.872 57.186 41.976 61.56 ; 
      RECT 41.44 57.186 41.544 61.56 ; 
      RECT 41.008 57.186 41.112 61.56 ; 
      RECT 40.576 57.186 40.68 61.56 ; 
      RECT 40.144 57.186 40.248 61.56 ; 
      RECT 39.712 57.186 39.816 61.56 ; 
      RECT 39.28 57.186 39.384 61.56 ; 
      RECT 38.848 57.186 38.952 61.56 ; 
      RECT 38.416 57.186 38.52 61.56 ; 
      RECT 37.984 57.186 38.088 61.56 ; 
      RECT 37.552 57.186 37.656 61.56 ; 
      RECT 36.7 57.186 37.008 61.56 ; 
      RECT 29.128 57.186 29.436 61.56 ; 
      RECT 28.48 57.186 28.584 61.56 ; 
      RECT 28.048 57.186 28.152 61.56 ; 
      RECT 27.616 57.186 27.72 61.56 ; 
      RECT 27.184 57.186 27.288 61.56 ; 
      RECT 26.752 57.186 26.856 61.56 ; 
      RECT 26.32 57.186 26.424 61.56 ; 
      RECT 25.888 57.186 25.992 61.56 ; 
      RECT 25.456 57.186 25.56 61.56 ; 
      RECT 25.024 57.186 25.128 61.56 ; 
      RECT 24.592 57.186 24.696 61.56 ; 
      RECT 24.16 57.186 24.264 61.56 ; 
      RECT 23.728 57.186 23.832 61.56 ; 
      RECT 23.296 57.186 23.4 61.56 ; 
      RECT 22.864 57.186 22.968 61.56 ; 
      RECT 22.432 57.186 22.536 61.56 ; 
      RECT 22 57.186 22.104 61.56 ; 
      RECT 21.568 57.186 21.672 61.56 ; 
      RECT 21.136 57.186 21.24 61.56 ; 
      RECT 20.704 57.186 20.808 61.56 ; 
      RECT 20.272 57.186 20.376 61.56 ; 
      RECT 19.84 57.186 19.944 61.56 ; 
      RECT 19.408 57.186 19.512 61.56 ; 
      RECT 18.976 57.186 19.08 61.56 ; 
      RECT 18.544 57.186 18.648 61.56 ; 
      RECT 18.112 57.186 18.216 61.56 ; 
      RECT 17.68 57.186 17.784 61.56 ; 
      RECT 17.248 57.186 17.352 61.56 ; 
      RECT 16.816 57.186 16.92 61.56 ; 
      RECT 16.384 57.186 16.488 61.56 ; 
      RECT 15.952 57.186 16.056 61.56 ; 
      RECT 15.52 57.186 15.624 61.56 ; 
      RECT 15.088 57.186 15.192 61.56 ; 
      RECT 14.656 57.186 14.76 61.56 ; 
      RECT 14.224 57.186 14.328 61.56 ; 
      RECT 13.792 57.186 13.896 61.56 ; 
      RECT 13.36 57.186 13.464 61.56 ; 
      RECT 12.928 57.186 13.032 61.56 ; 
      RECT 12.496 57.186 12.6 61.56 ; 
      RECT 12.064 57.186 12.168 61.56 ; 
      RECT 11.632 57.186 11.736 61.56 ; 
      RECT 11.2 57.186 11.304 61.56 ; 
      RECT 10.768 57.186 10.872 61.56 ; 
      RECT 10.336 57.186 10.44 61.56 ; 
      RECT 9.904 57.186 10.008 61.56 ; 
      RECT 9.472 57.186 9.576 61.56 ; 
      RECT 9.04 57.186 9.144 61.56 ; 
      RECT 8.608 57.186 8.712 61.56 ; 
      RECT 8.176 57.186 8.28 61.56 ; 
      RECT 7.744 57.186 7.848 61.56 ; 
      RECT 7.312 57.186 7.416 61.56 ; 
      RECT 6.88 57.186 6.984 61.56 ; 
      RECT 6.448 57.186 6.552 61.56 ; 
      RECT 6.016 57.186 6.12 61.56 ; 
      RECT 5.584 57.186 5.688 61.56 ; 
      RECT 5.152 57.186 5.256 61.56 ; 
      RECT 4.72 57.186 4.824 61.56 ; 
      RECT 4.288 57.186 4.392 61.56 ; 
      RECT 3.856 57.186 3.96 61.56 ; 
      RECT 3.424 57.186 3.528 61.56 ; 
      RECT 2.992 57.186 3.096 61.56 ; 
      RECT 2.56 57.186 2.664 61.56 ; 
      RECT 2.128 57.186 2.232 61.56 ; 
      RECT 1.696 57.186 1.8 61.56 ; 
      RECT 1.264 57.186 1.368 61.56 ; 
      RECT 0.832 57.186 0.936 61.56 ; 
      RECT 0.02 57.186 0.36 61.56 ; 
      RECT 34.564 61.506 35.076 65.88 ; 
      RECT 34.508 64.168 35.076 65.458 ; 
      RECT 33.916 63.076 34.164 65.88 ; 
      RECT 33.86 64.314 34.164 64.928 ; 
      RECT 33.916 61.506 34.02 65.88 ; 
      RECT 33.916 61.99 34.076 62.948 ; 
      RECT 33.916 61.506 34.164 61.862 ; 
      RECT 32.728 63.308 33.552 65.88 ; 
      RECT 33.448 61.506 33.552 65.88 ; 
      RECT 32.728 64.416 33.608 65.448 ; 
      RECT 32.728 61.506 33.12 65.88 ; 
      RECT 31.06 61.506 31.392 65.88 ; 
      RECT 31.06 61.86 31.448 65.602 ; 
      RECT 65.776 61.506 66.116 65.88 ; 
      RECT 65.2 61.506 65.304 65.88 ; 
      RECT 64.768 61.506 64.872 65.88 ; 
      RECT 64.336 61.506 64.44 65.88 ; 
      RECT 63.904 61.506 64.008 65.88 ; 
      RECT 63.472 61.506 63.576 65.88 ; 
      RECT 63.04 61.506 63.144 65.88 ; 
      RECT 62.608 61.506 62.712 65.88 ; 
      RECT 62.176 61.506 62.28 65.88 ; 
      RECT 61.744 61.506 61.848 65.88 ; 
      RECT 61.312 61.506 61.416 65.88 ; 
      RECT 60.88 61.506 60.984 65.88 ; 
      RECT 60.448 61.506 60.552 65.88 ; 
      RECT 60.016 61.506 60.12 65.88 ; 
      RECT 59.584 61.506 59.688 65.88 ; 
      RECT 59.152 61.506 59.256 65.88 ; 
      RECT 58.72 61.506 58.824 65.88 ; 
      RECT 58.288 61.506 58.392 65.88 ; 
      RECT 57.856 61.506 57.96 65.88 ; 
      RECT 57.424 61.506 57.528 65.88 ; 
      RECT 56.992 61.506 57.096 65.88 ; 
      RECT 56.56 61.506 56.664 65.88 ; 
      RECT 56.128 61.506 56.232 65.88 ; 
      RECT 55.696 61.506 55.8 65.88 ; 
      RECT 55.264 61.506 55.368 65.88 ; 
      RECT 54.832 61.506 54.936 65.88 ; 
      RECT 54.4 61.506 54.504 65.88 ; 
      RECT 53.968 61.506 54.072 65.88 ; 
      RECT 53.536 61.506 53.64 65.88 ; 
      RECT 53.104 61.506 53.208 65.88 ; 
      RECT 52.672 61.506 52.776 65.88 ; 
      RECT 52.24 61.506 52.344 65.88 ; 
      RECT 51.808 61.506 51.912 65.88 ; 
      RECT 51.376 61.506 51.48 65.88 ; 
      RECT 50.944 61.506 51.048 65.88 ; 
      RECT 50.512 61.506 50.616 65.88 ; 
      RECT 50.08 61.506 50.184 65.88 ; 
      RECT 49.648 61.506 49.752 65.88 ; 
      RECT 49.216 61.506 49.32 65.88 ; 
      RECT 48.784 61.506 48.888 65.88 ; 
      RECT 48.352 61.506 48.456 65.88 ; 
      RECT 47.92 61.506 48.024 65.88 ; 
      RECT 47.488 61.506 47.592 65.88 ; 
      RECT 47.056 61.506 47.16 65.88 ; 
      RECT 46.624 61.506 46.728 65.88 ; 
      RECT 46.192 61.506 46.296 65.88 ; 
      RECT 45.76 61.506 45.864 65.88 ; 
      RECT 45.328 61.506 45.432 65.88 ; 
      RECT 44.896 61.506 45 65.88 ; 
      RECT 44.464 61.506 44.568 65.88 ; 
      RECT 44.032 61.506 44.136 65.88 ; 
      RECT 43.6 61.506 43.704 65.88 ; 
      RECT 43.168 61.506 43.272 65.88 ; 
      RECT 42.736 61.506 42.84 65.88 ; 
      RECT 42.304 61.506 42.408 65.88 ; 
      RECT 41.872 61.506 41.976 65.88 ; 
      RECT 41.44 61.506 41.544 65.88 ; 
      RECT 41.008 61.506 41.112 65.88 ; 
      RECT 40.576 61.506 40.68 65.88 ; 
      RECT 40.144 61.506 40.248 65.88 ; 
      RECT 39.712 61.506 39.816 65.88 ; 
      RECT 39.28 61.506 39.384 65.88 ; 
      RECT 38.848 61.506 38.952 65.88 ; 
      RECT 38.416 61.506 38.52 65.88 ; 
      RECT 37.984 61.506 38.088 65.88 ; 
      RECT 37.552 61.506 37.656 65.88 ; 
      RECT 36.7 61.506 37.008 65.88 ; 
      RECT 29.128 61.506 29.436 65.88 ; 
      RECT 28.48 61.506 28.584 65.88 ; 
      RECT 28.048 61.506 28.152 65.88 ; 
      RECT 27.616 61.506 27.72 65.88 ; 
      RECT 27.184 61.506 27.288 65.88 ; 
      RECT 26.752 61.506 26.856 65.88 ; 
      RECT 26.32 61.506 26.424 65.88 ; 
      RECT 25.888 61.506 25.992 65.88 ; 
      RECT 25.456 61.506 25.56 65.88 ; 
      RECT 25.024 61.506 25.128 65.88 ; 
      RECT 24.592 61.506 24.696 65.88 ; 
      RECT 24.16 61.506 24.264 65.88 ; 
      RECT 23.728 61.506 23.832 65.88 ; 
      RECT 23.296 61.506 23.4 65.88 ; 
      RECT 22.864 61.506 22.968 65.88 ; 
      RECT 22.432 61.506 22.536 65.88 ; 
      RECT 22 61.506 22.104 65.88 ; 
      RECT 21.568 61.506 21.672 65.88 ; 
      RECT 21.136 61.506 21.24 65.88 ; 
      RECT 20.704 61.506 20.808 65.88 ; 
      RECT 20.272 61.506 20.376 65.88 ; 
      RECT 19.84 61.506 19.944 65.88 ; 
      RECT 19.408 61.506 19.512 65.88 ; 
      RECT 18.976 61.506 19.08 65.88 ; 
      RECT 18.544 61.506 18.648 65.88 ; 
      RECT 18.112 61.506 18.216 65.88 ; 
      RECT 17.68 61.506 17.784 65.88 ; 
      RECT 17.248 61.506 17.352 65.88 ; 
      RECT 16.816 61.506 16.92 65.88 ; 
      RECT 16.384 61.506 16.488 65.88 ; 
      RECT 15.952 61.506 16.056 65.88 ; 
      RECT 15.52 61.506 15.624 65.88 ; 
      RECT 15.088 61.506 15.192 65.88 ; 
      RECT 14.656 61.506 14.76 65.88 ; 
      RECT 14.224 61.506 14.328 65.88 ; 
      RECT 13.792 61.506 13.896 65.88 ; 
      RECT 13.36 61.506 13.464 65.88 ; 
      RECT 12.928 61.506 13.032 65.88 ; 
      RECT 12.496 61.506 12.6 65.88 ; 
      RECT 12.064 61.506 12.168 65.88 ; 
      RECT 11.632 61.506 11.736 65.88 ; 
      RECT 11.2 61.506 11.304 65.88 ; 
      RECT 10.768 61.506 10.872 65.88 ; 
      RECT 10.336 61.506 10.44 65.88 ; 
      RECT 9.904 61.506 10.008 65.88 ; 
      RECT 9.472 61.506 9.576 65.88 ; 
      RECT 9.04 61.506 9.144 65.88 ; 
      RECT 8.608 61.506 8.712 65.88 ; 
      RECT 8.176 61.506 8.28 65.88 ; 
      RECT 7.744 61.506 7.848 65.88 ; 
      RECT 7.312 61.506 7.416 65.88 ; 
      RECT 6.88 61.506 6.984 65.88 ; 
      RECT 6.448 61.506 6.552 65.88 ; 
      RECT 6.016 61.506 6.12 65.88 ; 
      RECT 5.584 61.506 5.688 65.88 ; 
      RECT 5.152 61.506 5.256 65.88 ; 
      RECT 4.72 61.506 4.824 65.88 ; 
      RECT 4.288 61.506 4.392 65.88 ; 
      RECT 3.856 61.506 3.96 65.88 ; 
      RECT 3.424 61.506 3.528 65.88 ; 
      RECT 2.992 61.506 3.096 65.88 ; 
      RECT 2.56 61.506 2.664 65.88 ; 
      RECT 2.128 61.506 2.232 65.88 ; 
      RECT 1.696 61.506 1.8 65.88 ; 
      RECT 1.264 61.506 1.368 65.88 ; 
      RECT 0.832 61.506 0.936 65.88 ; 
      RECT 0.02 61.506 0.36 65.88 ; 
      RECT 34.564 65.826 35.076 70.2 ; 
      RECT 34.508 68.488 35.076 69.778 ; 
      RECT 33.916 67.396 34.164 70.2 ; 
      RECT 33.86 68.634 34.164 69.248 ; 
      RECT 33.916 65.826 34.02 70.2 ; 
      RECT 33.916 66.31 34.076 67.268 ; 
      RECT 33.916 65.826 34.164 66.182 ; 
      RECT 32.728 67.628 33.552 70.2 ; 
      RECT 33.448 65.826 33.552 70.2 ; 
      RECT 32.728 68.736 33.608 69.768 ; 
      RECT 32.728 65.826 33.12 70.2 ; 
      RECT 31.06 65.826 31.392 70.2 ; 
      RECT 31.06 66.18 31.448 69.922 ; 
      RECT 65.776 65.826 66.116 70.2 ; 
      RECT 65.2 65.826 65.304 70.2 ; 
      RECT 64.768 65.826 64.872 70.2 ; 
      RECT 64.336 65.826 64.44 70.2 ; 
      RECT 63.904 65.826 64.008 70.2 ; 
      RECT 63.472 65.826 63.576 70.2 ; 
      RECT 63.04 65.826 63.144 70.2 ; 
      RECT 62.608 65.826 62.712 70.2 ; 
      RECT 62.176 65.826 62.28 70.2 ; 
      RECT 61.744 65.826 61.848 70.2 ; 
      RECT 61.312 65.826 61.416 70.2 ; 
      RECT 60.88 65.826 60.984 70.2 ; 
      RECT 60.448 65.826 60.552 70.2 ; 
      RECT 60.016 65.826 60.12 70.2 ; 
      RECT 59.584 65.826 59.688 70.2 ; 
      RECT 59.152 65.826 59.256 70.2 ; 
      RECT 58.72 65.826 58.824 70.2 ; 
      RECT 58.288 65.826 58.392 70.2 ; 
      RECT 57.856 65.826 57.96 70.2 ; 
      RECT 57.424 65.826 57.528 70.2 ; 
      RECT 56.992 65.826 57.096 70.2 ; 
      RECT 56.56 65.826 56.664 70.2 ; 
      RECT 56.128 65.826 56.232 70.2 ; 
      RECT 55.696 65.826 55.8 70.2 ; 
      RECT 55.264 65.826 55.368 70.2 ; 
      RECT 54.832 65.826 54.936 70.2 ; 
      RECT 54.4 65.826 54.504 70.2 ; 
      RECT 53.968 65.826 54.072 70.2 ; 
      RECT 53.536 65.826 53.64 70.2 ; 
      RECT 53.104 65.826 53.208 70.2 ; 
      RECT 52.672 65.826 52.776 70.2 ; 
      RECT 52.24 65.826 52.344 70.2 ; 
      RECT 51.808 65.826 51.912 70.2 ; 
      RECT 51.376 65.826 51.48 70.2 ; 
      RECT 50.944 65.826 51.048 70.2 ; 
      RECT 50.512 65.826 50.616 70.2 ; 
      RECT 50.08 65.826 50.184 70.2 ; 
      RECT 49.648 65.826 49.752 70.2 ; 
      RECT 49.216 65.826 49.32 70.2 ; 
      RECT 48.784 65.826 48.888 70.2 ; 
      RECT 48.352 65.826 48.456 70.2 ; 
      RECT 47.92 65.826 48.024 70.2 ; 
      RECT 47.488 65.826 47.592 70.2 ; 
      RECT 47.056 65.826 47.16 70.2 ; 
      RECT 46.624 65.826 46.728 70.2 ; 
      RECT 46.192 65.826 46.296 70.2 ; 
      RECT 45.76 65.826 45.864 70.2 ; 
      RECT 45.328 65.826 45.432 70.2 ; 
      RECT 44.896 65.826 45 70.2 ; 
      RECT 44.464 65.826 44.568 70.2 ; 
      RECT 44.032 65.826 44.136 70.2 ; 
      RECT 43.6 65.826 43.704 70.2 ; 
      RECT 43.168 65.826 43.272 70.2 ; 
      RECT 42.736 65.826 42.84 70.2 ; 
      RECT 42.304 65.826 42.408 70.2 ; 
      RECT 41.872 65.826 41.976 70.2 ; 
      RECT 41.44 65.826 41.544 70.2 ; 
      RECT 41.008 65.826 41.112 70.2 ; 
      RECT 40.576 65.826 40.68 70.2 ; 
      RECT 40.144 65.826 40.248 70.2 ; 
      RECT 39.712 65.826 39.816 70.2 ; 
      RECT 39.28 65.826 39.384 70.2 ; 
      RECT 38.848 65.826 38.952 70.2 ; 
      RECT 38.416 65.826 38.52 70.2 ; 
      RECT 37.984 65.826 38.088 70.2 ; 
      RECT 37.552 65.826 37.656 70.2 ; 
      RECT 36.7 65.826 37.008 70.2 ; 
      RECT 29.128 65.826 29.436 70.2 ; 
      RECT 28.48 65.826 28.584 70.2 ; 
      RECT 28.048 65.826 28.152 70.2 ; 
      RECT 27.616 65.826 27.72 70.2 ; 
      RECT 27.184 65.826 27.288 70.2 ; 
      RECT 26.752 65.826 26.856 70.2 ; 
      RECT 26.32 65.826 26.424 70.2 ; 
      RECT 25.888 65.826 25.992 70.2 ; 
      RECT 25.456 65.826 25.56 70.2 ; 
      RECT 25.024 65.826 25.128 70.2 ; 
      RECT 24.592 65.826 24.696 70.2 ; 
      RECT 24.16 65.826 24.264 70.2 ; 
      RECT 23.728 65.826 23.832 70.2 ; 
      RECT 23.296 65.826 23.4 70.2 ; 
      RECT 22.864 65.826 22.968 70.2 ; 
      RECT 22.432 65.826 22.536 70.2 ; 
      RECT 22 65.826 22.104 70.2 ; 
      RECT 21.568 65.826 21.672 70.2 ; 
      RECT 21.136 65.826 21.24 70.2 ; 
      RECT 20.704 65.826 20.808 70.2 ; 
      RECT 20.272 65.826 20.376 70.2 ; 
      RECT 19.84 65.826 19.944 70.2 ; 
      RECT 19.408 65.826 19.512 70.2 ; 
      RECT 18.976 65.826 19.08 70.2 ; 
      RECT 18.544 65.826 18.648 70.2 ; 
      RECT 18.112 65.826 18.216 70.2 ; 
      RECT 17.68 65.826 17.784 70.2 ; 
      RECT 17.248 65.826 17.352 70.2 ; 
      RECT 16.816 65.826 16.92 70.2 ; 
      RECT 16.384 65.826 16.488 70.2 ; 
      RECT 15.952 65.826 16.056 70.2 ; 
      RECT 15.52 65.826 15.624 70.2 ; 
      RECT 15.088 65.826 15.192 70.2 ; 
      RECT 14.656 65.826 14.76 70.2 ; 
      RECT 14.224 65.826 14.328 70.2 ; 
      RECT 13.792 65.826 13.896 70.2 ; 
      RECT 13.36 65.826 13.464 70.2 ; 
      RECT 12.928 65.826 13.032 70.2 ; 
      RECT 12.496 65.826 12.6 70.2 ; 
      RECT 12.064 65.826 12.168 70.2 ; 
      RECT 11.632 65.826 11.736 70.2 ; 
      RECT 11.2 65.826 11.304 70.2 ; 
      RECT 10.768 65.826 10.872 70.2 ; 
      RECT 10.336 65.826 10.44 70.2 ; 
      RECT 9.904 65.826 10.008 70.2 ; 
      RECT 9.472 65.826 9.576 70.2 ; 
      RECT 9.04 65.826 9.144 70.2 ; 
      RECT 8.608 65.826 8.712 70.2 ; 
      RECT 8.176 65.826 8.28 70.2 ; 
      RECT 7.744 65.826 7.848 70.2 ; 
      RECT 7.312 65.826 7.416 70.2 ; 
      RECT 6.88 65.826 6.984 70.2 ; 
      RECT 6.448 65.826 6.552 70.2 ; 
      RECT 6.016 65.826 6.12 70.2 ; 
      RECT 5.584 65.826 5.688 70.2 ; 
      RECT 5.152 65.826 5.256 70.2 ; 
      RECT 4.72 65.826 4.824 70.2 ; 
      RECT 4.288 65.826 4.392 70.2 ; 
      RECT 3.856 65.826 3.96 70.2 ; 
      RECT 3.424 65.826 3.528 70.2 ; 
      RECT 2.992 65.826 3.096 70.2 ; 
      RECT 2.56 65.826 2.664 70.2 ; 
      RECT 2.128 65.826 2.232 70.2 ; 
      RECT 1.696 65.826 1.8 70.2 ; 
      RECT 1.264 65.826 1.368 70.2 ; 
      RECT 0.832 65.826 0.936 70.2 ; 
      RECT 0.02 65.826 0.36 70.2 ; 
      RECT 34.564 70.146 35.076 74.52 ; 
      RECT 34.508 72.808 35.076 74.098 ; 
      RECT 33.916 71.716 34.164 74.52 ; 
      RECT 33.86 72.954 34.164 73.568 ; 
      RECT 33.916 70.146 34.02 74.52 ; 
      RECT 33.916 70.63 34.076 71.588 ; 
      RECT 33.916 70.146 34.164 70.502 ; 
      RECT 32.728 71.948 33.552 74.52 ; 
      RECT 33.448 70.146 33.552 74.52 ; 
      RECT 32.728 73.056 33.608 74.088 ; 
      RECT 32.728 70.146 33.12 74.52 ; 
      RECT 31.06 70.146 31.392 74.52 ; 
      RECT 31.06 70.5 31.448 74.242 ; 
      RECT 65.776 70.146 66.116 74.52 ; 
      RECT 65.2 70.146 65.304 74.52 ; 
      RECT 64.768 70.146 64.872 74.52 ; 
      RECT 64.336 70.146 64.44 74.52 ; 
      RECT 63.904 70.146 64.008 74.52 ; 
      RECT 63.472 70.146 63.576 74.52 ; 
      RECT 63.04 70.146 63.144 74.52 ; 
      RECT 62.608 70.146 62.712 74.52 ; 
      RECT 62.176 70.146 62.28 74.52 ; 
      RECT 61.744 70.146 61.848 74.52 ; 
      RECT 61.312 70.146 61.416 74.52 ; 
      RECT 60.88 70.146 60.984 74.52 ; 
      RECT 60.448 70.146 60.552 74.52 ; 
      RECT 60.016 70.146 60.12 74.52 ; 
      RECT 59.584 70.146 59.688 74.52 ; 
      RECT 59.152 70.146 59.256 74.52 ; 
      RECT 58.72 70.146 58.824 74.52 ; 
      RECT 58.288 70.146 58.392 74.52 ; 
      RECT 57.856 70.146 57.96 74.52 ; 
      RECT 57.424 70.146 57.528 74.52 ; 
      RECT 56.992 70.146 57.096 74.52 ; 
      RECT 56.56 70.146 56.664 74.52 ; 
      RECT 56.128 70.146 56.232 74.52 ; 
      RECT 55.696 70.146 55.8 74.52 ; 
      RECT 55.264 70.146 55.368 74.52 ; 
      RECT 54.832 70.146 54.936 74.52 ; 
      RECT 54.4 70.146 54.504 74.52 ; 
      RECT 53.968 70.146 54.072 74.52 ; 
      RECT 53.536 70.146 53.64 74.52 ; 
      RECT 53.104 70.146 53.208 74.52 ; 
      RECT 52.672 70.146 52.776 74.52 ; 
      RECT 52.24 70.146 52.344 74.52 ; 
      RECT 51.808 70.146 51.912 74.52 ; 
      RECT 51.376 70.146 51.48 74.52 ; 
      RECT 50.944 70.146 51.048 74.52 ; 
      RECT 50.512 70.146 50.616 74.52 ; 
      RECT 50.08 70.146 50.184 74.52 ; 
      RECT 49.648 70.146 49.752 74.52 ; 
      RECT 49.216 70.146 49.32 74.52 ; 
      RECT 48.784 70.146 48.888 74.52 ; 
      RECT 48.352 70.146 48.456 74.52 ; 
      RECT 47.92 70.146 48.024 74.52 ; 
      RECT 47.488 70.146 47.592 74.52 ; 
      RECT 47.056 70.146 47.16 74.52 ; 
      RECT 46.624 70.146 46.728 74.52 ; 
      RECT 46.192 70.146 46.296 74.52 ; 
      RECT 45.76 70.146 45.864 74.52 ; 
      RECT 45.328 70.146 45.432 74.52 ; 
      RECT 44.896 70.146 45 74.52 ; 
      RECT 44.464 70.146 44.568 74.52 ; 
      RECT 44.032 70.146 44.136 74.52 ; 
      RECT 43.6 70.146 43.704 74.52 ; 
      RECT 43.168 70.146 43.272 74.52 ; 
      RECT 42.736 70.146 42.84 74.52 ; 
      RECT 42.304 70.146 42.408 74.52 ; 
      RECT 41.872 70.146 41.976 74.52 ; 
      RECT 41.44 70.146 41.544 74.52 ; 
      RECT 41.008 70.146 41.112 74.52 ; 
      RECT 40.576 70.146 40.68 74.52 ; 
      RECT 40.144 70.146 40.248 74.52 ; 
      RECT 39.712 70.146 39.816 74.52 ; 
      RECT 39.28 70.146 39.384 74.52 ; 
      RECT 38.848 70.146 38.952 74.52 ; 
      RECT 38.416 70.146 38.52 74.52 ; 
      RECT 37.984 70.146 38.088 74.52 ; 
      RECT 37.552 70.146 37.656 74.52 ; 
      RECT 36.7 70.146 37.008 74.52 ; 
      RECT 29.128 70.146 29.436 74.52 ; 
      RECT 28.48 70.146 28.584 74.52 ; 
      RECT 28.048 70.146 28.152 74.52 ; 
      RECT 27.616 70.146 27.72 74.52 ; 
      RECT 27.184 70.146 27.288 74.52 ; 
      RECT 26.752 70.146 26.856 74.52 ; 
      RECT 26.32 70.146 26.424 74.52 ; 
      RECT 25.888 70.146 25.992 74.52 ; 
      RECT 25.456 70.146 25.56 74.52 ; 
      RECT 25.024 70.146 25.128 74.52 ; 
      RECT 24.592 70.146 24.696 74.52 ; 
      RECT 24.16 70.146 24.264 74.52 ; 
      RECT 23.728 70.146 23.832 74.52 ; 
      RECT 23.296 70.146 23.4 74.52 ; 
      RECT 22.864 70.146 22.968 74.52 ; 
      RECT 22.432 70.146 22.536 74.52 ; 
      RECT 22 70.146 22.104 74.52 ; 
      RECT 21.568 70.146 21.672 74.52 ; 
      RECT 21.136 70.146 21.24 74.52 ; 
      RECT 20.704 70.146 20.808 74.52 ; 
      RECT 20.272 70.146 20.376 74.52 ; 
      RECT 19.84 70.146 19.944 74.52 ; 
      RECT 19.408 70.146 19.512 74.52 ; 
      RECT 18.976 70.146 19.08 74.52 ; 
      RECT 18.544 70.146 18.648 74.52 ; 
      RECT 18.112 70.146 18.216 74.52 ; 
      RECT 17.68 70.146 17.784 74.52 ; 
      RECT 17.248 70.146 17.352 74.52 ; 
      RECT 16.816 70.146 16.92 74.52 ; 
      RECT 16.384 70.146 16.488 74.52 ; 
      RECT 15.952 70.146 16.056 74.52 ; 
      RECT 15.52 70.146 15.624 74.52 ; 
      RECT 15.088 70.146 15.192 74.52 ; 
      RECT 14.656 70.146 14.76 74.52 ; 
      RECT 14.224 70.146 14.328 74.52 ; 
      RECT 13.792 70.146 13.896 74.52 ; 
      RECT 13.36 70.146 13.464 74.52 ; 
      RECT 12.928 70.146 13.032 74.52 ; 
      RECT 12.496 70.146 12.6 74.52 ; 
      RECT 12.064 70.146 12.168 74.52 ; 
      RECT 11.632 70.146 11.736 74.52 ; 
      RECT 11.2 70.146 11.304 74.52 ; 
      RECT 10.768 70.146 10.872 74.52 ; 
      RECT 10.336 70.146 10.44 74.52 ; 
      RECT 9.904 70.146 10.008 74.52 ; 
      RECT 9.472 70.146 9.576 74.52 ; 
      RECT 9.04 70.146 9.144 74.52 ; 
      RECT 8.608 70.146 8.712 74.52 ; 
      RECT 8.176 70.146 8.28 74.52 ; 
      RECT 7.744 70.146 7.848 74.52 ; 
      RECT 7.312 70.146 7.416 74.52 ; 
      RECT 6.88 70.146 6.984 74.52 ; 
      RECT 6.448 70.146 6.552 74.52 ; 
      RECT 6.016 70.146 6.12 74.52 ; 
      RECT 5.584 70.146 5.688 74.52 ; 
      RECT 5.152 70.146 5.256 74.52 ; 
      RECT 4.72 70.146 4.824 74.52 ; 
      RECT 4.288 70.146 4.392 74.52 ; 
      RECT 3.856 70.146 3.96 74.52 ; 
      RECT 3.424 70.146 3.528 74.52 ; 
      RECT 2.992 70.146 3.096 74.52 ; 
      RECT 2.56 70.146 2.664 74.52 ; 
      RECT 2.128 70.146 2.232 74.52 ; 
      RECT 1.696 70.146 1.8 74.52 ; 
      RECT 1.264 70.146 1.368 74.52 ; 
      RECT 0.832 70.146 0.936 74.52 ; 
      RECT 0.02 70.146 0.36 74.52 ; 
      RECT 34.564 74.466 35.076 78.84 ; 
      RECT 34.508 77.128 35.076 78.418 ; 
      RECT 33.916 76.036 34.164 78.84 ; 
      RECT 33.86 77.274 34.164 77.888 ; 
      RECT 33.916 74.466 34.02 78.84 ; 
      RECT 33.916 74.95 34.076 75.908 ; 
      RECT 33.916 74.466 34.164 74.822 ; 
      RECT 32.728 76.268 33.552 78.84 ; 
      RECT 33.448 74.466 33.552 78.84 ; 
      RECT 32.728 77.376 33.608 78.408 ; 
      RECT 32.728 74.466 33.12 78.84 ; 
      RECT 31.06 74.466 31.392 78.84 ; 
      RECT 31.06 74.82 31.448 78.562 ; 
      RECT 65.776 74.466 66.116 78.84 ; 
      RECT 65.2 74.466 65.304 78.84 ; 
      RECT 64.768 74.466 64.872 78.84 ; 
      RECT 64.336 74.466 64.44 78.84 ; 
      RECT 63.904 74.466 64.008 78.84 ; 
      RECT 63.472 74.466 63.576 78.84 ; 
      RECT 63.04 74.466 63.144 78.84 ; 
      RECT 62.608 74.466 62.712 78.84 ; 
      RECT 62.176 74.466 62.28 78.84 ; 
      RECT 61.744 74.466 61.848 78.84 ; 
      RECT 61.312 74.466 61.416 78.84 ; 
      RECT 60.88 74.466 60.984 78.84 ; 
      RECT 60.448 74.466 60.552 78.84 ; 
      RECT 60.016 74.466 60.12 78.84 ; 
      RECT 59.584 74.466 59.688 78.84 ; 
      RECT 59.152 74.466 59.256 78.84 ; 
      RECT 58.72 74.466 58.824 78.84 ; 
      RECT 58.288 74.466 58.392 78.84 ; 
      RECT 57.856 74.466 57.96 78.84 ; 
      RECT 57.424 74.466 57.528 78.84 ; 
      RECT 56.992 74.466 57.096 78.84 ; 
      RECT 56.56 74.466 56.664 78.84 ; 
      RECT 56.128 74.466 56.232 78.84 ; 
      RECT 55.696 74.466 55.8 78.84 ; 
      RECT 55.264 74.466 55.368 78.84 ; 
      RECT 54.832 74.466 54.936 78.84 ; 
      RECT 54.4 74.466 54.504 78.84 ; 
      RECT 53.968 74.466 54.072 78.84 ; 
      RECT 53.536 74.466 53.64 78.84 ; 
      RECT 53.104 74.466 53.208 78.84 ; 
      RECT 52.672 74.466 52.776 78.84 ; 
      RECT 52.24 74.466 52.344 78.84 ; 
      RECT 51.808 74.466 51.912 78.84 ; 
      RECT 51.376 74.466 51.48 78.84 ; 
      RECT 50.944 74.466 51.048 78.84 ; 
      RECT 50.512 74.466 50.616 78.84 ; 
      RECT 50.08 74.466 50.184 78.84 ; 
      RECT 49.648 74.466 49.752 78.84 ; 
      RECT 49.216 74.466 49.32 78.84 ; 
      RECT 48.784 74.466 48.888 78.84 ; 
      RECT 48.352 74.466 48.456 78.84 ; 
      RECT 47.92 74.466 48.024 78.84 ; 
      RECT 47.488 74.466 47.592 78.84 ; 
      RECT 47.056 74.466 47.16 78.84 ; 
      RECT 46.624 74.466 46.728 78.84 ; 
      RECT 46.192 74.466 46.296 78.84 ; 
      RECT 45.76 74.466 45.864 78.84 ; 
      RECT 45.328 74.466 45.432 78.84 ; 
      RECT 44.896 74.466 45 78.84 ; 
      RECT 44.464 74.466 44.568 78.84 ; 
      RECT 44.032 74.466 44.136 78.84 ; 
      RECT 43.6 74.466 43.704 78.84 ; 
      RECT 43.168 74.466 43.272 78.84 ; 
      RECT 42.736 74.466 42.84 78.84 ; 
      RECT 42.304 74.466 42.408 78.84 ; 
      RECT 41.872 74.466 41.976 78.84 ; 
      RECT 41.44 74.466 41.544 78.84 ; 
      RECT 41.008 74.466 41.112 78.84 ; 
      RECT 40.576 74.466 40.68 78.84 ; 
      RECT 40.144 74.466 40.248 78.84 ; 
      RECT 39.712 74.466 39.816 78.84 ; 
      RECT 39.28 74.466 39.384 78.84 ; 
      RECT 38.848 74.466 38.952 78.84 ; 
      RECT 38.416 74.466 38.52 78.84 ; 
      RECT 37.984 74.466 38.088 78.84 ; 
      RECT 37.552 74.466 37.656 78.84 ; 
      RECT 36.7 74.466 37.008 78.84 ; 
      RECT 29.128 74.466 29.436 78.84 ; 
      RECT 28.48 74.466 28.584 78.84 ; 
      RECT 28.048 74.466 28.152 78.84 ; 
      RECT 27.616 74.466 27.72 78.84 ; 
      RECT 27.184 74.466 27.288 78.84 ; 
      RECT 26.752 74.466 26.856 78.84 ; 
      RECT 26.32 74.466 26.424 78.84 ; 
      RECT 25.888 74.466 25.992 78.84 ; 
      RECT 25.456 74.466 25.56 78.84 ; 
      RECT 25.024 74.466 25.128 78.84 ; 
      RECT 24.592 74.466 24.696 78.84 ; 
      RECT 24.16 74.466 24.264 78.84 ; 
      RECT 23.728 74.466 23.832 78.84 ; 
      RECT 23.296 74.466 23.4 78.84 ; 
      RECT 22.864 74.466 22.968 78.84 ; 
      RECT 22.432 74.466 22.536 78.84 ; 
      RECT 22 74.466 22.104 78.84 ; 
      RECT 21.568 74.466 21.672 78.84 ; 
      RECT 21.136 74.466 21.24 78.84 ; 
      RECT 20.704 74.466 20.808 78.84 ; 
      RECT 20.272 74.466 20.376 78.84 ; 
      RECT 19.84 74.466 19.944 78.84 ; 
      RECT 19.408 74.466 19.512 78.84 ; 
      RECT 18.976 74.466 19.08 78.84 ; 
      RECT 18.544 74.466 18.648 78.84 ; 
      RECT 18.112 74.466 18.216 78.84 ; 
      RECT 17.68 74.466 17.784 78.84 ; 
      RECT 17.248 74.466 17.352 78.84 ; 
      RECT 16.816 74.466 16.92 78.84 ; 
      RECT 16.384 74.466 16.488 78.84 ; 
      RECT 15.952 74.466 16.056 78.84 ; 
      RECT 15.52 74.466 15.624 78.84 ; 
      RECT 15.088 74.466 15.192 78.84 ; 
      RECT 14.656 74.466 14.76 78.84 ; 
      RECT 14.224 74.466 14.328 78.84 ; 
      RECT 13.792 74.466 13.896 78.84 ; 
      RECT 13.36 74.466 13.464 78.84 ; 
      RECT 12.928 74.466 13.032 78.84 ; 
      RECT 12.496 74.466 12.6 78.84 ; 
      RECT 12.064 74.466 12.168 78.84 ; 
      RECT 11.632 74.466 11.736 78.84 ; 
      RECT 11.2 74.466 11.304 78.84 ; 
      RECT 10.768 74.466 10.872 78.84 ; 
      RECT 10.336 74.466 10.44 78.84 ; 
      RECT 9.904 74.466 10.008 78.84 ; 
      RECT 9.472 74.466 9.576 78.84 ; 
      RECT 9.04 74.466 9.144 78.84 ; 
      RECT 8.608 74.466 8.712 78.84 ; 
      RECT 8.176 74.466 8.28 78.84 ; 
      RECT 7.744 74.466 7.848 78.84 ; 
      RECT 7.312 74.466 7.416 78.84 ; 
      RECT 6.88 74.466 6.984 78.84 ; 
      RECT 6.448 74.466 6.552 78.84 ; 
      RECT 6.016 74.466 6.12 78.84 ; 
      RECT 5.584 74.466 5.688 78.84 ; 
      RECT 5.152 74.466 5.256 78.84 ; 
      RECT 4.72 74.466 4.824 78.84 ; 
      RECT 4.288 74.466 4.392 78.84 ; 
      RECT 3.856 74.466 3.96 78.84 ; 
      RECT 3.424 74.466 3.528 78.84 ; 
      RECT 2.992 74.466 3.096 78.84 ; 
      RECT 2.56 74.466 2.664 78.84 ; 
      RECT 2.128 74.466 2.232 78.84 ; 
      RECT 1.696 74.466 1.8 78.84 ; 
      RECT 1.264 74.466 1.368 78.84 ; 
      RECT 0.832 74.466 0.936 78.84 ; 
      RECT 0.02 74.466 0.36 78.84 ; 
      RECT 34.564 78.786 35.076 83.16 ; 
      RECT 34.508 81.448 35.076 82.738 ; 
      RECT 33.916 80.356 34.164 83.16 ; 
      RECT 33.86 81.594 34.164 82.208 ; 
      RECT 33.916 78.786 34.02 83.16 ; 
      RECT 33.916 79.27 34.076 80.228 ; 
      RECT 33.916 78.786 34.164 79.142 ; 
      RECT 32.728 80.588 33.552 83.16 ; 
      RECT 33.448 78.786 33.552 83.16 ; 
      RECT 32.728 81.696 33.608 82.728 ; 
      RECT 32.728 78.786 33.12 83.16 ; 
      RECT 31.06 78.786 31.392 83.16 ; 
      RECT 31.06 79.14 31.448 82.882 ; 
      RECT 65.776 78.786 66.116 83.16 ; 
      RECT 65.2 78.786 65.304 83.16 ; 
      RECT 64.768 78.786 64.872 83.16 ; 
      RECT 64.336 78.786 64.44 83.16 ; 
      RECT 63.904 78.786 64.008 83.16 ; 
      RECT 63.472 78.786 63.576 83.16 ; 
      RECT 63.04 78.786 63.144 83.16 ; 
      RECT 62.608 78.786 62.712 83.16 ; 
      RECT 62.176 78.786 62.28 83.16 ; 
      RECT 61.744 78.786 61.848 83.16 ; 
      RECT 61.312 78.786 61.416 83.16 ; 
      RECT 60.88 78.786 60.984 83.16 ; 
      RECT 60.448 78.786 60.552 83.16 ; 
      RECT 60.016 78.786 60.12 83.16 ; 
      RECT 59.584 78.786 59.688 83.16 ; 
      RECT 59.152 78.786 59.256 83.16 ; 
      RECT 58.72 78.786 58.824 83.16 ; 
      RECT 58.288 78.786 58.392 83.16 ; 
      RECT 57.856 78.786 57.96 83.16 ; 
      RECT 57.424 78.786 57.528 83.16 ; 
      RECT 56.992 78.786 57.096 83.16 ; 
      RECT 56.56 78.786 56.664 83.16 ; 
      RECT 56.128 78.786 56.232 83.16 ; 
      RECT 55.696 78.786 55.8 83.16 ; 
      RECT 55.264 78.786 55.368 83.16 ; 
      RECT 54.832 78.786 54.936 83.16 ; 
      RECT 54.4 78.786 54.504 83.16 ; 
      RECT 53.968 78.786 54.072 83.16 ; 
      RECT 53.536 78.786 53.64 83.16 ; 
      RECT 53.104 78.786 53.208 83.16 ; 
      RECT 52.672 78.786 52.776 83.16 ; 
      RECT 52.24 78.786 52.344 83.16 ; 
      RECT 51.808 78.786 51.912 83.16 ; 
      RECT 51.376 78.786 51.48 83.16 ; 
      RECT 50.944 78.786 51.048 83.16 ; 
      RECT 50.512 78.786 50.616 83.16 ; 
      RECT 50.08 78.786 50.184 83.16 ; 
      RECT 49.648 78.786 49.752 83.16 ; 
      RECT 49.216 78.786 49.32 83.16 ; 
      RECT 48.784 78.786 48.888 83.16 ; 
      RECT 48.352 78.786 48.456 83.16 ; 
      RECT 47.92 78.786 48.024 83.16 ; 
      RECT 47.488 78.786 47.592 83.16 ; 
      RECT 47.056 78.786 47.16 83.16 ; 
      RECT 46.624 78.786 46.728 83.16 ; 
      RECT 46.192 78.786 46.296 83.16 ; 
      RECT 45.76 78.786 45.864 83.16 ; 
      RECT 45.328 78.786 45.432 83.16 ; 
      RECT 44.896 78.786 45 83.16 ; 
      RECT 44.464 78.786 44.568 83.16 ; 
      RECT 44.032 78.786 44.136 83.16 ; 
      RECT 43.6 78.786 43.704 83.16 ; 
      RECT 43.168 78.786 43.272 83.16 ; 
      RECT 42.736 78.786 42.84 83.16 ; 
      RECT 42.304 78.786 42.408 83.16 ; 
      RECT 41.872 78.786 41.976 83.16 ; 
      RECT 41.44 78.786 41.544 83.16 ; 
      RECT 41.008 78.786 41.112 83.16 ; 
      RECT 40.576 78.786 40.68 83.16 ; 
      RECT 40.144 78.786 40.248 83.16 ; 
      RECT 39.712 78.786 39.816 83.16 ; 
      RECT 39.28 78.786 39.384 83.16 ; 
      RECT 38.848 78.786 38.952 83.16 ; 
      RECT 38.416 78.786 38.52 83.16 ; 
      RECT 37.984 78.786 38.088 83.16 ; 
      RECT 37.552 78.786 37.656 83.16 ; 
      RECT 36.7 78.786 37.008 83.16 ; 
      RECT 29.128 78.786 29.436 83.16 ; 
      RECT 28.48 78.786 28.584 83.16 ; 
      RECT 28.048 78.786 28.152 83.16 ; 
      RECT 27.616 78.786 27.72 83.16 ; 
      RECT 27.184 78.786 27.288 83.16 ; 
      RECT 26.752 78.786 26.856 83.16 ; 
      RECT 26.32 78.786 26.424 83.16 ; 
      RECT 25.888 78.786 25.992 83.16 ; 
      RECT 25.456 78.786 25.56 83.16 ; 
      RECT 25.024 78.786 25.128 83.16 ; 
      RECT 24.592 78.786 24.696 83.16 ; 
      RECT 24.16 78.786 24.264 83.16 ; 
      RECT 23.728 78.786 23.832 83.16 ; 
      RECT 23.296 78.786 23.4 83.16 ; 
      RECT 22.864 78.786 22.968 83.16 ; 
      RECT 22.432 78.786 22.536 83.16 ; 
      RECT 22 78.786 22.104 83.16 ; 
      RECT 21.568 78.786 21.672 83.16 ; 
      RECT 21.136 78.786 21.24 83.16 ; 
      RECT 20.704 78.786 20.808 83.16 ; 
      RECT 20.272 78.786 20.376 83.16 ; 
      RECT 19.84 78.786 19.944 83.16 ; 
      RECT 19.408 78.786 19.512 83.16 ; 
      RECT 18.976 78.786 19.08 83.16 ; 
      RECT 18.544 78.786 18.648 83.16 ; 
      RECT 18.112 78.786 18.216 83.16 ; 
      RECT 17.68 78.786 17.784 83.16 ; 
      RECT 17.248 78.786 17.352 83.16 ; 
      RECT 16.816 78.786 16.92 83.16 ; 
      RECT 16.384 78.786 16.488 83.16 ; 
      RECT 15.952 78.786 16.056 83.16 ; 
      RECT 15.52 78.786 15.624 83.16 ; 
      RECT 15.088 78.786 15.192 83.16 ; 
      RECT 14.656 78.786 14.76 83.16 ; 
      RECT 14.224 78.786 14.328 83.16 ; 
      RECT 13.792 78.786 13.896 83.16 ; 
      RECT 13.36 78.786 13.464 83.16 ; 
      RECT 12.928 78.786 13.032 83.16 ; 
      RECT 12.496 78.786 12.6 83.16 ; 
      RECT 12.064 78.786 12.168 83.16 ; 
      RECT 11.632 78.786 11.736 83.16 ; 
      RECT 11.2 78.786 11.304 83.16 ; 
      RECT 10.768 78.786 10.872 83.16 ; 
      RECT 10.336 78.786 10.44 83.16 ; 
      RECT 9.904 78.786 10.008 83.16 ; 
      RECT 9.472 78.786 9.576 83.16 ; 
      RECT 9.04 78.786 9.144 83.16 ; 
      RECT 8.608 78.786 8.712 83.16 ; 
      RECT 8.176 78.786 8.28 83.16 ; 
      RECT 7.744 78.786 7.848 83.16 ; 
      RECT 7.312 78.786 7.416 83.16 ; 
      RECT 6.88 78.786 6.984 83.16 ; 
      RECT 6.448 78.786 6.552 83.16 ; 
      RECT 6.016 78.786 6.12 83.16 ; 
      RECT 5.584 78.786 5.688 83.16 ; 
      RECT 5.152 78.786 5.256 83.16 ; 
      RECT 4.72 78.786 4.824 83.16 ; 
      RECT 4.288 78.786 4.392 83.16 ; 
      RECT 3.856 78.786 3.96 83.16 ; 
      RECT 3.424 78.786 3.528 83.16 ; 
      RECT 2.992 78.786 3.096 83.16 ; 
      RECT 2.56 78.786 2.664 83.16 ; 
      RECT 2.128 78.786 2.232 83.16 ; 
      RECT 1.696 78.786 1.8 83.16 ; 
      RECT 1.264 78.786 1.368 83.16 ; 
      RECT 0.832 78.786 0.936 83.16 ; 
      RECT 0.02 78.786 0.36 83.16 ; 
      RECT 34.564 83.106 35.076 87.48 ; 
      RECT 34.508 85.768 35.076 87.058 ; 
      RECT 33.916 84.676 34.164 87.48 ; 
      RECT 33.86 85.914 34.164 86.528 ; 
      RECT 33.916 83.106 34.02 87.48 ; 
      RECT 33.916 83.59 34.076 84.548 ; 
      RECT 33.916 83.106 34.164 83.462 ; 
      RECT 32.728 84.908 33.552 87.48 ; 
      RECT 33.448 83.106 33.552 87.48 ; 
      RECT 32.728 86.016 33.608 87.048 ; 
      RECT 32.728 83.106 33.12 87.48 ; 
      RECT 31.06 83.106 31.392 87.48 ; 
      RECT 31.06 83.46 31.448 87.202 ; 
      RECT 65.776 83.106 66.116 87.48 ; 
      RECT 65.2 83.106 65.304 87.48 ; 
      RECT 64.768 83.106 64.872 87.48 ; 
      RECT 64.336 83.106 64.44 87.48 ; 
      RECT 63.904 83.106 64.008 87.48 ; 
      RECT 63.472 83.106 63.576 87.48 ; 
      RECT 63.04 83.106 63.144 87.48 ; 
      RECT 62.608 83.106 62.712 87.48 ; 
      RECT 62.176 83.106 62.28 87.48 ; 
      RECT 61.744 83.106 61.848 87.48 ; 
      RECT 61.312 83.106 61.416 87.48 ; 
      RECT 60.88 83.106 60.984 87.48 ; 
      RECT 60.448 83.106 60.552 87.48 ; 
      RECT 60.016 83.106 60.12 87.48 ; 
      RECT 59.584 83.106 59.688 87.48 ; 
      RECT 59.152 83.106 59.256 87.48 ; 
      RECT 58.72 83.106 58.824 87.48 ; 
      RECT 58.288 83.106 58.392 87.48 ; 
      RECT 57.856 83.106 57.96 87.48 ; 
      RECT 57.424 83.106 57.528 87.48 ; 
      RECT 56.992 83.106 57.096 87.48 ; 
      RECT 56.56 83.106 56.664 87.48 ; 
      RECT 56.128 83.106 56.232 87.48 ; 
      RECT 55.696 83.106 55.8 87.48 ; 
      RECT 55.264 83.106 55.368 87.48 ; 
      RECT 54.832 83.106 54.936 87.48 ; 
      RECT 54.4 83.106 54.504 87.48 ; 
      RECT 53.968 83.106 54.072 87.48 ; 
      RECT 53.536 83.106 53.64 87.48 ; 
      RECT 53.104 83.106 53.208 87.48 ; 
      RECT 52.672 83.106 52.776 87.48 ; 
      RECT 52.24 83.106 52.344 87.48 ; 
      RECT 51.808 83.106 51.912 87.48 ; 
      RECT 51.376 83.106 51.48 87.48 ; 
      RECT 50.944 83.106 51.048 87.48 ; 
      RECT 50.512 83.106 50.616 87.48 ; 
      RECT 50.08 83.106 50.184 87.48 ; 
      RECT 49.648 83.106 49.752 87.48 ; 
      RECT 49.216 83.106 49.32 87.48 ; 
      RECT 48.784 83.106 48.888 87.48 ; 
      RECT 48.352 83.106 48.456 87.48 ; 
      RECT 47.92 83.106 48.024 87.48 ; 
      RECT 47.488 83.106 47.592 87.48 ; 
      RECT 47.056 83.106 47.16 87.48 ; 
      RECT 46.624 83.106 46.728 87.48 ; 
      RECT 46.192 83.106 46.296 87.48 ; 
      RECT 45.76 83.106 45.864 87.48 ; 
      RECT 45.328 83.106 45.432 87.48 ; 
      RECT 44.896 83.106 45 87.48 ; 
      RECT 44.464 83.106 44.568 87.48 ; 
      RECT 44.032 83.106 44.136 87.48 ; 
      RECT 43.6 83.106 43.704 87.48 ; 
      RECT 43.168 83.106 43.272 87.48 ; 
      RECT 42.736 83.106 42.84 87.48 ; 
      RECT 42.304 83.106 42.408 87.48 ; 
      RECT 41.872 83.106 41.976 87.48 ; 
      RECT 41.44 83.106 41.544 87.48 ; 
      RECT 41.008 83.106 41.112 87.48 ; 
      RECT 40.576 83.106 40.68 87.48 ; 
      RECT 40.144 83.106 40.248 87.48 ; 
      RECT 39.712 83.106 39.816 87.48 ; 
      RECT 39.28 83.106 39.384 87.48 ; 
      RECT 38.848 83.106 38.952 87.48 ; 
      RECT 38.416 83.106 38.52 87.48 ; 
      RECT 37.984 83.106 38.088 87.48 ; 
      RECT 37.552 83.106 37.656 87.48 ; 
      RECT 36.7 83.106 37.008 87.48 ; 
      RECT 29.128 83.106 29.436 87.48 ; 
      RECT 28.48 83.106 28.584 87.48 ; 
      RECT 28.048 83.106 28.152 87.48 ; 
      RECT 27.616 83.106 27.72 87.48 ; 
      RECT 27.184 83.106 27.288 87.48 ; 
      RECT 26.752 83.106 26.856 87.48 ; 
      RECT 26.32 83.106 26.424 87.48 ; 
      RECT 25.888 83.106 25.992 87.48 ; 
      RECT 25.456 83.106 25.56 87.48 ; 
      RECT 25.024 83.106 25.128 87.48 ; 
      RECT 24.592 83.106 24.696 87.48 ; 
      RECT 24.16 83.106 24.264 87.48 ; 
      RECT 23.728 83.106 23.832 87.48 ; 
      RECT 23.296 83.106 23.4 87.48 ; 
      RECT 22.864 83.106 22.968 87.48 ; 
      RECT 22.432 83.106 22.536 87.48 ; 
      RECT 22 83.106 22.104 87.48 ; 
      RECT 21.568 83.106 21.672 87.48 ; 
      RECT 21.136 83.106 21.24 87.48 ; 
      RECT 20.704 83.106 20.808 87.48 ; 
      RECT 20.272 83.106 20.376 87.48 ; 
      RECT 19.84 83.106 19.944 87.48 ; 
      RECT 19.408 83.106 19.512 87.48 ; 
      RECT 18.976 83.106 19.08 87.48 ; 
      RECT 18.544 83.106 18.648 87.48 ; 
      RECT 18.112 83.106 18.216 87.48 ; 
      RECT 17.68 83.106 17.784 87.48 ; 
      RECT 17.248 83.106 17.352 87.48 ; 
      RECT 16.816 83.106 16.92 87.48 ; 
      RECT 16.384 83.106 16.488 87.48 ; 
      RECT 15.952 83.106 16.056 87.48 ; 
      RECT 15.52 83.106 15.624 87.48 ; 
      RECT 15.088 83.106 15.192 87.48 ; 
      RECT 14.656 83.106 14.76 87.48 ; 
      RECT 14.224 83.106 14.328 87.48 ; 
      RECT 13.792 83.106 13.896 87.48 ; 
      RECT 13.36 83.106 13.464 87.48 ; 
      RECT 12.928 83.106 13.032 87.48 ; 
      RECT 12.496 83.106 12.6 87.48 ; 
      RECT 12.064 83.106 12.168 87.48 ; 
      RECT 11.632 83.106 11.736 87.48 ; 
      RECT 11.2 83.106 11.304 87.48 ; 
      RECT 10.768 83.106 10.872 87.48 ; 
      RECT 10.336 83.106 10.44 87.48 ; 
      RECT 9.904 83.106 10.008 87.48 ; 
      RECT 9.472 83.106 9.576 87.48 ; 
      RECT 9.04 83.106 9.144 87.48 ; 
      RECT 8.608 83.106 8.712 87.48 ; 
      RECT 8.176 83.106 8.28 87.48 ; 
      RECT 7.744 83.106 7.848 87.48 ; 
      RECT 7.312 83.106 7.416 87.48 ; 
      RECT 6.88 83.106 6.984 87.48 ; 
      RECT 6.448 83.106 6.552 87.48 ; 
      RECT 6.016 83.106 6.12 87.48 ; 
      RECT 5.584 83.106 5.688 87.48 ; 
      RECT 5.152 83.106 5.256 87.48 ; 
      RECT 4.72 83.106 4.824 87.48 ; 
      RECT 4.288 83.106 4.392 87.48 ; 
      RECT 3.856 83.106 3.96 87.48 ; 
      RECT 3.424 83.106 3.528 87.48 ; 
      RECT 2.992 83.106 3.096 87.48 ; 
      RECT 2.56 83.106 2.664 87.48 ; 
      RECT 2.128 83.106 2.232 87.48 ; 
      RECT 1.696 83.106 1.8 87.48 ; 
      RECT 1.264 83.106 1.368 87.48 ; 
      RECT 0.832 83.106 0.936 87.48 ; 
      RECT 0.02 83.106 0.36 87.48 ; 
      RECT 34.564 87.426 35.076 91.8 ; 
      RECT 34.508 90.088 35.076 91.378 ; 
      RECT 33.916 88.996 34.164 91.8 ; 
      RECT 33.86 90.234 34.164 90.848 ; 
      RECT 33.916 87.426 34.02 91.8 ; 
      RECT 33.916 87.91 34.076 88.868 ; 
      RECT 33.916 87.426 34.164 87.782 ; 
      RECT 32.728 89.228 33.552 91.8 ; 
      RECT 33.448 87.426 33.552 91.8 ; 
      RECT 32.728 90.336 33.608 91.368 ; 
      RECT 32.728 87.426 33.12 91.8 ; 
      RECT 31.06 87.426 31.392 91.8 ; 
      RECT 31.06 87.78 31.448 91.522 ; 
      RECT 65.776 87.426 66.116 91.8 ; 
      RECT 65.2 87.426 65.304 91.8 ; 
      RECT 64.768 87.426 64.872 91.8 ; 
      RECT 64.336 87.426 64.44 91.8 ; 
      RECT 63.904 87.426 64.008 91.8 ; 
      RECT 63.472 87.426 63.576 91.8 ; 
      RECT 63.04 87.426 63.144 91.8 ; 
      RECT 62.608 87.426 62.712 91.8 ; 
      RECT 62.176 87.426 62.28 91.8 ; 
      RECT 61.744 87.426 61.848 91.8 ; 
      RECT 61.312 87.426 61.416 91.8 ; 
      RECT 60.88 87.426 60.984 91.8 ; 
      RECT 60.448 87.426 60.552 91.8 ; 
      RECT 60.016 87.426 60.12 91.8 ; 
      RECT 59.584 87.426 59.688 91.8 ; 
      RECT 59.152 87.426 59.256 91.8 ; 
      RECT 58.72 87.426 58.824 91.8 ; 
      RECT 58.288 87.426 58.392 91.8 ; 
      RECT 57.856 87.426 57.96 91.8 ; 
      RECT 57.424 87.426 57.528 91.8 ; 
      RECT 56.992 87.426 57.096 91.8 ; 
      RECT 56.56 87.426 56.664 91.8 ; 
      RECT 56.128 87.426 56.232 91.8 ; 
      RECT 55.696 87.426 55.8 91.8 ; 
      RECT 55.264 87.426 55.368 91.8 ; 
      RECT 54.832 87.426 54.936 91.8 ; 
      RECT 54.4 87.426 54.504 91.8 ; 
      RECT 53.968 87.426 54.072 91.8 ; 
      RECT 53.536 87.426 53.64 91.8 ; 
      RECT 53.104 87.426 53.208 91.8 ; 
      RECT 52.672 87.426 52.776 91.8 ; 
      RECT 52.24 87.426 52.344 91.8 ; 
      RECT 51.808 87.426 51.912 91.8 ; 
      RECT 51.376 87.426 51.48 91.8 ; 
      RECT 50.944 87.426 51.048 91.8 ; 
      RECT 50.512 87.426 50.616 91.8 ; 
      RECT 50.08 87.426 50.184 91.8 ; 
      RECT 49.648 87.426 49.752 91.8 ; 
      RECT 49.216 87.426 49.32 91.8 ; 
      RECT 48.784 87.426 48.888 91.8 ; 
      RECT 48.352 87.426 48.456 91.8 ; 
      RECT 47.92 87.426 48.024 91.8 ; 
      RECT 47.488 87.426 47.592 91.8 ; 
      RECT 47.056 87.426 47.16 91.8 ; 
      RECT 46.624 87.426 46.728 91.8 ; 
      RECT 46.192 87.426 46.296 91.8 ; 
      RECT 45.76 87.426 45.864 91.8 ; 
      RECT 45.328 87.426 45.432 91.8 ; 
      RECT 44.896 87.426 45 91.8 ; 
      RECT 44.464 87.426 44.568 91.8 ; 
      RECT 44.032 87.426 44.136 91.8 ; 
      RECT 43.6 87.426 43.704 91.8 ; 
      RECT 43.168 87.426 43.272 91.8 ; 
      RECT 42.736 87.426 42.84 91.8 ; 
      RECT 42.304 87.426 42.408 91.8 ; 
      RECT 41.872 87.426 41.976 91.8 ; 
      RECT 41.44 87.426 41.544 91.8 ; 
      RECT 41.008 87.426 41.112 91.8 ; 
      RECT 40.576 87.426 40.68 91.8 ; 
      RECT 40.144 87.426 40.248 91.8 ; 
      RECT 39.712 87.426 39.816 91.8 ; 
      RECT 39.28 87.426 39.384 91.8 ; 
      RECT 38.848 87.426 38.952 91.8 ; 
      RECT 38.416 87.426 38.52 91.8 ; 
      RECT 37.984 87.426 38.088 91.8 ; 
      RECT 37.552 87.426 37.656 91.8 ; 
      RECT 36.7 87.426 37.008 91.8 ; 
      RECT 29.128 87.426 29.436 91.8 ; 
      RECT 28.48 87.426 28.584 91.8 ; 
      RECT 28.048 87.426 28.152 91.8 ; 
      RECT 27.616 87.426 27.72 91.8 ; 
      RECT 27.184 87.426 27.288 91.8 ; 
      RECT 26.752 87.426 26.856 91.8 ; 
      RECT 26.32 87.426 26.424 91.8 ; 
      RECT 25.888 87.426 25.992 91.8 ; 
      RECT 25.456 87.426 25.56 91.8 ; 
      RECT 25.024 87.426 25.128 91.8 ; 
      RECT 24.592 87.426 24.696 91.8 ; 
      RECT 24.16 87.426 24.264 91.8 ; 
      RECT 23.728 87.426 23.832 91.8 ; 
      RECT 23.296 87.426 23.4 91.8 ; 
      RECT 22.864 87.426 22.968 91.8 ; 
      RECT 22.432 87.426 22.536 91.8 ; 
      RECT 22 87.426 22.104 91.8 ; 
      RECT 21.568 87.426 21.672 91.8 ; 
      RECT 21.136 87.426 21.24 91.8 ; 
      RECT 20.704 87.426 20.808 91.8 ; 
      RECT 20.272 87.426 20.376 91.8 ; 
      RECT 19.84 87.426 19.944 91.8 ; 
      RECT 19.408 87.426 19.512 91.8 ; 
      RECT 18.976 87.426 19.08 91.8 ; 
      RECT 18.544 87.426 18.648 91.8 ; 
      RECT 18.112 87.426 18.216 91.8 ; 
      RECT 17.68 87.426 17.784 91.8 ; 
      RECT 17.248 87.426 17.352 91.8 ; 
      RECT 16.816 87.426 16.92 91.8 ; 
      RECT 16.384 87.426 16.488 91.8 ; 
      RECT 15.952 87.426 16.056 91.8 ; 
      RECT 15.52 87.426 15.624 91.8 ; 
      RECT 15.088 87.426 15.192 91.8 ; 
      RECT 14.656 87.426 14.76 91.8 ; 
      RECT 14.224 87.426 14.328 91.8 ; 
      RECT 13.792 87.426 13.896 91.8 ; 
      RECT 13.36 87.426 13.464 91.8 ; 
      RECT 12.928 87.426 13.032 91.8 ; 
      RECT 12.496 87.426 12.6 91.8 ; 
      RECT 12.064 87.426 12.168 91.8 ; 
      RECT 11.632 87.426 11.736 91.8 ; 
      RECT 11.2 87.426 11.304 91.8 ; 
      RECT 10.768 87.426 10.872 91.8 ; 
      RECT 10.336 87.426 10.44 91.8 ; 
      RECT 9.904 87.426 10.008 91.8 ; 
      RECT 9.472 87.426 9.576 91.8 ; 
      RECT 9.04 87.426 9.144 91.8 ; 
      RECT 8.608 87.426 8.712 91.8 ; 
      RECT 8.176 87.426 8.28 91.8 ; 
      RECT 7.744 87.426 7.848 91.8 ; 
      RECT 7.312 87.426 7.416 91.8 ; 
      RECT 6.88 87.426 6.984 91.8 ; 
      RECT 6.448 87.426 6.552 91.8 ; 
      RECT 6.016 87.426 6.12 91.8 ; 
      RECT 5.584 87.426 5.688 91.8 ; 
      RECT 5.152 87.426 5.256 91.8 ; 
      RECT 4.72 87.426 4.824 91.8 ; 
      RECT 4.288 87.426 4.392 91.8 ; 
      RECT 3.856 87.426 3.96 91.8 ; 
      RECT 3.424 87.426 3.528 91.8 ; 
      RECT 2.992 87.426 3.096 91.8 ; 
      RECT 2.56 87.426 2.664 91.8 ; 
      RECT 2.128 87.426 2.232 91.8 ; 
      RECT 1.696 87.426 1.8 91.8 ; 
      RECT 1.264 87.426 1.368 91.8 ; 
      RECT 0.832 87.426 0.936 91.8 ; 
      RECT 0.02 87.426 0.36 91.8 ; 
      RECT 34.564 91.746 35.076 96.12 ; 
      RECT 34.508 94.408 35.076 95.698 ; 
      RECT 33.916 93.316 34.164 96.12 ; 
      RECT 33.86 94.554 34.164 95.168 ; 
      RECT 33.916 91.746 34.02 96.12 ; 
      RECT 33.916 92.23 34.076 93.188 ; 
      RECT 33.916 91.746 34.164 92.102 ; 
      RECT 32.728 93.548 33.552 96.12 ; 
      RECT 33.448 91.746 33.552 96.12 ; 
      RECT 32.728 94.656 33.608 95.688 ; 
      RECT 32.728 91.746 33.12 96.12 ; 
      RECT 31.06 91.746 31.392 96.12 ; 
      RECT 31.06 92.1 31.448 95.842 ; 
      RECT 65.776 91.746 66.116 96.12 ; 
      RECT 65.2 91.746 65.304 96.12 ; 
      RECT 64.768 91.746 64.872 96.12 ; 
      RECT 64.336 91.746 64.44 96.12 ; 
      RECT 63.904 91.746 64.008 96.12 ; 
      RECT 63.472 91.746 63.576 96.12 ; 
      RECT 63.04 91.746 63.144 96.12 ; 
      RECT 62.608 91.746 62.712 96.12 ; 
      RECT 62.176 91.746 62.28 96.12 ; 
      RECT 61.744 91.746 61.848 96.12 ; 
      RECT 61.312 91.746 61.416 96.12 ; 
      RECT 60.88 91.746 60.984 96.12 ; 
      RECT 60.448 91.746 60.552 96.12 ; 
      RECT 60.016 91.746 60.12 96.12 ; 
      RECT 59.584 91.746 59.688 96.12 ; 
      RECT 59.152 91.746 59.256 96.12 ; 
      RECT 58.72 91.746 58.824 96.12 ; 
      RECT 58.288 91.746 58.392 96.12 ; 
      RECT 57.856 91.746 57.96 96.12 ; 
      RECT 57.424 91.746 57.528 96.12 ; 
      RECT 56.992 91.746 57.096 96.12 ; 
      RECT 56.56 91.746 56.664 96.12 ; 
      RECT 56.128 91.746 56.232 96.12 ; 
      RECT 55.696 91.746 55.8 96.12 ; 
      RECT 55.264 91.746 55.368 96.12 ; 
      RECT 54.832 91.746 54.936 96.12 ; 
      RECT 54.4 91.746 54.504 96.12 ; 
      RECT 53.968 91.746 54.072 96.12 ; 
      RECT 53.536 91.746 53.64 96.12 ; 
      RECT 53.104 91.746 53.208 96.12 ; 
      RECT 52.672 91.746 52.776 96.12 ; 
      RECT 52.24 91.746 52.344 96.12 ; 
      RECT 51.808 91.746 51.912 96.12 ; 
      RECT 51.376 91.746 51.48 96.12 ; 
      RECT 50.944 91.746 51.048 96.12 ; 
      RECT 50.512 91.746 50.616 96.12 ; 
      RECT 50.08 91.746 50.184 96.12 ; 
      RECT 49.648 91.746 49.752 96.12 ; 
      RECT 49.216 91.746 49.32 96.12 ; 
      RECT 48.784 91.746 48.888 96.12 ; 
      RECT 48.352 91.746 48.456 96.12 ; 
      RECT 47.92 91.746 48.024 96.12 ; 
      RECT 47.488 91.746 47.592 96.12 ; 
      RECT 47.056 91.746 47.16 96.12 ; 
      RECT 46.624 91.746 46.728 96.12 ; 
      RECT 46.192 91.746 46.296 96.12 ; 
      RECT 45.76 91.746 45.864 96.12 ; 
      RECT 45.328 91.746 45.432 96.12 ; 
      RECT 44.896 91.746 45 96.12 ; 
      RECT 44.464 91.746 44.568 96.12 ; 
      RECT 44.032 91.746 44.136 96.12 ; 
      RECT 43.6 91.746 43.704 96.12 ; 
      RECT 43.168 91.746 43.272 96.12 ; 
      RECT 42.736 91.746 42.84 96.12 ; 
      RECT 42.304 91.746 42.408 96.12 ; 
      RECT 41.872 91.746 41.976 96.12 ; 
      RECT 41.44 91.746 41.544 96.12 ; 
      RECT 41.008 91.746 41.112 96.12 ; 
      RECT 40.576 91.746 40.68 96.12 ; 
      RECT 40.144 91.746 40.248 96.12 ; 
      RECT 39.712 91.746 39.816 96.12 ; 
      RECT 39.28 91.746 39.384 96.12 ; 
      RECT 38.848 91.746 38.952 96.12 ; 
      RECT 38.416 91.746 38.52 96.12 ; 
      RECT 37.984 91.746 38.088 96.12 ; 
      RECT 37.552 91.746 37.656 96.12 ; 
      RECT 36.7 91.746 37.008 96.12 ; 
      RECT 29.128 91.746 29.436 96.12 ; 
      RECT 28.48 91.746 28.584 96.12 ; 
      RECT 28.048 91.746 28.152 96.12 ; 
      RECT 27.616 91.746 27.72 96.12 ; 
      RECT 27.184 91.746 27.288 96.12 ; 
      RECT 26.752 91.746 26.856 96.12 ; 
      RECT 26.32 91.746 26.424 96.12 ; 
      RECT 25.888 91.746 25.992 96.12 ; 
      RECT 25.456 91.746 25.56 96.12 ; 
      RECT 25.024 91.746 25.128 96.12 ; 
      RECT 24.592 91.746 24.696 96.12 ; 
      RECT 24.16 91.746 24.264 96.12 ; 
      RECT 23.728 91.746 23.832 96.12 ; 
      RECT 23.296 91.746 23.4 96.12 ; 
      RECT 22.864 91.746 22.968 96.12 ; 
      RECT 22.432 91.746 22.536 96.12 ; 
      RECT 22 91.746 22.104 96.12 ; 
      RECT 21.568 91.746 21.672 96.12 ; 
      RECT 21.136 91.746 21.24 96.12 ; 
      RECT 20.704 91.746 20.808 96.12 ; 
      RECT 20.272 91.746 20.376 96.12 ; 
      RECT 19.84 91.746 19.944 96.12 ; 
      RECT 19.408 91.746 19.512 96.12 ; 
      RECT 18.976 91.746 19.08 96.12 ; 
      RECT 18.544 91.746 18.648 96.12 ; 
      RECT 18.112 91.746 18.216 96.12 ; 
      RECT 17.68 91.746 17.784 96.12 ; 
      RECT 17.248 91.746 17.352 96.12 ; 
      RECT 16.816 91.746 16.92 96.12 ; 
      RECT 16.384 91.746 16.488 96.12 ; 
      RECT 15.952 91.746 16.056 96.12 ; 
      RECT 15.52 91.746 15.624 96.12 ; 
      RECT 15.088 91.746 15.192 96.12 ; 
      RECT 14.656 91.746 14.76 96.12 ; 
      RECT 14.224 91.746 14.328 96.12 ; 
      RECT 13.792 91.746 13.896 96.12 ; 
      RECT 13.36 91.746 13.464 96.12 ; 
      RECT 12.928 91.746 13.032 96.12 ; 
      RECT 12.496 91.746 12.6 96.12 ; 
      RECT 12.064 91.746 12.168 96.12 ; 
      RECT 11.632 91.746 11.736 96.12 ; 
      RECT 11.2 91.746 11.304 96.12 ; 
      RECT 10.768 91.746 10.872 96.12 ; 
      RECT 10.336 91.746 10.44 96.12 ; 
      RECT 9.904 91.746 10.008 96.12 ; 
      RECT 9.472 91.746 9.576 96.12 ; 
      RECT 9.04 91.746 9.144 96.12 ; 
      RECT 8.608 91.746 8.712 96.12 ; 
      RECT 8.176 91.746 8.28 96.12 ; 
      RECT 7.744 91.746 7.848 96.12 ; 
      RECT 7.312 91.746 7.416 96.12 ; 
      RECT 6.88 91.746 6.984 96.12 ; 
      RECT 6.448 91.746 6.552 96.12 ; 
      RECT 6.016 91.746 6.12 96.12 ; 
      RECT 5.584 91.746 5.688 96.12 ; 
      RECT 5.152 91.746 5.256 96.12 ; 
      RECT 4.72 91.746 4.824 96.12 ; 
      RECT 4.288 91.746 4.392 96.12 ; 
      RECT 3.856 91.746 3.96 96.12 ; 
      RECT 3.424 91.746 3.528 96.12 ; 
      RECT 2.992 91.746 3.096 96.12 ; 
      RECT 2.56 91.746 2.664 96.12 ; 
      RECT 2.128 91.746 2.232 96.12 ; 
      RECT 1.696 91.746 1.8 96.12 ; 
      RECT 1.264 91.746 1.368 96.12 ; 
      RECT 0.832 91.746 0.936 96.12 ; 
      RECT 0.02 91.746 0.36 96.12 ; 
      RECT 34.564 96.066 35.076 100.44 ; 
      RECT 34.508 98.728 35.076 100.018 ; 
      RECT 33.916 97.636 34.164 100.44 ; 
      RECT 33.86 98.874 34.164 99.488 ; 
      RECT 33.916 96.066 34.02 100.44 ; 
      RECT 33.916 96.55 34.076 97.508 ; 
      RECT 33.916 96.066 34.164 96.422 ; 
      RECT 32.728 97.868 33.552 100.44 ; 
      RECT 33.448 96.066 33.552 100.44 ; 
      RECT 32.728 98.976 33.608 100.008 ; 
      RECT 32.728 96.066 33.12 100.44 ; 
      RECT 31.06 96.066 31.392 100.44 ; 
      RECT 31.06 96.42 31.448 100.162 ; 
      RECT 65.776 96.066 66.116 100.44 ; 
      RECT 65.2 96.066 65.304 100.44 ; 
      RECT 64.768 96.066 64.872 100.44 ; 
      RECT 64.336 96.066 64.44 100.44 ; 
      RECT 63.904 96.066 64.008 100.44 ; 
      RECT 63.472 96.066 63.576 100.44 ; 
      RECT 63.04 96.066 63.144 100.44 ; 
      RECT 62.608 96.066 62.712 100.44 ; 
      RECT 62.176 96.066 62.28 100.44 ; 
      RECT 61.744 96.066 61.848 100.44 ; 
      RECT 61.312 96.066 61.416 100.44 ; 
      RECT 60.88 96.066 60.984 100.44 ; 
      RECT 60.448 96.066 60.552 100.44 ; 
      RECT 60.016 96.066 60.12 100.44 ; 
      RECT 59.584 96.066 59.688 100.44 ; 
      RECT 59.152 96.066 59.256 100.44 ; 
      RECT 58.72 96.066 58.824 100.44 ; 
      RECT 58.288 96.066 58.392 100.44 ; 
      RECT 57.856 96.066 57.96 100.44 ; 
      RECT 57.424 96.066 57.528 100.44 ; 
      RECT 56.992 96.066 57.096 100.44 ; 
      RECT 56.56 96.066 56.664 100.44 ; 
      RECT 56.128 96.066 56.232 100.44 ; 
      RECT 55.696 96.066 55.8 100.44 ; 
      RECT 55.264 96.066 55.368 100.44 ; 
      RECT 54.832 96.066 54.936 100.44 ; 
      RECT 54.4 96.066 54.504 100.44 ; 
      RECT 53.968 96.066 54.072 100.44 ; 
      RECT 53.536 96.066 53.64 100.44 ; 
      RECT 53.104 96.066 53.208 100.44 ; 
      RECT 52.672 96.066 52.776 100.44 ; 
      RECT 52.24 96.066 52.344 100.44 ; 
      RECT 51.808 96.066 51.912 100.44 ; 
      RECT 51.376 96.066 51.48 100.44 ; 
      RECT 50.944 96.066 51.048 100.44 ; 
      RECT 50.512 96.066 50.616 100.44 ; 
      RECT 50.08 96.066 50.184 100.44 ; 
      RECT 49.648 96.066 49.752 100.44 ; 
      RECT 49.216 96.066 49.32 100.44 ; 
      RECT 48.784 96.066 48.888 100.44 ; 
      RECT 48.352 96.066 48.456 100.44 ; 
      RECT 47.92 96.066 48.024 100.44 ; 
      RECT 47.488 96.066 47.592 100.44 ; 
      RECT 47.056 96.066 47.16 100.44 ; 
      RECT 46.624 96.066 46.728 100.44 ; 
      RECT 46.192 96.066 46.296 100.44 ; 
      RECT 45.76 96.066 45.864 100.44 ; 
      RECT 45.328 96.066 45.432 100.44 ; 
      RECT 44.896 96.066 45 100.44 ; 
      RECT 44.464 96.066 44.568 100.44 ; 
      RECT 44.032 96.066 44.136 100.44 ; 
      RECT 43.6 96.066 43.704 100.44 ; 
      RECT 43.168 96.066 43.272 100.44 ; 
      RECT 42.736 96.066 42.84 100.44 ; 
      RECT 42.304 96.066 42.408 100.44 ; 
      RECT 41.872 96.066 41.976 100.44 ; 
      RECT 41.44 96.066 41.544 100.44 ; 
      RECT 41.008 96.066 41.112 100.44 ; 
      RECT 40.576 96.066 40.68 100.44 ; 
      RECT 40.144 96.066 40.248 100.44 ; 
      RECT 39.712 96.066 39.816 100.44 ; 
      RECT 39.28 96.066 39.384 100.44 ; 
      RECT 38.848 96.066 38.952 100.44 ; 
      RECT 38.416 96.066 38.52 100.44 ; 
      RECT 37.984 96.066 38.088 100.44 ; 
      RECT 37.552 96.066 37.656 100.44 ; 
      RECT 36.7 96.066 37.008 100.44 ; 
      RECT 29.128 96.066 29.436 100.44 ; 
      RECT 28.48 96.066 28.584 100.44 ; 
      RECT 28.048 96.066 28.152 100.44 ; 
      RECT 27.616 96.066 27.72 100.44 ; 
      RECT 27.184 96.066 27.288 100.44 ; 
      RECT 26.752 96.066 26.856 100.44 ; 
      RECT 26.32 96.066 26.424 100.44 ; 
      RECT 25.888 96.066 25.992 100.44 ; 
      RECT 25.456 96.066 25.56 100.44 ; 
      RECT 25.024 96.066 25.128 100.44 ; 
      RECT 24.592 96.066 24.696 100.44 ; 
      RECT 24.16 96.066 24.264 100.44 ; 
      RECT 23.728 96.066 23.832 100.44 ; 
      RECT 23.296 96.066 23.4 100.44 ; 
      RECT 22.864 96.066 22.968 100.44 ; 
      RECT 22.432 96.066 22.536 100.44 ; 
      RECT 22 96.066 22.104 100.44 ; 
      RECT 21.568 96.066 21.672 100.44 ; 
      RECT 21.136 96.066 21.24 100.44 ; 
      RECT 20.704 96.066 20.808 100.44 ; 
      RECT 20.272 96.066 20.376 100.44 ; 
      RECT 19.84 96.066 19.944 100.44 ; 
      RECT 19.408 96.066 19.512 100.44 ; 
      RECT 18.976 96.066 19.08 100.44 ; 
      RECT 18.544 96.066 18.648 100.44 ; 
      RECT 18.112 96.066 18.216 100.44 ; 
      RECT 17.68 96.066 17.784 100.44 ; 
      RECT 17.248 96.066 17.352 100.44 ; 
      RECT 16.816 96.066 16.92 100.44 ; 
      RECT 16.384 96.066 16.488 100.44 ; 
      RECT 15.952 96.066 16.056 100.44 ; 
      RECT 15.52 96.066 15.624 100.44 ; 
      RECT 15.088 96.066 15.192 100.44 ; 
      RECT 14.656 96.066 14.76 100.44 ; 
      RECT 14.224 96.066 14.328 100.44 ; 
      RECT 13.792 96.066 13.896 100.44 ; 
      RECT 13.36 96.066 13.464 100.44 ; 
      RECT 12.928 96.066 13.032 100.44 ; 
      RECT 12.496 96.066 12.6 100.44 ; 
      RECT 12.064 96.066 12.168 100.44 ; 
      RECT 11.632 96.066 11.736 100.44 ; 
      RECT 11.2 96.066 11.304 100.44 ; 
      RECT 10.768 96.066 10.872 100.44 ; 
      RECT 10.336 96.066 10.44 100.44 ; 
      RECT 9.904 96.066 10.008 100.44 ; 
      RECT 9.472 96.066 9.576 100.44 ; 
      RECT 9.04 96.066 9.144 100.44 ; 
      RECT 8.608 96.066 8.712 100.44 ; 
      RECT 8.176 96.066 8.28 100.44 ; 
      RECT 7.744 96.066 7.848 100.44 ; 
      RECT 7.312 96.066 7.416 100.44 ; 
      RECT 6.88 96.066 6.984 100.44 ; 
      RECT 6.448 96.066 6.552 100.44 ; 
      RECT 6.016 96.066 6.12 100.44 ; 
      RECT 5.584 96.066 5.688 100.44 ; 
      RECT 5.152 96.066 5.256 100.44 ; 
      RECT 4.72 96.066 4.824 100.44 ; 
      RECT 4.288 96.066 4.392 100.44 ; 
      RECT 3.856 96.066 3.96 100.44 ; 
      RECT 3.424 96.066 3.528 100.44 ; 
      RECT 2.992 96.066 3.096 100.44 ; 
      RECT 2.56 96.066 2.664 100.44 ; 
      RECT 2.128 96.066 2.232 100.44 ; 
      RECT 1.696 96.066 1.8 100.44 ; 
      RECT 1.264 96.066 1.368 100.44 ; 
      RECT 0.832 96.066 0.936 100.44 ; 
      RECT 0.02 96.066 0.36 100.44 ; 
      RECT 34.564 100.386 35.076 104.76 ; 
      RECT 34.508 103.048 35.076 104.338 ; 
      RECT 33.916 101.956 34.164 104.76 ; 
      RECT 33.86 103.194 34.164 103.808 ; 
      RECT 33.916 100.386 34.02 104.76 ; 
      RECT 33.916 100.87 34.076 101.828 ; 
      RECT 33.916 100.386 34.164 100.742 ; 
      RECT 32.728 102.188 33.552 104.76 ; 
      RECT 33.448 100.386 33.552 104.76 ; 
      RECT 32.728 103.296 33.608 104.328 ; 
      RECT 32.728 100.386 33.12 104.76 ; 
      RECT 31.06 100.386 31.392 104.76 ; 
      RECT 31.06 100.74 31.448 104.482 ; 
      RECT 65.776 100.386 66.116 104.76 ; 
      RECT 65.2 100.386 65.304 104.76 ; 
      RECT 64.768 100.386 64.872 104.76 ; 
      RECT 64.336 100.386 64.44 104.76 ; 
      RECT 63.904 100.386 64.008 104.76 ; 
      RECT 63.472 100.386 63.576 104.76 ; 
      RECT 63.04 100.386 63.144 104.76 ; 
      RECT 62.608 100.386 62.712 104.76 ; 
      RECT 62.176 100.386 62.28 104.76 ; 
      RECT 61.744 100.386 61.848 104.76 ; 
      RECT 61.312 100.386 61.416 104.76 ; 
      RECT 60.88 100.386 60.984 104.76 ; 
      RECT 60.448 100.386 60.552 104.76 ; 
      RECT 60.016 100.386 60.12 104.76 ; 
      RECT 59.584 100.386 59.688 104.76 ; 
      RECT 59.152 100.386 59.256 104.76 ; 
      RECT 58.72 100.386 58.824 104.76 ; 
      RECT 58.288 100.386 58.392 104.76 ; 
      RECT 57.856 100.386 57.96 104.76 ; 
      RECT 57.424 100.386 57.528 104.76 ; 
      RECT 56.992 100.386 57.096 104.76 ; 
      RECT 56.56 100.386 56.664 104.76 ; 
      RECT 56.128 100.386 56.232 104.76 ; 
      RECT 55.696 100.386 55.8 104.76 ; 
      RECT 55.264 100.386 55.368 104.76 ; 
      RECT 54.832 100.386 54.936 104.76 ; 
      RECT 54.4 100.386 54.504 104.76 ; 
      RECT 53.968 100.386 54.072 104.76 ; 
      RECT 53.536 100.386 53.64 104.76 ; 
      RECT 53.104 100.386 53.208 104.76 ; 
      RECT 52.672 100.386 52.776 104.76 ; 
      RECT 52.24 100.386 52.344 104.76 ; 
      RECT 51.808 100.386 51.912 104.76 ; 
      RECT 51.376 100.386 51.48 104.76 ; 
      RECT 50.944 100.386 51.048 104.76 ; 
      RECT 50.512 100.386 50.616 104.76 ; 
      RECT 50.08 100.386 50.184 104.76 ; 
      RECT 49.648 100.386 49.752 104.76 ; 
      RECT 49.216 100.386 49.32 104.76 ; 
      RECT 48.784 100.386 48.888 104.76 ; 
      RECT 48.352 100.386 48.456 104.76 ; 
      RECT 47.92 100.386 48.024 104.76 ; 
      RECT 47.488 100.386 47.592 104.76 ; 
      RECT 47.056 100.386 47.16 104.76 ; 
      RECT 46.624 100.386 46.728 104.76 ; 
      RECT 46.192 100.386 46.296 104.76 ; 
      RECT 45.76 100.386 45.864 104.76 ; 
      RECT 45.328 100.386 45.432 104.76 ; 
      RECT 44.896 100.386 45 104.76 ; 
      RECT 44.464 100.386 44.568 104.76 ; 
      RECT 44.032 100.386 44.136 104.76 ; 
      RECT 43.6 100.386 43.704 104.76 ; 
      RECT 43.168 100.386 43.272 104.76 ; 
      RECT 42.736 100.386 42.84 104.76 ; 
      RECT 42.304 100.386 42.408 104.76 ; 
      RECT 41.872 100.386 41.976 104.76 ; 
      RECT 41.44 100.386 41.544 104.76 ; 
      RECT 41.008 100.386 41.112 104.76 ; 
      RECT 40.576 100.386 40.68 104.76 ; 
      RECT 40.144 100.386 40.248 104.76 ; 
      RECT 39.712 100.386 39.816 104.76 ; 
      RECT 39.28 100.386 39.384 104.76 ; 
      RECT 38.848 100.386 38.952 104.76 ; 
      RECT 38.416 100.386 38.52 104.76 ; 
      RECT 37.984 100.386 38.088 104.76 ; 
      RECT 37.552 100.386 37.656 104.76 ; 
      RECT 36.7 100.386 37.008 104.76 ; 
      RECT 29.128 100.386 29.436 104.76 ; 
      RECT 28.48 100.386 28.584 104.76 ; 
      RECT 28.048 100.386 28.152 104.76 ; 
      RECT 27.616 100.386 27.72 104.76 ; 
      RECT 27.184 100.386 27.288 104.76 ; 
      RECT 26.752 100.386 26.856 104.76 ; 
      RECT 26.32 100.386 26.424 104.76 ; 
      RECT 25.888 100.386 25.992 104.76 ; 
      RECT 25.456 100.386 25.56 104.76 ; 
      RECT 25.024 100.386 25.128 104.76 ; 
      RECT 24.592 100.386 24.696 104.76 ; 
      RECT 24.16 100.386 24.264 104.76 ; 
      RECT 23.728 100.386 23.832 104.76 ; 
      RECT 23.296 100.386 23.4 104.76 ; 
      RECT 22.864 100.386 22.968 104.76 ; 
      RECT 22.432 100.386 22.536 104.76 ; 
      RECT 22 100.386 22.104 104.76 ; 
      RECT 21.568 100.386 21.672 104.76 ; 
      RECT 21.136 100.386 21.24 104.76 ; 
      RECT 20.704 100.386 20.808 104.76 ; 
      RECT 20.272 100.386 20.376 104.76 ; 
      RECT 19.84 100.386 19.944 104.76 ; 
      RECT 19.408 100.386 19.512 104.76 ; 
      RECT 18.976 100.386 19.08 104.76 ; 
      RECT 18.544 100.386 18.648 104.76 ; 
      RECT 18.112 100.386 18.216 104.76 ; 
      RECT 17.68 100.386 17.784 104.76 ; 
      RECT 17.248 100.386 17.352 104.76 ; 
      RECT 16.816 100.386 16.92 104.76 ; 
      RECT 16.384 100.386 16.488 104.76 ; 
      RECT 15.952 100.386 16.056 104.76 ; 
      RECT 15.52 100.386 15.624 104.76 ; 
      RECT 15.088 100.386 15.192 104.76 ; 
      RECT 14.656 100.386 14.76 104.76 ; 
      RECT 14.224 100.386 14.328 104.76 ; 
      RECT 13.792 100.386 13.896 104.76 ; 
      RECT 13.36 100.386 13.464 104.76 ; 
      RECT 12.928 100.386 13.032 104.76 ; 
      RECT 12.496 100.386 12.6 104.76 ; 
      RECT 12.064 100.386 12.168 104.76 ; 
      RECT 11.632 100.386 11.736 104.76 ; 
      RECT 11.2 100.386 11.304 104.76 ; 
      RECT 10.768 100.386 10.872 104.76 ; 
      RECT 10.336 100.386 10.44 104.76 ; 
      RECT 9.904 100.386 10.008 104.76 ; 
      RECT 9.472 100.386 9.576 104.76 ; 
      RECT 9.04 100.386 9.144 104.76 ; 
      RECT 8.608 100.386 8.712 104.76 ; 
      RECT 8.176 100.386 8.28 104.76 ; 
      RECT 7.744 100.386 7.848 104.76 ; 
      RECT 7.312 100.386 7.416 104.76 ; 
      RECT 6.88 100.386 6.984 104.76 ; 
      RECT 6.448 100.386 6.552 104.76 ; 
      RECT 6.016 100.386 6.12 104.76 ; 
      RECT 5.584 100.386 5.688 104.76 ; 
      RECT 5.152 100.386 5.256 104.76 ; 
      RECT 4.72 100.386 4.824 104.76 ; 
      RECT 4.288 100.386 4.392 104.76 ; 
      RECT 3.856 100.386 3.96 104.76 ; 
      RECT 3.424 100.386 3.528 104.76 ; 
      RECT 2.992 100.386 3.096 104.76 ; 
      RECT 2.56 100.386 2.664 104.76 ; 
      RECT 2.128 100.386 2.232 104.76 ; 
      RECT 1.696 100.386 1.8 104.76 ; 
      RECT 1.264 100.386 1.368 104.76 ; 
      RECT 0.832 100.386 0.936 104.76 ; 
      RECT 0.02 100.386 0.36 104.76 ; 
      RECT 0 137.478 66.096 139.242 ; 
      RECT 65.756 104.628 66.096 139.242 ; 
      RECT 37.532 110.644 65.284 139.242 ; 
      RECT 43.364 104.628 65.284 139.242 ; 
      RECT 28.892 137.448 37.204 139.242 ; 
      RECT 31.988 137.322 37.204 139.242 ; 
      RECT 0.812 109.864 28.564 139.242 ; 
      RECT 27.38 104.628 28.564 139.242 ; 
      RECT 0 104.628 0.34 139.242 ; 
      RECT 28.892 111.076 31.372 139.242 ; 
      RECT 31.988 137.304 37.06 139.242 ; 
      RECT 34.58 110.248 37.06 139.242 ; 
      RECT 34.544 136.276 37.06 139.242 ; 
      RECT 33.896 136.276 34.144 139.242 ; 
      RECT 31.988 136.276 33.532 139.242 ; 
      RECT 37.532 119.8 65.34 137.216 ; 
      RECT 0.756 119.8 28.564 137.216 ; 
      RECT 37.476 119.8 65.34 137.198 ; 
      RECT 0.756 119.8 28.62 137.198 ; 
      RECT 28.836 119.8 31.372 137.194 ; 
      RECT 32.708 107.368 33.388 139.242 ; 
      RECT 33.14 104.628 33.388 139.242 ; 
      RECT 29.972 106.312 31.516 135.688 ; 
      RECT 28.836 135.508 31.572 135.656 ; 
      RECT 34.524 131.212 37.06 135.644 ; 
      RECT 32.652 134.452 33.388 135.356 ; 
      RECT 32.708 132.148 33.444 133.196 ; 
      RECT 28.836 131.356 31.572 133.196 ; 
      RECT 32.652 129.196 33.388 131.036 ; 
      RECT 34.524 121.06 37.06 130.388 ; 
      RECT 28.836 123.652 31.572 128.228 ; 
      RECT 32.708 122.572 33.444 127.796 ; 
      RECT 32.652 124.876 33.444 126.716 ; 
      RECT 32.652 111.916 33.388 124.556 ; 
      RECT 32.652 111.916 33.444 122.396 ; 
      RECT 28.836 121.492 31.572 122.396 ; 
      RECT 34.58 110.248 37.204 119.672 ; 
      RECT 34.524 109.756 36.988 116.9 ; 
      RECT 28.892 113.644 31.572 115.124 ; 
      RECT 32.708 110.836 33.444 111.596 ; 
      RECT 29.108 110.692 31.572 111.452 ; 
      RECT 32.652 110.26 33.388 110.804 ; 
      RECT 29.108 107.692 31.516 135.688 ; 
      RECT 32.708 109.756 33.444 110.66 ; 
      RECT 38.18 109.876 65.284 139.242 ; 
      RECT 42.5 109.864 65.284 139.242 ; 
      RECT 37.532 104.628 37.852 139.242 ; 
      RECT 28.892 107.368 29.644 110.624 ; 
      RECT 37.532 104.628 38.716 110.24 ; 
      RECT 37.532 109.096 42.172 110.24 ; 
      RECT 42.5 104.628 43.036 139.242 ; 
      RECT 23.924 108.34 27.052 139.242 ; 
      RECT 0.812 104.628 23.596 139.242 ; 
      RECT 34.58 107.692 36.988 139.242 ; 
      RECT 34.724 105.334 37.204 109.628 ; 
      RECT 37.532 109.096 43.036 109.472 ; 
      RECT 41.636 104.628 65.284 109.46 ; 
      RECT 26.516 104.628 28.564 109.46 ; 
      RECT 32.652 109.18 33.444 109.436 ; 
      RECT 32.652 108.676 33.388 109.436 ; 
      RECT 40.772 107.56 65.284 109.46 ; 
      RECT 37.532 107.692 40.444 110.24 ; 
      RECT 32.708 107.596 33.444 108.644 ; 
      RECT 0.812 107.56 26.188 109.46 ; 
      RECT 25.652 104.628 26.188 139.242 ; 
      RECT 39.908 104.628 41.308 108.116 ; 
      RECT 37.532 107.368 39.58 110.24 ; 
      RECT 39.044 104.628 39.58 139.242 ; 
      RECT 24.788 107.368 26.188 139.242 ; 
      RECT 0.812 104.628 24.46 109.46 ; 
      RECT 32.708 104.628 32.812 139.242 ; 
      RECT 29.252 104.628 29.644 139.242 ; 
      RECT 24.788 104.628 25.324 139.242 ; 
      RECT 39.044 104.628 41.308 107.168 ; 
      RECT 34.58 104.628 36.988 107.168 ; 
      RECT 29.252 104.628 31.372 107.168 ; 
      RECT 25.652 104.628 28.564 107.168 ; 
      RECT 39.044 104.628 65.284 107.156 ; 
      RECT 0.812 104.628 25.324 107.156 ; 
      RECT 34.524 106.516 37.204 107.132 ; 
      RECT 37.532 104.628 65.284 106.1 ; 
      RECT 32.708 104.628 33.388 106.1 ; 
      RECT 28.892 104.628 31.372 106.1 ; 
      RECT 0.812 104.628 28.564 106.1 ; 
      RECT 31.988 104.628 33.388 105.688 ; 
      RECT 34.544 104.628 36.988 105.288 ; 
      RECT 31.988 104.628 33.532 105.288 ; 
      RECT 39.06 104.522 39.132 139.242 ; 
      RECT 38.628 104.522 38.7 139.242 ; 
      RECT 27.396 104.572 27.468 139.242 ; 
      RECT 26.964 104.572 27.036 139.242 ; 
      RECT 26.532 104.572 26.604 139.242 ; 
      RECT 26.1 104.572 26.172 139.242 ; 
      RECT 25.668 104.522 25.74 139.242 ; 
      RECT 25.236 104.522 25.308 139.242 ; 
      RECT 24.804 104.572 24.876 139.242 ; 
      RECT 24.372 104.572 24.444 139.242 ; 
      RECT 23.94 104.572 24.012 139.242 ; 
      RECT 23.508 104.572 23.58 139.242 ; 
      RECT 33.896 104.628 34.144 105.288 ; 
        RECT 34.564 137.214 35.076 141.588 ; 
        RECT 34.508 139.876 35.076 141.166 ; 
        RECT 33.916 138.784 34.164 141.588 ; 
        RECT 33.86 140.022 34.164 140.636 ; 
        RECT 33.916 137.214 34.02 141.588 ; 
        RECT 33.916 137.698 34.076 138.656 ; 
        RECT 33.916 137.214 34.164 137.57 ; 
        RECT 32.728 139.016 33.552 141.588 ; 
        RECT 33.448 137.214 33.552 141.588 ; 
        RECT 32.728 140.124 33.608 141.156 ; 
        RECT 32.728 137.214 33.12 141.588 ; 
        RECT 31.06 137.214 31.392 141.588 ; 
        RECT 31.06 137.568 31.448 141.31 ; 
        RECT 65.776 137.214 66.116 141.588 ; 
        RECT 65.2 137.214 65.304 141.588 ; 
        RECT 64.768 137.214 64.872 141.588 ; 
        RECT 64.336 137.214 64.44 141.588 ; 
        RECT 63.904 137.214 64.008 141.588 ; 
        RECT 63.472 137.214 63.576 141.588 ; 
        RECT 63.04 137.214 63.144 141.588 ; 
        RECT 62.608 137.214 62.712 141.588 ; 
        RECT 62.176 137.214 62.28 141.588 ; 
        RECT 61.744 137.214 61.848 141.588 ; 
        RECT 61.312 137.214 61.416 141.588 ; 
        RECT 60.88 137.214 60.984 141.588 ; 
        RECT 60.448 137.214 60.552 141.588 ; 
        RECT 60.016 137.214 60.12 141.588 ; 
        RECT 59.584 137.214 59.688 141.588 ; 
        RECT 59.152 137.214 59.256 141.588 ; 
        RECT 58.72 137.214 58.824 141.588 ; 
        RECT 58.288 137.214 58.392 141.588 ; 
        RECT 57.856 137.214 57.96 141.588 ; 
        RECT 57.424 137.214 57.528 141.588 ; 
        RECT 56.992 137.214 57.096 141.588 ; 
        RECT 56.56 137.214 56.664 141.588 ; 
        RECT 56.128 137.214 56.232 141.588 ; 
        RECT 55.696 137.214 55.8 141.588 ; 
        RECT 55.264 137.214 55.368 141.588 ; 
        RECT 54.832 137.214 54.936 141.588 ; 
        RECT 54.4 137.214 54.504 141.588 ; 
        RECT 53.968 137.214 54.072 141.588 ; 
        RECT 53.536 137.214 53.64 141.588 ; 
        RECT 53.104 137.214 53.208 141.588 ; 
        RECT 52.672 137.214 52.776 141.588 ; 
        RECT 52.24 137.214 52.344 141.588 ; 
        RECT 51.808 137.214 51.912 141.588 ; 
        RECT 51.376 137.214 51.48 141.588 ; 
        RECT 50.944 137.214 51.048 141.588 ; 
        RECT 50.512 137.214 50.616 141.588 ; 
        RECT 50.08 137.214 50.184 141.588 ; 
        RECT 49.648 137.214 49.752 141.588 ; 
        RECT 49.216 137.214 49.32 141.588 ; 
        RECT 48.784 137.214 48.888 141.588 ; 
        RECT 48.352 137.214 48.456 141.588 ; 
        RECT 47.92 137.214 48.024 141.588 ; 
        RECT 47.488 137.214 47.592 141.588 ; 
        RECT 47.056 137.214 47.16 141.588 ; 
        RECT 46.624 137.214 46.728 141.588 ; 
        RECT 46.192 137.214 46.296 141.588 ; 
        RECT 45.76 137.214 45.864 141.588 ; 
        RECT 45.328 137.214 45.432 141.588 ; 
        RECT 44.896 137.214 45 141.588 ; 
        RECT 44.464 137.214 44.568 141.588 ; 
        RECT 44.032 137.214 44.136 141.588 ; 
        RECT 43.6 137.214 43.704 141.588 ; 
        RECT 43.168 137.214 43.272 141.588 ; 
        RECT 42.736 137.214 42.84 141.588 ; 
        RECT 42.304 137.214 42.408 141.588 ; 
        RECT 41.872 137.214 41.976 141.588 ; 
        RECT 41.44 137.214 41.544 141.588 ; 
        RECT 41.008 137.214 41.112 141.588 ; 
        RECT 40.576 137.214 40.68 141.588 ; 
        RECT 40.144 137.214 40.248 141.588 ; 
        RECT 39.712 137.214 39.816 141.588 ; 
        RECT 39.28 137.214 39.384 141.588 ; 
        RECT 38.848 137.214 38.952 141.588 ; 
        RECT 38.416 137.214 38.52 141.588 ; 
        RECT 37.984 137.214 38.088 141.588 ; 
        RECT 37.552 137.214 37.656 141.588 ; 
        RECT 36.7 137.214 37.008 141.588 ; 
        RECT 29.128 137.214 29.436 141.588 ; 
        RECT 28.48 137.214 28.584 141.588 ; 
        RECT 28.048 137.214 28.152 141.588 ; 
        RECT 27.616 137.214 27.72 141.588 ; 
        RECT 27.184 137.214 27.288 141.588 ; 
        RECT 26.752 137.214 26.856 141.588 ; 
        RECT 26.32 137.214 26.424 141.588 ; 
        RECT 25.888 137.214 25.992 141.588 ; 
        RECT 25.456 137.214 25.56 141.588 ; 
        RECT 25.024 137.214 25.128 141.588 ; 
        RECT 24.592 137.214 24.696 141.588 ; 
        RECT 24.16 137.214 24.264 141.588 ; 
        RECT 23.728 137.214 23.832 141.588 ; 
        RECT 23.296 137.214 23.4 141.588 ; 
        RECT 22.864 137.214 22.968 141.588 ; 
        RECT 22.432 137.214 22.536 141.588 ; 
        RECT 22 137.214 22.104 141.588 ; 
        RECT 21.568 137.214 21.672 141.588 ; 
        RECT 21.136 137.214 21.24 141.588 ; 
        RECT 20.704 137.214 20.808 141.588 ; 
        RECT 20.272 137.214 20.376 141.588 ; 
        RECT 19.84 137.214 19.944 141.588 ; 
        RECT 19.408 137.214 19.512 141.588 ; 
        RECT 18.976 137.214 19.08 141.588 ; 
        RECT 18.544 137.214 18.648 141.588 ; 
        RECT 18.112 137.214 18.216 141.588 ; 
        RECT 17.68 137.214 17.784 141.588 ; 
        RECT 17.248 137.214 17.352 141.588 ; 
        RECT 16.816 137.214 16.92 141.588 ; 
        RECT 16.384 137.214 16.488 141.588 ; 
        RECT 15.952 137.214 16.056 141.588 ; 
        RECT 15.52 137.214 15.624 141.588 ; 
        RECT 15.088 137.214 15.192 141.588 ; 
        RECT 14.656 137.214 14.76 141.588 ; 
        RECT 14.224 137.214 14.328 141.588 ; 
        RECT 13.792 137.214 13.896 141.588 ; 
        RECT 13.36 137.214 13.464 141.588 ; 
        RECT 12.928 137.214 13.032 141.588 ; 
        RECT 12.496 137.214 12.6 141.588 ; 
        RECT 12.064 137.214 12.168 141.588 ; 
        RECT 11.632 137.214 11.736 141.588 ; 
        RECT 11.2 137.214 11.304 141.588 ; 
        RECT 10.768 137.214 10.872 141.588 ; 
        RECT 10.336 137.214 10.44 141.588 ; 
        RECT 9.904 137.214 10.008 141.588 ; 
        RECT 9.472 137.214 9.576 141.588 ; 
        RECT 9.04 137.214 9.144 141.588 ; 
        RECT 8.608 137.214 8.712 141.588 ; 
        RECT 8.176 137.214 8.28 141.588 ; 
        RECT 7.744 137.214 7.848 141.588 ; 
        RECT 7.312 137.214 7.416 141.588 ; 
        RECT 6.88 137.214 6.984 141.588 ; 
        RECT 6.448 137.214 6.552 141.588 ; 
        RECT 6.016 137.214 6.12 141.588 ; 
        RECT 5.584 137.214 5.688 141.588 ; 
        RECT 5.152 137.214 5.256 141.588 ; 
        RECT 4.72 137.214 4.824 141.588 ; 
        RECT 4.288 137.214 4.392 141.588 ; 
        RECT 3.856 137.214 3.96 141.588 ; 
        RECT 3.424 137.214 3.528 141.588 ; 
        RECT 2.992 137.214 3.096 141.588 ; 
        RECT 2.56 137.214 2.664 141.588 ; 
        RECT 2.128 137.214 2.232 141.588 ; 
        RECT 1.696 137.214 1.8 141.588 ; 
        RECT 1.264 137.214 1.368 141.588 ; 
        RECT 0.832 137.214 0.936 141.588 ; 
        RECT 0.02 137.214 0.36 141.588 ; 
        RECT 34.564 141.534 35.076 145.908 ; 
        RECT 34.508 144.196 35.076 145.486 ; 
        RECT 33.916 143.104 34.164 145.908 ; 
        RECT 33.86 144.342 34.164 144.956 ; 
        RECT 33.916 141.534 34.02 145.908 ; 
        RECT 33.916 142.018 34.076 142.976 ; 
        RECT 33.916 141.534 34.164 141.89 ; 
        RECT 32.728 143.336 33.552 145.908 ; 
        RECT 33.448 141.534 33.552 145.908 ; 
        RECT 32.728 144.444 33.608 145.476 ; 
        RECT 32.728 141.534 33.12 145.908 ; 
        RECT 31.06 141.534 31.392 145.908 ; 
        RECT 31.06 141.888 31.448 145.63 ; 
        RECT 65.776 141.534 66.116 145.908 ; 
        RECT 65.2 141.534 65.304 145.908 ; 
        RECT 64.768 141.534 64.872 145.908 ; 
        RECT 64.336 141.534 64.44 145.908 ; 
        RECT 63.904 141.534 64.008 145.908 ; 
        RECT 63.472 141.534 63.576 145.908 ; 
        RECT 63.04 141.534 63.144 145.908 ; 
        RECT 62.608 141.534 62.712 145.908 ; 
        RECT 62.176 141.534 62.28 145.908 ; 
        RECT 61.744 141.534 61.848 145.908 ; 
        RECT 61.312 141.534 61.416 145.908 ; 
        RECT 60.88 141.534 60.984 145.908 ; 
        RECT 60.448 141.534 60.552 145.908 ; 
        RECT 60.016 141.534 60.12 145.908 ; 
        RECT 59.584 141.534 59.688 145.908 ; 
        RECT 59.152 141.534 59.256 145.908 ; 
        RECT 58.72 141.534 58.824 145.908 ; 
        RECT 58.288 141.534 58.392 145.908 ; 
        RECT 57.856 141.534 57.96 145.908 ; 
        RECT 57.424 141.534 57.528 145.908 ; 
        RECT 56.992 141.534 57.096 145.908 ; 
        RECT 56.56 141.534 56.664 145.908 ; 
        RECT 56.128 141.534 56.232 145.908 ; 
        RECT 55.696 141.534 55.8 145.908 ; 
        RECT 55.264 141.534 55.368 145.908 ; 
        RECT 54.832 141.534 54.936 145.908 ; 
        RECT 54.4 141.534 54.504 145.908 ; 
        RECT 53.968 141.534 54.072 145.908 ; 
        RECT 53.536 141.534 53.64 145.908 ; 
        RECT 53.104 141.534 53.208 145.908 ; 
        RECT 52.672 141.534 52.776 145.908 ; 
        RECT 52.24 141.534 52.344 145.908 ; 
        RECT 51.808 141.534 51.912 145.908 ; 
        RECT 51.376 141.534 51.48 145.908 ; 
        RECT 50.944 141.534 51.048 145.908 ; 
        RECT 50.512 141.534 50.616 145.908 ; 
        RECT 50.08 141.534 50.184 145.908 ; 
        RECT 49.648 141.534 49.752 145.908 ; 
        RECT 49.216 141.534 49.32 145.908 ; 
        RECT 48.784 141.534 48.888 145.908 ; 
        RECT 48.352 141.534 48.456 145.908 ; 
        RECT 47.92 141.534 48.024 145.908 ; 
        RECT 47.488 141.534 47.592 145.908 ; 
        RECT 47.056 141.534 47.16 145.908 ; 
        RECT 46.624 141.534 46.728 145.908 ; 
        RECT 46.192 141.534 46.296 145.908 ; 
        RECT 45.76 141.534 45.864 145.908 ; 
        RECT 45.328 141.534 45.432 145.908 ; 
        RECT 44.896 141.534 45 145.908 ; 
        RECT 44.464 141.534 44.568 145.908 ; 
        RECT 44.032 141.534 44.136 145.908 ; 
        RECT 43.6 141.534 43.704 145.908 ; 
        RECT 43.168 141.534 43.272 145.908 ; 
        RECT 42.736 141.534 42.84 145.908 ; 
        RECT 42.304 141.534 42.408 145.908 ; 
        RECT 41.872 141.534 41.976 145.908 ; 
        RECT 41.44 141.534 41.544 145.908 ; 
        RECT 41.008 141.534 41.112 145.908 ; 
        RECT 40.576 141.534 40.68 145.908 ; 
        RECT 40.144 141.534 40.248 145.908 ; 
        RECT 39.712 141.534 39.816 145.908 ; 
        RECT 39.28 141.534 39.384 145.908 ; 
        RECT 38.848 141.534 38.952 145.908 ; 
        RECT 38.416 141.534 38.52 145.908 ; 
        RECT 37.984 141.534 38.088 145.908 ; 
        RECT 37.552 141.534 37.656 145.908 ; 
        RECT 36.7 141.534 37.008 145.908 ; 
        RECT 29.128 141.534 29.436 145.908 ; 
        RECT 28.48 141.534 28.584 145.908 ; 
        RECT 28.048 141.534 28.152 145.908 ; 
        RECT 27.616 141.534 27.72 145.908 ; 
        RECT 27.184 141.534 27.288 145.908 ; 
        RECT 26.752 141.534 26.856 145.908 ; 
        RECT 26.32 141.534 26.424 145.908 ; 
        RECT 25.888 141.534 25.992 145.908 ; 
        RECT 25.456 141.534 25.56 145.908 ; 
        RECT 25.024 141.534 25.128 145.908 ; 
        RECT 24.592 141.534 24.696 145.908 ; 
        RECT 24.16 141.534 24.264 145.908 ; 
        RECT 23.728 141.534 23.832 145.908 ; 
        RECT 23.296 141.534 23.4 145.908 ; 
        RECT 22.864 141.534 22.968 145.908 ; 
        RECT 22.432 141.534 22.536 145.908 ; 
        RECT 22 141.534 22.104 145.908 ; 
        RECT 21.568 141.534 21.672 145.908 ; 
        RECT 21.136 141.534 21.24 145.908 ; 
        RECT 20.704 141.534 20.808 145.908 ; 
        RECT 20.272 141.534 20.376 145.908 ; 
        RECT 19.84 141.534 19.944 145.908 ; 
        RECT 19.408 141.534 19.512 145.908 ; 
        RECT 18.976 141.534 19.08 145.908 ; 
        RECT 18.544 141.534 18.648 145.908 ; 
        RECT 18.112 141.534 18.216 145.908 ; 
        RECT 17.68 141.534 17.784 145.908 ; 
        RECT 17.248 141.534 17.352 145.908 ; 
        RECT 16.816 141.534 16.92 145.908 ; 
        RECT 16.384 141.534 16.488 145.908 ; 
        RECT 15.952 141.534 16.056 145.908 ; 
        RECT 15.52 141.534 15.624 145.908 ; 
        RECT 15.088 141.534 15.192 145.908 ; 
        RECT 14.656 141.534 14.76 145.908 ; 
        RECT 14.224 141.534 14.328 145.908 ; 
        RECT 13.792 141.534 13.896 145.908 ; 
        RECT 13.36 141.534 13.464 145.908 ; 
        RECT 12.928 141.534 13.032 145.908 ; 
        RECT 12.496 141.534 12.6 145.908 ; 
        RECT 12.064 141.534 12.168 145.908 ; 
        RECT 11.632 141.534 11.736 145.908 ; 
        RECT 11.2 141.534 11.304 145.908 ; 
        RECT 10.768 141.534 10.872 145.908 ; 
        RECT 10.336 141.534 10.44 145.908 ; 
        RECT 9.904 141.534 10.008 145.908 ; 
        RECT 9.472 141.534 9.576 145.908 ; 
        RECT 9.04 141.534 9.144 145.908 ; 
        RECT 8.608 141.534 8.712 145.908 ; 
        RECT 8.176 141.534 8.28 145.908 ; 
        RECT 7.744 141.534 7.848 145.908 ; 
        RECT 7.312 141.534 7.416 145.908 ; 
        RECT 6.88 141.534 6.984 145.908 ; 
        RECT 6.448 141.534 6.552 145.908 ; 
        RECT 6.016 141.534 6.12 145.908 ; 
        RECT 5.584 141.534 5.688 145.908 ; 
        RECT 5.152 141.534 5.256 145.908 ; 
        RECT 4.72 141.534 4.824 145.908 ; 
        RECT 4.288 141.534 4.392 145.908 ; 
        RECT 3.856 141.534 3.96 145.908 ; 
        RECT 3.424 141.534 3.528 145.908 ; 
        RECT 2.992 141.534 3.096 145.908 ; 
        RECT 2.56 141.534 2.664 145.908 ; 
        RECT 2.128 141.534 2.232 145.908 ; 
        RECT 1.696 141.534 1.8 145.908 ; 
        RECT 1.264 141.534 1.368 145.908 ; 
        RECT 0.832 141.534 0.936 145.908 ; 
        RECT 0.02 141.534 0.36 145.908 ; 
        RECT 34.564 145.854 35.076 150.228 ; 
        RECT 34.508 148.516 35.076 149.806 ; 
        RECT 33.916 147.424 34.164 150.228 ; 
        RECT 33.86 148.662 34.164 149.276 ; 
        RECT 33.916 145.854 34.02 150.228 ; 
        RECT 33.916 146.338 34.076 147.296 ; 
        RECT 33.916 145.854 34.164 146.21 ; 
        RECT 32.728 147.656 33.552 150.228 ; 
        RECT 33.448 145.854 33.552 150.228 ; 
        RECT 32.728 148.764 33.608 149.796 ; 
        RECT 32.728 145.854 33.12 150.228 ; 
        RECT 31.06 145.854 31.392 150.228 ; 
        RECT 31.06 146.208 31.448 149.95 ; 
        RECT 65.776 145.854 66.116 150.228 ; 
        RECT 65.2 145.854 65.304 150.228 ; 
        RECT 64.768 145.854 64.872 150.228 ; 
        RECT 64.336 145.854 64.44 150.228 ; 
        RECT 63.904 145.854 64.008 150.228 ; 
        RECT 63.472 145.854 63.576 150.228 ; 
        RECT 63.04 145.854 63.144 150.228 ; 
        RECT 62.608 145.854 62.712 150.228 ; 
        RECT 62.176 145.854 62.28 150.228 ; 
        RECT 61.744 145.854 61.848 150.228 ; 
        RECT 61.312 145.854 61.416 150.228 ; 
        RECT 60.88 145.854 60.984 150.228 ; 
        RECT 60.448 145.854 60.552 150.228 ; 
        RECT 60.016 145.854 60.12 150.228 ; 
        RECT 59.584 145.854 59.688 150.228 ; 
        RECT 59.152 145.854 59.256 150.228 ; 
        RECT 58.72 145.854 58.824 150.228 ; 
        RECT 58.288 145.854 58.392 150.228 ; 
        RECT 57.856 145.854 57.96 150.228 ; 
        RECT 57.424 145.854 57.528 150.228 ; 
        RECT 56.992 145.854 57.096 150.228 ; 
        RECT 56.56 145.854 56.664 150.228 ; 
        RECT 56.128 145.854 56.232 150.228 ; 
        RECT 55.696 145.854 55.8 150.228 ; 
        RECT 55.264 145.854 55.368 150.228 ; 
        RECT 54.832 145.854 54.936 150.228 ; 
        RECT 54.4 145.854 54.504 150.228 ; 
        RECT 53.968 145.854 54.072 150.228 ; 
        RECT 53.536 145.854 53.64 150.228 ; 
        RECT 53.104 145.854 53.208 150.228 ; 
        RECT 52.672 145.854 52.776 150.228 ; 
        RECT 52.24 145.854 52.344 150.228 ; 
        RECT 51.808 145.854 51.912 150.228 ; 
        RECT 51.376 145.854 51.48 150.228 ; 
        RECT 50.944 145.854 51.048 150.228 ; 
        RECT 50.512 145.854 50.616 150.228 ; 
        RECT 50.08 145.854 50.184 150.228 ; 
        RECT 49.648 145.854 49.752 150.228 ; 
        RECT 49.216 145.854 49.32 150.228 ; 
        RECT 48.784 145.854 48.888 150.228 ; 
        RECT 48.352 145.854 48.456 150.228 ; 
        RECT 47.92 145.854 48.024 150.228 ; 
        RECT 47.488 145.854 47.592 150.228 ; 
        RECT 47.056 145.854 47.16 150.228 ; 
        RECT 46.624 145.854 46.728 150.228 ; 
        RECT 46.192 145.854 46.296 150.228 ; 
        RECT 45.76 145.854 45.864 150.228 ; 
        RECT 45.328 145.854 45.432 150.228 ; 
        RECT 44.896 145.854 45 150.228 ; 
        RECT 44.464 145.854 44.568 150.228 ; 
        RECT 44.032 145.854 44.136 150.228 ; 
        RECT 43.6 145.854 43.704 150.228 ; 
        RECT 43.168 145.854 43.272 150.228 ; 
        RECT 42.736 145.854 42.84 150.228 ; 
        RECT 42.304 145.854 42.408 150.228 ; 
        RECT 41.872 145.854 41.976 150.228 ; 
        RECT 41.44 145.854 41.544 150.228 ; 
        RECT 41.008 145.854 41.112 150.228 ; 
        RECT 40.576 145.854 40.68 150.228 ; 
        RECT 40.144 145.854 40.248 150.228 ; 
        RECT 39.712 145.854 39.816 150.228 ; 
        RECT 39.28 145.854 39.384 150.228 ; 
        RECT 38.848 145.854 38.952 150.228 ; 
        RECT 38.416 145.854 38.52 150.228 ; 
        RECT 37.984 145.854 38.088 150.228 ; 
        RECT 37.552 145.854 37.656 150.228 ; 
        RECT 36.7 145.854 37.008 150.228 ; 
        RECT 29.128 145.854 29.436 150.228 ; 
        RECT 28.48 145.854 28.584 150.228 ; 
        RECT 28.048 145.854 28.152 150.228 ; 
        RECT 27.616 145.854 27.72 150.228 ; 
        RECT 27.184 145.854 27.288 150.228 ; 
        RECT 26.752 145.854 26.856 150.228 ; 
        RECT 26.32 145.854 26.424 150.228 ; 
        RECT 25.888 145.854 25.992 150.228 ; 
        RECT 25.456 145.854 25.56 150.228 ; 
        RECT 25.024 145.854 25.128 150.228 ; 
        RECT 24.592 145.854 24.696 150.228 ; 
        RECT 24.16 145.854 24.264 150.228 ; 
        RECT 23.728 145.854 23.832 150.228 ; 
        RECT 23.296 145.854 23.4 150.228 ; 
        RECT 22.864 145.854 22.968 150.228 ; 
        RECT 22.432 145.854 22.536 150.228 ; 
        RECT 22 145.854 22.104 150.228 ; 
        RECT 21.568 145.854 21.672 150.228 ; 
        RECT 21.136 145.854 21.24 150.228 ; 
        RECT 20.704 145.854 20.808 150.228 ; 
        RECT 20.272 145.854 20.376 150.228 ; 
        RECT 19.84 145.854 19.944 150.228 ; 
        RECT 19.408 145.854 19.512 150.228 ; 
        RECT 18.976 145.854 19.08 150.228 ; 
        RECT 18.544 145.854 18.648 150.228 ; 
        RECT 18.112 145.854 18.216 150.228 ; 
        RECT 17.68 145.854 17.784 150.228 ; 
        RECT 17.248 145.854 17.352 150.228 ; 
        RECT 16.816 145.854 16.92 150.228 ; 
        RECT 16.384 145.854 16.488 150.228 ; 
        RECT 15.952 145.854 16.056 150.228 ; 
        RECT 15.52 145.854 15.624 150.228 ; 
        RECT 15.088 145.854 15.192 150.228 ; 
        RECT 14.656 145.854 14.76 150.228 ; 
        RECT 14.224 145.854 14.328 150.228 ; 
        RECT 13.792 145.854 13.896 150.228 ; 
        RECT 13.36 145.854 13.464 150.228 ; 
        RECT 12.928 145.854 13.032 150.228 ; 
        RECT 12.496 145.854 12.6 150.228 ; 
        RECT 12.064 145.854 12.168 150.228 ; 
        RECT 11.632 145.854 11.736 150.228 ; 
        RECT 11.2 145.854 11.304 150.228 ; 
        RECT 10.768 145.854 10.872 150.228 ; 
        RECT 10.336 145.854 10.44 150.228 ; 
        RECT 9.904 145.854 10.008 150.228 ; 
        RECT 9.472 145.854 9.576 150.228 ; 
        RECT 9.04 145.854 9.144 150.228 ; 
        RECT 8.608 145.854 8.712 150.228 ; 
        RECT 8.176 145.854 8.28 150.228 ; 
        RECT 7.744 145.854 7.848 150.228 ; 
        RECT 7.312 145.854 7.416 150.228 ; 
        RECT 6.88 145.854 6.984 150.228 ; 
        RECT 6.448 145.854 6.552 150.228 ; 
        RECT 6.016 145.854 6.12 150.228 ; 
        RECT 5.584 145.854 5.688 150.228 ; 
        RECT 5.152 145.854 5.256 150.228 ; 
        RECT 4.72 145.854 4.824 150.228 ; 
        RECT 4.288 145.854 4.392 150.228 ; 
        RECT 3.856 145.854 3.96 150.228 ; 
        RECT 3.424 145.854 3.528 150.228 ; 
        RECT 2.992 145.854 3.096 150.228 ; 
        RECT 2.56 145.854 2.664 150.228 ; 
        RECT 2.128 145.854 2.232 150.228 ; 
        RECT 1.696 145.854 1.8 150.228 ; 
        RECT 1.264 145.854 1.368 150.228 ; 
        RECT 0.832 145.854 0.936 150.228 ; 
        RECT 0.02 145.854 0.36 150.228 ; 
        RECT 34.564 150.174 35.076 154.548 ; 
        RECT 34.508 152.836 35.076 154.126 ; 
        RECT 33.916 151.744 34.164 154.548 ; 
        RECT 33.86 152.982 34.164 153.596 ; 
        RECT 33.916 150.174 34.02 154.548 ; 
        RECT 33.916 150.658 34.076 151.616 ; 
        RECT 33.916 150.174 34.164 150.53 ; 
        RECT 32.728 151.976 33.552 154.548 ; 
        RECT 33.448 150.174 33.552 154.548 ; 
        RECT 32.728 153.084 33.608 154.116 ; 
        RECT 32.728 150.174 33.12 154.548 ; 
        RECT 31.06 150.174 31.392 154.548 ; 
        RECT 31.06 150.528 31.448 154.27 ; 
        RECT 65.776 150.174 66.116 154.548 ; 
        RECT 65.2 150.174 65.304 154.548 ; 
        RECT 64.768 150.174 64.872 154.548 ; 
        RECT 64.336 150.174 64.44 154.548 ; 
        RECT 63.904 150.174 64.008 154.548 ; 
        RECT 63.472 150.174 63.576 154.548 ; 
        RECT 63.04 150.174 63.144 154.548 ; 
        RECT 62.608 150.174 62.712 154.548 ; 
        RECT 62.176 150.174 62.28 154.548 ; 
        RECT 61.744 150.174 61.848 154.548 ; 
        RECT 61.312 150.174 61.416 154.548 ; 
        RECT 60.88 150.174 60.984 154.548 ; 
        RECT 60.448 150.174 60.552 154.548 ; 
        RECT 60.016 150.174 60.12 154.548 ; 
        RECT 59.584 150.174 59.688 154.548 ; 
        RECT 59.152 150.174 59.256 154.548 ; 
        RECT 58.72 150.174 58.824 154.548 ; 
        RECT 58.288 150.174 58.392 154.548 ; 
        RECT 57.856 150.174 57.96 154.548 ; 
        RECT 57.424 150.174 57.528 154.548 ; 
        RECT 56.992 150.174 57.096 154.548 ; 
        RECT 56.56 150.174 56.664 154.548 ; 
        RECT 56.128 150.174 56.232 154.548 ; 
        RECT 55.696 150.174 55.8 154.548 ; 
        RECT 55.264 150.174 55.368 154.548 ; 
        RECT 54.832 150.174 54.936 154.548 ; 
        RECT 54.4 150.174 54.504 154.548 ; 
        RECT 53.968 150.174 54.072 154.548 ; 
        RECT 53.536 150.174 53.64 154.548 ; 
        RECT 53.104 150.174 53.208 154.548 ; 
        RECT 52.672 150.174 52.776 154.548 ; 
        RECT 52.24 150.174 52.344 154.548 ; 
        RECT 51.808 150.174 51.912 154.548 ; 
        RECT 51.376 150.174 51.48 154.548 ; 
        RECT 50.944 150.174 51.048 154.548 ; 
        RECT 50.512 150.174 50.616 154.548 ; 
        RECT 50.08 150.174 50.184 154.548 ; 
        RECT 49.648 150.174 49.752 154.548 ; 
        RECT 49.216 150.174 49.32 154.548 ; 
        RECT 48.784 150.174 48.888 154.548 ; 
        RECT 48.352 150.174 48.456 154.548 ; 
        RECT 47.92 150.174 48.024 154.548 ; 
        RECT 47.488 150.174 47.592 154.548 ; 
        RECT 47.056 150.174 47.16 154.548 ; 
        RECT 46.624 150.174 46.728 154.548 ; 
        RECT 46.192 150.174 46.296 154.548 ; 
        RECT 45.76 150.174 45.864 154.548 ; 
        RECT 45.328 150.174 45.432 154.548 ; 
        RECT 44.896 150.174 45 154.548 ; 
        RECT 44.464 150.174 44.568 154.548 ; 
        RECT 44.032 150.174 44.136 154.548 ; 
        RECT 43.6 150.174 43.704 154.548 ; 
        RECT 43.168 150.174 43.272 154.548 ; 
        RECT 42.736 150.174 42.84 154.548 ; 
        RECT 42.304 150.174 42.408 154.548 ; 
        RECT 41.872 150.174 41.976 154.548 ; 
        RECT 41.44 150.174 41.544 154.548 ; 
        RECT 41.008 150.174 41.112 154.548 ; 
        RECT 40.576 150.174 40.68 154.548 ; 
        RECT 40.144 150.174 40.248 154.548 ; 
        RECT 39.712 150.174 39.816 154.548 ; 
        RECT 39.28 150.174 39.384 154.548 ; 
        RECT 38.848 150.174 38.952 154.548 ; 
        RECT 38.416 150.174 38.52 154.548 ; 
        RECT 37.984 150.174 38.088 154.548 ; 
        RECT 37.552 150.174 37.656 154.548 ; 
        RECT 36.7 150.174 37.008 154.548 ; 
        RECT 29.128 150.174 29.436 154.548 ; 
        RECT 28.48 150.174 28.584 154.548 ; 
        RECT 28.048 150.174 28.152 154.548 ; 
        RECT 27.616 150.174 27.72 154.548 ; 
        RECT 27.184 150.174 27.288 154.548 ; 
        RECT 26.752 150.174 26.856 154.548 ; 
        RECT 26.32 150.174 26.424 154.548 ; 
        RECT 25.888 150.174 25.992 154.548 ; 
        RECT 25.456 150.174 25.56 154.548 ; 
        RECT 25.024 150.174 25.128 154.548 ; 
        RECT 24.592 150.174 24.696 154.548 ; 
        RECT 24.16 150.174 24.264 154.548 ; 
        RECT 23.728 150.174 23.832 154.548 ; 
        RECT 23.296 150.174 23.4 154.548 ; 
        RECT 22.864 150.174 22.968 154.548 ; 
        RECT 22.432 150.174 22.536 154.548 ; 
        RECT 22 150.174 22.104 154.548 ; 
        RECT 21.568 150.174 21.672 154.548 ; 
        RECT 21.136 150.174 21.24 154.548 ; 
        RECT 20.704 150.174 20.808 154.548 ; 
        RECT 20.272 150.174 20.376 154.548 ; 
        RECT 19.84 150.174 19.944 154.548 ; 
        RECT 19.408 150.174 19.512 154.548 ; 
        RECT 18.976 150.174 19.08 154.548 ; 
        RECT 18.544 150.174 18.648 154.548 ; 
        RECT 18.112 150.174 18.216 154.548 ; 
        RECT 17.68 150.174 17.784 154.548 ; 
        RECT 17.248 150.174 17.352 154.548 ; 
        RECT 16.816 150.174 16.92 154.548 ; 
        RECT 16.384 150.174 16.488 154.548 ; 
        RECT 15.952 150.174 16.056 154.548 ; 
        RECT 15.52 150.174 15.624 154.548 ; 
        RECT 15.088 150.174 15.192 154.548 ; 
        RECT 14.656 150.174 14.76 154.548 ; 
        RECT 14.224 150.174 14.328 154.548 ; 
        RECT 13.792 150.174 13.896 154.548 ; 
        RECT 13.36 150.174 13.464 154.548 ; 
        RECT 12.928 150.174 13.032 154.548 ; 
        RECT 12.496 150.174 12.6 154.548 ; 
        RECT 12.064 150.174 12.168 154.548 ; 
        RECT 11.632 150.174 11.736 154.548 ; 
        RECT 11.2 150.174 11.304 154.548 ; 
        RECT 10.768 150.174 10.872 154.548 ; 
        RECT 10.336 150.174 10.44 154.548 ; 
        RECT 9.904 150.174 10.008 154.548 ; 
        RECT 9.472 150.174 9.576 154.548 ; 
        RECT 9.04 150.174 9.144 154.548 ; 
        RECT 8.608 150.174 8.712 154.548 ; 
        RECT 8.176 150.174 8.28 154.548 ; 
        RECT 7.744 150.174 7.848 154.548 ; 
        RECT 7.312 150.174 7.416 154.548 ; 
        RECT 6.88 150.174 6.984 154.548 ; 
        RECT 6.448 150.174 6.552 154.548 ; 
        RECT 6.016 150.174 6.12 154.548 ; 
        RECT 5.584 150.174 5.688 154.548 ; 
        RECT 5.152 150.174 5.256 154.548 ; 
        RECT 4.72 150.174 4.824 154.548 ; 
        RECT 4.288 150.174 4.392 154.548 ; 
        RECT 3.856 150.174 3.96 154.548 ; 
        RECT 3.424 150.174 3.528 154.548 ; 
        RECT 2.992 150.174 3.096 154.548 ; 
        RECT 2.56 150.174 2.664 154.548 ; 
        RECT 2.128 150.174 2.232 154.548 ; 
        RECT 1.696 150.174 1.8 154.548 ; 
        RECT 1.264 150.174 1.368 154.548 ; 
        RECT 0.832 150.174 0.936 154.548 ; 
        RECT 0.02 150.174 0.36 154.548 ; 
        RECT 34.564 154.494 35.076 158.868 ; 
        RECT 34.508 157.156 35.076 158.446 ; 
        RECT 33.916 156.064 34.164 158.868 ; 
        RECT 33.86 157.302 34.164 157.916 ; 
        RECT 33.916 154.494 34.02 158.868 ; 
        RECT 33.916 154.978 34.076 155.936 ; 
        RECT 33.916 154.494 34.164 154.85 ; 
        RECT 32.728 156.296 33.552 158.868 ; 
        RECT 33.448 154.494 33.552 158.868 ; 
        RECT 32.728 157.404 33.608 158.436 ; 
        RECT 32.728 154.494 33.12 158.868 ; 
        RECT 31.06 154.494 31.392 158.868 ; 
        RECT 31.06 154.848 31.448 158.59 ; 
        RECT 65.776 154.494 66.116 158.868 ; 
        RECT 65.2 154.494 65.304 158.868 ; 
        RECT 64.768 154.494 64.872 158.868 ; 
        RECT 64.336 154.494 64.44 158.868 ; 
        RECT 63.904 154.494 64.008 158.868 ; 
        RECT 63.472 154.494 63.576 158.868 ; 
        RECT 63.04 154.494 63.144 158.868 ; 
        RECT 62.608 154.494 62.712 158.868 ; 
        RECT 62.176 154.494 62.28 158.868 ; 
        RECT 61.744 154.494 61.848 158.868 ; 
        RECT 61.312 154.494 61.416 158.868 ; 
        RECT 60.88 154.494 60.984 158.868 ; 
        RECT 60.448 154.494 60.552 158.868 ; 
        RECT 60.016 154.494 60.12 158.868 ; 
        RECT 59.584 154.494 59.688 158.868 ; 
        RECT 59.152 154.494 59.256 158.868 ; 
        RECT 58.72 154.494 58.824 158.868 ; 
        RECT 58.288 154.494 58.392 158.868 ; 
        RECT 57.856 154.494 57.96 158.868 ; 
        RECT 57.424 154.494 57.528 158.868 ; 
        RECT 56.992 154.494 57.096 158.868 ; 
        RECT 56.56 154.494 56.664 158.868 ; 
        RECT 56.128 154.494 56.232 158.868 ; 
        RECT 55.696 154.494 55.8 158.868 ; 
        RECT 55.264 154.494 55.368 158.868 ; 
        RECT 54.832 154.494 54.936 158.868 ; 
        RECT 54.4 154.494 54.504 158.868 ; 
        RECT 53.968 154.494 54.072 158.868 ; 
        RECT 53.536 154.494 53.64 158.868 ; 
        RECT 53.104 154.494 53.208 158.868 ; 
        RECT 52.672 154.494 52.776 158.868 ; 
        RECT 52.24 154.494 52.344 158.868 ; 
        RECT 51.808 154.494 51.912 158.868 ; 
        RECT 51.376 154.494 51.48 158.868 ; 
        RECT 50.944 154.494 51.048 158.868 ; 
        RECT 50.512 154.494 50.616 158.868 ; 
        RECT 50.08 154.494 50.184 158.868 ; 
        RECT 49.648 154.494 49.752 158.868 ; 
        RECT 49.216 154.494 49.32 158.868 ; 
        RECT 48.784 154.494 48.888 158.868 ; 
        RECT 48.352 154.494 48.456 158.868 ; 
        RECT 47.92 154.494 48.024 158.868 ; 
        RECT 47.488 154.494 47.592 158.868 ; 
        RECT 47.056 154.494 47.16 158.868 ; 
        RECT 46.624 154.494 46.728 158.868 ; 
        RECT 46.192 154.494 46.296 158.868 ; 
        RECT 45.76 154.494 45.864 158.868 ; 
        RECT 45.328 154.494 45.432 158.868 ; 
        RECT 44.896 154.494 45 158.868 ; 
        RECT 44.464 154.494 44.568 158.868 ; 
        RECT 44.032 154.494 44.136 158.868 ; 
        RECT 43.6 154.494 43.704 158.868 ; 
        RECT 43.168 154.494 43.272 158.868 ; 
        RECT 42.736 154.494 42.84 158.868 ; 
        RECT 42.304 154.494 42.408 158.868 ; 
        RECT 41.872 154.494 41.976 158.868 ; 
        RECT 41.44 154.494 41.544 158.868 ; 
        RECT 41.008 154.494 41.112 158.868 ; 
        RECT 40.576 154.494 40.68 158.868 ; 
        RECT 40.144 154.494 40.248 158.868 ; 
        RECT 39.712 154.494 39.816 158.868 ; 
        RECT 39.28 154.494 39.384 158.868 ; 
        RECT 38.848 154.494 38.952 158.868 ; 
        RECT 38.416 154.494 38.52 158.868 ; 
        RECT 37.984 154.494 38.088 158.868 ; 
        RECT 37.552 154.494 37.656 158.868 ; 
        RECT 36.7 154.494 37.008 158.868 ; 
        RECT 29.128 154.494 29.436 158.868 ; 
        RECT 28.48 154.494 28.584 158.868 ; 
        RECT 28.048 154.494 28.152 158.868 ; 
        RECT 27.616 154.494 27.72 158.868 ; 
        RECT 27.184 154.494 27.288 158.868 ; 
        RECT 26.752 154.494 26.856 158.868 ; 
        RECT 26.32 154.494 26.424 158.868 ; 
        RECT 25.888 154.494 25.992 158.868 ; 
        RECT 25.456 154.494 25.56 158.868 ; 
        RECT 25.024 154.494 25.128 158.868 ; 
        RECT 24.592 154.494 24.696 158.868 ; 
        RECT 24.16 154.494 24.264 158.868 ; 
        RECT 23.728 154.494 23.832 158.868 ; 
        RECT 23.296 154.494 23.4 158.868 ; 
        RECT 22.864 154.494 22.968 158.868 ; 
        RECT 22.432 154.494 22.536 158.868 ; 
        RECT 22 154.494 22.104 158.868 ; 
        RECT 21.568 154.494 21.672 158.868 ; 
        RECT 21.136 154.494 21.24 158.868 ; 
        RECT 20.704 154.494 20.808 158.868 ; 
        RECT 20.272 154.494 20.376 158.868 ; 
        RECT 19.84 154.494 19.944 158.868 ; 
        RECT 19.408 154.494 19.512 158.868 ; 
        RECT 18.976 154.494 19.08 158.868 ; 
        RECT 18.544 154.494 18.648 158.868 ; 
        RECT 18.112 154.494 18.216 158.868 ; 
        RECT 17.68 154.494 17.784 158.868 ; 
        RECT 17.248 154.494 17.352 158.868 ; 
        RECT 16.816 154.494 16.92 158.868 ; 
        RECT 16.384 154.494 16.488 158.868 ; 
        RECT 15.952 154.494 16.056 158.868 ; 
        RECT 15.52 154.494 15.624 158.868 ; 
        RECT 15.088 154.494 15.192 158.868 ; 
        RECT 14.656 154.494 14.76 158.868 ; 
        RECT 14.224 154.494 14.328 158.868 ; 
        RECT 13.792 154.494 13.896 158.868 ; 
        RECT 13.36 154.494 13.464 158.868 ; 
        RECT 12.928 154.494 13.032 158.868 ; 
        RECT 12.496 154.494 12.6 158.868 ; 
        RECT 12.064 154.494 12.168 158.868 ; 
        RECT 11.632 154.494 11.736 158.868 ; 
        RECT 11.2 154.494 11.304 158.868 ; 
        RECT 10.768 154.494 10.872 158.868 ; 
        RECT 10.336 154.494 10.44 158.868 ; 
        RECT 9.904 154.494 10.008 158.868 ; 
        RECT 9.472 154.494 9.576 158.868 ; 
        RECT 9.04 154.494 9.144 158.868 ; 
        RECT 8.608 154.494 8.712 158.868 ; 
        RECT 8.176 154.494 8.28 158.868 ; 
        RECT 7.744 154.494 7.848 158.868 ; 
        RECT 7.312 154.494 7.416 158.868 ; 
        RECT 6.88 154.494 6.984 158.868 ; 
        RECT 6.448 154.494 6.552 158.868 ; 
        RECT 6.016 154.494 6.12 158.868 ; 
        RECT 5.584 154.494 5.688 158.868 ; 
        RECT 5.152 154.494 5.256 158.868 ; 
        RECT 4.72 154.494 4.824 158.868 ; 
        RECT 4.288 154.494 4.392 158.868 ; 
        RECT 3.856 154.494 3.96 158.868 ; 
        RECT 3.424 154.494 3.528 158.868 ; 
        RECT 2.992 154.494 3.096 158.868 ; 
        RECT 2.56 154.494 2.664 158.868 ; 
        RECT 2.128 154.494 2.232 158.868 ; 
        RECT 1.696 154.494 1.8 158.868 ; 
        RECT 1.264 154.494 1.368 158.868 ; 
        RECT 0.832 154.494 0.936 158.868 ; 
        RECT 0.02 154.494 0.36 158.868 ; 
        RECT 34.564 158.814 35.076 163.188 ; 
        RECT 34.508 161.476 35.076 162.766 ; 
        RECT 33.916 160.384 34.164 163.188 ; 
        RECT 33.86 161.622 34.164 162.236 ; 
        RECT 33.916 158.814 34.02 163.188 ; 
        RECT 33.916 159.298 34.076 160.256 ; 
        RECT 33.916 158.814 34.164 159.17 ; 
        RECT 32.728 160.616 33.552 163.188 ; 
        RECT 33.448 158.814 33.552 163.188 ; 
        RECT 32.728 161.724 33.608 162.756 ; 
        RECT 32.728 158.814 33.12 163.188 ; 
        RECT 31.06 158.814 31.392 163.188 ; 
        RECT 31.06 159.168 31.448 162.91 ; 
        RECT 65.776 158.814 66.116 163.188 ; 
        RECT 65.2 158.814 65.304 163.188 ; 
        RECT 64.768 158.814 64.872 163.188 ; 
        RECT 64.336 158.814 64.44 163.188 ; 
        RECT 63.904 158.814 64.008 163.188 ; 
        RECT 63.472 158.814 63.576 163.188 ; 
        RECT 63.04 158.814 63.144 163.188 ; 
        RECT 62.608 158.814 62.712 163.188 ; 
        RECT 62.176 158.814 62.28 163.188 ; 
        RECT 61.744 158.814 61.848 163.188 ; 
        RECT 61.312 158.814 61.416 163.188 ; 
        RECT 60.88 158.814 60.984 163.188 ; 
        RECT 60.448 158.814 60.552 163.188 ; 
        RECT 60.016 158.814 60.12 163.188 ; 
        RECT 59.584 158.814 59.688 163.188 ; 
        RECT 59.152 158.814 59.256 163.188 ; 
        RECT 58.72 158.814 58.824 163.188 ; 
        RECT 58.288 158.814 58.392 163.188 ; 
        RECT 57.856 158.814 57.96 163.188 ; 
        RECT 57.424 158.814 57.528 163.188 ; 
        RECT 56.992 158.814 57.096 163.188 ; 
        RECT 56.56 158.814 56.664 163.188 ; 
        RECT 56.128 158.814 56.232 163.188 ; 
        RECT 55.696 158.814 55.8 163.188 ; 
        RECT 55.264 158.814 55.368 163.188 ; 
        RECT 54.832 158.814 54.936 163.188 ; 
        RECT 54.4 158.814 54.504 163.188 ; 
        RECT 53.968 158.814 54.072 163.188 ; 
        RECT 53.536 158.814 53.64 163.188 ; 
        RECT 53.104 158.814 53.208 163.188 ; 
        RECT 52.672 158.814 52.776 163.188 ; 
        RECT 52.24 158.814 52.344 163.188 ; 
        RECT 51.808 158.814 51.912 163.188 ; 
        RECT 51.376 158.814 51.48 163.188 ; 
        RECT 50.944 158.814 51.048 163.188 ; 
        RECT 50.512 158.814 50.616 163.188 ; 
        RECT 50.08 158.814 50.184 163.188 ; 
        RECT 49.648 158.814 49.752 163.188 ; 
        RECT 49.216 158.814 49.32 163.188 ; 
        RECT 48.784 158.814 48.888 163.188 ; 
        RECT 48.352 158.814 48.456 163.188 ; 
        RECT 47.92 158.814 48.024 163.188 ; 
        RECT 47.488 158.814 47.592 163.188 ; 
        RECT 47.056 158.814 47.16 163.188 ; 
        RECT 46.624 158.814 46.728 163.188 ; 
        RECT 46.192 158.814 46.296 163.188 ; 
        RECT 45.76 158.814 45.864 163.188 ; 
        RECT 45.328 158.814 45.432 163.188 ; 
        RECT 44.896 158.814 45 163.188 ; 
        RECT 44.464 158.814 44.568 163.188 ; 
        RECT 44.032 158.814 44.136 163.188 ; 
        RECT 43.6 158.814 43.704 163.188 ; 
        RECT 43.168 158.814 43.272 163.188 ; 
        RECT 42.736 158.814 42.84 163.188 ; 
        RECT 42.304 158.814 42.408 163.188 ; 
        RECT 41.872 158.814 41.976 163.188 ; 
        RECT 41.44 158.814 41.544 163.188 ; 
        RECT 41.008 158.814 41.112 163.188 ; 
        RECT 40.576 158.814 40.68 163.188 ; 
        RECT 40.144 158.814 40.248 163.188 ; 
        RECT 39.712 158.814 39.816 163.188 ; 
        RECT 39.28 158.814 39.384 163.188 ; 
        RECT 38.848 158.814 38.952 163.188 ; 
        RECT 38.416 158.814 38.52 163.188 ; 
        RECT 37.984 158.814 38.088 163.188 ; 
        RECT 37.552 158.814 37.656 163.188 ; 
        RECT 36.7 158.814 37.008 163.188 ; 
        RECT 29.128 158.814 29.436 163.188 ; 
        RECT 28.48 158.814 28.584 163.188 ; 
        RECT 28.048 158.814 28.152 163.188 ; 
        RECT 27.616 158.814 27.72 163.188 ; 
        RECT 27.184 158.814 27.288 163.188 ; 
        RECT 26.752 158.814 26.856 163.188 ; 
        RECT 26.32 158.814 26.424 163.188 ; 
        RECT 25.888 158.814 25.992 163.188 ; 
        RECT 25.456 158.814 25.56 163.188 ; 
        RECT 25.024 158.814 25.128 163.188 ; 
        RECT 24.592 158.814 24.696 163.188 ; 
        RECT 24.16 158.814 24.264 163.188 ; 
        RECT 23.728 158.814 23.832 163.188 ; 
        RECT 23.296 158.814 23.4 163.188 ; 
        RECT 22.864 158.814 22.968 163.188 ; 
        RECT 22.432 158.814 22.536 163.188 ; 
        RECT 22 158.814 22.104 163.188 ; 
        RECT 21.568 158.814 21.672 163.188 ; 
        RECT 21.136 158.814 21.24 163.188 ; 
        RECT 20.704 158.814 20.808 163.188 ; 
        RECT 20.272 158.814 20.376 163.188 ; 
        RECT 19.84 158.814 19.944 163.188 ; 
        RECT 19.408 158.814 19.512 163.188 ; 
        RECT 18.976 158.814 19.08 163.188 ; 
        RECT 18.544 158.814 18.648 163.188 ; 
        RECT 18.112 158.814 18.216 163.188 ; 
        RECT 17.68 158.814 17.784 163.188 ; 
        RECT 17.248 158.814 17.352 163.188 ; 
        RECT 16.816 158.814 16.92 163.188 ; 
        RECT 16.384 158.814 16.488 163.188 ; 
        RECT 15.952 158.814 16.056 163.188 ; 
        RECT 15.52 158.814 15.624 163.188 ; 
        RECT 15.088 158.814 15.192 163.188 ; 
        RECT 14.656 158.814 14.76 163.188 ; 
        RECT 14.224 158.814 14.328 163.188 ; 
        RECT 13.792 158.814 13.896 163.188 ; 
        RECT 13.36 158.814 13.464 163.188 ; 
        RECT 12.928 158.814 13.032 163.188 ; 
        RECT 12.496 158.814 12.6 163.188 ; 
        RECT 12.064 158.814 12.168 163.188 ; 
        RECT 11.632 158.814 11.736 163.188 ; 
        RECT 11.2 158.814 11.304 163.188 ; 
        RECT 10.768 158.814 10.872 163.188 ; 
        RECT 10.336 158.814 10.44 163.188 ; 
        RECT 9.904 158.814 10.008 163.188 ; 
        RECT 9.472 158.814 9.576 163.188 ; 
        RECT 9.04 158.814 9.144 163.188 ; 
        RECT 8.608 158.814 8.712 163.188 ; 
        RECT 8.176 158.814 8.28 163.188 ; 
        RECT 7.744 158.814 7.848 163.188 ; 
        RECT 7.312 158.814 7.416 163.188 ; 
        RECT 6.88 158.814 6.984 163.188 ; 
        RECT 6.448 158.814 6.552 163.188 ; 
        RECT 6.016 158.814 6.12 163.188 ; 
        RECT 5.584 158.814 5.688 163.188 ; 
        RECT 5.152 158.814 5.256 163.188 ; 
        RECT 4.72 158.814 4.824 163.188 ; 
        RECT 4.288 158.814 4.392 163.188 ; 
        RECT 3.856 158.814 3.96 163.188 ; 
        RECT 3.424 158.814 3.528 163.188 ; 
        RECT 2.992 158.814 3.096 163.188 ; 
        RECT 2.56 158.814 2.664 163.188 ; 
        RECT 2.128 158.814 2.232 163.188 ; 
        RECT 1.696 158.814 1.8 163.188 ; 
        RECT 1.264 158.814 1.368 163.188 ; 
        RECT 0.832 158.814 0.936 163.188 ; 
        RECT 0.02 158.814 0.36 163.188 ; 
        RECT 34.564 163.134 35.076 167.508 ; 
        RECT 34.508 165.796 35.076 167.086 ; 
        RECT 33.916 164.704 34.164 167.508 ; 
        RECT 33.86 165.942 34.164 166.556 ; 
        RECT 33.916 163.134 34.02 167.508 ; 
        RECT 33.916 163.618 34.076 164.576 ; 
        RECT 33.916 163.134 34.164 163.49 ; 
        RECT 32.728 164.936 33.552 167.508 ; 
        RECT 33.448 163.134 33.552 167.508 ; 
        RECT 32.728 166.044 33.608 167.076 ; 
        RECT 32.728 163.134 33.12 167.508 ; 
        RECT 31.06 163.134 31.392 167.508 ; 
        RECT 31.06 163.488 31.448 167.23 ; 
        RECT 65.776 163.134 66.116 167.508 ; 
        RECT 65.2 163.134 65.304 167.508 ; 
        RECT 64.768 163.134 64.872 167.508 ; 
        RECT 64.336 163.134 64.44 167.508 ; 
        RECT 63.904 163.134 64.008 167.508 ; 
        RECT 63.472 163.134 63.576 167.508 ; 
        RECT 63.04 163.134 63.144 167.508 ; 
        RECT 62.608 163.134 62.712 167.508 ; 
        RECT 62.176 163.134 62.28 167.508 ; 
        RECT 61.744 163.134 61.848 167.508 ; 
        RECT 61.312 163.134 61.416 167.508 ; 
        RECT 60.88 163.134 60.984 167.508 ; 
        RECT 60.448 163.134 60.552 167.508 ; 
        RECT 60.016 163.134 60.12 167.508 ; 
        RECT 59.584 163.134 59.688 167.508 ; 
        RECT 59.152 163.134 59.256 167.508 ; 
        RECT 58.72 163.134 58.824 167.508 ; 
        RECT 58.288 163.134 58.392 167.508 ; 
        RECT 57.856 163.134 57.96 167.508 ; 
        RECT 57.424 163.134 57.528 167.508 ; 
        RECT 56.992 163.134 57.096 167.508 ; 
        RECT 56.56 163.134 56.664 167.508 ; 
        RECT 56.128 163.134 56.232 167.508 ; 
        RECT 55.696 163.134 55.8 167.508 ; 
        RECT 55.264 163.134 55.368 167.508 ; 
        RECT 54.832 163.134 54.936 167.508 ; 
        RECT 54.4 163.134 54.504 167.508 ; 
        RECT 53.968 163.134 54.072 167.508 ; 
        RECT 53.536 163.134 53.64 167.508 ; 
        RECT 53.104 163.134 53.208 167.508 ; 
        RECT 52.672 163.134 52.776 167.508 ; 
        RECT 52.24 163.134 52.344 167.508 ; 
        RECT 51.808 163.134 51.912 167.508 ; 
        RECT 51.376 163.134 51.48 167.508 ; 
        RECT 50.944 163.134 51.048 167.508 ; 
        RECT 50.512 163.134 50.616 167.508 ; 
        RECT 50.08 163.134 50.184 167.508 ; 
        RECT 49.648 163.134 49.752 167.508 ; 
        RECT 49.216 163.134 49.32 167.508 ; 
        RECT 48.784 163.134 48.888 167.508 ; 
        RECT 48.352 163.134 48.456 167.508 ; 
        RECT 47.92 163.134 48.024 167.508 ; 
        RECT 47.488 163.134 47.592 167.508 ; 
        RECT 47.056 163.134 47.16 167.508 ; 
        RECT 46.624 163.134 46.728 167.508 ; 
        RECT 46.192 163.134 46.296 167.508 ; 
        RECT 45.76 163.134 45.864 167.508 ; 
        RECT 45.328 163.134 45.432 167.508 ; 
        RECT 44.896 163.134 45 167.508 ; 
        RECT 44.464 163.134 44.568 167.508 ; 
        RECT 44.032 163.134 44.136 167.508 ; 
        RECT 43.6 163.134 43.704 167.508 ; 
        RECT 43.168 163.134 43.272 167.508 ; 
        RECT 42.736 163.134 42.84 167.508 ; 
        RECT 42.304 163.134 42.408 167.508 ; 
        RECT 41.872 163.134 41.976 167.508 ; 
        RECT 41.44 163.134 41.544 167.508 ; 
        RECT 41.008 163.134 41.112 167.508 ; 
        RECT 40.576 163.134 40.68 167.508 ; 
        RECT 40.144 163.134 40.248 167.508 ; 
        RECT 39.712 163.134 39.816 167.508 ; 
        RECT 39.28 163.134 39.384 167.508 ; 
        RECT 38.848 163.134 38.952 167.508 ; 
        RECT 38.416 163.134 38.52 167.508 ; 
        RECT 37.984 163.134 38.088 167.508 ; 
        RECT 37.552 163.134 37.656 167.508 ; 
        RECT 36.7 163.134 37.008 167.508 ; 
        RECT 29.128 163.134 29.436 167.508 ; 
        RECT 28.48 163.134 28.584 167.508 ; 
        RECT 28.048 163.134 28.152 167.508 ; 
        RECT 27.616 163.134 27.72 167.508 ; 
        RECT 27.184 163.134 27.288 167.508 ; 
        RECT 26.752 163.134 26.856 167.508 ; 
        RECT 26.32 163.134 26.424 167.508 ; 
        RECT 25.888 163.134 25.992 167.508 ; 
        RECT 25.456 163.134 25.56 167.508 ; 
        RECT 25.024 163.134 25.128 167.508 ; 
        RECT 24.592 163.134 24.696 167.508 ; 
        RECT 24.16 163.134 24.264 167.508 ; 
        RECT 23.728 163.134 23.832 167.508 ; 
        RECT 23.296 163.134 23.4 167.508 ; 
        RECT 22.864 163.134 22.968 167.508 ; 
        RECT 22.432 163.134 22.536 167.508 ; 
        RECT 22 163.134 22.104 167.508 ; 
        RECT 21.568 163.134 21.672 167.508 ; 
        RECT 21.136 163.134 21.24 167.508 ; 
        RECT 20.704 163.134 20.808 167.508 ; 
        RECT 20.272 163.134 20.376 167.508 ; 
        RECT 19.84 163.134 19.944 167.508 ; 
        RECT 19.408 163.134 19.512 167.508 ; 
        RECT 18.976 163.134 19.08 167.508 ; 
        RECT 18.544 163.134 18.648 167.508 ; 
        RECT 18.112 163.134 18.216 167.508 ; 
        RECT 17.68 163.134 17.784 167.508 ; 
        RECT 17.248 163.134 17.352 167.508 ; 
        RECT 16.816 163.134 16.92 167.508 ; 
        RECT 16.384 163.134 16.488 167.508 ; 
        RECT 15.952 163.134 16.056 167.508 ; 
        RECT 15.52 163.134 15.624 167.508 ; 
        RECT 15.088 163.134 15.192 167.508 ; 
        RECT 14.656 163.134 14.76 167.508 ; 
        RECT 14.224 163.134 14.328 167.508 ; 
        RECT 13.792 163.134 13.896 167.508 ; 
        RECT 13.36 163.134 13.464 167.508 ; 
        RECT 12.928 163.134 13.032 167.508 ; 
        RECT 12.496 163.134 12.6 167.508 ; 
        RECT 12.064 163.134 12.168 167.508 ; 
        RECT 11.632 163.134 11.736 167.508 ; 
        RECT 11.2 163.134 11.304 167.508 ; 
        RECT 10.768 163.134 10.872 167.508 ; 
        RECT 10.336 163.134 10.44 167.508 ; 
        RECT 9.904 163.134 10.008 167.508 ; 
        RECT 9.472 163.134 9.576 167.508 ; 
        RECT 9.04 163.134 9.144 167.508 ; 
        RECT 8.608 163.134 8.712 167.508 ; 
        RECT 8.176 163.134 8.28 167.508 ; 
        RECT 7.744 163.134 7.848 167.508 ; 
        RECT 7.312 163.134 7.416 167.508 ; 
        RECT 6.88 163.134 6.984 167.508 ; 
        RECT 6.448 163.134 6.552 167.508 ; 
        RECT 6.016 163.134 6.12 167.508 ; 
        RECT 5.584 163.134 5.688 167.508 ; 
        RECT 5.152 163.134 5.256 167.508 ; 
        RECT 4.72 163.134 4.824 167.508 ; 
        RECT 4.288 163.134 4.392 167.508 ; 
        RECT 3.856 163.134 3.96 167.508 ; 
        RECT 3.424 163.134 3.528 167.508 ; 
        RECT 2.992 163.134 3.096 167.508 ; 
        RECT 2.56 163.134 2.664 167.508 ; 
        RECT 2.128 163.134 2.232 167.508 ; 
        RECT 1.696 163.134 1.8 167.508 ; 
        RECT 1.264 163.134 1.368 167.508 ; 
        RECT 0.832 163.134 0.936 167.508 ; 
        RECT 0.02 163.134 0.36 167.508 ; 
        RECT 34.564 167.454 35.076 171.828 ; 
        RECT 34.508 170.116 35.076 171.406 ; 
        RECT 33.916 169.024 34.164 171.828 ; 
        RECT 33.86 170.262 34.164 170.876 ; 
        RECT 33.916 167.454 34.02 171.828 ; 
        RECT 33.916 167.938 34.076 168.896 ; 
        RECT 33.916 167.454 34.164 167.81 ; 
        RECT 32.728 169.256 33.552 171.828 ; 
        RECT 33.448 167.454 33.552 171.828 ; 
        RECT 32.728 170.364 33.608 171.396 ; 
        RECT 32.728 167.454 33.12 171.828 ; 
        RECT 31.06 167.454 31.392 171.828 ; 
        RECT 31.06 167.808 31.448 171.55 ; 
        RECT 65.776 167.454 66.116 171.828 ; 
        RECT 65.2 167.454 65.304 171.828 ; 
        RECT 64.768 167.454 64.872 171.828 ; 
        RECT 64.336 167.454 64.44 171.828 ; 
        RECT 63.904 167.454 64.008 171.828 ; 
        RECT 63.472 167.454 63.576 171.828 ; 
        RECT 63.04 167.454 63.144 171.828 ; 
        RECT 62.608 167.454 62.712 171.828 ; 
        RECT 62.176 167.454 62.28 171.828 ; 
        RECT 61.744 167.454 61.848 171.828 ; 
        RECT 61.312 167.454 61.416 171.828 ; 
        RECT 60.88 167.454 60.984 171.828 ; 
        RECT 60.448 167.454 60.552 171.828 ; 
        RECT 60.016 167.454 60.12 171.828 ; 
        RECT 59.584 167.454 59.688 171.828 ; 
        RECT 59.152 167.454 59.256 171.828 ; 
        RECT 58.72 167.454 58.824 171.828 ; 
        RECT 58.288 167.454 58.392 171.828 ; 
        RECT 57.856 167.454 57.96 171.828 ; 
        RECT 57.424 167.454 57.528 171.828 ; 
        RECT 56.992 167.454 57.096 171.828 ; 
        RECT 56.56 167.454 56.664 171.828 ; 
        RECT 56.128 167.454 56.232 171.828 ; 
        RECT 55.696 167.454 55.8 171.828 ; 
        RECT 55.264 167.454 55.368 171.828 ; 
        RECT 54.832 167.454 54.936 171.828 ; 
        RECT 54.4 167.454 54.504 171.828 ; 
        RECT 53.968 167.454 54.072 171.828 ; 
        RECT 53.536 167.454 53.64 171.828 ; 
        RECT 53.104 167.454 53.208 171.828 ; 
        RECT 52.672 167.454 52.776 171.828 ; 
        RECT 52.24 167.454 52.344 171.828 ; 
        RECT 51.808 167.454 51.912 171.828 ; 
        RECT 51.376 167.454 51.48 171.828 ; 
        RECT 50.944 167.454 51.048 171.828 ; 
        RECT 50.512 167.454 50.616 171.828 ; 
        RECT 50.08 167.454 50.184 171.828 ; 
        RECT 49.648 167.454 49.752 171.828 ; 
        RECT 49.216 167.454 49.32 171.828 ; 
        RECT 48.784 167.454 48.888 171.828 ; 
        RECT 48.352 167.454 48.456 171.828 ; 
        RECT 47.92 167.454 48.024 171.828 ; 
        RECT 47.488 167.454 47.592 171.828 ; 
        RECT 47.056 167.454 47.16 171.828 ; 
        RECT 46.624 167.454 46.728 171.828 ; 
        RECT 46.192 167.454 46.296 171.828 ; 
        RECT 45.76 167.454 45.864 171.828 ; 
        RECT 45.328 167.454 45.432 171.828 ; 
        RECT 44.896 167.454 45 171.828 ; 
        RECT 44.464 167.454 44.568 171.828 ; 
        RECT 44.032 167.454 44.136 171.828 ; 
        RECT 43.6 167.454 43.704 171.828 ; 
        RECT 43.168 167.454 43.272 171.828 ; 
        RECT 42.736 167.454 42.84 171.828 ; 
        RECT 42.304 167.454 42.408 171.828 ; 
        RECT 41.872 167.454 41.976 171.828 ; 
        RECT 41.44 167.454 41.544 171.828 ; 
        RECT 41.008 167.454 41.112 171.828 ; 
        RECT 40.576 167.454 40.68 171.828 ; 
        RECT 40.144 167.454 40.248 171.828 ; 
        RECT 39.712 167.454 39.816 171.828 ; 
        RECT 39.28 167.454 39.384 171.828 ; 
        RECT 38.848 167.454 38.952 171.828 ; 
        RECT 38.416 167.454 38.52 171.828 ; 
        RECT 37.984 167.454 38.088 171.828 ; 
        RECT 37.552 167.454 37.656 171.828 ; 
        RECT 36.7 167.454 37.008 171.828 ; 
        RECT 29.128 167.454 29.436 171.828 ; 
        RECT 28.48 167.454 28.584 171.828 ; 
        RECT 28.048 167.454 28.152 171.828 ; 
        RECT 27.616 167.454 27.72 171.828 ; 
        RECT 27.184 167.454 27.288 171.828 ; 
        RECT 26.752 167.454 26.856 171.828 ; 
        RECT 26.32 167.454 26.424 171.828 ; 
        RECT 25.888 167.454 25.992 171.828 ; 
        RECT 25.456 167.454 25.56 171.828 ; 
        RECT 25.024 167.454 25.128 171.828 ; 
        RECT 24.592 167.454 24.696 171.828 ; 
        RECT 24.16 167.454 24.264 171.828 ; 
        RECT 23.728 167.454 23.832 171.828 ; 
        RECT 23.296 167.454 23.4 171.828 ; 
        RECT 22.864 167.454 22.968 171.828 ; 
        RECT 22.432 167.454 22.536 171.828 ; 
        RECT 22 167.454 22.104 171.828 ; 
        RECT 21.568 167.454 21.672 171.828 ; 
        RECT 21.136 167.454 21.24 171.828 ; 
        RECT 20.704 167.454 20.808 171.828 ; 
        RECT 20.272 167.454 20.376 171.828 ; 
        RECT 19.84 167.454 19.944 171.828 ; 
        RECT 19.408 167.454 19.512 171.828 ; 
        RECT 18.976 167.454 19.08 171.828 ; 
        RECT 18.544 167.454 18.648 171.828 ; 
        RECT 18.112 167.454 18.216 171.828 ; 
        RECT 17.68 167.454 17.784 171.828 ; 
        RECT 17.248 167.454 17.352 171.828 ; 
        RECT 16.816 167.454 16.92 171.828 ; 
        RECT 16.384 167.454 16.488 171.828 ; 
        RECT 15.952 167.454 16.056 171.828 ; 
        RECT 15.52 167.454 15.624 171.828 ; 
        RECT 15.088 167.454 15.192 171.828 ; 
        RECT 14.656 167.454 14.76 171.828 ; 
        RECT 14.224 167.454 14.328 171.828 ; 
        RECT 13.792 167.454 13.896 171.828 ; 
        RECT 13.36 167.454 13.464 171.828 ; 
        RECT 12.928 167.454 13.032 171.828 ; 
        RECT 12.496 167.454 12.6 171.828 ; 
        RECT 12.064 167.454 12.168 171.828 ; 
        RECT 11.632 167.454 11.736 171.828 ; 
        RECT 11.2 167.454 11.304 171.828 ; 
        RECT 10.768 167.454 10.872 171.828 ; 
        RECT 10.336 167.454 10.44 171.828 ; 
        RECT 9.904 167.454 10.008 171.828 ; 
        RECT 9.472 167.454 9.576 171.828 ; 
        RECT 9.04 167.454 9.144 171.828 ; 
        RECT 8.608 167.454 8.712 171.828 ; 
        RECT 8.176 167.454 8.28 171.828 ; 
        RECT 7.744 167.454 7.848 171.828 ; 
        RECT 7.312 167.454 7.416 171.828 ; 
        RECT 6.88 167.454 6.984 171.828 ; 
        RECT 6.448 167.454 6.552 171.828 ; 
        RECT 6.016 167.454 6.12 171.828 ; 
        RECT 5.584 167.454 5.688 171.828 ; 
        RECT 5.152 167.454 5.256 171.828 ; 
        RECT 4.72 167.454 4.824 171.828 ; 
        RECT 4.288 167.454 4.392 171.828 ; 
        RECT 3.856 167.454 3.96 171.828 ; 
        RECT 3.424 167.454 3.528 171.828 ; 
        RECT 2.992 167.454 3.096 171.828 ; 
        RECT 2.56 167.454 2.664 171.828 ; 
        RECT 2.128 167.454 2.232 171.828 ; 
        RECT 1.696 167.454 1.8 171.828 ; 
        RECT 1.264 167.454 1.368 171.828 ; 
        RECT 0.832 167.454 0.936 171.828 ; 
        RECT 0.02 167.454 0.36 171.828 ; 
        RECT 34.564 171.774 35.076 176.148 ; 
        RECT 34.508 174.436 35.076 175.726 ; 
        RECT 33.916 173.344 34.164 176.148 ; 
        RECT 33.86 174.582 34.164 175.196 ; 
        RECT 33.916 171.774 34.02 176.148 ; 
        RECT 33.916 172.258 34.076 173.216 ; 
        RECT 33.916 171.774 34.164 172.13 ; 
        RECT 32.728 173.576 33.552 176.148 ; 
        RECT 33.448 171.774 33.552 176.148 ; 
        RECT 32.728 174.684 33.608 175.716 ; 
        RECT 32.728 171.774 33.12 176.148 ; 
        RECT 31.06 171.774 31.392 176.148 ; 
        RECT 31.06 172.128 31.448 175.87 ; 
        RECT 65.776 171.774 66.116 176.148 ; 
        RECT 65.2 171.774 65.304 176.148 ; 
        RECT 64.768 171.774 64.872 176.148 ; 
        RECT 64.336 171.774 64.44 176.148 ; 
        RECT 63.904 171.774 64.008 176.148 ; 
        RECT 63.472 171.774 63.576 176.148 ; 
        RECT 63.04 171.774 63.144 176.148 ; 
        RECT 62.608 171.774 62.712 176.148 ; 
        RECT 62.176 171.774 62.28 176.148 ; 
        RECT 61.744 171.774 61.848 176.148 ; 
        RECT 61.312 171.774 61.416 176.148 ; 
        RECT 60.88 171.774 60.984 176.148 ; 
        RECT 60.448 171.774 60.552 176.148 ; 
        RECT 60.016 171.774 60.12 176.148 ; 
        RECT 59.584 171.774 59.688 176.148 ; 
        RECT 59.152 171.774 59.256 176.148 ; 
        RECT 58.72 171.774 58.824 176.148 ; 
        RECT 58.288 171.774 58.392 176.148 ; 
        RECT 57.856 171.774 57.96 176.148 ; 
        RECT 57.424 171.774 57.528 176.148 ; 
        RECT 56.992 171.774 57.096 176.148 ; 
        RECT 56.56 171.774 56.664 176.148 ; 
        RECT 56.128 171.774 56.232 176.148 ; 
        RECT 55.696 171.774 55.8 176.148 ; 
        RECT 55.264 171.774 55.368 176.148 ; 
        RECT 54.832 171.774 54.936 176.148 ; 
        RECT 54.4 171.774 54.504 176.148 ; 
        RECT 53.968 171.774 54.072 176.148 ; 
        RECT 53.536 171.774 53.64 176.148 ; 
        RECT 53.104 171.774 53.208 176.148 ; 
        RECT 52.672 171.774 52.776 176.148 ; 
        RECT 52.24 171.774 52.344 176.148 ; 
        RECT 51.808 171.774 51.912 176.148 ; 
        RECT 51.376 171.774 51.48 176.148 ; 
        RECT 50.944 171.774 51.048 176.148 ; 
        RECT 50.512 171.774 50.616 176.148 ; 
        RECT 50.08 171.774 50.184 176.148 ; 
        RECT 49.648 171.774 49.752 176.148 ; 
        RECT 49.216 171.774 49.32 176.148 ; 
        RECT 48.784 171.774 48.888 176.148 ; 
        RECT 48.352 171.774 48.456 176.148 ; 
        RECT 47.92 171.774 48.024 176.148 ; 
        RECT 47.488 171.774 47.592 176.148 ; 
        RECT 47.056 171.774 47.16 176.148 ; 
        RECT 46.624 171.774 46.728 176.148 ; 
        RECT 46.192 171.774 46.296 176.148 ; 
        RECT 45.76 171.774 45.864 176.148 ; 
        RECT 45.328 171.774 45.432 176.148 ; 
        RECT 44.896 171.774 45 176.148 ; 
        RECT 44.464 171.774 44.568 176.148 ; 
        RECT 44.032 171.774 44.136 176.148 ; 
        RECT 43.6 171.774 43.704 176.148 ; 
        RECT 43.168 171.774 43.272 176.148 ; 
        RECT 42.736 171.774 42.84 176.148 ; 
        RECT 42.304 171.774 42.408 176.148 ; 
        RECT 41.872 171.774 41.976 176.148 ; 
        RECT 41.44 171.774 41.544 176.148 ; 
        RECT 41.008 171.774 41.112 176.148 ; 
        RECT 40.576 171.774 40.68 176.148 ; 
        RECT 40.144 171.774 40.248 176.148 ; 
        RECT 39.712 171.774 39.816 176.148 ; 
        RECT 39.28 171.774 39.384 176.148 ; 
        RECT 38.848 171.774 38.952 176.148 ; 
        RECT 38.416 171.774 38.52 176.148 ; 
        RECT 37.984 171.774 38.088 176.148 ; 
        RECT 37.552 171.774 37.656 176.148 ; 
        RECT 36.7 171.774 37.008 176.148 ; 
        RECT 29.128 171.774 29.436 176.148 ; 
        RECT 28.48 171.774 28.584 176.148 ; 
        RECT 28.048 171.774 28.152 176.148 ; 
        RECT 27.616 171.774 27.72 176.148 ; 
        RECT 27.184 171.774 27.288 176.148 ; 
        RECT 26.752 171.774 26.856 176.148 ; 
        RECT 26.32 171.774 26.424 176.148 ; 
        RECT 25.888 171.774 25.992 176.148 ; 
        RECT 25.456 171.774 25.56 176.148 ; 
        RECT 25.024 171.774 25.128 176.148 ; 
        RECT 24.592 171.774 24.696 176.148 ; 
        RECT 24.16 171.774 24.264 176.148 ; 
        RECT 23.728 171.774 23.832 176.148 ; 
        RECT 23.296 171.774 23.4 176.148 ; 
        RECT 22.864 171.774 22.968 176.148 ; 
        RECT 22.432 171.774 22.536 176.148 ; 
        RECT 22 171.774 22.104 176.148 ; 
        RECT 21.568 171.774 21.672 176.148 ; 
        RECT 21.136 171.774 21.24 176.148 ; 
        RECT 20.704 171.774 20.808 176.148 ; 
        RECT 20.272 171.774 20.376 176.148 ; 
        RECT 19.84 171.774 19.944 176.148 ; 
        RECT 19.408 171.774 19.512 176.148 ; 
        RECT 18.976 171.774 19.08 176.148 ; 
        RECT 18.544 171.774 18.648 176.148 ; 
        RECT 18.112 171.774 18.216 176.148 ; 
        RECT 17.68 171.774 17.784 176.148 ; 
        RECT 17.248 171.774 17.352 176.148 ; 
        RECT 16.816 171.774 16.92 176.148 ; 
        RECT 16.384 171.774 16.488 176.148 ; 
        RECT 15.952 171.774 16.056 176.148 ; 
        RECT 15.52 171.774 15.624 176.148 ; 
        RECT 15.088 171.774 15.192 176.148 ; 
        RECT 14.656 171.774 14.76 176.148 ; 
        RECT 14.224 171.774 14.328 176.148 ; 
        RECT 13.792 171.774 13.896 176.148 ; 
        RECT 13.36 171.774 13.464 176.148 ; 
        RECT 12.928 171.774 13.032 176.148 ; 
        RECT 12.496 171.774 12.6 176.148 ; 
        RECT 12.064 171.774 12.168 176.148 ; 
        RECT 11.632 171.774 11.736 176.148 ; 
        RECT 11.2 171.774 11.304 176.148 ; 
        RECT 10.768 171.774 10.872 176.148 ; 
        RECT 10.336 171.774 10.44 176.148 ; 
        RECT 9.904 171.774 10.008 176.148 ; 
        RECT 9.472 171.774 9.576 176.148 ; 
        RECT 9.04 171.774 9.144 176.148 ; 
        RECT 8.608 171.774 8.712 176.148 ; 
        RECT 8.176 171.774 8.28 176.148 ; 
        RECT 7.744 171.774 7.848 176.148 ; 
        RECT 7.312 171.774 7.416 176.148 ; 
        RECT 6.88 171.774 6.984 176.148 ; 
        RECT 6.448 171.774 6.552 176.148 ; 
        RECT 6.016 171.774 6.12 176.148 ; 
        RECT 5.584 171.774 5.688 176.148 ; 
        RECT 5.152 171.774 5.256 176.148 ; 
        RECT 4.72 171.774 4.824 176.148 ; 
        RECT 4.288 171.774 4.392 176.148 ; 
        RECT 3.856 171.774 3.96 176.148 ; 
        RECT 3.424 171.774 3.528 176.148 ; 
        RECT 2.992 171.774 3.096 176.148 ; 
        RECT 2.56 171.774 2.664 176.148 ; 
        RECT 2.128 171.774 2.232 176.148 ; 
        RECT 1.696 171.774 1.8 176.148 ; 
        RECT 1.264 171.774 1.368 176.148 ; 
        RECT 0.832 171.774 0.936 176.148 ; 
        RECT 0.02 171.774 0.36 176.148 ; 
        RECT 34.564 176.094 35.076 180.468 ; 
        RECT 34.508 178.756 35.076 180.046 ; 
        RECT 33.916 177.664 34.164 180.468 ; 
        RECT 33.86 178.902 34.164 179.516 ; 
        RECT 33.916 176.094 34.02 180.468 ; 
        RECT 33.916 176.578 34.076 177.536 ; 
        RECT 33.916 176.094 34.164 176.45 ; 
        RECT 32.728 177.896 33.552 180.468 ; 
        RECT 33.448 176.094 33.552 180.468 ; 
        RECT 32.728 179.004 33.608 180.036 ; 
        RECT 32.728 176.094 33.12 180.468 ; 
        RECT 31.06 176.094 31.392 180.468 ; 
        RECT 31.06 176.448 31.448 180.19 ; 
        RECT 65.776 176.094 66.116 180.468 ; 
        RECT 65.2 176.094 65.304 180.468 ; 
        RECT 64.768 176.094 64.872 180.468 ; 
        RECT 64.336 176.094 64.44 180.468 ; 
        RECT 63.904 176.094 64.008 180.468 ; 
        RECT 63.472 176.094 63.576 180.468 ; 
        RECT 63.04 176.094 63.144 180.468 ; 
        RECT 62.608 176.094 62.712 180.468 ; 
        RECT 62.176 176.094 62.28 180.468 ; 
        RECT 61.744 176.094 61.848 180.468 ; 
        RECT 61.312 176.094 61.416 180.468 ; 
        RECT 60.88 176.094 60.984 180.468 ; 
        RECT 60.448 176.094 60.552 180.468 ; 
        RECT 60.016 176.094 60.12 180.468 ; 
        RECT 59.584 176.094 59.688 180.468 ; 
        RECT 59.152 176.094 59.256 180.468 ; 
        RECT 58.72 176.094 58.824 180.468 ; 
        RECT 58.288 176.094 58.392 180.468 ; 
        RECT 57.856 176.094 57.96 180.468 ; 
        RECT 57.424 176.094 57.528 180.468 ; 
        RECT 56.992 176.094 57.096 180.468 ; 
        RECT 56.56 176.094 56.664 180.468 ; 
        RECT 56.128 176.094 56.232 180.468 ; 
        RECT 55.696 176.094 55.8 180.468 ; 
        RECT 55.264 176.094 55.368 180.468 ; 
        RECT 54.832 176.094 54.936 180.468 ; 
        RECT 54.4 176.094 54.504 180.468 ; 
        RECT 53.968 176.094 54.072 180.468 ; 
        RECT 53.536 176.094 53.64 180.468 ; 
        RECT 53.104 176.094 53.208 180.468 ; 
        RECT 52.672 176.094 52.776 180.468 ; 
        RECT 52.24 176.094 52.344 180.468 ; 
        RECT 51.808 176.094 51.912 180.468 ; 
        RECT 51.376 176.094 51.48 180.468 ; 
        RECT 50.944 176.094 51.048 180.468 ; 
        RECT 50.512 176.094 50.616 180.468 ; 
        RECT 50.08 176.094 50.184 180.468 ; 
        RECT 49.648 176.094 49.752 180.468 ; 
        RECT 49.216 176.094 49.32 180.468 ; 
        RECT 48.784 176.094 48.888 180.468 ; 
        RECT 48.352 176.094 48.456 180.468 ; 
        RECT 47.92 176.094 48.024 180.468 ; 
        RECT 47.488 176.094 47.592 180.468 ; 
        RECT 47.056 176.094 47.16 180.468 ; 
        RECT 46.624 176.094 46.728 180.468 ; 
        RECT 46.192 176.094 46.296 180.468 ; 
        RECT 45.76 176.094 45.864 180.468 ; 
        RECT 45.328 176.094 45.432 180.468 ; 
        RECT 44.896 176.094 45 180.468 ; 
        RECT 44.464 176.094 44.568 180.468 ; 
        RECT 44.032 176.094 44.136 180.468 ; 
        RECT 43.6 176.094 43.704 180.468 ; 
        RECT 43.168 176.094 43.272 180.468 ; 
        RECT 42.736 176.094 42.84 180.468 ; 
        RECT 42.304 176.094 42.408 180.468 ; 
        RECT 41.872 176.094 41.976 180.468 ; 
        RECT 41.44 176.094 41.544 180.468 ; 
        RECT 41.008 176.094 41.112 180.468 ; 
        RECT 40.576 176.094 40.68 180.468 ; 
        RECT 40.144 176.094 40.248 180.468 ; 
        RECT 39.712 176.094 39.816 180.468 ; 
        RECT 39.28 176.094 39.384 180.468 ; 
        RECT 38.848 176.094 38.952 180.468 ; 
        RECT 38.416 176.094 38.52 180.468 ; 
        RECT 37.984 176.094 38.088 180.468 ; 
        RECT 37.552 176.094 37.656 180.468 ; 
        RECT 36.7 176.094 37.008 180.468 ; 
        RECT 29.128 176.094 29.436 180.468 ; 
        RECT 28.48 176.094 28.584 180.468 ; 
        RECT 28.048 176.094 28.152 180.468 ; 
        RECT 27.616 176.094 27.72 180.468 ; 
        RECT 27.184 176.094 27.288 180.468 ; 
        RECT 26.752 176.094 26.856 180.468 ; 
        RECT 26.32 176.094 26.424 180.468 ; 
        RECT 25.888 176.094 25.992 180.468 ; 
        RECT 25.456 176.094 25.56 180.468 ; 
        RECT 25.024 176.094 25.128 180.468 ; 
        RECT 24.592 176.094 24.696 180.468 ; 
        RECT 24.16 176.094 24.264 180.468 ; 
        RECT 23.728 176.094 23.832 180.468 ; 
        RECT 23.296 176.094 23.4 180.468 ; 
        RECT 22.864 176.094 22.968 180.468 ; 
        RECT 22.432 176.094 22.536 180.468 ; 
        RECT 22 176.094 22.104 180.468 ; 
        RECT 21.568 176.094 21.672 180.468 ; 
        RECT 21.136 176.094 21.24 180.468 ; 
        RECT 20.704 176.094 20.808 180.468 ; 
        RECT 20.272 176.094 20.376 180.468 ; 
        RECT 19.84 176.094 19.944 180.468 ; 
        RECT 19.408 176.094 19.512 180.468 ; 
        RECT 18.976 176.094 19.08 180.468 ; 
        RECT 18.544 176.094 18.648 180.468 ; 
        RECT 18.112 176.094 18.216 180.468 ; 
        RECT 17.68 176.094 17.784 180.468 ; 
        RECT 17.248 176.094 17.352 180.468 ; 
        RECT 16.816 176.094 16.92 180.468 ; 
        RECT 16.384 176.094 16.488 180.468 ; 
        RECT 15.952 176.094 16.056 180.468 ; 
        RECT 15.52 176.094 15.624 180.468 ; 
        RECT 15.088 176.094 15.192 180.468 ; 
        RECT 14.656 176.094 14.76 180.468 ; 
        RECT 14.224 176.094 14.328 180.468 ; 
        RECT 13.792 176.094 13.896 180.468 ; 
        RECT 13.36 176.094 13.464 180.468 ; 
        RECT 12.928 176.094 13.032 180.468 ; 
        RECT 12.496 176.094 12.6 180.468 ; 
        RECT 12.064 176.094 12.168 180.468 ; 
        RECT 11.632 176.094 11.736 180.468 ; 
        RECT 11.2 176.094 11.304 180.468 ; 
        RECT 10.768 176.094 10.872 180.468 ; 
        RECT 10.336 176.094 10.44 180.468 ; 
        RECT 9.904 176.094 10.008 180.468 ; 
        RECT 9.472 176.094 9.576 180.468 ; 
        RECT 9.04 176.094 9.144 180.468 ; 
        RECT 8.608 176.094 8.712 180.468 ; 
        RECT 8.176 176.094 8.28 180.468 ; 
        RECT 7.744 176.094 7.848 180.468 ; 
        RECT 7.312 176.094 7.416 180.468 ; 
        RECT 6.88 176.094 6.984 180.468 ; 
        RECT 6.448 176.094 6.552 180.468 ; 
        RECT 6.016 176.094 6.12 180.468 ; 
        RECT 5.584 176.094 5.688 180.468 ; 
        RECT 5.152 176.094 5.256 180.468 ; 
        RECT 4.72 176.094 4.824 180.468 ; 
        RECT 4.288 176.094 4.392 180.468 ; 
        RECT 3.856 176.094 3.96 180.468 ; 
        RECT 3.424 176.094 3.528 180.468 ; 
        RECT 2.992 176.094 3.096 180.468 ; 
        RECT 2.56 176.094 2.664 180.468 ; 
        RECT 2.128 176.094 2.232 180.468 ; 
        RECT 1.696 176.094 1.8 180.468 ; 
        RECT 1.264 176.094 1.368 180.468 ; 
        RECT 0.832 176.094 0.936 180.468 ; 
        RECT 0.02 176.094 0.36 180.468 ; 
        RECT 34.564 180.414 35.076 184.788 ; 
        RECT 34.508 183.076 35.076 184.366 ; 
        RECT 33.916 181.984 34.164 184.788 ; 
        RECT 33.86 183.222 34.164 183.836 ; 
        RECT 33.916 180.414 34.02 184.788 ; 
        RECT 33.916 180.898 34.076 181.856 ; 
        RECT 33.916 180.414 34.164 180.77 ; 
        RECT 32.728 182.216 33.552 184.788 ; 
        RECT 33.448 180.414 33.552 184.788 ; 
        RECT 32.728 183.324 33.608 184.356 ; 
        RECT 32.728 180.414 33.12 184.788 ; 
        RECT 31.06 180.414 31.392 184.788 ; 
        RECT 31.06 180.768 31.448 184.51 ; 
        RECT 65.776 180.414 66.116 184.788 ; 
        RECT 65.2 180.414 65.304 184.788 ; 
        RECT 64.768 180.414 64.872 184.788 ; 
        RECT 64.336 180.414 64.44 184.788 ; 
        RECT 63.904 180.414 64.008 184.788 ; 
        RECT 63.472 180.414 63.576 184.788 ; 
        RECT 63.04 180.414 63.144 184.788 ; 
        RECT 62.608 180.414 62.712 184.788 ; 
        RECT 62.176 180.414 62.28 184.788 ; 
        RECT 61.744 180.414 61.848 184.788 ; 
        RECT 61.312 180.414 61.416 184.788 ; 
        RECT 60.88 180.414 60.984 184.788 ; 
        RECT 60.448 180.414 60.552 184.788 ; 
        RECT 60.016 180.414 60.12 184.788 ; 
        RECT 59.584 180.414 59.688 184.788 ; 
        RECT 59.152 180.414 59.256 184.788 ; 
        RECT 58.72 180.414 58.824 184.788 ; 
        RECT 58.288 180.414 58.392 184.788 ; 
        RECT 57.856 180.414 57.96 184.788 ; 
        RECT 57.424 180.414 57.528 184.788 ; 
        RECT 56.992 180.414 57.096 184.788 ; 
        RECT 56.56 180.414 56.664 184.788 ; 
        RECT 56.128 180.414 56.232 184.788 ; 
        RECT 55.696 180.414 55.8 184.788 ; 
        RECT 55.264 180.414 55.368 184.788 ; 
        RECT 54.832 180.414 54.936 184.788 ; 
        RECT 54.4 180.414 54.504 184.788 ; 
        RECT 53.968 180.414 54.072 184.788 ; 
        RECT 53.536 180.414 53.64 184.788 ; 
        RECT 53.104 180.414 53.208 184.788 ; 
        RECT 52.672 180.414 52.776 184.788 ; 
        RECT 52.24 180.414 52.344 184.788 ; 
        RECT 51.808 180.414 51.912 184.788 ; 
        RECT 51.376 180.414 51.48 184.788 ; 
        RECT 50.944 180.414 51.048 184.788 ; 
        RECT 50.512 180.414 50.616 184.788 ; 
        RECT 50.08 180.414 50.184 184.788 ; 
        RECT 49.648 180.414 49.752 184.788 ; 
        RECT 49.216 180.414 49.32 184.788 ; 
        RECT 48.784 180.414 48.888 184.788 ; 
        RECT 48.352 180.414 48.456 184.788 ; 
        RECT 47.92 180.414 48.024 184.788 ; 
        RECT 47.488 180.414 47.592 184.788 ; 
        RECT 47.056 180.414 47.16 184.788 ; 
        RECT 46.624 180.414 46.728 184.788 ; 
        RECT 46.192 180.414 46.296 184.788 ; 
        RECT 45.76 180.414 45.864 184.788 ; 
        RECT 45.328 180.414 45.432 184.788 ; 
        RECT 44.896 180.414 45 184.788 ; 
        RECT 44.464 180.414 44.568 184.788 ; 
        RECT 44.032 180.414 44.136 184.788 ; 
        RECT 43.6 180.414 43.704 184.788 ; 
        RECT 43.168 180.414 43.272 184.788 ; 
        RECT 42.736 180.414 42.84 184.788 ; 
        RECT 42.304 180.414 42.408 184.788 ; 
        RECT 41.872 180.414 41.976 184.788 ; 
        RECT 41.44 180.414 41.544 184.788 ; 
        RECT 41.008 180.414 41.112 184.788 ; 
        RECT 40.576 180.414 40.68 184.788 ; 
        RECT 40.144 180.414 40.248 184.788 ; 
        RECT 39.712 180.414 39.816 184.788 ; 
        RECT 39.28 180.414 39.384 184.788 ; 
        RECT 38.848 180.414 38.952 184.788 ; 
        RECT 38.416 180.414 38.52 184.788 ; 
        RECT 37.984 180.414 38.088 184.788 ; 
        RECT 37.552 180.414 37.656 184.788 ; 
        RECT 36.7 180.414 37.008 184.788 ; 
        RECT 29.128 180.414 29.436 184.788 ; 
        RECT 28.48 180.414 28.584 184.788 ; 
        RECT 28.048 180.414 28.152 184.788 ; 
        RECT 27.616 180.414 27.72 184.788 ; 
        RECT 27.184 180.414 27.288 184.788 ; 
        RECT 26.752 180.414 26.856 184.788 ; 
        RECT 26.32 180.414 26.424 184.788 ; 
        RECT 25.888 180.414 25.992 184.788 ; 
        RECT 25.456 180.414 25.56 184.788 ; 
        RECT 25.024 180.414 25.128 184.788 ; 
        RECT 24.592 180.414 24.696 184.788 ; 
        RECT 24.16 180.414 24.264 184.788 ; 
        RECT 23.728 180.414 23.832 184.788 ; 
        RECT 23.296 180.414 23.4 184.788 ; 
        RECT 22.864 180.414 22.968 184.788 ; 
        RECT 22.432 180.414 22.536 184.788 ; 
        RECT 22 180.414 22.104 184.788 ; 
        RECT 21.568 180.414 21.672 184.788 ; 
        RECT 21.136 180.414 21.24 184.788 ; 
        RECT 20.704 180.414 20.808 184.788 ; 
        RECT 20.272 180.414 20.376 184.788 ; 
        RECT 19.84 180.414 19.944 184.788 ; 
        RECT 19.408 180.414 19.512 184.788 ; 
        RECT 18.976 180.414 19.08 184.788 ; 
        RECT 18.544 180.414 18.648 184.788 ; 
        RECT 18.112 180.414 18.216 184.788 ; 
        RECT 17.68 180.414 17.784 184.788 ; 
        RECT 17.248 180.414 17.352 184.788 ; 
        RECT 16.816 180.414 16.92 184.788 ; 
        RECT 16.384 180.414 16.488 184.788 ; 
        RECT 15.952 180.414 16.056 184.788 ; 
        RECT 15.52 180.414 15.624 184.788 ; 
        RECT 15.088 180.414 15.192 184.788 ; 
        RECT 14.656 180.414 14.76 184.788 ; 
        RECT 14.224 180.414 14.328 184.788 ; 
        RECT 13.792 180.414 13.896 184.788 ; 
        RECT 13.36 180.414 13.464 184.788 ; 
        RECT 12.928 180.414 13.032 184.788 ; 
        RECT 12.496 180.414 12.6 184.788 ; 
        RECT 12.064 180.414 12.168 184.788 ; 
        RECT 11.632 180.414 11.736 184.788 ; 
        RECT 11.2 180.414 11.304 184.788 ; 
        RECT 10.768 180.414 10.872 184.788 ; 
        RECT 10.336 180.414 10.44 184.788 ; 
        RECT 9.904 180.414 10.008 184.788 ; 
        RECT 9.472 180.414 9.576 184.788 ; 
        RECT 9.04 180.414 9.144 184.788 ; 
        RECT 8.608 180.414 8.712 184.788 ; 
        RECT 8.176 180.414 8.28 184.788 ; 
        RECT 7.744 180.414 7.848 184.788 ; 
        RECT 7.312 180.414 7.416 184.788 ; 
        RECT 6.88 180.414 6.984 184.788 ; 
        RECT 6.448 180.414 6.552 184.788 ; 
        RECT 6.016 180.414 6.12 184.788 ; 
        RECT 5.584 180.414 5.688 184.788 ; 
        RECT 5.152 180.414 5.256 184.788 ; 
        RECT 4.72 180.414 4.824 184.788 ; 
        RECT 4.288 180.414 4.392 184.788 ; 
        RECT 3.856 180.414 3.96 184.788 ; 
        RECT 3.424 180.414 3.528 184.788 ; 
        RECT 2.992 180.414 3.096 184.788 ; 
        RECT 2.56 180.414 2.664 184.788 ; 
        RECT 2.128 180.414 2.232 184.788 ; 
        RECT 1.696 180.414 1.8 184.788 ; 
        RECT 1.264 180.414 1.368 184.788 ; 
        RECT 0.832 180.414 0.936 184.788 ; 
        RECT 0.02 180.414 0.36 184.788 ; 
        RECT 34.564 184.734 35.076 189.108 ; 
        RECT 34.508 187.396 35.076 188.686 ; 
        RECT 33.916 186.304 34.164 189.108 ; 
        RECT 33.86 187.542 34.164 188.156 ; 
        RECT 33.916 184.734 34.02 189.108 ; 
        RECT 33.916 185.218 34.076 186.176 ; 
        RECT 33.916 184.734 34.164 185.09 ; 
        RECT 32.728 186.536 33.552 189.108 ; 
        RECT 33.448 184.734 33.552 189.108 ; 
        RECT 32.728 187.644 33.608 188.676 ; 
        RECT 32.728 184.734 33.12 189.108 ; 
        RECT 31.06 184.734 31.392 189.108 ; 
        RECT 31.06 185.088 31.448 188.83 ; 
        RECT 65.776 184.734 66.116 189.108 ; 
        RECT 65.2 184.734 65.304 189.108 ; 
        RECT 64.768 184.734 64.872 189.108 ; 
        RECT 64.336 184.734 64.44 189.108 ; 
        RECT 63.904 184.734 64.008 189.108 ; 
        RECT 63.472 184.734 63.576 189.108 ; 
        RECT 63.04 184.734 63.144 189.108 ; 
        RECT 62.608 184.734 62.712 189.108 ; 
        RECT 62.176 184.734 62.28 189.108 ; 
        RECT 61.744 184.734 61.848 189.108 ; 
        RECT 61.312 184.734 61.416 189.108 ; 
        RECT 60.88 184.734 60.984 189.108 ; 
        RECT 60.448 184.734 60.552 189.108 ; 
        RECT 60.016 184.734 60.12 189.108 ; 
        RECT 59.584 184.734 59.688 189.108 ; 
        RECT 59.152 184.734 59.256 189.108 ; 
        RECT 58.72 184.734 58.824 189.108 ; 
        RECT 58.288 184.734 58.392 189.108 ; 
        RECT 57.856 184.734 57.96 189.108 ; 
        RECT 57.424 184.734 57.528 189.108 ; 
        RECT 56.992 184.734 57.096 189.108 ; 
        RECT 56.56 184.734 56.664 189.108 ; 
        RECT 56.128 184.734 56.232 189.108 ; 
        RECT 55.696 184.734 55.8 189.108 ; 
        RECT 55.264 184.734 55.368 189.108 ; 
        RECT 54.832 184.734 54.936 189.108 ; 
        RECT 54.4 184.734 54.504 189.108 ; 
        RECT 53.968 184.734 54.072 189.108 ; 
        RECT 53.536 184.734 53.64 189.108 ; 
        RECT 53.104 184.734 53.208 189.108 ; 
        RECT 52.672 184.734 52.776 189.108 ; 
        RECT 52.24 184.734 52.344 189.108 ; 
        RECT 51.808 184.734 51.912 189.108 ; 
        RECT 51.376 184.734 51.48 189.108 ; 
        RECT 50.944 184.734 51.048 189.108 ; 
        RECT 50.512 184.734 50.616 189.108 ; 
        RECT 50.08 184.734 50.184 189.108 ; 
        RECT 49.648 184.734 49.752 189.108 ; 
        RECT 49.216 184.734 49.32 189.108 ; 
        RECT 48.784 184.734 48.888 189.108 ; 
        RECT 48.352 184.734 48.456 189.108 ; 
        RECT 47.92 184.734 48.024 189.108 ; 
        RECT 47.488 184.734 47.592 189.108 ; 
        RECT 47.056 184.734 47.16 189.108 ; 
        RECT 46.624 184.734 46.728 189.108 ; 
        RECT 46.192 184.734 46.296 189.108 ; 
        RECT 45.76 184.734 45.864 189.108 ; 
        RECT 45.328 184.734 45.432 189.108 ; 
        RECT 44.896 184.734 45 189.108 ; 
        RECT 44.464 184.734 44.568 189.108 ; 
        RECT 44.032 184.734 44.136 189.108 ; 
        RECT 43.6 184.734 43.704 189.108 ; 
        RECT 43.168 184.734 43.272 189.108 ; 
        RECT 42.736 184.734 42.84 189.108 ; 
        RECT 42.304 184.734 42.408 189.108 ; 
        RECT 41.872 184.734 41.976 189.108 ; 
        RECT 41.44 184.734 41.544 189.108 ; 
        RECT 41.008 184.734 41.112 189.108 ; 
        RECT 40.576 184.734 40.68 189.108 ; 
        RECT 40.144 184.734 40.248 189.108 ; 
        RECT 39.712 184.734 39.816 189.108 ; 
        RECT 39.28 184.734 39.384 189.108 ; 
        RECT 38.848 184.734 38.952 189.108 ; 
        RECT 38.416 184.734 38.52 189.108 ; 
        RECT 37.984 184.734 38.088 189.108 ; 
        RECT 37.552 184.734 37.656 189.108 ; 
        RECT 36.7 184.734 37.008 189.108 ; 
        RECT 29.128 184.734 29.436 189.108 ; 
        RECT 28.48 184.734 28.584 189.108 ; 
        RECT 28.048 184.734 28.152 189.108 ; 
        RECT 27.616 184.734 27.72 189.108 ; 
        RECT 27.184 184.734 27.288 189.108 ; 
        RECT 26.752 184.734 26.856 189.108 ; 
        RECT 26.32 184.734 26.424 189.108 ; 
        RECT 25.888 184.734 25.992 189.108 ; 
        RECT 25.456 184.734 25.56 189.108 ; 
        RECT 25.024 184.734 25.128 189.108 ; 
        RECT 24.592 184.734 24.696 189.108 ; 
        RECT 24.16 184.734 24.264 189.108 ; 
        RECT 23.728 184.734 23.832 189.108 ; 
        RECT 23.296 184.734 23.4 189.108 ; 
        RECT 22.864 184.734 22.968 189.108 ; 
        RECT 22.432 184.734 22.536 189.108 ; 
        RECT 22 184.734 22.104 189.108 ; 
        RECT 21.568 184.734 21.672 189.108 ; 
        RECT 21.136 184.734 21.24 189.108 ; 
        RECT 20.704 184.734 20.808 189.108 ; 
        RECT 20.272 184.734 20.376 189.108 ; 
        RECT 19.84 184.734 19.944 189.108 ; 
        RECT 19.408 184.734 19.512 189.108 ; 
        RECT 18.976 184.734 19.08 189.108 ; 
        RECT 18.544 184.734 18.648 189.108 ; 
        RECT 18.112 184.734 18.216 189.108 ; 
        RECT 17.68 184.734 17.784 189.108 ; 
        RECT 17.248 184.734 17.352 189.108 ; 
        RECT 16.816 184.734 16.92 189.108 ; 
        RECT 16.384 184.734 16.488 189.108 ; 
        RECT 15.952 184.734 16.056 189.108 ; 
        RECT 15.52 184.734 15.624 189.108 ; 
        RECT 15.088 184.734 15.192 189.108 ; 
        RECT 14.656 184.734 14.76 189.108 ; 
        RECT 14.224 184.734 14.328 189.108 ; 
        RECT 13.792 184.734 13.896 189.108 ; 
        RECT 13.36 184.734 13.464 189.108 ; 
        RECT 12.928 184.734 13.032 189.108 ; 
        RECT 12.496 184.734 12.6 189.108 ; 
        RECT 12.064 184.734 12.168 189.108 ; 
        RECT 11.632 184.734 11.736 189.108 ; 
        RECT 11.2 184.734 11.304 189.108 ; 
        RECT 10.768 184.734 10.872 189.108 ; 
        RECT 10.336 184.734 10.44 189.108 ; 
        RECT 9.904 184.734 10.008 189.108 ; 
        RECT 9.472 184.734 9.576 189.108 ; 
        RECT 9.04 184.734 9.144 189.108 ; 
        RECT 8.608 184.734 8.712 189.108 ; 
        RECT 8.176 184.734 8.28 189.108 ; 
        RECT 7.744 184.734 7.848 189.108 ; 
        RECT 7.312 184.734 7.416 189.108 ; 
        RECT 6.88 184.734 6.984 189.108 ; 
        RECT 6.448 184.734 6.552 189.108 ; 
        RECT 6.016 184.734 6.12 189.108 ; 
        RECT 5.584 184.734 5.688 189.108 ; 
        RECT 5.152 184.734 5.256 189.108 ; 
        RECT 4.72 184.734 4.824 189.108 ; 
        RECT 4.288 184.734 4.392 189.108 ; 
        RECT 3.856 184.734 3.96 189.108 ; 
        RECT 3.424 184.734 3.528 189.108 ; 
        RECT 2.992 184.734 3.096 189.108 ; 
        RECT 2.56 184.734 2.664 189.108 ; 
        RECT 2.128 184.734 2.232 189.108 ; 
        RECT 1.696 184.734 1.8 189.108 ; 
        RECT 1.264 184.734 1.368 189.108 ; 
        RECT 0.832 184.734 0.936 189.108 ; 
        RECT 0.02 184.734 0.36 189.108 ; 
        RECT 34.564 189.054 35.076 193.428 ; 
        RECT 34.508 191.716 35.076 193.006 ; 
        RECT 33.916 190.624 34.164 193.428 ; 
        RECT 33.86 191.862 34.164 192.476 ; 
        RECT 33.916 189.054 34.02 193.428 ; 
        RECT 33.916 189.538 34.076 190.496 ; 
        RECT 33.916 189.054 34.164 189.41 ; 
        RECT 32.728 190.856 33.552 193.428 ; 
        RECT 33.448 189.054 33.552 193.428 ; 
        RECT 32.728 191.964 33.608 192.996 ; 
        RECT 32.728 189.054 33.12 193.428 ; 
        RECT 31.06 189.054 31.392 193.428 ; 
        RECT 31.06 189.408 31.448 193.15 ; 
        RECT 65.776 189.054 66.116 193.428 ; 
        RECT 65.2 189.054 65.304 193.428 ; 
        RECT 64.768 189.054 64.872 193.428 ; 
        RECT 64.336 189.054 64.44 193.428 ; 
        RECT 63.904 189.054 64.008 193.428 ; 
        RECT 63.472 189.054 63.576 193.428 ; 
        RECT 63.04 189.054 63.144 193.428 ; 
        RECT 62.608 189.054 62.712 193.428 ; 
        RECT 62.176 189.054 62.28 193.428 ; 
        RECT 61.744 189.054 61.848 193.428 ; 
        RECT 61.312 189.054 61.416 193.428 ; 
        RECT 60.88 189.054 60.984 193.428 ; 
        RECT 60.448 189.054 60.552 193.428 ; 
        RECT 60.016 189.054 60.12 193.428 ; 
        RECT 59.584 189.054 59.688 193.428 ; 
        RECT 59.152 189.054 59.256 193.428 ; 
        RECT 58.72 189.054 58.824 193.428 ; 
        RECT 58.288 189.054 58.392 193.428 ; 
        RECT 57.856 189.054 57.96 193.428 ; 
        RECT 57.424 189.054 57.528 193.428 ; 
        RECT 56.992 189.054 57.096 193.428 ; 
        RECT 56.56 189.054 56.664 193.428 ; 
        RECT 56.128 189.054 56.232 193.428 ; 
        RECT 55.696 189.054 55.8 193.428 ; 
        RECT 55.264 189.054 55.368 193.428 ; 
        RECT 54.832 189.054 54.936 193.428 ; 
        RECT 54.4 189.054 54.504 193.428 ; 
        RECT 53.968 189.054 54.072 193.428 ; 
        RECT 53.536 189.054 53.64 193.428 ; 
        RECT 53.104 189.054 53.208 193.428 ; 
        RECT 52.672 189.054 52.776 193.428 ; 
        RECT 52.24 189.054 52.344 193.428 ; 
        RECT 51.808 189.054 51.912 193.428 ; 
        RECT 51.376 189.054 51.48 193.428 ; 
        RECT 50.944 189.054 51.048 193.428 ; 
        RECT 50.512 189.054 50.616 193.428 ; 
        RECT 50.08 189.054 50.184 193.428 ; 
        RECT 49.648 189.054 49.752 193.428 ; 
        RECT 49.216 189.054 49.32 193.428 ; 
        RECT 48.784 189.054 48.888 193.428 ; 
        RECT 48.352 189.054 48.456 193.428 ; 
        RECT 47.92 189.054 48.024 193.428 ; 
        RECT 47.488 189.054 47.592 193.428 ; 
        RECT 47.056 189.054 47.16 193.428 ; 
        RECT 46.624 189.054 46.728 193.428 ; 
        RECT 46.192 189.054 46.296 193.428 ; 
        RECT 45.76 189.054 45.864 193.428 ; 
        RECT 45.328 189.054 45.432 193.428 ; 
        RECT 44.896 189.054 45 193.428 ; 
        RECT 44.464 189.054 44.568 193.428 ; 
        RECT 44.032 189.054 44.136 193.428 ; 
        RECT 43.6 189.054 43.704 193.428 ; 
        RECT 43.168 189.054 43.272 193.428 ; 
        RECT 42.736 189.054 42.84 193.428 ; 
        RECT 42.304 189.054 42.408 193.428 ; 
        RECT 41.872 189.054 41.976 193.428 ; 
        RECT 41.44 189.054 41.544 193.428 ; 
        RECT 41.008 189.054 41.112 193.428 ; 
        RECT 40.576 189.054 40.68 193.428 ; 
        RECT 40.144 189.054 40.248 193.428 ; 
        RECT 39.712 189.054 39.816 193.428 ; 
        RECT 39.28 189.054 39.384 193.428 ; 
        RECT 38.848 189.054 38.952 193.428 ; 
        RECT 38.416 189.054 38.52 193.428 ; 
        RECT 37.984 189.054 38.088 193.428 ; 
        RECT 37.552 189.054 37.656 193.428 ; 
        RECT 36.7 189.054 37.008 193.428 ; 
        RECT 29.128 189.054 29.436 193.428 ; 
        RECT 28.48 189.054 28.584 193.428 ; 
        RECT 28.048 189.054 28.152 193.428 ; 
        RECT 27.616 189.054 27.72 193.428 ; 
        RECT 27.184 189.054 27.288 193.428 ; 
        RECT 26.752 189.054 26.856 193.428 ; 
        RECT 26.32 189.054 26.424 193.428 ; 
        RECT 25.888 189.054 25.992 193.428 ; 
        RECT 25.456 189.054 25.56 193.428 ; 
        RECT 25.024 189.054 25.128 193.428 ; 
        RECT 24.592 189.054 24.696 193.428 ; 
        RECT 24.16 189.054 24.264 193.428 ; 
        RECT 23.728 189.054 23.832 193.428 ; 
        RECT 23.296 189.054 23.4 193.428 ; 
        RECT 22.864 189.054 22.968 193.428 ; 
        RECT 22.432 189.054 22.536 193.428 ; 
        RECT 22 189.054 22.104 193.428 ; 
        RECT 21.568 189.054 21.672 193.428 ; 
        RECT 21.136 189.054 21.24 193.428 ; 
        RECT 20.704 189.054 20.808 193.428 ; 
        RECT 20.272 189.054 20.376 193.428 ; 
        RECT 19.84 189.054 19.944 193.428 ; 
        RECT 19.408 189.054 19.512 193.428 ; 
        RECT 18.976 189.054 19.08 193.428 ; 
        RECT 18.544 189.054 18.648 193.428 ; 
        RECT 18.112 189.054 18.216 193.428 ; 
        RECT 17.68 189.054 17.784 193.428 ; 
        RECT 17.248 189.054 17.352 193.428 ; 
        RECT 16.816 189.054 16.92 193.428 ; 
        RECT 16.384 189.054 16.488 193.428 ; 
        RECT 15.952 189.054 16.056 193.428 ; 
        RECT 15.52 189.054 15.624 193.428 ; 
        RECT 15.088 189.054 15.192 193.428 ; 
        RECT 14.656 189.054 14.76 193.428 ; 
        RECT 14.224 189.054 14.328 193.428 ; 
        RECT 13.792 189.054 13.896 193.428 ; 
        RECT 13.36 189.054 13.464 193.428 ; 
        RECT 12.928 189.054 13.032 193.428 ; 
        RECT 12.496 189.054 12.6 193.428 ; 
        RECT 12.064 189.054 12.168 193.428 ; 
        RECT 11.632 189.054 11.736 193.428 ; 
        RECT 11.2 189.054 11.304 193.428 ; 
        RECT 10.768 189.054 10.872 193.428 ; 
        RECT 10.336 189.054 10.44 193.428 ; 
        RECT 9.904 189.054 10.008 193.428 ; 
        RECT 9.472 189.054 9.576 193.428 ; 
        RECT 9.04 189.054 9.144 193.428 ; 
        RECT 8.608 189.054 8.712 193.428 ; 
        RECT 8.176 189.054 8.28 193.428 ; 
        RECT 7.744 189.054 7.848 193.428 ; 
        RECT 7.312 189.054 7.416 193.428 ; 
        RECT 6.88 189.054 6.984 193.428 ; 
        RECT 6.448 189.054 6.552 193.428 ; 
        RECT 6.016 189.054 6.12 193.428 ; 
        RECT 5.584 189.054 5.688 193.428 ; 
        RECT 5.152 189.054 5.256 193.428 ; 
        RECT 4.72 189.054 4.824 193.428 ; 
        RECT 4.288 189.054 4.392 193.428 ; 
        RECT 3.856 189.054 3.96 193.428 ; 
        RECT 3.424 189.054 3.528 193.428 ; 
        RECT 2.992 189.054 3.096 193.428 ; 
        RECT 2.56 189.054 2.664 193.428 ; 
        RECT 2.128 189.054 2.232 193.428 ; 
        RECT 1.696 189.054 1.8 193.428 ; 
        RECT 1.264 189.054 1.368 193.428 ; 
        RECT 0.832 189.054 0.936 193.428 ; 
        RECT 0.02 189.054 0.36 193.428 ; 
        RECT 34.564 193.374 35.076 197.748 ; 
        RECT 34.508 196.036 35.076 197.326 ; 
        RECT 33.916 194.944 34.164 197.748 ; 
        RECT 33.86 196.182 34.164 196.796 ; 
        RECT 33.916 193.374 34.02 197.748 ; 
        RECT 33.916 193.858 34.076 194.816 ; 
        RECT 33.916 193.374 34.164 193.73 ; 
        RECT 32.728 195.176 33.552 197.748 ; 
        RECT 33.448 193.374 33.552 197.748 ; 
        RECT 32.728 196.284 33.608 197.316 ; 
        RECT 32.728 193.374 33.12 197.748 ; 
        RECT 31.06 193.374 31.392 197.748 ; 
        RECT 31.06 193.728 31.448 197.47 ; 
        RECT 65.776 193.374 66.116 197.748 ; 
        RECT 65.2 193.374 65.304 197.748 ; 
        RECT 64.768 193.374 64.872 197.748 ; 
        RECT 64.336 193.374 64.44 197.748 ; 
        RECT 63.904 193.374 64.008 197.748 ; 
        RECT 63.472 193.374 63.576 197.748 ; 
        RECT 63.04 193.374 63.144 197.748 ; 
        RECT 62.608 193.374 62.712 197.748 ; 
        RECT 62.176 193.374 62.28 197.748 ; 
        RECT 61.744 193.374 61.848 197.748 ; 
        RECT 61.312 193.374 61.416 197.748 ; 
        RECT 60.88 193.374 60.984 197.748 ; 
        RECT 60.448 193.374 60.552 197.748 ; 
        RECT 60.016 193.374 60.12 197.748 ; 
        RECT 59.584 193.374 59.688 197.748 ; 
        RECT 59.152 193.374 59.256 197.748 ; 
        RECT 58.72 193.374 58.824 197.748 ; 
        RECT 58.288 193.374 58.392 197.748 ; 
        RECT 57.856 193.374 57.96 197.748 ; 
        RECT 57.424 193.374 57.528 197.748 ; 
        RECT 56.992 193.374 57.096 197.748 ; 
        RECT 56.56 193.374 56.664 197.748 ; 
        RECT 56.128 193.374 56.232 197.748 ; 
        RECT 55.696 193.374 55.8 197.748 ; 
        RECT 55.264 193.374 55.368 197.748 ; 
        RECT 54.832 193.374 54.936 197.748 ; 
        RECT 54.4 193.374 54.504 197.748 ; 
        RECT 53.968 193.374 54.072 197.748 ; 
        RECT 53.536 193.374 53.64 197.748 ; 
        RECT 53.104 193.374 53.208 197.748 ; 
        RECT 52.672 193.374 52.776 197.748 ; 
        RECT 52.24 193.374 52.344 197.748 ; 
        RECT 51.808 193.374 51.912 197.748 ; 
        RECT 51.376 193.374 51.48 197.748 ; 
        RECT 50.944 193.374 51.048 197.748 ; 
        RECT 50.512 193.374 50.616 197.748 ; 
        RECT 50.08 193.374 50.184 197.748 ; 
        RECT 49.648 193.374 49.752 197.748 ; 
        RECT 49.216 193.374 49.32 197.748 ; 
        RECT 48.784 193.374 48.888 197.748 ; 
        RECT 48.352 193.374 48.456 197.748 ; 
        RECT 47.92 193.374 48.024 197.748 ; 
        RECT 47.488 193.374 47.592 197.748 ; 
        RECT 47.056 193.374 47.16 197.748 ; 
        RECT 46.624 193.374 46.728 197.748 ; 
        RECT 46.192 193.374 46.296 197.748 ; 
        RECT 45.76 193.374 45.864 197.748 ; 
        RECT 45.328 193.374 45.432 197.748 ; 
        RECT 44.896 193.374 45 197.748 ; 
        RECT 44.464 193.374 44.568 197.748 ; 
        RECT 44.032 193.374 44.136 197.748 ; 
        RECT 43.6 193.374 43.704 197.748 ; 
        RECT 43.168 193.374 43.272 197.748 ; 
        RECT 42.736 193.374 42.84 197.748 ; 
        RECT 42.304 193.374 42.408 197.748 ; 
        RECT 41.872 193.374 41.976 197.748 ; 
        RECT 41.44 193.374 41.544 197.748 ; 
        RECT 41.008 193.374 41.112 197.748 ; 
        RECT 40.576 193.374 40.68 197.748 ; 
        RECT 40.144 193.374 40.248 197.748 ; 
        RECT 39.712 193.374 39.816 197.748 ; 
        RECT 39.28 193.374 39.384 197.748 ; 
        RECT 38.848 193.374 38.952 197.748 ; 
        RECT 38.416 193.374 38.52 197.748 ; 
        RECT 37.984 193.374 38.088 197.748 ; 
        RECT 37.552 193.374 37.656 197.748 ; 
        RECT 36.7 193.374 37.008 197.748 ; 
        RECT 29.128 193.374 29.436 197.748 ; 
        RECT 28.48 193.374 28.584 197.748 ; 
        RECT 28.048 193.374 28.152 197.748 ; 
        RECT 27.616 193.374 27.72 197.748 ; 
        RECT 27.184 193.374 27.288 197.748 ; 
        RECT 26.752 193.374 26.856 197.748 ; 
        RECT 26.32 193.374 26.424 197.748 ; 
        RECT 25.888 193.374 25.992 197.748 ; 
        RECT 25.456 193.374 25.56 197.748 ; 
        RECT 25.024 193.374 25.128 197.748 ; 
        RECT 24.592 193.374 24.696 197.748 ; 
        RECT 24.16 193.374 24.264 197.748 ; 
        RECT 23.728 193.374 23.832 197.748 ; 
        RECT 23.296 193.374 23.4 197.748 ; 
        RECT 22.864 193.374 22.968 197.748 ; 
        RECT 22.432 193.374 22.536 197.748 ; 
        RECT 22 193.374 22.104 197.748 ; 
        RECT 21.568 193.374 21.672 197.748 ; 
        RECT 21.136 193.374 21.24 197.748 ; 
        RECT 20.704 193.374 20.808 197.748 ; 
        RECT 20.272 193.374 20.376 197.748 ; 
        RECT 19.84 193.374 19.944 197.748 ; 
        RECT 19.408 193.374 19.512 197.748 ; 
        RECT 18.976 193.374 19.08 197.748 ; 
        RECT 18.544 193.374 18.648 197.748 ; 
        RECT 18.112 193.374 18.216 197.748 ; 
        RECT 17.68 193.374 17.784 197.748 ; 
        RECT 17.248 193.374 17.352 197.748 ; 
        RECT 16.816 193.374 16.92 197.748 ; 
        RECT 16.384 193.374 16.488 197.748 ; 
        RECT 15.952 193.374 16.056 197.748 ; 
        RECT 15.52 193.374 15.624 197.748 ; 
        RECT 15.088 193.374 15.192 197.748 ; 
        RECT 14.656 193.374 14.76 197.748 ; 
        RECT 14.224 193.374 14.328 197.748 ; 
        RECT 13.792 193.374 13.896 197.748 ; 
        RECT 13.36 193.374 13.464 197.748 ; 
        RECT 12.928 193.374 13.032 197.748 ; 
        RECT 12.496 193.374 12.6 197.748 ; 
        RECT 12.064 193.374 12.168 197.748 ; 
        RECT 11.632 193.374 11.736 197.748 ; 
        RECT 11.2 193.374 11.304 197.748 ; 
        RECT 10.768 193.374 10.872 197.748 ; 
        RECT 10.336 193.374 10.44 197.748 ; 
        RECT 9.904 193.374 10.008 197.748 ; 
        RECT 9.472 193.374 9.576 197.748 ; 
        RECT 9.04 193.374 9.144 197.748 ; 
        RECT 8.608 193.374 8.712 197.748 ; 
        RECT 8.176 193.374 8.28 197.748 ; 
        RECT 7.744 193.374 7.848 197.748 ; 
        RECT 7.312 193.374 7.416 197.748 ; 
        RECT 6.88 193.374 6.984 197.748 ; 
        RECT 6.448 193.374 6.552 197.748 ; 
        RECT 6.016 193.374 6.12 197.748 ; 
        RECT 5.584 193.374 5.688 197.748 ; 
        RECT 5.152 193.374 5.256 197.748 ; 
        RECT 4.72 193.374 4.824 197.748 ; 
        RECT 4.288 193.374 4.392 197.748 ; 
        RECT 3.856 193.374 3.96 197.748 ; 
        RECT 3.424 193.374 3.528 197.748 ; 
        RECT 2.992 193.374 3.096 197.748 ; 
        RECT 2.56 193.374 2.664 197.748 ; 
        RECT 2.128 193.374 2.232 197.748 ; 
        RECT 1.696 193.374 1.8 197.748 ; 
        RECT 1.264 193.374 1.368 197.748 ; 
        RECT 0.832 193.374 0.936 197.748 ; 
        RECT 0.02 193.374 0.36 197.748 ; 
        RECT 34.564 197.694 35.076 202.068 ; 
        RECT 34.508 200.356 35.076 201.646 ; 
        RECT 33.916 199.264 34.164 202.068 ; 
        RECT 33.86 200.502 34.164 201.116 ; 
        RECT 33.916 197.694 34.02 202.068 ; 
        RECT 33.916 198.178 34.076 199.136 ; 
        RECT 33.916 197.694 34.164 198.05 ; 
        RECT 32.728 199.496 33.552 202.068 ; 
        RECT 33.448 197.694 33.552 202.068 ; 
        RECT 32.728 200.604 33.608 201.636 ; 
        RECT 32.728 197.694 33.12 202.068 ; 
        RECT 31.06 197.694 31.392 202.068 ; 
        RECT 31.06 198.048 31.448 201.79 ; 
        RECT 65.776 197.694 66.116 202.068 ; 
        RECT 65.2 197.694 65.304 202.068 ; 
        RECT 64.768 197.694 64.872 202.068 ; 
        RECT 64.336 197.694 64.44 202.068 ; 
        RECT 63.904 197.694 64.008 202.068 ; 
        RECT 63.472 197.694 63.576 202.068 ; 
        RECT 63.04 197.694 63.144 202.068 ; 
        RECT 62.608 197.694 62.712 202.068 ; 
        RECT 62.176 197.694 62.28 202.068 ; 
        RECT 61.744 197.694 61.848 202.068 ; 
        RECT 61.312 197.694 61.416 202.068 ; 
        RECT 60.88 197.694 60.984 202.068 ; 
        RECT 60.448 197.694 60.552 202.068 ; 
        RECT 60.016 197.694 60.12 202.068 ; 
        RECT 59.584 197.694 59.688 202.068 ; 
        RECT 59.152 197.694 59.256 202.068 ; 
        RECT 58.72 197.694 58.824 202.068 ; 
        RECT 58.288 197.694 58.392 202.068 ; 
        RECT 57.856 197.694 57.96 202.068 ; 
        RECT 57.424 197.694 57.528 202.068 ; 
        RECT 56.992 197.694 57.096 202.068 ; 
        RECT 56.56 197.694 56.664 202.068 ; 
        RECT 56.128 197.694 56.232 202.068 ; 
        RECT 55.696 197.694 55.8 202.068 ; 
        RECT 55.264 197.694 55.368 202.068 ; 
        RECT 54.832 197.694 54.936 202.068 ; 
        RECT 54.4 197.694 54.504 202.068 ; 
        RECT 53.968 197.694 54.072 202.068 ; 
        RECT 53.536 197.694 53.64 202.068 ; 
        RECT 53.104 197.694 53.208 202.068 ; 
        RECT 52.672 197.694 52.776 202.068 ; 
        RECT 52.24 197.694 52.344 202.068 ; 
        RECT 51.808 197.694 51.912 202.068 ; 
        RECT 51.376 197.694 51.48 202.068 ; 
        RECT 50.944 197.694 51.048 202.068 ; 
        RECT 50.512 197.694 50.616 202.068 ; 
        RECT 50.08 197.694 50.184 202.068 ; 
        RECT 49.648 197.694 49.752 202.068 ; 
        RECT 49.216 197.694 49.32 202.068 ; 
        RECT 48.784 197.694 48.888 202.068 ; 
        RECT 48.352 197.694 48.456 202.068 ; 
        RECT 47.92 197.694 48.024 202.068 ; 
        RECT 47.488 197.694 47.592 202.068 ; 
        RECT 47.056 197.694 47.16 202.068 ; 
        RECT 46.624 197.694 46.728 202.068 ; 
        RECT 46.192 197.694 46.296 202.068 ; 
        RECT 45.76 197.694 45.864 202.068 ; 
        RECT 45.328 197.694 45.432 202.068 ; 
        RECT 44.896 197.694 45 202.068 ; 
        RECT 44.464 197.694 44.568 202.068 ; 
        RECT 44.032 197.694 44.136 202.068 ; 
        RECT 43.6 197.694 43.704 202.068 ; 
        RECT 43.168 197.694 43.272 202.068 ; 
        RECT 42.736 197.694 42.84 202.068 ; 
        RECT 42.304 197.694 42.408 202.068 ; 
        RECT 41.872 197.694 41.976 202.068 ; 
        RECT 41.44 197.694 41.544 202.068 ; 
        RECT 41.008 197.694 41.112 202.068 ; 
        RECT 40.576 197.694 40.68 202.068 ; 
        RECT 40.144 197.694 40.248 202.068 ; 
        RECT 39.712 197.694 39.816 202.068 ; 
        RECT 39.28 197.694 39.384 202.068 ; 
        RECT 38.848 197.694 38.952 202.068 ; 
        RECT 38.416 197.694 38.52 202.068 ; 
        RECT 37.984 197.694 38.088 202.068 ; 
        RECT 37.552 197.694 37.656 202.068 ; 
        RECT 36.7 197.694 37.008 202.068 ; 
        RECT 29.128 197.694 29.436 202.068 ; 
        RECT 28.48 197.694 28.584 202.068 ; 
        RECT 28.048 197.694 28.152 202.068 ; 
        RECT 27.616 197.694 27.72 202.068 ; 
        RECT 27.184 197.694 27.288 202.068 ; 
        RECT 26.752 197.694 26.856 202.068 ; 
        RECT 26.32 197.694 26.424 202.068 ; 
        RECT 25.888 197.694 25.992 202.068 ; 
        RECT 25.456 197.694 25.56 202.068 ; 
        RECT 25.024 197.694 25.128 202.068 ; 
        RECT 24.592 197.694 24.696 202.068 ; 
        RECT 24.16 197.694 24.264 202.068 ; 
        RECT 23.728 197.694 23.832 202.068 ; 
        RECT 23.296 197.694 23.4 202.068 ; 
        RECT 22.864 197.694 22.968 202.068 ; 
        RECT 22.432 197.694 22.536 202.068 ; 
        RECT 22 197.694 22.104 202.068 ; 
        RECT 21.568 197.694 21.672 202.068 ; 
        RECT 21.136 197.694 21.24 202.068 ; 
        RECT 20.704 197.694 20.808 202.068 ; 
        RECT 20.272 197.694 20.376 202.068 ; 
        RECT 19.84 197.694 19.944 202.068 ; 
        RECT 19.408 197.694 19.512 202.068 ; 
        RECT 18.976 197.694 19.08 202.068 ; 
        RECT 18.544 197.694 18.648 202.068 ; 
        RECT 18.112 197.694 18.216 202.068 ; 
        RECT 17.68 197.694 17.784 202.068 ; 
        RECT 17.248 197.694 17.352 202.068 ; 
        RECT 16.816 197.694 16.92 202.068 ; 
        RECT 16.384 197.694 16.488 202.068 ; 
        RECT 15.952 197.694 16.056 202.068 ; 
        RECT 15.52 197.694 15.624 202.068 ; 
        RECT 15.088 197.694 15.192 202.068 ; 
        RECT 14.656 197.694 14.76 202.068 ; 
        RECT 14.224 197.694 14.328 202.068 ; 
        RECT 13.792 197.694 13.896 202.068 ; 
        RECT 13.36 197.694 13.464 202.068 ; 
        RECT 12.928 197.694 13.032 202.068 ; 
        RECT 12.496 197.694 12.6 202.068 ; 
        RECT 12.064 197.694 12.168 202.068 ; 
        RECT 11.632 197.694 11.736 202.068 ; 
        RECT 11.2 197.694 11.304 202.068 ; 
        RECT 10.768 197.694 10.872 202.068 ; 
        RECT 10.336 197.694 10.44 202.068 ; 
        RECT 9.904 197.694 10.008 202.068 ; 
        RECT 9.472 197.694 9.576 202.068 ; 
        RECT 9.04 197.694 9.144 202.068 ; 
        RECT 8.608 197.694 8.712 202.068 ; 
        RECT 8.176 197.694 8.28 202.068 ; 
        RECT 7.744 197.694 7.848 202.068 ; 
        RECT 7.312 197.694 7.416 202.068 ; 
        RECT 6.88 197.694 6.984 202.068 ; 
        RECT 6.448 197.694 6.552 202.068 ; 
        RECT 6.016 197.694 6.12 202.068 ; 
        RECT 5.584 197.694 5.688 202.068 ; 
        RECT 5.152 197.694 5.256 202.068 ; 
        RECT 4.72 197.694 4.824 202.068 ; 
        RECT 4.288 197.694 4.392 202.068 ; 
        RECT 3.856 197.694 3.96 202.068 ; 
        RECT 3.424 197.694 3.528 202.068 ; 
        RECT 2.992 197.694 3.096 202.068 ; 
        RECT 2.56 197.694 2.664 202.068 ; 
        RECT 2.128 197.694 2.232 202.068 ; 
        RECT 1.696 197.694 1.8 202.068 ; 
        RECT 1.264 197.694 1.368 202.068 ; 
        RECT 0.832 197.694 0.936 202.068 ; 
        RECT 0.02 197.694 0.36 202.068 ; 
        RECT 34.564 202.014 35.076 206.388 ; 
        RECT 34.508 204.676 35.076 205.966 ; 
        RECT 33.916 203.584 34.164 206.388 ; 
        RECT 33.86 204.822 34.164 205.436 ; 
        RECT 33.916 202.014 34.02 206.388 ; 
        RECT 33.916 202.498 34.076 203.456 ; 
        RECT 33.916 202.014 34.164 202.37 ; 
        RECT 32.728 203.816 33.552 206.388 ; 
        RECT 33.448 202.014 33.552 206.388 ; 
        RECT 32.728 204.924 33.608 205.956 ; 
        RECT 32.728 202.014 33.12 206.388 ; 
        RECT 31.06 202.014 31.392 206.388 ; 
        RECT 31.06 202.368 31.448 206.11 ; 
        RECT 65.776 202.014 66.116 206.388 ; 
        RECT 65.2 202.014 65.304 206.388 ; 
        RECT 64.768 202.014 64.872 206.388 ; 
        RECT 64.336 202.014 64.44 206.388 ; 
        RECT 63.904 202.014 64.008 206.388 ; 
        RECT 63.472 202.014 63.576 206.388 ; 
        RECT 63.04 202.014 63.144 206.388 ; 
        RECT 62.608 202.014 62.712 206.388 ; 
        RECT 62.176 202.014 62.28 206.388 ; 
        RECT 61.744 202.014 61.848 206.388 ; 
        RECT 61.312 202.014 61.416 206.388 ; 
        RECT 60.88 202.014 60.984 206.388 ; 
        RECT 60.448 202.014 60.552 206.388 ; 
        RECT 60.016 202.014 60.12 206.388 ; 
        RECT 59.584 202.014 59.688 206.388 ; 
        RECT 59.152 202.014 59.256 206.388 ; 
        RECT 58.72 202.014 58.824 206.388 ; 
        RECT 58.288 202.014 58.392 206.388 ; 
        RECT 57.856 202.014 57.96 206.388 ; 
        RECT 57.424 202.014 57.528 206.388 ; 
        RECT 56.992 202.014 57.096 206.388 ; 
        RECT 56.56 202.014 56.664 206.388 ; 
        RECT 56.128 202.014 56.232 206.388 ; 
        RECT 55.696 202.014 55.8 206.388 ; 
        RECT 55.264 202.014 55.368 206.388 ; 
        RECT 54.832 202.014 54.936 206.388 ; 
        RECT 54.4 202.014 54.504 206.388 ; 
        RECT 53.968 202.014 54.072 206.388 ; 
        RECT 53.536 202.014 53.64 206.388 ; 
        RECT 53.104 202.014 53.208 206.388 ; 
        RECT 52.672 202.014 52.776 206.388 ; 
        RECT 52.24 202.014 52.344 206.388 ; 
        RECT 51.808 202.014 51.912 206.388 ; 
        RECT 51.376 202.014 51.48 206.388 ; 
        RECT 50.944 202.014 51.048 206.388 ; 
        RECT 50.512 202.014 50.616 206.388 ; 
        RECT 50.08 202.014 50.184 206.388 ; 
        RECT 49.648 202.014 49.752 206.388 ; 
        RECT 49.216 202.014 49.32 206.388 ; 
        RECT 48.784 202.014 48.888 206.388 ; 
        RECT 48.352 202.014 48.456 206.388 ; 
        RECT 47.92 202.014 48.024 206.388 ; 
        RECT 47.488 202.014 47.592 206.388 ; 
        RECT 47.056 202.014 47.16 206.388 ; 
        RECT 46.624 202.014 46.728 206.388 ; 
        RECT 46.192 202.014 46.296 206.388 ; 
        RECT 45.76 202.014 45.864 206.388 ; 
        RECT 45.328 202.014 45.432 206.388 ; 
        RECT 44.896 202.014 45 206.388 ; 
        RECT 44.464 202.014 44.568 206.388 ; 
        RECT 44.032 202.014 44.136 206.388 ; 
        RECT 43.6 202.014 43.704 206.388 ; 
        RECT 43.168 202.014 43.272 206.388 ; 
        RECT 42.736 202.014 42.84 206.388 ; 
        RECT 42.304 202.014 42.408 206.388 ; 
        RECT 41.872 202.014 41.976 206.388 ; 
        RECT 41.44 202.014 41.544 206.388 ; 
        RECT 41.008 202.014 41.112 206.388 ; 
        RECT 40.576 202.014 40.68 206.388 ; 
        RECT 40.144 202.014 40.248 206.388 ; 
        RECT 39.712 202.014 39.816 206.388 ; 
        RECT 39.28 202.014 39.384 206.388 ; 
        RECT 38.848 202.014 38.952 206.388 ; 
        RECT 38.416 202.014 38.52 206.388 ; 
        RECT 37.984 202.014 38.088 206.388 ; 
        RECT 37.552 202.014 37.656 206.388 ; 
        RECT 36.7 202.014 37.008 206.388 ; 
        RECT 29.128 202.014 29.436 206.388 ; 
        RECT 28.48 202.014 28.584 206.388 ; 
        RECT 28.048 202.014 28.152 206.388 ; 
        RECT 27.616 202.014 27.72 206.388 ; 
        RECT 27.184 202.014 27.288 206.388 ; 
        RECT 26.752 202.014 26.856 206.388 ; 
        RECT 26.32 202.014 26.424 206.388 ; 
        RECT 25.888 202.014 25.992 206.388 ; 
        RECT 25.456 202.014 25.56 206.388 ; 
        RECT 25.024 202.014 25.128 206.388 ; 
        RECT 24.592 202.014 24.696 206.388 ; 
        RECT 24.16 202.014 24.264 206.388 ; 
        RECT 23.728 202.014 23.832 206.388 ; 
        RECT 23.296 202.014 23.4 206.388 ; 
        RECT 22.864 202.014 22.968 206.388 ; 
        RECT 22.432 202.014 22.536 206.388 ; 
        RECT 22 202.014 22.104 206.388 ; 
        RECT 21.568 202.014 21.672 206.388 ; 
        RECT 21.136 202.014 21.24 206.388 ; 
        RECT 20.704 202.014 20.808 206.388 ; 
        RECT 20.272 202.014 20.376 206.388 ; 
        RECT 19.84 202.014 19.944 206.388 ; 
        RECT 19.408 202.014 19.512 206.388 ; 
        RECT 18.976 202.014 19.08 206.388 ; 
        RECT 18.544 202.014 18.648 206.388 ; 
        RECT 18.112 202.014 18.216 206.388 ; 
        RECT 17.68 202.014 17.784 206.388 ; 
        RECT 17.248 202.014 17.352 206.388 ; 
        RECT 16.816 202.014 16.92 206.388 ; 
        RECT 16.384 202.014 16.488 206.388 ; 
        RECT 15.952 202.014 16.056 206.388 ; 
        RECT 15.52 202.014 15.624 206.388 ; 
        RECT 15.088 202.014 15.192 206.388 ; 
        RECT 14.656 202.014 14.76 206.388 ; 
        RECT 14.224 202.014 14.328 206.388 ; 
        RECT 13.792 202.014 13.896 206.388 ; 
        RECT 13.36 202.014 13.464 206.388 ; 
        RECT 12.928 202.014 13.032 206.388 ; 
        RECT 12.496 202.014 12.6 206.388 ; 
        RECT 12.064 202.014 12.168 206.388 ; 
        RECT 11.632 202.014 11.736 206.388 ; 
        RECT 11.2 202.014 11.304 206.388 ; 
        RECT 10.768 202.014 10.872 206.388 ; 
        RECT 10.336 202.014 10.44 206.388 ; 
        RECT 9.904 202.014 10.008 206.388 ; 
        RECT 9.472 202.014 9.576 206.388 ; 
        RECT 9.04 202.014 9.144 206.388 ; 
        RECT 8.608 202.014 8.712 206.388 ; 
        RECT 8.176 202.014 8.28 206.388 ; 
        RECT 7.744 202.014 7.848 206.388 ; 
        RECT 7.312 202.014 7.416 206.388 ; 
        RECT 6.88 202.014 6.984 206.388 ; 
        RECT 6.448 202.014 6.552 206.388 ; 
        RECT 6.016 202.014 6.12 206.388 ; 
        RECT 5.584 202.014 5.688 206.388 ; 
        RECT 5.152 202.014 5.256 206.388 ; 
        RECT 4.72 202.014 4.824 206.388 ; 
        RECT 4.288 202.014 4.392 206.388 ; 
        RECT 3.856 202.014 3.96 206.388 ; 
        RECT 3.424 202.014 3.528 206.388 ; 
        RECT 2.992 202.014 3.096 206.388 ; 
        RECT 2.56 202.014 2.664 206.388 ; 
        RECT 2.128 202.014 2.232 206.388 ; 
        RECT 1.696 202.014 1.8 206.388 ; 
        RECT 1.264 202.014 1.368 206.388 ; 
        RECT 0.832 202.014 0.936 206.388 ; 
        RECT 0.02 202.014 0.36 206.388 ; 
        RECT 34.564 206.334 35.076 210.708 ; 
        RECT 34.508 208.996 35.076 210.286 ; 
        RECT 33.916 207.904 34.164 210.708 ; 
        RECT 33.86 209.142 34.164 209.756 ; 
        RECT 33.916 206.334 34.02 210.708 ; 
        RECT 33.916 206.818 34.076 207.776 ; 
        RECT 33.916 206.334 34.164 206.69 ; 
        RECT 32.728 208.136 33.552 210.708 ; 
        RECT 33.448 206.334 33.552 210.708 ; 
        RECT 32.728 209.244 33.608 210.276 ; 
        RECT 32.728 206.334 33.12 210.708 ; 
        RECT 31.06 206.334 31.392 210.708 ; 
        RECT 31.06 206.688 31.448 210.43 ; 
        RECT 65.776 206.334 66.116 210.708 ; 
        RECT 65.2 206.334 65.304 210.708 ; 
        RECT 64.768 206.334 64.872 210.708 ; 
        RECT 64.336 206.334 64.44 210.708 ; 
        RECT 63.904 206.334 64.008 210.708 ; 
        RECT 63.472 206.334 63.576 210.708 ; 
        RECT 63.04 206.334 63.144 210.708 ; 
        RECT 62.608 206.334 62.712 210.708 ; 
        RECT 62.176 206.334 62.28 210.708 ; 
        RECT 61.744 206.334 61.848 210.708 ; 
        RECT 61.312 206.334 61.416 210.708 ; 
        RECT 60.88 206.334 60.984 210.708 ; 
        RECT 60.448 206.334 60.552 210.708 ; 
        RECT 60.016 206.334 60.12 210.708 ; 
        RECT 59.584 206.334 59.688 210.708 ; 
        RECT 59.152 206.334 59.256 210.708 ; 
        RECT 58.72 206.334 58.824 210.708 ; 
        RECT 58.288 206.334 58.392 210.708 ; 
        RECT 57.856 206.334 57.96 210.708 ; 
        RECT 57.424 206.334 57.528 210.708 ; 
        RECT 56.992 206.334 57.096 210.708 ; 
        RECT 56.56 206.334 56.664 210.708 ; 
        RECT 56.128 206.334 56.232 210.708 ; 
        RECT 55.696 206.334 55.8 210.708 ; 
        RECT 55.264 206.334 55.368 210.708 ; 
        RECT 54.832 206.334 54.936 210.708 ; 
        RECT 54.4 206.334 54.504 210.708 ; 
        RECT 53.968 206.334 54.072 210.708 ; 
        RECT 53.536 206.334 53.64 210.708 ; 
        RECT 53.104 206.334 53.208 210.708 ; 
        RECT 52.672 206.334 52.776 210.708 ; 
        RECT 52.24 206.334 52.344 210.708 ; 
        RECT 51.808 206.334 51.912 210.708 ; 
        RECT 51.376 206.334 51.48 210.708 ; 
        RECT 50.944 206.334 51.048 210.708 ; 
        RECT 50.512 206.334 50.616 210.708 ; 
        RECT 50.08 206.334 50.184 210.708 ; 
        RECT 49.648 206.334 49.752 210.708 ; 
        RECT 49.216 206.334 49.32 210.708 ; 
        RECT 48.784 206.334 48.888 210.708 ; 
        RECT 48.352 206.334 48.456 210.708 ; 
        RECT 47.92 206.334 48.024 210.708 ; 
        RECT 47.488 206.334 47.592 210.708 ; 
        RECT 47.056 206.334 47.16 210.708 ; 
        RECT 46.624 206.334 46.728 210.708 ; 
        RECT 46.192 206.334 46.296 210.708 ; 
        RECT 45.76 206.334 45.864 210.708 ; 
        RECT 45.328 206.334 45.432 210.708 ; 
        RECT 44.896 206.334 45 210.708 ; 
        RECT 44.464 206.334 44.568 210.708 ; 
        RECT 44.032 206.334 44.136 210.708 ; 
        RECT 43.6 206.334 43.704 210.708 ; 
        RECT 43.168 206.334 43.272 210.708 ; 
        RECT 42.736 206.334 42.84 210.708 ; 
        RECT 42.304 206.334 42.408 210.708 ; 
        RECT 41.872 206.334 41.976 210.708 ; 
        RECT 41.44 206.334 41.544 210.708 ; 
        RECT 41.008 206.334 41.112 210.708 ; 
        RECT 40.576 206.334 40.68 210.708 ; 
        RECT 40.144 206.334 40.248 210.708 ; 
        RECT 39.712 206.334 39.816 210.708 ; 
        RECT 39.28 206.334 39.384 210.708 ; 
        RECT 38.848 206.334 38.952 210.708 ; 
        RECT 38.416 206.334 38.52 210.708 ; 
        RECT 37.984 206.334 38.088 210.708 ; 
        RECT 37.552 206.334 37.656 210.708 ; 
        RECT 36.7 206.334 37.008 210.708 ; 
        RECT 29.128 206.334 29.436 210.708 ; 
        RECT 28.48 206.334 28.584 210.708 ; 
        RECT 28.048 206.334 28.152 210.708 ; 
        RECT 27.616 206.334 27.72 210.708 ; 
        RECT 27.184 206.334 27.288 210.708 ; 
        RECT 26.752 206.334 26.856 210.708 ; 
        RECT 26.32 206.334 26.424 210.708 ; 
        RECT 25.888 206.334 25.992 210.708 ; 
        RECT 25.456 206.334 25.56 210.708 ; 
        RECT 25.024 206.334 25.128 210.708 ; 
        RECT 24.592 206.334 24.696 210.708 ; 
        RECT 24.16 206.334 24.264 210.708 ; 
        RECT 23.728 206.334 23.832 210.708 ; 
        RECT 23.296 206.334 23.4 210.708 ; 
        RECT 22.864 206.334 22.968 210.708 ; 
        RECT 22.432 206.334 22.536 210.708 ; 
        RECT 22 206.334 22.104 210.708 ; 
        RECT 21.568 206.334 21.672 210.708 ; 
        RECT 21.136 206.334 21.24 210.708 ; 
        RECT 20.704 206.334 20.808 210.708 ; 
        RECT 20.272 206.334 20.376 210.708 ; 
        RECT 19.84 206.334 19.944 210.708 ; 
        RECT 19.408 206.334 19.512 210.708 ; 
        RECT 18.976 206.334 19.08 210.708 ; 
        RECT 18.544 206.334 18.648 210.708 ; 
        RECT 18.112 206.334 18.216 210.708 ; 
        RECT 17.68 206.334 17.784 210.708 ; 
        RECT 17.248 206.334 17.352 210.708 ; 
        RECT 16.816 206.334 16.92 210.708 ; 
        RECT 16.384 206.334 16.488 210.708 ; 
        RECT 15.952 206.334 16.056 210.708 ; 
        RECT 15.52 206.334 15.624 210.708 ; 
        RECT 15.088 206.334 15.192 210.708 ; 
        RECT 14.656 206.334 14.76 210.708 ; 
        RECT 14.224 206.334 14.328 210.708 ; 
        RECT 13.792 206.334 13.896 210.708 ; 
        RECT 13.36 206.334 13.464 210.708 ; 
        RECT 12.928 206.334 13.032 210.708 ; 
        RECT 12.496 206.334 12.6 210.708 ; 
        RECT 12.064 206.334 12.168 210.708 ; 
        RECT 11.632 206.334 11.736 210.708 ; 
        RECT 11.2 206.334 11.304 210.708 ; 
        RECT 10.768 206.334 10.872 210.708 ; 
        RECT 10.336 206.334 10.44 210.708 ; 
        RECT 9.904 206.334 10.008 210.708 ; 
        RECT 9.472 206.334 9.576 210.708 ; 
        RECT 9.04 206.334 9.144 210.708 ; 
        RECT 8.608 206.334 8.712 210.708 ; 
        RECT 8.176 206.334 8.28 210.708 ; 
        RECT 7.744 206.334 7.848 210.708 ; 
        RECT 7.312 206.334 7.416 210.708 ; 
        RECT 6.88 206.334 6.984 210.708 ; 
        RECT 6.448 206.334 6.552 210.708 ; 
        RECT 6.016 206.334 6.12 210.708 ; 
        RECT 5.584 206.334 5.688 210.708 ; 
        RECT 5.152 206.334 5.256 210.708 ; 
        RECT 4.72 206.334 4.824 210.708 ; 
        RECT 4.288 206.334 4.392 210.708 ; 
        RECT 3.856 206.334 3.96 210.708 ; 
        RECT 3.424 206.334 3.528 210.708 ; 
        RECT 2.992 206.334 3.096 210.708 ; 
        RECT 2.56 206.334 2.664 210.708 ; 
        RECT 2.128 206.334 2.232 210.708 ; 
        RECT 1.696 206.334 1.8 210.708 ; 
        RECT 1.264 206.334 1.368 210.708 ; 
        RECT 0.832 206.334 0.936 210.708 ; 
        RECT 0.02 206.334 0.36 210.708 ; 
        RECT 34.564 210.654 35.076 215.028 ; 
        RECT 34.508 213.316 35.076 214.606 ; 
        RECT 33.916 212.224 34.164 215.028 ; 
        RECT 33.86 213.462 34.164 214.076 ; 
        RECT 33.916 210.654 34.02 215.028 ; 
        RECT 33.916 211.138 34.076 212.096 ; 
        RECT 33.916 210.654 34.164 211.01 ; 
        RECT 32.728 212.456 33.552 215.028 ; 
        RECT 33.448 210.654 33.552 215.028 ; 
        RECT 32.728 213.564 33.608 214.596 ; 
        RECT 32.728 210.654 33.12 215.028 ; 
        RECT 31.06 210.654 31.392 215.028 ; 
        RECT 31.06 211.008 31.448 214.75 ; 
        RECT 65.776 210.654 66.116 215.028 ; 
        RECT 65.2 210.654 65.304 215.028 ; 
        RECT 64.768 210.654 64.872 215.028 ; 
        RECT 64.336 210.654 64.44 215.028 ; 
        RECT 63.904 210.654 64.008 215.028 ; 
        RECT 63.472 210.654 63.576 215.028 ; 
        RECT 63.04 210.654 63.144 215.028 ; 
        RECT 62.608 210.654 62.712 215.028 ; 
        RECT 62.176 210.654 62.28 215.028 ; 
        RECT 61.744 210.654 61.848 215.028 ; 
        RECT 61.312 210.654 61.416 215.028 ; 
        RECT 60.88 210.654 60.984 215.028 ; 
        RECT 60.448 210.654 60.552 215.028 ; 
        RECT 60.016 210.654 60.12 215.028 ; 
        RECT 59.584 210.654 59.688 215.028 ; 
        RECT 59.152 210.654 59.256 215.028 ; 
        RECT 58.72 210.654 58.824 215.028 ; 
        RECT 58.288 210.654 58.392 215.028 ; 
        RECT 57.856 210.654 57.96 215.028 ; 
        RECT 57.424 210.654 57.528 215.028 ; 
        RECT 56.992 210.654 57.096 215.028 ; 
        RECT 56.56 210.654 56.664 215.028 ; 
        RECT 56.128 210.654 56.232 215.028 ; 
        RECT 55.696 210.654 55.8 215.028 ; 
        RECT 55.264 210.654 55.368 215.028 ; 
        RECT 54.832 210.654 54.936 215.028 ; 
        RECT 54.4 210.654 54.504 215.028 ; 
        RECT 53.968 210.654 54.072 215.028 ; 
        RECT 53.536 210.654 53.64 215.028 ; 
        RECT 53.104 210.654 53.208 215.028 ; 
        RECT 52.672 210.654 52.776 215.028 ; 
        RECT 52.24 210.654 52.344 215.028 ; 
        RECT 51.808 210.654 51.912 215.028 ; 
        RECT 51.376 210.654 51.48 215.028 ; 
        RECT 50.944 210.654 51.048 215.028 ; 
        RECT 50.512 210.654 50.616 215.028 ; 
        RECT 50.08 210.654 50.184 215.028 ; 
        RECT 49.648 210.654 49.752 215.028 ; 
        RECT 49.216 210.654 49.32 215.028 ; 
        RECT 48.784 210.654 48.888 215.028 ; 
        RECT 48.352 210.654 48.456 215.028 ; 
        RECT 47.92 210.654 48.024 215.028 ; 
        RECT 47.488 210.654 47.592 215.028 ; 
        RECT 47.056 210.654 47.16 215.028 ; 
        RECT 46.624 210.654 46.728 215.028 ; 
        RECT 46.192 210.654 46.296 215.028 ; 
        RECT 45.76 210.654 45.864 215.028 ; 
        RECT 45.328 210.654 45.432 215.028 ; 
        RECT 44.896 210.654 45 215.028 ; 
        RECT 44.464 210.654 44.568 215.028 ; 
        RECT 44.032 210.654 44.136 215.028 ; 
        RECT 43.6 210.654 43.704 215.028 ; 
        RECT 43.168 210.654 43.272 215.028 ; 
        RECT 42.736 210.654 42.84 215.028 ; 
        RECT 42.304 210.654 42.408 215.028 ; 
        RECT 41.872 210.654 41.976 215.028 ; 
        RECT 41.44 210.654 41.544 215.028 ; 
        RECT 41.008 210.654 41.112 215.028 ; 
        RECT 40.576 210.654 40.68 215.028 ; 
        RECT 40.144 210.654 40.248 215.028 ; 
        RECT 39.712 210.654 39.816 215.028 ; 
        RECT 39.28 210.654 39.384 215.028 ; 
        RECT 38.848 210.654 38.952 215.028 ; 
        RECT 38.416 210.654 38.52 215.028 ; 
        RECT 37.984 210.654 38.088 215.028 ; 
        RECT 37.552 210.654 37.656 215.028 ; 
        RECT 36.7 210.654 37.008 215.028 ; 
        RECT 29.128 210.654 29.436 215.028 ; 
        RECT 28.48 210.654 28.584 215.028 ; 
        RECT 28.048 210.654 28.152 215.028 ; 
        RECT 27.616 210.654 27.72 215.028 ; 
        RECT 27.184 210.654 27.288 215.028 ; 
        RECT 26.752 210.654 26.856 215.028 ; 
        RECT 26.32 210.654 26.424 215.028 ; 
        RECT 25.888 210.654 25.992 215.028 ; 
        RECT 25.456 210.654 25.56 215.028 ; 
        RECT 25.024 210.654 25.128 215.028 ; 
        RECT 24.592 210.654 24.696 215.028 ; 
        RECT 24.16 210.654 24.264 215.028 ; 
        RECT 23.728 210.654 23.832 215.028 ; 
        RECT 23.296 210.654 23.4 215.028 ; 
        RECT 22.864 210.654 22.968 215.028 ; 
        RECT 22.432 210.654 22.536 215.028 ; 
        RECT 22 210.654 22.104 215.028 ; 
        RECT 21.568 210.654 21.672 215.028 ; 
        RECT 21.136 210.654 21.24 215.028 ; 
        RECT 20.704 210.654 20.808 215.028 ; 
        RECT 20.272 210.654 20.376 215.028 ; 
        RECT 19.84 210.654 19.944 215.028 ; 
        RECT 19.408 210.654 19.512 215.028 ; 
        RECT 18.976 210.654 19.08 215.028 ; 
        RECT 18.544 210.654 18.648 215.028 ; 
        RECT 18.112 210.654 18.216 215.028 ; 
        RECT 17.68 210.654 17.784 215.028 ; 
        RECT 17.248 210.654 17.352 215.028 ; 
        RECT 16.816 210.654 16.92 215.028 ; 
        RECT 16.384 210.654 16.488 215.028 ; 
        RECT 15.952 210.654 16.056 215.028 ; 
        RECT 15.52 210.654 15.624 215.028 ; 
        RECT 15.088 210.654 15.192 215.028 ; 
        RECT 14.656 210.654 14.76 215.028 ; 
        RECT 14.224 210.654 14.328 215.028 ; 
        RECT 13.792 210.654 13.896 215.028 ; 
        RECT 13.36 210.654 13.464 215.028 ; 
        RECT 12.928 210.654 13.032 215.028 ; 
        RECT 12.496 210.654 12.6 215.028 ; 
        RECT 12.064 210.654 12.168 215.028 ; 
        RECT 11.632 210.654 11.736 215.028 ; 
        RECT 11.2 210.654 11.304 215.028 ; 
        RECT 10.768 210.654 10.872 215.028 ; 
        RECT 10.336 210.654 10.44 215.028 ; 
        RECT 9.904 210.654 10.008 215.028 ; 
        RECT 9.472 210.654 9.576 215.028 ; 
        RECT 9.04 210.654 9.144 215.028 ; 
        RECT 8.608 210.654 8.712 215.028 ; 
        RECT 8.176 210.654 8.28 215.028 ; 
        RECT 7.744 210.654 7.848 215.028 ; 
        RECT 7.312 210.654 7.416 215.028 ; 
        RECT 6.88 210.654 6.984 215.028 ; 
        RECT 6.448 210.654 6.552 215.028 ; 
        RECT 6.016 210.654 6.12 215.028 ; 
        RECT 5.584 210.654 5.688 215.028 ; 
        RECT 5.152 210.654 5.256 215.028 ; 
        RECT 4.72 210.654 4.824 215.028 ; 
        RECT 4.288 210.654 4.392 215.028 ; 
        RECT 3.856 210.654 3.96 215.028 ; 
        RECT 3.424 210.654 3.528 215.028 ; 
        RECT 2.992 210.654 3.096 215.028 ; 
        RECT 2.56 210.654 2.664 215.028 ; 
        RECT 2.128 210.654 2.232 215.028 ; 
        RECT 1.696 210.654 1.8 215.028 ; 
        RECT 1.264 210.654 1.368 215.028 ; 
        RECT 0.832 210.654 0.936 215.028 ; 
        RECT 0.02 210.654 0.36 215.028 ; 
        RECT 34.564 214.974 35.076 219.348 ; 
        RECT 34.508 217.636 35.076 218.926 ; 
        RECT 33.916 216.544 34.164 219.348 ; 
        RECT 33.86 217.782 34.164 218.396 ; 
        RECT 33.916 214.974 34.02 219.348 ; 
        RECT 33.916 215.458 34.076 216.416 ; 
        RECT 33.916 214.974 34.164 215.33 ; 
        RECT 32.728 216.776 33.552 219.348 ; 
        RECT 33.448 214.974 33.552 219.348 ; 
        RECT 32.728 217.884 33.608 218.916 ; 
        RECT 32.728 214.974 33.12 219.348 ; 
        RECT 31.06 214.974 31.392 219.348 ; 
        RECT 31.06 215.328 31.448 219.07 ; 
        RECT 65.776 214.974 66.116 219.348 ; 
        RECT 65.2 214.974 65.304 219.348 ; 
        RECT 64.768 214.974 64.872 219.348 ; 
        RECT 64.336 214.974 64.44 219.348 ; 
        RECT 63.904 214.974 64.008 219.348 ; 
        RECT 63.472 214.974 63.576 219.348 ; 
        RECT 63.04 214.974 63.144 219.348 ; 
        RECT 62.608 214.974 62.712 219.348 ; 
        RECT 62.176 214.974 62.28 219.348 ; 
        RECT 61.744 214.974 61.848 219.348 ; 
        RECT 61.312 214.974 61.416 219.348 ; 
        RECT 60.88 214.974 60.984 219.348 ; 
        RECT 60.448 214.974 60.552 219.348 ; 
        RECT 60.016 214.974 60.12 219.348 ; 
        RECT 59.584 214.974 59.688 219.348 ; 
        RECT 59.152 214.974 59.256 219.348 ; 
        RECT 58.72 214.974 58.824 219.348 ; 
        RECT 58.288 214.974 58.392 219.348 ; 
        RECT 57.856 214.974 57.96 219.348 ; 
        RECT 57.424 214.974 57.528 219.348 ; 
        RECT 56.992 214.974 57.096 219.348 ; 
        RECT 56.56 214.974 56.664 219.348 ; 
        RECT 56.128 214.974 56.232 219.348 ; 
        RECT 55.696 214.974 55.8 219.348 ; 
        RECT 55.264 214.974 55.368 219.348 ; 
        RECT 54.832 214.974 54.936 219.348 ; 
        RECT 54.4 214.974 54.504 219.348 ; 
        RECT 53.968 214.974 54.072 219.348 ; 
        RECT 53.536 214.974 53.64 219.348 ; 
        RECT 53.104 214.974 53.208 219.348 ; 
        RECT 52.672 214.974 52.776 219.348 ; 
        RECT 52.24 214.974 52.344 219.348 ; 
        RECT 51.808 214.974 51.912 219.348 ; 
        RECT 51.376 214.974 51.48 219.348 ; 
        RECT 50.944 214.974 51.048 219.348 ; 
        RECT 50.512 214.974 50.616 219.348 ; 
        RECT 50.08 214.974 50.184 219.348 ; 
        RECT 49.648 214.974 49.752 219.348 ; 
        RECT 49.216 214.974 49.32 219.348 ; 
        RECT 48.784 214.974 48.888 219.348 ; 
        RECT 48.352 214.974 48.456 219.348 ; 
        RECT 47.92 214.974 48.024 219.348 ; 
        RECT 47.488 214.974 47.592 219.348 ; 
        RECT 47.056 214.974 47.16 219.348 ; 
        RECT 46.624 214.974 46.728 219.348 ; 
        RECT 46.192 214.974 46.296 219.348 ; 
        RECT 45.76 214.974 45.864 219.348 ; 
        RECT 45.328 214.974 45.432 219.348 ; 
        RECT 44.896 214.974 45 219.348 ; 
        RECT 44.464 214.974 44.568 219.348 ; 
        RECT 44.032 214.974 44.136 219.348 ; 
        RECT 43.6 214.974 43.704 219.348 ; 
        RECT 43.168 214.974 43.272 219.348 ; 
        RECT 42.736 214.974 42.84 219.348 ; 
        RECT 42.304 214.974 42.408 219.348 ; 
        RECT 41.872 214.974 41.976 219.348 ; 
        RECT 41.44 214.974 41.544 219.348 ; 
        RECT 41.008 214.974 41.112 219.348 ; 
        RECT 40.576 214.974 40.68 219.348 ; 
        RECT 40.144 214.974 40.248 219.348 ; 
        RECT 39.712 214.974 39.816 219.348 ; 
        RECT 39.28 214.974 39.384 219.348 ; 
        RECT 38.848 214.974 38.952 219.348 ; 
        RECT 38.416 214.974 38.52 219.348 ; 
        RECT 37.984 214.974 38.088 219.348 ; 
        RECT 37.552 214.974 37.656 219.348 ; 
        RECT 36.7 214.974 37.008 219.348 ; 
        RECT 29.128 214.974 29.436 219.348 ; 
        RECT 28.48 214.974 28.584 219.348 ; 
        RECT 28.048 214.974 28.152 219.348 ; 
        RECT 27.616 214.974 27.72 219.348 ; 
        RECT 27.184 214.974 27.288 219.348 ; 
        RECT 26.752 214.974 26.856 219.348 ; 
        RECT 26.32 214.974 26.424 219.348 ; 
        RECT 25.888 214.974 25.992 219.348 ; 
        RECT 25.456 214.974 25.56 219.348 ; 
        RECT 25.024 214.974 25.128 219.348 ; 
        RECT 24.592 214.974 24.696 219.348 ; 
        RECT 24.16 214.974 24.264 219.348 ; 
        RECT 23.728 214.974 23.832 219.348 ; 
        RECT 23.296 214.974 23.4 219.348 ; 
        RECT 22.864 214.974 22.968 219.348 ; 
        RECT 22.432 214.974 22.536 219.348 ; 
        RECT 22 214.974 22.104 219.348 ; 
        RECT 21.568 214.974 21.672 219.348 ; 
        RECT 21.136 214.974 21.24 219.348 ; 
        RECT 20.704 214.974 20.808 219.348 ; 
        RECT 20.272 214.974 20.376 219.348 ; 
        RECT 19.84 214.974 19.944 219.348 ; 
        RECT 19.408 214.974 19.512 219.348 ; 
        RECT 18.976 214.974 19.08 219.348 ; 
        RECT 18.544 214.974 18.648 219.348 ; 
        RECT 18.112 214.974 18.216 219.348 ; 
        RECT 17.68 214.974 17.784 219.348 ; 
        RECT 17.248 214.974 17.352 219.348 ; 
        RECT 16.816 214.974 16.92 219.348 ; 
        RECT 16.384 214.974 16.488 219.348 ; 
        RECT 15.952 214.974 16.056 219.348 ; 
        RECT 15.52 214.974 15.624 219.348 ; 
        RECT 15.088 214.974 15.192 219.348 ; 
        RECT 14.656 214.974 14.76 219.348 ; 
        RECT 14.224 214.974 14.328 219.348 ; 
        RECT 13.792 214.974 13.896 219.348 ; 
        RECT 13.36 214.974 13.464 219.348 ; 
        RECT 12.928 214.974 13.032 219.348 ; 
        RECT 12.496 214.974 12.6 219.348 ; 
        RECT 12.064 214.974 12.168 219.348 ; 
        RECT 11.632 214.974 11.736 219.348 ; 
        RECT 11.2 214.974 11.304 219.348 ; 
        RECT 10.768 214.974 10.872 219.348 ; 
        RECT 10.336 214.974 10.44 219.348 ; 
        RECT 9.904 214.974 10.008 219.348 ; 
        RECT 9.472 214.974 9.576 219.348 ; 
        RECT 9.04 214.974 9.144 219.348 ; 
        RECT 8.608 214.974 8.712 219.348 ; 
        RECT 8.176 214.974 8.28 219.348 ; 
        RECT 7.744 214.974 7.848 219.348 ; 
        RECT 7.312 214.974 7.416 219.348 ; 
        RECT 6.88 214.974 6.984 219.348 ; 
        RECT 6.448 214.974 6.552 219.348 ; 
        RECT 6.016 214.974 6.12 219.348 ; 
        RECT 5.584 214.974 5.688 219.348 ; 
        RECT 5.152 214.974 5.256 219.348 ; 
        RECT 4.72 214.974 4.824 219.348 ; 
        RECT 4.288 214.974 4.392 219.348 ; 
        RECT 3.856 214.974 3.96 219.348 ; 
        RECT 3.424 214.974 3.528 219.348 ; 
        RECT 2.992 214.974 3.096 219.348 ; 
        RECT 2.56 214.974 2.664 219.348 ; 
        RECT 2.128 214.974 2.232 219.348 ; 
        RECT 1.696 214.974 1.8 219.348 ; 
        RECT 1.264 214.974 1.368 219.348 ; 
        RECT 0.832 214.974 0.936 219.348 ; 
        RECT 0.02 214.974 0.36 219.348 ; 
        RECT 34.564 219.294 35.076 223.668 ; 
        RECT 34.508 221.956 35.076 223.246 ; 
        RECT 33.916 220.864 34.164 223.668 ; 
        RECT 33.86 222.102 34.164 222.716 ; 
        RECT 33.916 219.294 34.02 223.668 ; 
        RECT 33.916 219.778 34.076 220.736 ; 
        RECT 33.916 219.294 34.164 219.65 ; 
        RECT 32.728 221.096 33.552 223.668 ; 
        RECT 33.448 219.294 33.552 223.668 ; 
        RECT 32.728 222.204 33.608 223.236 ; 
        RECT 32.728 219.294 33.12 223.668 ; 
        RECT 31.06 219.294 31.392 223.668 ; 
        RECT 31.06 219.648 31.448 223.39 ; 
        RECT 65.776 219.294 66.116 223.668 ; 
        RECT 65.2 219.294 65.304 223.668 ; 
        RECT 64.768 219.294 64.872 223.668 ; 
        RECT 64.336 219.294 64.44 223.668 ; 
        RECT 63.904 219.294 64.008 223.668 ; 
        RECT 63.472 219.294 63.576 223.668 ; 
        RECT 63.04 219.294 63.144 223.668 ; 
        RECT 62.608 219.294 62.712 223.668 ; 
        RECT 62.176 219.294 62.28 223.668 ; 
        RECT 61.744 219.294 61.848 223.668 ; 
        RECT 61.312 219.294 61.416 223.668 ; 
        RECT 60.88 219.294 60.984 223.668 ; 
        RECT 60.448 219.294 60.552 223.668 ; 
        RECT 60.016 219.294 60.12 223.668 ; 
        RECT 59.584 219.294 59.688 223.668 ; 
        RECT 59.152 219.294 59.256 223.668 ; 
        RECT 58.72 219.294 58.824 223.668 ; 
        RECT 58.288 219.294 58.392 223.668 ; 
        RECT 57.856 219.294 57.96 223.668 ; 
        RECT 57.424 219.294 57.528 223.668 ; 
        RECT 56.992 219.294 57.096 223.668 ; 
        RECT 56.56 219.294 56.664 223.668 ; 
        RECT 56.128 219.294 56.232 223.668 ; 
        RECT 55.696 219.294 55.8 223.668 ; 
        RECT 55.264 219.294 55.368 223.668 ; 
        RECT 54.832 219.294 54.936 223.668 ; 
        RECT 54.4 219.294 54.504 223.668 ; 
        RECT 53.968 219.294 54.072 223.668 ; 
        RECT 53.536 219.294 53.64 223.668 ; 
        RECT 53.104 219.294 53.208 223.668 ; 
        RECT 52.672 219.294 52.776 223.668 ; 
        RECT 52.24 219.294 52.344 223.668 ; 
        RECT 51.808 219.294 51.912 223.668 ; 
        RECT 51.376 219.294 51.48 223.668 ; 
        RECT 50.944 219.294 51.048 223.668 ; 
        RECT 50.512 219.294 50.616 223.668 ; 
        RECT 50.08 219.294 50.184 223.668 ; 
        RECT 49.648 219.294 49.752 223.668 ; 
        RECT 49.216 219.294 49.32 223.668 ; 
        RECT 48.784 219.294 48.888 223.668 ; 
        RECT 48.352 219.294 48.456 223.668 ; 
        RECT 47.92 219.294 48.024 223.668 ; 
        RECT 47.488 219.294 47.592 223.668 ; 
        RECT 47.056 219.294 47.16 223.668 ; 
        RECT 46.624 219.294 46.728 223.668 ; 
        RECT 46.192 219.294 46.296 223.668 ; 
        RECT 45.76 219.294 45.864 223.668 ; 
        RECT 45.328 219.294 45.432 223.668 ; 
        RECT 44.896 219.294 45 223.668 ; 
        RECT 44.464 219.294 44.568 223.668 ; 
        RECT 44.032 219.294 44.136 223.668 ; 
        RECT 43.6 219.294 43.704 223.668 ; 
        RECT 43.168 219.294 43.272 223.668 ; 
        RECT 42.736 219.294 42.84 223.668 ; 
        RECT 42.304 219.294 42.408 223.668 ; 
        RECT 41.872 219.294 41.976 223.668 ; 
        RECT 41.44 219.294 41.544 223.668 ; 
        RECT 41.008 219.294 41.112 223.668 ; 
        RECT 40.576 219.294 40.68 223.668 ; 
        RECT 40.144 219.294 40.248 223.668 ; 
        RECT 39.712 219.294 39.816 223.668 ; 
        RECT 39.28 219.294 39.384 223.668 ; 
        RECT 38.848 219.294 38.952 223.668 ; 
        RECT 38.416 219.294 38.52 223.668 ; 
        RECT 37.984 219.294 38.088 223.668 ; 
        RECT 37.552 219.294 37.656 223.668 ; 
        RECT 36.7 219.294 37.008 223.668 ; 
        RECT 29.128 219.294 29.436 223.668 ; 
        RECT 28.48 219.294 28.584 223.668 ; 
        RECT 28.048 219.294 28.152 223.668 ; 
        RECT 27.616 219.294 27.72 223.668 ; 
        RECT 27.184 219.294 27.288 223.668 ; 
        RECT 26.752 219.294 26.856 223.668 ; 
        RECT 26.32 219.294 26.424 223.668 ; 
        RECT 25.888 219.294 25.992 223.668 ; 
        RECT 25.456 219.294 25.56 223.668 ; 
        RECT 25.024 219.294 25.128 223.668 ; 
        RECT 24.592 219.294 24.696 223.668 ; 
        RECT 24.16 219.294 24.264 223.668 ; 
        RECT 23.728 219.294 23.832 223.668 ; 
        RECT 23.296 219.294 23.4 223.668 ; 
        RECT 22.864 219.294 22.968 223.668 ; 
        RECT 22.432 219.294 22.536 223.668 ; 
        RECT 22 219.294 22.104 223.668 ; 
        RECT 21.568 219.294 21.672 223.668 ; 
        RECT 21.136 219.294 21.24 223.668 ; 
        RECT 20.704 219.294 20.808 223.668 ; 
        RECT 20.272 219.294 20.376 223.668 ; 
        RECT 19.84 219.294 19.944 223.668 ; 
        RECT 19.408 219.294 19.512 223.668 ; 
        RECT 18.976 219.294 19.08 223.668 ; 
        RECT 18.544 219.294 18.648 223.668 ; 
        RECT 18.112 219.294 18.216 223.668 ; 
        RECT 17.68 219.294 17.784 223.668 ; 
        RECT 17.248 219.294 17.352 223.668 ; 
        RECT 16.816 219.294 16.92 223.668 ; 
        RECT 16.384 219.294 16.488 223.668 ; 
        RECT 15.952 219.294 16.056 223.668 ; 
        RECT 15.52 219.294 15.624 223.668 ; 
        RECT 15.088 219.294 15.192 223.668 ; 
        RECT 14.656 219.294 14.76 223.668 ; 
        RECT 14.224 219.294 14.328 223.668 ; 
        RECT 13.792 219.294 13.896 223.668 ; 
        RECT 13.36 219.294 13.464 223.668 ; 
        RECT 12.928 219.294 13.032 223.668 ; 
        RECT 12.496 219.294 12.6 223.668 ; 
        RECT 12.064 219.294 12.168 223.668 ; 
        RECT 11.632 219.294 11.736 223.668 ; 
        RECT 11.2 219.294 11.304 223.668 ; 
        RECT 10.768 219.294 10.872 223.668 ; 
        RECT 10.336 219.294 10.44 223.668 ; 
        RECT 9.904 219.294 10.008 223.668 ; 
        RECT 9.472 219.294 9.576 223.668 ; 
        RECT 9.04 219.294 9.144 223.668 ; 
        RECT 8.608 219.294 8.712 223.668 ; 
        RECT 8.176 219.294 8.28 223.668 ; 
        RECT 7.744 219.294 7.848 223.668 ; 
        RECT 7.312 219.294 7.416 223.668 ; 
        RECT 6.88 219.294 6.984 223.668 ; 
        RECT 6.448 219.294 6.552 223.668 ; 
        RECT 6.016 219.294 6.12 223.668 ; 
        RECT 5.584 219.294 5.688 223.668 ; 
        RECT 5.152 219.294 5.256 223.668 ; 
        RECT 4.72 219.294 4.824 223.668 ; 
        RECT 4.288 219.294 4.392 223.668 ; 
        RECT 3.856 219.294 3.96 223.668 ; 
        RECT 3.424 219.294 3.528 223.668 ; 
        RECT 2.992 219.294 3.096 223.668 ; 
        RECT 2.56 219.294 2.664 223.668 ; 
        RECT 2.128 219.294 2.232 223.668 ; 
        RECT 1.696 219.294 1.8 223.668 ; 
        RECT 1.264 219.294 1.368 223.668 ; 
        RECT 0.832 219.294 0.936 223.668 ; 
        RECT 0.02 219.294 0.36 223.668 ; 
        RECT 34.564 223.614 35.076 227.988 ; 
        RECT 34.508 226.276 35.076 227.566 ; 
        RECT 33.916 225.184 34.164 227.988 ; 
        RECT 33.86 226.422 34.164 227.036 ; 
        RECT 33.916 223.614 34.02 227.988 ; 
        RECT 33.916 224.098 34.076 225.056 ; 
        RECT 33.916 223.614 34.164 223.97 ; 
        RECT 32.728 225.416 33.552 227.988 ; 
        RECT 33.448 223.614 33.552 227.988 ; 
        RECT 32.728 226.524 33.608 227.556 ; 
        RECT 32.728 223.614 33.12 227.988 ; 
        RECT 31.06 223.614 31.392 227.988 ; 
        RECT 31.06 223.968 31.448 227.71 ; 
        RECT 65.776 223.614 66.116 227.988 ; 
        RECT 65.2 223.614 65.304 227.988 ; 
        RECT 64.768 223.614 64.872 227.988 ; 
        RECT 64.336 223.614 64.44 227.988 ; 
        RECT 63.904 223.614 64.008 227.988 ; 
        RECT 63.472 223.614 63.576 227.988 ; 
        RECT 63.04 223.614 63.144 227.988 ; 
        RECT 62.608 223.614 62.712 227.988 ; 
        RECT 62.176 223.614 62.28 227.988 ; 
        RECT 61.744 223.614 61.848 227.988 ; 
        RECT 61.312 223.614 61.416 227.988 ; 
        RECT 60.88 223.614 60.984 227.988 ; 
        RECT 60.448 223.614 60.552 227.988 ; 
        RECT 60.016 223.614 60.12 227.988 ; 
        RECT 59.584 223.614 59.688 227.988 ; 
        RECT 59.152 223.614 59.256 227.988 ; 
        RECT 58.72 223.614 58.824 227.988 ; 
        RECT 58.288 223.614 58.392 227.988 ; 
        RECT 57.856 223.614 57.96 227.988 ; 
        RECT 57.424 223.614 57.528 227.988 ; 
        RECT 56.992 223.614 57.096 227.988 ; 
        RECT 56.56 223.614 56.664 227.988 ; 
        RECT 56.128 223.614 56.232 227.988 ; 
        RECT 55.696 223.614 55.8 227.988 ; 
        RECT 55.264 223.614 55.368 227.988 ; 
        RECT 54.832 223.614 54.936 227.988 ; 
        RECT 54.4 223.614 54.504 227.988 ; 
        RECT 53.968 223.614 54.072 227.988 ; 
        RECT 53.536 223.614 53.64 227.988 ; 
        RECT 53.104 223.614 53.208 227.988 ; 
        RECT 52.672 223.614 52.776 227.988 ; 
        RECT 52.24 223.614 52.344 227.988 ; 
        RECT 51.808 223.614 51.912 227.988 ; 
        RECT 51.376 223.614 51.48 227.988 ; 
        RECT 50.944 223.614 51.048 227.988 ; 
        RECT 50.512 223.614 50.616 227.988 ; 
        RECT 50.08 223.614 50.184 227.988 ; 
        RECT 49.648 223.614 49.752 227.988 ; 
        RECT 49.216 223.614 49.32 227.988 ; 
        RECT 48.784 223.614 48.888 227.988 ; 
        RECT 48.352 223.614 48.456 227.988 ; 
        RECT 47.92 223.614 48.024 227.988 ; 
        RECT 47.488 223.614 47.592 227.988 ; 
        RECT 47.056 223.614 47.16 227.988 ; 
        RECT 46.624 223.614 46.728 227.988 ; 
        RECT 46.192 223.614 46.296 227.988 ; 
        RECT 45.76 223.614 45.864 227.988 ; 
        RECT 45.328 223.614 45.432 227.988 ; 
        RECT 44.896 223.614 45 227.988 ; 
        RECT 44.464 223.614 44.568 227.988 ; 
        RECT 44.032 223.614 44.136 227.988 ; 
        RECT 43.6 223.614 43.704 227.988 ; 
        RECT 43.168 223.614 43.272 227.988 ; 
        RECT 42.736 223.614 42.84 227.988 ; 
        RECT 42.304 223.614 42.408 227.988 ; 
        RECT 41.872 223.614 41.976 227.988 ; 
        RECT 41.44 223.614 41.544 227.988 ; 
        RECT 41.008 223.614 41.112 227.988 ; 
        RECT 40.576 223.614 40.68 227.988 ; 
        RECT 40.144 223.614 40.248 227.988 ; 
        RECT 39.712 223.614 39.816 227.988 ; 
        RECT 39.28 223.614 39.384 227.988 ; 
        RECT 38.848 223.614 38.952 227.988 ; 
        RECT 38.416 223.614 38.52 227.988 ; 
        RECT 37.984 223.614 38.088 227.988 ; 
        RECT 37.552 223.614 37.656 227.988 ; 
        RECT 36.7 223.614 37.008 227.988 ; 
        RECT 29.128 223.614 29.436 227.988 ; 
        RECT 28.48 223.614 28.584 227.988 ; 
        RECT 28.048 223.614 28.152 227.988 ; 
        RECT 27.616 223.614 27.72 227.988 ; 
        RECT 27.184 223.614 27.288 227.988 ; 
        RECT 26.752 223.614 26.856 227.988 ; 
        RECT 26.32 223.614 26.424 227.988 ; 
        RECT 25.888 223.614 25.992 227.988 ; 
        RECT 25.456 223.614 25.56 227.988 ; 
        RECT 25.024 223.614 25.128 227.988 ; 
        RECT 24.592 223.614 24.696 227.988 ; 
        RECT 24.16 223.614 24.264 227.988 ; 
        RECT 23.728 223.614 23.832 227.988 ; 
        RECT 23.296 223.614 23.4 227.988 ; 
        RECT 22.864 223.614 22.968 227.988 ; 
        RECT 22.432 223.614 22.536 227.988 ; 
        RECT 22 223.614 22.104 227.988 ; 
        RECT 21.568 223.614 21.672 227.988 ; 
        RECT 21.136 223.614 21.24 227.988 ; 
        RECT 20.704 223.614 20.808 227.988 ; 
        RECT 20.272 223.614 20.376 227.988 ; 
        RECT 19.84 223.614 19.944 227.988 ; 
        RECT 19.408 223.614 19.512 227.988 ; 
        RECT 18.976 223.614 19.08 227.988 ; 
        RECT 18.544 223.614 18.648 227.988 ; 
        RECT 18.112 223.614 18.216 227.988 ; 
        RECT 17.68 223.614 17.784 227.988 ; 
        RECT 17.248 223.614 17.352 227.988 ; 
        RECT 16.816 223.614 16.92 227.988 ; 
        RECT 16.384 223.614 16.488 227.988 ; 
        RECT 15.952 223.614 16.056 227.988 ; 
        RECT 15.52 223.614 15.624 227.988 ; 
        RECT 15.088 223.614 15.192 227.988 ; 
        RECT 14.656 223.614 14.76 227.988 ; 
        RECT 14.224 223.614 14.328 227.988 ; 
        RECT 13.792 223.614 13.896 227.988 ; 
        RECT 13.36 223.614 13.464 227.988 ; 
        RECT 12.928 223.614 13.032 227.988 ; 
        RECT 12.496 223.614 12.6 227.988 ; 
        RECT 12.064 223.614 12.168 227.988 ; 
        RECT 11.632 223.614 11.736 227.988 ; 
        RECT 11.2 223.614 11.304 227.988 ; 
        RECT 10.768 223.614 10.872 227.988 ; 
        RECT 10.336 223.614 10.44 227.988 ; 
        RECT 9.904 223.614 10.008 227.988 ; 
        RECT 9.472 223.614 9.576 227.988 ; 
        RECT 9.04 223.614 9.144 227.988 ; 
        RECT 8.608 223.614 8.712 227.988 ; 
        RECT 8.176 223.614 8.28 227.988 ; 
        RECT 7.744 223.614 7.848 227.988 ; 
        RECT 7.312 223.614 7.416 227.988 ; 
        RECT 6.88 223.614 6.984 227.988 ; 
        RECT 6.448 223.614 6.552 227.988 ; 
        RECT 6.016 223.614 6.12 227.988 ; 
        RECT 5.584 223.614 5.688 227.988 ; 
        RECT 5.152 223.614 5.256 227.988 ; 
        RECT 4.72 223.614 4.824 227.988 ; 
        RECT 4.288 223.614 4.392 227.988 ; 
        RECT 3.856 223.614 3.96 227.988 ; 
        RECT 3.424 223.614 3.528 227.988 ; 
        RECT 2.992 223.614 3.096 227.988 ; 
        RECT 2.56 223.614 2.664 227.988 ; 
        RECT 2.128 223.614 2.232 227.988 ; 
        RECT 1.696 223.614 1.8 227.988 ; 
        RECT 1.264 223.614 1.368 227.988 ; 
        RECT 0.832 223.614 0.936 227.988 ; 
        RECT 0.02 223.614 0.36 227.988 ; 
        RECT 34.564 227.934 35.076 232.308 ; 
        RECT 34.508 230.596 35.076 231.886 ; 
        RECT 33.916 229.504 34.164 232.308 ; 
        RECT 33.86 230.742 34.164 231.356 ; 
        RECT 33.916 227.934 34.02 232.308 ; 
        RECT 33.916 228.418 34.076 229.376 ; 
        RECT 33.916 227.934 34.164 228.29 ; 
        RECT 32.728 229.736 33.552 232.308 ; 
        RECT 33.448 227.934 33.552 232.308 ; 
        RECT 32.728 230.844 33.608 231.876 ; 
        RECT 32.728 227.934 33.12 232.308 ; 
        RECT 31.06 227.934 31.392 232.308 ; 
        RECT 31.06 228.288 31.448 232.03 ; 
        RECT 65.776 227.934 66.116 232.308 ; 
        RECT 65.2 227.934 65.304 232.308 ; 
        RECT 64.768 227.934 64.872 232.308 ; 
        RECT 64.336 227.934 64.44 232.308 ; 
        RECT 63.904 227.934 64.008 232.308 ; 
        RECT 63.472 227.934 63.576 232.308 ; 
        RECT 63.04 227.934 63.144 232.308 ; 
        RECT 62.608 227.934 62.712 232.308 ; 
        RECT 62.176 227.934 62.28 232.308 ; 
        RECT 61.744 227.934 61.848 232.308 ; 
        RECT 61.312 227.934 61.416 232.308 ; 
        RECT 60.88 227.934 60.984 232.308 ; 
        RECT 60.448 227.934 60.552 232.308 ; 
        RECT 60.016 227.934 60.12 232.308 ; 
        RECT 59.584 227.934 59.688 232.308 ; 
        RECT 59.152 227.934 59.256 232.308 ; 
        RECT 58.72 227.934 58.824 232.308 ; 
        RECT 58.288 227.934 58.392 232.308 ; 
        RECT 57.856 227.934 57.96 232.308 ; 
        RECT 57.424 227.934 57.528 232.308 ; 
        RECT 56.992 227.934 57.096 232.308 ; 
        RECT 56.56 227.934 56.664 232.308 ; 
        RECT 56.128 227.934 56.232 232.308 ; 
        RECT 55.696 227.934 55.8 232.308 ; 
        RECT 55.264 227.934 55.368 232.308 ; 
        RECT 54.832 227.934 54.936 232.308 ; 
        RECT 54.4 227.934 54.504 232.308 ; 
        RECT 53.968 227.934 54.072 232.308 ; 
        RECT 53.536 227.934 53.64 232.308 ; 
        RECT 53.104 227.934 53.208 232.308 ; 
        RECT 52.672 227.934 52.776 232.308 ; 
        RECT 52.24 227.934 52.344 232.308 ; 
        RECT 51.808 227.934 51.912 232.308 ; 
        RECT 51.376 227.934 51.48 232.308 ; 
        RECT 50.944 227.934 51.048 232.308 ; 
        RECT 50.512 227.934 50.616 232.308 ; 
        RECT 50.08 227.934 50.184 232.308 ; 
        RECT 49.648 227.934 49.752 232.308 ; 
        RECT 49.216 227.934 49.32 232.308 ; 
        RECT 48.784 227.934 48.888 232.308 ; 
        RECT 48.352 227.934 48.456 232.308 ; 
        RECT 47.92 227.934 48.024 232.308 ; 
        RECT 47.488 227.934 47.592 232.308 ; 
        RECT 47.056 227.934 47.16 232.308 ; 
        RECT 46.624 227.934 46.728 232.308 ; 
        RECT 46.192 227.934 46.296 232.308 ; 
        RECT 45.76 227.934 45.864 232.308 ; 
        RECT 45.328 227.934 45.432 232.308 ; 
        RECT 44.896 227.934 45 232.308 ; 
        RECT 44.464 227.934 44.568 232.308 ; 
        RECT 44.032 227.934 44.136 232.308 ; 
        RECT 43.6 227.934 43.704 232.308 ; 
        RECT 43.168 227.934 43.272 232.308 ; 
        RECT 42.736 227.934 42.84 232.308 ; 
        RECT 42.304 227.934 42.408 232.308 ; 
        RECT 41.872 227.934 41.976 232.308 ; 
        RECT 41.44 227.934 41.544 232.308 ; 
        RECT 41.008 227.934 41.112 232.308 ; 
        RECT 40.576 227.934 40.68 232.308 ; 
        RECT 40.144 227.934 40.248 232.308 ; 
        RECT 39.712 227.934 39.816 232.308 ; 
        RECT 39.28 227.934 39.384 232.308 ; 
        RECT 38.848 227.934 38.952 232.308 ; 
        RECT 38.416 227.934 38.52 232.308 ; 
        RECT 37.984 227.934 38.088 232.308 ; 
        RECT 37.552 227.934 37.656 232.308 ; 
        RECT 36.7 227.934 37.008 232.308 ; 
        RECT 29.128 227.934 29.436 232.308 ; 
        RECT 28.48 227.934 28.584 232.308 ; 
        RECT 28.048 227.934 28.152 232.308 ; 
        RECT 27.616 227.934 27.72 232.308 ; 
        RECT 27.184 227.934 27.288 232.308 ; 
        RECT 26.752 227.934 26.856 232.308 ; 
        RECT 26.32 227.934 26.424 232.308 ; 
        RECT 25.888 227.934 25.992 232.308 ; 
        RECT 25.456 227.934 25.56 232.308 ; 
        RECT 25.024 227.934 25.128 232.308 ; 
        RECT 24.592 227.934 24.696 232.308 ; 
        RECT 24.16 227.934 24.264 232.308 ; 
        RECT 23.728 227.934 23.832 232.308 ; 
        RECT 23.296 227.934 23.4 232.308 ; 
        RECT 22.864 227.934 22.968 232.308 ; 
        RECT 22.432 227.934 22.536 232.308 ; 
        RECT 22 227.934 22.104 232.308 ; 
        RECT 21.568 227.934 21.672 232.308 ; 
        RECT 21.136 227.934 21.24 232.308 ; 
        RECT 20.704 227.934 20.808 232.308 ; 
        RECT 20.272 227.934 20.376 232.308 ; 
        RECT 19.84 227.934 19.944 232.308 ; 
        RECT 19.408 227.934 19.512 232.308 ; 
        RECT 18.976 227.934 19.08 232.308 ; 
        RECT 18.544 227.934 18.648 232.308 ; 
        RECT 18.112 227.934 18.216 232.308 ; 
        RECT 17.68 227.934 17.784 232.308 ; 
        RECT 17.248 227.934 17.352 232.308 ; 
        RECT 16.816 227.934 16.92 232.308 ; 
        RECT 16.384 227.934 16.488 232.308 ; 
        RECT 15.952 227.934 16.056 232.308 ; 
        RECT 15.52 227.934 15.624 232.308 ; 
        RECT 15.088 227.934 15.192 232.308 ; 
        RECT 14.656 227.934 14.76 232.308 ; 
        RECT 14.224 227.934 14.328 232.308 ; 
        RECT 13.792 227.934 13.896 232.308 ; 
        RECT 13.36 227.934 13.464 232.308 ; 
        RECT 12.928 227.934 13.032 232.308 ; 
        RECT 12.496 227.934 12.6 232.308 ; 
        RECT 12.064 227.934 12.168 232.308 ; 
        RECT 11.632 227.934 11.736 232.308 ; 
        RECT 11.2 227.934 11.304 232.308 ; 
        RECT 10.768 227.934 10.872 232.308 ; 
        RECT 10.336 227.934 10.44 232.308 ; 
        RECT 9.904 227.934 10.008 232.308 ; 
        RECT 9.472 227.934 9.576 232.308 ; 
        RECT 9.04 227.934 9.144 232.308 ; 
        RECT 8.608 227.934 8.712 232.308 ; 
        RECT 8.176 227.934 8.28 232.308 ; 
        RECT 7.744 227.934 7.848 232.308 ; 
        RECT 7.312 227.934 7.416 232.308 ; 
        RECT 6.88 227.934 6.984 232.308 ; 
        RECT 6.448 227.934 6.552 232.308 ; 
        RECT 6.016 227.934 6.12 232.308 ; 
        RECT 5.584 227.934 5.688 232.308 ; 
        RECT 5.152 227.934 5.256 232.308 ; 
        RECT 4.72 227.934 4.824 232.308 ; 
        RECT 4.288 227.934 4.392 232.308 ; 
        RECT 3.856 227.934 3.96 232.308 ; 
        RECT 3.424 227.934 3.528 232.308 ; 
        RECT 2.992 227.934 3.096 232.308 ; 
        RECT 2.56 227.934 2.664 232.308 ; 
        RECT 2.128 227.934 2.232 232.308 ; 
        RECT 1.696 227.934 1.8 232.308 ; 
        RECT 1.264 227.934 1.368 232.308 ; 
        RECT 0.832 227.934 0.936 232.308 ; 
        RECT 0.02 227.934 0.36 232.308 ; 
        RECT 34.564 232.254 35.076 236.628 ; 
        RECT 34.508 234.916 35.076 236.206 ; 
        RECT 33.916 233.824 34.164 236.628 ; 
        RECT 33.86 235.062 34.164 235.676 ; 
        RECT 33.916 232.254 34.02 236.628 ; 
        RECT 33.916 232.738 34.076 233.696 ; 
        RECT 33.916 232.254 34.164 232.61 ; 
        RECT 32.728 234.056 33.552 236.628 ; 
        RECT 33.448 232.254 33.552 236.628 ; 
        RECT 32.728 235.164 33.608 236.196 ; 
        RECT 32.728 232.254 33.12 236.628 ; 
        RECT 31.06 232.254 31.392 236.628 ; 
        RECT 31.06 232.608 31.448 236.35 ; 
        RECT 65.776 232.254 66.116 236.628 ; 
        RECT 65.2 232.254 65.304 236.628 ; 
        RECT 64.768 232.254 64.872 236.628 ; 
        RECT 64.336 232.254 64.44 236.628 ; 
        RECT 63.904 232.254 64.008 236.628 ; 
        RECT 63.472 232.254 63.576 236.628 ; 
        RECT 63.04 232.254 63.144 236.628 ; 
        RECT 62.608 232.254 62.712 236.628 ; 
        RECT 62.176 232.254 62.28 236.628 ; 
        RECT 61.744 232.254 61.848 236.628 ; 
        RECT 61.312 232.254 61.416 236.628 ; 
        RECT 60.88 232.254 60.984 236.628 ; 
        RECT 60.448 232.254 60.552 236.628 ; 
        RECT 60.016 232.254 60.12 236.628 ; 
        RECT 59.584 232.254 59.688 236.628 ; 
        RECT 59.152 232.254 59.256 236.628 ; 
        RECT 58.72 232.254 58.824 236.628 ; 
        RECT 58.288 232.254 58.392 236.628 ; 
        RECT 57.856 232.254 57.96 236.628 ; 
        RECT 57.424 232.254 57.528 236.628 ; 
        RECT 56.992 232.254 57.096 236.628 ; 
        RECT 56.56 232.254 56.664 236.628 ; 
        RECT 56.128 232.254 56.232 236.628 ; 
        RECT 55.696 232.254 55.8 236.628 ; 
        RECT 55.264 232.254 55.368 236.628 ; 
        RECT 54.832 232.254 54.936 236.628 ; 
        RECT 54.4 232.254 54.504 236.628 ; 
        RECT 53.968 232.254 54.072 236.628 ; 
        RECT 53.536 232.254 53.64 236.628 ; 
        RECT 53.104 232.254 53.208 236.628 ; 
        RECT 52.672 232.254 52.776 236.628 ; 
        RECT 52.24 232.254 52.344 236.628 ; 
        RECT 51.808 232.254 51.912 236.628 ; 
        RECT 51.376 232.254 51.48 236.628 ; 
        RECT 50.944 232.254 51.048 236.628 ; 
        RECT 50.512 232.254 50.616 236.628 ; 
        RECT 50.08 232.254 50.184 236.628 ; 
        RECT 49.648 232.254 49.752 236.628 ; 
        RECT 49.216 232.254 49.32 236.628 ; 
        RECT 48.784 232.254 48.888 236.628 ; 
        RECT 48.352 232.254 48.456 236.628 ; 
        RECT 47.92 232.254 48.024 236.628 ; 
        RECT 47.488 232.254 47.592 236.628 ; 
        RECT 47.056 232.254 47.16 236.628 ; 
        RECT 46.624 232.254 46.728 236.628 ; 
        RECT 46.192 232.254 46.296 236.628 ; 
        RECT 45.76 232.254 45.864 236.628 ; 
        RECT 45.328 232.254 45.432 236.628 ; 
        RECT 44.896 232.254 45 236.628 ; 
        RECT 44.464 232.254 44.568 236.628 ; 
        RECT 44.032 232.254 44.136 236.628 ; 
        RECT 43.6 232.254 43.704 236.628 ; 
        RECT 43.168 232.254 43.272 236.628 ; 
        RECT 42.736 232.254 42.84 236.628 ; 
        RECT 42.304 232.254 42.408 236.628 ; 
        RECT 41.872 232.254 41.976 236.628 ; 
        RECT 41.44 232.254 41.544 236.628 ; 
        RECT 41.008 232.254 41.112 236.628 ; 
        RECT 40.576 232.254 40.68 236.628 ; 
        RECT 40.144 232.254 40.248 236.628 ; 
        RECT 39.712 232.254 39.816 236.628 ; 
        RECT 39.28 232.254 39.384 236.628 ; 
        RECT 38.848 232.254 38.952 236.628 ; 
        RECT 38.416 232.254 38.52 236.628 ; 
        RECT 37.984 232.254 38.088 236.628 ; 
        RECT 37.552 232.254 37.656 236.628 ; 
        RECT 36.7 232.254 37.008 236.628 ; 
        RECT 29.128 232.254 29.436 236.628 ; 
        RECT 28.48 232.254 28.584 236.628 ; 
        RECT 28.048 232.254 28.152 236.628 ; 
        RECT 27.616 232.254 27.72 236.628 ; 
        RECT 27.184 232.254 27.288 236.628 ; 
        RECT 26.752 232.254 26.856 236.628 ; 
        RECT 26.32 232.254 26.424 236.628 ; 
        RECT 25.888 232.254 25.992 236.628 ; 
        RECT 25.456 232.254 25.56 236.628 ; 
        RECT 25.024 232.254 25.128 236.628 ; 
        RECT 24.592 232.254 24.696 236.628 ; 
        RECT 24.16 232.254 24.264 236.628 ; 
        RECT 23.728 232.254 23.832 236.628 ; 
        RECT 23.296 232.254 23.4 236.628 ; 
        RECT 22.864 232.254 22.968 236.628 ; 
        RECT 22.432 232.254 22.536 236.628 ; 
        RECT 22 232.254 22.104 236.628 ; 
        RECT 21.568 232.254 21.672 236.628 ; 
        RECT 21.136 232.254 21.24 236.628 ; 
        RECT 20.704 232.254 20.808 236.628 ; 
        RECT 20.272 232.254 20.376 236.628 ; 
        RECT 19.84 232.254 19.944 236.628 ; 
        RECT 19.408 232.254 19.512 236.628 ; 
        RECT 18.976 232.254 19.08 236.628 ; 
        RECT 18.544 232.254 18.648 236.628 ; 
        RECT 18.112 232.254 18.216 236.628 ; 
        RECT 17.68 232.254 17.784 236.628 ; 
        RECT 17.248 232.254 17.352 236.628 ; 
        RECT 16.816 232.254 16.92 236.628 ; 
        RECT 16.384 232.254 16.488 236.628 ; 
        RECT 15.952 232.254 16.056 236.628 ; 
        RECT 15.52 232.254 15.624 236.628 ; 
        RECT 15.088 232.254 15.192 236.628 ; 
        RECT 14.656 232.254 14.76 236.628 ; 
        RECT 14.224 232.254 14.328 236.628 ; 
        RECT 13.792 232.254 13.896 236.628 ; 
        RECT 13.36 232.254 13.464 236.628 ; 
        RECT 12.928 232.254 13.032 236.628 ; 
        RECT 12.496 232.254 12.6 236.628 ; 
        RECT 12.064 232.254 12.168 236.628 ; 
        RECT 11.632 232.254 11.736 236.628 ; 
        RECT 11.2 232.254 11.304 236.628 ; 
        RECT 10.768 232.254 10.872 236.628 ; 
        RECT 10.336 232.254 10.44 236.628 ; 
        RECT 9.904 232.254 10.008 236.628 ; 
        RECT 9.472 232.254 9.576 236.628 ; 
        RECT 9.04 232.254 9.144 236.628 ; 
        RECT 8.608 232.254 8.712 236.628 ; 
        RECT 8.176 232.254 8.28 236.628 ; 
        RECT 7.744 232.254 7.848 236.628 ; 
        RECT 7.312 232.254 7.416 236.628 ; 
        RECT 6.88 232.254 6.984 236.628 ; 
        RECT 6.448 232.254 6.552 236.628 ; 
        RECT 6.016 232.254 6.12 236.628 ; 
        RECT 5.584 232.254 5.688 236.628 ; 
        RECT 5.152 232.254 5.256 236.628 ; 
        RECT 4.72 232.254 4.824 236.628 ; 
        RECT 4.288 232.254 4.392 236.628 ; 
        RECT 3.856 232.254 3.96 236.628 ; 
        RECT 3.424 232.254 3.528 236.628 ; 
        RECT 2.992 232.254 3.096 236.628 ; 
        RECT 2.56 232.254 2.664 236.628 ; 
        RECT 2.128 232.254 2.232 236.628 ; 
        RECT 1.696 232.254 1.8 236.628 ; 
        RECT 1.264 232.254 1.368 236.628 ; 
        RECT 0.832 232.254 0.936 236.628 ; 
        RECT 0.02 232.254 0.36 236.628 ; 
        RECT 34.564 236.574 35.076 240.948 ; 
        RECT 34.508 239.236 35.076 240.526 ; 
        RECT 33.916 238.144 34.164 240.948 ; 
        RECT 33.86 239.382 34.164 239.996 ; 
        RECT 33.916 236.574 34.02 240.948 ; 
        RECT 33.916 237.058 34.076 238.016 ; 
        RECT 33.916 236.574 34.164 236.93 ; 
        RECT 32.728 238.376 33.552 240.948 ; 
        RECT 33.448 236.574 33.552 240.948 ; 
        RECT 32.728 239.484 33.608 240.516 ; 
        RECT 32.728 236.574 33.12 240.948 ; 
        RECT 31.06 236.574 31.392 240.948 ; 
        RECT 31.06 236.928 31.448 240.67 ; 
        RECT 65.776 236.574 66.116 240.948 ; 
        RECT 65.2 236.574 65.304 240.948 ; 
        RECT 64.768 236.574 64.872 240.948 ; 
        RECT 64.336 236.574 64.44 240.948 ; 
        RECT 63.904 236.574 64.008 240.948 ; 
        RECT 63.472 236.574 63.576 240.948 ; 
        RECT 63.04 236.574 63.144 240.948 ; 
        RECT 62.608 236.574 62.712 240.948 ; 
        RECT 62.176 236.574 62.28 240.948 ; 
        RECT 61.744 236.574 61.848 240.948 ; 
        RECT 61.312 236.574 61.416 240.948 ; 
        RECT 60.88 236.574 60.984 240.948 ; 
        RECT 60.448 236.574 60.552 240.948 ; 
        RECT 60.016 236.574 60.12 240.948 ; 
        RECT 59.584 236.574 59.688 240.948 ; 
        RECT 59.152 236.574 59.256 240.948 ; 
        RECT 58.72 236.574 58.824 240.948 ; 
        RECT 58.288 236.574 58.392 240.948 ; 
        RECT 57.856 236.574 57.96 240.948 ; 
        RECT 57.424 236.574 57.528 240.948 ; 
        RECT 56.992 236.574 57.096 240.948 ; 
        RECT 56.56 236.574 56.664 240.948 ; 
        RECT 56.128 236.574 56.232 240.948 ; 
        RECT 55.696 236.574 55.8 240.948 ; 
        RECT 55.264 236.574 55.368 240.948 ; 
        RECT 54.832 236.574 54.936 240.948 ; 
        RECT 54.4 236.574 54.504 240.948 ; 
        RECT 53.968 236.574 54.072 240.948 ; 
        RECT 53.536 236.574 53.64 240.948 ; 
        RECT 53.104 236.574 53.208 240.948 ; 
        RECT 52.672 236.574 52.776 240.948 ; 
        RECT 52.24 236.574 52.344 240.948 ; 
        RECT 51.808 236.574 51.912 240.948 ; 
        RECT 51.376 236.574 51.48 240.948 ; 
        RECT 50.944 236.574 51.048 240.948 ; 
        RECT 50.512 236.574 50.616 240.948 ; 
        RECT 50.08 236.574 50.184 240.948 ; 
        RECT 49.648 236.574 49.752 240.948 ; 
        RECT 49.216 236.574 49.32 240.948 ; 
        RECT 48.784 236.574 48.888 240.948 ; 
        RECT 48.352 236.574 48.456 240.948 ; 
        RECT 47.92 236.574 48.024 240.948 ; 
        RECT 47.488 236.574 47.592 240.948 ; 
        RECT 47.056 236.574 47.16 240.948 ; 
        RECT 46.624 236.574 46.728 240.948 ; 
        RECT 46.192 236.574 46.296 240.948 ; 
        RECT 45.76 236.574 45.864 240.948 ; 
        RECT 45.328 236.574 45.432 240.948 ; 
        RECT 44.896 236.574 45 240.948 ; 
        RECT 44.464 236.574 44.568 240.948 ; 
        RECT 44.032 236.574 44.136 240.948 ; 
        RECT 43.6 236.574 43.704 240.948 ; 
        RECT 43.168 236.574 43.272 240.948 ; 
        RECT 42.736 236.574 42.84 240.948 ; 
        RECT 42.304 236.574 42.408 240.948 ; 
        RECT 41.872 236.574 41.976 240.948 ; 
        RECT 41.44 236.574 41.544 240.948 ; 
        RECT 41.008 236.574 41.112 240.948 ; 
        RECT 40.576 236.574 40.68 240.948 ; 
        RECT 40.144 236.574 40.248 240.948 ; 
        RECT 39.712 236.574 39.816 240.948 ; 
        RECT 39.28 236.574 39.384 240.948 ; 
        RECT 38.848 236.574 38.952 240.948 ; 
        RECT 38.416 236.574 38.52 240.948 ; 
        RECT 37.984 236.574 38.088 240.948 ; 
        RECT 37.552 236.574 37.656 240.948 ; 
        RECT 36.7 236.574 37.008 240.948 ; 
        RECT 29.128 236.574 29.436 240.948 ; 
        RECT 28.48 236.574 28.584 240.948 ; 
        RECT 28.048 236.574 28.152 240.948 ; 
        RECT 27.616 236.574 27.72 240.948 ; 
        RECT 27.184 236.574 27.288 240.948 ; 
        RECT 26.752 236.574 26.856 240.948 ; 
        RECT 26.32 236.574 26.424 240.948 ; 
        RECT 25.888 236.574 25.992 240.948 ; 
        RECT 25.456 236.574 25.56 240.948 ; 
        RECT 25.024 236.574 25.128 240.948 ; 
        RECT 24.592 236.574 24.696 240.948 ; 
        RECT 24.16 236.574 24.264 240.948 ; 
        RECT 23.728 236.574 23.832 240.948 ; 
        RECT 23.296 236.574 23.4 240.948 ; 
        RECT 22.864 236.574 22.968 240.948 ; 
        RECT 22.432 236.574 22.536 240.948 ; 
        RECT 22 236.574 22.104 240.948 ; 
        RECT 21.568 236.574 21.672 240.948 ; 
        RECT 21.136 236.574 21.24 240.948 ; 
        RECT 20.704 236.574 20.808 240.948 ; 
        RECT 20.272 236.574 20.376 240.948 ; 
        RECT 19.84 236.574 19.944 240.948 ; 
        RECT 19.408 236.574 19.512 240.948 ; 
        RECT 18.976 236.574 19.08 240.948 ; 
        RECT 18.544 236.574 18.648 240.948 ; 
        RECT 18.112 236.574 18.216 240.948 ; 
        RECT 17.68 236.574 17.784 240.948 ; 
        RECT 17.248 236.574 17.352 240.948 ; 
        RECT 16.816 236.574 16.92 240.948 ; 
        RECT 16.384 236.574 16.488 240.948 ; 
        RECT 15.952 236.574 16.056 240.948 ; 
        RECT 15.52 236.574 15.624 240.948 ; 
        RECT 15.088 236.574 15.192 240.948 ; 
        RECT 14.656 236.574 14.76 240.948 ; 
        RECT 14.224 236.574 14.328 240.948 ; 
        RECT 13.792 236.574 13.896 240.948 ; 
        RECT 13.36 236.574 13.464 240.948 ; 
        RECT 12.928 236.574 13.032 240.948 ; 
        RECT 12.496 236.574 12.6 240.948 ; 
        RECT 12.064 236.574 12.168 240.948 ; 
        RECT 11.632 236.574 11.736 240.948 ; 
        RECT 11.2 236.574 11.304 240.948 ; 
        RECT 10.768 236.574 10.872 240.948 ; 
        RECT 10.336 236.574 10.44 240.948 ; 
        RECT 9.904 236.574 10.008 240.948 ; 
        RECT 9.472 236.574 9.576 240.948 ; 
        RECT 9.04 236.574 9.144 240.948 ; 
        RECT 8.608 236.574 8.712 240.948 ; 
        RECT 8.176 236.574 8.28 240.948 ; 
        RECT 7.744 236.574 7.848 240.948 ; 
        RECT 7.312 236.574 7.416 240.948 ; 
        RECT 6.88 236.574 6.984 240.948 ; 
        RECT 6.448 236.574 6.552 240.948 ; 
        RECT 6.016 236.574 6.12 240.948 ; 
        RECT 5.584 236.574 5.688 240.948 ; 
        RECT 5.152 236.574 5.256 240.948 ; 
        RECT 4.72 236.574 4.824 240.948 ; 
        RECT 4.288 236.574 4.392 240.948 ; 
        RECT 3.856 236.574 3.96 240.948 ; 
        RECT 3.424 236.574 3.528 240.948 ; 
        RECT 2.992 236.574 3.096 240.948 ; 
        RECT 2.56 236.574 2.664 240.948 ; 
        RECT 2.128 236.574 2.232 240.948 ; 
        RECT 1.696 236.574 1.8 240.948 ; 
        RECT 1.264 236.574 1.368 240.948 ; 
        RECT 0.832 236.574 0.936 240.948 ; 
        RECT 0.02 236.574 0.36 240.948 ; 
  LAYER V3 SPACING 0.072 ; 
      RECT 0.02 4.88 66.116 5.4 ; 
      RECT 65.648 1.026 66.116 5.4 ; 
      RECT 37.208 4.496 65.576 5.4 ; 
      RECT 31.88 4.496 37.136 5.4 ; 
      RECT 29 1.026 31.52 5.4 ; 
      RECT 0.56 4.496 28.928 5.4 ; 
      RECT 0.02 1.026 0.488 5.4 ; 
      RECT 65.504 1.026 66.116 4.688 ; 
      RECT 37.424 1.026 65.432 5.4 ; 
      RECT 34.436 1.026 37.352 4.688 ; 
      RECT 33.788 1.808 34.292 5.4 ; 
      RECT 28.784 1.424 33.68 4.688 ; 
      RECT 0.704 1.026 28.712 5.4 ; 
      RECT 0.02 1.026 0.632 4.688 ; 
      RECT 34.22 1.026 66.116 4.304 ; 
      RECT 0.02 1.424 34.148 4.304 ; 
      RECT 33.32 1.026 66.116 1.712 ; 
      RECT 0.02 1.026 33.248 4.304 ; 
      RECT 0.02 1.026 66.116 1.328 ; 
      RECT 0.02 9.2 66.116 9.72 ; 
      RECT 65.648 5.346 66.116 9.72 ; 
      RECT 37.208 8.816 65.576 9.72 ; 
      RECT 31.88 8.816 37.136 9.72 ; 
      RECT 29 5.346 31.52 9.72 ; 
      RECT 0.56 8.816 28.928 9.72 ; 
      RECT 0.02 5.346 0.488 9.72 ; 
      RECT 65.504 5.346 66.116 9.008 ; 
      RECT 37.424 5.346 65.432 9.72 ; 
      RECT 34.436 5.346 37.352 9.008 ; 
      RECT 33.788 6.128 34.292 9.72 ; 
      RECT 28.784 5.744 33.68 9.008 ; 
      RECT 0.704 5.346 28.712 9.72 ; 
      RECT 0.02 5.346 0.632 9.008 ; 
      RECT 34.22 5.346 66.116 8.624 ; 
      RECT 0.02 5.744 34.148 8.624 ; 
      RECT 33.32 5.346 66.116 6.032 ; 
      RECT 0.02 5.346 33.248 8.624 ; 
      RECT 0.02 5.346 66.116 5.648 ; 
      RECT 0.02 13.52 66.116 14.04 ; 
      RECT 65.648 9.666 66.116 14.04 ; 
      RECT 37.208 13.136 65.576 14.04 ; 
      RECT 31.88 13.136 37.136 14.04 ; 
      RECT 29 9.666 31.52 14.04 ; 
      RECT 0.56 13.136 28.928 14.04 ; 
      RECT 0.02 9.666 0.488 14.04 ; 
      RECT 65.504 9.666 66.116 13.328 ; 
      RECT 37.424 9.666 65.432 14.04 ; 
      RECT 34.436 9.666 37.352 13.328 ; 
      RECT 33.788 10.448 34.292 14.04 ; 
      RECT 28.784 10.064 33.68 13.328 ; 
      RECT 0.704 9.666 28.712 14.04 ; 
      RECT 0.02 9.666 0.632 13.328 ; 
      RECT 34.22 9.666 66.116 12.944 ; 
      RECT 0.02 10.064 34.148 12.944 ; 
      RECT 33.32 9.666 66.116 10.352 ; 
      RECT 0.02 9.666 33.248 12.944 ; 
      RECT 0.02 9.666 66.116 9.968 ; 
      RECT 0.02 17.84 66.116 18.36 ; 
      RECT 65.648 13.986 66.116 18.36 ; 
      RECT 37.208 17.456 65.576 18.36 ; 
      RECT 31.88 17.456 37.136 18.36 ; 
      RECT 29 13.986 31.52 18.36 ; 
      RECT 0.56 17.456 28.928 18.36 ; 
      RECT 0.02 13.986 0.488 18.36 ; 
      RECT 65.504 13.986 66.116 17.648 ; 
      RECT 37.424 13.986 65.432 18.36 ; 
      RECT 34.436 13.986 37.352 17.648 ; 
      RECT 33.788 14.768 34.292 18.36 ; 
      RECT 28.784 14.384 33.68 17.648 ; 
      RECT 0.704 13.986 28.712 18.36 ; 
      RECT 0.02 13.986 0.632 17.648 ; 
      RECT 34.22 13.986 66.116 17.264 ; 
      RECT 0.02 14.384 34.148 17.264 ; 
      RECT 33.32 13.986 66.116 14.672 ; 
      RECT 0.02 13.986 33.248 17.264 ; 
      RECT 0.02 13.986 66.116 14.288 ; 
      RECT 0.02 22.16 66.116 22.68 ; 
      RECT 65.648 18.306 66.116 22.68 ; 
      RECT 37.208 21.776 65.576 22.68 ; 
      RECT 31.88 21.776 37.136 22.68 ; 
      RECT 29 18.306 31.52 22.68 ; 
      RECT 0.56 21.776 28.928 22.68 ; 
      RECT 0.02 18.306 0.488 22.68 ; 
      RECT 65.504 18.306 66.116 21.968 ; 
      RECT 37.424 18.306 65.432 22.68 ; 
      RECT 34.436 18.306 37.352 21.968 ; 
      RECT 33.788 19.088 34.292 22.68 ; 
      RECT 28.784 18.704 33.68 21.968 ; 
      RECT 0.704 18.306 28.712 22.68 ; 
      RECT 0.02 18.306 0.632 21.968 ; 
      RECT 34.22 18.306 66.116 21.584 ; 
      RECT 0.02 18.704 34.148 21.584 ; 
      RECT 33.32 18.306 66.116 18.992 ; 
      RECT 0.02 18.306 33.248 21.584 ; 
      RECT 0.02 18.306 66.116 18.608 ; 
      RECT 0.02 26.48 66.116 27 ; 
      RECT 65.648 22.626 66.116 27 ; 
      RECT 37.208 26.096 65.576 27 ; 
      RECT 31.88 26.096 37.136 27 ; 
      RECT 29 22.626 31.52 27 ; 
      RECT 0.56 26.096 28.928 27 ; 
      RECT 0.02 22.626 0.488 27 ; 
      RECT 65.504 22.626 66.116 26.288 ; 
      RECT 37.424 22.626 65.432 27 ; 
      RECT 34.436 22.626 37.352 26.288 ; 
      RECT 33.788 23.408 34.292 27 ; 
      RECT 28.784 23.024 33.68 26.288 ; 
      RECT 0.704 22.626 28.712 27 ; 
      RECT 0.02 22.626 0.632 26.288 ; 
      RECT 34.22 22.626 66.116 25.904 ; 
      RECT 0.02 23.024 34.148 25.904 ; 
      RECT 33.32 22.626 66.116 23.312 ; 
      RECT 0.02 22.626 33.248 25.904 ; 
      RECT 0.02 22.626 66.116 22.928 ; 
      RECT 0.02 30.8 66.116 31.32 ; 
      RECT 65.648 26.946 66.116 31.32 ; 
      RECT 37.208 30.416 65.576 31.32 ; 
      RECT 31.88 30.416 37.136 31.32 ; 
      RECT 29 26.946 31.52 31.32 ; 
      RECT 0.56 30.416 28.928 31.32 ; 
      RECT 0.02 26.946 0.488 31.32 ; 
      RECT 65.504 26.946 66.116 30.608 ; 
      RECT 37.424 26.946 65.432 31.32 ; 
      RECT 34.436 26.946 37.352 30.608 ; 
      RECT 33.788 27.728 34.292 31.32 ; 
      RECT 28.784 27.344 33.68 30.608 ; 
      RECT 0.704 26.946 28.712 31.32 ; 
      RECT 0.02 26.946 0.632 30.608 ; 
      RECT 34.22 26.946 66.116 30.224 ; 
      RECT 0.02 27.344 34.148 30.224 ; 
      RECT 33.32 26.946 66.116 27.632 ; 
      RECT 0.02 26.946 33.248 30.224 ; 
      RECT 0.02 26.946 66.116 27.248 ; 
      RECT 0.02 35.12 66.116 35.64 ; 
      RECT 65.648 31.266 66.116 35.64 ; 
      RECT 37.208 34.736 65.576 35.64 ; 
      RECT 31.88 34.736 37.136 35.64 ; 
      RECT 29 31.266 31.52 35.64 ; 
      RECT 0.56 34.736 28.928 35.64 ; 
      RECT 0.02 31.266 0.488 35.64 ; 
      RECT 65.504 31.266 66.116 34.928 ; 
      RECT 37.424 31.266 65.432 35.64 ; 
      RECT 34.436 31.266 37.352 34.928 ; 
      RECT 33.788 32.048 34.292 35.64 ; 
      RECT 28.784 31.664 33.68 34.928 ; 
      RECT 0.704 31.266 28.712 35.64 ; 
      RECT 0.02 31.266 0.632 34.928 ; 
      RECT 34.22 31.266 66.116 34.544 ; 
      RECT 0.02 31.664 34.148 34.544 ; 
      RECT 33.32 31.266 66.116 31.952 ; 
      RECT 0.02 31.266 33.248 34.544 ; 
      RECT 0.02 31.266 66.116 31.568 ; 
      RECT 0.02 39.44 66.116 39.96 ; 
      RECT 65.648 35.586 66.116 39.96 ; 
      RECT 37.208 39.056 65.576 39.96 ; 
      RECT 31.88 39.056 37.136 39.96 ; 
      RECT 29 35.586 31.52 39.96 ; 
      RECT 0.56 39.056 28.928 39.96 ; 
      RECT 0.02 35.586 0.488 39.96 ; 
      RECT 65.504 35.586 66.116 39.248 ; 
      RECT 37.424 35.586 65.432 39.96 ; 
      RECT 34.436 35.586 37.352 39.248 ; 
      RECT 33.788 36.368 34.292 39.96 ; 
      RECT 28.784 35.984 33.68 39.248 ; 
      RECT 0.704 35.586 28.712 39.96 ; 
      RECT 0.02 35.586 0.632 39.248 ; 
      RECT 34.22 35.586 66.116 38.864 ; 
      RECT 0.02 35.984 34.148 38.864 ; 
      RECT 33.32 35.586 66.116 36.272 ; 
      RECT 0.02 35.586 33.248 38.864 ; 
      RECT 0.02 35.586 66.116 35.888 ; 
      RECT 0.02 43.76 66.116 44.28 ; 
      RECT 65.648 39.906 66.116 44.28 ; 
      RECT 37.208 43.376 65.576 44.28 ; 
      RECT 31.88 43.376 37.136 44.28 ; 
      RECT 29 39.906 31.52 44.28 ; 
      RECT 0.56 43.376 28.928 44.28 ; 
      RECT 0.02 39.906 0.488 44.28 ; 
      RECT 65.504 39.906 66.116 43.568 ; 
      RECT 37.424 39.906 65.432 44.28 ; 
      RECT 34.436 39.906 37.352 43.568 ; 
      RECT 33.788 40.688 34.292 44.28 ; 
      RECT 28.784 40.304 33.68 43.568 ; 
      RECT 0.704 39.906 28.712 44.28 ; 
      RECT 0.02 39.906 0.632 43.568 ; 
      RECT 34.22 39.906 66.116 43.184 ; 
      RECT 0.02 40.304 34.148 43.184 ; 
      RECT 33.32 39.906 66.116 40.592 ; 
      RECT 0.02 39.906 33.248 43.184 ; 
      RECT 0.02 39.906 66.116 40.208 ; 
      RECT 0.02 48.08 66.116 48.6 ; 
      RECT 65.648 44.226 66.116 48.6 ; 
      RECT 37.208 47.696 65.576 48.6 ; 
      RECT 31.88 47.696 37.136 48.6 ; 
      RECT 29 44.226 31.52 48.6 ; 
      RECT 0.56 47.696 28.928 48.6 ; 
      RECT 0.02 44.226 0.488 48.6 ; 
      RECT 65.504 44.226 66.116 47.888 ; 
      RECT 37.424 44.226 65.432 48.6 ; 
      RECT 34.436 44.226 37.352 47.888 ; 
      RECT 33.788 45.008 34.292 48.6 ; 
      RECT 28.784 44.624 33.68 47.888 ; 
      RECT 0.704 44.226 28.712 48.6 ; 
      RECT 0.02 44.226 0.632 47.888 ; 
      RECT 34.22 44.226 66.116 47.504 ; 
      RECT 0.02 44.624 34.148 47.504 ; 
      RECT 33.32 44.226 66.116 44.912 ; 
      RECT 0.02 44.226 33.248 47.504 ; 
      RECT 0.02 44.226 66.116 44.528 ; 
      RECT 0.02 52.4 66.116 52.92 ; 
      RECT 65.648 48.546 66.116 52.92 ; 
      RECT 37.208 52.016 65.576 52.92 ; 
      RECT 31.88 52.016 37.136 52.92 ; 
      RECT 29 48.546 31.52 52.92 ; 
      RECT 0.56 52.016 28.928 52.92 ; 
      RECT 0.02 48.546 0.488 52.92 ; 
      RECT 65.504 48.546 66.116 52.208 ; 
      RECT 37.424 48.546 65.432 52.92 ; 
      RECT 34.436 48.546 37.352 52.208 ; 
      RECT 33.788 49.328 34.292 52.92 ; 
      RECT 28.784 48.944 33.68 52.208 ; 
      RECT 0.704 48.546 28.712 52.92 ; 
      RECT 0.02 48.546 0.632 52.208 ; 
      RECT 34.22 48.546 66.116 51.824 ; 
      RECT 0.02 48.944 34.148 51.824 ; 
      RECT 33.32 48.546 66.116 49.232 ; 
      RECT 0.02 48.546 33.248 51.824 ; 
      RECT 0.02 48.546 66.116 48.848 ; 
      RECT 0.02 56.72 66.116 57.24 ; 
      RECT 65.648 52.866 66.116 57.24 ; 
      RECT 37.208 56.336 65.576 57.24 ; 
      RECT 31.88 56.336 37.136 57.24 ; 
      RECT 29 52.866 31.52 57.24 ; 
      RECT 0.56 56.336 28.928 57.24 ; 
      RECT 0.02 52.866 0.488 57.24 ; 
      RECT 65.504 52.866 66.116 56.528 ; 
      RECT 37.424 52.866 65.432 57.24 ; 
      RECT 34.436 52.866 37.352 56.528 ; 
      RECT 33.788 53.648 34.292 57.24 ; 
      RECT 28.784 53.264 33.68 56.528 ; 
      RECT 0.704 52.866 28.712 57.24 ; 
      RECT 0.02 52.866 0.632 56.528 ; 
      RECT 34.22 52.866 66.116 56.144 ; 
      RECT 0.02 53.264 34.148 56.144 ; 
      RECT 33.32 52.866 66.116 53.552 ; 
      RECT 0.02 52.866 33.248 56.144 ; 
      RECT 0.02 52.866 66.116 53.168 ; 
      RECT 0.02 61.04 66.116 61.56 ; 
      RECT 65.648 57.186 66.116 61.56 ; 
      RECT 37.208 60.656 65.576 61.56 ; 
      RECT 31.88 60.656 37.136 61.56 ; 
      RECT 29 57.186 31.52 61.56 ; 
      RECT 0.56 60.656 28.928 61.56 ; 
      RECT 0.02 57.186 0.488 61.56 ; 
      RECT 65.504 57.186 66.116 60.848 ; 
      RECT 37.424 57.186 65.432 61.56 ; 
      RECT 34.436 57.186 37.352 60.848 ; 
      RECT 33.788 57.968 34.292 61.56 ; 
      RECT 28.784 57.584 33.68 60.848 ; 
      RECT 0.704 57.186 28.712 61.56 ; 
      RECT 0.02 57.186 0.632 60.848 ; 
      RECT 34.22 57.186 66.116 60.464 ; 
      RECT 0.02 57.584 34.148 60.464 ; 
      RECT 33.32 57.186 66.116 57.872 ; 
      RECT 0.02 57.186 33.248 60.464 ; 
      RECT 0.02 57.186 66.116 57.488 ; 
      RECT 0.02 65.36 66.116 65.88 ; 
      RECT 65.648 61.506 66.116 65.88 ; 
      RECT 37.208 64.976 65.576 65.88 ; 
      RECT 31.88 64.976 37.136 65.88 ; 
      RECT 29 61.506 31.52 65.88 ; 
      RECT 0.56 64.976 28.928 65.88 ; 
      RECT 0.02 61.506 0.488 65.88 ; 
      RECT 65.504 61.506 66.116 65.168 ; 
      RECT 37.424 61.506 65.432 65.88 ; 
      RECT 34.436 61.506 37.352 65.168 ; 
      RECT 33.788 62.288 34.292 65.88 ; 
      RECT 28.784 61.904 33.68 65.168 ; 
      RECT 0.704 61.506 28.712 65.88 ; 
      RECT 0.02 61.506 0.632 65.168 ; 
      RECT 34.22 61.506 66.116 64.784 ; 
      RECT 0.02 61.904 34.148 64.784 ; 
      RECT 33.32 61.506 66.116 62.192 ; 
      RECT 0.02 61.506 33.248 64.784 ; 
      RECT 0.02 61.506 66.116 61.808 ; 
      RECT 0.02 69.68 66.116 70.2 ; 
      RECT 65.648 65.826 66.116 70.2 ; 
      RECT 37.208 69.296 65.576 70.2 ; 
      RECT 31.88 69.296 37.136 70.2 ; 
      RECT 29 65.826 31.52 70.2 ; 
      RECT 0.56 69.296 28.928 70.2 ; 
      RECT 0.02 65.826 0.488 70.2 ; 
      RECT 65.504 65.826 66.116 69.488 ; 
      RECT 37.424 65.826 65.432 70.2 ; 
      RECT 34.436 65.826 37.352 69.488 ; 
      RECT 33.788 66.608 34.292 70.2 ; 
      RECT 28.784 66.224 33.68 69.488 ; 
      RECT 0.704 65.826 28.712 70.2 ; 
      RECT 0.02 65.826 0.632 69.488 ; 
      RECT 34.22 65.826 66.116 69.104 ; 
      RECT 0.02 66.224 34.148 69.104 ; 
      RECT 33.32 65.826 66.116 66.512 ; 
      RECT 0.02 65.826 33.248 69.104 ; 
      RECT 0.02 65.826 66.116 66.128 ; 
      RECT 0.02 74 66.116 74.52 ; 
      RECT 65.648 70.146 66.116 74.52 ; 
      RECT 37.208 73.616 65.576 74.52 ; 
      RECT 31.88 73.616 37.136 74.52 ; 
      RECT 29 70.146 31.52 74.52 ; 
      RECT 0.56 73.616 28.928 74.52 ; 
      RECT 0.02 70.146 0.488 74.52 ; 
      RECT 65.504 70.146 66.116 73.808 ; 
      RECT 37.424 70.146 65.432 74.52 ; 
      RECT 34.436 70.146 37.352 73.808 ; 
      RECT 33.788 70.928 34.292 74.52 ; 
      RECT 28.784 70.544 33.68 73.808 ; 
      RECT 0.704 70.146 28.712 74.52 ; 
      RECT 0.02 70.146 0.632 73.808 ; 
      RECT 34.22 70.146 66.116 73.424 ; 
      RECT 0.02 70.544 34.148 73.424 ; 
      RECT 33.32 70.146 66.116 70.832 ; 
      RECT 0.02 70.146 33.248 73.424 ; 
      RECT 0.02 70.146 66.116 70.448 ; 
      RECT 0.02 78.32 66.116 78.84 ; 
      RECT 65.648 74.466 66.116 78.84 ; 
      RECT 37.208 77.936 65.576 78.84 ; 
      RECT 31.88 77.936 37.136 78.84 ; 
      RECT 29 74.466 31.52 78.84 ; 
      RECT 0.56 77.936 28.928 78.84 ; 
      RECT 0.02 74.466 0.488 78.84 ; 
      RECT 65.504 74.466 66.116 78.128 ; 
      RECT 37.424 74.466 65.432 78.84 ; 
      RECT 34.436 74.466 37.352 78.128 ; 
      RECT 33.788 75.248 34.292 78.84 ; 
      RECT 28.784 74.864 33.68 78.128 ; 
      RECT 0.704 74.466 28.712 78.84 ; 
      RECT 0.02 74.466 0.632 78.128 ; 
      RECT 34.22 74.466 66.116 77.744 ; 
      RECT 0.02 74.864 34.148 77.744 ; 
      RECT 33.32 74.466 66.116 75.152 ; 
      RECT 0.02 74.466 33.248 77.744 ; 
      RECT 0.02 74.466 66.116 74.768 ; 
      RECT 0.02 82.64 66.116 83.16 ; 
      RECT 65.648 78.786 66.116 83.16 ; 
      RECT 37.208 82.256 65.576 83.16 ; 
      RECT 31.88 82.256 37.136 83.16 ; 
      RECT 29 78.786 31.52 83.16 ; 
      RECT 0.56 82.256 28.928 83.16 ; 
      RECT 0.02 78.786 0.488 83.16 ; 
      RECT 65.504 78.786 66.116 82.448 ; 
      RECT 37.424 78.786 65.432 83.16 ; 
      RECT 34.436 78.786 37.352 82.448 ; 
      RECT 33.788 79.568 34.292 83.16 ; 
      RECT 28.784 79.184 33.68 82.448 ; 
      RECT 0.704 78.786 28.712 83.16 ; 
      RECT 0.02 78.786 0.632 82.448 ; 
      RECT 34.22 78.786 66.116 82.064 ; 
      RECT 0.02 79.184 34.148 82.064 ; 
      RECT 33.32 78.786 66.116 79.472 ; 
      RECT 0.02 78.786 33.248 82.064 ; 
      RECT 0.02 78.786 66.116 79.088 ; 
      RECT 0.02 86.96 66.116 87.48 ; 
      RECT 65.648 83.106 66.116 87.48 ; 
      RECT 37.208 86.576 65.576 87.48 ; 
      RECT 31.88 86.576 37.136 87.48 ; 
      RECT 29 83.106 31.52 87.48 ; 
      RECT 0.56 86.576 28.928 87.48 ; 
      RECT 0.02 83.106 0.488 87.48 ; 
      RECT 65.504 83.106 66.116 86.768 ; 
      RECT 37.424 83.106 65.432 87.48 ; 
      RECT 34.436 83.106 37.352 86.768 ; 
      RECT 33.788 83.888 34.292 87.48 ; 
      RECT 28.784 83.504 33.68 86.768 ; 
      RECT 0.704 83.106 28.712 87.48 ; 
      RECT 0.02 83.106 0.632 86.768 ; 
      RECT 34.22 83.106 66.116 86.384 ; 
      RECT 0.02 83.504 34.148 86.384 ; 
      RECT 33.32 83.106 66.116 83.792 ; 
      RECT 0.02 83.106 33.248 86.384 ; 
      RECT 0.02 83.106 66.116 83.408 ; 
      RECT 0.02 91.28 66.116 91.8 ; 
      RECT 65.648 87.426 66.116 91.8 ; 
      RECT 37.208 90.896 65.576 91.8 ; 
      RECT 31.88 90.896 37.136 91.8 ; 
      RECT 29 87.426 31.52 91.8 ; 
      RECT 0.56 90.896 28.928 91.8 ; 
      RECT 0.02 87.426 0.488 91.8 ; 
      RECT 65.504 87.426 66.116 91.088 ; 
      RECT 37.424 87.426 65.432 91.8 ; 
      RECT 34.436 87.426 37.352 91.088 ; 
      RECT 33.788 88.208 34.292 91.8 ; 
      RECT 28.784 87.824 33.68 91.088 ; 
      RECT 0.704 87.426 28.712 91.8 ; 
      RECT 0.02 87.426 0.632 91.088 ; 
      RECT 34.22 87.426 66.116 90.704 ; 
      RECT 0.02 87.824 34.148 90.704 ; 
      RECT 33.32 87.426 66.116 88.112 ; 
      RECT 0.02 87.426 33.248 90.704 ; 
      RECT 0.02 87.426 66.116 87.728 ; 
      RECT 0.02 95.6 66.116 96.12 ; 
      RECT 65.648 91.746 66.116 96.12 ; 
      RECT 37.208 95.216 65.576 96.12 ; 
      RECT 31.88 95.216 37.136 96.12 ; 
      RECT 29 91.746 31.52 96.12 ; 
      RECT 0.56 95.216 28.928 96.12 ; 
      RECT 0.02 91.746 0.488 96.12 ; 
      RECT 65.504 91.746 66.116 95.408 ; 
      RECT 37.424 91.746 65.432 96.12 ; 
      RECT 34.436 91.746 37.352 95.408 ; 
      RECT 33.788 92.528 34.292 96.12 ; 
      RECT 28.784 92.144 33.68 95.408 ; 
      RECT 0.704 91.746 28.712 96.12 ; 
      RECT 0.02 91.746 0.632 95.408 ; 
      RECT 34.22 91.746 66.116 95.024 ; 
      RECT 0.02 92.144 34.148 95.024 ; 
      RECT 33.32 91.746 66.116 92.432 ; 
      RECT 0.02 91.746 33.248 95.024 ; 
      RECT 0.02 91.746 66.116 92.048 ; 
      RECT 0.02 99.92 66.116 100.44 ; 
      RECT 65.648 96.066 66.116 100.44 ; 
      RECT 37.208 99.536 65.576 100.44 ; 
      RECT 31.88 99.536 37.136 100.44 ; 
      RECT 29 96.066 31.52 100.44 ; 
      RECT 0.56 99.536 28.928 100.44 ; 
      RECT 0.02 96.066 0.488 100.44 ; 
      RECT 65.504 96.066 66.116 99.728 ; 
      RECT 37.424 96.066 65.432 100.44 ; 
      RECT 34.436 96.066 37.352 99.728 ; 
      RECT 33.788 96.848 34.292 100.44 ; 
      RECT 28.784 96.464 33.68 99.728 ; 
      RECT 0.704 96.066 28.712 100.44 ; 
      RECT 0.02 96.066 0.632 99.728 ; 
      RECT 34.22 96.066 66.116 99.344 ; 
      RECT 0.02 96.464 34.148 99.344 ; 
      RECT 33.32 96.066 66.116 96.752 ; 
      RECT 0.02 96.066 33.248 99.344 ; 
      RECT 0.02 96.066 66.116 96.368 ; 
      RECT 0.02 104.24 66.116 104.76 ; 
      RECT 65.648 100.386 66.116 104.76 ; 
      RECT 37.208 103.856 65.576 104.76 ; 
      RECT 31.88 103.856 37.136 104.76 ; 
      RECT 29 100.386 31.52 104.76 ; 
      RECT 0.56 103.856 28.928 104.76 ; 
      RECT 0.02 100.386 0.488 104.76 ; 
      RECT 65.504 100.386 66.116 104.048 ; 
      RECT 37.424 100.386 65.432 104.76 ; 
      RECT 34.436 100.386 37.352 104.048 ; 
      RECT 33.788 101.168 34.292 104.76 ; 
      RECT 28.784 100.784 33.68 104.048 ; 
      RECT 0.704 100.386 28.712 104.76 ; 
      RECT 0.02 100.386 0.632 104.048 ; 
      RECT 34.22 100.386 66.116 103.664 ; 
      RECT 0.02 100.784 34.148 103.664 ; 
      RECT 33.32 100.386 66.116 101.072 ; 
      RECT 0.02 100.386 33.248 103.664 ; 
      RECT 0.02 100.386 66.116 100.688 ; 
      RECT 0 133.908 66.096 139.242 ; 
      RECT 43.236 104.628 66.096 139.242 ; 
      RECT 34.436 120.084 66.096 139.242 ; 
      RECT 38.052 109.716 66.096 139.242 ; 
      RECT 34.228 104.628 34.364 139.242 ; 
      RECT 34.02 104.628 34.156 139.242 ; 
      RECT 33.812 104.628 33.948 139.242 ; 
      RECT 33.604 104.628 33.74 139.242 ; 
      RECT 0 132.18 33.532 139.242 ; 
      RECT 32.564 121.236 66.096 133.044 ; 
      RECT 32.356 104.628 32.492 139.242 ; 
      RECT 32.148 104.628 32.284 139.242 ; 
      RECT 31.94 104.628 32.076 139.242 ; 
      RECT 31.732 104.628 31.868 139.242 ; 
      RECT 0 110.868 31.66 139.242 ; 
      RECT 0 119.508 33.532 131.316 ; 
      RECT 32.564 108.564 37.116 120.372 ; 
      RECT 37.26 110.484 66.096 139.242 ; 
      RECT 0 119.508 37.188 120.372 ; 
      RECT 32.564 110.484 66.096 119.988 ; 
      RECT 29.844 106.836 32.94 118.644 ; 
      RECT 28.98 107.412 31.66 139.242 ; 
      RECT 0 109.716 28.908 139.242 ; 
      RECT 27.252 104.628 29.052 110.772 ; 
      RECT 0 110.1 37.98 110.772 ; 
      RECT 37.188 109.716 66.096 110.388 ; 
      RECT 42.372 104.628 43.164 139.242 ; 
      RECT 27.252 108.948 42.3 110.004 ; 
      RECT 23.796 107.412 27.18 139.242 ; 
      RECT 0 104.628 23.724 139.242 ; 
      RECT 41.508 104.628 66.096 109.62 ; 
      RECT 40.644 107.412 66.096 109.62 ; 
      RECT 0 108.566 40.572 109.62 ; 
      RECT 39.78 104.628 41.436 108.852 ; 
      RECT 37.404 107.412 66.096 108.852 ; 
      RECT 34.436 107.412 37.332 110.004 ; 
      RECT 32.564 107.22 33.532 139.242 ; 
      RECT 33.012 104.628 34.524 107.7 ; 
      RECT 34.596 107.22 39.708 107.702 ; 
      RECT 26.388 107.22 29.772 109.62 ; 
      RECT 24.66 107.22 26.316 139.242 ; 
      RECT 0 104.628 24.588 109.62 ; 
      RECT 38.916 104.628 66.096 107.316 ; 
      RECT 33.012 104.948 38.844 107.316 ; 
      RECT 29.124 106.836 32.94 107.316 ; 
      RECT 25.524 104.628 29.052 107.316 ; 
      RECT 0 104.628 25.452 107.316 ; 
      RECT 37.188 104.628 66.096 107.124 ; 
      RECT 32.564 104.948 66.096 107.124 ; 
      RECT 0 104.628 31.66 107.124 ; 
      RECT 0 104.628 37.116 105.972 ; 
      RECT 0 104.628 66.096 104.852 ; 
        RECT 0.02 141.068 66.116 141.588 ; 
        RECT 65.648 137.214 66.116 141.588 ; 
        RECT 37.208 140.684 65.576 141.588 ; 
        RECT 31.88 140.684 37.136 141.588 ; 
        RECT 29 137.214 31.52 141.588 ; 
        RECT 0.56 140.684 28.928 141.588 ; 
        RECT 0.02 137.214 0.488 141.588 ; 
        RECT 65.504 137.214 66.116 140.876 ; 
        RECT 37.424 137.214 65.432 141.588 ; 
        RECT 34.436 137.214 37.352 140.876 ; 
        RECT 33.788 137.996 34.292 141.588 ; 
        RECT 28.784 137.612 33.68 140.876 ; 
        RECT 0.704 137.214 28.712 141.588 ; 
        RECT 0.02 137.214 0.632 140.876 ; 
        RECT 34.22 137.214 66.116 140.492 ; 
        RECT 0.02 137.612 34.148 140.492 ; 
        RECT 33.32 137.214 66.116 137.9 ; 
        RECT 0.02 137.214 33.248 140.492 ; 
        RECT 0.02 137.214 66.116 137.516 ; 
        RECT 0.02 145.388 66.116 145.908 ; 
        RECT 65.648 141.534 66.116 145.908 ; 
        RECT 37.208 145.004 65.576 145.908 ; 
        RECT 31.88 145.004 37.136 145.908 ; 
        RECT 29 141.534 31.52 145.908 ; 
        RECT 0.56 145.004 28.928 145.908 ; 
        RECT 0.02 141.534 0.488 145.908 ; 
        RECT 65.504 141.534 66.116 145.196 ; 
        RECT 37.424 141.534 65.432 145.908 ; 
        RECT 34.436 141.534 37.352 145.196 ; 
        RECT 33.788 142.316 34.292 145.908 ; 
        RECT 28.784 141.932 33.68 145.196 ; 
        RECT 0.704 141.534 28.712 145.908 ; 
        RECT 0.02 141.534 0.632 145.196 ; 
        RECT 34.22 141.534 66.116 144.812 ; 
        RECT 0.02 141.932 34.148 144.812 ; 
        RECT 33.32 141.534 66.116 142.22 ; 
        RECT 0.02 141.534 33.248 144.812 ; 
        RECT 0.02 141.534 66.116 141.836 ; 
        RECT 0.02 149.708 66.116 150.228 ; 
        RECT 65.648 145.854 66.116 150.228 ; 
        RECT 37.208 149.324 65.576 150.228 ; 
        RECT 31.88 149.324 37.136 150.228 ; 
        RECT 29 145.854 31.52 150.228 ; 
        RECT 0.56 149.324 28.928 150.228 ; 
        RECT 0.02 145.854 0.488 150.228 ; 
        RECT 65.504 145.854 66.116 149.516 ; 
        RECT 37.424 145.854 65.432 150.228 ; 
        RECT 34.436 145.854 37.352 149.516 ; 
        RECT 33.788 146.636 34.292 150.228 ; 
        RECT 28.784 146.252 33.68 149.516 ; 
        RECT 0.704 145.854 28.712 150.228 ; 
        RECT 0.02 145.854 0.632 149.516 ; 
        RECT 34.22 145.854 66.116 149.132 ; 
        RECT 0.02 146.252 34.148 149.132 ; 
        RECT 33.32 145.854 66.116 146.54 ; 
        RECT 0.02 145.854 33.248 149.132 ; 
        RECT 0.02 145.854 66.116 146.156 ; 
        RECT 0.02 154.028 66.116 154.548 ; 
        RECT 65.648 150.174 66.116 154.548 ; 
        RECT 37.208 153.644 65.576 154.548 ; 
        RECT 31.88 153.644 37.136 154.548 ; 
        RECT 29 150.174 31.52 154.548 ; 
        RECT 0.56 153.644 28.928 154.548 ; 
        RECT 0.02 150.174 0.488 154.548 ; 
        RECT 65.504 150.174 66.116 153.836 ; 
        RECT 37.424 150.174 65.432 154.548 ; 
        RECT 34.436 150.174 37.352 153.836 ; 
        RECT 33.788 150.956 34.292 154.548 ; 
        RECT 28.784 150.572 33.68 153.836 ; 
        RECT 0.704 150.174 28.712 154.548 ; 
        RECT 0.02 150.174 0.632 153.836 ; 
        RECT 34.22 150.174 66.116 153.452 ; 
        RECT 0.02 150.572 34.148 153.452 ; 
        RECT 33.32 150.174 66.116 150.86 ; 
        RECT 0.02 150.174 33.248 153.452 ; 
        RECT 0.02 150.174 66.116 150.476 ; 
        RECT 0.02 158.348 66.116 158.868 ; 
        RECT 65.648 154.494 66.116 158.868 ; 
        RECT 37.208 157.964 65.576 158.868 ; 
        RECT 31.88 157.964 37.136 158.868 ; 
        RECT 29 154.494 31.52 158.868 ; 
        RECT 0.56 157.964 28.928 158.868 ; 
        RECT 0.02 154.494 0.488 158.868 ; 
        RECT 65.504 154.494 66.116 158.156 ; 
        RECT 37.424 154.494 65.432 158.868 ; 
        RECT 34.436 154.494 37.352 158.156 ; 
        RECT 33.788 155.276 34.292 158.868 ; 
        RECT 28.784 154.892 33.68 158.156 ; 
        RECT 0.704 154.494 28.712 158.868 ; 
        RECT 0.02 154.494 0.632 158.156 ; 
        RECT 34.22 154.494 66.116 157.772 ; 
        RECT 0.02 154.892 34.148 157.772 ; 
        RECT 33.32 154.494 66.116 155.18 ; 
        RECT 0.02 154.494 33.248 157.772 ; 
        RECT 0.02 154.494 66.116 154.796 ; 
        RECT 0.02 162.668 66.116 163.188 ; 
        RECT 65.648 158.814 66.116 163.188 ; 
        RECT 37.208 162.284 65.576 163.188 ; 
        RECT 31.88 162.284 37.136 163.188 ; 
        RECT 29 158.814 31.52 163.188 ; 
        RECT 0.56 162.284 28.928 163.188 ; 
        RECT 0.02 158.814 0.488 163.188 ; 
        RECT 65.504 158.814 66.116 162.476 ; 
        RECT 37.424 158.814 65.432 163.188 ; 
        RECT 34.436 158.814 37.352 162.476 ; 
        RECT 33.788 159.596 34.292 163.188 ; 
        RECT 28.784 159.212 33.68 162.476 ; 
        RECT 0.704 158.814 28.712 163.188 ; 
        RECT 0.02 158.814 0.632 162.476 ; 
        RECT 34.22 158.814 66.116 162.092 ; 
        RECT 0.02 159.212 34.148 162.092 ; 
        RECT 33.32 158.814 66.116 159.5 ; 
        RECT 0.02 158.814 33.248 162.092 ; 
        RECT 0.02 158.814 66.116 159.116 ; 
        RECT 0.02 166.988 66.116 167.508 ; 
        RECT 65.648 163.134 66.116 167.508 ; 
        RECT 37.208 166.604 65.576 167.508 ; 
        RECT 31.88 166.604 37.136 167.508 ; 
        RECT 29 163.134 31.52 167.508 ; 
        RECT 0.56 166.604 28.928 167.508 ; 
        RECT 0.02 163.134 0.488 167.508 ; 
        RECT 65.504 163.134 66.116 166.796 ; 
        RECT 37.424 163.134 65.432 167.508 ; 
        RECT 34.436 163.134 37.352 166.796 ; 
        RECT 33.788 163.916 34.292 167.508 ; 
        RECT 28.784 163.532 33.68 166.796 ; 
        RECT 0.704 163.134 28.712 167.508 ; 
        RECT 0.02 163.134 0.632 166.796 ; 
        RECT 34.22 163.134 66.116 166.412 ; 
        RECT 0.02 163.532 34.148 166.412 ; 
        RECT 33.32 163.134 66.116 163.82 ; 
        RECT 0.02 163.134 33.248 166.412 ; 
        RECT 0.02 163.134 66.116 163.436 ; 
        RECT 0.02 171.308 66.116 171.828 ; 
        RECT 65.648 167.454 66.116 171.828 ; 
        RECT 37.208 170.924 65.576 171.828 ; 
        RECT 31.88 170.924 37.136 171.828 ; 
        RECT 29 167.454 31.52 171.828 ; 
        RECT 0.56 170.924 28.928 171.828 ; 
        RECT 0.02 167.454 0.488 171.828 ; 
        RECT 65.504 167.454 66.116 171.116 ; 
        RECT 37.424 167.454 65.432 171.828 ; 
        RECT 34.436 167.454 37.352 171.116 ; 
        RECT 33.788 168.236 34.292 171.828 ; 
        RECT 28.784 167.852 33.68 171.116 ; 
        RECT 0.704 167.454 28.712 171.828 ; 
        RECT 0.02 167.454 0.632 171.116 ; 
        RECT 34.22 167.454 66.116 170.732 ; 
        RECT 0.02 167.852 34.148 170.732 ; 
        RECT 33.32 167.454 66.116 168.14 ; 
        RECT 0.02 167.454 33.248 170.732 ; 
        RECT 0.02 167.454 66.116 167.756 ; 
        RECT 0.02 175.628 66.116 176.148 ; 
        RECT 65.648 171.774 66.116 176.148 ; 
        RECT 37.208 175.244 65.576 176.148 ; 
        RECT 31.88 175.244 37.136 176.148 ; 
        RECT 29 171.774 31.52 176.148 ; 
        RECT 0.56 175.244 28.928 176.148 ; 
        RECT 0.02 171.774 0.488 176.148 ; 
        RECT 65.504 171.774 66.116 175.436 ; 
        RECT 37.424 171.774 65.432 176.148 ; 
        RECT 34.436 171.774 37.352 175.436 ; 
        RECT 33.788 172.556 34.292 176.148 ; 
        RECT 28.784 172.172 33.68 175.436 ; 
        RECT 0.704 171.774 28.712 176.148 ; 
        RECT 0.02 171.774 0.632 175.436 ; 
        RECT 34.22 171.774 66.116 175.052 ; 
        RECT 0.02 172.172 34.148 175.052 ; 
        RECT 33.32 171.774 66.116 172.46 ; 
        RECT 0.02 171.774 33.248 175.052 ; 
        RECT 0.02 171.774 66.116 172.076 ; 
        RECT 0.02 179.948 66.116 180.468 ; 
        RECT 65.648 176.094 66.116 180.468 ; 
        RECT 37.208 179.564 65.576 180.468 ; 
        RECT 31.88 179.564 37.136 180.468 ; 
        RECT 29 176.094 31.52 180.468 ; 
        RECT 0.56 179.564 28.928 180.468 ; 
        RECT 0.02 176.094 0.488 180.468 ; 
        RECT 65.504 176.094 66.116 179.756 ; 
        RECT 37.424 176.094 65.432 180.468 ; 
        RECT 34.436 176.094 37.352 179.756 ; 
        RECT 33.788 176.876 34.292 180.468 ; 
        RECT 28.784 176.492 33.68 179.756 ; 
        RECT 0.704 176.094 28.712 180.468 ; 
        RECT 0.02 176.094 0.632 179.756 ; 
        RECT 34.22 176.094 66.116 179.372 ; 
        RECT 0.02 176.492 34.148 179.372 ; 
        RECT 33.32 176.094 66.116 176.78 ; 
        RECT 0.02 176.094 33.248 179.372 ; 
        RECT 0.02 176.094 66.116 176.396 ; 
        RECT 0.02 184.268 66.116 184.788 ; 
        RECT 65.648 180.414 66.116 184.788 ; 
        RECT 37.208 183.884 65.576 184.788 ; 
        RECT 31.88 183.884 37.136 184.788 ; 
        RECT 29 180.414 31.52 184.788 ; 
        RECT 0.56 183.884 28.928 184.788 ; 
        RECT 0.02 180.414 0.488 184.788 ; 
        RECT 65.504 180.414 66.116 184.076 ; 
        RECT 37.424 180.414 65.432 184.788 ; 
        RECT 34.436 180.414 37.352 184.076 ; 
        RECT 33.788 181.196 34.292 184.788 ; 
        RECT 28.784 180.812 33.68 184.076 ; 
        RECT 0.704 180.414 28.712 184.788 ; 
        RECT 0.02 180.414 0.632 184.076 ; 
        RECT 34.22 180.414 66.116 183.692 ; 
        RECT 0.02 180.812 34.148 183.692 ; 
        RECT 33.32 180.414 66.116 181.1 ; 
        RECT 0.02 180.414 33.248 183.692 ; 
        RECT 0.02 180.414 66.116 180.716 ; 
        RECT 0.02 188.588 66.116 189.108 ; 
        RECT 65.648 184.734 66.116 189.108 ; 
        RECT 37.208 188.204 65.576 189.108 ; 
        RECT 31.88 188.204 37.136 189.108 ; 
        RECT 29 184.734 31.52 189.108 ; 
        RECT 0.56 188.204 28.928 189.108 ; 
        RECT 0.02 184.734 0.488 189.108 ; 
        RECT 65.504 184.734 66.116 188.396 ; 
        RECT 37.424 184.734 65.432 189.108 ; 
        RECT 34.436 184.734 37.352 188.396 ; 
        RECT 33.788 185.516 34.292 189.108 ; 
        RECT 28.784 185.132 33.68 188.396 ; 
        RECT 0.704 184.734 28.712 189.108 ; 
        RECT 0.02 184.734 0.632 188.396 ; 
        RECT 34.22 184.734 66.116 188.012 ; 
        RECT 0.02 185.132 34.148 188.012 ; 
        RECT 33.32 184.734 66.116 185.42 ; 
        RECT 0.02 184.734 33.248 188.012 ; 
        RECT 0.02 184.734 66.116 185.036 ; 
        RECT 0.02 192.908 66.116 193.428 ; 
        RECT 65.648 189.054 66.116 193.428 ; 
        RECT 37.208 192.524 65.576 193.428 ; 
        RECT 31.88 192.524 37.136 193.428 ; 
        RECT 29 189.054 31.52 193.428 ; 
        RECT 0.56 192.524 28.928 193.428 ; 
        RECT 0.02 189.054 0.488 193.428 ; 
        RECT 65.504 189.054 66.116 192.716 ; 
        RECT 37.424 189.054 65.432 193.428 ; 
        RECT 34.436 189.054 37.352 192.716 ; 
        RECT 33.788 189.836 34.292 193.428 ; 
        RECT 28.784 189.452 33.68 192.716 ; 
        RECT 0.704 189.054 28.712 193.428 ; 
        RECT 0.02 189.054 0.632 192.716 ; 
        RECT 34.22 189.054 66.116 192.332 ; 
        RECT 0.02 189.452 34.148 192.332 ; 
        RECT 33.32 189.054 66.116 189.74 ; 
        RECT 0.02 189.054 33.248 192.332 ; 
        RECT 0.02 189.054 66.116 189.356 ; 
        RECT 0.02 197.228 66.116 197.748 ; 
        RECT 65.648 193.374 66.116 197.748 ; 
        RECT 37.208 196.844 65.576 197.748 ; 
        RECT 31.88 196.844 37.136 197.748 ; 
        RECT 29 193.374 31.52 197.748 ; 
        RECT 0.56 196.844 28.928 197.748 ; 
        RECT 0.02 193.374 0.488 197.748 ; 
        RECT 65.504 193.374 66.116 197.036 ; 
        RECT 37.424 193.374 65.432 197.748 ; 
        RECT 34.436 193.374 37.352 197.036 ; 
        RECT 33.788 194.156 34.292 197.748 ; 
        RECT 28.784 193.772 33.68 197.036 ; 
        RECT 0.704 193.374 28.712 197.748 ; 
        RECT 0.02 193.374 0.632 197.036 ; 
        RECT 34.22 193.374 66.116 196.652 ; 
        RECT 0.02 193.772 34.148 196.652 ; 
        RECT 33.32 193.374 66.116 194.06 ; 
        RECT 0.02 193.374 33.248 196.652 ; 
        RECT 0.02 193.374 66.116 193.676 ; 
        RECT 0.02 201.548 66.116 202.068 ; 
        RECT 65.648 197.694 66.116 202.068 ; 
        RECT 37.208 201.164 65.576 202.068 ; 
        RECT 31.88 201.164 37.136 202.068 ; 
        RECT 29 197.694 31.52 202.068 ; 
        RECT 0.56 201.164 28.928 202.068 ; 
        RECT 0.02 197.694 0.488 202.068 ; 
        RECT 65.504 197.694 66.116 201.356 ; 
        RECT 37.424 197.694 65.432 202.068 ; 
        RECT 34.436 197.694 37.352 201.356 ; 
        RECT 33.788 198.476 34.292 202.068 ; 
        RECT 28.784 198.092 33.68 201.356 ; 
        RECT 0.704 197.694 28.712 202.068 ; 
        RECT 0.02 197.694 0.632 201.356 ; 
        RECT 34.22 197.694 66.116 200.972 ; 
        RECT 0.02 198.092 34.148 200.972 ; 
        RECT 33.32 197.694 66.116 198.38 ; 
        RECT 0.02 197.694 33.248 200.972 ; 
        RECT 0.02 197.694 66.116 197.996 ; 
        RECT 0.02 205.868 66.116 206.388 ; 
        RECT 65.648 202.014 66.116 206.388 ; 
        RECT 37.208 205.484 65.576 206.388 ; 
        RECT 31.88 205.484 37.136 206.388 ; 
        RECT 29 202.014 31.52 206.388 ; 
        RECT 0.56 205.484 28.928 206.388 ; 
        RECT 0.02 202.014 0.488 206.388 ; 
        RECT 65.504 202.014 66.116 205.676 ; 
        RECT 37.424 202.014 65.432 206.388 ; 
        RECT 34.436 202.014 37.352 205.676 ; 
        RECT 33.788 202.796 34.292 206.388 ; 
        RECT 28.784 202.412 33.68 205.676 ; 
        RECT 0.704 202.014 28.712 206.388 ; 
        RECT 0.02 202.014 0.632 205.676 ; 
        RECT 34.22 202.014 66.116 205.292 ; 
        RECT 0.02 202.412 34.148 205.292 ; 
        RECT 33.32 202.014 66.116 202.7 ; 
        RECT 0.02 202.014 33.248 205.292 ; 
        RECT 0.02 202.014 66.116 202.316 ; 
        RECT 0.02 210.188 66.116 210.708 ; 
        RECT 65.648 206.334 66.116 210.708 ; 
        RECT 37.208 209.804 65.576 210.708 ; 
        RECT 31.88 209.804 37.136 210.708 ; 
        RECT 29 206.334 31.52 210.708 ; 
        RECT 0.56 209.804 28.928 210.708 ; 
        RECT 0.02 206.334 0.488 210.708 ; 
        RECT 65.504 206.334 66.116 209.996 ; 
        RECT 37.424 206.334 65.432 210.708 ; 
        RECT 34.436 206.334 37.352 209.996 ; 
        RECT 33.788 207.116 34.292 210.708 ; 
        RECT 28.784 206.732 33.68 209.996 ; 
        RECT 0.704 206.334 28.712 210.708 ; 
        RECT 0.02 206.334 0.632 209.996 ; 
        RECT 34.22 206.334 66.116 209.612 ; 
        RECT 0.02 206.732 34.148 209.612 ; 
        RECT 33.32 206.334 66.116 207.02 ; 
        RECT 0.02 206.334 33.248 209.612 ; 
        RECT 0.02 206.334 66.116 206.636 ; 
        RECT 0.02 214.508 66.116 215.028 ; 
        RECT 65.648 210.654 66.116 215.028 ; 
        RECT 37.208 214.124 65.576 215.028 ; 
        RECT 31.88 214.124 37.136 215.028 ; 
        RECT 29 210.654 31.52 215.028 ; 
        RECT 0.56 214.124 28.928 215.028 ; 
        RECT 0.02 210.654 0.488 215.028 ; 
        RECT 65.504 210.654 66.116 214.316 ; 
        RECT 37.424 210.654 65.432 215.028 ; 
        RECT 34.436 210.654 37.352 214.316 ; 
        RECT 33.788 211.436 34.292 215.028 ; 
        RECT 28.784 211.052 33.68 214.316 ; 
        RECT 0.704 210.654 28.712 215.028 ; 
        RECT 0.02 210.654 0.632 214.316 ; 
        RECT 34.22 210.654 66.116 213.932 ; 
        RECT 0.02 211.052 34.148 213.932 ; 
        RECT 33.32 210.654 66.116 211.34 ; 
        RECT 0.02 210.654 33.248 213.932 ; 
        RECT 0.02 210.654 66.116 210.956 ; 
        RECT 0.02 218.828 66.116 219.348 ; 
        RECT 65.648 214.974 66.116 219.348 ; 
        RECT 37.208 218.444 65.576 219.348 ; 
        RECT 31.88 218.444 37.136 219.348 ; 
        RECT 29 214.974 31.52 219.348 ; 
        RECT 0.56 218.444 28.928 219.348 ; 
        RECT 0.02 214.974 0.488 219.348 ; 
        RECT 65.504 214.974 66.116 218.636 ; 
        RECT 37.424 214.974 65.432 219.348 ; 
        RECT 34.436 214.974 37.352 218.636 ; 
        RECT 33.788 215.756 34.292 219.348 ; 
        RECT 28.784 215.372 33.68 218.636 ; 
        RECT 0.704 214.974 28.712 219.348 ; 
        RECT 0.02 214.974 0.632 218.636 ; 
        RECT 34.22 214.974 66.116 218.252 ; 
        RECT 0.02 215.372 34.148 218.252 ; 
        RECT 33.32 214.974 66.116 215.66 ; 
        RECT 0.02 214.974 33.248 218.252 ; 
        RECT 0.02 214.974 66.116 215.276 ; 
        RECT 0.02 223.148 66.116 223.668 ; 
        RECT 65.648 219.294 66.116 223.668 ; 
        RECT 37.208 222.764 65.576 223.668 ; 
        RECT 31.88 222.764 37.136 223.668 ; 
        RECT 29 219.294 31.52 223.668 ; 
        RECT 0.56 222.764 28.928 223.668 ; 
        RECT 0.02 219.294 0.488 223.668 ; 
        RECT 65.504 219.294 66.116 222.956 ; 
        RECT 37.424 219.294 65.432 223.668 ; 
        RECT 34.436 219.294 37.352 222.956 ; 
        RECT 33.788 220.076 34.292 223.668 ; 
        RECT 28.784 219.692 33.68 222.956 ; 
        RECT 0.704 219.294 28.712 223.668 ; 
        RECT 0.02 219.294 0.632 222.956 ; 
        RECT 34.22 219.294 66.116 222.572 ; 
        RECT 0.02 219.692 34.148 222.572 ; 
        RECT 33.32 219.294 66.116 219.98 ; 
        RECT 0.02 219.294 33.248 222.572 ; 
        RECT 0.02 219.294 66.116 219.596 ; 
        RECT 0.02 227.468 66.116 227.988 ; 
        RECT 65.648 223.614 66.116 227.988 ; 
        RECT 37.208 227.084 65.576 227.988 ; 
        RECT 31.88 227.084 37.136 227.988 ; 
        RECT 29 223.614 31.52 227.988 ; 
        RECT 0.56 227.084 28.928 227.988 ; 
        RECT 0.02 223.614 0.488 227.988 ; 
        RECT 65.504 223.614 66.116 227.276 ; 
        RECT 37.424 223.614 65.432 227.988 ; 
        RECT 34.436 223.614 37.352 227.276 ; 
        RECT 33.788 224.396 34.292 227.988 ; 
        RECT 28.784 224.012 33.68 227.276 ; 
        RECT 0.704 223.614 28.712 227.988 ; 
        RECT 0.02 223.614 0.632 227.276 ; 
        RECT 34.22 223.614 66.116 226.892 ; 
        RECT 0.02 224.012 34.148 226.892 ; 
        RECT 33.32 223.614 66.116 224.3 ; 
        RECT 0.02 223.614 33.248 226.892 ; 
        RECT 0.02 223.614 66.116 223.916 ; 
        RECT 0.02 231.788 66.116 232.308 ; 
        RECT 65.648 227.934 66.116 232.308 ; 
        RECT 37.208 231.404 65.576 232.308 ; 
        RECT 31.88 231.404 37.136 232.308 ; 
        RECT 29 227.934 31.52 232.308 ; 
        RECT 0.56 231.404 28.928 232.308 ; 
        RECT 0.02 227.934 0.488 232.308 ; 
        RECT 65.504 227.934 66.116 231.596 ; 
        RECT 37.424 227.934 65.432 232.308 ; 
        RECT 34.436 227.934 37.352 231.596 ; 
        RECT 33.788 228.716 34.292 232.308 ; 
        RECT 28.784 228.332 33.68 231.596 ; 
        RECT 0.704 227.934 28.712 232.308 ; 
        RECT 0.02 227.934 0.632 231.596 ; 
        RECT 34.22 227.934 66.116 231.212 ; 
        RECT 0.02 228.332 34.148 231.212 ; 
        RECT 33.32 227.934 66.116 228.62 ; 
        RECT 0.02 227.934 33.248 231.212 ; 
        RECT 0.02 227.934 66.116 228.236 ; 
        RECT 0.02 236.108 66.116 236.628 ; 
        RECT 65.648 232.254 66.116 236.628 ; 
        RECT 37.208 235.724 65.576 236.628 ; 
        RECT 31.88 235.724 37.136 236.628 ; 
        RECT 29 232.254 31.52 236.628 ; 
        RECT 0.56 235.724 28.928 236.628 ; 
        RECT 0.02 232.254 0.488 236.628 ; 
        RECT 65.504 232.254 66.116 235.916 ; 
        RECT 37.424 232.254 65.432 236.628 ; 
        RECT 34.436 232.254 37.352 235.916 ; 
        RECT 33.788 233.036 34.292 236.628 ; 
        RECT 28.784 232.652 33.68 235.916 ; 
        RECT 0.704 232.254 28.712 236.628 ; 
        RECT 0.02 232.254 0.632 235.916 ; 
        RECT 34.22 232.254 66.116 235.532 ; 
        RECT 0.02 232.652 34.148 235.532 ; 
        RECT 33.32 232.254 66.116 232.94 ; 
        RECT 0.02 232.254 33.248 235.532 ; 
        RECT 0.02 232.254 66.116 232.556 ; 
        RECT 0.02 240.428 66.116 240.948 ; 
        RECT 65.648 236.574 66.116 240.948 ; 
        RECT 37.208 240.044 65.576 240.948 ; 
        RECT 31.88 240.044 37.136 240.948 ; 
        RECT 29 236.574 31.52 240.948 ; 
        RECT 0.56 240.044 28.928 240.948 ; 
        RECT 0.02 236.574 0.488 240.948 ; 
        RECT 65.504 236.574 66.116 240.236 ; 
        RECT 37.424 236.574 65.432 240.948 ; 
        RECT 34.436 236.574 37.352 240.236 ; 
        RECT 33.788 237.356 34.292 240.948 ; 
        RECT 28.784 236.972 33.68 240.236 ; 
        RECT 0.704 236.574 28.712 240.948 ; 
        RECT 0.02 236.574 0.632 240.236 ; 
        RECT 34.22 236.574 66.116 239.852 ; 
        RECT 0.02 236.972 34.148 239.852 ; 
        RECT 33.32 236.574 66.116 237.26 ; 
        RECT 0.02 236.574 33.248 239.852 ; 
        RECT 0.02 236.574 66.116 236.876 ; 
  LAYER M4 ; 
      RECT 6.276 111.48 60.038 111.576 ; 
      RECT 6.276 112.632 60.038 112.728 ; 
      RECT 6.276 114.168 60.038 114.264 ; 
      RECT 6.276 114.552 60.038 114.648 ; 
      RECT 6.276 115.896 60.038 115.992 ; 
      RECT 6.276 117.432 60.038 117.528 ; 
      RECT 43.82 107.316 44.156 107.412 ; 
      RECT 43.068 109.044 43.588 109.14 ; 
      RECT 43.1 111.674 43.568 111.77 ; 
      RECT 43.1 112.824 43.568 112.92 ; 
      RECT 40.544 109.044 42.828 109.14 ; 
      RECT 40.784 112.152 41.216 112.248 ; 
      RECT 35.452 113.652 39.824 113.748 ; 
      RECT 38.204 111.924 38.54 112.02 ; 
      RECT 35.068 116.724 38.54 116.82 ; 
      RECT 38.204 117.108 38.54 117.204 ; 
      RECT 37.492 110.004 37.828 110.1 ; 
      RECT 37.34 115.38 37.676 115.476 ; 
      RECT 37.34 118.26 37.676 118.356 ; 
      RECT 36.628 109.62 36.964 109.716 ; 
      RECT 35.772 104.468 36.824 104.564 ; 
      RECT 35.772 138.964 36.824 139.06 ; 
      RECT 35.836 115.572 36.812 115.668 ; 
      RECT 36.476 116.148 36.812 116.244 ; 
      RECT 30.652 117.108 36.812 117.204 ; 
      RECT 36.476 118.26 36.812 118.356 ; 
      RECT 35.54 138.58 36.592 138.676 ; 
      RECT 35.536 104.084 36.588 104.18 ; 
      RECT 35.384 103.7 36.436 103.796 ; 
      RECT 35.384 137.812 36.436 137.908 ; 
      RECT 36.044 119.988 36.38 120.084 ; 
      RECT 32.956 121.524 36.38 121.62 ; 
      RECT 34.492 130.548 36.38 130.644 ; 
      RECT 36.044 130.932 36.38 131.028 ; 
      RECT 35.192 103.316 36.244 103.412 ; 
      RECT 35.192 137.428 36.244 137.524 ; 
      RECT 34.3 126.9 36.08 126.996 ; 
      RECT 35.016 102.932 36.068 103.028 ; 
      RECT 35.016 138.772 36.068 138.868 ; 
      RECT 34.82 104.276 35.872 104.372 ; 
      RECT 34.82 138.388 35.872 138.484 ; 
      RECT 35.344 116.148 35.828 116.244 ; 
      RECT 35.26 124.596 35.792 124.692 ; 
      RECT 34.632 103.892 35.684 103.988 ; 
      RECT 34.632 138.004 35.684 138.1 ; 
      RECT 34.492 102.74 35.544 102.836 ; 
      RECT 34.492 137.62 35.544 137.716 ; 
      RECT 31.228 130.932 35.504 131.028 ; 
      RECT 35.168 135.54 35.504 135.636 ; 
      RECT 34.268 102.164 35.32 102.26 ; 
      RECT 34.268 137.236 35.32 137.332 ; 
      RECT 34.876 119.988 35.216 120.084 ; 
      RECT 30.46 122.292 34.928 122.388 ; 
      RECT 33.04 113.652 34.868 113.748 ; 
      RECT 32.348 105.044 33.416 105.14 ; 
      RECT 32.348 136.66 33.416 136.756 ; 
      RECT 32.896 119.796 33.332 119.892 ; 
      RECT 32.256 104.66 33.224 104.756 ; 
      RECT 32.256 139.156 33.224 139.252 ; 
      RECT 32.032 102.74 33 102.836 ; 
      RECT 32.148 139.54 33 139.636 ; 
      RECT 32.612 118.26 32.948 118.356 ; 
      RECT 31.816 103.124 32.808 103.22 ; 
      RECT 31.816 138.964 32.808 139.06 ; 
      RECT 30.88 128.628 32.564 128.724 ; 
      RECT 30.752 104.468 31.82 104.564 ; 
      RECT 30.752 139.54 31.82 139.636 ; 
      RECT 31.312 122.868 31.796 122.964 ; 
      RECT 31.28 135.54 31.616 135.636 ; 
      RECT 30.616 104.084 31.604 104.18 ; 
      RECT 30.348 137.812 31.604 137.908 ; 
      RECT 30.512 103.7 31.432 103.796 ; 
      RECT 30.464 139.156 31.432 139.252 ; 
      RECT 30.3 103.316 31.22 103.412 ; 
      RECT 30.884 129.204 31.22 129.3 ; 
      RECT 30.1 137.428 31.22 137.524 ; 
      RECT 30.12 102.932 31.04 103.028 ; 
      RECT 30.12 138.772 31.04 138.868 ; 
      RECT 26.272 118.26 31.028 118.356 ; 
      RECT 29.968 103.892 30.888 103.988 ; 
      RECT 29.968 138.388 30.888 138.484 ; 
      RECT 29.896 103.508 30.668 103.604 ; 
      RECT 29.896 138.004 30.668 138.1 ; 
      RECT 29.7 103.124 30.472 103.22 ; 
      RECT 29.7 137.62 30.472 137.716 ; 
      RECT 29.716 121.908 30.452 122.004 ; 
      RECT 29.492 102.74 30.264 102.836 ; 
      RECT 29.492 137.236 30.264 137.332 ; 
      RECT 27.556 111.156 30.26 111.252 ; 
      RECT 29.716 122.292 30.052 122.388 ; 
      RECT 28.64 104.852 29.692 104.948 ; 
      RECT 28.77 119.988 29.304 120.084 ; 
      RECT 27.404 111.924 27.74 112.02 ; 
  LAYER V4 ; 
      RECT 44.016 107.316 44.112 107.412 ; 
      RECT 44.016 111.48 44.112 111.576 ; 
      RECT 43.344 109.044 43.44 109.14 ; 
      RECT 43.344 111.674 43.44 111.77 ; 
      RECT 43.344 112.824 43.44 112.92 ; 
      RECT 40.848 109.044 40.944 109.14 ; 
      RECT 40.848 112.152 40.944 112.248 ; 
      RECT 38.4 111.924 38.496 112.02 ; 
      RECT 38.4 112.632 38.496 112.728 ; 
      RECT 38.4 116.724 38.496 116.82 ; 
      RECT 38.4 117.108 38.496 117.204 ; 
      RECT 37.536 110.004 37.632 110.1 ; 
      RECT 37.536 114.168 37.632 114.264 ; 
      RECT 37.536 115.38 37.632 115.476 ; 
      RECT 37.536 115.896 37.632 115.992 ; 
      RECT 37.536 117.432 37.632 117.528 ; 
      RECT 37.536 118.26 37.632 118.356 ; 
      RECT 36.672 109.62 36.768 109.716 ; 
      RECT 36.672 114.552 36.768 114.648 ; 
      RECT 36.672 115.572 36.768 115.668 ; 
      RECT 36.672 116.148 36.768 116.244 ; 
      RECT 36.672 117.108 36.768 117.204 ; 
      RECT 36.672 118.26 36.768 118.356 ; 
      RECT 36.24 119.988 36.336 120.084 ; 
      RECT 36.24 121.524 36.336 121.62 ; 
      RECT 36.24 130.548 36.336 130.644 ; 
      RECT 36.24 130.932 36.336 131.028 ; 
      RECT 35.88 104.468 35.976 104.564 ; 
      RECT 35.88 115.572 35.976 115.668 ; 
      RECT 35.88 138.964 35.976 139.06 ; 
      RECT 35.688 104.084 35.784 104.18 ; 
      RECT 35.688 116.148 35.784 116.244 ; 
      RECT 35.688 138.58 35.784 138.676 ; 
      RECT 35.496 103.7 35.592 103.796 ; 
      RECT 35.496 113.652 35.592 113.748 ; 
      RECT 35.496 137.812 35.592 137.908 ; 
      RECT 35.304 103.316 35.4 103.412 ; 
      RECT 35.304 124.596 35.4 124.692 ; 
      RECT 35.304 135.54 35.4 135.636 ; 
      RECT 35.304 137.428 35.4 137.524 ; 
      RECT 35.112 102.932 35.208 103.028 ; 
      RECT 35.112 116.724 35.208 116.82 ; 
      RECT 35.112 138.772 35.208 138.868 ; 
      RECT 34.92 104.276 35.016 104.372 ; 
      RECT 34.92 119.988 35.016 120.084 ; 
      RECT 34.92 138.388 35.016 138.484 ; 
      RECT 34.728 103.892 34.824 103.988 ; 
      RECT 34.728 113.652 34.824 113.748 ; 
      RECT 34.728 138.004 34.824 138.1 ; 
      RECT 34.536 102.74 34.632 102.836 ; 
      RECT 34.536 130.548 34.632 130.644 ; 
      RECT 34.536 137.62 34.632 137.716 ; 
      RECT 34.344 102.164 34.44 102.26 ; 
      RECT 34.344 126.9 34.44 126.996 ; 
      RECT 34.344 137.236 34.44 137.332 ; 
      RECT 33.192 105.044 33.288 105.14 ; 
      RECT 33.192 119.796 33.288 119.892 ; 
      RECT 33.192 136.66 33.288 136.756 ; 
      RECT 33 104.66 33.096 104.756 ; 
      RECT 33 121.524 33.096 121.62 ; 
      RECT 33 139.156 33.096 139.252 ; 
      RECT 32.808 102.74 32.904 102.836 ; 
      RECT 32.808 118.26 32.904 118.356 ; 
      RECT 32.808 139.54 32.904 139.636 ; 
      RECT 32.424 103.124 32.52 103.22 ; 
      RECT 32.424 128.628 32.52 128.724 ; 
      RECT 32.424 138.964 32.52 139.06 ; 
      RECT 31.656 104.468 31.752 104.564 ; 
      RECT 31.656 122.868 31.752 122.964 ; 
      RECT 31.656 139.54 31.752 139.636 ; 
      RECT 31.464 104.084 31.56 104.18 ; 
      RECT 31.464 135.54 31.56 135.636 ; 
      RECT 31.464 137.812 31.56 137.908 ; 
      RECT 31.272 103.7 31.368 103.796 ; 
      RECT 31.272 130.932 31.368 131.028 ; 
      RECT 31.272 139.156 31.368 139.252 ; 
      RECT 31.08 103.316 31.176 103.412 ; 
      RECT 31.08 129.204 31.176 129.3 ; 
      RECT 31.08 137.428 31.176 137.524 ; 
      RECT 30.888 102.932 30.984 103.028 ; 
      RECT 30.888 118.26 30.984 118.356 ; 
      RECT 30.888 138.772 30.984 138.868 ; 
      RECT 30.696 103.892 30.792 103.988 ; 
      RECT 30.696 117.108 30.792 117.204 ; 
      RECT 30.696 138.388 30.792 138.484 ; 
      RECT 30.504 103.508 30.6 103.604 ; 
      RECT 30.504 122.292 30.6 122.388 ; 
      RECT 30.504 138.004 30.6 138.1 ; 
      RECT 30.312 103.124 30.408 103.22 ; 
      RECT 30.312 121.908 30.408 122.004 ; 
      RECT 30.312 137.62 30.408 137.716 ; 
      RECT 30.12 102.74 30.216 102.836 ; 
      RECT 30.12 111.156 30.216 111.252 ; 
      RECT 30.12 137.236 30.216 137.332 ; 
      RECT 29.76 121.908 29.856 122.004 ; 
      RECT 29.76 122.292 29.856 122.388 ; 
      RECT 29.088 104.852 29.184 104.948 ; 
      RECT 29.088 119.988 29.184 120.084 ; 
      RECT 27.6 111.156 27.696 111.252 ; 
      RECT 27.6 111.924 27.696 112.02 ; 
  LAYER M5 ; 
      RECT 44.016 107.272 44.112 111.62 ; 
      RECT 43.344 108.932 43.44 113.174 ; 
      RECT 40.848 108.966 40.944 112.296 ; 
      RECT 38.4 111.88 38.496 112.772 ; 
      RECT 38.4 116.68 38.496 117.248 ; 
      RECT 37.536 109.96 37.632 114.308 ; 
      RECT 37.536 115.336 37.632 116.036 ; 
      RECT 37.536 117.388 37.632 118.4 ; 
      RECT 36.672 109.576 36.768 114.692 ; 
      RECT 36.672 115.528 36.768 116.288 ; 
      RECT 36.672 117.064 36.768 118.4 ; 
      RECT 36.24 119.944 36.336 121.664 ; 
      RECT 36.24 130.504 36.336 131.072 ; 
      RECT 35.88 105.816 35.976 136.148 ; 
      RECT 35.688 105.816 35.784 136.148 ; 
      RECT 35.496 105.816 35.592 136.148 ; 
      RECT 35.304 105.816 35.4 136.148 ; 
      RECT 35.112 105.816 35.208 136.148 ; 
      RECT 34.92 105.816 35.016 136.148 ; 
      RECT 34.728 105.816 34.824 136.148 ; 
      RECT 34.536 105.816 34.632 136.148 ; 
      RECT 34.344 105.816 34.44 136.148 ; 
      RECT 33.192 105.816 33.288 136.148 ; 
      RECT 33 105.816 33.096 136.148 ; 
      RECT 32.808 105.816 32.904 136.148 ; 
      RECT 32.424 105.816 32.52 136.148 ; 
      RECT 31.656 105.816 31.752 136.148 ; 
      RECT 31.464 105.816 31.56 136.148 ; 
      RECT 31.272 105.816 31.368 136.148 ; 
      RECT 31.08 105.816 31.176 136.148 ; 
      RECT 30.888 105.816 30.984 136.148 ; 
      RECT 30.696 105.816 30.792 136.148 ; 
      RECT 30.504 102.448 30.6 138.668 ; 
      RECT 30.312 102.3 30.408 138.484 ; 
      RECT 30.12 102.084 30.216 138.268 ; 
      RECT 29.76 121.864 29.856 122.432 ; 
      RECT 29.088 104.78 29.184 120.156 ; 
      RECT 27.6 111.112 27.696 112.064 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 63.568 241.776 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 63.568 241.776 ; 
  END 
END srambank_128x4x48_6t122 
