VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_128x4x74_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_128x4x74_6t122 0 0 ;
  SIZE 16.0 BY 88.56 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.1720 16.4420 1.2200 ;
        RECT 0.0940 2.2520 16.4420 2.3000 ;
        RECT 0.0940 3.3320 16.4420 3.3800 ;
        RECT 0.0940 4.4120 16.4420 4.4600 ;
        RECT 0.0940 5.4920 16.4420 5.5400 ;
        RECT 0.0940 6.5720 16.4420 6.6200 ;
        RECT 0.0940 7.6520 16.4420 7.7000 ;
        RECT 0.0940 8.7320 16.4420 8.7800 ;
        RECT 0.0940 9.8120 16.4420 9.8600 ;
        RECT 0.0940 10.8920 16.4420 10.9400 ;
        RECT 0.0940 11.9720 16.4420 12.0200 ;
        RECT 0.0940 13.0520 16.4420 13.1000 ;
        RECT 0.0940 14.1320 16.4420 14.1800 ;
        RECT 0.0940 15.2120 16.4420 15.2600 ;
        RECT 0.0940 16.2920 16.4420 16.3400 ;
        RECT 0.0940 17.3720 16.4420 17.4200 ;
        RECT 0.0940 18.4520 16.4420 18.5000 ;
        RECT 0.0940 19.5320 16.4420 19.5800 ;
        RECT 0.0940 20.6120 16.4420 20.6600 ;
        RECT 0.0940 21.6920 16.4420 21.7400 ;
        RECT 0.0940 22.7720 16.4420 22.8200 ;
        RECT 0.0940 23.8520 16.4420 23.9000 ;
        RECT 0.0940 24.9320 16.4420 24.9800 ;
        RECT 0.0940 26.0120 16.4420 26.0600 ;
        RECT 0.0940 27.0920 16.4420 27.1400 ;
        RECT 0.0940 28.1720 16.4420 28.2200 ;
        RECT 0.0940 29.2520 16.4420 29.3000 ;
        RECT 0.0940 30.3320 16.4420 30.3800 ;
        RECT 0.0940 31.4120 16.4420 31.4600 ;
        RECT 0.0940 32.4920 16.4420 32.5400 ;
        RECT 0.0940 33.5720 16.4420 33.6200 ;
        RECT 0.0940 34.6520 16.4420 34.7000 ;
        RECT 0.0940 35.7320 16.4420 35.7800 ;
        RECT 0.0940 36.8120 16.4420 36.8600 ;
        RECT 0.0940 37.8920 16.4420 37.9400 ;
        RECT 0.0940 38.9720 16.4420 39.0200 ;
        RECT 0.0940 40.0520 16.4420 40.1000 ;
        RECT 3.5640 40.5330 12.9600 40.7490 ;
        RECT 9.1970 44.0370 9.3380 44.0610 ;
        RECT 9.0660 40.2530 9.3290 40.2770 ;
        RECT 7.3980 43.7010 9.1260 43.9170 ;
        RECT 7.3980 46.8690 9.1260 47.0850 ;
        RECT 0.0940 49.2590 16.4420 49.3070 ;
        RECT 0.0940 50.3390 16.4420 50.3870 ;
        RECT 0.0940 51.4190 16.4420 51.4670 ;
        RECT 0.0940 52.4990 16.4420 52.5470 ;
        RECT 0.0940 53.5790 16.4420 53.6270 ;
        RECT 0.0940 54.6590 16.4420 54.7070 ;
        RECT 0.0940 55.7390 16.4420 55.7870 ;
        RECT 0.0940 56.8190 16.4420 56.8670 ;
        RECT 0.0940 57.8990 16.4420 57.9470 ;
        RECT 0.0940 58.9790 16.4420 59.0270 ;
        RECT 0.0940 60.0590 16.4420 60.1070 ;
        RECT 0.0940 61.1390 16.4420 61.1870 ;
        RECT 0.0940 62.2190 16.4420 62.2670 ;
        RECT 0.0940 63.2990 16.4420 63.3470 ;
        RECT 0.0940 64.3790 16.4420 64.4270 ;
        RECT 0.0940 65.4590 16.4420 65.5070 ;
        RECT 0.0940 66.5390 16.4420 66.5870 ;
        RECT 0.0940 67.6190 16.4420 67.6670 ;
        RECT 0.0940 68.6990 16.4420 68.7470 ;
        RECT 0.0940 69.7790 16.4420 69.8270 ;
        RECT 0.0940 70.8590 16.4420 70.9070 ;
        RECT 0.0940 71.9390 16.4420 71.9870 ;
        RECT 0.0940 73.0190 16.4420 73.0670 ;
        RECT 0.0940 74.0990 16.4420 74.1470 ;
        RECT 0.0940 75.1790 16.4420 75.2270 ;
        RECT 0.0940 76.2590 16.4420 76.3070 ;
        RECT 0.0940 77.3390 16.4420 77.3870 ;
        RECT 0.0940 78.4190 16.4420 78.4670 ;
        RECT 0.0940 79.4990 16.4420 79.5470 ;
        RECT 0.0940 80.5790 16.4420 80.6270 ;
        RECT 0.0940 81.6590 16.4420 81.7070 ;
        RECT 0.0940 82.7390 16.4420 82.7870 ;
        RECT 0.0940 83.8190 16.4420 83.8670 ;
        RECT 0.0940 84.8990 16.4420 84.9470 ;
        RECT 0.0940 85.9790 16.4420 86.0270 ;
        RECT 0.0940 87.0590 16.4420 87.1070 ;
        RECT 0.0940 88.1390 16.4420 88.1870 ;
      LAYER M3  ;
        RECT 16.3940 0.2165 16.4120 1.3765 ;
        RECT 9.2840 0.2170 9.3020 1.3760 ;
        RECT 7.8800 0.2570 7.9700 1.3710 ;
        RECT 7.2320 0.2170 7.2500 1.3760 ;
        RECT 0.1220 0.2165 0.1400 1.3765 ;
        RECT 16.3940 1.2965 16.4120 2.4565 ;
        RECT 9.2840 1.2970 9.3020 2.4560 ;
        RECT 7.8800 1.3370 7.9700 2.4510 ;
        RECT 7.2320 1.2970 7.2500 2.4560 ;
        RECT 0.1220 1.2965 0.1400 2.4565 ;
        RECT 16.3940 2.3765 16.4120 3.5365 ;
        RECT 9.2840 2.3770 9.3020 3.5360 ;
        RECT 7.8800 2.4170 7.9700 3.5310 ;
        RECT 7.2320 2.3770 7.2500 3.5360 ;
        RECT 0.1220 2.3765 0.1400 3.5365 ;
        RECT 16.3940 3.4565 16.4120 4.6165 ;
        RECT 9.2840 3.4570 9.3020 4.6160 ;
        RECT 7.8800 3.4970 7.9700 4.6110 ;
        RECT 7.2320 3.4570 7.2500 4.6160 ;
        RECT 0.1220 3.4565 0.1400 4.6165 ;
        RECT 16.3940 4.5365 16.4120 5.6965 ;
        RECT 9.2840 4.5370 9.3020 5.6960 ;
        RECT 7.8800 4.5770 7.9700 5.6910 ;
        RECT 7.2320 4.5370 7.2500 5.6960 ;
        RECT 0.1220 4.5365 0.1400 5.6965 ;
        RECT 16.3940 5.6165 16.4120 6.7765 ;
        RECT 9.2840 5.6170 9.3020 6.7760 ;
        RECT 7.8800 5.6570 7.9700 6.7710 ;
        RECT 7.2320 5.6170 7.2500 6.7760 ;
        RECT 0.1220 5.6165 0.1400 6.7765 ;
        RECT 16.3940 6.6965 16.4120 7.8565 ;
        RECT 9.2840 6.6970 9.3020 7.8560 ;
        RECT 7.8800 6.7370 7.9700 7.8510 ;
        RECT 7.2320 6.6970 7.2500 7.8560 ;
        RECT 0.1220 6.6965 0.1400 7.8565 ;
        RECT 16.3940 7.7765 16.4120 8.9365 ;
        RECT 9.2840 7.7770 9.3020 8.9360 ;
        RECT 7.8800 7.8170 7.9700 8.9310 ;
        RECT 7.2320 7.7770 7.2500 8.9360 ;
        RECT 0.1220 7.7765 0.1400 8.9365 ;
        RECT 16.3940 8.8565 16.4120 10.0165 ;
        RECT 9.2840 8.8570 9.3020 10.0160 ;
        RECT 7.8800 8.8970 7.9700 10.0110 ;
        RECT 7.2320 8.8570 7.2500 10.0160 ;
        RECT 0.1220 8.8565 0.1400 10.0165 ;
        RECT 16.3940 9.9365 16.4120 11.0965 ;
        RECT 9.2840 9.9370 9.3020 11.0960 ;
        RECT 7.8800 9.9770 7.9700 11.0910 ;
        RECT 7.2320 9.9370 7.2500 11.0960 ;
        RECT 0.1220 9.9365 0.1400 11.0965 ;
        RECT 16.3940 11.0165 16.4120 12.1765 ;
        RECT 9.2840 11.0170 9.3020 12.1760 ;
        RECT 7.8800 11.0570 7.9700 12.1710 ;
        RECT 7.2320 11.0170 7.2500 12.1760 ;
        RECT 0.1220 11.0165 0.1400 12.1765 ;
        RECT 16.3940 12.0965 16.4120 13.2565 ;
        RECT 9.2840 12.0970 9.3020 13.2560 ;
        RECT 7.8800 12.1370 7.9700 13.2510 ;
        RECT 7.2320 12.0970 7.2500 13.2560 ;
        RECT 0.1220 12.0965 0.1400 13.2565 ;
        RECT 16.3940 13.1765 16.4120 14.3365 ;
        RECT 9.2840 13.1770 9.3020 14.3360 ;
        RECT 7.8800 13.2170 7.9700 14.3310 ;
        RECT 7.2320 13.1770 7.2500 14.3360 ;
        RECT 0.1220 13.1765 0.1400 14.3365 ;
        RECT 16.3940 14.2565 16.4120 15.4165 ;
        RECT 9.2840 14.2570 9.3020 15.4160 ;
        RECT 7.8800 14.2970 7.9700 15.4110 ;
        RECT 7.2320 14.2570 7.2500 15.4160 ;
        RECT 0.1220 14.2565 0.1400 15.4165 ;
        RECT 16.3940 15.3365 16.4120 16.4965 ;
        RECT 9.2840 15.3370 9.3020 16.4960 ;
        RECT 7.8800 15.3770 7.9700 16.4910 ;
        RECT 7.2320 15.3370 7.2500 16.4960 ;
        RECT 0.1220 15.3365 0.1400 16.4965 ;
        RECT 16.3940 16.4165 16.4120 17.5765 ;
        RECT 9.2840 16.4170 9.3020 17.5760 ;
        RECT 7.8800 16.4570 7.9700 17.5710 ;
        RECT 7.2320 16.4170 7.2500 17.5760 ;
        RECT 0.1220 16.4165 0.1400 17.5765 ;
        RECT 16.3940 17.4965 16.4120 18.6565 ;
        RECT 9.2840 17.4970 9.3020 18.6560 ;
        RECT 7.8800 17.5370 7.9700 18.6510 ;
        RECT 7.2320 17.4970 7.2500 18.6560 ;
        RECT 0.1220 17.4965 0.1400 18.6565 ;
        RECT 16.3940 18.5765 16.4120 19.7365 ;
        RECT 9.2840 18.5770 9.3020 19.7360 ;
        RECT 7.8800 18.6170 7.9700 19.7310 ;
        RECT 7.2320 18.5770 7.2500 19.7360 ;
        RECT 0.1220 18.5765 0.1400 19.7365 ;
        RECT 16.3940 19.6565 16.4120 20.8165 ;
        RECT 9.2840 19.6570 9.3020 20.8160 ;
        RECT 7.8800 19.6970 7.9700 20.8110 ;
        RECT 7.2320 19.6570 7.2500 20.8160 ;
        RECT 0.1220 19.6565 0.1400 20.8165 ;
        RECT 16.3940 20.7365 16.4120 21.8965 ;
        RECT 9.2840 20.7370 9.3020 21.8960 ;
        RECT 7.8800 20.7770 7.9700 21.8910 ;
        RECT 7.2320 20.7370 7.2500 21.8960 ;
        RECT 0.1220 20.7365 0.1400 21.8965 ;
        RECT 16.3940 21.8165 16.4120 22.9765 ;
        RECT 9.2840 21.8170 9.3020 22.9760 ;
        RECT 7.8800 21.8570 7.9700 22.9710 ;
        RECT 7.2320 21.8170 7.2500 22.9760 ;
        RECT 0.1220 21.8165 0.1400 22.9765 ;
        RECT 16.3940 22.8965 16.4120 24.0565 ;
        RECT 9.2840 22.8970 9.3020 24.0560 ;
        RECT 7.8800 22.9370 7.9700 24.0510 ;
        RECT 7.2320 22.8970 7.2500 24.0560 ;
        RECT 0.1220 22.8965 0.1400 24.0565 ;
        RECT 16.3940 23.9765 16.4120 25.1365 ;
        RECT 9.2840 23.9770 9.3020 25.1360 ;
        RECT 7.8800 24.0170 7.9700 25.1310 ;
        RECT 7.2320 23.9770 7.2500 25.1360 ;
        RECT 0.1220 23.9765 0.1400 25.1365 ;
        RECT 16.3940 25.0565 16.4120 26.2165 ;
        RECT 9.2840 25.0570 9.3020 26.2160 ;
        RECT 7.8800 25.0970 7.9700 26.2110 ;
        RECT 7.2320 25.0570 7.2500 26.2160 ;
        RECT 0.1220 25.0565 0.1400 26.2165 ;
        RECT 16.3940 26.1365 16.4120 27.2965 ;
        RECT 9.2840 26.1370 9.3020 27.2960 ;
        RECT 7.8800 26.1770 7.9700 27.2910 ;
        RECT 7.2320 26.1370 7.2500 27.2960 ;
        RECT 0.1220 26.1365 0.1400 27.2965 ;
        RECT 16.3940 27.2165 16.4120 28.3765 ;
        RECT 9.2840 27.2170 9.3020 28.3760 ;
        RECT 7.8800 27.2570 7.9700 28.3710 ;
        RECT 7.2320 27.2170 7.2500 28.3760 ;
        RECT 0.1220 27.2165 0.1400 28.3765 ;
        RECT 16.3940 28.2965 16.4120 29.4565 ;
        RECT 9.2840 28.2970 9.3020 29.4560 ;
        RECT 7.8800 28.3370 7.9700 29.4510 ;
        RECT 7.2320 28.2970 7.2500 29.4560 ;
        RECT 0.1220 28.2965 0.1400 29.4565 ;
        RECT 16.3940 29.3765 16.4120 30.5365 ;
        RECT 9.2840 29.3770 9.3020 30.5360 ;
        RECT 7.8800 29.4170 7.9700 30.5310 ;
        RECT 7.2320 29.3770 7.2500 30.5360 ;
        RECT 0.1220 29.3765 0.1400 30.5365 ;
        RECT 16.3940 30.4565 16.4120 31.6165 ;
        RECT 9.2840 30.4570 9.3020 31.6160 ;
        RECT 7.8800 30.4970 7.9700 31.6110 ;
        RECT 7.2320 30.4570 7.2500 31.6160 ;
        RECT 0.1220 30.4565 0.1400 31.6165 ;
        RECT 16.3940 31.5365 16.4120 32.6965 ;
        RECT 9.2840 31.5370 9.3020 32.6960 ;
        RECT 7.8800 31.5770 7.9700 32.6910 ;
        RECT 7.2320 31.5370 7.2500 32.6960 ;
        RECT 0.1220 31.5365 0.1400 32.6965 ;
        RECT 16.3940 32.6165 16.4120 33.7765 ;
        RECT 9.2840 32.6170 9.3020 33.7760 ;
        RECT 7.8800 32.6570 7.9700 33.7710 ;
        RECT 7.2320 32.6170 7.2500 33.7760 ;
        RECT 0.1220 32.6165 0.1400 33.7765 ;
        RECT 16.3940 33.6965 16.4120 34.8565 ;
        RECT 9.2840 33.6970 9.3020 34.8560 ;
        RECT 7.8800 33.7370 7.9700 34.8510 ;
        RECT 7.2320 33.6970 7.2500 34.8560 ;
        RECT 0.1220 33.6965 0.1400 34.8565 ;
        RECT 16.3940 34.7765 16.4120 35.9365 ;
        RECT 9.2840 34.7770 9.3020 35.9360 ;
        RECT 7.8800 34.8170 7.9700 35.9310 ;
        RECT 7.2320 34.7770 7.2500 35.9360 ;
        RECT 0.1220 34.7765 0.1400 35.9365 ;
        RECT 16.3940 35.8565 16.4120 37.0165 ;
        RECT 9.2840 35.8570 9.3020 37.0160 ;
        RECT 7.8800 35.8970 7.9700 37.0110 ;
        RECT 7.2320 35.8570 7.2500 37.0160 ;
        RECT 0.1220 35.8565 0.1400 37.0165 ;
        RECT 16.3940 36.9365 16.4120 38.0965 ;
        RECT 9.2840 36.9370 9.3020 38.0960 ;
        RECT 7.8800 36.9770 7.9700 38.0910 ;
        RECT 7.2320 36.9370 7.2500 38.0960 ;
        RECT 0.1220 36.9365 0.1400 38.0965 ;
        RECT 16.3940 38.0165 16.4120 39.1765 ;
        RECT 9.2840 38.0170 9.3020 39.1760 ;
        RECT 7.8800 38.0570 7.9700 39.1710 ;
        RECT 7.2320 38.0170 7.2500 39.1760 ;
        RECT 0.1220 38.0165 0.1400 39.1765 ;
        RECT 16.3940 39.0965 16.4120 40.2565 ;
        RECT 9.2840 39.0970 9.3020 40.2560 ;
        RECT 7.8800 39.1370 7.9700 40.2510 ;
        RECT 7.2320 39.0970 7.2500 40.2560 ;
        RECT 0.1220 39.0965 0.1400 40.2565 ;
        RECT 16.3890 40.1705 16.4070 48.3775 ;
        RECT 9.2970 43.9900 9.3150 48.3385 ;
        RECT 9.2790 40.2035 9.2970 40.3415 ;
        RECT 7.9110 40.4940 8.1450 48.0770 ;
        RECT 7.8750 47.9940 7.9650 48.3700 ;
        RECT 7.8750 40.2100 7.9650 40.5860 ;
        RECT 0.1170 40.1705 0.1350 48.3775 ;
        RECT 16.3940 48.3035 16.4120 49.4635 ;
        RECT 9.2840 48.3040 9.3020 49.4630 ;
        RECT 7.8800 48.3440 7.9700 49.4580 ;
        RECT 7.2320 48.3040 7.2500 49.4630 ;
        RECT 0.1220 48.3035 0.1400 49.4635 ;
        RECT 16.3940 49.3835 16.4120 50.5435 ;
        RECT 9.2840 49.3840 9.3020 50.5430 ;
        RECT 7.8800 49.4240 7.9700 50.5380 ;
        RECT 7.2320 49.3840 7.2500 50.5430 ;
        RECT 0.1220 49.3835 0.1400 50.5435 ;
        RECT 16.3940 50.4635 16.4120 51.6235 ;
        RECT 9.2840 50.4640 9.3020 51.6230 ;
        RECT 7.8800 50.5040 7.9700 51.6180 ;
        RECT 7.2320 50.4640 7.2500 51.6230 ;
        RECT 0.1220 50.4635 0.1400 51.6235 ;
        RECT 16.3940 51.5435 16.4120 52.7035 ;
        RECT 9.2840 51.5440 9.3020 52.7030 ;
        RECT 7.8800 51.5840 7.9700 52.6980 ;
        RECT 7.2320 51.5440 7.2500 52.7030 ;
        RECT 0.1220 51.5435 0.1400 52.7035 ;
        RECT 16.3940 52.6235 16.4120 53.7835 ;
        RECT 9.2840 52.6240 9.3020 53.7830 ;
        RECT 7.8800 52.6640 7.9700 53.7780 ;
        RECT 7.2320 52.6240 7.2500 53.7830 ;
        RECT 0.1220 52.6235 0.1400 53.7835 ;
        RECT 16.3940 53.7035 16.4120 54.8635 ;
        RECT 9.2840 53.7040 9.3020 54.8630 ;
        RECT 7.8800 53.7440 7.9700 54.8580 ;
        RECT 7.2320 53.7040 7.2500 54.8630 ;
        RECT 0.1220 53.7035 0.1400 54.8635 ;
        RECT 16.3940 54.7835 16.4120 55.9435 ;
        RECT 9.2840 54.7840 9.3020 55.9430 ;
        RECT 7.8800 54.8240 7.9700 55.9380 ;
        RECT 7.2320 54.7840 7.2500 55.9430 ;
        RECT 0.1220 54.7835 0.1400 55.9435 ;
        RECT 16.3940 55.8635 16.4120 57.0235 ;
        RECT 9.2840 55.8640 9.3020 57.0230 ;
        RECT 7.8800 55.9040 7.9700 57.0180 ;
        RECT 7.2320 55.8640 7.2500 57.0230 ;
        RECT 0.1220 55.8635 0.1400 57.0235 ;
        RECT 16.3940 56.9435 16.4120 58.1035 ;
        RECT 9.2840 56.9440 9.3020 58.1030 ;
        RECT 7.8800 56.9840 7.9700 58.0980 ;
        RECT 7.2320 56.9440 7.2500 58.1030 ;
        RECT 0.1220 56.9435 0.1400 58.1035 ;
        RECT 16.3940 58.0235 16.4120 59.1835 ;
        RECT 9.2840 58.0240 9.3020 59.1830 ;
        RECT 7.8800 58.0640 7.9700 59.1780 ;
        RECT 7.2320 58.0240 7.2500 59.1830 ;
        RECT 0.1220 58.0235 0.1400 59.1835 ;
        RECT 16.3940 59.1035 16.4120 60.2635 ;
        RECT 9.2840 59.1040 9.3020 60.2630 ;
        RECT 7.8800 59.1440 7.9700 60.2580 ;
        RECT 7.2320 59.1040 7.2500 60.2630 ;
        RECT 0.1220 59.1035 0.1400 60.2635 ;
        RECT 16.3940 60.1835 16.4120 61.3435 ;
        RECT 9.2840 60.1840 9.3020 61.3430 ;
        RECT 7.8800 60.2240 7.9700 61.3380 ;
        RECT 7.2320 60.1840 7.2500 61.3430 ;
        RECT 0.1220 60.1835 0.1400 61.3435 ;
        RECT 16.3940 61.2635 16.4120 62.4235 ;
        RECT 9.2840 61.2640 9.3020 62.4230 ;
        RECT 7.8800 61.3040 7.9700 62.4180 ;
        RECT 7.2320 61.2640 7.2500 62.4230 ;
        RECT 0.1220 61.2635 0.1400 62.4235 ;
        RECT 16.3940 62.3435 16.4120 63.5035 ;
        RECT 9.2840 62.3440 9.3020 63.5030 ;
        RECT 7.8800 62.3840 7.9700 63.4980 ;
        RECT 7.2320 62.3440 7.2500 63.5030 ;
        RECT 0.1220 62.3435 0.1400 63.5035 ;
        RECT 16.3940 63.4235 16.4120 64.5835 ;
        RECT 9.2840 63.4240 9.3020 64.5830 ;
        RECT 7.8800 63.4640 7.9700 64.5780 ;
        RECT 7.2320 63.4240 7.2500 64.5830 ;
        RECT 0.1220 63.4235 0.1400 64.5835 ;
        RECT 16.3940 64.5035 16.4120 65.6635 ;
        RECT 9.2840 64.5040 9.3020 65.6630 ;
        RECT 7.8800 64.5440 7.9700 65.6580 ;
        RECT 7.2320 64.5040 7.2500 65.6630 ;
        RECT 0.1220 64.5035 0.1400 65.6635 ;
        RECT 16.3940 65.5835 16.4120 66.7435 ;
        RECT 9.2840 65.5840 9.3020 66.7430 ;
        RECT 7.8800 65.6240 7.9700 66.7380 ;
        RECT 7.2320 65.5840 7.2500 66.7430 ;
        RECT 0.1220 65.5835 0.1400 66.7435 ;
        RECT 16.3940 66.6635 16.4120 67.8235 ;
        RECT 9.2840 66.6640 9.3020 67.8230 ;
        RECT 7.8800 66.7040 7.9700 67.8180 ;
        RECT 7.2320 66.6640 7.2500 67.8230 ;
        RECT 0.1220 66.6635 0.1400 67.8235 ;
        RECT 16.3940 67.7435 16.4120 68.9035 ;
        RECT 9.2840 67.7440 9.3020 68.9030 ;
        RECT 7.8800 67.7840 7.9700 68.8980 ;
        RECT 7.2320 67.7440 7.2500 68.9030 ;
        RECT 0.1220 67.7435 0.1400 68.9035 ;
        RECT 16.3940 68.8235 16.4120 69.9835 ;
        RECT 9.2840 68.8240 9.3020 69.9830 ;
        RECT 7.8800 68.8640 7.9700 69.9780 ;
        RECT 7.2320 68.8240 7.2500 69.9830 ;
        RECT 0.1220 68.8235 0.1400 69.9835 ;
        RECT 16.3940 69.9035 16.4120 71.0635 ;
        RECT 9.2840 69.9040 9.3020 71.0630 ;
        RECT 7.8800 69.9440 7.9700 71.0580 ;
        RECT 7.2320 69.9040 7.2500 71.0630 ;
        RECT 0.1220 69.9035 0.1400 71.0635 ;
        RECT 16.3940 70.9835 16.4120 72.1435 ;
        RECT 9.2840 70.9840 9.3020 72.1430 ;
        RECT 7.8800 71.0240 7.9700 72.1380 ;
        RECT 7.2320 70.9840 7.2500 72.1430 ;
        RECT 0.1220 70.9835 0.1400 72.1435 ;
        RECT 16.3940 72.0635 16.4120 73.2235 ;
        RECT 9.2840 72.0640 9.3020 73.2230 ;
        RECT 7.8800 72.1040 7.9700 73.2180 ;
        RECT 7.2320 72.0640 7.2500 73.2230 ;
        RECT 0.1220 72.0635 0.1400 73.2235 ;
        RECT 16.3940 73.1435 16.4120 74.3035 ;
        RECT 9.2840 73.1440 9.3020 74.3030 ;
        RECT 7.8800 73.1840 7.9700 74.2980 ;
        RECT 7.2320 73.1440 7.2500 74.3030 ;
        RECT 0.1220 73.1435 0.1400 74.3035 ;
        RECT 16.3940 74.2235 16.4120 75.3835 ;
        RECT 9.2840 74.2240 9.3020 75.3830 ;
        RECT 7.8800 74.2640 7.9700 75.3780 ;
        RECT 7.2320 74.2240 7.2500 75.3830 ;
        RECT 0.1220 74.2235 0.1400 75.3835 ;
        RECT 16.3940 75.3035 16.4120 76.4635 ;
        RECT 9.2840 75.3040 9.3020 76.4630 ;
        RECT 7.8800 75.3440 7.9700 76.4580 ;
        RECT 7.2320 75.3040 7.2500 76.4630 ;
        RECT 0.1220 75.3035 0.1400 76.4635 ;
        RECT 16.3940 76.3835 16.4120 77.5435 ;
        RECT 9.2840 76.3840 9.3020 77.5430 ;
        RECT 7.8800 76.4240 7.9700 77.5380 ;
        RECT 7.2320 76.3840 7.2500 77.5430 ;
        RECT 0.1220 76.3835 0.1400 77.5435 ;
        RECT 16.3940 77.4635 16.4120 78.6235 ;
        RECT 9.2840 77.4640 9.3020 78.6230 ;
        RECT 7.8800 77.5040 7.9700 78.6180 ;
        RECT 7.2320 77.4640 7.2500 78.6230 ;
        RECT 0.1220 77.4635 0.1400 78.6235 ;
        RECT 16.3940 78.5435 16.4120 79.7035 ;
        RECT 9.2840 78.5440 9.3020 79.7030 ;
        RECT 7.8800 78.5840 7.9700 79.6980 ;
        RECT 7.2320 78.5440 7.2500 79.7030 ;
        RECT 0.1220 78.5435 0.1400 79.7035 ;
        RECT 16.3940 79.6235 16.4120 80.7835 ;
        RECT 9.2840 79.6240 9.3020 80.7830 ;
        RECT 7.8800 79.6640 7.9700 80.7780 ;
        RECT 7.2320 79.6240 7.2500 80.7830 ;
        RECT 0.1220 79.6235 0.1400 80.7835 ;
        RECT 16.3940 80.7035 16.4120 81.8635 ;
        RECT 9.2840 80.7040 9.3020 81.8630 ;
        RECT 7.8800 80.7440 7.9700 81.8580 ;
        RECT 7.2320 80.7040 7.2500 81.8630 ;
        RECT 0.1220 80.7035 0.1400 81.8635 ;
        RECT 16.3940 81.7835 16.4120 82.9435 ;
        RECT 9.2840 81.7840 9.3020 82.9430 ;
        RECT 7.8800 81.8240 7.9700 82.9380 ;
        RECT 7.2320 81.7840 7.2500 82.9430 ;
        RECT 0.1220 81.7835 0.1400 82.9435 ;
        RECT 16.3940 82.8635 16.4120 84.0235 ;
        RECT 9.2840 82.8640 9.3020 84.0230 ;
        RECT 7.8800 82.9040 7.9700 84.0180 ;
        RECT 7.2320 82.8640 7.2500 84.0230 ;
        RECT 0.1220 82.8635 0.1400 84.0235 ;
        RECT 16.3940 83.9435 16.4120 85.1035 ;
        RECT 9.2840 83.9440 9.3020 85.1030 ;
        RECT 7.8800 83.9840 7.9700 85.0980 ;
        RECT 7.2320 83.9440 7.2500 85.1030 ;
        RECT 0.1220 83.9435 0.1400 85.1035 ;
        RECT 16.3940 85.0235 16.4120 86.1835 ;
        RECT 9.2840 85.0240 9.3020 86.1830 ;
        RECT 7.8800 85.0640 7.9700 86.1780 ;
        RECT 7.2320 85.0240 7.2500 86.1830 ;
        RECT 0.1220 85.0235 0.1400 86.1835 ;
        RECT 16.3940 86.1035 16.4120 87.2635 ;
        RECT 9.2840 86.1040 9.3020 87.2630 ;
        RECT 7.8800 86.1440 7.9700 87.2580 ;
        RECT 7.2320 86.1040 7.2500 87.2630 ;
        RECT 0.1220 86.1035 0.1400 87.2635 ;
        RECT 16.3940 87.1835 16.4120 88.3435 ;
        RECT 9.2840 87.1840 9.3020 88.3430 ;
        RECT 7.8800 87.2240 7.9700 88.3380 ;
        RECT 7.2320 87.1840 7.2500 88.3430 ;
        RECT 0.1220 87.1835 0.1400 88.3435 ;
      LAYER V3  ;
        RECT 0.1220 1.1720 0.1400 1.2200 ;
        RECT 7.2320 1.1720 7.2500 1.2200 ;
        RECT 7.8800 1.1720 7.9700 1.2200 ;
        RECT 9.2840 1.1720 9.3020 1.2200 ;
        RECT 16.3940 1.1720 16.4120 1.2200 ;
        RECT 0.1220 2.2520 0.1400 2.3000 ;
        RECT 7.2320 2.2520 7.2500 2.3000 ;
        RECT 7.8800 2.2520 7.9700 2.3000 ;
        RECT 9.2840 2.2520 9.3020 2.3000 ;
        RECT 16.3940 2.2520 16.4120 2.3000 ;
        RECT 0.1220 3.3320 0.1400 3.3800 ;
        RECT 7.2320 3.3320 7.2500 3.3800 ;
        RECT 7.8800 3.3320 7.9700 3.3800 ;
        RECT 9.2840 3.3320 9.3020 3.3800 ;
        RECT 16.3940 3.3320 16.4120 3.3800 ;
        RECT 0.1220 4.4120 0.1400 4.4600 ;
        RECT 7.2320 4.4120 7.2500 4.4600 ;
        RECT 7.8800 4.4120 7.9700 4.4600 ;
        RECT 9.2840 4.4120 9.3020 4.4600 ;
        RECT 16.3940 4.4120 16.4120 4.4600 ;
        RECT 0.1220 5.4920 0.1400 5.5400 ;
        RECT 7.2320 5.4920 7.2500 5.5400 ;
        RECT 7.8800 5.4920 7.9700 5.5400 ;
        RECT 9.2840 5.4920 9.3020 5.5400 ;
        RECT 16.3940 5.4920 16.4120 5.5400 ;
        RECT 0.1220 6.5720 0.1400 6.6200 ;
        RECT 7.2320 6.5720 7.2500 6.6200 ;
        RECT 7.8800 6.5720 7.9700 6.6200 ;
        RECT 9.2840 6.5720 9.3020 6.6200 ;
        RECT 16.3940 6.5720 16.4120 6.6200 ;
        RECT 0.1220 7.6520 0.1400 7.7000 ;
        RECT 7.2320 7.6520 7.2500 7.7000 ;
        RECT 7.8800 7.6520 7.9700 7.7000 ;
        RECT 9.2840 7.6520 9.3020 7.7000 ;
        RECT 16.3940 7.6520 16.4120 7.7000 ;
        RECT 0.1220 8.7320 0.1400 8.7800 ;
        RECT 7.2320 8.7320 7.2500 8.7800 ;
        RECT 7.8800 8.7320 7.9700 8.7800 ;
        RECT 9.2840 8.7320 9.3020 8.7800 ;
        RECT 16.3940 8.7320 16.4120 8.7800 ;
        RECT 0.1220 9.8120 0.1400 9.8600 ;
        RECT 7.2320 9.8120 7.2500 9.8600 ;
        RECT 7.8800 9.8120 7.9700 9.8600 ;
        RECT 9.2840 9.8120 9.3020 9.8600 ;
        RECT 16.3940 9.8120 16.4120 9.8600 ;
        RECT 0.1220 10.8920 0.1400 10.9400 ;
        RECT 7.2320 10.8920 7.2500 10.9400 ;
        RECT 7.8800 10.8920 7.9700 10.9400 ;
        RECT 9.2840 10.8920 9.3020 10.9400 ;
        RECT 16.3940 10.8920 16.4120 10.9400 ;
        RECT 0.1220 11.9720 0.1400 12.0200 ;
        RECT 7.2320 11.9720 7.2500 12.0200 ;
        RECT 7.8800 11.9720 7.9700 12.0200 ;
        RECT 9.2840 11.9720 9.3020 12.0200 ;
        RECT 16.3940 11.9720 16.4120 12.0200 ;
        RECT 0.1220 13.0520 0.1400 13.1000 ;
        RECT 7.2320 13.0520 7.2500 13.1000 ;
        RECT 7.8800 13.0520 7.9700 13.1000 ;
        RECT 9.2840 13.0520 9.3020 13.1000 ;
        RECT 16.3940 13.0520 16.4120 13.1000 ;
        RECT 0.1220 14.1320 0.1400 14.1800 ;
        RECT 7.2320 14.1320 7.2500 14.1800 ;
        RECT 7.8800 14.1320 7.9700 14.1800 ;
        RECT 9.2840 14.1320 9.3020 14.1800 ;
        RECT 16.3940 14.1320 16.4120 14.1800 ;
        RECT 0.1220 15.2120 0.1400 15.2600 ;
        RECT 7.2320 15.2120 7.2500 15.2600 ;
        RECT 7.8800 15.2120 7.9700 15.2600 ;
        RECT 9.2840 15.2120 9.3020 15.2600 ;
        RECT 16.3940 15.2120 16.4120 15.2600 ;
        RECT 0.1220 16.2920 0.1400 16.3400 ;
        RECT 7.2320 16.2920 7.2500 16.3400 ;
        RECT 7.8800 16.2920 7.9700 16.3400 ;
        RECT 9.2840 16.2920 9.3020 16.3400 ;
        RECT 16.3940 16.2920 16.4120 16.3400 ;
        RECT 0.1220 17.3720 0.1400 17.4200 ;
        RECT 7.2320 17.3720 7.2500 17.4200 ;
        RECT 7.8800 17.3720 7.9700 17.4200 ;
        RECT 9.2840 17.3720 9.3020 17.4200 ;
        RECT 16.3940 17.3720 16.4120 17.4200 ;
        RECT 0.1220 18.4520 0.1400 18.5000 ;
        RECT 7.2320 18.4520 7.2500 18.5000 ;
        RECT 7.8800 18.4520 7.9700 18.5000 ;
        RECT 9.2840 18.4520 9.3020 18.5000 ;
        RECT 16.3940 18.4520 16.4120 18.5000 ;
        RECT 0.1220 19.5320 0.1400 19.5800 ;
        RECT 7.2320 19.5320 7.2500 19.5800 ;
        RECT 7.8800 19.5320 7.9700 19.5800 ;
        RECT 9.2840 19.5320 9.3020 19.5800 ;
        RECT 16.3940 19.5320 16.4120 19.5800 ;
        RECT 0.1220 20.6120 0.1400 20.6600 ;
        RECT 7.2320 20.6120 7.2500 20.6600 ;
        RECT 7.8800 20.6120 7.9700 20.6600 ;
        RECT 9.2840 20.6120 9.3020 20.6600 ;
        RECT 16.3940 20.6120 16.4120 20.6600 ;
        RECT 0.1220 21.6920 0.1400 21.7400 ;
        RECT 7.2320 21.6920 7.2500 21.7400 ;
        RECT 7.8800 21.6920 7.9700 21.7400 ;
        RECT 9.2840 21.6920 9.3020 21.7400 ;
        RECT 16.3940 21.6920 16.4120 21.7400 ;
        RECT 0.1220 22.7720 0.1400 22.8200 ;
        RECT 7.2320 22.7720 7.2500 22.8200 ;
        RECT 7.8800 22.7720 7.9700 22.8200 ;
        RECT 9.2840 22.7720 9.3020 22.8200 ;
        RECT 16.3940 22.7720 16.4120 22.8200 ;
        RECT 0.1220 23.8520 0.1400 23.9000 ;
        RECT 7.2320 23.8520 7.2500 23.9000 ;
        RECT 7.8800 23.8520 7.9700 23.9000 ;
        RECT 9.2840 23.8520 9.3020 23.9000 ;
        RECT 16.3940 23.8520 16.4120 23.9000 ;
        RECT 0.1220 24.9320 0.1400 24.9800 ;
        RECT 7.2320 24.9320 7.2500 24.9800 ;
        RECT 7.8800 24.9320 7.9700 24.9800 ;
        RECT 9.2840 24.9320 9.3020 24.9800 ;
        RECT 16.3940 24.9320 16.4120 24.9800 ;
        RECT 0.1220 26.0120 0.1400 26.0600 ;
        RECT 7.2320 26.0120 7.2500 26.0600 ;
        RECT 7.8800 26.0120 7.9700 26.0600 ;
        RECT 9.2840 26.0120 9.3020 26.0600 ;
        RECT 16.3940 26.0120 16.4120 26.0600 ;
        RECT 0.1220 27.0920 0.1400 27.1400 ;
        RECT 7.2320 27.0920 7.2500 27.1400 ;
        RECT 7.8800 27.0920 7.9700 27.1400 ;
        RECT 9.2840 27.0920 9.3020 27.1400 ;
        RECT 16.3940 27.0920 16.4120 27.1400 ;
        RECT 0.1220 28.1720 0.1400 28.2200 ;
        RECT 7.2320 28.1720 7.2500 28.2200 ;
        RECT 7.8800 28.1720 7.9700 28.2200 ;
        RECT 9.2840 28.1720 9.3020 28.2200 ;
        RECT 16.3940 28.1720 16.4120 28.2200 ;
        RECT 0.1220 29.2520 0.1400 29.3000 ;
        RECT 7.2320 29.2520 7.2500 29.3000 ;
        RECT 7.8800 29.2520 7.9700 29.3000 ;
        RECT 9.2840 29.2520 9.3020 29.3000 ;
        RECT 16.3940 29.2520 16.4120 29.3000 ;
        RECT 0.1220 30.3320 0.1400 30.3800 ;
        RECT 7.2320 30.3320 7.2500 30.3800 ;
        RECT 7.8800 30.3320 7.9700 30.3800 ;
        RECT 9.2840 30.3320 9.3020 30.3800 ;
        RECT 16.3940 30.3320 16.4120 30.3800 ;
        RECT 0.1220 31.4120 0.1400 31.4600 ;
        RECT 7.2320 31.4120 7.2500 31.4600 ;
        RECT 7.8800 31.4120 7.9700 31.4600 ;
        RECT 9.2840 31.4120 9.3020 31.4600 ;
        RECT 16.3940 31.4120 16.4120 31.4600 ;
        RECT 0.1220 32.4920 0.1400 32.5400 ;
        RECT 7.2320 32.4920 7.2500 32.5400 ;
        RECT 7.8800 32.4920 7.9700 32.5400 ;
        RECT 9.2840 32.4920 9.3020 32.5400 ;
        RECT 16.3940 32.4920 16.4120 32.5400 ;
        RECT 0.1220 33.5720 0.1400 33.6200 ;
        RECT 7.2320 33.5720 7.2500 33.6200 ;
        RECT 7.8800 33.5720 7.9700 33.6200 ;
        RECT 9.2840 33.5720 9.3020 33.6200 ;
        RECT 16.3940 33.5720 16.4120 33.6200 ;
        RECT 0.1220 34.6520 0.1400 34.7000 ;
        RECT 7.2320 34.6520 7.2500 34.7000 ;
        RECT 7.8800 34.6520 7.9700 34.7000 ;
        RECT 9.2840 34.6520 9.3020 34.7000 ;
        RECT 16.3940 34.6520 16.4120 34.7000 ;
        RECT 0.1220 35.7320 0.1400 35.7800 ;
        RECT 7.2320 35.7320 7.2500 35.7800 ;
        RECT 7.8800 35.7320 7.9700 35.7800 ;
        RECT 9.2840 35.7320 9.3020 35.7800 ;
        RECT 16.3940 35.7320 16.4120 35.7800 ;
        RECT 0.1220 36.8120 0.1400 36.8600 ;
        RECT 7.2320 36.8120 7.2500 36.8600 ;
        RECT 7.8800 36.8120 7.9700 36.8600 ;
        RECT 9.2840 36.8120 9.3020 36.8600 ;
        RECT 16.3940 36.8120 16.4120 36.8600 ;
        RECT 0.1220 37.8920 0.1400 37.9400 ;
        RECT 7.2320 37.8920 7.2500 37.9400 ;
        RECT 7.8800 37.8920 7.9700 37.9400 ;
        RECT 9.2840 37.8920 9.3020 37.9400 ;
        RECT 16.3940 37.8920 16.4120 37.9400 ;
        RECT 0.1220 38.9720 0.1400 39.0200 ;
        RECT 7.2320 38.9720 7.2500 39.0200 ;
        RECT 7.8800 38.9720 7.9700 39.0200 ;
        RECT 9.2840 38.9720 9.3020 39.0200 ;
        RECT 16.3940 38.9720 16.4120 39.0200 ;
        RECT 0.1220 40.0520 0.1400 40.1000 ;
        RECT 7.2320 40.0520 7.2500 40.1000 ;
        RECT 7.8800 40.0520 7.9700 40.1000 ;
        RECT 9.2840 40.0520 9.3020 40.1000 ;
        RECT 16.3940 40.0520 16.4120 40.1000 ;
        RECT 7.9150 46.8690 7.9330 47.0850 ;
        RECT 7.9150 43.7010 7.9330 43.9170 ;
        RECT 7.9150 40.5330 7.9330 40.7490 ;
        RECT 7.9670 46.8690 7.9850 47.0850 ;
        RECT 7.9670 43.7010 7.9850 43.9170 ;
        RECT 7.9670 40.5330 7.9850 40.7490 ;
        RECT 8.0190 46.8690 8.0370 47.0850 ;
        RECT 8.0190 43.7010 8.0370 43.9170 ;
        RECT 8.0190 40.5330 8.0370 40.7490 ;
        RECT 8.0710 46.8690 8.0890 47.0850 ;
        RECT 8.0710 43.7010 8.0890 43.9170 ;
        RECT 8.0710 40.5330 8.0890 40.7490 ;
        RECT 8.1230 46.8690 8.1410 47.0850 ;
        RECT 8.1230 43.7010 8.1410 43.9170 ;
        RECT 8.1230 40.5330 8.1410 40.7490 ;
        RECT 9.2790 40.2530 9.2970 40.2770 ;
        RECT 9.2970 44.0370 9.3150 44.0610 ;
        RECT 0.1220 49.2590 0.1400 49.3070 ;
        RECT 7.2320 49.2590 7.2500 49.3070 ;
        RECT 7.8800 49.2590 7.9700 49.3070 ;
        RECT 9.2840 49.2590 9.3020 49.3070 ;
        RECT 16.3940 49.2590 16.4120 49.3070 ;
        RECT 0.1220 50.3390 0.1400 50.3870 ;
        RECT 7.2320 50.3390 7.2500 50.3870 ;
        RECT 7.8800 50.3390 7.9700 50.3870 ;
        RECT 9.2840 50.3390 9.3020 50.3870 ;
        RECT 16.3940 50.3390 16.4120 50.3870 ;
        RECT 0.1220 51.4190 0.1400 51.4670 ;
        RECT 7.2320 51.4190 7.2500 51.4670 ;
        RECT 7.8800 51.4190 7.9700 51.4670 ;
        RECT 9.2840 51.4190 9.3020 51.4670 ;
        RECT 16.3940 51.4190 16.4120 51.4670 ;
        RECT 0.1220 52.4990 0.1400 52.5470 ;
        RECT 7.2320 52.4990 7.2500 52.5470 ;
        RECT 7.8800 52.4990 7.9700 52.5470 ;
        RECT 9.2840 52.4990 9.3020 52.5470 ;
        RECT 16.3940 52.4990 16.4120 52.5470 ;
        RECT 0.1220 53.5790 0.1400 53.6270 ;
        RECT 7.2320 53.5790 7.2500 53.6270 ;
        RECT 7.8800 53.5790 7.9700 53.6270 ;
        RECT 9.2840 53.5790 9.3020 53.6270 ;
        RECT 16.3940 53.5790 16.4120 53.6270 ;
        RECT 0.1220 54.6590 0.1400 54.7070 ;
        RECT 7.2320 54.6590 7.2500 54.7070 ;
        RECT 7.8800 54.6590 7.9700 54.7070 ;
        RECT 9.2840 54.6590 9.3020 54.7070 ;
        RECT 16.3940 54.6590 16.4120 54.7070 ;
        RECT 0.1220 55.7390 0.1400 55.7870 ;
        RECT 7.2320 55.7390 7.2500 55.7870 ;
        RECT 7.8800 55.7390 7.9700 55.7870 ;
        RECT 9.2840 55.7390 9.3020 55.7870 ;
        RECT 16.3940 55.7390 16.4120 55.7870 ;
        RECT 0.1220 56.8190 0.1400 56.8670 ;
        RECT 7.2320 56.8190 7.2500 56.8670 ;
        RECT 7.8800 56.8190 7.9700 56.8670 ;
        RECT 9.2840 56.8190 9.3020 56.8670 ;
        RECT 16.3940 56.8190 16.4120 56.8670 ;
        RECT 0.1220 57.8990 0.1400 57.9470 ;
        RECT 7.2320 57.8990 7.2500 57.9470 ;
        RECT 7.8800 57.8990 7.9700 57.9470 ;
        RECT 9.2840 57.8990 9.3020 57.9470 ;
        RECT 16.3940 57.8990 16.4120 57.9470 ;
        RECT 0.1220 58.9790 0.1400 59.0270 ;
        RECT 7.2320 58.9790 7.2500 59.0270 ;
        RECT 7.8800 58.9790 7.9700 59.0270 ;
        RECT 9.2840 58.9790 9.3020 59.0270 ;
        RECT 16.3940 58.9790 16.4120 59.0270 ;
        RECT 0.1220 60.0590 0.1400 60.1070 ;
        RECT 7.2320 60.0590 7.2500 60.1070 ;
        RECT 7.8800 60.0590 7.9700 60.1070 ;
        RECT 9.2840 60.0590 9.3020 60.1070 ;
        RECT 16.3940 60.0590 16.4120 60.1070 ;
        RECT 0.1220 61.1390 0.1400 61.1870 ;
        RECT 7.2320 61.1390 7.2500 61.1870 ;
        RECT 7.8800 61.1390 7.9700 61.1870 ;
        RECT 9.2840 61.1390 9.3020 61.1870 ;
        RECT 16.3940 61.1390 16.4120 61.1870 ;
        RECT 0.1220 62.2190 0.1400 62.2670 ;
        RECT 7.2320 62.2190 7.2500 62.2670 ;
        RECT 7.8800 62.2190 7.9700 62.2670 ;
        RECT 9.2840 62.2190 9.3020 62.2670 ;
        RECT 16.3940 62.2190 16.4120 62.2670 ;
        RECT 0.1220 63.2990 0.1400 63.3470 ;
        RECT 7.2320 63.2990 7.2500 63.3470 ;
        RECT 7.8800 63.2990 7.9700 63.3470 ;
        RECT 9.2840 63.2990 9.3020 63.3470 ;
        RECT 16.3940 63.2990 16.4120 63.3470 ;
        RECT 0.1220 64.3790 0.1400 64.4270 ;
        RECT 7.2320 64.3790 7.2500 64.4270 ;
        RECT 7.8800 64.3790 7.9700 64.4270 ;
        RECT 9.2840 64.3790 9.3020 64.4270 ;
        RECT 16.3940 64.3790 16.4120 64.4270 ;
        RECT 0.1220 65.4590 0.1400 65.5070 ;
        RECT 7.2320 65.4590 7.2500 65.5070 ;
        RECT 7.8800 65.4590 7.9700 65.5070 ;
        RECT 9.2840 65.4590 9.3020 65.5070 ;
        RECT 16.3940 65.4590 16.4120 65.5070 ;
        RECT 0.1220 66.5390 0.1400 66.5870 ;
        RECT 7.2320 66.5390 7.2500 66.5870 ;
        RECT 7.8800 66.5390 7.9700 66.5870 ;
        RECT 9.2840 66.5390 9.3020 66.5870 ;
        RECT 16.3940 66.5390 16.4120 66.5870 ;
        RECT 0.1220 67.6190 0.1400 67.6670 ;
        RECT 7.2320 67.6190 7.2500 67.6670 ;
        RECT 7.8800 67.6190 7.9700 67.6670 ;
        RECT 9.2840 67.6190 9.3020 67.6670 ;
        RECT 16.3940 67.6190 16.4120 67.6670 ;
        RECT 0.1220 68.6990 0.1400 68.7470 ;
        RECT 7.2320 68.6990 7.2500 68.7470 ;
        RECT 7.8800 68.6990 7.9700 68.7470 ;
        RECT 9.2840 68.6990 9.3020 68.7470 ;
        RECT 16.3940 68.6990 16.4120 68.7470 ;
        RECT 0.1220 69.7790 0.1400 69.8270 ;
        RECT 7.2320 69.7790 7.2500 69.8270 ;
        RECT 7.8800 69.7790 7.9700 69.8270 ;
        RECT 9.2840 69.7790 9.3020 69.8270 ;
        RECT 16.3940 69.7790 16.4120 69.8270 ;
        RECT 0.1220 70.8590 0.1400 70.9070 ;
        RECT 7.2320 70.8590 7.2500 70.9070 ;
        RECT 7.8800 70.8590 7.9700 70.9070 ;
        RECT 9.2840 70.8590 9.3020 70.9070 ;
        RECT 16.3940 70.8590 16.4120 70.9070 ;
        RECT 0.1220 71.9390 0.1400 71.9870 ;
        RECT 7.2320 71.9390 7.2500 71.9870 ;
        RECT 7.8800 71.9390 7.9700 71.9870 ;
        RECT 9.2840 71.9390 9.3020 71.9870 ;
        RECT 16.3940 71.9390 16.4120 71.9870 ;
        RECT 0.1220 73.0190 0.1400 73.0670 ;
        RECT 7.2320 73.0190 7.2500 73.0670 ;
        RECT 7.8800 73.0190 7.9700 73.0670 ;
        RECT 9.2840 73.0190 9.3020 73.0670 ;
        RECT 16.3940 73.0190 16.4120 73.0670 ;
        RECT 0.1220 74.0990 0.1400 74.1470 ;
        RECT 7.2320 74.0990 7.2500 74.1470 ;
        RECT 7.8800 74.0990 7.9700 74.1470 ;
        RECT 9.2840 74.0990 9.3020 74.1470 ;
        RECT 16.3940 74.0990 16.4120 74.1470 ;
        RECT 0.1220 75.1790 0.1400 75.2270 ;
        RECT 7.2320 75.1790 7.2500 75.2270 ;
        RECT 7.8800 75.1790 7.9700 75.2270 ;
        RECT 9.2840 75.1790 9.3020 75.2270 ;
        RECT 16.3940 75.1790 16.4120 75.2270 ;
        RECT 0.1220 76.2590 0.1400 76.3070 ;
        RECT 7.2320 76.2590 7.2500 76.3070 ;
        RECT 7.8800 76.2590 7.9700 76.3070 ;
        RECT 9.2840 76.2590 9.3020 76.3070 ;
        RECT 16.3940 76.2590 16.4120 76.3070 ;
        RECT 0.1220 77.3390 0.1400 77.3870 ;
        RECT 7.2320 77.3390 7.2500 77.3870 ;
        RECT 7.8800 77.3390 7.9700 77.3870 ;
        RECT 9.2840 77.3390 9.3020 77.3870 ;
        RECT 16.3940 77.3390 16.4120 77.3870 ;
        RECT 0.1220 78.4190 0.1400 78.4670 ;
        RECT 7.2320 78.4190 7.2500 78.4670 ;
        RECT 7.8800 78.4190 7.9700 78.4670 ;
        RECT 9.2840 78.4190 9.3020 78.4670 ;
        RECT 16.3940 78.4190 16.4120 78.4670 ;
        RECT 0.1220 79.4990 0.1400 79.5470 ;
        RECT 7.2320 79.4990 7.2500 79.5470 ;
        RECT 7.8800 79.4990 7.9700 79.5470 ;
        RECT 9.2840 79.4990 9.3020 79.5470 ;
        RECT 16.3940 79.4990 16.4120 79.5470 ;
        RECT 0.1220 80.5790 0.1400 80.6270 ;
        RECT 7.2320 80.5790 7.2500 80.6270 ;
        RECT 7.8800 80.5790 7.9700 80.6270 ;
        RECT 9.2840 80.5790 9.3020 80.6270 ;
        RECT 16.3940 80.5790 16.4120 80.6270 ;
        RECT 0.1220 81.6590 0.1400 81.7070 ;
        RECT 7.2320 81.6590 7.2500 81.7070 ;
        RECT 7.8800 81.6590 7.9700 81.7070 ;
        RECT 9.2840 81.6590 9.3020 81.7070 ;
        RECT 16.3940 81.6590 16.4120 81.7070 ;
        RECT 0.1220 82.7390 0.1400 82.7870 ;
        RECT 7.2320 82.7390 7.2500 82.7870 ;
        RECT 7.8800 82.7390 7.9700 82.7870 ;
        RECT 9.2840 82.7390 9.3020 82.7870 ;
        RECT 16.3940 82.7390 16.4120 82.7870 ;
        RECT 0.1220 83.8190 0.1400 83.8670 ;
        RECT 7.2320 83.8190 7.2500 83.8670 ;
        RECT 7.8800 83.8190 7.9700 83.8670 ;
        RECT 9.2840 83.8190 9.3020 83.8670 ;
        RECT 16.3940 83.8190 16.4120 83.8670 ;
        RECT 0.1220 84.8990 0.1400 84.9470 ;
        RECT 7.2320 84.8990 7.2500 84.9470 ;
        RECT 7.8800 84.8990 7.9700 84.9470 ;
        RECT 9.2840 84.8990 9.3020 84.9470 ;
        RECT 16.3940 84.8990 16.4120 84.9470 ;
        RECT 0.1220 85.9790 0.1400 86.0270 ;
        RECT 7.2320 85.9790 7.2500 86.0270 ;
        RECT 7.8800 85.9790 7.9700 86.0270 ;
        RECT 9.2840 85.9790 9.3020 86.0270 ;
        RECT 16.3940 85.9790 16.4120 86.0270 ;
        RECT 0.1220 87.0590 0.1400 87.1070 ;
        RECT 7.2320 87.0590 7.2500 87.1070 ;
        RECT 7.8800 87.0590 7.9700 87.1070 ;
        RECT 9.2840 87.0590 9.3020 87.1070 ;
        RECT 16.3940 87.0590 16.4120 87.1070 ;
        RECT 0.1220 88.1390 0.1400 88.1870 ;
        RECT 7.2320 88.1390 7.2500 88.1870 ;
        RECT 7.8800 88.1390 7.9700 88.1870 ;
        RECT 9.2840 88.1390 9.3020 88.1870 ;
        RECT 16.3940 88.1390 16.4120 88.1870 ;
      LAYER M5  ;
        RECT 9.2160 40.2350 9.2400 44.0790 ;
      LAYER V4  ;
        RECT 9.2160 44.0370 9.2400 44.0610 ;
        RECT 9.2160 40.5330 9.2400 40.7490 ;
        RECT 9.2160 40.2530 9.2400 40.2770 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.0760 16.4370 1.1240 ;
        RECT 0.0940 2.1560 16.4370 2.2040 ;
        RECT 0.0940 3.2360 16.4370 3.2840 ;
        RECT 0.0940 4.3160 16.4370 4.3640 ;
        RECT 0.0940 5.3960 16.4370 5.4440 ;
        RECT 0.0940 6.4760 16.4370 6.5240 ;
        RECT 0.0940 7.5560 16.4370 7.6040 ;
        RECT 0.0940 8.6360 16.4370 8.6840 ;
        RECT 0.0940 9.7160 16.4370 9.7640 ;
        RECT 0.0940 10.7960 16.4370 10.8440 ;
        RECT 0.0940 11.8760 16.4370 11.9240 ;
        RECT 0.0940 12.9560 16.4370 13.0040 ;
        RECT 0.0940 14.0360 16.4370 14.0840 ;
        RECT 0.0940 15.1160 16.4370 15.1640 ;
        RECT 0.0940 16.1960 16.4370 16.2440 ;
        RECT 0.0940 17.2760 16.4370 17.3240 ;
        RECT 0.0940 18.3560 16.4370 18.4040 ;
        RECT 0.0940 19.4360 16.4370 19.4840 ;
        RECT 0.0940 20.5160 16.4370 20.5640 ;
        RECT 0.0940 21.5960 16.4370 21.6440 ;
        RECT 0.0940 22.6760 16.4370 22.7240 ;
        RECT 0.0940 23.7560 16.4370 23.8040 ;
        RECT 0.0940 24.8360 16.4370 24.8840 ;
        RECT 0.0940 25.9160 16.4370 25.9640 ;
        RECT 0.0940 26.9960 16.4370 27.0440 ;
        RECT 0.0940 28.0760 16.4370 28.1240 ;
        RECT 0.0940 29.1560 16.4370 29.2040 ;
        RECT 0.0940 30.2360 16.4370 30.2840 ;
        RECT 0.0940 31.3160 16.4370 31.3640 ;
        RECT 0.0940 32.3960 16.4370 32.4440 ;
        RECT 0.0940 33.4760 16.4370 33.5240 ;
        RECT 0.0940 34.5560 16.4370 34.6040 ;
        RECT 0.0940 35.6360 16.4370 35.6840 ;
        RECT 0.0940 36.7160 16.4370 36.7640 ;
        RECT 0.0940 37.7960 16.4370 37.8440 ;
        RECT 0.0940 38.8760 16.4370 38.9240 ;
        RECT 0.0940 39.9560 16.4370 40.0040 ;
        RECT 3.5640 40.9650 12.9600 41.1810 ;
        RECT 7.3980 44.1330 9.1260 44.3490 ;
        RECT 7.3980 47.3010 9.1260 47.5170 ;
        RECT 0.0940 49.1630 16.4370 49.2110 ;
        RECT 0.0940 50.2430 16.4370 50.2910 ;
        RECT 0.0940 51.3230 16.4370 51.3710 ;
        RECT 0.0940 52.4030 16.4370 52.4510 ;
        RECT 0.0940 53.4830 16.4370 53.5310 ;
        RECT 0.0940 54.5630 16.4370 54.6110 ;
        RECT 0.0940 55.6430 16.4370 55.6910 ;
        RECT 0.0940 56.7230 16.4370 56.7710 ;
        RECT 0.0940 57.8030 16.4370 57.8510 ;
        RECT 0.0940 58.8830 16.4370 58.9310 ;
        RECT 0.0940 59.9630 16.4370 60.0110 ;
        RECT 0.0940 61.0430 16.4370 61.0910 ;
        RECT 0.0940 62.1230 16.4370 62.1710 ;
        RECT 0.0940 63.2030 16.4370 63.2510 ;
        RECT 0.0940 64.2830 16.4370 64.3310 ;
        RECT 0.0940 65.3630 16.4370 65.4110 ;
        RECT 0.0940 66.4430 16.4370 66.4910 ;
        RECT 0.0940 67.5230 16.4370 67.5710 ;
        RECT 0.0940 68.6030 16.4370 68.6510 ;
        RECT 0.0940 69.6830 16.4370 69.7310 ;
        RECT 0.0940 70.7630 16.4370 70.8110 ;
        RECT 0.0940 71.8430 16.4370 71.8910 ;
        RECT 0.0940 72.9230 16.4370 72.9710 ;
        RECT 0.0940 74.0030 16.4370 74.0510 ;
        RECT 0.0940 75.0830 16.4370 75.1310 ;
        RECT 0.0940 76.1630 16.4370 76.2110 ;
        RECT 0.0940 77.2430 16.4370 77.2910 ;
        RECT 0.0940 78.3230 16.4370 78.3710 ;
        RECT 0.0940 79.4030 16.4370 79.4510 ;
        RECT 0.0940 80.4830 16.4370 80.5310 ;
        RECT 0.0940 81.5630 16.4370 81.6110 ;
        RECT 0.0940 82.6430 16.4370 82.6910 ;
        RECT 0.0940 83.7230 16.4370 83.7710 ;
        RECT 0.0940 84.8030 16.4370 84.8510 ;
        RECT 0.0940 85.8830 16.4370 85.9310 ;
        RECT 0.0940 86.9630 16.4370 87.0110 ;
        RECT 0.0940 88.0430 16.4370 88.0910 ;
      LAYER M3  ;
        RECT 16.3580 0.2165 16.3760 1.3765 ;
        RECT 9.3380 0.2165 9.3560 1.3765 ;
        RECT 8.5730 0.2530 8.6090 1.3670 ;
        RECT 8.4200 0.2530 8.4470 1.3670 ;
        RECT 7.1780 0.2165 7.1960 1.3765 ;
        RECT 0.1580 0.2165 0.1760 1.3765 ;
        RECT 16.3580 1.2965 16.3760 2.4565 ;
        RECT 9.3380 1.2965 9.3560 2.4565 ;
        RECT 8.5730 1.3330 8.6090 2.4470 ;
        RECT 8.4200 1.3330 8.4470 2.4470 ;
        RECT 7.1780 1.2965 7.1960 2.4565 ;
        RECT 0.1580 1.2965 0.1760 2.4565 ;
        RECT 16.3580 2.3765 16.3760 3.5365 ;
        RECT 9.3380 2.3765 9.3560 3.5365 ;
        RECT 8.5730 2.4130 8.6090 3.5270 ;
        RECT 8.4200 2.4130 8.4470 3.5270 ;
        RECT 7.1780 2.3765 7.1960 3.5365 ;
        RECT 0.1580 2.3765 0.1760 3.5365 ;
        RECT 16.3580 3.4565 16.3760 4.6165 ;
        RECT 9.3380 3.4565 9.3560 4.6165 ;
        RECT 8.5730 3.4930 8.6090 4.6070 ;
        RECT 8.4200 3.4930 8.4470 4.6070 ;
        RECT 7.1780 3.4565 7.1960 4.6165 ;
        RECT 0.1580 3.4565 0.1760 4.6165 ;
        RECT 16.3580 4.5365 16.3760 5.6965 ;
        RECT 9.3380 4.5365 9.3560 5.6965 ;
        RECT 8.5730 4.5730 8.6090 5.6870 ;
        RECT 8.4200 4.5730 8.4470 5.6870 ;
        RECT 7.1780 4.5365 7.1960 5.6965 ;
        RECT 0.1580 4.5365 0.1760 5.6965 ;
        RECT 16.3580 5.6165 16.3760 6.7765 ;
        RECT 9.3380 5.6165 9.3560 6.7765 ;
        RECT 8.5730 5.6530 8.6090 6.7670 ;
        RECT 8.4200 5.6530 8.4470 6.7670 ;
        RECT 7.1780 5.6165 7.1960 6.7765 ;
        RECT 0.1580 5.6165 0.1760 6.7765 ;
        RECT 16.3580 6.6965 16.3760 7.8565 ;
        RECT 9.3380 6.6965 9.3560 7.8565 ;
        RECT 8.5730 6.7330 8.6090 7.8470 ;
        RECT 8.4200 6.7330 8.4470 7.8470 ;
        RECT 7.1780 6.6965 7.1960 7.8565 ;
        RECT 0.1580 6.6965 0.1760 7.8565 ;
        RECT 16.3580 7.7765 16.3760 8.9365 ;
        RECT 9.3380 7.7765 9.3560 8.9365 ;
        RECT 8.5730 7.8130 8.6090 8.9270 ;
        RECT 8.4200 7.8130 8.4470 8.9270 ;
        RECT 7.1780 7.7765 7.1960 8.9365 ;
        RECT 0.1580 7.7765 0.1760 8.9365 ;
        RECT 16.3580 8.8565 16.3760 10.0165 ;
        RECT 9.3380 8.8565 9.3560 10.0165 ;
        RECT 8.5730 8.8930 8.6090 10.0070 ;
        RECT 8.4200 8.8930 8.4470 10.0070 ;
        RECT 7.1780 8.8565 7.1960 10.0165 ;
        RECT 0.1580 8.8565 0.1760 10.0165 ;
        RECT 16.3580 9.9365 16.3760 11.0965 ;
        RECT 9.3380 9.9365 9.3560 11.0965 ;
        RECT 8.5730 9.9730 8.6090 11.0870 ;
        RECT 8.4200 9.9730 8.4470 11.0870 ;
        RECT 7.1780 9.9365 7.1960 11.0965 ;
        RECT 0.1580 9.9365 0.1760 11.0965 ;
        RECT 16.3580 11.0165 16.3760 12.1765 ;
        RECT 9.3380 11.0165 9.3560 12.1765 ;
        RECT 8.5730 11.0530 8.6090 12.1670 ;
        RECT 8.4200 11.0530 8.4470 12.1670 ;
        RECT 7.1780 11.0165 7.1960 12.1765 ;
        RECT 0.1580 11.0165 0.1760 12.1765 ;
        RECT 16.3580 12.0965 16.3760 13.2565 ;
        RECT 9.3380 12.0965 9.3560 13.2565 ;
        RECT 8.5730 12.1330 8.6090 13.2470 ;
        RECT 8.4200 12.1330 8.4470 13.2470 ;
        RECT 7.1780 12.0965 7.1960 13.2565 ;
        RECT 0.1580 12.0965 0.1760 13.2565 ;
        RECT 16.3580 13.1765 16.3760 14.3365 ;
        RECT 9.3380 13.1765 9.3560 14.3365 ;
        RECT 8.5730 13.2130 8.6090 14.3270 ;
        RECT 8.4200 13.2130 8.4470 14.3270 ;
        RECT 7.1780 13.1765 7.1960 14.3365 ;
        RECT 0.1580 13.1765 0.1760 14.3365 ;
        RECT 16.3580 14.2565 16.3760 15.4165 ;
        RECT 9.3380 14.2565 9.3560 15.4165 ;
        RECT 8.5730 14.2930 8.6090 15.4070 ;
        RECT 8.4200 14.2930 8.4470 15.4070 ;
        RECT 7.1780 14.2565 7.1960 15.4165 ;
        RECT 0.1580 14.2565 0.1760 15.4165 ;
        RECT 16.3580 15.3365 16.3760 16.4965 ;
        RECT 9.3380 15.3365 9.3560 16.4965 ;
        RECT 8.5730 15.3730 8.6090 16.4870 ;
        RECT 8.4200 15.3730 8.4470 16.4870 ;
        RECT 7.1780 15.3365 7.1960 16.4965 ;
        RECT 0.1580 15.3365 0.1760 16.4965 ;
        RECT 16.3580 16.4165 16.3760 17.5765 ;
        RECT 9.3380 16.4165 9.3560 17.5765 ;
        RECT 8.5730 16.4530 8.6090 17.5670 ;
        RECT 8.4200 16.4530 8.4470 17.5670 ;
        RECT 7.1780 16.4165 7.1960 17.5765 ;
        RECT 0.1580 16.4165 0.1760 17.5765 ;
        RECT 16.3580 17.4965 16.3760 18.6565 ;
        RECT 9.3380 17.4965 9.3560 18.6565 ;
        RECT 8.5730 17.5330 8.6090 18.6470 ;
        RECT 8.4200 17.5330 8.4470 18.6470 ;
        RECT 7.1780 17.4965 7.1960 18.6565 ;
        RECT 0.1580 17.4965 0.1760 18.6565 ;
        RECT 16.3580 18.5765 16.3760 19.7365 ;
        RECT 9.3380 18.5765 9.3560 19.7365 ;
        RECT 8.5730 18.6130 8.6090 19.7270 ;
        RECT 8.4200 18.6130 8.4470 19.7270 ;
        RECT 7.1780 18.5765 7.1960 19.7365 ;
        RECT 0.1580 18.5765 0.1760 19.7365 ;
        RECT 16.3580 19.6565 16.3760 20.8165 ;
        RECT 9.3380 19.6565 9.3560 20.8165 ;
        RECT 8.5730 19.6930 8.6090 20.8070 ;
        RECT 8.4200 19.6930 8.4470 20.8070 ;
        RECT 7.1780 19.6565 7.1960 20.8165 ;
        RECT 0.1580 19.6565 0.1760 20.8165 ;
        RECT 16.3580 20.7365 16.3760 21.8965 ;
        RECT 9.3380 20.7365 9.3560 21.8965 ;
        RECT 8.5730 20.7730 8.6090 21.8870 ;
        RECT 8.4200 20.7730 8.4470 21.8870 ;
        RECT 7.1780 20.7365 7.1960 21.8965 ;
        RECT 0.1580 20.7365 0.1760 21.8965 ;
        RECT 16.3580 21.8165 16.3760 22.9765 ;
        RECT 9.3380 21.8165 9.3560 22.9765 ;
        RECT 8.5730 21.8530 8.6090 22.9670 ;
        RECT 8.4200 21.8530 8.4470 22.9670 ;
        RECT 7.1780 21.8165 7.1960 22.9765 ;
        RECT 0.1580 21.8165 0.1760 22.9765 ;
        RECT 16.3580 22.8965 16.3760 24.0565 ;
        RECT 9.3380 22.8965 9.3560 24.0565 ;
        RECT 8.5730 22.9330 8.6090 24.0470 ;
        RECT 8.4200 22.9330 8.4470 24.0470 ;
        RECT 7.1780 22.8965 7.1960 24.0565 ;
        RECT 0.1580 22.8965 0.1760 24.0565 ;
        RECT 16.3580 23.9765 16.3760 25.1365 ;
        RECT 9.3380 23.9765 9.3560 25.1365 ;
        RECT 8.5730 24.0130 8.6090 25.1270 ;
        RECT 8.4200 24.0130 8.4470 25.1270 ;
        RECT 7.1780 23.9765 7.1960 25.1365 ;
        RECT 0.1580 23.9765 0.1760 25.1365 ;
        RECT 16.3580 25.0565 16.3760 26.2165 ;
        RECT 9.3380 25.0565 9.3560 26.2165 ;
        RECT 8.5730 25.0930 8.6090 26.2070 ;
        RECT 8.4200 25.0930 8.4470 26.2070 ;
        RECT 7.1780 25.0565 7.1960 26.2165 ;
        RECT 0.1580 25.0565 0.1760 26.2165 ;
        RECT 16.3580 26.1365 16.3760 27.2965 ;
        RECT 9.3380 26.1365 9.3560 27.2965 ;
        RECT 8.5730 26.1730 8.6090 27.2870 ;
        RECT 8.4200 26.1730 8.4470 27.2870 ;
        RECT 7.1780 26.1365 7.1960 27.2965 ;
        RECT 0.1580 26.1365 0.1760 27.2965 ;
        RECT 16.3580 27.2165 16.3760 28.3765 ;
        RECT 9.3380 27.2165 9.3560 28.3765 ;
        RECT 8.5730 27.2530 8.6090 28.3670 ;
        RECT 8.4200 27.2530 8.4470 28.3670 ;
        RECT 7.1780 27.2165 7.1960 28.3765 ;
        RECT 0.1580 27.2165 0.1760 28.3765 ;
        RECT 16.3580 28.2965 16.3760 29.4565 ;
        RECT 9.3380 28.2965 9.3560 29.4565 ;
        RECT 8.5730 28.3330 8.6090 29.4470 ;
        RECT 8.4200 28.3330 8.4470 29.4470 ;
        RECT 7.1780 28.2965 7.1960 29.4565 ;
        RECT 0.1580 28.2965 0.1760 29.4565 ;
        RECT 16.3580 29.3765 16.3760 30.5365 ;
        RECT 9.3380 29.3765 9.3560 30.5365 ;
        RECT 8.5730 29.4130 8.6090 30.5270 ;
        RECT 8.4200 29.4130 8.4470 30.5270 ;
        RECT 7.1780 29.3765 7.1960 30.5365 ;
        RECT 0.1580 29.3765 0.1760 30.5365 ;
        RECT 16.3580 30.4565 16.3760 31.6165 ;
        RECT 9.3380 30.4565 9.3560 31.6165 ;
        RECT 8.5730 30.4930 8.6090 31.6070 ;
        RECT 8.4200 30.4930 8.4470 31.6070 ;
        RECT 7.1780 30.4565 7.1960 31.6165 ;
        RECT 0.1580 30.4565 0.1760 31.6165 ;
        RECT 16.3580 31.5365 16.3760 32.6965 ;
        RECT 9.3380 31.5365 9.3560 32.6965 ;
        RECT 8.5730 31.5730 8.6090 32.6870 ;
        RECT 8.4200 31.5730 8.4470 32.6870 ;
        RECT 7.1780 31.5365 7.1960 32.6965 ;
        RECT 0.1580 31.5365 0.1760 32.6965 ;
        RECT 16.3580 32.6165 16.3760 33.7765 ;
        RECT 9.3380 32.6165 9.3560 33.7765 ;
        RECT 8.5730 32.6530 8.6090 33.7670 ;
        RECT 8.4200 32.6530 8.4470 33.7670 ;
        RECT 7.1780 32.6165 7.1960 33.7765 ;
        RECT 0.1580 32.6165 0.1760 33.7765 ;
        RECT 16.3580 33.6965 16.3760 34.8565 ;
        RECT 9.3380 33.6965 9.3560 34.8565 ;
        RECT 8.5730 33.7330 8.6090 34.8470 ;
        RECT 8.4200 33.7330 8.4470 34.8470 ;
        RECT 7.1780 33.6965 7.1960 34.8565 ;
        RECT 0.1580 33.6965 0.1760 34.8565 ;
        RECT 16.3580 34.7765 16.3760 35.9365 ;
        RECT 9.3380 34.7765 9.3560 35.9365 ;
        RECT 8.5730 34.8130 8.6090 35.9270 ;
        RECT 8.4200 34.8130 8.4470 35.9270 ;
        RECT 7.1780 34.7765 7.1960 35.9365 ;
        RECT 0.1580 34.7765 0.1760 35.9365 ;
        RECT 16.3580 35.8565 16.3760 37.0165 ;
        RECT 9.3380 35.8565 9.3560 37.0165 ;
        RECT 8.5730 35.8930 8.6090 37.0070 ;
        RECT 8.4200 35.8930 8.4470 37.0070 ;
        RECT 7.1780 35.8565 7.1960 37.0165 ;
        RECT 0.1580 35.8565 0.1760 37.0165 ;
        RECT 16.3580 36.9365 16.3760 38.0965 ;
        RECT 9.3380 36.9365 9.3560 38.0965 ;
        RECT 8.5730 36.9730 8.6090 38.0870 ;
        RECT 8.4200 36.9730 8.4470 38.0870 ;
        RECT 7.1780 36.9365 7.1960 38.0965 ;
        RECT 0.1580 36.9365 0.1760 38.0965 ;
        RECT 16.3580 38.0165 16.3760 39.1765 ;
        RECT 9.3380 38.0165 9.3560 39.1765 ;
        RECT 8.5730 38.0530 8.6090 39.1670 ;
        RECT 8.4200 38.0530 8.4470 39.1670 ;
        RECT 7.1780 38.0165 7.1960 39.1765 ;
        RECT 0.1580 38.0165 0.1760 39.1765 ;
        RECT 16.3580 39.0965 16.3760 40.2565 ;
        RECT 9.3380 39.0965 9.3560 40.2565 ;
        RECT 8.5730 39.1330 8.6090 40.2470 ;
        RECT 8.4200 39.1330 8.4470 40.2470 ;
        RECT 7.1780 39.0965 7.1960 40.2565 ;
        RECT 0.1580 39.0965 0.1760 40.2565 ;
        RECT 16.3530 40.1705 16.3710 48.3775 ;
        RECT 9.3330 40.1705 9.3510 48.3775 ;
        RECT 8.3790 40.3940 8.6130 48.0770 ;
        RECT 8.5680 40.2145 8.6040 48.3340 ;
        RECT 8.4150 40.2140 8.4420 48.3340 ;
        RECT 7.1730 40.1705 7.1910 48.3775 ;
        RECT 0.1530 40.1705 0.1710 48.3775 ;
        RECT 16.3580 48.3035 16.3760 49.4635 ;
        RECT 9.3380 48.3035 9.3560 49.4635 ;
        RECT 8.5730 48.3400 8.6090 49.4540 ;
        RECT 8.4200 48.3400 8.4470 49.4540 ;
        RECT 7.1780 48.3035 7.1960 49.4635 ;
        RECT 0.1580 48.3035 0.1760 49.4635 ;
        RECT 16.3580 49.3835 16.3760 50.5435 ;
        RECT 9.3380 49.3835 9.3560 50.5435 ;
        RECT 8.5730 49.4200 8.6090 50.5340 ;
        RECT 8.4200 49.4200 8.4470 50.5340 ;
        RECT 7.1780 49.3835 7.1960 50.5435 ;
        RECT 0.1580 49.3835 0.1760 50.5435 ;
        RECT 16.3580 50.4635 16.3760 51.6235 ;
        RECT 9.3380 50.4635 9.3560 51.6235 ;
        RECT 8.5730 50.5000 8.6090 51.6140 ;
        RECT 8.4200 50.5000 8.4470 51.6140 ;
        RECT 7.1780 50.4635 7.1960 51.6235 ;
        RECT 0.1580 50.4635 0.1760 51.6235 ;
        RECT 16.3580 51.5435 16.3760 52.7035 ;
        RECT 9.3380 51.5435 9.3560 52.7035 ;
        RECT 8.5730 51.5800 8.6090 52.6940 ;
        RECT 8.4200 51.5800 8.4470 52.6940 ;
        RECT 7.1780 51.5435 7.1960 52.7035 ;
        RECT 0.1580 51.5435 0.1760 52.7035 ;
        RECT 16.3580 52.6235 16.3760 53.7835 ;
        RECT 9.3380 52.6235 9.3560 53.7835 ;
        RECT 8.5730 52.6600 8.6090 53.7740 ;
        RECT 8.4200 52.6600 8.4470 53.7740 ;
        RECT 7.1780 52.6235 7.1960 53.7835 ;
        RECT 0.1580 52.6235 0.1760 53.7835 ;
        RECT 16.3580 53.7035 16.3760 54.8635 ;
        RECT 9.3380 53.7035 9.3560 54.8635 ;
        RECT 8.5730 53.7400 8.6090 54.8540 ;
        RECT 8.4200 53.7400 8.4470 54.8540 ;
        RECT 7.1780 53.7035 7.1960 54.8635 ;
        RECT 0.1580 53.7035 0.1760 54.8635 ;
        RECT 16.3580 54.7835 16.3760 55.9435 ;
        RECT 9.3380 54.7835 9.3560 55.9435 ;
        RECT 8.5730 54.8200 8.6090 55.9340 ;
        RECT 8.4200 54.8200 8.4470 55.9340 ;
        RECT 7.1780 54.7835 7.1960 55.9435 ;
        RECT 0.1580 54.7835 0.1760 55.9435 ;
        RECT 16.3580 55.8635 16.3760 57.0235 ;
        RECT 9.3380 55.8635 9.3560 57.0235 ;
        RECT 8.5730 55.9000 8.6090 57.0140 ;
        RECT 8.4200 55.9000 8.4470 57.0140 ;
        RECT 7.1780 55.8635 7.1960 57.0235 ;
        RECT 0.1580 55.8635 0.1760 57.0235 ;
        RECT 16.3580 56.9435 16.3760 58.1035 ;
        RECT 9.3380 56.9435 9.3560 58.1035 ;
        RECT 8.5730 56.9800 8.6090 58.0940 ;
        RECT 8.4200 56.9800 8.4470 58.0940 ;
        RECT 7.1780 56.9435 7.1960 58.1035 ;
        RECT 0.1580 56.9435 0.1760 58.1035 ;
        RECT 16.3580 58.0235 16.3760 59.1835 ;
        RECT 9.3380 58.0235 9.3560 59.1835 ;
        RECT 8.5730 58.0600 8.6090 59.1740 ;
        RECT 8.4200 58.0600 8.4470 59.1740 ;
        RECT 7.1780 58.0235 7.1960 59.1835 ;
        RECT 0.1580 58.0235 0.1760 59.1835 ;
        RECT 16.3580 59.1035 16.3760 60.2635 ;
        RECT 9.3380 59.1035 9.3560 60.2635 ;
        RECT 8.5730 59.1400 8.6090 60.2540 ;
        RECT 8.4200 59.1400 8.4470 60.2540 ;
        RECT 7.1780 59.1035 7.1960 60.2635 ;
        RECT 0.1580 59.1035 0.1760 60.2635 ;
        RECT 16.3580 60.1835 16.3760 61.3435 ;
        RECT 9.3380 60.1835 9.3560 61.3435 ;
        RECT 8.5730 60.2200 8.6090 61.3340 ;
        RECT 8.4200 60.2200 8.4470 61.3340 ;
        RECT 7.1780 60.1835 7.1960 61.3435 ;
        RECT 0.1580 60.1835 0.1760 61.3435 ;
        RECT 16.3580 61.2635 16.3760 62.4235 ;
        RECT 9.3380 61.2635 9.3560 62.4235 ;
        RECT 8.5730 61.3000 8.6090 62.4140 ;
        RECT 8.4200 61.3000 8.4470 62.4140 ;
        RECT 7.1780 61.2635 7.1960 62.4235 ;
        RECT 0.1580 61.2635 0.1760 62.4235 ;
        RECT 16.3580 62.3435 16.3760 63.5035 ;
        RECT 9.3380 62.3435 9.3560 63.5035 ;
        RECT 8.5730 62.3800 8.6090 63.4940 ;
        RECT 8.4200 62.3800 8.4470 63.4940 ;
        RECT 7.1780 62.3435 7.1960 63.5035 ;
        RECT 0.1580 62.3435 0.1760 63.5035 ;
        RECT 16.3580 63.4235 16.3760 64.5835 ;
        RECT 9.3380 63.4235 9.3560 64.5835 ;
        RECT 8.5730 63.4600 8.6090 64.5740 ;
        RECT 8.4200 63.4600 8.4470 64.5740 ;
        RECT 7.1780 63.4235 7.1960 64.5835 ;
        RECT 0.1580 63.4235 0.1760 64.5835 ;
        RECT 16.3580 64.5035 16.3760 65.6635 ;
        RECT 9.3380 64.5035 9.3560 65.6635 ;
        RECT 8.5730 64.5400 8.6090 65.6540 ;
        RECT 8.4200 64.5400 8.4470 65.6540 ;
        RECT 7.1780 64.5035 7.1960 65.6635 ;
        RECT 0.1580 64.5035 0.1760 65.6635 ;
        RECT 16.3580 65.5835 16.3760 66.7435 ;
        RECT 9.3380 65.5835 9.3560 66.7435 ;
        RECT 8.5730 65.6200 8.6090 66.7340 ;
        RECT 8.4200 65.6200 8.4470 66.7340 ;
        RECT 7.1780 65.5835 7.1960 66.7435 ;
        RECT 0.1580 65.5835 0.1760 66.7435 ;
        RECT 16.3580 66.6635 16.3760 67.8235 ;
        RECT 9.3380 66.6635 9.3560 67.8235 ;
        RECT 8.5730 66.7000 8.6090 67.8140 ;
        RECT 8.4200 66.7000 8.4470 67.8140 ;
        RECT 7.1780 66.6635 7.1960 67.8235 ;
        RECT 0.1580 66.6635 0.1760 67.8235 ;
        RECT 16.3580 67.7435 16.3760 68.9035 ;
        RECT 9.3380 67.7435 9.3560 68.9035 ;
        RECT 8.5730 67.7800 8.6090 68.8940 ;
        RECT 8.4200 67.7800 8.4470 68.8940 ;
        RECT 7.1780 67.7435 7.1960 68.9035 ;
        RECT 0.1580 67.7435 0.1760 68.9035 ;
        RECT 16.3580 68.8235 16.3760 69.9835 ;
        RECT 9.3380 68.8235 9.3560 69.9835 ;
        RECT 8.5730 68.8600 8.6090 69.9740 ;
        RECT 8.4200 68.8600 8.4470 69.9740 ;
        RECT 7.1780 68.8235 7.1960 69.9835 ;
        RECT 0.1580 68.8235 0.1760 69.9835 ;
        RECT 16.3580 69.9035 16.3760 71.0635 ;
        RECT 9.3380 69.9035 9.3560 71.0635 ;
        RECT 8.5730 69.9400 8.6090 71.0540 ;
        RECT 8.4200 69.9400 8.4470 71.0540 ;
        RECT 7.1780 69.9035 7.1960 71.0635 ;
        RECT 0.1580 69.9035 0.1760 71.0635 ;
        RECT 16.3580 70.9835 16.3760 72.1435 ;
        RECT 9.3380 70.9835 9.3560 72.1435 ;
        RECT 8.5730 71.0200 8.6090 72.1340 ;
        RECT 8.4200 71.0200 8.4470 72.1340 ;
        RECT 7.1780 70.9835 7.1960 72.1435 ;
        RECT 0.1580 70.9835 0.1760 72.1435 ;
        RECT 16.3580 72.0635 16.3760 73.2235 ;
        RECT 9.3380 72.0635 9.3560 73.2235 ;
        RECT 8.5730 72.1000 8.6090 73.2140 ;
        RECT 8.4200 72.1000 8.4470 73.2140 ;
        RECT 7.1780 72.0635 7.1960 73.2235 ;
        RECT 0.1580 72.0635 0.1760 73.2235 ;
        RECT 16.3580 73.1435 16.3760 74.3035 ;
        RECT 9.3380 73.1435 9.3560 74.3035 ;
        RECT 8.5730 73.1800 8.6090 74.2940 ;
        RECT 8.4200 73.1800 8.4470 74.2940 ;
        RECT 7.1780 73.1435 7.1960 74.3035 ;
        RECT 0.1580 73.1435 0.1760 74.3035 ;
        RECT 16.3580 74.2235 16.3760 75.3835 ;
        RECT 9.3380 74.2235 9.3560 75.3835 ;
        RECT 8.5730 74.2600 8.6090 75.3740 ;
        RECT 8.4200 74.2600 8.4470 75.3740 ;
        RECT 7.1780 74.2235 7.1960 75.3835 ;
        RECT 0.1580 74.2235 0.1760 75.3835 ;
        RECT 16.3580 75.3035 16.3760 76.4635 ;
        RECT 9.3380 75.3035 9.3560 76.4635 ;
        RECT 8.5730 75.3400 8.6090 76.4540 ;
        RECT 8.4200 75.3400 8.4470 76.4540 ;
        RECT 7.1780 75.3035 7.1960 76.4635 ;
        RECT 0.1580 75.3035 0.1760 76.4635 ;
        RECT 16.3580 76.3835 16.3760 77.5435 ;
        RECT 9.3380 76.3835 9.3560 77.5435 ;
        RECT 8.5730 76.4200 8.6090 77.5340 ;
        RECT 8.4200 76.4200 8.4470 77.5340 ;
        RECT 7.1780 76.3835 7.1960 77.5435 ;
        RECT 0.1580 76.3835 0.1760 77.5435 ;
        RECT 16.3580 77.4635 16.3760 78.6235 ;
        RECT 9.3380 77.4635 9.3560 78.6235 ;
        RECT 8.5730 77.5000 8.6090 78.6140 ;
        RECT 8.4200 77.5000 8.4470 78.6140 ;
        RECT 7.1780 77.4635 7.1960 78.6235 ;
        RECT 0.1580 77.4635 0.1760 78.6235 ;
        RECT 16.3580 78.5435 16.3760 79.7035 ;
        RECT 9.3380 78.5435 9.3560 79.7035 ;
        RECT 8.5730 78.5800 8.6090 79.6940 ;
        RECT 8.4200 78.5800 8.4470 79.6940 ;
        RECT 7.1780 78.5435 7.1960 79.7035 ;
        RECT 0.1580 78.5435 0.1760 79.7035 ;
        RECT 16.3580 79.6235 16.3760 80.7835 ;
        RECT 9.3380 79.6235 9.3560 80.7835 ;
        RECT 8.5730 79.6600 8.6090 80.7740 ;
        RECT 8.4200 79.6600 8.4470 80.7740 ;
        RECT 7.1780 79.6235 7.1960 80.7835 ;
        RECT 0.1580 79.6235 0.1760 80.7835 ;
        RECT 16.3580 80.7035 16.3760 81.8635 ;
        RECT 9.3380 80.7035 9.3560 81.8635 ;
        RECT 8.5730 80.7400 8.6090 81.8540 ;
        RECT 8.4200 80.7400 8.4470 81.8540 ;
        RECT 7.1780 80.7035 7.1960 81.8635 ;
        RECT 0.1580 80.7035 0.1760 81.8635 ;
        RECT 16.3580 81.7835 16.3760 82.9435 ;
        RECT 9.3380 81.7835 9.3560 82.9435 ;
        RECT 8.5730 81.8200 8.6090 82.9340 ;
        RECT 8.4200 81.8200 8.4470 82.9340 ;
        RECT 7.1780 81.7835 7.1960 82.9435 ;
        RECT 0.1580 81.7835 0.1760 82.9435 ;
        RECT 16.3580 82.8635 16.3760 84.0235 ;
        RECT 9.3380 82.8635 9.3560 84.0235 ;
        RECT 8.5730 82.9000 8.6090 84.0140 ;
        RECT 8.4200 82.9000 8.4470 84.0140 ;
        RECT 7.1780 82.8635 7.1960 84.0235 ;
        RECT 0.1580 82.8635 0.1760 84.0235 ;
        RECT 16.3580 83.9435 16.3760 85.1035 ;
        RECT 9.3380 83.9435 9.3560 85.1035 ;
        RECT 8.5730 83.9800 8.6090 85.0940 ;
        RECT 8.4200 83.9800 8.4470 85.0940 ;
        RECT 7.1780 83.9435 7.1960 85.1035 ;
        RECT 0.1580 83.9435 0.1760 85.1035 ;
        RECT 16.3580 85.0235 16.3760 86.1835 ;
        RECT 9.3380 85.0235 9.3560 86.1835 ;
        RECT 8.5730 85.0600 8.6090 86.1740 ;
        RECT 8.4200 85.0600 8.4470 86.1740 ;
        RECT 7.1780 85.0235 7.1960 86.1835 ;
        RECT 0.1580 85.0235 0.1760 86.1835 ;
        RECT 16.3580 86.1035 16.3760 87.2635 ;
        RECT 9.3380 86.1035 9.3560 87.2635 ;
        RECT 8.5730 86.1400 8.6090 87.2540 ;
        RECT 8.4200 86.1400 8.4470 87.2540 ;
        RECT 7.1780 86.1035 7.1960 87.2635 ;
        RECT 0.1580 86.1035 0.1760 87.2635 ;
        RECT 16.3580 87.1835 16.3760 88.3435 ;
        RECT 9.3380 87.1835 9.3560 88.3435 ;
        RECT 8.5730 87.2200 8.6090 88.3340 ;
        RECT 8.4200 87.2200 8.4470 88.3340 ;
        RECT 7.1780 87.1835 7.1960 88.3435 ;
        RECT 0.1580 87.1835 0.1760 88.3435 ;
      LAYER V3  ;
        RECT 0.1580 1.0760 0.1760 1.1240 ;
        RECT 7.1780 1.0760 7.1960 1.1240 ;
        RECT 8.4200 1.0760 8.4470 1.1240 ;
        RECT 8.5730 1.0760 8.6090 1.1240 ;
        RECT 9.3380 1.0760 9.3560 1.1240 ;
        RECT 16.3580 1.0760 16.3760 1.1240 ;
        RECT 0.1580 2.1560 0.1760 2.2040 ;
        RECT 7.1780 2.1560 7.1960 2.2040 ;
        RECT 8.4200 2.1560 8.4470 2.2040 ;
        RECT 8.5730 2.1560 8.6090 2.2040 ;
        RECT 9.3380 2.1560 9.3560 2.2040 ;
        RECT 16.3580 2.1560 16.3760 2.2040 ;
        RECT 0.1580 3.2360 0.1760 3.2840 ;
        RECT 7.1780 3.2360 7.1960 3.2840 ;
        RECT 8.4200 3.2360 8.4470 3.2840 ;
        RECT 8.5730 3.2360 8.6090 3.2840 ;
        RECT 9.3380 3.2360 9.3560 3.2840 ;
        RECT 16.3580 3.2360 16.3760 3.2840 ;
        RECT 0.1580 4.3160 0.1760 4.3640 ;
        RECT 7.1780 4.3160 7.1960 4.3640 ;
        RECT 8.4200 4.3160 8.4470 4.3640 ;
        RECT 8.5730 4.3160 8.6090 4.3640 ;
        RECT 9.3380 4.3160 9.3560 4.3640 ;
        RECT 16.3580 4.3160 16.3760 4.3640 ;
        RECT 0.1580 5.3960 0.1760 5.4440 ;
        RECT 7.1780 5.3960 7.1960 5.4440 ;
        RECT 8.4200 5.3960 8.4470 5.4440 ;
        RECT 8.5730 5.3960 8.6090 5.4440 ;
        RECT 9.3380 5.3960 9.3560 5.4440 ;
        RECT 16.3580 5.3960 16.3760 5.4440 ;
        RECT 0.1580 6.4760 0.1760 6.5240 ;
        RECT 7.1780 6.4760 7.1960 6.5240 ;
        RECT 8.4200 6.4760 8.4470 6.5240 ;
        RECT 8.5730 6.4760 8.6090 6.5240 ;
        RECT 9.3380 6.4760 9.3560 6.5240 ;
        RECT 16.3580 6.4760 16.3760 6.5240 ;
        RECT 0.1580 7.5560 0.1760 7.6040 ;
        RECT 7.1780 7.5560 7.1960 7.6040 ;
        RECT 8.4200 7.5560 8.4470 7.6040 ;
        RECT 8.5730 7.5560 8.6090 7.6040 ;
        RECT 9.3380 7.5560 9.3560 7.6040 ;
        RECT 16.3580 7.5560 16.3760 7.6040 ;
        RECT 0.1580 8.6360 0.1760 8.6840 ;
        RECT 7.1780 8.6360 7.1960 8.6840 ;
        RECT 8.4200 8.6360 8.4470 8.6840 ;
        RECT 8.5730 8.6360 8.6090 8.6840 ;
        RECT 9.3380 8.6360 9.3560 8.6840 ;
        RECT 16.3580 8.6360 16.3760 8.6840 ;
        RECT 0.1580 9.7160 0.1760 9.7640 ;
        RECT 7.1780 9.7160 7.1960 9.7640 ;
        RECT 8.4200 9.7160 8.4470 9.7640 ;
        RECT 8.5730 9.7160 8.6090 9.7640 ;
        RECT 9.3380 9.7160 9.3560 9.7640 ;
        RECT 16.3580 9.7160 16.3760 9.7640 ;
        RECT 0.1580 10.7960 0.1760 10.8440 ;
        RECT 7.1780 10.7960 7.1960 10.8440 ;
        RECT 8.4200 10.7960 8.4470 10.8440 ;
        RECT 8.5730 10.7960 8.6090 10.8440 ;
        RECT 9.3380 10.7960 9.3560 10.8440 ;
        RECT 16.3580 10.7960 16.3760 10.8440 ;
        RECT 0.1580 11.8760 0.1760 11.9240 ;
        RECT 7.1780 11.8760 7.1960 11.9240 ;
        RECT 8.4200 11.8760 8.4470 11.9240 ;
        RECT 8.5730 11.8760 8.6090 11.9240 ;
        RECT 9.3380 11.8760 9.3560 11.9240 ;
        RECT 16.3580 11.8760 16.3760 11.9240 ;
        RECT 0.1580 12.9560 0.1760 13.0040 ;
        RECT 7.1780 12.9560 7.1960 13.0040 ;
        RECT 8.4200 12.9560 8.4470 13.0040 ;
        RECT 8.5730 12.9560 8.6090 13.0040 ;
        RECT 9.3380 12.9560 9.3560 13.0040 ;
        RECT 16.3580 12.9560 16.3760 13.0040 ;
        RECT 0.1580 14.0360 0.1760 14.0840 ;
        RECT 7.1780 14.0360 7.1960 14.0840 ;
        RECT 8.4200 14.0360 8.4470 14.0840 ;
        RECT 8.5730 14.0360 8.6090 14.0840 ;
        RECT 9.3380 14.0360 9.3560 14.0840 ;
        RECT 16.3580 14.0360 16.3760 14.0840 ;
        RECT 0.1580 15.1160 0.1760 15.1640 ;
        RECT 7.1780 15.1160 7.1960 15.1640 ;
        RECT 8.4200 15.1160 8.4470 15.1640 ;
        RECT 8.5730 15.1160 8.6090 15.1640 ;
        RECT 9.3380 15.1160 9.3560 15.1640 ;
        RECT 16.3580 15.1160 16.3760 15.1640 ;
        RECT 0.1580 16.1960 0.1760 16.2440 ;
        RECT 7.1780 16.1960 7.1960 16.2440 ;
        RECT 8.4200 16.1960 8.4470 16.2440 ;
        RECT 8.5730 16.1960 8.6090 16.2440 ;
        RECT 9.3380 16.1960 9.3560 16.2440 ;
        RECT 16.3580 16.1960 16.3760 16.2440 ;
        RECT 0.1580 17.2760 0.1760 17.3240 ;
        RECT 7.1780 17.2760 7.1960 17.3240 ;
        RECT 8.4200 17.2760 8.4470 17.3240 ;
        RECT 8.5730 17.2760 8.6090 17.3240 ;
        RECT 9.3380 17.2760 9.3560 17.3240 ;
        RECT 16.3580 17.2760 16.3760 17.3240 ;
        RECT 0.1580 18.3560 0.1760 18.4040 ;
        RECT 7.1780 18.3560 7.1960 18.4040 ;
        RECT 8.4200 18.3560 8.4470 18.4040 ;
        RECT 8.5730 18.3560 8.6090 18.4040 ;
        RECT 9.3380 18.3560 9.3560 18.4040 ;
        RECT 16.3580 18.3560 16.3760 18.4040 ;
        RECT 0.1580 19.4360 0.1760 19.4840 ;
        RECT 7.1780 19.4360 7.1960 19.4840 ;
        RECT 8.4200 19.4360 8.4470 19.4840 ;
        RECT 8.5730 19.4360 8.6090 19.4840 ;
        RECT 9.3380 19.4360 9.3560 19.4840 ;
        RECT 16.3580 19.4360 16.3760 19.4840 ;
        RECT 0.1580 20.5160 0.1760 20.5640 ;
        RECT 7.1780 20.5160 7.1960 20.5640 ;
        RECT 8.4200 20.5160 8.4470 20.5640 ;
        RECT 8.5730 20.5160 8.6090 20.5640 ;
        RECT 9.3380 20.5160 9.3560 20.5640 ;
        RECT 16.3580 20.5160 16.3760 20.5640 ;
        RECT 0.1580 21.5960 0.1760 21.6440 ;
        RECT 7.1780 21.5960 7.1960 21.6440 ;
        RECT 8.4200 21.5960 8.4470 21.6440 ;
        RECT 8.5730 21.5960 8.6090 21.6440 ;
        RECT 9.3380 21.5960 9.3560 21.6440 ;
        RECT 16.3580 21.5960 16.3760 21.6440 ;
        RECT 0.1580 22.6760 0.1760 22.7240 ;
        RECT 7.1780 22.6760 7.1960 22.7240 ;
        RECT 8.4200 22.6760 8.4470 22.7240 ;
        RECT 8.5730 22.6760 8.6090 22.7240 ;
        RECT 9.3380 22.6760 9.3560 22.7240 ;
        RECT 16.3580 22.6760 16.3760 22.7240 ;
        RECT 0.1580 23.7560 0.1760 23.8040 ;
        RECT 7.1780 23.7560 7.1960 23.8040 ;
        RECT 8.4200 23.7560 8.4470 23.8040 ;
        RECT 8.5730 23.7560 8.6090 23.8040 ;
        RECT 9.3380 23.7560 9.3560 23.8040 ;
        RECT 16.3580 23.7560 16.3760 23.8040 ;
        RECT 0.1580 24.8360 0.1760 24.8840 ;
        RECT 7.1780 24.8360 7.1960 24.8840 ;
        RECT 8.4200 24.8360 8.4470 24.8840 ;
        RECT 8.5730 24.8360 8.6090 24.8840 ;
        RECT 9.3380 24.8360 9.3560 24.8840 ;
        RECT 16.3580 24.8360 16.3760 24.8840 ;
        RECT 0.1580 25.9160 0.1760 25.9640 ;
        RECT 7.1780 25.9160 7.1960 25.9640 ;
        RECT 8.4200 25.9160 8.4470 25.9640 ;
        RECT 8.5730 25.9160 8.6090 25.9640 ;
        RECT 9.3380 25.9160 9.3560 25.9640 ;
        RECT 16.3580 25.9160 16.3760 25.9640 ;
        RECT 0.1580 26.9960 0.1760 27.0440 ;
        RECT 7.1780 26.9960 7.1960 27.0440 ;
        RECT 8.4200 26.9960 8.4470 27.0440 ;
        RECT 8.5730 26.9960 8.6090 27.0440 ;
        RECT 9.3380 26.9960 9.3560 27.0440 ;
        RECT 16.3580 26.9960 16.3760 27.0440 ;
        RECT 0.1580 28.0760 0.1760 28.1240 ;
        RECT 7.1780 28.0760 7.1960 28.1240 ;
        RECT 8.4200 28.0760 8.4470 28.1240 ;
        RECT 8.5730 28.0760 8.6090 28.1240 ;
        RECT 9.3380 28.0760 9.3560 28.1240 ;
        RECT 16.3580 28.0760 16.3760 28.1240 ;
        RECT 0.1580 29.1560 0.1760 29.2040 ;
        RECT 7.1780 29.1560 7.1960 29.2040 ;
        RECT 8.4200 29.1560 8.4470 29.2040 ;
        RECT 8.5730 29.1560 8.6090 29.2040 ;
        RECT 9.3380 29.1560 9.3560 29.2040 ;
        RECT 16.3580 29.1560 16.3760 29.2040 ;
        RECT 0.1580 30.2360 0.1760 30.2840 ;
        RECT 7.1780 30.2360 7.1960 30.2840 ;
        RECT 8.4200 30.2360 8.4470 30.2840 ;
        RECT 8.5730 30.2360 8.6090 30.2840 ;
        RECT 9.3380 30.2360 9.3560 30.2840 ;
        RECT 16.3580 30.2360 16.3760 30.2840 ;
        RECT 0.1580 31.3160 0.1760 31.3640 ;
        RECT 7.1780 31.3160 7.1960 31.3640 ;
        RECT 8.4200 31.3160 8.4470 31.3640 ;
        RECT 8.5730 31.3160 8.6090 31.3640 ;
        RECT 9.3380 31.3160 9.3560 31.3640 ;
        RECT 16.3580 31.3160 16.3760 31.3640 ;
        RECT 0.1580 32.3960 0.1760 32.4440 ;
        RECT 7.1780 32.3960 7.1960 32.4440 ;
        RECT 8.4200 32.3960 8.4470 32.4440 ;
        RECT 8.5730 32.3960 8.6090 32.4440 ;
        RECT 9.3380 32.3960 9.3560 32.4440 ;
        RECT 16.3580 32.3960 16.3760 32.4440 ;
        RECT 0.1580 33.4760 0.1760 33.5240 ;
        RECT 7.1780 33.4760 7.1960 33.5240 ;
        RECT 8.4200 33.4760 8.4470 33.5240 ;
        RECT 8.5730 33.4760 8.6090 33.5240 ;
        RECT 9.3380 33.4760 9.3560 33.5240 ;
        RECT 16.3580 33.4760 16.3760 33.5240 ;
        RECT 0.1580 34.5560 0.1760 34.6040 ;
        RECT 7.1780 34.5560 7.1960 34.6040 ;
        RECT 8.4200 34.5560 8.4470 34.6040 ;
        RECT 8.5730 34.5560 8.6090 34.6040 ;
        RECT 9.3380 34.5560 9.3560 34.6040 ;
        RECT 16.3580 34.5560 16.3760 34.6040 ;
        RECT 0.1580 35.6360 0.1760 35.6840 ;
        RECT 7.1780 35.6360 7.1960 35.6840 ;
        RECT 8.4200 35.6360 8.4470 35.6840 ;
        RECT 8.5730 35.6360 8.6090 35.6840 ;
        RECT 9.3380 35.6360 9.3560 35.6840 ;
        RECT 16.3580 35.6360 16.3760 35.6840 ;
        RECT 0.1580 36.7160 0.1760 36.7640 ;
        RECT 7.1780 36.7160 7.1960 36.7640 ;
        RECT 8.4200 36.7160 8.4470 36.7640 ;
        RECT 8.5730 36.7160 8.6090 36.7640 ;
        RECT 9.3380 36.7160 9.3560 36.7640 ;
        RECT 16.3580 36.7160 16.3760 36.7640 ;
        RECT 0.1580 37.7960 0.1760 37.8440 ;
        RECT 7.1780 37.7960 7.1960 37.8440 ;
        RECT 8.4200 37.7960 8.4470 37.8440 ;
        RECT 8.5730 37.7960 8.6090 37.8440 ;
        RECT 9.3380 37.7960 9.3560 37.8440 ;
        RECT 16.3580 37.7960 16.3760 37.8440 ;
        RECT 0.1580 38.8760 0.1760 38.9240 ;
        RECT 7.1780 38.8760 7.1960 38.9240 ;
        RECT 8.4200 38.8760 8.4470 38.9240 ;
        RECT 8.5730 38.8760 8.6090 38.9240 ;
        RECT 9.3380 38.8760 9.3560 38.9240 ;
        RECT 16.3580 38.8760 16.3760 38.9240 ;
        RECT 0.1580 39.9560 0.1760 40.0040 ;
        RECT 7.1780 39.9560 7.1960 40.0040 ;
        RECT 8.4200 39.9560 8.4470 40.0040 ;
        RECT 8.5730 39.9560 8.6090 40.0040 ;
        RECT 9.3380 39.9560 9.3560 40.0040 ;
        RECT 16.3580 39.9560 16.3760 40.0040 ;
        RECT 8.3830 47.3010 8.4010 47.5170 ;
        RECT 8.3830 44.1330 8.4010 44.3490 ;
        RECT 8.3830 40.9650 8.4010 41.1810 ;
        RECT 8.4350 47.3010 8.4530 47.5170 ;
        RECT 8.4350 44.1330 8.4530 44.3490 ;
        RECT 8.4350 40.9650 8.4530 41.1810 ;
        RECT 8.4870 47.3010 8.5050 47.5170 ;
        RECT 8.4870 44.1330 8.5050 44.3490 ;
        RECT 8.4870 40.9650 8.5050 41.1810 ;
        RECT 8.5390 47.3010 8.5570 47.5170 ;
        RECT 8.5390 44.1330 8.5570 44.3490 ;
        RECT 8.5390 40.9650 8.5570 41.1810 ;
        RECT 8.5910 47.3010 8.6090 47.5170 ;
        RECT 8.5910 44.1330 8.6090 44.3490 ;
        RECT 8.5910 40.9650 8.6090 41.1810 ;
        RECT 9.3330 40.9655 9.3510 41.1815 ;
        RECT 0.1580 49.1630 0.1760 49.2110 ;
        RECT 7.1780 49.1630 7.1960 49.2110 ;
        RECT 8.4200 49.1630 8.4470 49.2110 ;
        RECT 8.5730 49.1630 8.6090 49.2110 ;
        RECT 9.3380 49.1630 9.3560 49.2110 ;
        RECT 16.3580 49.1630 16.3760 49.2110 ;
        RECT 0.1580 50.2430 0.1760 50.2910 ;
        RECT 7.1780 50.2430 7.1960 50.2910 ;
        RECT 8.4200 50.2430 8.4470 50.2910 ;
        RECT 8.5730 50.2430 8.6090 50.2910 ;
        RECT 9.3380 50.2430 9.3560 50.2910 ;
        RECT 16.3580 50.2430 16.3760 50.2910 ;
        RECT 0.1580 51.3230 0.1760 51.3710 ;
        RECT 7.1780 51.3230 7.1960 51.3710 ;
        RECT 8.4200 51.3230 8.4470 51.3710 ;
        RECT 8.5730 51.3230 8.6090 51.3710 ;
        RECT 9.3380 51.3230 9.3560 51.3710 ;
        RECT 16.3580 51.3230 16.3760 51.3710 ;
        RECT 0.1580 52.4030 0.1760 52.4510 ;
        RECT 7.1780 52.4030 7.1960 52.4510 ;
        RECT 8.4200 52.4030 8.4470 52.4510 ;
        RECT 8.5730 52.4030 8.6090 52.4510 ;
        RECT 9.3380 52.4030 9.3560 52.4510 ;
        RECT 16.3580 52.4030 16.3760 52.4510 ;
        RECT 0.1580 53.4830 0.1760 53.5310 ;
        RECT 7.1780 53.4830 7.1960 53.5310 ;
        RECT 8.4200 53.4830 8.4470 53.5310 ;
        RECT 8.5730 53.4830 8.6090 53.5310 ;
        RECT 9.3380 53.4830 9.3560 53.5310 ;
        RECT 16.3580 53.4830 16.3760 53.5310 ;
        RECT 0.1580 54.5630 0.1760 54.6110 ;
        RECT 7.1780 54.5630 7.1960 54.6110 ;
        RECT 8.4200 54.5630 8.4470 54.6110 ;
        RECT 8.5730 54.5630 8.6090 54.6110 ;
        RECT 9.3380 54.5630 9.3560 54.6110 ;
        RECT 16.3580 54.5630 16.3760 54.6110 ;
        RECT 0.1580 55.6430 0.1760 55.6910 ;
        RECT 7.1780 55.6430 7.1960 55.6910 ;
        RECT 8.4200 55.6430 8.4470 55.6910 ;
        RECT 8.5730 55.6430 8.6090 55.6910 ;
        RECT 9.3380 55.6430 9.3560 55.6910 ;
        RECT 16.3580 55.6430 16.3760 55.6910 ;
        RECT 0.1580 56.7230 0.1760 56.7710 ;
        RECT 7.1780 56.7230 7.1960 56.7710 ;
        RECT 8.4200 56.7230 8.4470 56.7710 ;
        RECT 8.5730 56.7230 8.6090 56.7710 ;
        RECT 9.3380 56.7230 9.3560 56.7710 ;
        RECT 16.3580 56.7230 16.3760 56.7710 ;
        RECT 0.1580 57.8030 0.1760 57.8510 ;
        RECT 7.1780 57.8030 7.1960 57.8510 ;
        RECT 8.4200 57.8030 8.4470 57.8510 ;
        RECT 8.5730 57.8030 8.6090 57.8510 ;
        RECT 9.3380 57.8030 9.3560 57.8510 ;
        RECT 16.3580 57.8030 16.3760 57.8510 ;
        RECT 0.1580 58.8830 0.1760 58.9310 ;
        RECT 7.1780 58.8830 7.1960 58.9310 ;
        RECT 8.4200 58.8830 8.4470 58.9310 ;
        RECT 8.5730 58.8830 8.6090 58.9310 ;
        RECT 9.3380 58.8830 9.3560 58.9310 ;
        RECT 16.3580 58.8830 16.3760 58.9310 ;
        RECT 0.1580 59.9630 0.1760 60.0110 ;
        RECT 7.1780 59.9630 7.1960 60.0110 ;
        RECT 8.4200 59.9630 8.4470 60.0110 ;
        RECT 8.5730 59.9630 8.6090 60.0110 ;
        RECT 9.3380 59.9630 9.3560 60.0110 ;
        RECT 16.3580 59.9630 16.3760 60.0110 ;
        RECT 0.1580 61.0430 0.1760 61.0910 ;
        RECT 7.1780 61.0430 7.1960 61.0910 ;
        RECT 8.4200 61.0430 8.4470 61.0910 ;
        RECT 8.5730 61.0430 8.6090 61.0910 ;
        RECT 9.3380 61.0430 9.3560 61.0910 ;
        RECT 16.3580 61.0430 16.3760 61.0910 ;
        RECT 0.1580 62.1230 0.1760 62.1710 ;
        RECT 7.1780 62.1230 7.1960 62.1710 ;
        RECT 8.4200 62.1230 8.4470 62.1710 ;
        RECT 8.5730 62.1230 8.6090 62.1710 ;
        RECT 9.3380 62.1230 9.3560 62.1710 ;
        RECT 16.3580 62.1230 16.3760 62.1710 ;
        RECT 0.1580 63.2030 0.1760 63.2510 ;
        RECT 7.1780 63.2030 7.1960 63.2510 ;
        RECT 8.4200 63.2030 8.4470 63.2510 ;
        RECT 8.5730 63.2030 8.6090 63.2510 ;
        RECT 9.3380 63.2030 9.3560 63.2510 ;
        RECT 16.3580 63.2030 16.3760 63.2510 ;
        RECT 0.1580 64.2830 0.1760 64.3310 ;
        RECT 7.1780 64.2830 7.1960 64.3310 ;
        RECT 8.4200 64.2830 8.4470 64.3310 ;
        RECT 8.5730 64.2830 8.6090 64.3310 ;
        RECT 9.3380 64.2830 9.3560 64.3310 ;
        RECT 16.3580 64.2830 16.3760 64.3310 ;
        RECT 0.1580 65.3630 0.1760 65.4110 ;
        RECT 7.1780 65.3630 7.1960 65.4110 ;
        RECT 8.4200 65.3630 8.4470 65.4110 ;
        RECT 8.5730 65.3630 8.6090 65.4110 ;
        RECT 9.3380 65.3630 9.3560 65.4110 ;
        RECT 16.3580 65.3630 16.3760 65.4110 ;
        RECT 0.1580 66.4430 0.1760 66.4910 ;
        RECT 7.1780 66.4430 7.1960 66.4910 ;
        RECT 8.4200 66.4430 8.4470 66.4910 ;
        RECT 8.5730 66.4430 8.6090 66.4910 ;
        RECT 9.3380 66.4430 9.3560 66.4910 ;
        RECT 16.3580 66.4430 16.3760 66.4910 ;
        RECT 0.1580 67.5230 0.1760 67.5710 ;
        RECT 7.1780 67.5230 7.1960 67.5710 ;
        RECT 8.4200 67.5230 8.4470 67.5710 ;
        RECT 8.5730 67.5230 8.6090 67.5710 ;
        RECT 9.3380 67.5230 9.3560 67.5710 ;
        RECT 16.3580 67.5230 16.3760 67.5710 ;
        RECT 0.1580 68.6030 0.1760 68.6510 ;
        RECT 7.1780 68.6030 7.1960 68.6510 ;
        RECT 8.4200 68.6030 8.4470 68.6510 ;
        RECT 8.5730 68.6030 8.6090 68.6510 ;
        RECT 9.3380 68.6030 9.3560 68.6510 ;
        RECT 16.3580 68.6030 16.3760 68.6510 ;
        RECT 0.1580 69.6830 0.1760 69.7310 ;
        RECT 7.1780 69.6830 7.1960 69.7310 ;
        RECT 8.4200 69.6830 8.4470 69.7310 ;
        RECT 8.5730 69.6830 8.6090 69.7310 ;
        RECT 9.3380 69.6830 9.3560 69.7310 ;
        RECT 16.3580 69.6830 16.3760 69.7310 ;
        RECT 0.1580 70.7630 0.1760 70.8110 ;
        RECT 7.1780 70.7630 7.1960 70.8110 ;
        RECT 8.4200 70.7630 8.4470 70.8110 ;
        RECT 8.5730 70.7630 8.6090 70.8110 ;
        RECT 9.3380 70.7630 9.3560 70.8110 ;
        RECT 16.3580 70.7630 16.3760 70.8110 ;
        RECT 0.1580 71.8430 0.1760 71.8910 ;
        RECT 7.1780 71.8430 7.1960 71.8910 ;
        RECT 8.4200 71.8430 8.4470 71.8910 ;
        RECT 8.5730 71.8430 8.6090 71.8910 ;
        RECT 9.3380 71.8430 9.3560 71.8910 ;
        RECT 16.3580 71.8430 16.3760 71.8910 ;
        RECT 0.1580 72.9230 0.1760 72.9710 ;
        RECT 7.1780 72.9230 7.1960 72.9710 ;
        RECT 8.4200 72.9230 8.4470 72.9710 ;
        RECT 8.5730 72.9230 8.6090 72.9710 ;
        RECT 9.3380 72.9230 9.3560 72.9710 ;
        RECT 16.3580 72.9230 16.3760 72.9710 ;
        RECT 0.1580 74.0030 0.1760 74.0510 ;
        RECT 7.1780 74.0030 7.1960 74.0510 ;
        RECT 8.4200 74.0030 8.4470 74.0510 ;
        RECT 8.5730 74.0030 8.6090 74.0510 ;
        RECT 9.3380 74.0030 9.3560 74.0510 ;
        RECT 16.3580 74.0030 16.3760 74.0510 ;
        RECT 0.1580 75.0830 0.1760 75.1310 ;
        RECT 7.1780 75.0830 7.1960 75.1310 ;
        RECT 8.4200 75.0830 8.4470 75.1310 ;
        RECT 8.5730 75.0830 8.6090 75.1310 ;
        RECT 9.3380 75.0830 9.3560 75.1310 ;
        RECT 16.3580 75.0830 16.3760 75.1310 ;
        RECT 0.1580 76.1630 0.1760 76.2110 ;
        RECT 7.1780 76.1630 7.1960 76.2110 ;
        RECT 8.4200 76.1630 8.4470 76.2110 ;
        RECT 8.5730 76.1630 8.6090 76.2110 ;
        RECT 9.3380 76.1630 9.3560 76.2110 ;
        RECT 16.3580 76.1630 16.3760 76.2110 ;
        RECT 0.1580 77.2430 0.1760 77.2910 ;
        RECT 7.1780 77.2430 7.1960 77.2910 ;
        RECT 8.4200 77.2430 8.4470 77.2910 ;
        RECT 8.5730 77.2430 8.6090 77.2910 ;
        RECT 9.3380 77.2430 9.3560 77.2910 ;
        RECT 16.3580 77.2430 16.3760 77.2910 ;
        RECT 0.1580 78.3230 0.1760 78.3710 ;
        RECT 7.1780 78.3230 7.1960 78.3710 ;
        RECT 8.4200 78.3230 8.4470 78.3710 ;
        RECT 8.5730 78.3230 8.6090 78.3710 ;
        RECT 9.3380 78.3230 9.3560 78.3710 ;
        RECT 16.3580 78.3230 16.3760 78.3710 ;
        RECT 0.1580 79.4030 0.1760 79.4510 ;
        RECT 7.1780 79.4030 7.1960 79.4510 ;
        RECT 8.4200 79.4030 8.4470 79.4510 ;
        RECT 8.5730 79.4030 8.6090 79.4510 ;
        RECT 9.3380 79.4030 9.3560 79.4510 ;
        RECT 16.3580 79.4030 16.3760 79.4510 ;
        RECT 0.1580 80.4830 0.1760 80.5310 ;
        RECT 7.1780 80.4830 7.1960 80.5310 ;
        RECT 8.4200 80.4830 8.4470 80.5310 ;
        RECT 8.5730 80.4830 8.6090 80.5310 ;
        RECT 9.3380 80.4830 9.3560 80.5310 ;
        RECT 16.3580 80.4830 16.3760 80.5310 ;
        RECT 0.1580 81.5630 0.1760 81.6110 ;
        RECT 7.1780 81.5630 7.1960 81.6110 ;
        RECT 8.4200 81.5630 8.4470 81.6110 ;
        RECT 8.5730 81.5630 8.6090 81.6110 ;
        RECT 9.3380 81.5630 9.3560 81.6110 ;
        RECT 16.3580 81.5630 16.3760 81.6110 ;
        RECT 0.1580 82.6430 0.1760 82.6910 ;
        RECT 7.1780 82.6430 7.1960 82.6910 ;
        RECT 8.4200 82.6430 8.4470 82.6910 ;
        RECT 8.5730 82.6430 8.6090 82.6910 ;
        RECT 9.3380 82.6430 9.3560 82.6910 ;
        RECT 16.3580 82.6430 16.3760 82.6910 ;
        RECT 0.1580 83.7230 0.1760 83.7710 ;
        RECT 7.1780 83.7230 7.1960 83.7710 ;
        RECT 8.4200 83.7230 8.4470 83.7710 ;
        RECT 8.5730 83.7230 8.6090 83.7710 ;
        RECT 9.3380 83.7230 9.3560 83.7710 ;
        RECT 16.3580 83.7230 16.3760 83.7710 ;
        RECT 0.1580 84.8030 0.1760 84.8510 ;
        RECT 7.1780 84.8030 7.1960 84.8510 ;
        RECT 8.4200 84.8030 8.4470 84.8510 ;
        RECT 8.5730 84.8030 8.6090 84.8510 ;
        RECT 9.3380 84.8030 9.3560 84.8510 ;
        RECT 16.3580 84.8030 16.3760 84.8510 ;
        RECT 0.1580 85.8830 0.1760 85.9310 ;
        RECT 7.1780 85.8830 7.1960 85.9310 ;
        RECT 8.4200 85.8830 8.4470 85.9310 ;
        RECT 8.5730 85.8830 8.6090 85.9310 ;
        RECT 9.3380 85.8830 9.3560 85.9310 ;
        RECT 16.3580 85.8830 16.3760 85.9310 ;
        RECT 0.1580 86.9630 0.1760 87.0110 ;
        RECT 7.1780 86.9630 7.1960 87.0110 ;
        RECT 8.4200 86.9630 8.4470 87.0110 ;
        RECT 8.5730 86.9630 8.6090 87.0110 ;
        RECT 9.3380 86.9630 9.3560 87.0110 ;
        RECT 16.3580 86.9630 16.3760 87.0110 ;
        RECT 0.1580 88.0430 0.1760 88.0910 ;
        RECT 7.1780 88.0430 7.1960 88.0910 ;
        RECT 8.4200 88.0430 8.4470 88.0910 ;
        RECT 8.5730 88.0430 8.6090 88.0910 ;
        RECT 9.3380 88.0430 9.3560 88.0910 ;
        RECT 16.3580 88.0430 16.3760 88.0910 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.7910 41.4370 10.8090 41.4740 ;
      LAYER M4  ;
        RECT 10.7390 41.4450 10.8230 41.4690 ;
      LAYER M5  ;
        RECT 10.7880 40.4940 10.8120 43.7340 ;
      LAYER V3  ;
        RECT 10.7910 41.4450 10.8090 41.4690 ;
      LAYER V4  ;
        RECT 10.7880 41.4450 10.8120 41.4690 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.5750 41.4400 10.5930 41.4770 ;
      LAYER M4  ;
        RECT 10.5230 41.4450 10.6070 41.4690 ;
      LAYER M5  ;
        RECT 10.5720 40.4940 10.5960 43.7340 ;
      LAYER V3  ;
        RECT 10.5750 41.4450 10.5930 41.4690 ;
      LAYER V4  ;
        RECT 10.5720 41.4450 10.5960 41.4690 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.3590 40.8610 10.3770 40.8980 ;
      LAYER M4  ;
        RECT 10.3070 40.8690 10.3910 40.8930 ;
      LAYER M5  ;
        RECT 10.3560 40.4940 10.3800 43.7340 ;
      LAYER V3  ;
        RECT 10.3590 40.8690 10.3770 40.8930 ;
      LAYER V4  ;
        RECT 10.3560 40.8690 10.3800 40.8930 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.1430 41.1010 10.1610 41.2820 ;
      LAYER M4  ;
        RECT 10.0910 41.2530 10.1750 41.2770 ;
      LAYER M5  ;
        RECT 10.1400 40.4940 10.1640 43.7340 ;
      LAYER V3  ;
        RECT 10.1430 41.2530 10.1610 41.2770 ;
      LAYER V4  ;
        RECT 10.1400 41.2530 10.1640 41.2770 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.9270 40.8640 9.9450 40.9310 ;
      LAYER M4  ;
        RECT 9.8750 40.8690 9.9590 40.8930 ;
      LAYER M5  ;
        RECT 9.9240 40.4940 9.9480 43.7340 ;
      LAYER V3  ;
        RECT 9.9270 40.8690 9.9450 40.8930 ;
      LAYER V4  ;
        RECT 9.9240 40.8690 9.9480 40.8930 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.7110 40.5970 9.7290 40.8500 ;
      LAYER M4  ;
        RECT 9.6590 40.8210 9.7430 40.8450 ;
      LAYER M5  ;
        RECT 9.7080 40.4940 9.7320 43.7340 ;
      LAYER V3  ;
        RECT 9.7110 40.8210 9.7290 40.8450 ;
      LAYER V4  ;
        RECT 9.7080 40.8210 9.7320 40.8450 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.4950 41.6320 9.5130 41.6690 ;
      LAYER M4  ;
        RECT 9.4430 41.6370 9.5270 41.6610 ;
      LAYER M5  ;
        RECT 9.4920 40.4940 9.5160 43.7340 ;
      LAYER V3  ;
        RECT 9.4950 41.6370 9.5130 41.6610 ;
      LAYER V4  ;
        RECT 9.4920 41.6370 9.5160 41.6610 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.2790 41.4790 9.2970 41.5700 ;
      LAYER M4  ;
        RECT 9.2270 41.5410 9.3110 41.5650 ;
      LAYER M5  ;
        RECT 9.2760 40.4940 9.3000 43.7340 ;
      LAYER V3  ;
        RECT 9.2790 41.5410 9.2970 41.5650 ;
      LAYER V4  ;
        RECT 9.2760 41.5410 9.3000 41.5650 ;
    END
  END ADDRESS[7]
  PIN ADDRESS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.6310 40.8640 8.6490 40.9310 ;
      LAYER M4  ;
        RECT 8.3470 40.8690 8.6600 40.8930 ;
      LAYER M5  ;
        RECT 8.3580 40.4940 8.3820 43.7340 ;
      LAYER V3  ;
        RECT 8.6310 40.8690 8.6490 40.8930 ;
      LAYER V4  ;
        RECT 8.3580 40.8690 8.3820 40.8930 ;
    END
  END ADDRESS[8]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.2350 40.5970 8.2530 40.8500 ;
      LAYER M4  ;
        RECT 8.0230 40.8210 8.2640 40.8450 ;
      LAYER M5  ;
        RECT 8.0340 40.4940 8.0580 43.7340 ;
      LAYER V3  ;
        RECT 8.2350 40.8210 8.2530 40.8450 ;
      LAYER V4  ;
        RECT 8.0340 40.8210 8.0580 40.8450 ;
    END
  END banksel
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.4430 40.8640 7.4610 40.9310 ;
      LAYER M4  ;
        RECT 7.3910 40.8690 7.4750 40.8930 ;
      LAYER M5  ;
        RECT 7.4400 40.4940 7.4640 43.7340 ;
      LAYER V3  ;
        RECT 7.4430 40.8690 7.4610 40.8930 ;
      LAYER V4  ;
        RECT 7.4400 40.8690 7.4640 40.8930 ;
    END
  END write
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2270 41.7280 7.2450 41.7770 ;
      LAYER M4  ;
        RECT 7.1750 41.7330 7.2590 41.7570 ;
      LAYER M5  ;
        RECT 7.2240 40.4940 7.2480 43.7340 ;
      LAYER V3  ;
        RECT 7.2270 41.7330 7.2450 41.7570 ;
      LAYER V4  ;
        RECT 7.2240 41.7330 7.2480 41.7570 ;
    END
  END clk
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2630 40.5970 7.2810 40.8500 ;
      LAYER M4  ;
        RECT 6.9970 40.8210 7.2920 40.8450 ;
      LAYER M5  ;
        RECT 7.0080 40.4940 7.0320 43.7340 ;
      LAYER V3  ;
        RECT 7.2630 40.8210 7.2810 40.8450 ;
      LAYER V4  ;
        RECT 7.0080 40.8210 7.0320 40.8450 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.7950 41.4370 6.8130 41.4740 ;
      LAYER M4  ;
        RECT 6.7430 41.4450 6.8270 41.4690 ;
      LAYER M5  ;
        RECT 6.7920 40.4940 6.8160 43.7340 ;
      LAYER V3  ;
        RECT 6.7950 41.4450 6.8130 41.4690 ;
      LAYER V4  ;
        RECT 6.7920 41.4450 6.8160 41.4690 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.5790 40.8640 6.5970 41.0930 ;
      LAYER M4  ;
        RECT 6.5270 40.8690 6.6110 40.8930 ;
      LAYER M5  ;
        RECT 6.5760 40.4940 6.6000 43.7340 ;
      LAYER V3  ;
        RECT 6.5790 40.8690 6.5970 40.8930 ;
      LAYER V4  ;
        RECT 6.5760 40.8690 6.6000 40.8930 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.3630 40.5970 6.3810 40.8500 ;
      LAYER M4  ;
        RECT 6.3110 40.8210 6.3950 40.8450 ;
      LAYER M5  ;
        RECT 6.3600 40.4940 6.3840 43.7340 ;
      LAYER V3  ;
        RECT 6.3630 40.8210 6.3810 40.8450 ;
      LAYER V4  ;
        RECT 6.3600 40.8210 6.3840 40.8450 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.1470 40.8610 6.1650 40.8980 ;
      LAYER M4  ;
        RECT 6.0950 40.8690 6.1790 40.8930 ;
      LAYER M5  ;
        RECT 6.1440 40.4940 6.1680 43.7340 ;
      LAYER V3  ;
        RECT 6.1470 40.8690 6.1650 40.8930 ;
      LAYER V4  ;
        RECT 6.1440 40.8690 6.1680 40.8930 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 5.9310 41.4370 5.9490 41.4740 ;
      LAYER M4  ;
        RECT 5.8790 41.4450 5.9630 41.4690 ;
      LAYER M5  ;
        RECT 5.9280 40.4940 5.9520 43.7340 ;
      LAYER V3  ;
        RECT 5.9310 41.4450 5.9490 41.4690 ;
      LAYER V4  ;
        RECT 5.9280 41.4450 5.9520 41.4690 ;
    END
  END sdel[4]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.4280 8.5970 0.4520 ;
      LAYER M3  ;
        RECT 8.5370 0.3775 8.5550 0.6170 ;
      LAYER V3  ;
        RECT 8.5370 0.4280 8.5550 0.4520 ;
    END
  END dataout[0]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.3320 8.6650 0.3560 ;
      LAYER M3  ;
        RECT 8.3120 0.2700 8.3300 0.6750 ;
      LAYER V3  ;
        RECT 8.3120 0.3320 8.3300 0.3560 ;
    END
  END wd[0]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.5080 8.5970 1.5320 ;
      LAYER M3  ;
        RECT 8.5370 1.4575 8.5550 1.6970 ;
      LAYER V3  ;
        RECT 8.5370 1.5080 8.5550 1.5320 ;
    END
  END dataout[1]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.4120 8.6650 1.4360 ;
      LAYER M3  ;
        RECT 8.3120 1.3500 8.3300 1.7550 ;
      LAYER V3  ;
        RECT 8.3120 1.4120 8.3300 1.4360 ;
    END
  END wd[1]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.5880 8.5970 2.6120 ;
      LAYER M3  ;
        RECT 8.5370 2.5375 8.5550 2.7770 ;
      LAYER V3  ;
        RECT 8.5370 2.5880 8.5550 2.6120 ;
    END
  END dataout[2]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.4920 8.6650 2.5160 ;
      LAYER M3  ;
        RECT 8.3120 2.4300 8.3300 2.8350 ;
      LAYER V3  ;
        RECT 8.3120 2.4920 8.3300 2.5160 ;
    END
  END wd[2]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.6680 8.5970 3.6920 ;
      LAYER M3  ;
        RECT 8.5370 3.6175 8.5550 3.8570 ;
      LAYER V3  ;
        RECT 8.5370 3.6680 8.5550 3.6920 ;
    END
  END dataout[3]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.5720 8.6650 3.5960 ;
      LAYER M3  ;
        RECT 8.3120 3.5100 8.3300 3.9150 ;
      LAYER V3  ;
        RECT 8.3120 3.5720 8.3300 3.5960 ;
    END
  END wd[3]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.7480 8.5970 4.7720 ;
      LAYER M3  ;
        RECT 8.5370 4.6975 8.5550 4.9370 ;
      LAYER V3  ;
        RECT 8.5370 4.7480 8.5550 4.7720 ;
    END
  END dataout[4]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.6520 8.6650 4.6760 ;
      LAYER M3  ;
        RECT 8.3120 4.5900 8.3300 4.9950 ;
      LAYER V3  ;
        RECT 8.3120 4.6520 8.3300 4.6760 ;
    END
  END wd[4]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.8280 8.5970 5.8520 ;
      LAYER M3  ;
        RECT 8.5370 5.7775 8.5550 6.0170 ;
      LAYER V3  ;
        RECT 8.5370 5.8280 8.5550 5.8520 ;
    END
  END dataout[5]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.7320 8.6650 5.7560 ;
      LAYER M3  ;
        RECT 8.3120 5.6700 8.3300 6.0750 ;
      LAYER V3  ;
        RECT 8.3120 5.7320 8.3300 5.7560 ;
    END
  END wd[5]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.9080 8.5970 6.9320 ;
      LAYER M3  ;
        RECT 8.5370 6.8575 8.5550 7.0970 ;
      LAYER V3  ;
        RECT 8.5370 6.9080 8.5550 6.9320 ;
    END
  END dataout[6]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.8120 8.6650 6.8360 ;
      LAYER M3  ;
        RECT 8.3120 6.7500 8.3300 7.1550 ;
      LAYER V3  ;
        RECT 8.3120 6.8120 8.3300 6.8360 ;
    END
  END wd[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.9880 8.5970 8.0120 ;
      LAYER M3  ;
        RECT 8.5370 7.9375 8.5550 8.1770 ;
      LAYER V3  ;
        RECT 8.5370 7.9880 8.5550 8.0120 ;
    END
  END dataout[7]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.8920 8.6650 7.9160 ;
      LAYER M3  ;
        RECT 8.3120 7.8300 8.3300 8.2350 ;
      LAYER V3  ;
        RECT 8.3120 7.8920 8.3300 7.9160 ;
    END
  END wd[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 9.0680 8.5970 9.0920 ;
      LAYER M3  ;
        RECT 8.5370 9.0175 8.5550 9.2570 ;
      LAYER V3  ;
        RECT 8.5370 9.0680 8.5550 9.0920 ;
    END
  END dataout[8]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 8.9720 8.6650 8.9960 ;
      LAYER M3  ;
        RECT 8.3120 8.9100 8.3300 9.3150 ;
      LAYER V3  ;
        RECT 8.3120 8.9720 8.3300 8.9960 ;
    END
  END wd[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 10.1480 8.5970 10.1720 ;
      LAYER M3  ;
        RECT 8.5370 10.0975 8.5550 10.3370 ;
      LAYER V3  ;
        RECT 8.5370 10.1480 8.5550 10.1720 ;
    END
  END dataout[9]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 10.0520 8.6650 10.0760 ;
      LAYER M3  ;
        RECT 8.3120 9.9900 8.3300 10.3950 ;
      LAYER V3  ;
        RECT 8.3120 10.0520 8.3300 10.0760 ;
    END
  END wd[9]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 11.2280 8.5970 11.2520 ;
      LAYER M3  ;
        RECT 8.5370 11.1775 8.5550 11.4170 ;
      LAYER V3  ;
        RECT 8.5370 11.2280 8.5550 11.2520 ;
    END
  END dataout[10]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 11.1320 8.6650 11.1560 ;
      LAYER M3  ;
        RECT 8.3120 11.0700 8.3300 11.4750 ;
      LAYER V3  ;
        RECT 8.3120 11.1320 8.3300 11.1560 ;
    END
  END wd[10]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 12.3080 8.5970 12.3320 ;
      LAYER M3  ;
        RECT 8.5370 12.2575 8.5550 12.4970 ;
      LAYER V3  ;
        RECT 8.5370 12.3080 8.5550 12.3320 ;
    END
  END dataout[11]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 12.2120 8.6650 12.2360 ;
      LAYER M3  ;
        RECT 8.3120 12.1500 8.3300 12.5550 ;
      LAYER V3  ;
        RECT 8.3120 12.2120 8.3300 12.2360 ;
    END
  END wd[11]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 13.3880 8.5970 13.4120 ;
      LAYER M3  ;
        RECT 8.5370 13.3375 8.5550 13.5770 ;
      LAYER V3  ;
        RECT 8.5370 13.3880 8.5550 13.4120 ;
    END
  END dataout[12]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 13.2920 8.6650 13.3160 ;
      LAYER M3  ;
        RECT 8.3120 13.2300 8.3300 13.6350 ;
      LAYER V3  ;
        RECT 8.3120 13.2920 8.3300 13.3160 ;
    END
  END wd[12]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 14.4680 8.5970 14.4920 ;
      LAYER M3  ;
        RECT 8.5370 14.4175 8.5550 14.6570 ;
      LAYER V3  ;
        RECT 8.5370 14.4680 8.5550 14.4920 ;
    END
  END dataout[13]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 14.3720 8.6650 14.3960 ;
      LAYER M3  ;
        RECT 8.3120 14.3100 8.3300 14.7150 ;
      LAYER V3  ;
        RECT 8.3120 14.3720 8.3300 14.3960 ;
    END
  END wd[13]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 15.5480 8.5970 15.5720 ;
      LAYER M3  ;
        RECT 8.5370 15.4975 8.5550 15.7370 ;
      LAYER V3  ;
        RECT 8.5370 15.5480 8.5550 15.5720 ;
    END
  END dataout[14]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 15.4520 8.6650 15.4760 ;
      LAYER M3  ;
        RECT 8.3120 15.3900 8.3300 15.7950 ;
      LAYER V3  ;
        RECT 8.3120 15.4520 8.3300 15.4760 ;
    END
  END wd[14]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 16.6280 8.5970 16.6520 ;
      LAYER M3  ;
        RECT 8.5370 16.5775 8.5550 16.8170 ;
      LAYER V3  ;
        RECT 8.5370 16.6280 8.5550 16.6520 ;
    END
  END dataout[15]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 16.5320 8.6650 16.5560 ;
      LAYER M3  ;
        RECT 8.3120 16.4700 8.3300 16.8750 ;
      LAYER V3  ;
        RECT 8.3120 16.5320 8.3300 16.5560 ;
    END
  END wd[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 17.7080 8.5970 17.7320 ;
      LAYER M3  ;
        RECT 8.5370 17.6575 8.5550 17.8970 ;
      LAYER V3  ;
        RECT 8.5370 17.7080 8.5550 17.7320 ;
    END
  END dataout[16]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 17.6120 8.6650 17.6360 ;
      LAYER M3  ;
        RECT 8.3120 17.5500 8.3300 17.9550 ;
      LAYER V3  ;
        RECT 8.3120 17.6120 8.3300 17.6360 ;
    END
  END wd[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 18.7880 8.5970 18.8120 ;
      LAYER M3  ;
        RECT 8.5370 18.7375 8.5550 18.9770 ;
      LAYER V3  ;
        RECT 8.5370 18.7880 8.5550 18.8120 ;
    END
  END dataout[17]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 18.6920 8.6650 18.7160 ;
      LAYER M3  ;
        RECT 8.3120 18.6300 8.3300 19.0350 ;
      LAYER V3  ;
        RECT 8.3120 18.6920 8.3300 18.7160 ;
    END
  END wd[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.8680 8.5970 19.8920 ;
      LAYER M3  ;
        RECT 8.5370 19.8175 8.5550 20.0570 ;
      LAYER V3  ;
        RECT 8.5370 19.8680 8.5550 19.8920 ;
    END
  END dataout[18]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.7720 8.6650 19.7960 ;
      LAYER M3  ;
        RECT 8.3120 19.7100 8.3300 20.1150 ;
      LAYER V3  ;
        RECT 8.3120 19.7720 8.3300 19.7960 ;
    END
  END wd[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.9480 8.5970 20.9720 ;
      LAYER M3  ;
        RECT 8.5370 20.8975 8.5550 21.1370 ;
      LAYER V3  ;
        RECT 8.5370 20.9480 8.5550 20.9720 ;
    END
  END dataout[19]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.8520 8.6650 20.8760 ;
      LAYER M3  ;
        RECT 8.3120 20.7900 8.3300 21.1950 ;
      LAYER V3  ;
        RECT 8.3120 20.8520 8.3300 20.8760 ;
    END
  END wd[19]
  PIN dataout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 22.0280 8.5970 22.0520 ;
      LAYER M3  ;
        RECT 8.5370 21.9775 8.5550 22.2170 ;
      LAYER V3  ;
        RECT 8.5370 22.0280 8.5550 22.0520 ;
    END
  END dataout[20]
  PIN wd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 21.9320 8.6650 21.9560 ;
      LAYER M3  ;
        RECT 8.3120 21.8700 8.3300 22.2750 ;
      LAYER V3  ;
        RECT 8.3120 21.9320 8.3300 21.9560 ;
    END
  END wd[20]
  PIN dataout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.1080 8.5970 23.1320 ;
      LAYER M3  ;
        RECT 8.5370 23.0575 8.5550 23.2970 ;
      LAYER V3  ;
        RECT 8.5370 23.1080 8.5550 23.1320 ;
    END
  END dataout[21]
  PIN wd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.0120 8.6650 23.0360 ;
      LAYER M3  ;
        RECT 8.3120 22.9500 8.3300 23.3550 ;
      LAYER V3  ;
        RECT 8.3120 23.0120 8.3300 23.0360 ;
    END
  END wd[21]
  PIN dataout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.1880 8.5970 24.2120 ;
      LAYER M3  ;
        RECT 8.5370 24.1375 8.5550 24.3770 ;
      LAYER V3  ;
        RECT 8.5370 24.1880 8.5550 24.2120 ;
    END
  END dataout[22]
  PIN wd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.0920 8.6650 24.1160 ;
      LAYER M3  ;
        RECT 8.3120 24.0300 8.3300 24.4350 ;
      LAYER V3  ;
        RECT 8.3120 24.0920 8.3300 24.1160 ;
    END
  END wd[22]
  PIN dataout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.2680 8.5970 25.2920 ;
      LAYER M3  ;
        RECT 8.5370 25.2175 8.5550 25.4570 ;
      LAYER V3  ;
        RECT 8.5370 25.2680 8.5550 25.2920 ;
    END
  END dataout[23]
  PIN wd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.1720 8.6650 25.1960 ;
      LAYER M3  ;
        RECT 8.3120 25.1100 8.3300 25.5150 ;
      LAYER V3  ;
        RECT 8.3120 25.1720 8.3300 25.1960 ;
    END
  END wd[23]
  PIN dataout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 26.3480 8.5970 26.3720 ;
      LAYER M3  ;
        RECT 8.5370 26.2975 8.5550 26.5370 ;
      LAYER V3  ;
        RECT 8.5370 26.3480 8.5550 26.3720 ;
    END
  END dataout[24]
  PIN wd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 26.2520 8.6650 26.2760 ;
      LAYER M3  ;
        RECT 8.3120 26.1900 8.3300 26.5950 ;
      LAYER V3  ;
        RECT 8.3120 26.2520 8.3300 26.2760 ;
    END
  END wd[24]
  PIN dataout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 27.4280 8.5970 27.4520 ;
      LAYER M3  ;
        RECT 8.5370 27.3775 8.5550 27.6170 ;
      LAYER V3  ;
        RECT 8.5370 27.4280 8.5550 27.4520 ;
    END
  END dataout[25]
  PIN wd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 27.3320 8.6650 27.3560 ;
      LAYER M3  ;
        RECT 8.3120 27.2700 8.3300 27.6750 ;
      LAYER V3  ;
        RECT 8.3120 27.3320 8.3300 27.3560 ;
    END
  END wd[25]
  PIN dataout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 28.5080 8.5970 28.5320 ;
      LAYER M3  ;
        RECT 8.5370 28.4575 8.5550 28.6970 ;
      LAYER V3  ;
        RECT 8.5370 28.5080 8.5550 28.5320 ;
    END
  END dataout[26]
  PIN wd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 28.4120 8.6650 28.4360 ;
      LAYER M3  ;
        RECT 8.3120 28.3500 8.3300 28.7550 ;
      LAYER V3  ;
        RECT 8.3120 28.4120 8.3300 28.4360 ;
    END
  END wd[26]
  PIN dataout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 29.5880 8.5970 29.6120 ;
      LAYER M3  ;
        RECT 8.5370 29.5375 8.5550 29.7770 ;
      LAYER V3  ;
        RECT 8.5370 29.5880 8.5550 29.6120 ;
    END
  END dataout[27]
  PIN wd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 29.4920 8.6650 29.5160 ;
      LAYER M3  ;
        RECT 8.3120 29.4300 8.3300 29.8350 ;
      LAYER V3  ;
        RECT 8.3120 29.4920 8.3300 29.5160 ;
    END
  END wd[27]
  PIN dataout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 30.6680 8.5970 30.6920 ;
      LAYER M3  ;
        RECT 8.5370 30.6175 8.5550 30.8570 ;
      LAYER V3  ;
        RECT 8.5370 30.6680 8.5550 30.6920 ;
    END
  END dataout[28]
  PIN wd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 30.5720 8.6650 30.5960 ;
      LAYER M3  ;
        RECT 8.3120 30.5100 8.3300 30.9150 ;
      LAYER V3  ;
        RECT 8.3120 30.5720 8.3300 30.5960 ;
    END
  END wd[28]
  PIN dataout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 31.7480 8.5970 31.7720 ;
      LAYER M3  ;
        RECT 8.5370 31.6975 8.5550 31.9370 ;
      LAYER V3  ;
        RECT 8.5370 31.7480 8.5550 31.7720 ;
    END
  END dataout[29]
  PIN wd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 31.6520 8.6650 31.6760 ;
      LAYER M3  ;
        RECT 8.3120 31.5900 8.3300 31.9950 ;
      LAYER V3  ;
        RECT 8.3120 31.6520 8.3300 31.6760 ;
    END
  END wd[29]
  PIN dataout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 32.8280 8.5970 32.8520 ;
      LAYER M3  ;
        RECT 8.5370 32.7775 8.5550 33.0170 ;
      LAYER V3  ;
        RECT 8.5370 32.8280 8.5550 32.8520 ;
    END
  END dataout[30]
  PIN wd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 32.7320 8.6650 32.7560 ;
      LAYER M3  ;
        RECT 8.3120 32.6700 8.3300 33.0750 ;
      LAYER V3  ;
        RECT 8.3120 32.7320 8.3300 32.7560 ;
    END
  END wd[30]
  PIN dataout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 33.9080 8.5970 33.9320 ;
      LAYER M3  ;
        RECT 8.5370 33.8575 8.5550 34.0970 ;
      LAYER V3  ;
        RECT 8.5370 33.9080 8.5550 33.9320 ;
    END
  END dataout[31]
  PIN wd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 33.8120 8.6650 33.8360 ;
      LAYER M3  ;
        RECT 8.3120 33.7500 8.3300 34.1550 ;
      LAYER V3  ;
        RECT 8.3120 33.8120 8.3300 33.8360 ;
    END
  END wd[31]
  PIN dataout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 34.9880 8.5970 35.0120 ;
      LAYER M3  ;
        RECT 8.5370 34.9375 8.5550 35.1770 ;
      LAYER V3  ;
        RECT 8.5370 34.9880 8.5550 35.0120 ;
    END
  END dataout[32]
  PIN wd[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 34.8920 8.6650 34.9160 ;
      LAYER M3  ;
        RECT 8.3120 34.8300 8.3300 35.2350 ;
      LAYER V3  ;
        RECT 8.3120 34.8920 8.3300 34.9160 ;
    END
  END wd[32]
  PIN dataout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 36.0680 8.5970 36.0920 ;
      LAYER M3  ;
        RECT 8.5370 36.0175 8.5550 36.2570 ;
      LAYER V3  ;
        RECT 8.5370 36.0680 8.5550 36.0920 ;
    END
  END dataout[33]
  PIN wd[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 35.9720 8.6650 35.9960 ;
      LAYER M3  ;
        RECT 8.3120 35.9100 8.3300 36.3150 ;
      LAYER V3  ;
        RECT 8.3120 35.9720 8.3300 35.9960 ;
    END
  END wd[33]
  PIN dataout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 37.1480 8.5970 37.1720 ;
      LAYER M3  ;
        RECT 8.5370 37.0975 8.5550 37.3370 ;
      LAYER V3  ;
        RECT 8.5370 37.1480 8.5550 37.1720 ;
    END
  END dataout[34]
  PIN wd[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 37.0520 8.6650 37.0760 ;
      LAYER M3  ;
        RECT 8.3120 36.9900 8.3300 37.3950 ;
      LAYER V3  ;
        RECT 8.3120 37.0520 8.3300 37.0760 ;
    END
  END wd[34]
  PIN dataout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 38.2280 8.5970 38.2520 ;
      LAYER M3  ;
        RECT 8.5370 38.1775 8.5550 38.4170 ;
      LAYER V3  ;
        RECT 8.5370 38.2280 8.5550 38.2520 ;
    END
  END dataout[35]
  PIN wd[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 38.1320 8.6650 38.1560 ;
      LAYER M3  ;
        RECT 8.3120 38.0700 8.3300 38.4750 ;
      LAYER V3  ;
        RECT 8.3120 38.1320 8.3300 38.1560 ;
    END
  END wd[35]
  PIN dataout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 39.3080 8.5970 39.3320 ;
      LAYER M3  ;
        RECT 8.5370 39.2575 8.5550 39.4970 ;
      LAYER V3  ;
        RECT 8.5370 39.3080 8.5550 39.3320 ;
    END
  END dataout[36]
  PIN wd[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 39.2120 8.6650 39.2360 ;
      LAYER M3  ;
        RECT 8.3120 39.1500 8.3300 39.5550 ;
      LAYER V3  ;
        RECT 8.3120 39.2120 8.3300 39.2360 ;
    END
  END wd[36]
  PIN dataout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 48.5150 8.5970 48.5390 ;
      LAYER M3  ;
        RECT 8.5370 48.4645 8.5550 48.7040 ;
      LAYER V3  ;
        RECT 8.5370 48.5150 8.5550 48.5390 ;
    END
  END dataout[37]
  PIN wd[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 48.4190 8.6650 48.4430 ;
      LAYER M3  ;
        RECT 8.3120 48.3570 8.3300 48.7620 ;
      LAYER V3  ;
        RECT 8.3120 48.4190 8.3300 48.4430 ;
    END
  END wd[37]
  PIN dataout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 49.5950 8.5970 49.6190 ;
      LAYER M3  ;
        RECT 8.5370 49.5445 8.5550 49.7840 ;
      LAYER V3  ;
        RECT 8.5370 49.5950 8.5550 49.6190 ;
    END
  END dataout[38]
  PIN wd[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 49.4990 8.6650 49.5230 ;
      LAYER M3  ;
        RECT 8.3120 49.4370 8.3300 49.8420 ;
      LAYER V3  ;
        RECT 8.3120 49.4990 8.3300 49.5230 ;
    END
  END wd[38]
  PIN dataout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 50.6750 8.5970 50.6990 ;
      LAYER M3  ;
        RECT 8.5370 50.6245 8.5550 50.8640 ;
      LAYER V3  ;
        RECT 8.5370 50.6750 8.5550 50.6990 ;
    END
  END dataout[39]
  PIN wd[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 50.5790 8.6650 50.6030 ;
      LAYER M3  ;
        RECT 8.3120 50.5170 8.3300 50.9220 ;
      LAYER V3  ;
        RECT 8.3120 50.5790 8.3300 50.6030 ;
    END
  END wd[39]
  PIN dataout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 51.7550 8.5970 51.7790 ;
      LAYER M3  ;
        RECT 8.5370 51.7045 8.5550 51.9440 ;
      LAYER V3  ;
        RECT 8.5370 51.7550 8.5550 51.7790 ;
    END
  END dataout[40]
  PIN wd[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 51.6590 8.6650 51.6830 ;
      LAYER M3  ;
        RECT 8.3120 51.5970 8.3300 52.0020 ;
      LAYER V3  ;
        RECT 8.3120 51.6590 8.3300 51.6830 ;
    END
  END wd[40]
  PIN dataout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 52.8350 8.5970 52.8590 ;
      LAYER M3  ;
        RECT 8.5370 52.7845 8.5550 53.0240 ;
      LAYER V3  ;
        RECT 8.5370 52.8350 8.5550 52.8590 ;
    END
  END dataout[41]
  PIN wd[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 52.7390 8.6650 52.7630 ;
      LAYER M3  ;
        RECT 8.3120 52.6770 8.3300 53.0820 ;
      LAYER V3  ;
        RECT 8.3120 52.7390 8.3300 52.7630 ;
    END
  END wd[41]
  PIN dataout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 53.9150 8.5970 53.9390 ;
      LAYER M3  ;
        RECT 8.5370 53.8645 8.5550 54.1040 ;
      LAYER V3  ;
        RECT 8.5370 53.9150 8.5550 53.9390 ;
    END
  END dataout[42]
  PIN wd[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 53.8190 8.6650 53.8430 ;
      LAYER M3  ;
        RECT 8.3120 53.7570 8.3300 54.1620 ;
      LAYER V3  ;
        RECT 8.3120 53.8190 8.3300 53.8430 ;
    END
  END wd[42]
  PIN dataout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 54.9950 8.5970 55.0190 ;
      LAYER M3  ;
        RECT 8.5370 54.9445 8.5550 55.1840 ;
      LAYER V3  ;
        RECT 8.5370 54.9950 8.5550 55.0190 ;
    END
  END dataout[43]
  PIN wd[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 54.8990 8.6650 54.9230 ;
      LAYER M3  ;
        RECT 8.3120 54.8370 8.3300 55.2420 ;
      LAYER V3  ;
        RECT 8.3120 54.8990 8.3300 54.9230 ;
    END
  END wd[43]
  PIN dataout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 56.0750 8.5970 56.0990 ;
      LAYER M3  ;
        RECT 8.5370 56.0245 8.5550 56.2640 ;
      LAYER V3  ;
        RECT 8.5370 56.0750 8.5550 56.0990 ;
    END
  END dataout[44]
  PIN wd[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 55.9790 8.6650 56.0030 ;
      LAYER M3  ;
        RECT 8.3120 55.9170 8.3300 56.3220 ;
      LAYER V3  ;
        RECT 8.3120 55.9790 8.3300 56.0030 ;
    END
  END wd[44]
  PIN dataout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 57.1550 8.5970 57.1790 ;
      LAYER M3  ;
        RECT 8.5370 57.1045 8.5550 57.3440 ;
      LAYER V3  ;
        RECT 8.5370 57.1550 8.5550 57.1790 ;
    END
  END dataout[45]
  PIN wd[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 57.0590 8.6650 57.0830 ;
      LAYER M3  ;
        RECT 8.3120 56.9970 8.3300 57.4020 ;
      LAYER V3  ;
        RECT 8.3120 57.0590 8.3300 57.0830 ;
    END
  END wd[45]
  PIN dataout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 58.2350 8.5970 58.2590 ;
      LAYER M3  ;
        RECT 8.5370 58.1845 8.5550 58.4240 ;
      LAYER V3  ;
        RECT 8.5370 58.2350 8.5550 58.2590 ;
    END
  END dataout[46]
  PIN wd[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 58.1390 8.6650 58.1630 ;
      LAYER M3  ;
        RECT 8.3120 58.0770 8.3300 58.4820 ;
      LAYER V3  ;
        RECT 8.3120 58.1390 8.3300 58.1630 ;
    END
  END wd[46]
  PIN dataout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 59.3150 8.5970 59.3390 ;
      LAYER M3  ;
        RECT 8.5370 59.2645 8.5550 59.5040 ;
      LAYER V3  ;
        RECT 8.5370 59.3150 8.5550 59.3390 ;
    END
  END dataout[47]
  PIN wd[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 59.2190 8.6650 59.2430 ;
      LAYER M3  ;
        RECT 8.3120 59.1570 8.3300 59.5620 ;
      LAYER V3  ;
        RECT 8.3120 59.2190 8.3300 59.2430 ;
    END
  END wd[47]
  PIN dataout[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 60.3950 8.5970 60.4190 ;
      LAYER M3  ;
        RECT 8.5370 60.3445 8.5550 60.5840 ;
      LAYER V3  ;
        RECT 8.5370 60.3950 8.5550 60.4190 ;
    END
  END dataout[48]
  PIN wd[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 60.2990 8.6650 60.3230 ;
      LAYER M3  ;
        RECT 8.3120 60.2370 8.3300 60.6420 ;
      LAYER V3  ;
        RECT 8.3120 60.2990 8.3300 60.3230 ;
    END
  END wd[48]
  PIN dataout[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 61.4750 8.5970 61.4990 ;
      LAYER M3  ;
        RECT 8.5370 61.4245 8.5550 61.6640 ;
      LAYER V3  ;
        RECT 8.5370 61.4750 8.5550 61.4990 ;
    END
  END dataout[49]
  PIN wd[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 61.3790 8.6650 61.4030 ;
      LAYER M3  ;
        RECT 8.3120 61.3170 8.3300 61.7220 ;
      LAYER V3  ;
        RECT 8.3120 61.3790 8.3300 61.4030 ;
    END
  END wd[49]
  PIN dataout[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 62.5550 8.5970 62.5790 ;
      LAYER M3  ;
        RECT 8.5370 62.5045 8.5550 62.7440 ;
      LAYER V3  ;
        RECT 8.5370 62.5550 8.5550 62.5790 ;
    END
  END dataout[50]
  PIN wd[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 62.4590 8.6650 62.4830 ;
      LAYER M3  ;
        RECT 8.3120 62.3970 8.3300 62.8020 ;
      LAYER V3  ;
        RECT 8.3120 62.4590 8.3300 62.4830 ;
    END
  END wd[50]
  PIN dataout[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 63.6350 8.5970 63.6590 ;
      LAYER M3  ;
        RECT 8.5370 63.5845 8.5550 63.8240 ;
      LAYER V3  ;
        RECT 8.5370 63.6350 8.5550 63.6590 ;
    END
  END dataout[51]
  PIN wd[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 63.5390 8.6650 63.5630 ;
      LAYER M3  ;
        RECT 8.3120 63.4770 8.3300 63.8820 ;
      LAYER V3  ;
        RECT 8.3120 63.5390 8.3300 63.5630 ;
    END
  END wd[51]
  PIN dataout[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 64.7150 8.5970 64.7390 ;
      LAYER M3  ;
        RECT 8.5370 64.6645 8.5550 64.9040 ;
      LAYER V3  ;
        RECT 8.5370 64.7150 8.5550 64.7390 ;
    END
  END dataout[52]
  PIN wd[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 64.6190 8.6650 64.6430 ;
      LAYER M3  ;
        RECT 8.3120 64.5570 8.3300 64.9620 ;
      LAYER V3  ;
        RECT 8.3120 64.6190 8.3300 64.6430 ;
    END
  END wd[52]
  PIN dataout[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 65.7950 8.5970 65.8190 ;
      LAYER M3  ;
        RECT 8.5370 65.7445 8.5550 65.9840 ;
      LAYER V3  ;
        RECT 8.5370 65.7950 8.5550 65.8190 ;
    END
  END dataout[53]
  PIN wd[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 65.6990 8.6650 65.7230 ;
      LAYER M3  ;
        RECT 8.3120 65.6370 8.3300 66.0420 ;
      LAYER V3  ;
        RECT 8.3120 65.6990 8.3300 65.7230 ;
    END
  END wd[53]
  PIN dataout[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 66.8750 8.5970 66.8990 ;
      LAYER M3  ;
        RECT 8.5370 66.8245 8.5550 67.0640 ;
      LAYER V3  ;
        RECT 8.5370 66.8750 8.5550 66.8990 ;
    END
  END dataout[54]
  PIN wd[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 66.7790 8.6650 66.8030 ;
      LAYER M3  ;
        RECT 8.3120 66.7170 8.3300 67.1220 ;
      LAYER V3  ;
        RECT 8.3120 66.7790 8.3300 66.8030 ;
    END
  END wd[54]
  PIN dataout[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 67.9550 8.5970 67.9790 ;
      LAYER M3  ;
        RECT 8.5370 67.9045 8.5550 68.1440 ;
      LAYER V3  ;
        RECT 8.5370 67.9550 8.5550 67.9790 ;
    END
  END dataout[55]
  PIN wd[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 67.8590 8.6650 67.8830 ;
      LAYER M3  ;
        RECT 8.3120 67.7970 8.3300 68.2020 ;
      LAYER V3  ;
        RECT 8.3120 67.8590 8.3300 67.8830 ;
    END
  END wd[55]
  PIN dataout[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 69.0350 8.5970 69.0590 ;
      LAYER M3  ;
        RECT 8.5370 68.9845 8.5550 69.2240 ;
      LAYER V3  ;
        RECT 8.5370 69.0350 8.5550 69.0590 ;
    END
  END dataout[56]
  PIN wd[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 68.9390 8.6650 68.9630 ;
      LAYER M3  ;
        RECT 8.3120 68.8770 8.3300 69.2820 ;
      LAYER V3  ;
        RECT 8.3120 68.9390 8.3300 68.9630 ;
    END
  END wd[56]
  PIN dataout[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 70.1150 8.5970 70.1390 ;
      LAYER M3  ;
        RECT 8.5370 70.0645 8.5550 70.3040 ;
      LAYER V3  ;
        RECT 8.5370 70.1150 8.5550 70.1390 ;
    END
  END dataout[57]
  PIN wd[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 70.0190 8.6650 70.0430 ;
      LAYER M3  ;
        RECT 8.3120 69.9570 8.3300 70.3620 ;
      LAYER V3  ;
        RECT 8.3120 70.0190 8.3300 70.0430 ;
    END
  END wd[57]
  PIN dataout[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 71.1950 8.5970 71.2190 ;
      LAYER M3  ;
        RECT 8.5370 71.1445 8.5550 71.3840 ;
      LAYER V3  ;
        RECT 8.5370 71.1950 8.5550 71.2190 ;
    END
  END dataout[58]
  PIN wd[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 71.0990 8.6650 71.1230 ;
      LAYER M3  ;
        RECT 8.3120 71.0370 8.3300 71.4420 ;
      LAYER V3  ;
        RECT 8.3120 71.0990 8.3300 71.1230 ;
    END
  END wd[58]
  PIN dataout[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 72.2750 8.5970 72.2990 ;
      LAYER M3  ;
        RECT 8.5370 72.2245 8.5550 72.4640 ;
      LAYER V3  ;
        RECT 8.5370 72.2750 8.5550 72.2990 ;
    END
  END dataout[59]
  PIN wd[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 72.1790 8.6650 72.2030 ;
      LAYER M3  ;
        RECT 8.3120 72.1170 8.3300 72.5220 ;
      LAYER V3  ;
        RECT 8.3120 72.1790 8.3300 72.2030 ;
    END
  END wd[59]
  PIN dataout[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 73.3550 8.5970 73.3790 ;
      LAYER M3  ;
        RECT 8.5370 73.3045 8.5550 73.5440 ;
      LAYER V3  ;
        RECT 8.5370 73.3550 8.5550 73.3790 ;
    END
  END dataout[60]
  PIN wd[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 73.2590 8.6650 73.2830 ;
      LAYER M3  ;
        RECT 8.3120 73.1970 8.3300 73.6020 ;
      LAYER V3  ;
        RECT 8.3120 73.2590 8.3300 73.2830 ;
    END
  END wd[60]
  PIN dataout[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 74.4350 8.5970 74.4590 ;
      LAYER M3  ;
        RECT 8.5370 74.3845 8.5550 74.6240 ;
      LAYER V3  ;
        RECT 8.5370 74.4350 8.5550 74.4590 ;
    END
  END dataout[61]
  PIN wd[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 74.3390 8.6650 74.3630 ;
      LAYER M3  ;
        RECT 8.3120 74.2770 8.3300 74.6820 ;
      LAYER V3  ;
        RECT 8.3120 74.3390 8.3300 74.3630 ;
    END
  END wd[61]
  PIN dataout[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 75.5150 8.5970 75.5390 ;
      LAYER M3  ;
        RECT 8.5370 75.4645 8.5550 75.7040 ;
      LAYER V3  ;
        RECT 8.5370 75.5150 8.5550 75.5390 ;
    END
  END dataout[62]
  PIN wd[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 75.4190 8.6650 75.4430 ;
      LAYER M3  ;
        RECT 8.3120 75.3570 8.3300 75.7620 ;
      LAYER V3  ;
        RECT 8.3120 75.4190 8.3300 75.4430 ;
    END
  END wd[62]
  PIN dataout[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 76.5950 8.5970 76.6190 ;
      LAYER M3  ;
        RECT 8.5370 76.5445 8.5550 76.7840 ;
      LAYER V3  ;
        RECT 8.5370 76.5950 8.5550 76.6190 ;
    END
  END dataout[63]
  PIN wd[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 76.4990 8.6650 76.5230 ;
      LAYER M3  ;
        RECT 8.3120 76.4370 8.3300 76.8420 ;
      LAYER V3  ;
        RECT 8.3120 76.4990 8.3300 76.5230 ;
    END
  END wd[63]
  PIN dataout[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 77.6750 8.5970 77.6990 ;
      LAYER M3  ;
        RECT 8.5370 77.6245 8.5550 77.8640 ;
      LAYER V3  ;
        RECT 8.5370 77.6750 8.5550 77.6990 ;
    END
  END dataout[64]
  PIN wd[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 77.5790 8.6650 77.6030 ;
      LAYER M3  ;
        RECT 8.3120 77.5170 8.3300 77.9220 ;
      LAYER V3  ;
        RECT 8.3120 77.5790 8.3300 77.6030 ;
    END
  END wd[64]
  PIN dataout[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 78.7550 8.5970 78.7790 ;
      LAYER M3  ;
        RECT 8.5370 78.7045 8.5550 78.9440 ;
      LAYER V3  ;
        RECT 8.5370 78.7550 8.5550 78.7790 ;
    END
  END dataout[65]
  PIN wd[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 78.6590 8.6650 78.6830 ;
      LAYER M3  ;
        RECT 8.3120 78.5970 8.3300 79.0020 ;
      LAYER V3  ;
        RECT 8.3120 78.6590 8.3300 78.6830 ;
    END
  END wd[65]
  PIN dataout[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 79.8350 8.5970 79.8590 ;
      LAYER M3  ;
        RECT 8.5370 79.7845 8.5550 80.0240 ;
      LAYER V3  ;
        RECT 8.5370 79.8350 8.5550 79.8590 ;
    END
  END dataout[66]
  PIN wd[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 79.7390 8.6650 79.7630 ;
      LAYER M3  ;
        RECT 8.3120 79.6770 8.3300 80.0820 ;
      LAYER V3  ;
        RECT 8.3120 79.7390 8.3300 79.7630 ;
    END
  END wd[66]
  PIN dataout[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 80.9150 8.5970 80.9390 ;
      LAYER M3  ;
        RECT 8.5370 80.8645 8.5550 81.1040 ;
      LAYER V3  ;
        RECT 8.5370 80.9150 8.5550 80.9390 ;
    END
  END dataout[67]
  PIN wd[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 80.8190 8.6650 80.8430 ;
      LAYER M3  ;
        RECT 8.3120 80.7570 8.3300 81.1620 ;
      LAYER V3  ;
        RECT 8.3120 80.8190 8.3300 80.8430 ;
    END
  END wd[67]
  PIN dataout[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 81.9950 8.5970 82.0190 ;
      LAYER M3  ;
        RECT 8.5370 81.9445 8.5550 82.1840 ;
      LAYER V3  ;
        RECT 8.5370 81.9950 8.5550 82.0190 ;
    END
  END dataout[68]
  PIN wd[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 81.8990 8.6650 81.9230 ;
      LAYER M3  ;
        RECT 8.3120 81.8370 8.3300 82.2420 ;
      LAYER V3  ;
        RECT 8.3120 81.8990 8.3300 81.9230 ;
    END
  END wd[68]
  PIN dataout[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 83.0750 8.5970 83.0990 ;
      LAYER M3  ;
        RECT 8.5370 83.0245 8.5550 83.2640 ;
      LAYER V3  ;
        RECT 8.5370 83.0750 8.5550 83.0990 ;
    END
  END dataout[69]
  PIN wd[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 82.9790 8.6650 83.0030 ;
      LAYER M3  ;
        RECT 8.3120 82.9170 8.3300 83.3220 ;
      LAYER V3  ;
        RECT 8.3120 82.9790 8.3300 83.0030 ;
    END
  END wd[69]
  PIN dataout[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 84.1550 8.5970 84.1790 ;
      LAYER M3  ;
        RECT 8.5370 84.1045 8.5550 84.3440 ;
      LAYER V3  ;
        RECT 8.5370 84.1550 8.5550 84.1790 ;
    END
  END dataout[70]
  PIN wd[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 84.0590 8.6650 84.0830 ;
      LAYER M3  ;
        RECT 8.3120 83.9970 8.3300 84.4020 ;
      LAYER V3  ;
        RECT 8.3120 84.0590 8.3300 84.0830 ;
    END
  END wd[70]
  PIN dataout[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 85.2350 8.5970 85.2590 ;
      LAYER M3  ;
        RECT 8.5370 85.1845 8.5550 85.4240 ;
      LAYER V3  ;
        RECT 8.5370 85.2350 8.5550 85.2590 ;
    END
  END dataout[71]
  PIN wd[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 85.1390 8.6650 85.1630 ;
      LAYER M3  ;
        RECT 8.3120 85.0770 8.3300 85.4820 ;
      LAYER V3  ;
        RECT 8.3120 85.1390 8.3300 85.1630 ;
    END
  END wd[71]
  PIN dataout[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 86.3150 8.5970 86.3390 ;
      LAYER M3  ;
        RECT 8.5370 86.2645 8.5550 86.5040 ;
      LAYER V3  ;
        RECT 8.5370 86.3150 8.5550 86.3390 ;
    END
  END dataout[72]
  PIN wd[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 86.2190 8.6650 86.2430 ;
      LAYER M3  ;
        RECT 8.3120 86.1570 8.3300 86.5620 ;
      LAYER V3  ;
        RECT 8.3120 86.2190 8.3300 86.2430 ;
    END
  END wd[72]
  PIN dataout[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 87.3950 8.5970 87.4190 ;
      LAYER M3  ;
        RECT 8.5370 87.3445 8.5550 87.5840 ;
      LAYER V3  ;
        RECT 8.5370 87.3950 8.5550 87.4190 ;
    END
  END dataout[73]
  PIN wd[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 87.2990 8.6650 87.3230 ;
      LAYER M3  ;
        RECT 8.3120 87.2370 8.3300 87.6420 ;
      LAYER V3  ;
        RECT 8.3120 87.2990 8.3300 87.3230 ;
    END
  END wd[73]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0050 26.1765 16.5290 27.2700 ;
      RECT 0.0050 27.2565 16.5290 28.3500 ;
      RECT 0.0050 28.3365 16.5290 29.4300 ;
      RECT 0.0050 29.4165 16.5290 30.5100 ;
      RECT 0.0050 30.4965 16.5290 31.5900 ;
      RECT 0.0050 31.5765 16.5290 32.6700 ;
      RECT 0.0050 32.6565 16.5290 33.7500 ;
      RECT 0.0050 33.7365 16.5290 34.8300 ;
      RECT 0.0050 34.8165 16.5290 35.9100 ;
      RECT 0.0050 35.8965 16.5290 36.9900 ;
      RECT 0.0050 36.9765 16.5290 38.0700 ;
      RECT 0.0050 38.0565 16.5290 39.1500 ;
      RECT 0.0050 39.1365 16.5290 40.2300 ;
      RECT 0.0000 40.1970 16.5240 48.8505 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
        RECT 0.0050 60.2235 16.5290 61.3170 ;
        RECT 0.0050 61.3035 16.5290 62.3970 ;
        RECT 0.0050 62.3835 16.5290 63.4770 ;
        RECT 0.0050 63.4635 16.5290 64.5570 ;
        RECT 0.0050 64.5435 16.5290 65.6370 ;
        RECT 0.0050 65.6235 16.5290 66.7170 ;
        RECT 0.0050 66.7035 16.5290 67.7970 ;
        RECT 0.0050 67.7835 16.5290 68.8770 ;
        RECT 0.0050 68.8635 16.5290 69.9570 ;
        RECT 0.0050 69.9435 16.5290 71.0370 ;
        RECT 0.0050 71.0235 16.5290 72.1170 ;
        RECT 0.0050 72.1035 16.5290 73.1970 ;
        RECT 0.0050 73.1835 16.5290 74.2770 ;
        RECT 0.0050 74.2635 16.5290 75.3570 ;
        RECT 0.0050 75.3435 16.5290 76.4370 ;
        RECT 0.0050 76.4235 16.5290 77.5170 ;
        RECT 0.0050 77.5035 16.5290 78.5970 ;
        RECT 0.0050 78.5835 16.5290 79.6770 ;
        RECT 0.0050 79.6635 16.5290 80.7570 ;
        RECT 0.0050 80.7435 16.5290 81.8370 ;
        RECT 0.0050 81.8235 16.5290 82.9170 ;
        RECT 0.0050 82.9035 16.5290 83.9970 ;
        RECT 0.0050 83.9835 16.5290 85.0770 ;
        RECT 0.0050 85.0635 16.5290 86.1570 ;
        RECT 0.0050 86.1435 16.5290 87.2370 ;
        RECT 0.0050 87.2235 16.5290 88.3170 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0050 26.1765 16.5290 27.2700 ;
      RECT 0.0050 27.2565 16.5290 28.3500 ;
      RECT 0.0050 28.3365 16.5290 29.4300 ;
      RECT 0.0050 29.4165 16.5290 30.5100 ;
      RECT 0.0050 30.4965 16.5290 31.5900 ;
      RECT 0.0050 31.5765 16.5290 32.6700 ;
      RECT 0.0050 32.6565 16.5290 33.7500 ;
      RECT 0.0050 33.7365 16.5290 34.8300 ;
      RECT 0.0050 34.8165 16.5290 35.9100 ;
      RECT 0.0050 35.8965 16.5290 36.9900 ;
      RECT 0.0050 36.9765 16.5290 38.0700 ;
      RECT 0.0050 38.0565 16.5290 39.1500 ;
      RECT 0.0050 39.1365 16.5290 40.2300 ;
      RECT 0.0000 40.1970 16.5240 48.8505 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
        RECT 0.0050 60.2235 16.5290 61.3170 ;
        RECT 0.0050 61.3035 16.5290 62.3970 ;
        RECT 0.0050 62.3835 16.5290 63.4770 ;
        RECT 0.0050 63.4635 16.5290 64.5570 ;
        RECT 0.0050 64.5435 16.5290 65.6370 ;
        RECT 0.0050 65.6235 16.5290 66.7170 ;
        RECT 0.0050 66.7035 16.5290 67.7970 ;
        RECT 0.0050 67.7835 16.5290 68.8770 ;
        RECT 0.0050 68.8635 16.5290 69.9570 ;
        RECT 0.0050 69.9435 16.5290 71.0370 ;
        RECT 0.0050 71.0235 16.5290 72.1170 ;
        RECT 0.0050 72.1035 16.5290 73.1970 ;
        RECT 0.0050 73.1835 16.5290 74.2770 ;
        RECT 0.0050 74.2635 16.5290 75.3570 ;
        RECT 0.0050 75.3435 16.5290 76.4370 ;
        RECT 0.0050 76.4235 16.5290 77.5170 ;
        RECT 0.0050 77.5035 16.5290 78.5970 ;
        RECT 0.0050 78.5835 16.5290 79.6770 ;
        RECT 0.0050 79.6635 16.5290 80.7570 ;
        RECT 0.0050 80.7435 16.5290 81.8370 ;
        RECT 0.0050 81.8235 16.5290 82.9170 ;
        RECT 0.0050 82.9035 16.5290 83.9970 ;
        RECT 0.0050 83.9835 16.5290 85.0770 ;
        RECT 0.0050 85.0635 16.5290 86.1570 ;
        RECT 0.0050 86.1435 16.5290 87.2370 ;
        RECT 0.0050 87.2235 16.5290 88.3170 ;
  LAYER V1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0050 26.1765 16.5290 27.2700 ;
      RECT 0.0050 27.2565 16.5290 28.3500 ;
      RECT 0.0050 28.3365 16.5290 29.4300 ;
      RECT 0.0050 29.4165 16.5290 30.5100 ;
      RECT 0.0050 30.4965 16.5290 31.5900 ;
      RECT 0.0050 31.5765 16.5290 32.6700 ;
      RECT 0.0050 32.6565 16.5290 33.7500 ;
      RECT 0.0050 33.7365 16.5290 34.8300 ;
      RECT 0.0050 34.8165 16.5290 35.9100 ;
      RECT 0.0050 35.8965 16.5290 36.9900 ;
      RECT 0.0050 36.9765 16.5290 38.0700 ;
      RECT 0.0050 38.0565 16.5290 39.1500 ;
      RECT 0.0050 39.1365 16.5290 40.2300 ;
      RECT 0.0000 40.1970 16.5240 48.8505 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
        RECT 0.0050 60.2235 16.5290 61.3170 ;
        RECT 0.0050 61.3035 16.5290 62.3970 ;
        RECT 0.0050 62.3835 16.5290 63.4770 ;
        RECT 0.0050 63.4635 16.5290 64.5570 ;
        RECT 0.0050 64.5435 16.5290 65.6370 ;
        RECT 0.0050 65.6235 16.5290 66.7170 ;
        RECT 0.0050 66.7035 16.5290 67.7970 ;
        RECT 0.0050 67.7835 16.5290 68.8770 ;
        RECT 0.0050 68.8635 16.5290 69.9570 ;
        RECT 0.0050 69.9435 16.5290 71.0370 ;
        RECT 0.0050 71.0235 16.5290 72.1170 ;
        RECT 0.0050 72.1035 16.5290 73.1970 ;
        RECT 0.0050 73.1835 16.5290 74.2770 ;
        RECT 0.0050 74.2635 16.5290 75.3570 ;
        RECT 0.0050 75.3435 16.5290 76.4370 ;
        RECT 0.0050 76.4235 16.5290 77.5170 ;
        RECT 0.0050 77.5035 16.5290 78.5970 ;
        RECT 0.0050 78.5835 16.5290 79.6770 ;
        RECT 0.0050 79.6635 16.5290 80.7570 ;
        RECT 0.0050 80.7435 16.5290 81.8370 ;
        RECT 0.0050 81.8235 16.5290 82.9170 ;
        RECT 0.0050 82.9035 16.5290 83.9970 ;
        RECT 0.0050 83.9835 16.5290 85.0770 ;
        RECT 0.0050 85.0635 16.5290 86.1570 ;
        RECT 0.0050 86.1435 16.5290 87.2370 ;
        RECT 0.0050 87.2235 16.5290 88.3170 ;
  LAYER V2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0050 26.1765 16.5290 27.2700 ;
      RECT 0.0050 27.2565 16.5290 28.3500 ;
      RECT 0.0050 28.3365 16.5290 29.4300 ;
      RECT 0.0050 29.4165 16.5290 30.5100 ;
      RECT 0.0050 30.4965 16.5290 31.5900 ;
      RECT 0.0050 31.5765 16.5290 32.6700 ;
      RECT 0.0050 32.6565 16.5290 33.7500 ;
      RECT 0.0050 33.7365 16.5290 34.8300 ;
      RECT 0.0050 34.8165 16.5290 35.9100 ;
      RECT 0.0050 35.8965 16.5290 36.9900 ;
      RECT 0.0050 36.9765 16.5290 38.0700 ;
      RECT 0.0050 38.0565 16.5290 39.1500 ;
      RECT 0.0050 39.1365 16.5290 40.2300 ;
      RECT 0.0000 40.1970 16.5240 48.8505 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
        RECT 0.0050 60.2235 16.5290 61.3170 ;
        RECT 0.0050 61.3035 16.5290 62.3970 ;
        RECT 0.0050 62.3835 16.5290 63.4770 ;
        RECT 0.0050 63.4635 16.5290 64.5570 ;
        RECT 0.0050 64.5435 16.5290 65.6370 ;
        RECT 0.0050 65.6235 16.5290 66.7170 ;
        RECT 0.0050 66.7035 16.5290 67.7970 ;
        RECT 0.0050 67.7835 16.5290 68.8770 ;
        RECT 0.0050 68.8635 16.5290 69.9570 ;
        RECT 0.0050 69.9435 16.5290 71.0370 ;
        RECT 0.0050 71.0235 16.5290 72.1170 ;
        RECT 0.0050 72.1035 16.5290 73.1970 ;
        RECT 0.0050 73.1835 16.5290 74.2770 ;
        RECT 0.0050 74.2635 16.5290 75.3570 ;
        RECT 0.0050 75.3435 16.5290 76.4370 ;
        RECT 0.0050 76.4235 16.5290 77.5170 ;
        RECT 0.0050 77.5035 16.5290 78.5970 ;
        RECT 0.0050 78.5835 16.5290 79.6770 ;
        RECT 0.0050 79.6635 16.5290 80.7570 ;
        RECT 0.0050 80.7435 16.5290 81.8370 ;
        RECT 0.0050 81.8235 16.5290 82.9170 ;
        RECT 0.0050 82.9035 16.5290 83.9970 ;
        RECT 0.0050 83.9835 16.5290 85.0770 ;
        RECT 0.0050 85.0635 16.5290 86.1570 ;
        RECT 0.0050 86.1435 16.5290 87.2370 ;
        RECT 0.0050 87.2235 16.5290 88.3170 ;
  LAYER M3  ;
      RECT 8.6990 0.3450 8.7170 1.2805 ;
      RECT 8.6630 0.3450 8.6810 1.2805 ;
      RECT 8.6270 0.9220 8.6450 1.2445 ;
      RECT 8.5100 1.1190 8.5280 1.2285 ;
      RECT 8.5010 0.3775 8.5190 0.6170 ;
      RECT 8.4650 0.9585 8.4830 1.1120 ;
      RECT 8.3840 0.9840 8.4020 1.2420 ;
      RECT 7.8440 0.3450 7.8620 1.2805 ;
      RECT 7.8080 0.3450 7.8260 1.2805 ;
      RECT 7.7720 0.5260 7.7900 1.0940 ;
      RECT 8.6990 1.4250 8.7170 2.3605 ;
      RECT 8.6630 1.4250 8.6810 2.3605 ;
      RECT 8.6270 2.0020 8.6450 2.3245 ;
      RECT 8.5100 2.1990 8.5280 2.3085 ;
      RECT 8.5010 1.4575 8.5190 1.6970 ;
      RECT 8.4650 2.0385 8.4830 2.1920 ;
      RECT 8.3840 2.0640 8.4020 2.3220 ;
      RECT 7.8440 1.4250 7.8620 2.3605 ;
      RECT 7.8080 1.4250 7.8260 2.3605 ;
      RECT 7.7720 1.6060 7.7900 2.1740 ;
      RECT 8.6990 2.5050 8.7170 3.4405 ;
      RECT 8.6630 2.5050 8.6810 3.4405 ;
      RECT 8.6270 3.0820 8.6450 3.4045 ;
      RECT 8.5100 3.2790 8.5280 3.3885 ;
      RECT 8.5010 2.5375 8.5190 2.7770 ;
      RECT 8.4650 3.1185 8.4830 3.2720 ;
      RECT 8.3840 3.1440 8.4020 3.4020 ;
      RECT 7.8440 2.5050 7.8620 3.4405 ;
      RECT 7.8080 2.5050 7.8260 3.4405 ;
      RECT 7.7720 2.6860 7.7900 3.2540 ;
      RECT 8.6990 3.5850 8.7170 4.5205 ;
      RECT 8.6630 3.5850 8.6810 4.5205 ;
      RECT 8.6270 4.1620 8.6450 4.4845 ;
      RECT 8.5100 4.3590 8.5280 4.4685 ;
      RECT 8.5010 3.6175 8.5190 3.8570 ;
      RECT 8.4650 4.1985 8.4830 4.3520 ;
      RECT 8.3840 4.2240 8.4020 4.4820 ;
      RECT 7.8440 3.5850 7.8620 4.5205 ;
      RECT 7.8080 3.5850 7.8260 4.5205 ;
      RECT 7.7720 3.7660 7.7900 4.3340 ;
      RECT 8.6990 4.6650 8.7170 5.6005 ;
      RECT 8.6630 4.6650 8.6810 5.6005 ;
      RECT 8.6270 5.2420 8.6450 5.5645 ;
      RECT 8.5100 5.4390 8.5280 5.5485 ;
      RECT 8.5010 4.6975 8.5190 4.9370 ;
      RECT 8.4650 5.2785 8.4830 5.4320 ;
      RECT 8.3840 5.3040 8.4020 5.5620 ;
      RECT 7.8440 4.6650 7.8620 5.6005 ;
      RECT 7.8080 4.6650 7.8260 5.6005 ;
      RECT 7.7720 4.8460 7.7900 5.4140 ;
      RECT 8.6990 5.7450 8.7170 6.6805 ;
      RECT 8.6630 5.7450 8.6810 6.6805 ;
      RECT 8.6270 6.3220 8.6450 6.6445 ;
      RECT 8.5100 6.5190 8.5280 6.6285 ;
      RECT 8.5010 5.7775 8.5190 6.0170 ;
      RECT 8.4650 6.3585 8.4830 6.5120 ;
      RECT 8.3840 6.3840 8.4020 6.6420 ;
      RECT 7.8440 5.7450 7.8620 6.6805 ;
      RECT 7.8080 5.7450 7.8260 6.6805 ;
      RECT 7.7720 5.9260 7.7900 6.4940 ;
      RECT 8.6990 6.8250 8.7170 7.7605 ;
      RECT 8.6630 6.8250 8.6810 7.7605 ;
      RECT 8.6270 7.4020 8.6450 7.7245 ;
      RECT 8.5100 7.5990 8.5280 7.7085 ;
      RECT 8.5010 6.8575 8.5190 7.0970 ;
      RECT 8.4650 7.4385 8.4830 7.5920 ;
      RECT 8.3840 7.4640 8.4020 7.7220 ;
      RECT 7.8440 6.8250 7.8620 7.7605 ;
      RECT 7.8080 6.8250 7.8260 7.7605 ;
      RECT 7.7720 7.0060 7.7900 7.5740 ;
      RECT 8.6990 7.9050 8.7170 8.8405 ;
      RECT 8.6630 7.9050 8.6810 8.8405 ;
      RECT 8.6270 8.4820 8.6450 8.8045 ;
      RECT 8.5100 8.6790 8.5280 8.7885 ;
      RECT 8.5010 7.9375 8.5190 8.1770 ;
      RECT 8.4650 8.5185 8.4830 8.6720 ;
      RECT 8.3840 8.5440 8.4020 8.8020 ;
      RECT 7.8440 7.9050 7.8620 8.8405 ;
      RECT 7.8080 7.9050 7.8260 8.8405 ;
      RECT 7.7720 8.0860 7.7900 8.6540 ;
      RECT 8.6990 8.9850 8.7170 9.9205 ;
      RECT 8.6630 8.9850 8.6810 9.9205 ;
      RECT 8.6270 9.5620 8.6450 9.8845 ;
      RECT 8.5100 9.7590 8.5280 9.8685 ;
      RECT 8.5010 9.0175 8.5190 9.2570 ;
      RECT 8.4650 9.5985 8.4830 9.7520 ;
      RECT 8.3840 9.6240 8.4020 9.8820 ;
      RECT 7.8440 8.9850 7.8620 9.9205 ;
      RECT 7.8080 8.9850 7.8260 9.9205 ;
      RECT 7.7720 9.1660 7.7900 9.7340 ;
      RECT 8.6990 10.0650 8.7170 11.0005 ;
      RECT 8.6630 10.0650 8.6810 11.0005 ;
      RECT 8.6270 10.6420 8.6450 10.9645 ;
      RECT 8.5100 10.8390 8.5280 10.9485 ;
      RECT 8.5010 10.0975 8.5190 10.3370 ;
      RECT 8.4650 10.6785 8.4830 10.8320 ;
      RECT 8.3840 10.7040 8.4020 10.9620 ;
      RECT 7.8440 10.0650 7.8620 11.0005 ;
      RECT 7.8080 10.0650 7.8260 11.0005 ;
      RECT 7.7720 10.2460 7.7900 10.8140 ;
      RECT 8.6990 11.1450 8.7170 12.0805 ;
      RECT 8.6630 11.1450 8.6810 12.0805 ;
      RECT 8.6270 11.7220 8.6450 12.0445 ;
      RECT 8.5100 11.9190 8.5280 12.0285 ;
      RECT 8.5010 11.1775 8.5190 11.4170 ;
      RECT 8.4650 11.7585 8.4830 11.9120 ;
      RECT 8.3840 11.7840 8.4020 12.0420 ;
      RECT 7.8440 11.1450 7.8620 12.0805 ;
      RECT 7.8080 11.1450 7.8260 12.0805 ;
      RECT 7.7720 11.3260 7.7900 11.8940 ;
      RECT 8.6990 12.2250 8.7170 13.1605 ;
      RECT 8.6630 12.2250 8.6810 13.1605 ;
      RECT 8.6270 12.8020 8.6450 13.1245 ;
      RECT 8.5100 12.9990 8.5280 13.1085 ;
      RECT 8.5010 12.2575 8.5190 12.4970 ;
      RECT 8.4650 12.8385 8.4830 12.9920 ;
      RECT 8.3840 12.8640 8.4020 13.1220 ;
      RECT 7.8440 12.2250 7.8620 13.1605 ;
      RECT 7.8080 12.2250 7.8260 13.1605 ;
      RECT 7.7720 12.4060 7.7900 12.9740 ;
      RECT 8.6990 13.3050 8.7170 14.2405 ;
      RECT 8.6630 13.3050 8.6810 14.2405 ;
      RECT 8.6270 13.8820 8.6450 14.2045 ;
      RECT 8.5100 14.0790 8.5280 14.1885 ;
      RECT 8.5010 13.3375 8.5190 13.5770 ;
      RECT 8.4650 13.9185 8.4830 14.0720 ;
      RECT 8.3840 13.9440 8.4020 14.2020 ;
      RECT 7.8440 13.3050 7.8620 14.2405 ;
      RECT 7.8080 13.3050 7.8260 14.2405 ;
      RECT 7.7720 13.4860 7.7900 14.0540 ;
      RECT 8.6990 14.3850 8.7170 15.3205 ;
      RECT 8.6630 14.3850 8.6810 15.3205 ;
      RECT 8.6270 14.9620 8.6450 15.2845 ;
      RECT 8.5100 15.1590 8.5280 15.2685 ;
      RECT 8.5010 14.4175 8.5190 14.6570 ;
      RECT 8.4650 14.9985 8.4830 15.1520 ;
      RECT 8.3840 15.0240 8.4020 15.2820 ;
      RECT 7.8440 14.3850 7.8620 15.3205 ;
      RECT 7.8080 14.3850 7.8260 15.3205 ;
      RECT 7.7720 14.5660 7.7900 15.1340 ;
      RECT 8.6990 15.4650 8.7170 16.4005 ;
      RECT 8.6630 15.4650 8.6810 16.4005 ;
      RECT 8.6270 16.0420 8.6450 16.3645 ;
      RECT 8.5100 16.2390 8.5280 16.3485 ;
      RECT 8.5010 15.4975 8.5190 15.7370 ;
      RECT 8.4650 16.0785 8.4830 16.2320 ;
      RECT 8.3840 16.1040 8.4020 16.3620 ;
      RECT 7.8440 15.4650 7.8620 16.4005 ;
      RECT 7.8080 15.4650 7.8260 16.4005 ;
      RECT 7.7720 15.6460 7.7900 16.2140 ;
      RECT 8.6990 16.5450 8.7170 17.4805 ;
      RECT 8.6630 16.5450 8.6810 17.4805 ;
      RECT 8.6270 17.1220 8.6450 17.4445 ;
      RECT 8.5100 17.3190 8.5280 17.4285 ;
      RECT 8.5010 16.5775 8.5190 16.8170 ;
      RECT 8.4650 17.1585 8.4830 17.3120 ;
      RECT 8.3840 17.1840 8.4020 17.4420 ;
      RECT 7.8440 16.5450 7.8620 17.4805 ;
      RECT 7.8080 16.5450 7.8260 17.4805 ;
      RECT 7.7720 16.7260 7.7900 17.2940 ;
      RECT 8.6990 17.6250 8.7170 18.5605 ;
      RECT 8.6630 17.6250 8.6810 18.5605 ;
      RECT 8.6270 18.2020 8.6450 18.5245 ;
      RECT 8.5100 18.3990 8.5280 18.5085 ;
      RECT 8.5010 17.6575 8.5190 17.8970 ;
      RECT 8.4650 18.2385 8.4830 18.3920 ;
      RECT 8.3840 18.2640 8.4020 18.5220 ;
      RECT 7.8440 17.6250 7.8620 18.5605 ;
      RECT 7.8080 17.6250 7.8260 18.5605 ;
      RECT 7.7720 17.8060 7.7900 18.3740 ;
      RECT 8.6990 18.7050 8.7170 19.6405 ;
      RECT 8.6630 18.7050 8.6810 19.6405 ;
      RECT 8.6270 19.2820 8.6450 19.6045 ;
      RECT 8.5100 19.4790 8.5280 19.5885 ;
      RECT 8.5010 18.7375 8.5190 18.9770 ;
      RECT 8.4650 19.3185 8.4830 19.4720 ;
      RECT 8.3840 19.3440 8.4020 19.6020 ;
      RECT 7.8440 18.7050 7.8620 19.6405 ;
      RECT 7.8080 18.7050 7.8260 19.6405 ;
      RECT 7.7720 18.8860 7.7900 19.4540 ;
      RECT 8.6990 19.7850 8.7170 20.7205 ;
      RECT 8.6630 19.7850 8.6810 20.7205 ;
      RECT 8.6270 20.3620 8.6450 20.6845 ;
      RECT 8.5100 20.5590 8.5280 20.6685 ;
      RECT 8.5010 19.8175 8.5190 20.0570 ;
      RECT 8.4650 20.3985 8.4830 20.5520 ;
      RECT 8.3840 20.4240 8.4020 20.6820 ;
      RECT 7.8440 19.7850 7.8620 20.7205 ;
      RECT 7.8080 19.7850 7.8260 20.7205 ;
      RECT 7.7720 19.9660 7.7900 20.5340 ;
      RECT 8.6990 20.8650 8.7170 21.8005 ;
      RECT 8.6630 20.8650 8.6810 21.8005 ;
      RECT 8.6270 21.4420 8.6450 21.7645 ;
      RECT 8.5100 21.6390 8.5280 21.7485 ;
      RECT 8.5010 20.8975 8.5190 21.1370 ;
      RECT 8.4650 21.4785 8.4830 21.6320 ;
      RECT 8.3840 21.5040 8.4020 21.7620 ;
      RECT 7.8440 20.8650 7.8620 21.8005 ;
      RECT 7.8080 20.8650 7.8260 21.8005 ;
      RECT 7.7720 21.0460 7.7900 21.6140 ;
      RECT 8.6990 21.9450 8.7170 22.8805 ;
      RECT 8.6630 21.9450 8.6810 22.8805 ;
      RECT 8.6270 22.5220 8.6450 22.8445 ;
      RECT 8.5100 22.7190 8.5280 22.8285 ;
      RECT 8.5010 21.9775 8.5190 22.2170 ;
      RECT 8.4650 22.5585 8.4830 22.7120 ;
      RECT 8.3840 22.5840 8.4020 22.8420 ;
      RECT 7.8440 21.9450 7.8620 22.8805 ;
      RECT 7.8080 21.9450 7.8260 22.8805 ;
      RECT 7.7720 22.1260 7.7900 22.6940 ;
      RECT 8.6990 23.0250 8.7170 23.9605 ;
      RECT 8.6630 23.0250 8.6810 23.9605 ;
      RECT 8.6270 23.6020 8.6450 23.9245 ;
      RECT 8.5100 23.7990 8.5280 23.9085 ;
      RECT 8.5010 23.0575 8.5190 23.2970 ;
      RECT 8.4650 23.6385 8.4830 23.7920 ;
      RECT 8.3840 23.6640 8.4020 23.9220 ;
      RECT 7.8440 23.0250 7.8620 23.9605 ;
      RECT 7.8080 23.0250 7.8260 23.9605 ;
      RECT 7.7720 23.2060 7.7900 23.7740 ;
      RECT 8.6990 24.1050 8.7170 25.0405 ;
      RECT 8.6630 24.1050 8.6810 25.0405 ;
      RECT 8.6270 24.6820 8.6450 25.0045 ;
      RECT 8.5100 24.8790 8.5280 24.9885 ;
      RECT 8.5010 24.1375 8.5190 24.3770 ;
      RECT 8.4650 24.7185 8.4830 24.8720 ;
      RECT 8.3840 24.7440 8.4020 25.0020 ;
      RECT 7.8440 24.1050 7.8620 25.0405 ;
      RECT 7.8080 24.1050 7.8260 25.0405 ;
      RECT 7.7720 24.2860 7.7900 24.8540 ;
      RECT 8.6990 25.1850 8.7170 26.1205 ;
      RECT 8.6630 25.1850 8.6810 26.1205 ;
      RECT 8.6270 25.7620 8.6450 26.0845 ;
      RECT 8.5100 25.9590 8.5280 26.0685 ;
      RECT 8.5010 25.2175 8.5190 25.4570 ;
      RECT 8.4650 25.7985 8.4830 25.9520 ;
      RECT 8.3840 25.8240 8.4020 26.0820 ;
      RECT 7.8440 25.1850 7.8620 26.1205 ;
      RECT 7.8080 25.1850 7.8260 26.1205 ;
      RECT 7.7720 25.3660 7.7900 25.9340 ;
      RECT 8.6990 26.2650 8.7170 27.2005 ;
      RECT 8.6630 26.2650 8.6810 27.2005 ;
      RECT 8.6270 26.8420 8.6450 27.1645 ;
      RECT 8.5100 27.0390 8.5280 27.1485 ;
      RECT 8.5010 26.2975 8.5190 26.5370 ;
      RECT 8.4650 26.8785 8.4830 27.0320 ;
      RECT 8.3840 26.9040 8.4020 27.1620 ;
      RECT 7.8440 26.2650 7.8620 27.2005 ;
      RECT 7.8080 26.2650 7.8260 27.2005 ;
      RECT 7.7720 26.4460 7.7900 27.0140 ;
      RECT 8.6990 27.3450 8.7170 28.2805 ;
      RECT 8.6630 27.3450 8.6810 28.2805 ;
      RECT 8.6270 27.9220 8.6450 28.2445 ;
      RECT 8.5100 28.1190 8.5280 28.2285 ;
      RECT 8.5010 27.3775 8.5190 27.6170 ;
      RECT 8.4650 27.9585 8.4830 28.1120 ;
      RECT 8.3840 27.9840 8.4020 28.2420 ;
      RECT 7.8440 27.3450 7.8620 28.2805 ;
      RECT 7.8080 27.3450 7.8260 28.2805 ;
      RECT 7.7720 27.5260 7.7900 28.0940 ;
      RECT 8.6990 28.4250 8.7170 29.3605 ;
      RECT 8.6630 28.4250 8.6810 29.3605 ;
      RECT 8.6270 29.0020 8.6450 29.3245 ;
      RECT 8.5100 29.1990 8.5280 29.3085 ;
      RECT 8.5010 28.4575 8.5190 28.6970 ;
      RECT 8.4650 29.0385 8.4830 29.1920 ;
      RECT 8.3840 29.0640 8.4020 29.3220 ;
      RECT 7.8440 28.4250 7.8620 29.3605 ;
      RECT 7.8080 28.4250 7.8260 29.3605 ;
      RECT 7.7720 28.6060 7.7900 29.1740 ;
      RECT 8.6990 29.5050 8.7170 30.4405 ;
      RECT 8.6630 29.5050 8.6810 30.4405 ;
      RECT 8.6270 30.0820 8.6450 30.4045 ;
      RECT 8.5100 30.2790 8.5280 30.3885 ;
      RECT 8.5010 29.5375 8.5190 29.7770 ;
      RECT 8.4650 30.1185 8.4830 30.2720 ;
      RECT 8.3840 30.1440 8.4020 30.4020 ;
      RECT 7.8440 29.5050 7.8620 30.4405 ;
      RECT 7.8080 29.5050 7.8260 30.4405 ;
      RECT 7.7720 29.6860 7.7900 30.2540 ;
      RECT 8.6990 30.5850 8.7170 31.5205 ;
      RECT 8.6630 30.5850 8.6810 31.5205 ;
      RECT 8.6270 31.1620 8.6450 31.4845 ;
      RECT 8.5100 31.3590 8.5280 31.4685 ;
      RECT 8.5010 30.6175 8.5190 30.8570 ;
      RECT 8.4650 31.1985 8.4830 31.3520 ;
      RECT 8.3840 31.2240 8.4020 31.4820 ;
      RECT 7.8440 30.5850 7.8620 31.5205 ;
      RECT 7.8080 30.5850 7.8260 31.5205 ;
      RECT 7.7720 30.7660 7.7900 31.3340 ;
      RECT 8.6990 31.6650 8.7170 32.6005 ;
      RECT 8.6630 31.6650 8.6810 32.6005 ;
      RECT 8.6270 32.2420 8.6450 32.5645 ;
      RECT 8.5100 32.4390 8.5280 32.5485 ;
      RECT 8.5010 31.6975 8.5190 31.9370 ;
      RECT 8.4650 32.2785 8.4830 32.4320 ;
      RECT 8.3840 32.3040 8.4020 32.5620 ;
      RECT 7.8440 31.6650 7.8620 32.6005 ;
      RECT 7.8080 31.6650 7.8260 32.6005 ;
      RECT 7.7720 31.8460 7.7900 32.4140 ;
      RECT 8.6990 32.7450 8.7170 33.6805 ;
      RECT 8.6630 32.7450 8.6810 33.6805 ;
      RECT 8.6270 33.3220 8.6450 33.6445 ;
      RECT 8.5100 33.5190 8.5280 33.6285 ;
      RECT 8.5010 32.7775 8.5190 33.0170 ;
      RECT 8.4650 33.3585 8.4830 33.5120 ;
      RECT 8.3840 33.3840 8.4020 33.6420 ;
      RECT 7.8440 32.7450 7.8620 33.6805 ;
      RECT 7.8080 32.7450 7.8260 33.6805 ;
      RECT 7.7720 32.9260 7.7900 33.4940 ;
      RECT 8.6990 33.8250 8.7170 34.7605 ;
      RECT 8.6630 33.8250 8.6810 34.7605 ;
      RECT 8.6270 34.4020 8.6450 34.7245 ;
      RECT 8.5100 34.5990 8.5280 34.7085 ;
      RECT 8.5010 33.8575 8.5190 34.0970 ;
      RECT 8.4650 34.4385 8.4830 34.5920 ;
      RECT 8.3840 34.4640 8.4020 34.7220 ;
      RECT 7.8440 33.8250 7.8620 34.7605 ;
      RECT 7.8080 33.8250 7.8260 34.7605 ;
      RECT 7.7720 34.0060 7.7900 34.5740 ;
      RECT 8.6990 34.9050 8.7170 35.8405 ;
      RECT 8.6630 34.9050 8.6810 35.8405 ;
      RECT 8.6270 35.4820 8.6450 35.8045 ;
      RECT 8.5100 35.6790 8.5280 35.7885 ;
      RECT 8.5010 34.9375 8.5190 35.1770 ;
      RECT 8.4650 35.5185 8.4830 35.6720 ;
      RECT 8.3840 35.5440 8.4020 35.8020 ;
      RECT 7.8440 34.9050 7.8620 35.8405 ;
      RECT 7.8080 34.9050 7.8260 35.8405 ;
      RECT 7.7720 35.0860 7.7900 35.6540 ;
      RECT 8.6990 35.9850 8.7170 36.9205 ;
      RECT 8.6630 35.9850 8.6810 36.9205 ;
      RECT 8.6270 36.5620 8.6450 36.8845 ;
      RECT 8.5100 36.7590 8.5280 36.8685 ;
      RECT 8.5010 36.0175 8.5190 36.2570 ;
      RECT 8.4650 36.5985 8.4830 36.7520 ;
      RECT 8.3840 36.6240 8.4020 36.8820 ;
      RECT 7.8440 35.9850 7.8620 36.9205 ;
      RECT 7.8080 35.9850 7.8260 36.9205 ;
      RECT 7.7720 36.1660 7.7900 36.7340 ;
      RECT 8.6990 37.0650 8.7170 38.0005 ;
      RECT 8.6630 37.0650 8.6810 38.0005 ;
      RECT 8.6270 37.6420 8.6450 37.9645 ;
      RECT 8.5100 37.8390 8.5280 37.9485 ;
      RECT 8.5010 37.0975 8.5190 37.3370 ;
      RECT 8.4650 37.6785 8.4830 37.8320 ;
      RECT 8.3840 37.7040 8.4020 37.9620 ;
      RECT 7.8440 37.0650 7.8620 38.0005 ;
      RECT 7.8080 37.0650 7.8260 38.0005 ;
      RECT 7.7720 37.2460 7.7900 37.8140 ;
      RECT 8.6990 38.1450 8.7170 39.0805 ;
      RECT 8.6630 38.1450 8.6810 39.0805 ;
      RECT 8.6270 38.7220 8.6450 39.0445 ;
      RECT 8.5100 38.9190 8.5280 39.0285 ;
      RECT 8.5010 38.1775 8.5190 38.4170 ;
      RECT 8.4650 38.7585 8.4830 38.9120 ;
      RECT 8.3840 38.7840 8.4020 39.0420 ;
      RECT 7.8440 38.1450 7.8620 39.0805 ;
      RECT 7.8080 38.1450 7.8260 39.0805 ;
      RECT 7.7720 38.3260 7.7900 38.8940 ;
      RECT 8.6990 39.2250 8.7170 40.1605 ;
      RECT 8.6630 39.2250 8.6810 40.1605 ;
      RECT 8.6270 39.8020 8.6450 40.1245 ;
      RECT 8.5100 39.9990 8.5280 40.1085 ;
      RECT 8.5010 39.2575 8.5190 39.4970 ;
      RECT 8.4650 39.8385 8.4830 39.9920 ;
      RECT 8.3840 39.8640 8.4020 40.1220 ;
      RECT 7.8440 39.2250 7.8620 40.1605 ;
      RECT 7.8080 39.2250 7.8260 40.1605 ;
      RECT 7.7720 39.4060 7.7900 39.9740 ;
      RECT 16.3170 43.9900 16.3350 48.3440 ;
      RECT 16.2810 42.6750 16.2990 42.7440 ;
      RECT 16.2810 44.2950 16.2990 44.3780 ;
      RECT 16.2450 40.1705 16.2630 48.3775 ;
      RECT 16.2090 44.0225 16.2270 44.7125 ;
      RECT 16.2090 44.7635 16.2270 45.7500 ;
      RECT 16.2090 45.7900 16.2270 46.4070 ;
      RECT 16.1730 43.9590 16.1910 44.6637 ;
      RECT 16.1730 45.4170 16.1910 46.5870 ;
      RECT 16.1370 40.1705 16.1550 43.7670 ;
      RECT 16.0290 40.1705 16.0470 43.7670 ;
      RECT 15.9210 40.1705 15.9390 43.7670 ;
      RECT 15.8130 40.1705 15.8310 43.7670 ;
      RECT 15.7050 40.1705 15.7230 43.7670 ;
      RECT 15.5970 40.1705 15.6150 43.7670 ;
      RECT 15.4890 40.1705 15.5070 43.7670 ;
      RECT 15.3810 40.1705 15.3990 43.7670 ;
      RECT 15.2730 40.1705 15.2910 43.7670 ;
      RECT 15.1650 40.1705 15.1830 43.7670 ;
      RECT 15.0570 40.1705 15.0750 43.7670 ;
      RECT 14.9490 40.1705 14.9670 43.7670 ;
      RECT 14.8410 40.1705 14.8590 43.7670 ;
      RECT 14.7330 40.1705 14.7510 43.7670 ;
      RECT 14.6250 40.1705 14.6430 43.7670 ;
      RECT 14.5170 40.1705 14.5350 43.7670 ;
      RECT 14.4090 40.1705 14.4270 43.7670 ;
      RECT 14.3010 40.1705 14.3190 43.7670 ;
      RECT 14.1930 40.1705 14.2110 43.7670 ;
      RECT 14.0850 40.1705 14.1030 43.7670 ;
      RECT 13.9770 40.1705 13.9950 43.7670 ;
      RECT 13.8690 40.1705 13.8870 43.7670 ;
      RECT 13.7610 40.1705 13.7790 43.7670 ;
      RECT 13.6530 40.1705 13.6710 43.7670 ;
      RECT 13.5450 40.1705 13.5630 43.7670 ;
      RECT 13.4370 40.1705 13.4550 43.7670 ;
      RECT 13.3290 40.1705 13.3470 43.7670 ;
      RECT 13.2210 40.1705 13.2390 43.7670 ;
      RECT 13.1130 40.1705 13.1310 43.7670 ;
      RECT 13.0050 40.1705 13.0230 43.7670 ;
      RECT 12.8970 40.1705 12.9150 43.7670 ;
      RECT 12.7890 40.1705 12.8070 43.7670 ;
      RECT 12.6810 40.1705 12.6990 43.7670 ;
      RECT 12.5730 40.1705 12.5910 43.7670 ;
      RECT 12.4650 40.1705 12.4830 43.7670 ;
      RECT 12.3570 40.1705 12.3750 43.7670 ;
      RECT 12.2490 40.1705 12.2670 43.7670 ;
      RECT 12.1410 40.1705 12.1590 43.7670 ;
      RECT 12.0330 40.1705 12.0510 43.7670 ;
      RECT 11.9250 40.1705 11.9430 43.7670 ;
      RECT 11.8170 40.1705 11.8350 43.7670 ;
      RECT 11.7090 40.1705 11.7270 43.7670 ;
      RECT 11.6010 40.1705 11.6190 43.7670 ;
      RECT 11.4930 40.1705 11.5110 43.7670 ;
      RECT 11.3850 40.1705 11.4030 43.7670 ;
      RECT 11.2770 40.1705 11.2950 43.7670 ;
      RECT 11.1690 40.1705 11.1870 43.7670 ;
      RECT 11.0610 40.1705 11.0790 43.7670 ;
      RECT 10.9530 40.1705 10.9710 43.7670 ;
      RECT 10.8450 40.1705 10.8630 43.7670 ;
      RECT 10.7370 40.1705 10.7550 43.7670 ;
      RECT 10.6290 40.1705 10.6470 43.7670 ;
      RECT 10.5210 40.1705 10.5390 43.7670 ;
      RECT 10.4130 40.1705 10.4310 43.7670 ;
      RECT 10.3050 40.1705 10.3230 43.7670 ;
      RECT 10.1970 40.1705 10.2150 43.7670 ;
      RECT 10.0890 40.1705 10.1070 43.7670 ;
      RECT 9.9810 40.1705 9.9990 43.7670 ;
      RECT 9.8730 40.1705 9.8910 43.7670 ;
      RECT 9.7650 40.1705 9.7830 43.7670 ;
      RECT 9.6570 40.1705 9.6750 43.7670 ;
      RECT 9.5490 40.1705 9.5670 43.7670 ;
      RECT 9.5130 44.0255 9.5310 44.6675 ;
      RECT 9.5130 45.3450 9.5310 45.8770 ;
      RECT 9.4950 40.8310 9.5130 41.5070 ;
      RECT 9.4950 42.2530 9.5130 42.5510 ;
      RECT 9.4950 43.3690 9.5130 43.6310 ;
      RECT 9.4770 43.9400 9.4950 44.7125 ;
      RECT 9.4770 44.7637 9.4950 45.2550 ;
      RECT 9.4770 45.3000 9.4950 45.6710 ;
      RECT 9.4770 45.7470 9.4950 46.4070 ;
      RECT 9.4410 40.1705 9.4590 48.3775 ;
      RECT 9.4050 44.4830 9.4230 44.9475 ;
      RECT 9.3870 40.9390 9.4050 41.5700 ;
      RECT 9.3870 41.9830 9.4050 42.1730 ;
      RECT 9.3870 42.8650 9.4050 42.9140 ;
      RECT 9.3870 43.5970 9.4050 43.6340 ;
      RECT 9.3690 43.9900 9.3870 48.3395 ;
      RECT 9.2790 40.5610 9.2970 41.3630 ;
      RECT 9.2790 41.9110 9.2970 42.4790 ;
      RECT 9.2430 41.9830 9.2610 42.3530 ;
      RECT 9.2070 41.3350 9.2250 41.4710 ;
      RECT 9.2070 42.3250 9.2250 42.5510 ;
      RECT 9.2070 43.5670 9.2250 43.6310 ;
      RECT 9.1710 41.4370 9.1890 41.4740 ;
      RECT 9.1710 43.0630 9.1890 43.1060 ;
      RECT 9.1710 43.5970 9.1890 43.6340 ;
      RECT 9.1350 41.7490 9.1530 42.2450 ;
      RECT 9.1350 42.2890 9.1530 42.4790 ;
      RECT 9.1350 43.2490 9.1530 43.5590 ;
      RECT 9.0990 41.6410 9.1170 42.8880 ;
      RECT 9.0990 45.5290 9.1170 46.2590 ;
      RECT 9.0990 46.6090 9.1170 47.3390 ;
      RECT 8.7750 41.3710 8.7930 41.6690 ;
      RECT 8.7750 42.5590 8.7930 42.6230 ;
      RECT 8.7750 42.8290 8.7930 43.2890 ;
      RECT 8.7750 44.0290 8.7930 44.0660 ;
      RECT 8.7750 46.0690 8.7930 46.3670 ;
      RECT 8.7390 41.4430 8.7570 41.9480 ;
      RECT 8.7390 42.2170 8.7570 43.0190 ;
      RECT 8.7390 44.0620 8.7570 44.3330 ;
      RECT 8.7390 44.4130 8.7570 44.6390 ;
      RECT 8.7030 41.3710 8.7210 42.0470 ;
      RECT 8.7030 42.1450 8.7210 42.4790 ;
      RECT 8.7030 42.6850 8.7210 42.8210 ;
      RECT 8.7030 43.3690 8.7210 44.1710 ;
      RECT 8.7030 44.6050 8.7210 44.6420 ;
      RECT 8.7030 46.7710 8.7210 47.1050 ;
      RECT 8.6670 41.6050 8.6850 41.7410 ;
      RECT 8.6670 43.4950 8.6850 44.4770 ;
      RECT 8.6670 44.9170 8.6850 45.2150 ;
      RECT 8.6670 46.6090 8.6850 46.8710 ;
      RECT 8.6310 40.6690 8.6490 40.8230 ;
      RECT 8.6310 41.4790 8.6490 43.2650 ;
      RECT 8.6310 44.3050 8.6490 46.6370 ;
      RECT 8.6310 46.8430 8.6490 47.9510 ;
      RECT 8.3430 40.9390 8.3610 41.2010 ;
      RECT 8.3430 41.3350 8.3610 41.3990 ;
      RECT 8.3430 41.4790 8.3610 41.7050 ;
      RECT 8.3430 41.7490 8.3610 41.9390 ;
      RECT 8.3430 42.0190 8.3610 44.6390 ;
      RECT 8.3430 44.6830 8.3610 45.9890 ;
      RECT 8.3430 47.0770 8.3610 47.3390 ;
      RECT 8.3070 41.9380 8.3250 42.2090 ;
      RECT 8.3070 42.2890 8.3250 43.1270 ;
      RECT 8.3070 43.2970 8.3250 44.1350 ;
      RECT 8.3070 44.1790 8.3250 45.4490 ;
      RECT 8.3070 45.6550 8.3250 45.8270 ;
      RECT 8.3070 46.5370 8.3250 47.6090 ;
      RECT 8.2710 42.0190 8.2890 42.2900 ;
      RECT 8.2710 42.4450 8.2890 42.4820 ;
      RECT 8.2710 43.2250 8.2890 44.2070 ;
      RECT 8.2710 44.4490 8.2890 44.9090 ;
      RECT 8.2710 45.2590 8.2890 45.9980 ;
      RECT 8.2350 41.1370 8.2530 42.2090 ;
      RECT 8.2350 43.8010 8.2530 44.0180 ;
      RECT 8.2350 45.1870 8.2530 45.4850 ;
      RECT 8.1990 41.7850 8.2170 42.2450 ;
      RECT 8.1990 43.3690 8.2170 43.5590 ;
      RECT 8.1990 43.6000 8.2170 43.6370 ;
      RECT 8.1990 43.8730 8.2170 44.2070 ;
      RECT 8.1990 44.3410 8.2170 45.6830 ;
      RECT 8.1990 45.7900 8.2170 46.9070 ;
      RECT 8.1630 41.2090 8.1810 41.3990 ;
      RECT 8.1630 41.6050 8.1810 41.7410 ;
      RECT 8.1630 42.0190 8.1810 45.1790 ;
      RECT 8.1630 45.2590 8.1810 45.7190 ;
      RECT 8.1630 46.3390 8.1810 46.7990 ;
      RECT 8.1630 47.6530 8.1810 47.8790 ;
      RECT 8.1270 40.1970 8.1450 40.3510 ;
      RECT 8.1270 48.1920 8.1450 48.3580 ;
      RECT 8.0910 40.1970 8.1090 40.2470 ;
      RECT 8.0190 40.1970 8.0370 40.2685 ;
      RECT 8.0190 48.2615 8.0370 48.3775 ;
      RECT 7.8750 41.7130 7.8930 41.9030 ;
      RECT 7.8750 42.4510 7.8930 42.8210 ;
      RECT 7.8750 44.4130 7.8930 44.6390 ;
      RECT 7.8750 44.9530 7.8930 46.0970 ;
      RECT 7.8750 46.8790 7.8930 47.3390 ;
      RECT 7.8750 47.9170 7.8930 47.9540 ;
      RECT 7.8390 40.6690 7.8570 41.1650 ;
      RECT 7.8390 44.7490 7.8570 44.7860 ;
      RECT 7.8390 45.8260 7.8570 46.6370 ;
      RECT 7.8030 41.1370 7.8210 41.3990 ;
      RECT 7.8030 41.6770 7.8210 42.0110 ;
      RECT 7.8030 42.2170 7.8210 42.3170 ;
      RECT 7.8030 43.0990 7.8210 45.8630 ;
      RECT 7.8030 45.9970 7.8210 46.2230 ;
      RECT 7.7670 40.7950 7.7850 41.9390 ;
      RECT 7.7670 45.5290 7.7850 45.7190 ;
      RECT 7.7670 46.3330 7.7850 46.3700 ;
      RECT 7.7670 46.6090 7.7850 47.4110 ;
      RECT 7.7310 41.7490 7.7490 42.7490 ;
      RECT 7.7310 46.1890 7.7490 46.2260 ;
      RECT 7.3710 41.3350 7.3890 41.7410 ;
      RECT 7.2990 41.3710 7.3170 41.9750 ;
      RECT 7.2630 41.2090 7.2810 41.2730 ;
      RECT 7.2270 40.2500 7.2450 40.3010 ;
      RECT 7.2270 43.3690 7.2450 43.5590 ;
      RECT 7.2090 43.9900 7.2270 48.3385 ;
      RECT 7.1370 43.9900 7.1550 48.3395 ;
      RECT 7.1190 40.6690 7.1370 40.8590 ;
      RECT 7.1190 41.4430 7.1370 43.7030 ;
      RECT 7.1010 44.4830 7.1190 44.9475 ;
      RECT 7.0650 40.1705 7.0830 48.3775 ;
      RECT 7.0290 43.9400 7.0470 44.7125 ;
      RECT 7.0290 44.7637 7.0470 45.2550 ;
      RECT 7.0290 45.3000 7.0470 45.6710 ;
      RECT 7.0290 45.7470 7.0470 46.4070 ;
      RECT 7.0110 40.6690 7.0290 41.1650 ;
      RECT 7.0110 41.9470 7.0290 42.5150 ;
      RECT 7.0110 42.8290 7.0290 43.5590 ;
      RECT 6.9930 44.0255 7.0110 44.6675 ;
      RECT 6.9930 45.3450 7.0110 45.8770 ;
      RECT 6.9570 40.1705 6.9750 43.7670 ;
      RECT 6.8490 40.1705 6.8670 43.7670 ;
      RECT 6.7410 40.1705 6.7590 43.7670 ;
      RECT 6.6330 40.1705 6.6510 43.7670 ;
      RECT 6.5250 40.1705 6.5430 43.7670 ;
      RECT 6.4170 40.1705 6.4350 43.7670 ;
      RECT 6.3090 40.1705 6.3270 43.7670 ;
      RECT 6.2010 40.1705 6.2190 43.7670 ;
      RECT 6.0930 40.1705 6.1110 43.7670 ;
      RECT 5.9850 40.1705 6.0030 43.7670 ;
      RECT 5.8770 40.1705 5.8950 43.7670 ;
      RECT 5.7690 40.1705 5.7870 43.7670 ;
      RECT 5.6610 40.1705 5.6790 43.7670 ;
      RECT 5.5530 40.1705 5.5710 43.7670 ;
      RECT 5.4450 40.1705 5.4630 43.7670 ;
      RECT 5.3370 40.1705 5.3550 43.7670 ;
      RECT 5.2290 40.1705 5.2470 43.7670 ;
      RECT 5.1210 40.1705 5.1390 43.7670 ;
      RECT 5.0130 40.1705 5.0310 43.7670 ;
      RECT 4.9050 40.1705 4.9230 43.7670 ;
      RECT 4.7970 40.1705 4.8150 43.7670 ;
      RECT 4.6890 40.1705 4.7070 43.7670 ;
      RECT 4.5810 40.1705 4.5990 43.7670 ;
      RECT 4.4730 40.1705 4.4910 43.7670 ;
      RECT 4.3650 40.1705 4.3830 43.7670 ;
      RECT 4.2570 40.1705 4.2750 43.7670 ;
      RECT 4.1490 40.1705 4.1670 43.7670 ;
      RECT 4.0410 40.1705 4.0590 43.7670 ;
      RECT 3.9330 40.1705 3.9510 43.7670 ;
      RECT 3.8250 40.1705 3.8430 43.7670 ;
      RECT 3.7170 40.1705 3.7350 43.7670 ;
      RECT 3.6090 40.1705 3.6270 43.7670 ;
      RECT 3.5010 40.1705 3.5190 43.7670 ;
      RECT 3.3930 40.1705 3.4110 43.7670 ;
      RECT 3.2850 40.1705 3.3030 43.7670 ;
      RECT 3.1770 40.1705 3.1950 43.7670 ;
      RECT 3.0690 40.1705 3.0870 43.7670 ;
      RECT 2.9610 40.1705 2.9790 43.7670 ;
      RECT 2.8530 40.1705 2.8710 43.7670 ;
      RECT 2.7450 40.1705 2.7630 43.7670 ;
      RECT 2.6370 40.1705 2.6550 43.7670 ;
      RECT 2.5290 40.1705 2.5470 43.7670 ;
      RECT 2.4210 40.1705 2.4390 43.7670 ;
      RECT 2.3130 40.1705 2.3310 43.7670 ;
      RECT 2.2050 40.1705 2.2230 43.7670 ;
      RECT 2.0970 40.1705 2.1150 43.7670 ;
      RECT 1.9890 40.1705 2.0070 43.7670 ;
      RECT 1.8810 40.1705 1.8990 43.7670 ;
      RECT 1.7730 40.1705 1.7910 43.7670 ;
      RECT 1.6650 40.1705 1.6830 43.7670 ;
      RECT 1.5570 40.1705 1.5750 43.7670 ;
      RECT 1.4490 40.1705 1.4670 43.7670 ;
      RECT 1.3410 40.1705 1.3590 43.7670 ;
      RECT 1.2330 40.1705 1.2510 43.7670 ;
      RECT 1.1250 40.1705 1.1430 43.7670 ;
      RECT 1.0170 40.1705 1.0350 43.7670 ;
      RECT 0.9090 40.1705 0.9270 43.7670 ;
      RECT 0.8010 40.1705 0.8190 43.7670 ;
      RECT 0.6930 40.1705 0.7110 43.7670 ;
      RECT 0.5850 40.1705 0.6030 43.7670 ;
      RECT 0.4770 40.1705 0.4950 43.7670 ;
      RECT 0.3690 40.1705 0.3870 43.7670 ;
      RECT 0.3330 43.9590 0.3510 44.6637 ;
      RECT 0.3330 45.4170 0.3510 46.5870 ;
      RECT 0.2970 44.0225 0.3150 44.7125 ;
      RECT 0.2970 44.7635 0.3150 45.7500 ;
      RECT 0.2970 45.7900 0.3150 46.4070 ;
      RECT 0.2610 40.1705 0.2790 48.3775 ;
      RECT 0.2250 42.6750 0.2430 42.7440 ;
      RECT 0.2250 44.2950 0.2430 44.3780 ;
      RECT 0.1890 43.9900 0.2070 48.3440 ;
        RECT 8.6990 48.4320 8.7170 49.3675 ;
        RECT 8.6630 48.4320 8.6810 49.3675 ;
        RECT 8.6270 49.0090 8.6450 49.3315 ;
        RECT 8.5100 49.2060 8.5280 49.3155 ;
        RECT 8.5010 48.4645 8.5190 48.7040 ;
        RECT 8.4650 49.0455 8.4830 49.1990 ;
        RECT 8.3840 49.0710 8.4020 49.3290 ;
        RECT 7.8440 48.4320 7.8620 49.3675 ;
        RECT 7.8080 48.4320 7.8260 49.3675 ;
        RECT 7.7720 48.6130 7.7900 49.1810 ;
        RECT 8.6990 49.5120 8.7170 50.4475 ;
        RECT 8.6630 49.5120 8.6810 50.4475 ;
        RECT 8.6270 50.0890 8.6450 50.4115 ;
        RECT 8.5100 50.2860 8.5280 50.3955 ;
        RECT 8.5010 49.5445 8.5190 49.7840 ;
        RECT 8.4650 50.1255 8.4830 50.2790 ;
        RECT 8.3840 50.1510 8.4020 50.4090 ;
        RECT 7.8440 49.5120 7.8620 50.4475 ;
        RECT 7.8080 49.5120 7.8260 50.4475 ;
        RECT 7.7720 49.6930 7.7900 50.2610 ;
        RECT 8.6990 50.5920 8.7170 51.5275 ;
        RECT 8.6630 50.5920 8.6810 51.5275 ;
        RECT 8.6270 51.1690 8.6450 51.4915 ;
        RECT 8.5100 51.3660 8.5280 51.4755 ;
        RECT 8.5010 50.6245 8.5190 50.8640 ;
        RECT 8.4650 51.2055 8.4830 51.3590 ;
        RECT 8.3840 51.2310 8.4020 51.4890 ;
        RECT 7.8440 50.5920 7.8620 51.5275 ;
        RECT 7.8080 50.5920 7.8260 51.5275 ;
        RECT 7.7720 50.7730 7.7900 51.3410 ;
        RECT 8.6990 51.6720 8.7170 52.6075 ;
        RECT 8.6630 51.6720 8.6810 52.6075 ;
        RECT 8.6270 52.2490 8.6450 52.5715 ;
        RECT 8.5100 52.4460 8.5280 52.5555 ;
        RECT 8.5010 51.7045 8.5190 51.9440 ;
        RECT 8.4650 52.2855 8.4830 52.4390 ;
        RECT 8.3840 52.3110 8.4020 52.5690 ;
        RECT 7.8440 51.6720 7.8620 52.6075 ;
        RECT 7.8080 51.6720 7.8260 52.6075 ;
        RECT 7.7720 51.8530 7.7900 52.4210 ;
        RECT 8.6990 52.7520 8.7170 53.6875 ;
        RECT 8.6630 52.7520 8.6810 53.6875 ;
        RECT 8.6270 53.3290 8.6450 53.6515 ;
        RECT 8.5100 53.5260 8.5280 53.6355 ;
        RECT 8.5010 52.7845 8.5190 53.0240 ;
        RECT 8.4650 53.3655 8.4830 53.5190 ;
        RECT 8.3840 53.3910 8.4020 53.6490 ;
        RECT 7.8440 52.7520 7.8620 53.6875 ;
        RECT 7.8080 52.7520 7.8260 53.6875 ;
        RECT 7.7720 52.9330 7.7900 53.5010 ;
        RECT 8.6990 53.8320 8.7170 54.7675 ;
        RECT 8.6630 53.8320 8.6810 54.7675 ;
        RECT 8.6270 54.4090 8.6450 54.7315 ;
        RECT 8.5100 54.6060 8.5280 54.7155 ;
        RECT 8.5010 53.8645 8.5190 54.1040 ;
        RECT 8.4650 54.4455 8.4830 54.5990 ;
        RECT 8.3840 54.4710 8.4020 54.7290 ;
        RECT 7.8440 53.8320 7.8620 54.7675 ;
        RECT 7.8080 53.8320 7.8260 54.7675 ;
        RECT 7.7720 54.0130 7.7900 54.5810 ;
        RECT 8.6990 54.9120 8.7170 55.8475 ;
        RECT 8.6630 54.9120 8.6810 55.8475 ;
        RECT 8.6270 55.4890 8.6450 55.8115 ;
        RECT 8.5100 55.6860 8.5280 55.7955 ;
        RECT 8.5010 54.9445 8.5190 55.1840 ;
        RECT 8.4650 55.5255 8.4830 55.6790 ;
        RECT 8.3840 55.5510 8.4020 55.8090 ;
        RECT 7.8440 54.9120 7.8620 55.8475 ;
        RECT 7.8080 54.9120 7.8260 55.8475 ;
        RECT 7.7720 55.0930 7.7900 55.6610 ;
        RECT 8.6990 55.9920 8.7170 56.9275 ;
        RECT 8.6630 55.9920 8.6810 56.9275 ;
        RECT 8.6270 56.5690 8.6450 56.8915 ;
        RECT 8.5100 56.7660 8.5280 56.8755 ;
        RECT 8.5010 56.0245 8.5190 56.2640 ;
        RECT 8.4650 56.6055 8.4830 56.7590 ;
        RECT 8.3840 56.6310 8.4020 56.8890 ;
        RECT 7.8440 55.9920 7.8620 56.9275 ;
        RECT 7.8080 55.9920 7.8260 56.9275 ;
        RECT 7.7720 56.1730 7.7900 56.7410 ;
        RECT 8.6990 57.0720 8.7170 58.0075 ;
        RECT 8.6630 57.0720 8.6810 58.0075 ;
        RECT 8.6270 57.6490 8.6450 57.9715 ;
        RECT 8.5100 57.8460 8.5280 57.9555 ;
        RECT 8.5010 57.1045 8.5190 57.3440 ;
        RECT 8.4650 57.6855 8.4830 57.8390 ;
        RECT 8.3840 57.7110 8.4020 57.9690 ;
        RECT 7.8440 57.0720 7.8620 58.0075 ;
        RECT 7.8080 57.0720 7.8260 58.0075 ;
        RECT 7.7720 57.2530 7.7900 57.8210 ;
        RECT 8.6990 58.1520 8.7170 59.0875 ;
        RECT 8.6630 58.1520 8.6810 59.0875 ;
        RECT 8.6270 58.7290 8.6450 59.0515 ;
        RECT 8.5100 58.9260 8.5280 59.0355 ;
        RECT 8.5010 58.1845 8.5190 58.4240 ;
        RECT 8.4650 58.7655 8.4830 58.9190 ;
        RECT 8.3840 58.7910 8.4020 59.0490 ;
        RECT 7.8440 58.1520 7.8620 59.0875 ;
        RECT 7.8080 58.1520 7.8260 59.0875 ;
        RECT 7.7720 58.3330 7.7900 58.9010 ;
        RECT 8.6990 59.2320 8.7170 60.1675 ;
        RECT 8.6630 59.2320 8.6810 60.1675 ;
        RECT 8.6270 59.8090 8.6450 60.1315 ;
        RECT 8.5100 60.0060 8.5280 60.1155 ;
        RECT 8.5010 59.2645 8.5190 59.5040 ;
        RECT 8.4650 59.8455 8.4830 59.9990 ;
        RECT 8.3840 59.8710 8.4020 60.1290 ;
        RECT 7.8440 59.2320 7.8620 60.1675 ;
        RECT 7.8080 59.2320 7.8260 60.1675 ;
        RECT 7.7720 59.4130 7.7900 59.9810 ;
        RECT 8.6990 60.3120 8.7170 61.2475 ;
        RECT 8.6630 60.3120 8.6810 61.2475 ;
        RECT 8.6270 60.8890 8.6450 61.2115 ;
        RECT 8.5100 61.0860 8.5280 61.1955 ;
        RECT 8.5010 60.3445 8.5190 60.5840 ;
        RECT 8.4650 60.9255 8.4830 61.0790 ;
        RECT 8.3840 60.9510 8.4020 61.2090 ;
        RECT 7.8440 60.3120 7.8620 61.2475 ;
        RECT 7.8080 60.3120 7.8260 61.2475 ;
        RECT 7.7720 60.4930 7.7900 61.0610 ;
        RECT 8.6990 61.3920 8.7170 62.3275 ;
        RECT 8.6630 61.3920 8.6810 62.3275 ;
        RECT 8.6270 61.9690 8.6450 62.2915 ;
        RECT 8.5100 62.1660 8.5280 62.2755 ;
        RECT 8.5010 61.4245 8.5190 61.6640 ;
        RECT 8.4650 62.0055 8.4830 62.1590 ;
        RECT 8.3840 62.0310 8.4020 62.2890 ;
        RECT 7.8440 61.3920 7.8620 62.3275 ;
        RECT 7.8080 61.3920 7.8260 62.3275 ;
        RECT 7.7720 61.5730 7.7900 62.1410 ;
        RECT 8.6990 62.4720 8.7170 63.4075 ;
        RECT 8.6630 62.4720 8.6810 63.4075 ;
        RECT 8.6270 63.0490 8.6450 63.3715 ;
        RECT 8.5100 63.2460 8.5280 63.3555 ;
        RECT 8.5010 62.5045 8.5190 62.7440 ;
        RECT 8.4650 63.0855 8.4830 63.2390 ;
        RECT 8.3840 63.1110 8.4020 63.3690 ;
        RECT 7.8440 62.4720 7.8620 63.4075 ;
        RECT 7.8080 62.4720 7.8260 63.4075 ;
        RECT 7.7720 62.6530 7.7900 63.2210 ;
        RECT 8.6990 63.5520 8.7170 64.4875 ;
        RECT 8.6630 63.5520 8.6810 64.4875 ;
        RECT 8.6270 64.1290 8.6450 64.4515 ;
        RECT 8.5100 64.3260 8.5280 64.4355 ;
        RECT 8.5010 63.5845 8.5190 63.8240 ;
        RECT 8.4650 64.1655 8.4830 64.3190 ;
        RECT 8.3840 64.1910 8.4020 64.4490 ;
        RECT 7.8440 63.5520 7.8620 64.4875 ;
        RECT 7.8080 63.5520 7.8260 64.4875 ;
        RECT 7.7720 63.7330 7.7900 64.3010 ;
        RECT 8.6990 64.6320 8.7170 65.5675 ;
        RECT 8.6630 64.6320 8.6810 65.5675 ;
        RECT 8.6270 65.2090 8.6450 65.5315 ;
        RECT 8.5100 65.4060 8.5280 65.5155 ;
        RECT 8.5010 64.6645 8.5190 64.9040 ;
        RECT 8.4650 65.2455 8.4830 65.3990 ;
        RECT 8.3840 65.2710 8.4020 65.5290 ;
        RECT 7.8440 64.6320 7.8620 65.5675 ;
        RECT 7.8080 64.6320 7.8260 65.5675 ;
        RECT 7.7720 64.8130 7.7900 65.3810 ;
        RECT 8.6990 65.7120 8.7170 66.6475 ;
        RECT 8.6630 65.7120 8.6810 66.6475 ;
        RECT 8.6270 66.2890 8.6450 66.6115 ;
        RECT 8.5100 66.4860 8.5280 66.5955 ;
        RECT 8.5010 65.7445 8.5190 65.9840 ;
        RECT 8.4650 66.3255 8.4830 66.4790 ;
        RECT 8.3840 66.3510 8.4020 66.6090 ;
        RECT 7.8440 65.7120 7.8620 66.6475 ;
        RECT 7.8080 65.7120 7.8260 66.6475 ;
        RECT 7.7720 65.8930 7.7900 66.4610 ;
        RECT 8.6990 66.7920 8.7170 67.7275 ;
        RECT 8.6630 66.7920 8.6810 67.7275 ;
        RECT 8.6270 67.3690 8.6450 67.6915 ;
        RECT 8.5100 67.5660 8.5280 67.6755 ;
        RECT 8.5010 66.8245 8.5190 67.0640 ;
        RECT 8.4650 67.4055 8.4830 67.5590 ;
        RECT 8.3840 67.4310 8.4020 67.6890 ;
        RECT 7.8440 66.7920 7.8620 67.7275 ;
        RECT 7.8080 66.7920 7.8260 67.7275 ;
        RECT 7.7720 66.9730 7.7900 67.5410 ;
        RECT 8.6990 67.8720 8.7170 68.8075 ;
        RECT 8.6630 67.8720 8.6810 68.8075 ;
        RECT 8.6270 68.4490 8.6450 68.7715 ;
        RECT 8.5100 68.6460 8.5280 68.7555 ;
        RECT 8.5010 67.9045 8.5190 68.1440 ;
        RECT 8.4650 68.4855 8.4830 68.6390 ;
        RECT 8.3840 68.5110 8.4020 68.7690 ;
        RECT 7.8440 67.8720 7.8620 68.8075 ;
        RECT 7.8080 67.8720 7.8260 68.8075 ;
        RECT 7.7720 68.0530 7.7900 68.6210 ;
        RECT 8.6990 68.9520 8.7170 69.8875 ;
        RECT 8.6630 68.9520 8.6810 69.8875 ;
        RECT 8.6270 69.5290 8.6450 69.8515 ;
        RECT 8.5100 69.7260 8.5280 69.8355 ;
        RECT 8.5010 68.9845 8.5190 69.2240 ;
        RECT 8.4650 69.5655 8.4830 69.7190 ;
        RECT 8.3840 69.5910 8.4020 69.8490 ;
        RECT 7.8440 68.9520 7.8620 69.8875 ;
        RECT 7.8080 68.9520 7.8260 69.8875 ;
        RECT 7.7720 69.1330 7.7900 69.7010 ;
        RECT 8.6990 70.0320 8.7170 70.9675 ;
        RECT 8.6630 70.0320 8.6810 70.9675 ;
        RECT 8.6270 70.6090 8.6450 70.9315 ;
        RECT 8.5100 70.8060 8.5280 70.9155 ;
        RECT 8.5010 70.0645 8.5190 70.3040 ;
        RECT 8.4650 70.6455 8.4830 70.7990 ;
        RECT 8.3840 70.6710 8.4020 70.9290 ;
        RECT 7.8440 70.0320 7.8620 70.9675 ;
        RECT 7.8080 70.0320 7.8260 70.9675 ;
        RECT 7.7720 70.2130 7.7900 70.7810 ;
        RECT 8.6990 71.1120 8.7170 72.0475 ;
        RECT 8.6630 71.1120 8.6810 72.0475 ;
        RECT 8.6270 71.6890 8.6450 72.0115 ;
        RECT 8.5100 71.8860 8.5280 71.9955 ;
        RECT 8.5010 71.1445 8.5190 71.3840 ;
        RECT 8.4650 71.7255 8.4830 71.8790 ;
        RECT 8.3840 71.7510 8.4020 72.0090 ;
        RECT 7.8440 71.1120 7.8620 72.0475 ;
        RECT 7.8080 71.1120 7.8260 72.0475 ;
        RECT 7.7720 71.2930 7.7900 71.8610 ;
        RECT 8.6990 72.1920 8.7170 73.1275 ;
        RECT 8.6630 72.1920 8.6810 73.1275 ;
        RECT 8.6270 72.7690 8.6450 73.0915 ;
        RECT 8.5100 72.9660 8.5280 73.0755 ;
        RECT 8.5010 72.2245 8.5190 72.4640 ;
        RECT 8.4650 72.8055 8.4830 72.9590 ;
        RECT 8.3840 72.8310 8.4020 73.0890 ;
        RECT 7.8440 72.1920 7.8620 73.1275 ;
        RECT 7.8080 72.1920 7.8260 73.1275 ;
        RECT 7.7720 72.3730 7.7900 72.9410 ;
        RECT 8.6990 73.2720 8.7170 74.2075 ;
        RECT 8.6630 73.2720 8.6810 74.2075 ;
        RECT 8.6270 73.8490 8.6450 74.1715 ;
        RECT 8.5100 74.0460 8.5280 74.1555 ;
        RECT 8.5010 73.3045 8.5190 73.5440 ;
        RECT 8.4650 73.8855 8.4830 74.0390 ;
        RECT 8.3840 73.9110 8.4020 74.1690 ;
        RECT 7.8440 73.2720 7.8620 74.2075 ;
        RECT 7.8080 73.2720 7.8260 74.2075 ;
        RECT 7.7720 73.4530 7.7900 74.0210 ;
        RECT 8.6990 74.3520 8.7170 75.2875 ;
        RECT 8.6630 74.3520 8.6810 75.2875 ;
        RECT 8.6270 74.9290 8.6450 75.2515 ;
        RECT 8.5100 75.1260 8.5280 75.2355 ;
        RECT 8.5010 74.3845 8.5190 74.6240 ;
        RECT 8.4650 74.9655 8.4830 75.1190 ;
        RECT 8.3840 74.9910 8.4020 75.2490 ;
        RECT 7.8440 74.3520 7.8620 75.2875 ;
        RECT 7.8080 74.3520 7.8260 75.2875 ;
        RECT 7.7720 74.5330 7.7900 75.1010 ;
        RECT 8.6990 75.4320 8.7170 76.3675 ;
        RECT 8.6630 75.4320 8.6810 76.3675 ;
        RECT 8.6270 76.0090 8.6450 76.3315 ;
        RECT 8.5100 76.2060 8.5280 76.3155 ;
        RECT 8.5010 75.4645 8.5190 75.7040 ;
        RECT 8.4650 76.0455 8.4830 76.1990 ;
        RECT 8.3840 76.0710 8.4020 76.3290 ;
        RECT 7.8440 75.4320 7.8620 76.3675 ;
        RECT 7.8080 75.4320 7.8260 76.3675 ;
        RECT 7.7720 75.6130 7.7900 76.1810 ;
        RECT 8.6990 76.5120 8.7170 77.4475 ;
        RECT 8.6630 76.5120 8.6810 77.4475 ;
        RECT 8.6270 77.0890 8.6450 77.4115 ;
        RECT 8.5100 77.2860 8.5280 77.3955 ;
        RECT 8.5010 76.5445 8.5190 76.7840 ;
        RECT 8.4650 77.1255 8.4830 77.2790 ;
        RECT 8.3840 77.1510 8.4020 77.4090 ;
        RECT 7.8440 76.5120 7.8620 77.4475 ;
        RECT 7.8080 76.5120 7.8260 77.4475 ;
        RECT 7.7720 76.6930 7.7900 77.2610 ;
        RECT 8.6990 77.5920 8.7170 78.5275 ;
        RECT 8.6630 77.5920 8.6810 78.5275 ;
        RECT 8.6270 78.1690 8.6450 78.4915 ;
        RECT 8.5100 78.3660 8.5280 78.4755 ;
        RECT 8.5010 77.6245 8.5190 77.8640 ;
        RECT 8.4650 78.2055 8.4830 78.3590 ;
        RECT 8.3840 78.2310 8.4020 78.4890 ;
        RECT 7.8440 77.5920 7.8620 78.5275 ;
        RECT 7.8080 77.5920 7.8260 78.5275 ;
        RECT 7.7720 77.7730 7.7900 78.3410 ;
        RECT 8.6990 78.6720 8.7170 79.6075 ;
        RECT 8.6630 78.6720 8.6810 79.6075 ;
        RECT 8.6270 79.2490 8.6450 79.5715 ;
        RECT 8.5100 79.4460 8.5280 79.5555 ;
        RECT 8.5010 78.7045 8.5190 78.9440 ;
        RECT 8.4650 79.2855 8.4830 79.4390 ;
        RECT 8.3840 79.3110 8.4020 79.5690 ;
        RECT 7.8440 78.6720 7.8620 79.6075 ;
        RECT 7.8080 78.6720 7.8260 79.6075 ;
        RECT 7.7720 78.8530 7.7900 79.4210 ;
        RECT 8.6990 79.7520 8.7170 80.6875 ;
        RECT 8.6630 79.7520 8.6810 80.6875 ;
        RECT 8.6270 80.3290 8.6450 80.6515 ;
        RECT 8.5100 80.5260 8.5280 80.6355 ;
        RECT 8.5010 79.7845 8.5190 80.0240 ;
        RECT 8.4650 80.3655 8.4830 80.5190 ;
        RECT 8.3840 80.3910 8.4020 80.6490 ;
        RECT 7.8440 79.7520 7.8620 80.6875 ;
        RECT 7.8080 79.7520 7.8260 80.6875 ;
        RECT 7.7720 79.9330 7.7900 80.5010 ;
        RECT 8.6990 80.8320 8.7170 81.7675 ;
        RECT 8.6630 80.8320 8.6810 81.7675 ;
        RECT 8.6270 81.4090 8.6450 81.7315 ;
        RECT 8.5100 81.6060 8.5280 81.7155 ;
        RECT 8.5010 80.8645 8.5190 81.1040 ;
        RECT 8.4650 81.4455 8.4830 81.5990 ;
        RECT 8.3840 81.4710 8.4020 81.7290 ;
        RECT 7.8440 80.8320 7.8620 81.7675 ;
        RECT 7.8080 80.8320 7.8260 81.7675 ;
        RECT 7.7720 81.0130 7.7900 81.5810 ;
        RECT 8.6990 81.9120 8.7170 82.8475 ;
        RECT 8.6630 81.9120 8.6810 82.8475 ;
        RECT 8.6270 82.4890 8.6450 82.8115 ;
        RECT 8.5100 82.6860 8.5280 82.7955 ;
        RECT 8.5010 81.9445 8.5190 82.1840 ;
        RECT 8.4650 82.5255 8.4830 82.6790 ;
        RECT 8.3840 82.5510 8.4020 82.8090 ;
        RECT 7.8440 81.9120 7.8620 82.8475 ;
        RECT 7.8080 81.9120 7.8260 82.8475 ;
        RECT 7.7720 82.0930 7.7900 82.6610 ;
        RECT 8.6990 82.9920 8.7170 83.9275 ;
        RECT 8.6630 82.9920 8.6810 83.9275 ;
        RECT 8.6270 83.5690 8.6450 83.8915 ;
        RECT 8.5100 83.7660 8.5280 83.8755 ;
        RECT 8.5010 83.0245 8.5190 83.2640 ;
        RECT 8.4650 83.6055 8.4830 83.7590 ;
        RECT 8.3840 83.6310 8.4020 83.8890 ;
        RECT 7.8440 82.9920 7.8620 83.9275 ;
        RECT 7.8080 82.9920 7.8260 83.9275 ;
        RECT 7.7720 83.1730 7.7900 83.7410 ;
        RECT 8.6990 84.0720 8.7170 85.0075 ;
        RECT 8.6630 84.0720 8.6810 85.0075 ;
        RECT 8.6270 84.6490 8.6450 84.9715 ;
        RECT 8.5100 84.8460 8.5280 84.9555 ;
        RECT 8.5010 84.1045 8.5190 84.3440 ;
        RECT 8.4650 84.6855 8.4830 84.8390 ;
        RECT 8.3840 84.7110 8.4020 84.9690 ;
        RECT 7.8440 84.0720 7.8620 85.0075 ;
        RECT 7.8080 84.0720 7.8260 85.0075 ;
        RECT 7.7720 84.2530 7.7900 84.8210 ;
        RECT 8.6990 85.1520 8.7170 86.0875 ;
        RECT 8.6630 85.1520 8.6810 86.0875 ;
        RECT 8.6270 85.7290 8.6450 86.0515 ;
        RECT 8.5100 85.9260 8.5280 86.0355 ;
        RECT 8.5010 85.1845 8.5190 85.4240 ;
        RECT 8.4650 85.7655 8.4830 85.9190 ;
        RECT 8.3840 85.7910 8.4020 86.0490 ;
        RECT 7.8440 85.1520 7.8620 86.0875 ;
        RECT 7.8080 85.1520 7.8260 86.0875 ;
        RECT 7.7720 85.3330 7.7900 85.9010 ;
        RECT 8.6990 86.2320 8.7170 87.1675 ;
        RECT 8.6630 86.2320 8.6810 87.1675 ;
        RECT 8.6270 86.8090 8.6450 87.1315 ;
        RECT 8.5100 87.0060 8.5280 87.1155 ;
        RECT 8.5010 86.2645 8.5190 86.5040 ;
        RECT 8.4650 86.8455 8.4830 86.9990 ;
        RECT 8.3840 86.8710 8.4020 87.1290 ;
        RECT 7.8440 86.2320 7.8620 87.1675 ;
        RECT 7.8080 86.2320 7.8260 87.1675 ;
        RECT 7.7720 86.4130 7.7900 86.9810 ;
        RECT 8.6990 87.3120 8.7170 88.2475 ;
        RECT 8.6630 87.3120 8.6810 88.2475 ;
        RECT 8.6270 87.8890 8.6450 88.2115 ;
        RECT 8.5100 88.0860 8.5280 88.1955 ;
        RECT 8.5010 87.3445 8.5190 87.5840 ;
        RECT 8.4650 87.9255 8.4830 88.0790 ;
        RECT 8.3840 87.9510 8.4020 88.2090 ;
        RECT 7.8440 87.3120 7.8620 88.2475 ;
        RECT 7.8080 87.3120 7.8260 88.2475 ;
        RECT 7.7720 87.4930 7.7900 88.0610 ;
  LAYER M3 SPACING 0.018  ;
      RECT 8.6410 0.2565 8.7690 1.3500 ;
      RECT 8.6270 0.9220 8.7690 1.2445 ;
      RECT 8.4790 0.6490 8.5410 1.3500 ;
      RECT 8.4650 0.9585 8.5410 1.1120 ;
      RECT 8.4790 0.2565 8.5050 1.3500 ;
      RECT 8.4790 0.3775 8.5190 0.6170 ;
      RECT 8.4790 0.2565 8.5410 0.3455 ;
      RECT 8.1820 0.7070 8.3880 1.3500 ;
      RECT 8.3620 0.2565 8.3880 1.3500 ;
      RECT 8.1820 0.9840 8.4020 1.2420 ;
      RECT 8.1820 0.2565 8.2800 1.3500 ;
      RECT 7.7650 0.2565 7.8480 1.3500 ;
      RECT 7.7650 0.3450 7.8620 1.2805 ;
      RECT 16.4440 0.2565 16.5290 1.3500 ;
      RECT 16.3000 0.2565 16.3260 1.3500 ;
      RECT 16.1920 0.2565 16.2180 1.3500 ;
      RECT 16.0840 0.2565 16.1100 1.3500 ;
      RECT 15.9760 0.2565 16.0020 1.3500 ;
      RECT 15.8680 0.2565 15.8940 1.3500 ;
      RECT 15.7600 0.2565 15.7860 1.3500 ;
      RECT 15.6520 0.2565 15.6780 1.3500 ;
      RECT 15.5440 0.2565 15.5700 1.3500 ;
      RECT 15.4360 0.2565 15.4620 1.3500 ;
      RECT 15.3280 0.2565 15.3540 1.3500 ;
      RECT 15.2200 0.2565 15.2460 1.3500 ;
      RECT 15.1120 0.2565 15.1380 1.3500 ;
      RECT 15.0040 0.2565 15.0300 1.3500 ;
      RECT 14.8960 0.2565 14.9220 1.3500 ;
      RECT 14.7880 0.2565 14.8140 1.3500 ;
      RECT 14.6800 0.2565 14.7060 1.3500 ;
      RECT 14.5720 0.2565 14.5980 1.3500 ;
      RECT 14.4640 0.2565 14.4900 1.3500 ;
      RECT 14.3560 0.2565 14.3820 1.3500 ;
      RECT 14.2480 0.2565 14.2740 1.3500 ;
      RECT 14.1400 0.2565 14.1660 1.3500 ;
      RECT 14.0320 0.2565 14.0580 1.3500 ;
      RECT 13.9240 0.2565 13.9500 1.3500 ;
      RECT 13.8160 0.2565 13.8420 1.3500 ;
      RECT 13.7080 0.2565 13.7340 1.3500 ;
      RECT 13.6000 0.2565 13.6260 1.3500 ;
      RECT 13.4920 0.2565 13.5180 1.3500 ;
      RECT 13.3840 0.2565 13.4100 1.3500 ;
      RECT 13.2760 0.2565 13.3020 1.3500 ;
      RECT 13.1680 0.2565 13.1940 1.3500 ;
      RECT 13.0600 0.2565 13.0860 1.3500 ;
      RECT 12.9520 0.2565 12.9780 1.3500 ;
      RECT 12.8440 0.2565 12.8700 1.3500 ;
      RECT 12.7360 0.2565 12.7620 1.3500 ;
      RECT 12.6280 0.2565 12.6540 1.3500 ;
      RECT 12.5200 0.2565 12.5460 1.3500 ;
      RECT 12.4120 0.2565 12.4380 1.3500 ;
      RECT 12.3040 0.2565 12.3300 1.3500 ;
      RECT 12.1960 0.2565 12.2220 1.3500 ;
      RECT 12.0880 0.2565 12.1140 1.3500 ;
      RECT 11.9800 0.2565 12.0060 1.3500 ;
      RECT 11.8720 0.2565 11.8980 1.3500 ;
      RECT 11.7640 0.2565 11.7900 1.3500 ;
      RECT 11.6560 0.2565 11.6820 1.3500 ;
      RECT 11.5480 0.2565 11.5740 1.3500 ;
      RECT 11.4400 0.2565 11.4660 1.3500 ;
      RECT 11.3320 0.2565 11.3580 1.3500 ;
      RECT 11.2240 0.2565 11.2500 1.3500 ;
      RECT 11.1160 0.2565 11.1420 1.3500 ;
      RECT 11.0080 0.2565 11.0340 1.3500 ;
      RECT 10.9000 0.2565 10.9260 1.3500 ;
      RECT 10.7920 0.2565 10.8180 1.3500 ;
      RECT 10.6840 0.2565 10.7100 1.3500 ;
      RECT 10.5760 0.2565 10.6020 1.3500 ;
      RECT 10.4680 0.2565 10.4940 1.3500 ;
      RECT 10.3600 0.2565 10.3860 1.3500 ;
      RECT 10.2520 0.2565 10.2780 1.3500 ;
      RECT 10.1440 0.2565 10.1700 1.3500 ;
      RECT 10.0360 0.2565 10.0620 1.3500 ;
      RECT 9.9280 0.2565 9.9540 1.3500 ;
      RECT 9.8200 0.2565 9.8460 1.3500 ;
      RECT 9.7120 0.2565 9.7380 1.3500 ;
      RECT 9.6040 0.2565 9.6300 1.3500 ;
      RECT 9.4960 0.2565 9.5220 1.3500 ;
      RECT 9.3880 0.2565 9.4140 1.3500 ;
      RECT 9.1750 0.2565 9.2520 1.3500 ;
      RECT 7.2820 0.2565 7.3590 1.3500 ;
      RECT 7.1200 0.2565 7.1460 1.3500 ;
      RECT 7.0120 0.2565 7.0380 1.3500 ;
      RECT 6.9040 0.2565 6.9300 1.3500 ;
      RECT 6.7960 0.2565 6.8220 1.3500 ;
      RECT 6.6880 0.2565 6.7140 1.3500 ;
      RECT 6.5800 0.2565 6.6060 1.3500 ;
      RECT 6.4720 0.2565 6.4980 1.3500 ;
      RECT 6.3640 0.2565 6.3900 1.3500 ;
      RECT 6.2560 0.2565 6.2820 1.3500 ;
      RECT 6.1480 0.2565 6.1740 1.3500 ;
      RECT 6.0400 0.2565 6.0660 1.3500 ;
      RECT 5.9320 0.2565 5.9580 1.3500 ;
      RECT 5.8240 0.2565 5.8500 1.3500 ;
      RECT 5.7160 0.2565 5.7420 1.3500 ;
      RECT 5.6080 0.2565 5.6340 1.3500 ;
      RECT 5.5000 0.2565 5.5260 1.3500 ;
      RECT 5.3920 0.2565 5.4180 1.3500 ;
      RECT 5.2840 0.2565 5.3100 1.3500 ;
      RECT 5.1760 0.2565 5.2020 1.3500 ;
      RECT 5.0680 0.2565 5.0940 1.3500 ;
      RECT 4.9600 0.2565 4.9860 1.3500 ;
      RECT 4.8520 0.2565 4.8780 1.3500 ;
      RECT 4.7440 0.2565 4.7700 1.3500 ;
      RECT 4.6360 0.2565 4.6620 1.3500 ;
      RECT 4.5280 0.2565 4.5540 1.3500 ;
      RECT 4.4200 0.2565 4.4460 1.3500 ;
      RECT 4.3120 0.2565 4.3380 1.3500 ;
      RECT 4.2040 0.2565 4.2300 1.3500 ;
      RECT 4.0960 0.2565 4.1220 1.3500 ;
      RECT 3.9880 0.2565 4.0140 1.3500 ;
      RECT 3.8800 0.2565 3.9060 1.3500 ;
      RECT 3.7720 0.2565 3.7980 1.3500 ;
      RECT 3.6640 0.2565 3.6900 1.3500 ;
      RECT 3.5560 0.2565 3.5820 1.3500 ;
      RECT 3.4480 0.2565 3.4740 1.3500 ;
      RECT 3.3400 0.2565 3.3660 1.3500 ;
      RECT 3.2320 0.2565 3.2580 1.3500 ;
      RECT 3.1240 0.2565 3.1500 1.3500 ;
      RECT 3.0160 0.2565 3.0420 1.3500 ;
      RECT 2.9080 0.2565 2.9340 1.3500 ;
      RECT 2.8000 0.2565 2.8260 1.3500 ;
      RECT 2.6920 0.2565 2.7180 1.3500 ;
      RECT 2.5840 0.2565 2.6100 1.3500 ;
      RECT 2.4760 0.2565 2.5020 1.3500 ;
      RECT 2.3680 0.2565 2.3940 1.3500 ;
      RECT 2.2600 0.2565 2.2860 1.3500 ;
      RECT 2.1520 0.2565 2.1780 1.3500 ;
      RECT 2.0440 0.2565 2.0700 1.3500 ;
      RECT 1.9360 0.2565 1.9620 1.3500 ;
      RECT 1.8280 0.2565 1.8540 1.3500 ;
      RECT 1.7200 0.2565 1.7460 1.3500 ;
      RECT 1.6120 0.2565 1.6380 1.3500 ;
      RECT 1.5040 0.2565 1.5300 1.3500 ;
      RECT 1.3960 0.2565 1.4220 1.3500 ;
      RECT 1.2880 0.2565 1.3140 1.3500 ;
      RECT 1.1800 0.2565 1.2060 1.3500 ;
      RECT 1.0720 0.2565 1.0980 1.3500 ;
      RECT 0.9640 0.2565 0.9900 1.3500 ;
      RECT 0.8560 0.2565 0.8820 1.3500 ;
      RECT 0.7480 0.2565 0.7740 1.3500 ;
      RECT 0.6400 0.2565 0.6660 1.3500 ;
      RECT 0.5320 0.2565 0.5580 1.3500 ;
      RECT 0.4240 0.2565 0.4500 1.3500 ;
      RECT 0.3160 0.2565 0.3420 1.3500 ;
      RECT 0.2080 0.2565 0.2340 1.3500 ;
      RECT 0.0050 0.2565 0.0900 1.3500 ;
      RECT 8.6410 1.3365 8.7690 2.4300 ;
      RECT 8.6270 2.0020 8.7690 2.3245 ;
      RECT 8.4790 1.7290 8.5410 2.4300 ;
      RECT 8.4650 2.0385 8.5410 2.1920 ;
      RECT 8.4790 1.3365 8.5050 2.4300 ;
      RECT 8.4790 1.4575 8.5190 1.6970 ;
      RECT 8.4790 1.3365 8.5410 1.4255 ;
      RECT 8.1820 1.7870 8.3880 2.4300 ;
      RECT 8.3620 1.3365 8.3880 2.4300 ;
      RECT 8.1820 2.0640 8.4020 2.3220 ;
      RECT 8.1820 1.3365 8.2800 2.4300 ;
      RECT 7.7650 1.3365 7.8480 2.4300 ;
      RECT 7.7650 1.4250 7.8620 2.3605 ;
      RECT 16.4440 1.3365 16.5290 2.4300 ;
      RECT 16.3000 1.3365 16.3260 2.4300 ;
      RECT 16.1920 1.3365 16.2180 2.4300 ;
      RECT 16.0840 1.3365 16.1100 2.4300 ;
      RECT 15.9760 1.3365 16.0020 2.4300 ;
      RECT 15.8680 1.3365 15.8940 2.4300 ;
      RECT 15.7600 1.3365 15.7860 2.4300 ;
      RECT 15.6520 1.3365 15.6780 2.4300 ;
      RECT 15.5440 1.3365 15.5700 2.4300 ;
      RECT 15.4360 1.3365 15.4620 2.4300 ;
      RECT 15.3280 1.3365 15.3540 2.4300 ;
      RECT 15.2200 1.3365 15.2460 2.4300 ;
      RECT 15.1120 1.3365 15.1380 2.4300 ;
      RECT 15.0040 1.3365 15.0300 2.4300 ;
      RECT 14.8960 1.3365 14.9220 2.4300 ;
      RECT 14.7880 1.3365 14.8140 2.4300 ;
      RECT 14.6800 1.3365 14.7060 2.4300 ;
      RECT 14.5720 1.3365 14.5980 2.4300 ;
      RECT 14.4640 1.3365 14.4900 2.4300 ;
      RECT 14.3560 1.3365 14.3820 2.4300 ;
      RECT 14.2480 1.3365 14.2740 2.4300 ;
      RECT 14.1400 1.3365 14.1660 2.4300 ;
      RECT 14.0320 1.3365 14.0580 2.4300 ;
      RECT 13.9240 1.3365 13.9500 2.4300 ;
      RECT 13.8160 1.3365 13.8420 2.4300 ;
      RECT 13.7080 1.3365 13.7340 2.4300 ;
      RECT 13.6000 1.3365 13.6260 2.4300 ;
      RECT 13.4920 1.3365 13.5180 2.4300 ;
      RECT 13.3840 1.3365 13.4100 2.4300 ;
      RECT 13.2760 1.3365 13.3020 2.4300 ;
      RECT 13.1680 1.3365 13.1940 2.4300 ;
      RECT 13.0600 1.3365 13.0860 2.4300 ;
      RECT 12.9520 1.3365 12.9780 2.4300 ;
      RECT 12.8440 1.3365 12.8700 2.4300 ;
      RECT 12.7360 1.3365 12.7620 2.4300 ;
      RECT 12.6280 1.3365 12.6540 2.4300 ;
      RECT 12.5200 1.3365 12.5460 2.4300 ;
      RECT 12.4120 1.3365 12.4380 2.4300 ;
      RECT 12.3040 1.3365 12.3300 2.4300 ;
      RECT 12.1960 1.3365 12.2220 2.4300 ;
      RECT 12.0880 1.3365 12.1140 2.4300 ;
      RECT 11.9800 1.3365 12.0060 2.4300 ;
      RECT 11.8720 1.3365 11.8980 2.4300 ;
      RECT 11.7640 1.3365 11.7900 2.4300 ;
      RECT 11.6560 1.3365 11.6820 2.4300 ;
      RECT 11.5480 1.3365 11.5740 2.4300 ;
      RECT 11.4400 1.3365 11.4660 2.4300 ;
      RECT 11.3320 1.3365 11.3580 2.4300 ;
      RECT 11.2240 1.3365 11.2500 2.4300 ;
      RECT 11.1160 1.3365 11.1420 2.4300 ;
      RECT 11.0080 1.3365 11.0340 2.4300 ;
      RECT 10.9000 1.3365 10.9260 2.4300 ;
      RECT 10.7920 1.3365 10.8180 2.4300 ;
      RECT 10.6840 1.3365 10.7100 2.4300 ;
      RECT 10.5760 1.3365 10.6020 2.4300 ;
      RECT 10.4680 1.3365 10.4940 2.4300 ;
      RECT 10.3600 1.3365 10.3860 2.4300 ;
      RECT 10.2520 1.3365 10.2780 2.4300 ;
      RECT 10.1440 1.3365 10.1700 2.4300 ;
      RECT 10.0360 1.3365 10.0620 2.4300 ;
      RECT 9.9280 1.3365 9.9540 2.4300 ;
      RECT 9.8200 1.3365 9.8460 2.4300 ;
      RECT 9.7120 1.3365 9.7380 2.4300 ;
      RECT 9.6040 1.3365 9.6300 2.4300 ;
      RECT 9.4960 1.3365 9.5220 2.4300 ;
      RECT 9.3880 1.3365 9.4140 2.4300 ;
      RECT 9.1750 1.3365 9.2520 2.4300 ;
      RECT 7.2820 1.3365 7.3590 2.4300 ;
      RECT 7.1200 1.3365 7.1460 2.4300 ;
      RECT 7.0120 1.3365 7.0380 2.4300 ;
      RECT 6.9040 1.3365 6.9300 2.4300 ;
      RECT 6.7960 1.3365 6.8220 2.4300 ;
      RECT 6.6880 1.3365 6.7140 2.4300 ;
      RECT 6.5800 1.3365 6.6060 2.4300 ;
      RECT 6.4720 1.3365 6.4980 2.4300 ;
      RECT 6.3640 1.3365 6.3900 2.4300 ;
      RECT 6.2560 1.3365 6.2820 2.4300 ;
      RECT 6.1480 1.3365 6.1740 2.4300 ;
      RECT 6.0400 1.3365 6.0660 2.4300 ;
      RECT 5.9320 1.3365 5.9580 2.4300 ;
      RECT 5.8240 1.3365 5.8500 2.4300 ;
      RECT 5.7160 1.3365 5.7420 2.4300 ;
      RECT 5.6080 1.3365 5.6340 2.4300 ;
      RECT 5.5000 1.3365 5.5260 2.4300 ;
      RECT 5.3920 1.3365 5.4180 2.4300 ;
      RECT 5.2840 1.3365 5.3100 2.4300 ;
      RECT 5.1760 1.3365 5.2020 2.4300 ;
      RECT 5.0680 1.3365 5.0940 2.4300 ;
      RECT 4.9600 1.3365 4.9860 2.4300 ;
      RECT 4.8520 1.3365 4.8780 2.4300 ;
      RECT 4.7440 1.3365 4.7700 2.4300 ;
      RECT 4.6360 1.3365 4.6620 2.4300 ;
      RECT 4.5280 1.3365 4.5540 2.4300 ;
      RECT 4.4200 1.3365 4.4460 2.4300 ;
      RECT 4.3120 1.3365 4.3380 2.4300 ;
      RECT 4.2040 1.3365 4.2300 2.4300 ;
      RECT 4.0960 1.3365 4.1220 2.4300 ;
      RECT 3.9880 1.3365 4.0140 2.4300 ;
      RECT 3.8800 1.3365 3.9060 2.4300 ;
      RECT 3.7720 1.3365 3.7980 2.4300 ;
      RECT 3.6640 1.3365 3.6900 2.4300 ;
      RECT 3.5560 1.3365 3.5820 2.4300 ;
      RECT 3.4480 1.3365 3.4740 2.4300 ;
      RECT 3.3400 1.3365 3.3660 2.4300 ;
      RECT 3.2320 1.3365 3.2580 2.4300 ;
      RECT 3.1240 1.3365 3.1500 2.4300 ;
      RECT 3.0160 1.3365 3.0420 2.4300 ;
      RECT 2.9080 1.3365 2.9340 2.4300 ;
      RECT 2.8000 1.3365 2.8260 2.4300 ;
      RECT 2.6920 1.3365 2.7180 2.4300 ;
      RECT 2.5840 1.3365 2.6100 2.4300 ;
      RECT 2.4760 1.3365 2.5020 2.4300 ;
      RECT 2.3680 1.3365 2.3940 2.4300 ;
      RECT 2.2600 1.3365 2.2860 2.4300 ;
      RECT 2.1520 1.3365 2.1780 2.4300 ;
      RECT 2.0440 1.3365 2.0700 2.4300 ;
      RECT 1.9360 1.3365 1.9620 2.4300 ;
      RECT 1.8280 1.3365 1.8540 2.4300 ;
      RECT 1.7200 1.3365 1.7460 2.4300 ;
      RECT 1.6120 1.3365 1.6380 2.4300 ;
      RECT 1.5040 1.3365 1.5300 2.4300 ;
      RECT 1.3960 1.3365 1.4220 2.4300 ;
      RECT 1.2880 1.3365 1.3140 2.4300 ;
      RECT 1.1800 1.3365 1.2060 2.4300 ;
      RECT 1.0720 1.3365 1.0980 2.4300 ;
      RECT 0.9640 1.3365 0.9900 2.4300 ;
      RECT 0.8560 1.3365 0.8820 2.4300 ;
      RECT 0.7480 1.3365 0.7740 2.4300 ;
      RECT 0.6400 1.3365 0.6660 2.4300 ;
      RECT 0.5320 1.3365 0.5580 2.4300 ;
      RECT 0.4240 1.3365 0.4500 2.4300 ;
      RECT 0.3160 1.3365 0.3420 2.4300 ;
      RECT 0.2080 1.3365 0.2340 2.4300 ;
      RECT 0.0050 1.3365 0.0900 2.4300 ;
      RECT 8.6410 2.4165 8.7690 3.5100 ;
      RECT 8.6270 3.0820 8.7690 3.4045 ;
      RECT 8.4790 2.8090 8.5410 3.5100 ;
      RECT 8.4650 3.1185 8.5410 3.2720 ;
      RECT 8.4790 2.4165 8.5050 3.5100 ;
      RECT 8.4790 2.5375 8.5190 2.7770 ;
      RECT 8.4790 2.4165 8.5410 2.5055 ;
      RECT 8.1820 2.8670 8.3880 3.5100 ;
      RECT 8.3620 2.4165 8.3880 3.5100 ;
      RECT 8.1820 3.1440 8.4020 3.4020 ;
      RECT 8.1820 2.4165 8.2800 3.5100 ;
      RECT 7.7650 2.4165 7.8480 3.5100 ;
      RECT 7.7650 2.5050 7.8620 3.4405 ;
      RECT 16.4440 2.4165 16.5290 3.5100 ;
      RECT 16.3000 2.4165 16.3260 3.5100 ;
      RECT 16.1920 2.4165 16.2180 3.5100 ;
      RECT 16.0840 2.4165 16.1100 3.5100 ;
      RECT 15.9760 2.4165 16.0020 3.5100 ;
      RECT 15.8680 2.4165 15.8940 3.5100 ;
      RECT 15.7600 2.4165 15.7860 3.5100 ;
      RECT 15.6520 2.4165 15.6780 3.5100 ;
      RECT 15.5440 2.4165 15.5700 3.5100 ;
      RECT 15.4360 2.4165 15.4620 3.5100 ;
      RECT 15.3280 2.4165 15.3540 3.5100 ;
      RECT 15.2200 2.4165 15.2460 3.5100 ;
      RECT 15.1120 2.4165 15.1380 3.5100 ;
      RECT 15.0040 2.4165 15.0300 3.5100 ;
      RECT 14.8960 2.4165 14.9220 3.5100 ;
      RECT 14.7880 2.4165 14.8140 3.5100 ;
      RECT 14.6800 2.4165 14.7060 3.5100 ;
      RECT 14.5720 2.4165 14.5980 3.5100 ;
      RECT 14.4640 2.4165 14.4900 3.5100 ;
      RECT 14.3560 2.4165 14.3820 3.5100 ;
      RECT 14.2480 2.4165 14.2740 3.5100 ;
      RECT 14.1400 2.4165 14.1660 3.5100 ;
      RECT 14.0320 2.4165 14.0580 3.5100 ;
      RECT 13.9240 2.4165 13.9500 3.5100 ;
      RECT 13.8160 2.4165 13.8420 3.5100 ;
      RECT 13.7080 2.4165 13.7340 3.5100 ;
      RECT 13.6000 2.4165 13.6260 3.5100 ;
      RECT 13.4920 2.4165 13.5180 3.5100 ;
      RECT 13.3840 2.4165 13.4100 3.5100 ;
      RECT 13.2760 2.4165 13.3020 3.5100 ;
      RECT 13.1680 2.4165 13.1940 3.5100 ;
      RECT 13.0600 2.4165 13.0860 3.5100 ;
      RECT 12.9520 2.4165 12.9780 3.5100 ;
      RECT 12.8440 2.4165 12.8700 3.5100 ;
      RECT 12.7360 2.4165 12.7620 3.5100 ;
      RECT 12.6280 2.4165 12.6540 3.5100 ;
      RECT 12.5200 2.4165 12.5460 3.5100 ;
      RECT 12.4120 2.4165 12.4380 3.5100 ;
      RECT 12.3040 2.4165 12.3300 3.5100 ;
      RECT 12.1960 2.4165 12.2220 3.5100 ;
      RECT 12.0880 2.4165 12.1140 3.5100 ;
      RECT 11.9800 2.4165 12.0060 3.5100 ;
      RECT 11.8720 2.4165 11.8980 3.5100 ;
      RECT 11.7640 2.4165 11.7900 3.5100 ;
      RECT 11.6560 2.4165 11.6820 3.5100 ;
      RECT 11.5480 2.4165 11.5740 3.5100 ;
      RECT 11.4400 2.4165 11.4660 3.5100 ;
      RECT 11.3320 2.4165 11.3580 3.5100 ;
      RECT 11.2240 2.4165 11.2500 3.5100 ;
      RECT 11.1160 2.4165 11.1420 3.5100 ;
      RECT 11.0080 2.4165 11.0340 3.5100 ;
      RECT 10.9000 2.4165 10.9260 3.5100 ;
      RECT 10.7920 2.4165 10.8180 3.5100 ;
      RECT 10.6840 2.4165 10.7100 3.5100 ;
      RECT 10.5760 2.4165 10.6020 3.5100 ;
      RECT 10.4680 2.4165 10.4940 3.5100 ;
      RECT 10.3600 2.4165 10.3860 3.5100 ;
      RECT 10.2520 2.4165 10.2780 3.5100 ;
      RECT 10.1440 2.4165 10.1700 3.5100 ;
      RECT 10.0360 2.4165 10.0620 3.5100 ;
      RECT 9.9280 2.4165 9.9540 3.5100 ;
      RECT 9.8200 2.4165 9.8460 3.5100 ;
      RECT 9.7120 2.4165 9.7380 3.5100 ;
      RECT 9.6040 2.4165 9.6300 3.5100 ;
      RECT 9.4960 2.4165 9.5220 3.5100 ;
      RECT 9.3880 2.4165 9.4140 3.5100 ;
      RECT 9.1750 2.4165 9.2520 3.5100 ;
      RECT 7.2820 2.4165 7.3590 3.5100 ;
      RECT 7.1200 2.4165 7.1460 3.5100 ;
      RECT 7.0120 2.4165 7.0380 3.5100 ;
      RECT 6.9040 2.4165 6.9300 3.5100 ;
      RECT 6.7960 2.4165 6.8220 3.5100 ;
      RECT 6.6880 2.4165 6.7140 3.5100 ;
      RECT 6.5800 2.4165 6.6060 3.5100 ;
      RECT 6.4720 2.4165 6.4980 3.5100 ;
      RECT 6.3640 2.4165 6.3900 3.5100 ;
      RECT 6.2560 2.4165 6.2820 3.5100 ;
      RECT 6.1480 2.4165 6.1740 3.5100 ;
      RECT 6.0400 2.4165 6.0660 3.5100 ;
      RECT 5.9320 2.4165 5.9580 3.5100 ;
      RECT 5.8240 2.4165 5.8500 3.5100 ;
      RECT 5.7160 2.4165 5.7420 3.5100 ;
      RECT 5.6080 2.4165 5.6340 3.5100 ;
      RECT 5.5000 2.4165 5.5260 3.5100 ;
      RECT 5.3920 2.4165 5.4180 3.5100 ;
      RECT 5.2840 2.4165 5.3100 3.5100 ;
      RECT 5.1760 2.4165 5.2020 3.5100 ;
      RECT 5.0680 2.4165 5.0940 3.5100 ;
      RECT 4.9600 2.4165 4.9860 3.5100 ;
      RECT 4.8520 2.4165 4.8780 3.5100 ;
      RECT 4.7440 2.4165 4.7700 3.5100 ;
      RECT 4.6360 2.4165 4.6620 3.5100 ;
      RECT 4.5280 2.4165 4.5540 3.5100 ;
      RECT 4.4200 2.4165 4.4460 3.5100 ;
      RECT 4.3120 2.4165 4.3380 3.5100 ;
      RECT 4.2040 2.4165 4.2300 3.5100 ;
      RECT 4.0960 2.4165 4.1220 3.5100 ;
      RECT 3.9880 2.4165 4.0140 3.5100 ;
      RECT 3.8800 2.4165 3.9060 3.5100 ;
      RECT 3.7720 2.4165 3.7980 3.5100 ;
      RECT 3.6640 2.4165 3.6900 3.5100 ;
      RECT 3.5560 2.4165 3.5820 3.5100 ;
      RECT 3.4480 2.4165 3.4740 3.5100 ;
      RECT 3.3400 2.4165 3.3660 3.5100 ;
      RECT 3.2320 2.4165 3.2580 3.5100 ;
      RECT 3.1240 2.4165 3.1500 3.5100 ;
      RECT 3.0160 2.4165 3.0420 3.5100 ;
      RECT 2.9080 2.4165 2.9340 3.5100 ;
      RECT 2.8000 2.4165 2.8260 3.5100 ;
      RECT 2.6920 2.4165 2.7180 3.5100 ;
      RECT 2.5840 2.4165 2.6100 3.5100 ;
      RECT 2.4760 2.4165 2.5020 3.5100 ;
      RECT 2.3680 2.4165 2.3940 3.5100 ;
      RECT 2.2600 2.4165 2.2860 3.5100 ;
      RECT 2.1520 2.4165 2.1780 3.5100 ;
      RECT 2.0440 2.4165 2.0700 3.5100 ;
      RECT 1.9360 2.4165 1.9620 3.5100 ;
      RECT 1.8280 2.4165 1.8540 3.5100 ;
      RECT 1.7200 2.4165 1.7460 3.5100 ;
      RECT 1.6120 2.4165 1.6380 3.5100 ;
      RECT 1.5040 2.4165 1.5300 3.5100 ;
      RECT 1.3960 2.4165 1.4220 3.5100 ;
      RECT 1.2880 2.4165 1.3140 3.5100 ;
      RECT 1.1800 2.4165 1.2060 3.5100 ;
      RECT 1.0720 2.4165 1.0980 3.5100 ;
      RECT 0.9640 2.4165 0.9900 3.5100 ;
      RECT 0.8560 2.4165 0.8820 3.5100 ;
      RECT 0.7480 2.4165 0.7740 3.5100 ;
      RECT 0.6400 2.4165 0.6660 3.5100 ;
      RECT 0.5320 2.4165 0.5580 3.5100 ;
      RECT 0.4240 2.4165 0.4500 3.5100 ;
      RECT 0.3160 2.4165 0.3420 3.5100 ;
      RECT 0.2080 2.4165 0.2340 3.5100 ;
      RECT 0.0050 2.4165 0.0900 3.5100 ;
      RECT 8.6410 3.4965 8.7690 4.5900 ;
      RECT 8.6270 4.1620 8.7690 4.4845 ;
      RECT 8.4790 3.8890 8.5410 4.5900 ;
      RECT 8.4650 4.1985 8.5410 4.3520 ;
      RECT 8.4790 3.4965 8.5050 4.5900 ;
      RECT 8.4790 3.6175 8.5190 3.8570 ;
      RECT 8.4790 3.4965 8.5410 3.5855 ;
      RECT 8.1820 3.9470 8.3880 4.5900 ;
      RECT 8.3620 3.4965 8.3880 4.5900 ;
      RECT 8.1820 4.2240 8.4020 4.4820 ;
      RECT 8.1820 3.4965 8.2800 4.5900 ;
      RECT 7.7650 3.4965 7.8480 4.5900 ;
      RECT 7.7650 3.5850 7.8620 4.5205 ;
      RECT 16.4440 3.4965 16.5290 4.5900 ;
      RECT 16.3000 3.4965 16.3260 4.5900 ;
      RECT 16.1920 3.4965 16.2180 4.5900 ;
      RECT 16.0840 3.4965 16.1100 4.5900 ;
      RECT 15.9760 3.4965 16.0020 4.5900 ;
      RECT 15.8680 3.4965 15.8940 4.5900 ;
      RECT 15.7600 3.4965 15.7860 4.5900 ;
      RECT 15.6520 3.4965 15.6780 4.5900 ;
      RECT 15.5440 3.4965 15.5700 4.5900 ;
      RECT 15.4360 3.4965 15.4620 4.5900 ;
      RECT 15.3280 3.4965 15.3540 4.5900 ;
      RECT 15.2200 3.4965 15.2460 4.5900 ;
      RECT 15.1120 3.4965 15.1380 4.5900 ;
      RECT 15.0040 3.4965 15.0300 4.5900 ;
      RECT 14.8960 3.4965 14.9220 4.5900 ;
      RECT 14.7880 3.4965 14.8140 4.5900 ;
      RECT 14.6800 3.4965 14.7060 4.5900 ;
      RECT 14.5720 3.4965 14.5980 4.5900 ;
      RECT 14.4640 3.4965 14.4900 4.5900 ;
      RECT 14.3560 3.4965 14.3820 4.5900 ;
      RECT 14.2480 3.4965 14.2740 4.5900 ;
      RECT 14.1400 3.4965 14.1660 4.5900 ;
      RECT 14.0320 3.4965 14.0580 4.5900 ;
      RECT 13.9240 3.4965 13.9500 4.5900 ;
      RECT 13.8160 3.4965 13.8420 4.5900 ;
      RECT 13.7080 3.4965 13.7340 4.5900 ;
      RECT 13.6000 3.4965 13.6260 4.5900 ;
      RECT 13.4920 3.4965 13.5180 4.5900 ;
      RECT 13.3840 3.4965 13.4100 4.5900 ;
      RECT 13.2760 3.4965 13.3020 4.5900 ;
      RECT 13.1680 3.4965 13.1940 4.5900 ;
      RECT 13.0600 3.4965 13.0860 4.5900 ;
      RECT 12.9520 3.4965 12.9780 4.5900 ;
      RECT 12.8440 3.4965 12.8700 4.5900 ;
      RECT 12.7360 3.4965 12.7620 4.5900 ;
      RECT 12.6280 3.4965 12.6540 4.5900 ;
      RECT 12.5200 3.4965 12.5460 4.5900 ;
      RECT 12.4120 3.4965 12.4380 4.5900 ;
      RECT 12.3040 3.4965 12.3300 4.5900 ;
      RECT 12.1960 3.4965 12.2220 4.5900 ;
      RECT 12.0880 3.4965 12.1140 4.5900 ;
      RECT 11.9800 3.4965 12.0060 4.5900 ;
      RECT 11.8720 3.4965 11.8980 4.5900 ;
      RECT 11.7640 3.4965 11.7900 4.5900 ;
      RECT 11.6560 3.4965 11.6820 4.5900 ;
      RECT 11.5480 3.4965 11.5740 4.5900 ;
      RECT 11.4400 3.4965 11.4660 4.5900 ;
      RECT 11.3320 3.4965 11.3580 4.5900 ;
      RECT 11.2240 3.4965 11.2500 4.5900 ;
      RECT 11.1160 3.4965 11.1420 4.5900 ;
      RECT 11.0080 3.4965 11.0340 4.5900 ;
      RECT 10.9000 3.4965 10.9260 4.5900 ;
      RECT 10.7920 3.4965 10.8180 4.5900 ;
      RECT 10.6840 3.4965 10.7100 4.5900 ;
      RECT 10.5760 3.4965 10.6020 4.5900 ;
      RECT 10.4680 3.4965 10.4940 4.5900 ;
      RECT 10.3600 3.4965 10.3860 4.5900 ;
      RECT 10.2520 3.4965 10.2780 4.5900 ;
      RECT 10.1440 3.4965 10.1700 4.5900 ;
      RECT 10.0360 3.4965 10.0620 4.5900 ;
      RECT 9.9280 3.4965 9.9540 4.5900 ;
      RECT 9.8200 3.4965 9.8460 4.5900 ;
      RECT 9.7120 3.4965 9.7380 4.5900 ;
      RECT 9.6040 3.4965 9.6300 4.5900 ;
      RECT 9.4960 3.4965 9.5220 4.5900 ;
      RECT 9.3880 3.4965 9.4140 4.5900 ;
      RECT 9.1750 3.4965 9.2520 4.5900 ;
      RECT 7.2820 3.4965 7.3590 4.5900 ;
      RECT 7.1200 3.4965 7.1460 4.5900 ;
      RECT 7.0120 3.4965 7.0380 4.5900 ;
      RECT 6.9040 3.4965 6.9300 4.5900 ;
      RECT 6.7960 3.4965 6.8220 4.5900 ;
      RECT 6.6880 3.4965 6.7140 4.5900 ;
      RECT 6.5800 3.4965 6.6060 4.5900 ;
      RECT 6.4720 3.4965 6.4980 4.5900 ;
      RECT 6.3640 3.4965 6.3900 4.5900 ;
      RECT 6.2560 3.4965 6.2820 4.5900 ;
      RECT 6.1480 3.4965 6.1740 4.5900 ;
      RECT 6.0400 3.4965 6.0660 4.5900 ;
      RECT 5.9320 3.4965 5.9580 4.5900 ;
      RECT 5.8240 3.4965 5.8500 4.5900 ;
      RECT 5.7160 3.4965 5.7420 4.5900 ;
      RECT 5.6080 3.4965 5.6340 4.5900 ;
      RECT 5.5000 3.4965 5.5260 4.5900 ;
      RECT 5.3920 3.4965 5.4180 4.5900 ;
      RECT 5.2840 3.4965 5.3100 4.5900 ;
      RECT 5.1760 3.4965 5.2020 4.5900 ;
      RECT 5.0680 3.4965 5.0940 4.5900 ;
      RECT 4.9600 3.4965 4.9860 4.5900 ;
      RECT 4.8520 3.4965 4.8780 4.5900 ;
      RECT 4.7440 3.4965 4.7700 4.5900 ;
      RECT 4.6360 3.4965 4.6620 4.5900 ;
      RECT 4.5280 3.4965 4.5540 4.5900 ;
      RECT 4.4200 3.4965 4.4460 4.5900 ;
      RECT 4.3120 3.4965 4.3380 4.5900 ;
      RECT 4.2040 3.4965 4.2300 4.5900 ;
      RECT 4.0960 3.4965 4.1220 4.5900 ;
      RECT 3.9880 3.4965 4.0140 4.5900 ;
      RECT 3.8800 3.4965 3.9060 4.5900 ;
      RECT 3.7720 3.4965 3.7980 4.5900 ;
      RECT 3.6640 3.4965 3.6900 4.5900 ;
      RECT 3.5560 3.4965 3.5820 4.5900 ;
      RECT 3.4480 3.4965 3.4740 4.5900 ;
      RECT 3.3400 3.4965 3.3660 4.5900 ;
      RECT 3.2320 3.4965 3.2580 4.5900 ;
      RECT 3.1240 3.4965 3.1500 4.5900 ;
      RECT 3.0160 3.4965 3.0420 4.5900 ;
      RECT 2.9080 3.4965 2.9340 4.5900 ;
      RECT 2.8000 3.4965 2.8260 4.5900 ;
      RECT 2.6920 3.4965 2.7180 4.5900 ;
      RECT 2.5840 3.4965 2.6100 4.5900 ;
      RECT 2.4760 3.4965 2.5020 4.5900 ;
      RECT 2.3680 3.4965 2.3940 4.5900 ;
      RECT 2.2600 3.4965 2.2860 4.5900 ;
      RECT 2.1520 3.4965 2.1780 4.5900 ;
      RECT 2.0440 3.4965 2.0700 4.5900 ;
      RECT 1.9360 3.4965 1.9620 4.5900 ;
      RECT 1.8280 3.4965 1.8540 4.5900 ;
      RECT 1.7200 3.4965 1.7460 4.5900 ;
      RECT 1.6120 3.4965 1.6380 4.5900 ;
      RECT 1.5040 3.4965 1.5300 4.5900 ;
      RECT 1.3960 3.4965 1.4220 4.5900 ;
      RECT 1.2880 3.4965 1.3140 4.5900 ;
      RECT 1.1800 3.4965 1.2060 4.5900 ;
      RECT 1.0720 3.4965 1.0980 4.5900 ;
      RECT 0.9640 3.4965 0.9900 4.5900 ;
      RECT 0.8560 3.4965 0.8820 4.5900 ;
      RECT 0.7480 3.4965 0.7740 4.5900 ;
      RECT 0.6400 3.4965 0.6660 4.5900 ;
      RECT 0.5320 3.4965 0.5580 4.5900 ;
      RECT 0.4240 3.4965 0.4500 4.5900 ;
      RECT 0.3160 3.4965 0.3420 4.5900 ;
      RECT 0.2080 3.4965 0.2340 4.5900 ;
      RECT 0.0050 3.4965 0.0900 4.5900 ;
      RECT 8.6410 4.5765 8.7690 5.6700 ;
      RECT 8.6270 5.2420 8.7690 5.5645 ;
      RECT 8.4790 4.9690 8.5410 5.6700 ;
      RECT 8.4650 5.2785 8.5410 5.4320 ;
      RECT 8.4790 4.5765 8.5050 5.6700 ;
      RECT 8.4790 4.6975 8.5190 4.9370 ;
      RECT 8.4790 4.5765 8.5410 4.6655 ;
      RECT 8.1820 5.0270 8.3880 5.6700 ;
      RECT 8.3620 4.5765 8.3880 5.6700 ;
      RECT 8.1820 5.3040 8.4020 5.5620 ;
      RECT 8.1820 4.5765 8.2800 5.6700 ;
      RECT 7.7650 4.5765 7.8480 5.6700 ;
      RECT 7.7650 4.6650 7.8620 5.6005 ;
      RECT 16.4440 4.5765 16.5290 5.6700 ;
      RECT 16.3000 4.5765 16.3260 5.6700 ;
      RECT 16.1920 4.5765 16.2180 5.6700 ;
      RECT 16.0840 4.5765 16.1100 5.6700 ;
      RECT 15.9760 4.5765 16.0020 5.6700 ;
      RECT 15.8680 4.5765 15.8940 5.6700 ;
      RECT 15.7600 4.5765 15.7860 5.6700 ;
      RECT 15.6520 4.5765 15.6780 5.6700 ;
      RECT 15.5440 4.5765 15.5700 5.6700 ;
      RECT 15.4360 4.5765 15.4620 5.6700 ;
      RECT 15.3280 4.5765 15.3540 5.6700 ;
      RECT 15.2200 4.5765 15.2460 5.6700 ;
      RECT 15.1120 4.5765 15.1380 5.6700 ;
      RECT 15.0040 4.5765 15.0300 5.6700 ;
      RECT 14.8960 4.5765 14.9220 5.6700 ;
      RECT 14.7880 4.5765 14.8140 5.6700 ;
      RECT 14.6800 4.5765 14.7060 5.6700 ;
      RECT 14.5720 4.5765 14.5980 5.6700 ;
      RECT 14.4640 4.5765 14.4900 5.6700 ;
      RECT 14.3560 4.5765 14.3820 5.6700 ;
      RECT 14.2480 4.5765 14.2740 5.6700 ;
      RECT 14.1400 4.5765 14.1660 5.6700 ;
      RECT 14.0320 4.5765 14.0580 5.6700 ;
      RECT 13.9240 4.5765 13.9500 5.6700 ;
      RECT 13.8160 4.5765 13.8420 5.6700 ;
      RECT 13.7080 4.5765 13.7340 5.6700 ;
      RECT 13.6000 4.5765 13.6260 5.6700 ;
      RECT 13.4920 4.5765 13.5180 5.6700 ;
      RECT 13.3840 4.5765 13.4100 5.6700 ;
      RECT 13.2760 4.5765 13.3020 5.6700 ;
      RECT 13.1680 4.5765 13.1940 5.6700 ;
      RECT 13.0600 4.5765 13.0860 5.6700 ;
      RECT 12.9520 4.5765 12.9780 5.6700 ;
      RECT 12.8440 4.5765 12.8700 5.6700 ;
      RECT 12.7360 4.5765 12.7620 5.6700 ;
      RECT 12.6280 4.5765 12.6540 5.6700 ;
      RECT 12.5200 4.5765 12.5460 5.6700 ;
      RECT 12.4120 4.5765 12.4380 5.6700 ;
      RECT 12.3040 4.5765 12.3300 5.6700 ;
      RECT 12.1960 4.5765 12.2220 5.6700 ;
      RECT 12.0880 4.5765 12.1140 5.6700 ;
      RECT 11.9800 4.5765 12.0060 5.6700 ;
      RECT 11.8720 4.5765 11.8980 5.6700 ;
      RECT 11.7640 4.5765 11.7900 5.6700 ;
      RECT 11.6560 4.5765 11.6820 5.6700 ;
      RECT 11.5480 4.5765 11.5740 5.6700 ;
      RECT 11.4400 4.5765 11.4660 5.6700 ;
      RECT 11.3320 4.5765 11.3580 5.6700 ;
      RECT 11.2240 4.5765 11.2500 5.6700 ;
      RECT 11.1160 4.5765 11.1420 5.6700 ;
      RECT 11.0080 4.5765 11.0340 5.6700 ;
      RECT 10.9000 4.5765 10.9260 5.6700 ;
      RECT 10.7920 4.5765 10.8180 5.6700 ;
      RECT 10.6840 4.5765 10.7100 5.6700 ;
      RECT 10.5760 4.5765 10.6020 5.6700 ;
      RECT 10.4680 4.5765 10.4940 5.6700 ;
      RECT 10.3600 4.5765 10.3860 5.6700 ;
      RECT 10.2520 4.5765 10.2780 5.6700 ;
      RECT 10.1440 4.5765 10.1700 5.6700 ;
      RECT 10.0360 4.5765 10.0620 5.6700 ;
      RECT 9.9280 4.5765 9.9540 5.6700 ;
      RECT 9.8200 4.5765 9.8460 5.6700 ;
      RECT 9.7120 4.5765 9.7380 5.6700 ;
      RECT 9.6040 4.5765 9.6300 5.6700 ;
      RECT 9.4960 4.5765 9.5220 5.6700 ;
      RECT 9.3880 4.5765 9.4140 5.6700 ;
      RECT 9.1750 4.5765 9.2520 5.6700 ;
      RECT 7.2820 4.5765 7.3590 5.6700 ;
      RECT 7.1200 4.5765 7.1460 5.6700 ;
      RECT 7.0120 4.5765 7.0380 5.6700 ;
      RECT 6.9040 4.5765 6.9300 5.6700 ;
      RECT 6.7960 4.5765 6.8220 5.6700 ;
      RECT 6.6880 4.5765 6.7140 5.6700 ;
      RECT 6.5800 4.5765 6.6060 5.6700 ;
      RECT 6.4720 4.5765 6.4980 5.6700 ;
      RECT 6.3640 4.5765 6.3900 5.6700 ;
      RECT 6.2560 4.5765 6.2820 5.6700 ;
      RECT 6.1480 4.5765 6.1740 5.6700 ;
      RECT 6.0400 4.5765 6.0660 5.6700 ;
      RECT 5.9320 4.5765 5.9580 5.6700 ;
      RECT 5.8240 4.5765 5.8500 5.6700 ;
      RECT 5.7160 4.5765 5.7420 5.6700 ;
      RECT 5.6080 4.5765 5.6340 5.6700 ;
      RECT 5.5000 4.5765 5.5260 5.6700 ;
      RECT 5.3920 4.5765 5.4180 5.6700 ;
      RECT 5.2840 4.5765 5.3100 5.6700 ;
      RECT 5.1760 4.5765 5.2020 5.6700 ;
      RECT 5.0680 4.5765 5.0940 5.6700 ;
      RECT 4.9600 4.5765 4.9860 5.6700 ;
      RECT 4.8520 4.5765 4.8780 5.6700 ;
      RECT 4.7440 4.5765 4.7700 5.6700 ;
      RECT 4.6360 4.5765 4.6620 5.6700 ;
      RECT 4.5280 4.5765 4.5540 5.6700 ;
      RECT 4.4200 4.5765 4.4460 5.6700 ;
      RECT 4.3120 4.5765 4.3380 5.6700 ;
      RECT 4.2040 4.5765 4.2300 5.6700 ;
      RECT 4.0960 4.5765 4.1220 5.6700 ;
      RECT 3.9880 4.5765 4.0140 5.6700 ;
      RECT 3.8800 4.5765 3.9060 5.6700 ;
      RECT 3.7720 4.5765 3.7980 5.6700 ;
      RECT 3.6640 4.5765 3.6900 5.6700 ;
      RECT 3.5560 4.5765 3.5820 5.6700 ;
      RECT 3.4480 4.5765 3.4740 5.6700 ;
      RECT 3.3400 4.5765 3.3660 5.6700 ;
      RECT 3.2320 4.5765 3.2580 5.6700 ;
      RECT 3.1240 4.5765 3.1500 5.6700 ;
      RECT 3.0160 4.5765 3.0420 5.6700 ;
      RECT 2.9080 4.5765 2.9340 5.6700 ;
      RECT 2.8000 4.5765 2.8260 5.6700 ;
      RECT 2.6920 4.5765 2.7180 5.6700 ;
      RECT 2.5840 4.5765 2.6100 5.6700 ;
      RECT 2.4760 4.5765 2.5020 5.6700 ;
      RECT 2.3680 4.5765 2.3940 5.6700 ;
      RECT 2.2600 4.5765 2.2860 5.6700 ;
      RECT 2.1520 4.5765 2.1780 5.6700 ;
      RECT 2.0440 4.5765 2.0700 5.6700 ;
      RECT 1.9360 4.5765 1.9620 5.6700 ;
      RECT 1.8280 4.5765 1.8540 5.6700 ;
      RECT 1.7200 4.5765 1.7460 5.6700 ;
      RECT 1.6120 4.5765 1.6380 5.6700 ;
      RECT 1.5040 4.5765 1.5300 5.6700 ;
      RECT 1.3960 4.5765 1.4220 5.6700 ;
      RECT 1.2880 4.5765 1.3140 5.6700 ;
      RECT 1.1800 4.5765 1.2060 5.6700 ;
      RECT 1.0720 4.5765 1.0980 5.6700 ;
      RECT 0.9640 4.5765 0.9900 5.6700 ;
      RECT 0.8560 4.5765 0.8820 5.6700 ;
      RECT 0.7480 4.5765 0.7740 5.6700 ;
      RECT 0.6400 4.5765 0.6660 5.6700 ;
      RECT 0.5320 4.5765 0.5580 5.6700 ;
      RECT 0.4240 4.5765 0.4500 5.6700 ;
      RECT 0.3160 4.5765 0.3420 5.6700 ;
      RECT 0.2080 4.5765 0.2340 5.6700 ;
      RECT 0.0050 4.5765 0.0900 5.6700 ;
      RECT 8.6410 5.6565 8.7690 6.7500 ;
      RECT 8.6270 6.3220 8.7690 6.6445 ;
      RECT 8.4790 6.0490 8.5410 6.7500 ;
      RECT 8.4650 6.3585 8.5410 6.5120 ;
      RECT 8.4790 5.6565 8.5050 6.7500 ;
      RECT 8.4790 5.7775 8.5190 6.0170 ;
      RECT 8.4790 5.6565 8.5410 5.7455 ;
      RECT 8.1820 6.1070 8.3880 6.7500 ;
      RECT 8.3620 5.6565 8.3880 6.7500 ;
      RECT 8.1820 6.3840 8.4020 6.6420 ;
      RECT 8.1820 5.6565 8.2800 6.7500 ;
      RECT 7.7650 5.6565 7.8480 6.7500 ;
      RECT 7.7650 5.7450 7.8620 6.6805 ;
      RECT 16.4440 5.6565 16.5290 6.7500 ;
      RECT 16.3000 5.6565 16.3260 6.7500 ;
      RECT 16.1920 5.6565 16.2180 6.7500 ;
      RECT 16.0840 5.6565 16.1100 6.7500 ;
      RECT 15.9760 5.6565 16.0020 6.7500 ;
      RECT 15.8680 5.6565 15.8940 6.7500 ;
      RECT 15.7600 5.6565 15.7860 6.7500 ;
      RECT 15.6520 5.6565 15.6780 6.7500 ;
      RECT 15.5440 5.6565 15.5700 6.7500 ;
      RECT 15.4360 5.6565 15.4620 6.7500 ;
      RECT 15.3280 5.6565 15.3540 6.7500 ;
      RECT 15.2200 5.6565 15.2460 6.7500 ;
      RECT 15.1120 5.6565 15.1380 6.7500 ;
      RECT 15.0040 5.6565 15.0300 6.7500 ;
      RECT 14.8960 5.6565 14.9220 6.7500 ;
      RECT 14.7880 5.6565 14.8140 6.7500 ;
      RECT 14.6800 5.6565 14.7060 6.7500 ;
      RECT 14.5720 5.6565 14.5980 6.7500 ;
      RECT 14.4640 5.6565 14.4900 6.7500 ;
      RECT 14.3560 5.6565 14.3820 6.7500 ;
      RECT 14.2480 5.6565 14.2740 6.7500 ;
      RECT 14.1400 5.6565 14.1660 6.7500 ;
      RECT 14.0320 5.6565 14.0580 6.7500 ;
      RECT 13.9240 5.6565 13.9500 6.7500 ;
      RECT 13.8160 5.6565 13.8420 6.7500 ;
      RECT 13.7080 5.6565 13.7340 6.7500 ;
      RECT 13.6000 5.6565 13.6260 6.7500 ;
      RECT 13.4920 5.6565 13.5180 6.7500 ;
      RECT 13.3840 5.6565 13.4100 6.7500 ;
      RECT 13.2760 5.6565 13.3020 6.7500 ;
      RECT 13.1680 5.6565 13.1940 6.7500 ;
      RECT 13.0600 5.6565 13.0860 6.7500 ;
      RECT 12.9520 5.6565 12.9780 6.7500 ;
      RECT 12.8440 5.6565 12.8700 6.7500 ;
      RECT 12.7360 5.6565 12.7620 6.7500 ;
      RECT 12.6280 5.6565 12.6540 6.7500 ;
      RECT 12.5200 5.6565 12.5460 6.7500 ;
      RECT 12.4120 5.6565 12.4380 6.7500 ;
      RECT 12.3040 5.6565 12.3300 6.7500 ;
      RECT 12.1960 5.6565 12.2220 6.7500 ;
      RECT 12.0880 5.6565 12.1140 6.7500 ;
      RECT 11.9800 5.6565 12.0060 6.7500 ;
      RECT 11.8720 5.6565 11.8980 6.7500 ;
      RECT 11.7640 5.6565 11.7900 6.7500 ;
      RECT 11.6560 5.6565 11.6820 6.7500 ;
      RECT 11.5480 5.6565 11.5740 6.7500 ;
      RECT 11.4400 5.6565 11.4660 6.7500 ;
      RECT 11.3320 5.6565 11.3580 6.7500 ;
      RECT 11.2240 5.6565 11.2500 6.7500 ;
      RECT 11.1160 5.6565 11.1420 6.7500 ;
      RECT 11.0080 5.6565 11.0340 6.7500 ;
      RECT 10.9000 5.6565 10.9260 6.7500 ;
      RECT 10.7920 5.6565 10.8180 6.7500 ;
      RECT 10.6840 5.6565 10.7100 6.7500 ;
      RECT 10.5760 5.6565 10.6020 6.7500 ;
      RECT 10.4680 5.6565 10.4940 6.7500 ;
      RECT 10.3600 5.6565 10.3860 6.7500 ;
      RECT 10.2520 5.6565 10.2780 6.7500 ;
      RECT 10.1440 5.6565 10.1700 6.7500 ;
      RECT 10.0360 5.6565 10.0620 6.7500 ;
      RECT 9.9280 5.6565 9.9540 6.7500 ;
      RECT 9.8200 5.6565 9.8460 6.7500 ;
      RECT 9.7120 5.6565 9.7380 6.7500 ;
      RECT 9.6040 5.6565 9.6300 6.7500 ;
      RECT 9.4960 5.6565 9.5220 6.7500 ;
      RECT 9.3880 5.6565 9.4140 6.7500 ;
      RECT 9.1750 5.6565 9.2520 6.7500 ;
      RECT 7.2820 5.6565 7.3590 6.7500 ;
      RECT 7.1200 5.6565 7.1460 6.7500 ;
      RECT 7.0120 5.6565 7.0380 6.7500 ;
      RECT 6.9040 5.6565 6.9300 6.7500 ;
      RECT 6.7960 5.6565 6.8220 6.7500 ;
      RECT 6.6880 5.6565 6.7140 6.7500 ;
      RECT 6.5800 5.6565 6.6060 6.7500 ;
      RECT 6.4720 5.6565 6.4980 6.7500 ;
      RECT 6.3640 5.6565 6.3900 6.7500 ;
      RECT 6.2560 5.6565 6.2820 6.7500 ;
      RECT 6.1480 5.6565 6.1740 6.7500 ;
      RECT 6.0400 5.6565 6.0660 6.7500 ;
      RECT 5.9320 5.6565 5.9580 6.7500 ;
      RECT 5.8240 5.6565 5.8500 6.7500 ;
      RECT 5.7160 5.6565 5.7420 6.7500 ;
      RECT 5.6080 5.6565 5.6340 6.7500 ;
      RECT 5.5000 5.6565 5.5260 6.7500 ;
      RECT 5.3920 5.6565 5.4180 6.7500 ;
      RECT 5.2840 5.6565 5.3100 6.7500 ;
      RECT 5.1760 5.6565 5.2020 6.7500 ;
      RECT 5.0680 5.6565 5.0940 6.7500 ;
      RECT 4.9600 5.6565 4.9860 6.7500 ;
      RECT 4.8520 5.6565 4.8780 6.7500 ;
      RECT 4.7440 5.6565 4.7700 6.7500 ;
      RECT 4.6360 5.6565 4.6620 6.7500 ;
      RECT 4.5280 5.6565 4.5540 6.7500 ;
      RECT 4.4200 5.6565 4.4460 6.7500 ;
      RECT 4.3120 5.6565 4.3380 6.7500 ;
      RECT 4.2040 5.6565 4.2300 6.7500 ;
      RECT 4.0960 5.6565 4.1220 6.7500 ;
      RECT 3.9880 5.6565 4.0140 6.7500 ;
      RECT 3.8800 5.6565 3.9060 6.7500 ;
      RECT 3.7720 5.6565 3.7980 6.7500 ;
      RECT 3.6640 5.6565 3.6900 6.7500 ;
      RECT 3.5560 5.6565 3.5820 6.7500 ;
      RECT 3.4480 5.6565 3.4740 6.7500 ;
      RECT 3.3400 5.6565 3.3660 6.7500 ;
      RECT 3.2320 5.6565 3.2580 6.7500 ;
      RECT 3.1240 5.6565 3.1500 6.7500 ;
      RECT 3.0160 5.6565 3.0420 6.7500 ;
      RECT 2.9080 5.6565 2.9340 6.7500 ;
      RECT 2.8000 5.6565 2.8260 6.7500 ;
      RECT 2.6920 5.6565 2.7180 6.7500 ;
      RECT 2.5840 5.6565 2.6100 6.7500 ;
      RECT 2.4760 5.6565 2.5020 6.7500 ;
      RECT 2.3680 5.6565 2.3940 6.7500 ;
      RECT 2.2600 5.6565 2.2860 6.7500 ;
      RECT 2.1520 5.6565 2.1780 6.7500 ;
      RECT 2.0440 5.6565 2.0700 6.7500 ;
      RECT 1.9360 5.6565 1.9620 6.7500 ;
      RECT 1.8280 5.6565 1.8540 6.7500 ;
      RECT 1.7200 5.6565 1.7460 6.7500 ;
      RECT 1.6120 5.6565 1.6380 6.7500 ;
      RECT 1.5040 5.6565 1.5300 6.7500 ;
      RECT 1.3960 5.6565 1.4220 6.7500 ;
      RECT 1.2880 5.6565 1.3140 6.7500 ;
      RECT 1.1800 5.6565 1.2060 6.7500 ;
      RECT 1.0720 5.6565 1.0980 6.7500 ;
      RECT 0.9640 5.6565 0.9900 6.7500 ;
      RECT 0.8560 5.6565 0.8820 6.7500 ;
      RECT 0.7480 5.6565 0.7740 6.7500 ;
      RECT 0.6400 5.6565 0.6660 6.7500 ;
      RECT 0.5320 5.6565 0.5580 6.7500 ;
      RECT 0.4240 5.6565 0.4500 6.7500 ;
      RECT 0.3160 5.6565 0.3420 6.7500 ;
      RECT 0.2080 5.6565 0.2340 6.7500 ;
      RECT 0.0050 5.6565 0.0900 6.7500 ;
      RECT 8.6410 6.7365 8.7690 7.8300 ;
      RECT 8.6270 7.4020 8.7690 7.7245 ;
      RECT 8.4790 7.1290 8.5410 7.8300 ;
      RECT 8.4650 7.4385 8.5410 7.5920 ;
      RECT 8.4790 6.7365 8.5050 7.8300 ;
      RECT 8.4790 6.8575 8.5190 7.0970 ;
      RECT 8.4790 6.7365 8.5410 6.8255 ;
      RECT 8.1820 7.1870 8.3880 7.8300 ;
      RECT 8.3620 6.7365 8.3880 7.8300 ;
      RECT 8.1820 7.4640 8.4020 7.7220 ;
      RECT 8.1820 6.7365 8.2800 7.8300 ;
      RECT 7.7650 6.7365 7.8480 7.8300 ;
      RECT 7.7650 6.8250 7.8620 7.7605 ;
      RECT 16.4440 6.7365 16.5290 7.8300 ;
      RECT 16.3000 6.7365 16.3260 7.8300 ;
      RECT 16.1920 6.7365 16.2180 7.8300 ;
      RECT 16.0840 6.7365 16.1100 7.8300 ;
      RECT 15.9760 6.7365 16.0020 7.8300 ;
      RECT 15.8680 6.7365 15.8940 7.8300 ;
      RECT 15.7600 6.7365 15.7860 7.8300 ;
      RECT 15.6520 6.7365 15.6780 7.8300 ;
      RECT 15.5440 6.7365 15.5700 7.8300 ;
      RECT 15.4360 6.7365 15.4620 7.8300 ;
      RECT 15.3280 6.7365 15.3540 7.8300 ;
      RECT 15.2200 6.7365 15.2460 7.8300 ;
      RECT 15.1120 6.7365 15.1380 7.8300 ;
      RECT 15.0040 6.7365 15.0300 7.8300 ;
      RECT 14.8960 6.7365 14.9220 7.8300 ;
      RECT 14.7880 6.7365 14.8140 7.8300 ;
      RECT 14.6800 6.7365 14.7060 7.8300 ;
      RECT 14.5720 6.7365 14.5980 7.8300 ;
      RECT 14.4640 6.7365 14.4900 7.8300 ;
      RECT 14.3560 6.7365 14.3820 7.8300 ;
      RECT 14.2480 6.7365 14.2740 7.8300 ;
      RECT 14.1400 6.7365 14.1660 7.8300 ;
      RECT 14.0320 6.7365 14.0580 7.8300 ;
      RECT 13.9240 6.7365 13.9500 7.8300 ;
      RECT 13.8160 6.7365 13.8420 7.8300 ;
      RECT 13.7080 6.7365 13.7340 7.8300 ;
      RECT 13.6000 6.7365 13.6260 7.8300 ;
      RECT 13.4920 6.7365 13.5180 7.8300 ;
      RECT 13.3840 6.7365 13.4100 7.8300 ;
      RECT 13.2760 6.7365 13.3020 7.8300 ;
      RECT 13.1680 6.7365 13.1940 7.8300 ;
      RECT 13.0600 6.7365 13.0860 7.8300 ;
      RECT 12.9520 6.7365 12.9780 7.8300 ;
      RECT 12.8440 6.7365 12.8700 7.8300 ;
      RECT 12.7360 6.7365 12.7620 7.8300 ;
      RECT 12.6280 6.7365 12.6540 7.8300 ;
      RECT 12.5200 6.7365 12.5460 7.8300 ;
      RECT 12.4120 6.7365 12.4380 7.8300 ;
      RECT 12.3040 6.7365 12.3300 7.8300 ;
      RECT 12.1960 6.7365 12.2220 7.8300 ;
      RECT 12.0880 6.7365 12.1140 7.8300 ;
      RECT 11.9800 6.7365 12.0060 7.8300 ;
      RECT 11.8720 6.7365 11.8980 7.8300 ;
      RECT 11.7640 6.7365 11.7900 7.8300 ;
      RECT 11.6560 6.7365 11.6820 7.8300 ;
      RECT 11.5480 6.7365 11.5740 7.8300 ;
      RECT 11.4400 6.7365 11.4660 7.8300 ;
      RECT 11.3320 6.7365 11.3580 7.8300 ;
      RECT 11.2240 6.7365 11.2500 7.8300 ;
      RECT 11.1160 6.7365 11.1420 7.8300 ;
      RECT 11.0080 6.7365 11.0340 7.8300 ;
      RECT 10.9000 6.7365 10.9260 7.8300 ;
      RECT 10.7920 6.7365 10.8180 7.8300 ;
      RECT 10.6840 6.7365 10.7100 7.8300 ;
      RECT 10.5760 6.7365 10.6020 7.8300 ;
      RECT 10.4680 6.7365 10.4940 7.8300 ;
      RECT 10.3600 6.7365 10.3860 7.8300 ;
      RECT 10.2520 6.7365 10.2780 7.8300 ;
      RECT 10.1440 6.7365 10.1700 7.8300 ;
      RECT 10.0360 6.7365 10.0620 7.8300 ;
      RECT 9.9280 6.7365 9.9540 7.8300 ;
      RECT 9.8200 6.7365 9.8460 7.8300 ;
      RECT 9.7120 6.7365 9.7380 7.8300 ;
      RECT 9.6040 6.7365 9.6300 7.8300 ;
      RECT 9.4960 6.7365 9.5220 7.8300 ;
      RECT 9.3880 6.7365 9.4140 7.8300 ;
      RECT 9.1750 6.7365 9.2520 7.8300 ;
      RECT 7.2820 6.7365 7.3590 7.8300 ;
      RECT 7.1200 6.7365 7.1460 7.8300 ;
      RECT 7.0120 6.7365 7.0380 7.8300 ;
      RECT 6.9040 6.7365 6.9300 7.8300 ;
      RECT 6.7960 6.7365 6.8220 7.8300 ;
      RECT 6.6880 6.7365 6.7140 7.8300 ;
      RECT 6.5800 6.7365 6.6060 7.8300 ;
      RECT 6.4720 6.7365 6.4980 7.8300 ;
      RECT 6.3640 6.7365 6.3900 7.8300 ;
      RECT 6.2560 6.7365 6.2820 7.8300 ;
      RECT 6.1480 6.7365 6.1740 7.8300 ;
      RECT 6.0400 6.7365 6.0660 7.8300 ;
      RECT 5.9320 6.7365 5.9580 7.8300 ;
      RECT 5.8240 6.7365 5.8500 7.8300 ;
      RECT 5.7160 6.7365 5.7420 7.8300 ;
      RECT 5.6080 6.7365 5.6340 7.8300 ;
      RECT 5.5000 6.7365 5.5260 7.8300 ;
      RECT 5.3920 6.7365 5.4180 7.8300 ;
      RECT 5.2840 6.7365 5.3100 7.8300 ;
      RECT 5.1760 6.7365 5.2020 7.8300 ;
      RECT 5.0680 6.7365 5.0940 7.8300 ;
      RECT 4.9600 6.7365 4.9860 7.8300 ;
      RECT 4.8520 6.7365 4.8780 7.8300 ;
      RECT 4.7440 6.7365 4.7700 7.8300 ;
      RECT 4.6360 6.7365 4.6620 7.8300 ;
      RECT 4.5280 6.7365 4.5540 7.8300 ;
      RECT 4.4200 6.7365 4.4460 7.8300 ;
      RECT 4.3120 6.7365 4.3380 7.8300 ;
      RECT 4.2040 6.7365 4.2300 7.8300 ;
      RECT 4.0960 6.7365 4.1220 7.8300 ;
      RECT 3.9880 6.7365 4.0140 7.8300 ;
      RECT 3.8800 6.7365 3.9060 7.8300 ;
      RECT 3.7720 6.7365 3.7980 7.8300 ;
      RECT 3.6640 6.7365 3.6900 7.8300 ;
      RECT 3.5560 6.7365 3.5820 7.8300 ;
      RECT 3.4480 6.7365 3.4740 7.8300 ;
      RECT 3.3400 6.7365 3.3660 7.8300 ;
      RECT 3.2320 6.7365 3.2580 7.8300 ;
      RECT 3.1240 6.7365 3.1500 7.8300 ;
      RECT 3.0160 6.7365 3.0420 7.8300 ;
      RECT 2.9080 6.7365 2.9340 7.8300 ;
      RECT 2.8000 6.7365 2.8260 7.8300 ;
      RECT 2.6920 6.7365 2.7180 7.8300 ;
      RECT 2.5840 6.7365 2.6100 7.8300 ;
      RECT 2.4760 6.7365 2.5020 7.8300 ;
      RECT 2.3680 6.7365 2.3940 7.8300 ;
      RECT 2.2600 6.7365 2.2860 7.8300 ;
      RECT 2.1520 6.7365 2.1780 7.8300 ;
      RECT 2.0440 6.7365 2.0700 7.8300 ;
      RECT 1.9360 6.7365 1.9620 7.8300 ;
      RECT 1.8280 6.7365 1.8540 7.8300 ;
      RECT 1.7200 6.7365 1.7460 7.8300 ;
      RECT 1.6120 6.7365 1.6380 7.8300 ;
      RECT 1.5040 6.7365 1.5300 7.8300 ;
      RECT 1.3960 6.7365 1.4220 7.8300 ;
      RECT 1.2880 6.7365 1.3140 7.8300 ;
      RECT 1.1800 6.7365 1.2060 7.8300 ;
      RECT 1.0720 6.7365 1.0980 7.8300 ;
      RECT 0.9640 6.7365 0.9900 7.8300 ;
      RECT 0.8560 6.7365 0.8820 7.8300 ;
      RECT 0.7480 6.7365 0.7740 7.8300 ;
      RECT 0.6400 6.7365 0.6660 7.8300 ;
      RECT 0.5320 6.7365 0.5580 7.8300 ;
      RECT 0.4240 6.7365 0.4500 7.8300 ;
      RECT 0.3160 6.7365 0.3420 7.8300 ;
      RECT 0.2080 6.7365 0.2340 7.8300 ;
      RECT 0.0050 6.7365 0.0900 7.8300 ;
      RECT 8.6410 7.8165 8.7690 8.9100 ;
      RECT 8.6270 8.4820 8.7690 8.8045 ;
      RECT 8.4790 8.2090 8.5410 8.9100 ;
      RECT 8.4650 8.5185 8.5410 8.6720 ;
      RECT 8.4790 7.8165 8.5050 8.9100 ;
      RECT 8.4790 7.9375 8.5190 8.1770 ;
      RECT 8.4790 7.8165 8.5410 7.9055 ;
      RECT 8.1820 8.2670 8.3880 8.9100 ;
      RECT 8.3620 7.8165 8.3880 8.9100 ;
      RECT 8.1820 8.5440 8.4020 8.8020 ;
      RECT 8.1820 7.8165 8.2800 8.9100 ;
      RECT 7.7650 7.8165 7.8480 8.9100 ;
      RECT 7.7650 7.9050 7.8620 8.8405 ;
      RECT 16.4440 7.8165 16.5290 8.9100 ;
      RECT 16.3000 7.8165 16.3260 8.9100 ;
      RECT 16.1920 7.8165 16.2180 8.9100 ;
      RECT 16.0840 7.8165 16.1100 8.9100 ;
      RECT 15.9760 7.8165 16.0020 8.9100 ;
      RECT 15.8680 7.8165 15.8940 8.9100 ;
      RECT 15.7600 7.8165 15.7860 8.9100 ;
      RECT 15.6520 7.8165 15.6780 8.9100 ;
      RECT 15.5440 7.8165 15.5700 8.9100 ;
      RECT 15.4360 7.8165 15.4620 8.9100 ;
      RECT 15.3280 7.8165 15.3540 8.9100 ;
      RECT 15.2200 7.8165 15.2460 8.9100 ;
      RECT 15.1120 7.8165 15.1380 8.9100 ;
      RECT 15.0040 7.8165 15.0300 8.9100 ;
      RECT 14.8960 7.8165 14.9220 8.9100 ;
      RECT 14.7880 7.8165 14.8140 8.9100 ;
      RECT 14.6800 7.8165 14.7060 8.9100 ;
      RECT 14.5720 7.8165 14.5980 8.9100 ;
      RECT 14.4640 7.8165 14.4900 8.9100 ;
      RECT 14.3560 7.8165 14.3820 8.9100 ;
      RECT 14.2480 7.8165 14.2740 8.9100 ;
      RECT 14.1400 7.8165 14.1660 8.9100 ;
      RECT 14.0320 7.8165 14.0580 8.9100 ;
      RECT 13.9240 7.8165 13.9500 8.9100 ;
      RECT 13.8160 7.8165 13.8420 8.9100 ;
      RECT 13.7080 7.8165 13.7340 8.9100 ;
      RECT 13.6000 7.8165 13.6260 8.9100 ;
      RECT 13.4920 7.8165 13.5180 8.9100 ;
      RECT 13.3840 7.8165 13.4100 8.9100 ;
      RECT 13.2760 7.8165 13.3020 8.9100 ;
      RECT 13.1680 7.8165 13.1940 8.9100 ;
      RECT 13.0600 7.8165 13.0860 8.9100 ;
      RECT 12.9520 7.8165 12.9780 8.9100 ;
      RECT 12.8440 7.8165 12.8700 8.9100 ;
      RECT 12.7360 7.8165 12.7620 8.9100 ;
      RECT 12.6280 7.8165 12.6540 8.9100 ;
      RECT 12.5200 7.8165 12.5460 8.9100 ;
      RECT 12.4120 7.8165 12.4380 8.9100 ;
      RECT 12.3040 7.8165 12.3300 8.9100 ;
      RECT 12.1960 7.8165 12.2220 8.9100 ;
      RECT 12.0880 7.8165 12.1140 8.9100 ;
      RECT 11.9800 7.8165 12.0060 8.9100 ;
      RECT 11.8720 7.8165 11.8980 8.9100 ;
      RECT 11.7640 7.8165 11.7900 8.9100 ;
      RECT 11.6560 7.8165 11.6820 8.9100 ;
      RECT 11.5480 7.8165 11.5740 8.9100 ;
      RECT 11.4400 7.8165 11.4660 8.9100 ;
      RECT 11.3320 7.8165 11.3580 8.9100 ;
      RECT 11.2240 7.8165 11.2500 8.9100 ;
      RECT 11.1160 7.8165 11.1420 8.9100 ;
      RECT 11.0080 7.8165 11.0340 8.9100 ;
      RECT 10.9000 7.8165 10.9260 8.9100 ;
      RECT 10.7920 7.8165 10.8180 8.9100 ;
      RECT 10.6840 7.8165 10.7100 8.9100 ;
      RECT 10.5760 7.8165 10.6020 8.9100 ;
      RECT 10.4680 7.8165 10.4940 8.9100 ;
      RECT 10.3600 7.8165 10.3860 8.9100 ;
      RECT 10.2520 7.8165 10.2780 8.9100 ;
      RECT 10.1440 7.8165 10.1700 8.9100 ;
      RECT 10.0360 7.8165 10.0620 8.9100 ;
      RECT 9.9280 7.8165 9.9540 8.9100 ;
      RECT 9.8200 7.8165 9.8460 8.9100 ;
      RECT 9.7120 7.8165 9.7380 8.9100 ;
      RECT 9.6040 7.8165 9.6300 8.9100 ;
      RECT 9.4960 7.8165 9.5220 8.9100 ;
      RECT 9.3880 7.8165 9.4140 8.9100 ;
      RECT 9.1750 7.8165 9.2520 8.9100 ;
      RECT 7.2820 7.8165 7.3590 8.9100 ;
      RECT 7.1200 7.8165 7.1460 8.9100 ;
      RECT 7.0120 7.8165 7.0380 8.9100 ;
      RECT 6.9040 7.8165 6.9300 8.9100 ;
      RECT 6.7960 7.8165 6.8220 8.9100 ;
      RECT 6.6880 7.8165 6.7140 8.9100 ;
      RECT 6.5800 7.8165 6.6060 8.9100 ;
      RECT 6.4720 7.8165 6.4980 8.9100 ;
      RECT 6.3640 7.8165 6.3900 8.9100 ;
      RECT 6.2560 7.8165 6.2820 8.9100 ;
      RECT 6.1480 7.8165 6.1740 8.9100 ;
      RECT 6.0400 7.8165 6.0660 8.9100 ;
      RECT 5.9320 7.8165 5.9580 8.9100 ;
      RECT 5.8240 7.8165 5.8500 8.9100 ;
      RECT 5.7160 7.8165 5.7420 8.9100 ;
      RECT 5.6080 7.8165 5.6340 8.9100 ;
      RECT 5.5000 7.8165 5.5260 8.9100 ;
      RECT 5.3920 7.8165 5.4180 8.9100 ;
      RECT 5.2840 7.8165 5.3100 8.9100 ;
      RECT 5.1760 7.8165 5.2020 8.9100 ;
      RECT 5.0680 7.8165 5.0940 8.9100 ;
      RECT 4.9600 7.8165 4.9860 8.9100 ;
      RECT 4.8520 7.8165 4.8780 8.9100 ;
      RECT 4.7440 7.8165 4.7700 8.9100 ;
      RECT 4.6360 7.8165 4.6620 8.9100 ;
      RECT 4.5280 7.8165 4.5540 8.9100 ;
      RECT 4.4200 7.8165 4.4460 8.9100 ;
      RECT 4.3120 7.8165 4.3380 8.9100 ;
      RECT 4.2040 7.8165 4.2300 8.9100 ;
      RECT 4.0960 7.8165 4.1220 8.9100 ;
      RECT 3.9880 7.8165 4.0140 8.9100 ;
      RECT 3.8800 7.8165 3.9060 8.9100 ;
      RECT 3.7720 7.8165 3.7980 8.9100 ;
      RECT 3.6640 7.8165 3.6900 8.9100 ;
      RECT 3.5560 7.8165 3.5820 8.9100 ;
      RECT 3.4480 7.8165 3.4740 8.9100 ;
      RECT 3.3400 7.8165 3.3660 8.9100 ;
      RECT 3.2320 7.8165 3.2580 8.9100 ;
      RECT 3.1240 7.8165 3.1500 8.9100 ;
      RECT 3.0160 7.8165 3.0420 8.9100 ;
      RECT 2.9080 7.8165 2.9340 8.9100 ;
      RECT 2.8000 7.8165 2.8260 8.9100 ;
      RECT 2.6920 7.8165 2.7180 8.9100 ;
      RECT 2.5840 7.8165 2.6100 8.9100 ;
      RECT 2.4760 7.8165 2.5020 8.9100 ;
      RECT 2.3680 7.8165 2.3940 8.9100 ;
      RECT 2.2600 7.8165 2.2860 8.9100 ;
      RECT 2.1520 7.8165 2.1780 8.9100 ;
      RECT 2.0440 7.8165 2.0700 8.9100 ;
      RECT 1.9360 7.8165 1.9620 8.9100 ;
      RECT 1.8280 7.8165 1.8540 8.9100 ;
      RECT 1.7200 7.8165 1.7460 8.9100 ;
      RECT 1.6120 7.8165 1.6380 8.9100 ;
      RECT 1.5040 7.8165 1.5300 8.9100 ;
      RECT 1.3960 7.8165 1.4220 8.9100 ;
      RECT 1.2880 7.8165 1.3140 8.9100 ;
      RECT 1.1800 7.8165 1.2060 8.9100 ;
      RECT 1.0720 7.8165 1.0980 8.9100 ;
      RECT 0.9640 7.8165 0.9900 8.9100 ;
      RECT 0.8560 7.8165 0.8820 8.9100 ;
      RECT 0.7480 7.8165 0.7740 8.9100 ;
      RECT 0.6400 7.8165 0.6660 8.9100 ;
      RECT 0.5320 7.8165 0.5580 8.9100 ;
      RECT 0.4240 7.8165 0.4500 8.9100 ;
      RECT 0.3160 7.8165 0.3420 8.9100 ;
      RECT 0.2080 7.8165 0.2340 8.9100 ;
      RECT 0.0050 7.8165 0.0900 8.9100 ;
      RECT 8.6410 8.8965 8.7690 9.9900 ;
      RECT 8.6270 9.5620 8.7690 9.8845 ;
      RECT 8.4790 9.2890 8.5410 9.9900 ;
      RECT 8.4650 9.5985 8.5410 9.7520 ;
      RECT 8.4790 8.8965 8.5050 9.9900 ;
      RECT 8.4790 9.0175 8.5190 9.2570 ;
      RECT 8.4790 8.8965 8.5410 8.9855 ;
      RECT 8.1820 9.3470 8.3880 9.9900 ;
      RECT 8.3620 8.8965 8.3880 9.9900 ;
      RECT 8.1820 9.6240 8.4020 9.8820 ;
      RECT 8.1820 8.8965 8.2800 9.9900 ;
      RECT 7.7650 8.8965 7.8480 9.9900 ;
      RECT 7.7650 8.9850 7.8620 9.9205 ;
      RECT 16.4440 8.8965 16.5290 9.9900 ;
      RECT 16.3000 8.8965 16.3260 9.9900 ;
      RECT 16.1920 8.8965 16.2180 9.9900 ;
      RECT 16.0840 8.8965 16.1100 9.9900 ;
      RECT 15.9760 8.8965 16.0020 9.9900 ;
      RECT 15.8680 8.8965 15.8940 9.9900 ;
      RECT 15.7600 8.8965 15.7860 9.9900 ;
      RECT 15.6520 8.8965 15.6780 9.9900 ;
      RECT 15.5440 8.8965 15.5700 9.9900 ;
      RECT 15.4360 8.8965 15.4620 9.9900 ;
      RECT 15.3280 8.8965 15.3540 9.9900 ;
      RECT 15.2200 8.8965 15.2460 9.9900 ;
      RECT 15.1120 8.8965 15.1380 9.9900 ;
      RECT 15.0040 8.8965 15.0300 9.9900 ;
      RECT 14.8960 8.8965 14.9220 9.9900 ;
      RECT 14.7880 8.8965 14.8140 9.9900 ;
      RECT 14.6800 8.8965 14.7060 9.9900 ;
      RECT 14.5720 8.8965 14.5980 9.9900 ;
      RECT 14.4640 8.8965 14.4900 9.9900 ;
      RECT 14.3560 8.8965 14.3820 9.9900 ;
      RECT 14.2480 8.8965 14.2740 9.9900 ;
      RECT 14.1400 8.8965 14.1660 9.9900 ;
      RECT 14.0320 8.8965 14.0580 9.9900 ;
      RECT 13.9240 8.8965 13.9500 9.9900 ;
      RECT 13.8160 8.8965 13.8420 9.9900 ;
      RECT 13.7080 8.8965 13.7340 9.9900 ;
      RECT 13.6000 8.8965 13.6260 9.9900 ;
      RECT 13.4920 8.8965 13.5180 9.9900 ;
      RECT 13.3840 8.8965 13.4100 9.9900 ;
      RECT 13.2760 8.8965 13.3020 9.9900 ;
      RECT 13.1680 8.8965 13.1940 9.9900 ;
      RECT 13.0600 8.8965 13.0860 9.9900 ;
      RECT 12.9520 8.8965 12.9780 9.9900 ;
      RECT 12.8440 8.8965 12.8700 9.9900 ;
      RECT 12.7360 8.8965 12.7620 9.9900 ;
      RECT 12.6280 8.8965 12.6540 9.9900 ;
      RECT 12.5200 8.8965 12.5460 9.9900 ;
      RECT 12.4120 8.8965 12.4380 9.9900 ;
      RECT 12.3040 8.8965 12.3300 9.9900 ;
      RECT 12.1960 8.8965 12.2220 9.9900 ;
      RECT 12.0880 8.8965 12.1140 9.9900 ;
      RECT 11.9800 8.8965 12.0060 9.9900 ;
      RECT 11.8720 8.8965 11.8980 9.9900 ;
      RECT 11.7640 8.8965 11.7900 9.9900 ;
      RECT 11.6560 8.8965 11.6820 9.9900 ;
      RECT 11.5480 8.8965 11.5740 9.9900 ;
      RECT 11.4400 8.8965 11.4660 9.9900 ;
      RECT 11.3320 8.8965 11.3580 9.9900 ;
      RECT 11.2240 8.8965 11.2500 9.9900 ;
      RECT 11.1160 8.8965 11.1420 9.9900 ;
      RECT 11.0080 8.8965 11.0340 9.9900 ;
      RECT 10.9000 8.8965 10.9260 9.9900 ;
      RECT 10.7920 8.8965 10.8180 9.9900 ;
      RECT 10.6840 8.8965 10.7100 9.9900 ;
      RECT 10.5760 8.8965 10.6020 9.9900 ;
      RECT 10.4680 8.8965 10.4940 9.9900 ;
      RECT 10.3600 8.8965 10.3860 9.9900 ;
      RECT 10.2520 8.8965 10.2780 9.9900 ;
      RECT 10.1440 8.8965 10.1700 9.9900 ;
      RECT 10.0360 8.8965 10.0620 9.9900 ;
      RECT 9.9280 8.8965 9.9540 9.9900 ;
      RECT 9.8200 8.8965 9.8460 9.9900 ;
      RECT 9.7120 8.8965 9.7380 9.9900 ;
      RECT 9.6040 8.8965 9.6300 9.9900 ;
      RECT 9.4960 8.8965 9.5220 9.9900 ;
      RECT 9.3880 8.8965 9.4140 9.9900 ;
      RECT 9.1750 8.8965 9.2520 9.9900 ;
      RECT 7.2820 8.8965 7.3590 9.9900 ;
      RECT 7.1200 8.8965 7.1460 9.9900 ;
      RECT 7.0120 8.8965 7.0380 9.9900 ;
      RECT 6.9040 8.8965 6.9300 9.9900 ;
      RECT 6.7960 8.8965 6.8220 9.9900 ;
      RECT 6.6880 8.8965 6.7140 9.9900 ;
      RECT 6.5800 8.8965 6.6060 9.9900 ;
      RECT 6.4720 8.8965 6.4980 9.9900 ;
      RECT 6.3640 8.8965 6.3900 9.9900 ;
      RECT 6.2560 8.8965 6.2820 9.9900 ;
      RECT 6.1480 8.8965 6.1740 9.9900 ;
      RECT 6.0400 8.8965 6.0660 9.9900 ;
      RECT 5.9320 8.8965 5.9580 9.9900 ;
      RECT 5.8240 8.8965 5.8500 9.9900 ;
      RECT 5.7160 8.8965 5.7420 9.9900 ;
      RECT 5.6080 8.8965 5.6340 9.9900 ;
      RECT 5.5000 8.8965 5.5260 9.9900 ;
      RECT 5.3920 8.8965 5.4180 9.9900 ;
      RECT 5.2840 8.8965 5.3100 9.9900 ;
      RECT 5.1760 8.8965 5.2020 9.9900 ;
      RECT 5.0680 8.8965 5.0940 9.9900 ;
      RECT 4.9600 8.8965 4.9860 9.9900 ;
      RECT 4.8520 8.8965 4.8780 9.9900 ;
      RECT 4.7440 8.8965 4.7700 9.9900 ;
      RECT 4.6360 8.8965 4.6620 9.9900 ;
      RECT 4.5280 8.8965 4.5540 9.9900 ;
      RECT 4.4200 8.8965 4.4460 9.9900 ;
      RECT 4.3120 8.8965 4.3380 9.9900 ;
      RECT 4.2040 8.8965 4.2300 9.9900 ;
      RECT 4.0960 8.8965 4.1220 9.9900 ;
      RECT 3.9880 8.8965 4.0140 9.9900 ;
      RECT 3.8800 8.8965 3.9060 9.9900 ;
      RECT 3.7720 8.8965 3.7980 9.9900 ;
      RECT 3.6640 8.8965 3.6900 9.9900 ;
      RECT 3.5560 8.8965 3.5820 9.9900 ;
      RECT 3.4480 8.8965 3.4740 9.9900 ;
      RECT 3.3400 8.8965 3.3660 9.9900 ;
      RECT 3.2320 8.8965 3.2580 9.9900 ;
      RECT 3.1240 8.8965 3.1500 9.9900 ;
      RECT 3.0160 8.8965 3.0420 9.9900 ;
      RECT 2.9080 8.8965 2.9340 9.9900 ;
      RECT 2.8000 8.8965 2.8260 9.9900 ;
      RECT 2.6920 8.8965 2.7180 9.9900 ;
      RECT 2.5840 8.8965 2.6100 9.9900 ;
      RECT 2.4760 8.8965 2.5020 9.9900 ;
      RECT 2.3680 8.8965 2.3940 9.9900 ;
      RECT 2.2600 8.8965 2.2860 9.9900 ;
      RECT 2.1520 8.8965 2.1780 9.9900 ;
      RECT 2.0440 8.8965 2.0700 9.9900 ;
      RECT 1.9360 8.8965 1.9620 9.9900 ;
      RECT 1.8280 8.8965 1.8540 9.9900 ;
      RECT 1.7200 8.8965 1.7460 9.9900 ;
      RECT 1.6120 8.8965 1.6380 9.9900 ;
      RECT 1.5040 8.8965 1.5300 9.9900 ;
      RECT 1.3960 8.8965 1.4220 9.9900 ;
      RECT 1.2880 8.8965 1.3140 9.9900 ;
      RECT 1.1800 8.8965 1.2060 9.9900 ;
      RECT 1.0720 8.8965 1.0980 9.9900 ;
      RECT 0.9640 8.8965 0.9900 9.9900 ;
      RECT 0.8560 8.8965 0.8820 9.9900 ;
      RECT 0.7480 8.8965 0.7740 9.9900 ;
      RECT 0.6400 8.8965 0.6660 9.9900 ;
      RECT 0.5320 8.8965 0.5580 9.9900 ;
      RECT 0.4240 8.8965 0.4500 9.9900 ;
      RECT 0.3160 8.8965 0.3420 9.9900 ;
      RECT 0.2080 8.8965 0.2340 9.9900 ;
      RECT 0.0050 8.8965 0.0900 9.9900 ;
      RECT 8.6410 9.9765 8.7690 11.0700 ;
      RECT 8.6270 10.6420 8.7690 10.9645 ;
      RECT 8.4790 10.3690 8.5410 11.0700 ;
      RECT 8.4650 10.6785 8.5410 10.8320 ;
      RECT 8.4790 9.9765 8.5050 11.0700 ;
      RECT 8.4790 10.0975 8.5190 10.3370 ;
      RECT 8.4790 9.9765 8.5410 10.0655 ;
      RECT 8.1820 10.4270 8.3880 11.0700 ;
      RECT 8.3620 9.9765 8.3880 11.0700 ;
      RECT 8.1820 10.7040 8.4020 10.9620 ;
      RECT 8.1820 9.9765 8.2800 11.0700 ;
      RECT 7.7650 9.9765 7.8480 11.0700 ;
      RECT 7.7650 10.0650 7.8620 11.0005 ;
      RECT 16.4440 9.9765 16.5290 11.0700 ;
      RECT 16.3000 9.9765 16.3260 11.0700 ;
      RECT 16.1920 9.9765 16.2180 11.0700 ;
      RECT 16.0840 9.9765 16.1100 11.0700 ;
      RECT 15.9760 9.9765 16.0020 11.0700 ;
      RECT 15.8680 9.9765 15.8940 11.0700 ;
      RECT 15.7600 9.9765 15.7860 11.0700 ;
      RECT 15.6520 9.9765 15.6780 11.0700 ;
      RECT 15.5440 9.9765 15.5700 11.0700 ;
      RECT 15.4360 9.9765 15.4620 11.0700 ;
      RECT 15.3280 9.9765 15.3540 11.0700 ;
      RECT 15.2200 9.9765 15.2460 11.0700 ;
      RECT 15.1120 9.9765 15.1380 11.0700 ;
      RECT 15.0040 9.9765 15.0300 11.0700 ;
      RECT 14.8960 9.9765 14.9220 11.0700 ;
      RECT 14.7880 9.9765 14.8140 11.0700 ;
      RECT 14.6800 9.9765 14.7060 11.0700 ;
      RECT 14.5720 9.9765 14.5980 11.0700 ;
      RECT 14.4640 9.9765 14.4900 11.0700 ;
      RECT 14.3560 9.9765 14.3820 11.0700 ;
      RECT 14.2480 9.9765 14.2740 11.0700 ;
      RECT 14.1400 9.9765 14.1660 11.0700 ;
      RECT 14.0320 9.9765 14.0580 11.0700 ;
      RECT 13.9240 9.9765 13.9500 11.0700 ;
      RECT 13.8160 9.9765 13.8420 11.0700 ;
      RECT 13.7080 9.9765 13.7340 11.0700 ;
      RECT 13.6000 9.9765 13.6260 11.0700 ;
      RECT 13.4920 9.9765 13.5180 11.0700 ;
      RECT 13.3840 9.9765 13.4100 11.0700 ;
      RECT 13.2760 9.9765 13.3020 11.0700 ;
      RECT 13.1680 9.9765 13.1940 11.0700 ;
      RECT 13.0600 9.9765 13.0860 11.0700 ;
      RECT 12.9520 9.9765 12.9780 11.0700 ;
      RECT 12.8440 9.9765 12.8700 11.0700 ;
      RECT 12.7360 9.9765 12.7620 11.0700 ;
      RECT 12.6280 9.9765 12.6540 11.0700 ;
      RECT 12.5200 9.9765 12.5460 11.0700 ;
      RECT 12.4120 9.9765 12.4380 11.0700 ;
      RECT 12.3040 9.9765 12.3300 11.0700 ;
      RECT 12.1960 9.9765 12.2220 11.0700 ;
      RECT 12.0880 9.9765 12.1140 11.0700 ;
      RECT 11.9800 9.9765 12.0060 11.0700 ;
      RECT 11.8720 9.9765 11.8980 11.0700 ;
      RECT 11.7640 9.9765 11.7900 11.0700 ;
      RECT 11.6560 9.9765 11.6820 11.0700 ;
      RECT 11.5480 9.9765 11.5740 11.0700 ;
      RECT 11.4400 9.9765 11.4660 11.0700 ;
      RECT 11.3320 9.9765 11.3580 11.0700 ;
      RECT 11.2240 9.9765 11.2500 11.0700 ;
      RECT 11.1160 9.9765 11.1420 11.0700 ;
      RECT 11.0080 9.9765 11.0340 11.0700 ;
      RECT 10.9000 9.9765 10.9260 11.0700 ;
      RECT 10.7920 9.9765 10.8180 11.0700 ;
      RECT 10.6840 9.9765 10.7100 11.0700 ;
      RECT 10.5760 9.9765 10.6020 11.0700 ;
      RECT 10.4680 9.9765 10.4940 11.0700 ;
      RECT 10.3600 9.9765 10.3860 11.0700 ;
      RECT 10.2520 9.9765 10.2780 11.0700 ;
      RECT 10.1440 9.9765 10.1700 11.0700 ;
      RECT 10.0360 9.9765 10.0620 11.0700 ;
      RECT 9.9280 9.9765 9.9540 11.0700 ;
      RECT 9.8200 9.9765 9.8460 11.0700 ;
      RECT 9.7120 9.9765 9.7380 11.0700 ;
      RECT 9.6040 9.9765 9.6300 11.0700 ;
      RECT 9.4960 9.9765 9.5220 11.0700 ;
      RECT 9.3880 9.9765 9.4140 11.0700 ;
      RECT 9.1750 9.9765 9.2520 11.0700 ;
      RECT 7.2820 9.9765 7.3590 11.0700 ;
      RECT 7.1200 9.9765 7.1460 11.0700 ;
      RECT 7.0120 9.9765 7.0380 11.0700 ;
      RECT 6.9040 9.9765 6.9300 11.0700 ;
      RECT 6.7960 9.9765 6.8220 11.0700 ;
      RECT 6.6880 9.9765 6.7140 11.0700 ;
      RECT 6.5800 9.9765 6.6060 11.0700 ;
      RECT 6.4720 9.9765 6.4980 11.0700 ;
      RECT 6.3640 9.9765 6.3900 11.0700 ;
      RECT 6.2560 9.9765 6.2820 11.0700 ;
      RECT 6.1480 9.9765 6.1740 11.0700 ;
      RECT 6.0400 9.9765 6.0660 11.0700 ;
      RECT 5.9320 9.9765 5.9580 11.0700 ;
      RECT 5.8240 9.9765 5.8500 11.0700 ;
      RECT 5.7160 9.9765 5.7420 11.0700 ;
      RECT 5.6080 9.9765 5.6340 11.0700 ;
      RECT 5.5000 9.9765 5.5260 11.0700 ;
      RECT 5.3920 9.9765 5.4180 11.0700 ;
      RECT 5.2840 9.9765 5.3100 11.0700 ;
      RECT 5.1760 9.9765 5.2020 11.0700 ;
      RECT 5.0680 9.9765 5.0940 11.0700 ;
      RECT 4.9600 9.9765 4.9860 11.0700 ;
      RECT 4.8520 9.9765 4.8780 11.0700 ;
      RECT 4.7440 9.9765 4.7700 11.0700 ;
      RECT 4.6360 9.9765 4.6620 11.0700 ;
      RECT 4.5280 9.9765 4.5540 11.0700 ;
      RECT 4.4200 9.9765 4.4460 11.0700 ;
      RECT 4.3120 9.9765 4.3380 11.0700 ;
      RECT 4.2040 9.9765 4.2300 11.0700 ;
      RECT 4.0960 9.9765 4.1220 11.0700 ;
      RECT 3.9880 9.9765 4.0140 11.0700 ;
      RECT 3.8800 9.9765 3.9060 11.0700 ;
      RECT 3.7720 9.9765 3.7980 11.0700 ;
      RECT 3.6640 9.9765 3.6900 11.0700 ;
      RECT 3.5560 9.9765 3.5820 11.0700 ;
      RECT 3.4480 9.9765 3.4740 11.0700 ;
      RECT 3.3400 9.9765 3.3660 11.0700 ;
      RECT 3.2320 9.9765 3.2580 11.0700 ;
      RECT 3.1240 9.9765 3.1500 11.0700 ;
      RECT 3.0160 9.9765 3.0420 11.0700 ;
      RECT 2.9080 9.9765 2.9340 11.0700 ;
      RECT 2.8000 9.9765 2.8260 11.0700 ;
      RECT 2.6920 9.9765 2.7180 11.0700 ;
      RECT 2.5840 9.9765 2.6100 11.0700 ;
      RECT 2.4760 9.9765 2.5020 11.0700 ;
      RECT 2.3680 9.9765 2.3940 11.0700 ;
      RECT 2.2600 9.9765 2.2860 11.0700 ;
      RECT 2.1520 9.9765 2.1780 11.0700 ;
      RECT 2.0440 9.9765 2.0700 11.0700 ;
      RECT 1.9360 9.9765 1.9620 11.0700 ;
      RECT 1.8280 9.9765 1.8540 11.0700 ;
      RECT 1.7200 9.9765 1.7460 11.0700 ;
      RECT 1.6120 9.9765 1.6380 11.0700 ;
      RECT 1.5040 9.9765 1.5300 11.0700 ;
      RECT 1.3960 9.9765 1.4220 11.0700 ;
      RECT 1.2880 9.9765 1.3140 11.0700 ;
      RECT 1.1800 9.9765 1.2060 11.0700 ;
      RECT 1.0720 9.9765 1.0980 11.0700 ;
      RECT 0.9640 9.9765 0.9900 11.0700 ;
      RECT 0.8560 9.9765 0.8820 11.0700 ;
      RECT 0.7480 9.9765 0.7740 11.0700 ;
      RECT 0.6400 9.9765 0.6660 11.0700 ;
      RECT 0.5320 9.9765 0.5580 11.0700 ;
      RECT 0.4240 9.9765 0.4500 11.0700 ;
      RECT 0.3160 9.9765 0.3420 11.0700 ;
      RECT 0.2080 9.9765 0.2340 11.0700 ;
      RECT 0.0050 9.9765 0.0900 11.0700 ;
      RECT 8.6410 11.0565 8.7690 12.1500 ;
      RECT 8.6270 11.7220 8.7690 12.0445 ;
      RECT 8.4790 11.4490 8.5410 12.1500 ;
      RECT 8.4650 11.7585 8.5410 11.9120 ;
      RECT 8.4790 11.0565 8.5050 12.1500 ;
      RECT 8.4790 11.1775 8.5190 11.4170 ;
      RECT 8.4790 11.0565 8.5410 11.1455 ;
      RECT 8.1820 11.5070 8.3880 12.1500 ;
      RECT 8.3620 11.0565 8.3880 12.1500 ;
      RECT 8.1820 11.7840 8.4020 12.0420 ;
      RECT 8.1820 11.0565 8.2800 12.1500 ;
      RECT 7.7650 11.0565 7.8480 12.1500 ;
      RECT 7.7650 11.1450 7.8620 12.0805 ;
      RECT 16.4440 11.0565 16.5290 12.1500 ;
      RECT 16.3000 11.0565 16.3260 12.1500 ;
      RECT 16.1920 11.0565 16.2180 12.1500 ;
      RECT 16.0840 11.0565 16.1100 12.1500 ;
      RECT 15.9760 11.0565 16.0020 12.1500 ;
      RECT 15.8680 11.0565 15.8940 12.1500 ;
      RECT 15.7600 11.0565 15.7860 12.1500 ;
      RECT 15.6520 11.0565 15.6780 12.1500 ;
      RECT 15.5440 11.0565 15.5700 12.1500 ;
      RECT 15.4360 11.0565 15.4620 12.1500 ;
      RECT 15.3280 11.0565 15.3540 12.1500 ;
      RECT 15.2200 11.0565 15.2460 12.1500 ;
      RECT 15.1120 11.0565 15.1380 12.1500 ;
      RECT 15.0040 11.0565 15.0300 12.1500 ;
      RECT 14.8960 11.0565 14.9220 12.1500 ;
      RECT 14.7880 11.0565 14.8140 12.1500 ;
      RECT 14.6800 11.0565 14.7060 12.1500 ;
      RECT 14.5720 11.0565 14.5980 12.1500 ;
      RECT 14.4640 11.0565 14.4900 12.1500 ;
      RECT 14.3560 11.0565 14.3820 12.1500 ;
      RECT 14.2480 11.0565 14.2740 12.1500 ;
      RECT 14.1400 11.0565 14.1660 12.1500 ;
      RECT 14.0320 11.0565 14.0580 12.1500 ;
      RECT 13.9240 11.0565 13.9500 12.1500 ;
      RECT 13.8160 11.0565 13.8420 12.1500 ;
      RECT 13.7080 11.0565 13.7340 12.1500 ;
      RECT 13.6000 11.0565 13.6260 12.1500 ;
      RECT 13.4920 11.0565 13.5180 12.1500 ;
      RECT 13.3840 11.0565 13.4100 12.1500 ;
      RECT 13.2760 11.0565 13.3020 12.1500 ;
      RECT 13.1680 11.0565 13.1940 12.1500 ;
      RECT 13.0600 11.0565 13.0860 12.1500 ;
      RECT 12.9520 11.0565 12.9780 12.1500 ;
      RECT 12.8440 11.0565 12.8700 12.1500 ;
      RECT 12.7360 11.0565 12.7620 12.1500 ;
      RECT 12.6280 11.0565 12.6540 12.1500 ;
      RECT 12.5200 11.0565 12.5460 12.1500 ;
      RECT 12.4120 11.0565 12.4380 12.1500 ;
      RECT 12.3040 11.0565 12.3300 12.1500 ;
      RECT 12.1960 11.0565 12.2220 12.1500 ;
      RECT 12.0880 11.0565 12.1140 12.1500 ;
      RECT 11.9800 11.0565 12.0060 12.1500 ;
      RECT 11.8720 11.0565 11.8980 12.1500 ;
      RECT 11.7640 11.0565 11.7900 12.1500 ;
      RECT 11.6560 11.0565 11.6820 12.1500 ;
      RECT 11.5480 11.0565 11.5740 12.1500 ;
      RECT 11.4400 11.0565 11.4660 12.1500 ;
      RECT 11.3320 11.0565 11.3580 12.1500 ;
      RECT 11.2240 11.0565 11.2500 12.1500 ;
      RECT 11.1160 11.0565 11.1420 12.1500 ;
      RECT 11.0080 11.0565 11.0340 12.1500 ;
      RECT 10.9000 11.0565 10.9260 12.1500 ;
      RECT 10.7920 11.0565 10.8180 12.1500 ;
      RECT 10.6840 11.0565 10.7100 12.1500 ;
      RECT 10.5760 11.0565 10.6020 12.1500 ;
      RECT 10.4680 11.0565 10.4940 12.1500 ;
      RECT 10.3600 11.0565 10.3860 12.1500 ;
      RECT 10.2520 11.0565 10.2780 12.1500 ;
      RECT 10.1440 11.0565 10.1700 12.1500 ;
      RECT 10.0360 11.0565 10.0620 12.1500 ;
      RECT 9.9280 11.0565 9.9540 12.1500 ;
      RECT 9.8200 11.0565 9.8460 12.1500 ;
      RECT 9.7120 11.0565 9.7380 12.1500 ;
      RECT 9.6040 11.0565 9.6300 12.1500 ;
      RECT 9.4960 11.0565 9.5220 12.1500 ;
      RECT 9.3880 11.0565 9.4140 12.1500 ;
      RECT 9.1750 11.0565 9.2520 12.1500 ;
      RECT 7.2820 11.0565 7.3590 12.1500 ;
      RECT 7.1200 11.0565 7.1460 12.1500 ;
      RECT 7.0120 11.0565 7.0380 12.1500 ;
      RECT 6.9040 11.0565 6.9300 12.1500 ;
      RECT 6.7960 11.0565 6.8220 12.1500 ;
      RECT 6.6880 11.0565 6.7140 12.1500 ;
      RECT 6.5800 11.0565 6.6060 12.1500 ;
      RECT 6.4720 11.0565 6.4980 12.1500 ;
      RECT 6.3640 11.0565 6.3900 12.1500 ;
      RECT 6.2560 11.0565 6.2820 12.1500 ;
      RECT 6.1480 11.0565 6.1740 12.1500 ;
      RECT 6.0400 11.0565 6.0660 12.1500 ;
      RECT 5.9320 11.0565 5.9580 12.1500 ;
      RECT 5.8240 11.0565 5.8500 12.1500 ;
      RECT 5.7160 11.0565 5.7420 12.1500 ;
      RECT 5.6080 11.0565 5.6340 12.1500 ;
      RECT 5.5000 11.0565 5.5260 12.1500 ;
      RECT 5.3920 11.0565 5.4180 12.1500 ;
      RECT 5.2840 11.0565 5.3100 12.1500 ;
      RECT 5.1760 11.0565 5.2020 12.1500 ;
      RECT 5.0680 11.0565 5.0940 12.1500 ;
      RECT 4.9600 11.0565 4.9860 12.1500 ;
      RECT 4.8520 11.0565 4.8780 12.1500 ;
      RECT 4.7440 11.0565 4.7700 12.1500 ;
      RECT 4.6360 11.0565 4.6620 12.1500 ;
      RECT 4.5280 11.0565 4.5540 12.1500 ;
      RECT 4.4200 11.0565 4.4460 12.1500 ;
      RECT 4.3120 11.0565 4.3380 12.1500 ;
      RECT 4.2040 11.0565 4.2300 12.1500 ;
      RECT 4.0960 11.0565 4.1220 12.1500 ;
      RECT 3.9880 11.0565 4.0140 12.1500 ;
      RECT 3.8800 11.0565 3.9060 12.1500 ;
      RECT 3.7720 11.0565 3.7980 12.1500 ;
      RECT 3.6640 11.0565 3.6900 12.1500 ;
      RECT 3.5560 11.0565 3.5820 12.1500 ;
      RECT 3.4480 11.0565 3.4740 12.1500 ;
      RECT 3.3400 11.0565 3.3660 12.1500 ;
      RECT 3.2320 11.0565 3.2580 12.1500 ;
      RECT 3.1240 11.0565 3.1500 12.1500 ;
      RECT 3.0160 11.0565 3.0420 12.1500 ;
      RECT 2.9080 11.0565 2.9340 12.1500 ;
      RECT 2.8000 11.0565 2.8260 12.1500 ;
      RECT 2.6920 11.0565 2.7180 12.1500 ;
      RECT 2.5840 11.0565 2.6100 12.1500 ;
      RECT 2.4760 11.0565 2.5020 12.1500 ;
      RECT 2.3680 11.0565 2.3940 12.1500 ;
      RECT 2.2600 11.0565 2.2860 12.1500 ;
      RECT 2.1520 11.0565 2.1780 12.1500 ;
      RECT 2.0440 11.0565 2.0700 12.1500 ;
      RECT 1.9360 11.0565 1.9620 12.1500 ;
      RECT 1.8280 11.0565 1.8540 12.1500 ;
      RECT 1.7200 11.0565 1.7460 12.1500 ;
      RECT 1.6120 11.0565 1.6380 12.1500 ;
      RECT 1.5040 11.0565 1.5300 12.1500 ;
      RECT 1.3960 11.0565 1.4220 12.1500 ;
      RECT 1.2880 11.0565 1.3140 12.1500 ;
      RECT 1.1800 11.0565 1.2060 12.1500 ;
      RECT 1.0720 11.0565 1.0980 12.1500 ;
      RECT 0.9640 11.0565 0.9900 12.1500 ;
      RECT 0.8560 11.0565 0.8820 12.1500 ;
      RECT 0.7480 11.0565 0.7740 12.1500 ;
      RECT 0.6400 11.0565 0.6660 12.1500 ;
      RECT 0.5320 11.0565 0.5580 12.1500 ;
      RECT 0.4240 11.0565 0.4500 12.1500 ;
      RECT 0.3160 11.0565 0.3420 12.1500 ;
      RECT 0.2080 11.0565 0.2340 12.1500 ;
      RECT 0.0050 11.0565 0.0900 12.1500 ;
      RECT 8.6410 12.1365 8.7690 13.2300 ;
      RECT 8.6270 12.8020 8.7690 13.1245 ;
      RECT 8.4790 12.5290 8.5410 13.2300 ;
      RECT 8.4650 12.8385 8.5410 12.9920 ;
      RECT 8.4790 12.1365 8.5050 13.2300 ;
      RECT 8.4790 12.2575 8.5190 12.4970 ;
      RECT 8.4790 12.1365 8.5410 12.2255 ;
      RECT 8.1820 12.5870 8.3880 13.2300 ;
      RECT 8.3620 12.1365 8.3880 13.2300 ;
      RECT 8.1820 12.8640 8.4020 13.1220 ;
      RECT 8.1820 12.1365 8.2800 13.2300 ;
      RECT 7.7650 12.1365 7.8480 13.2300 ;
      RECT 7.7650 12.2250 7.8620 13.1605 ;
      RECT 16.4440 12.1365 16.5290 13.2300 ;
      RECT 16.3000 12.1365 16.3260 13.2300 ;
      RECT 16.1920 12.1365 16.2180 13.2300 ;
      RECT 16.0840 12.1365 16.1100 13.2300 ;
      RECT 15.9760 12.1365 16.0020 13.2300 ;
      RECT 15.8680 12.1365 15.8940 13.2300 ;
      RECT 15.7600 12.1365 15.7860 13.2300 ;
      RECT 15.6520 12.1365 15.6780 13.2300 ;
      RECT 15.5440 12.1365 15.5700 13.2300 ;
      RECT 15.4360 12.1365 15.4620 13.2300 ;
      RECT 15.3280 12.1365 15.3540 13.2300 ;
      RECT 15.2200 12.1365 15.2460 13.2300 ;
      RECT 15.1120 12.1365 15.1380 13.2300 ;
      RECT 15.0040 12.1365 15.0300 13.2300 ;
      RECT 14.8960 12.1365 14.9220 13.2300 ;
      RECT 14.7880 12.1365 14.8140 13.2300 ;
      RECT 14.6800 12.1365 14.7060 13.2300 ;
      RECT 14.5720 12.1365 14.5980 13.2300 ;
      RECT 14.4640 12.1365 14.4900 13.2300 ;
      RECT 14.3560 12.1365 14.3820 13.2300 ;
      RECT 14.2480 12.1365 14.2740 13.2300 ;
      RECT 14.1400 12.1365 14.1660 13.2300 ;
      RECT 14.0320 12.1365 14.0580 13.2300 ;
      RECT 13.9240 12.1365 13.9500 13.2300 ;
      RECT 13.8160 12.1365 13.8420 13.2300 ;
      RECT 13.7080 12.1365 13.7340 13.2300 ;
      RECT 13.6000 12.1365 13.6260 13.2300 ;
      RECT 13.4920 12.1365 13.5180 13.2300 ;
      RECT 13.3840 12.1365 13.4100 13.2300 ;
      RECT 13.2760 12.1365 13.3020 13.2300 ;
      RECT 13.1680 12.1365 13.1940 13.2300 ;
      RECT 13.0600 12.1365 13.0860 13.2300 ;
      RECT 12.9520 12.1365 12.9780 13.2300 ;
      RECT 12.8440 12.1365 12.8700 13.2300 ;
      RECT 12.7360 12.1365 12.7620 13.2300 ;
      RECT 12.6280 12.1365 12.6540 13.2300 ;
      RECT 12.5200 12.1365 12.5460 13.2300 ;
      RECT 12.4120 12.1365 12.4380 13.2300 ;
      RECT 12.3040 12.1365 12.3300 13.2300 ;
      RECT 12.1960 12.1365 12.2220 13.2300 ;
      RECT 12.0880 12.1365 12.1140 13.2300 ;
      RECT 11.9800 12.1365 12.0060 13.2300 ;
      RECT 11.8720 12.1365 11.8980 13.2300 ;
      RECT 11.7640 12.1365 11.7900 13.2300 ;
      RECT 11.6560 12.1365 11.6820 13.2300 ;
      RECT 11.5480 12.1365 11.5740 13.2300 ;
      RECT 11.4400 12.1365 11.4660 13.2300 ;
      RECT 11.3320 12.1365 11.3580 13.2300 ;
      RECT 11.2240 12.1365 11.2500 13.2300 ;
      RECT 11.1160 12.1365 11.1420 13.2300 ;
      RECT 11.0080 12.1365 11.0340 13.2300 ;
      RECT 10.9000 12.1365 10.9260 13.2300 ;
      RECT 10.7920 12.1365 10.8180 13.2300 ;
      RECT 10.6840 12.1365 10.7100 13.2300 ;
      RECT 10.5760 12.1365 10.6020 13.2300 ;
      RECT 10.4680 12.1365 10.4940 13.2300 ;
      RECT 10.3600 12.1365 10.3860 13.2300 ;
      RECT 10.2520 12.1365 10.2780 13.2300 ;
      RECT 10.1440 12.1365 10.1700 13.2300 ;
      RECT 10.0360 12.1365 10.0620 13.2300 ;
      RECT 9.9280 12.1365 9.9540 13.2300 ;
      RECT 9.8200 12.1365 9.8460 13.2300 ;
      RECT 9.7120 12.1365 9.7380 13.2300 ;
      RECT 9.6040 12.1365 9.6300 13.2300 ;
      RECT 9.4960 12.1365 9.5220 13.2300 ;
      RECT 9.3880 12.1365 9.4140 13.2300 ;
      RECT 9.1750 12.1365 9.2520 13.2300 ;
      RECT 7.2820 12.1365 7.3590 13.2300 ;
      RECT 7.1200 12.1365 7.1460 13.2300 ;
      RECT 7.0120 12.1365 7.0380 13.2300 ;
      RECT 6.9040 12.1365 6.9300 13.2300 ;
      RECT 6.7960 12.1365 6.8220 13.2300 ;
      RECT 6.6880 12.1365 6.7140 13.2300 ;
      RECT 6.5800 12.1365 6.6060 13.2300 ;
      RECT 6.4720 12.1365 6.4980 13.2300 ;
      RECT 6.3640 12.1365 6.3900 13.2300 ;
      RECT 6.2560 12.1365 6.2820 13.2300 ;
      RECT 6.1480 12.1365 6.1740 13.2300 ;
      RECT 6.0400 12.1365 6.0660 13.2300 ;
      RECT 5.9320 12.1365 5.9580 13.2300 ;
      RECT 5.8240 12.1365 5.8500 13.2300 ;
      RECT 5.7160 12.1365 5.7420 13.2300 ;
      RECT 5.6080 12.1365 5.6340 13.2300 ;
      RECT 5.5000 12.1365 5.5260 13.2300 ;
      RECT 5.3920 12.1365 5.4180 13.2300 ;
      RECT 5.2840 12.1365 5.3100 13.2300 ;
      RECT 5.1760 12.1365 5.2020 13.2300 ;
      RECT 5.0680 12.1365 5.0940 13.2300 ;
      RECT 4.9600 12.1365 4.9860 13.2300 ;
      RECT 4.8520 12.1365 4.8780 13.2300 ;
      RECT 4.7440 12.1365 4.7700 13.2300 ;
      RECT 4.6360 12.1365 4.6620 13.2300 ;
      RECT 4.5280 12.1365 4.5540 13.2300 ;
      RECT 4.4200 12.1365 4.4460 13.2300 ;
      RECT 4.3120 12.1365 4.3380 13.2300 ;
      RECT 4.2040 12.1365 4.2300 13.2300 ;
      RECT 4.0960 12.1365 4.1220 13.2300 ;
      RECT 3.9880 12.1365 4.0140 13.2300 ;
      RECT 3.8800 12.1365 3.9060 13.2300 ;
      RECT 3.7720 12.1365 3.7980 13.2300 ;
      RECT 3.6640 12.1365 3.6900 13.2300 ;
      RECT 3.5560 12.1365 3.5820 13.2300 ;
      RECT 3.4480 12.1365 3.4740 13.2300 ;
      RECT 3.3400 12.1365 3.3660 13.2300 ;
      RECT 3.2320 12.1365 3.2580 13.2300 ;
      RECT 3.1240 12.1365 3.1500 13.2300 ;
      RECT 3.0160 12.1365 3.0420 13.2300 ;
      RECT 2.9080 12.1365 2.9340 13.2300 ;
      RECT 2.8000 12.1365 2.8260 13.2300 ;
      RECT 2.6920 12.1365 2.7180 13.2300 ;
      RECT 2.5840 12.1365 2.6100 13.2300 ;
      RECT 2.4760 12.1365 2.5020 13.2300 ;
      RECT 2.3680 12.1365 2.3940 13.2300 ;
      RECT 2.2600 12.1365 2.2860 13.2300 ;
      RECT 2.1520 12.1365 2.1780 13.2300 ;
      RECT 2.0440 12.1365 2.0700 13.2300 ;
      RECT 1.9360 12.1365 1.9620 13.2300 ;
      RECT 1.8280 12.1365 1.8540 13.2300 ;
      RECT 1.7200 12.1365 1.7460 13.2300 ;
      RECT 1.6120 12.1365 1.6380 13.2300 ;
      RECT 1.5040 12.1365 1.5300 13.2300 ;
      RECT 1.3960 12.1365 1.4220 13.2300 ;
      RECT 1.2880 12.1365 1.3140 13.2300 ;
      RECT 1.1800 12.1365 1.2060 13.2300 ;
      RECT 1.0720 12.1365 1.0980 13.2300 ;
      RECT 0.9640 12.1365 0.9900 13.2300 ;
      RECT 0.8560 12.1365 0.8820 13.2300 ;
      RECT 0.7480 12.1365 0.7740 13.2300 ;
      RECT 0.6400 12.1365 0.6660 13.2300 ;
      RECT 0.5320 12.1365 0.5580 13.2300 ;
      RECT 0.4240 12.1365 0.4500 13.2300 ;
      RECT 0.3160 12.1365 0.3420 13.2300 ;
      RECT 0.2080 12.1365 0.2340 13.2300 ;
      RECT 0.0050 12.1365 0.0900 13.2300 ;
      RECT 8.6410 13.2165 8.7690 14.3100 ;
      RECT 8.6270 13.8820 8.7690 14.2045 ;
      RECT 8.4790 13.6090 8.5410 14.3100 ;
      RECT 8.4650 13.9185 8.5410 14.0720 ;
      RECT 8.4790 13.2165 8.5050 14.3100 ;
      RECT 8.4790 13.3375 8.5190 13.5770 ;
      RECT 8.4790 13.2165 8.5410 13.3055 ;
      RECT 8.1820 13.6670 8.3880 14.3100 ;
      RECT 8.3620 13.2165 8.3880 14.3100 ;
      RECT 8.1820 13.9440 8.4020 14.2020 ;
      RECT 8.1820 13.2165 8.2800 14.3100 ;
      RECT 7.7650 13.2165 7.8480 14.3100 ;
      RECT 7.7650 13.3050 7.8620 14.2405 ;
      RECT 16.4440 13.2165 16.5290 14.3100 ;
      RECT 16.3000 13.2165 16.3260 14.3100 ;
      RECT 16.1920 13.2165 16.2180 14.3100 ;
      RECT 16.0840 13.2165 16.1100 14.3100 ;
      RECT 15.9760 13.2165 16.0020 14.3100 ;
      RECT 15.8680 13.2165 15.8940 14.3100 ;
      RECT 15.7600 13.2165 15.7860 14.3100 ;
      RECT 15.6520 13.2165 15.6780 14.3100 ;
      RECT 15.5440 13.2165 15.5700 14.3100 ;
      RECT 15.4360 13.2165 15.4620 14.3100 ;
      RECT 15.3280 13.2165 15.3540 14.3100 ;
      RECT 15.2200 13.2165 15.2460 14.3100 ;
      RECT 15.1120 13.2165 15.1380 14.3100 ;
      RECT 15.0040 13.2165 15.0300 14.3100 ;
      RECT 14.8960 13.2165 14.9220 14.3100 ;
      RECT 14.7880 13.2165 14.8140 14.3100 ;
      RECT 14.6800 13.2165 14.7060 14.3100 ;
      RECT 14.5720 13.2165 14.5980 14.3100 ;
      RECT 14.4640 13.2165 14.4900 14.3100 ;
      RECT 14.3560 13.2165 14.3820 14.3100 ;
      RECT 14.2480 13.2165 14.2740 14.3100 ;
      RECT 14.1400 13.2165 14.1660 14.3100 ;
      RECT 14.0320 13.2165 14.0580 14.3100 ;
      RECT 13.9240 13.2165 13.9500 14.3100 ;
      RECT 13.8160 13.2165 13.8420 14.3100 ;
      RECT 13.7080 13.2165 13.7340 14.3100 ;
      RECT 13.6000 13.2165 13.6260 14.3100 ;
      RECT 13.4920 13.2165 13.5180 14.3100 ;
      RECT 13.3840 13.2165 13.4100 14.3100 ;
      RECT 13.2760 13.2165 13.3020 14.3100 ;
      RECT 13.1680 13.2165 13.1940 14.3100 ;
      RECT 13.0600 13.2165 13.0860 14.3100 ;
      RECT 12.9520 13.2165 12.9780 14.3100 ;
      RECT 12.8440 13.2165 12.8700 14.3100 ;
      RECT 12.7360 13.2165 12.7620 14.3100 ;
      RECT 12.6280 13.2165 12.6540 14.3100 ;
      RECT 12.5200 13.2165 12.5460 14.3100 ;
      RECT 12.4120 13.2165 12.4380 14.3100 ;
      RECT 12.3040 13.2165 12.3300 14.3100 ;
      RECT 12.1960 13.2165 12.2220 14.3100 ;
      RECT 12.0880 13.2165 12.1140 14.3100 ;
      RECT 11.9800 13.2165 12.0060 14.3100 ;
      RECT 11.8720 13.2165 11.8980 14.3100 ;
      RECT 11.7640 13.2165 11.7900 14.3100 ;
      RECT 11.6560 13.2165 11.6820 14.3100 ;
      RECT 11.5480 13.2165 11.5740 14.3100 ;
      RECT 11.4400 13.2165 11.4660 14.3100 ;
      RECT 11.3320 13.2165 11.3580 14.3100 ;
      RECT 11.2240 13.2165 11.2500 14.3100 ;
      RECT 11.1160 13.2165 11.1420 14.3100 ;
      RECT 11.0080 13.2165 11.0340 14.3100 ;
      RECT 10.9000 13.2165 10.9260 14.3100 ;
      RECT 10.7920 13.2165 10.8180 14.3100 ;
      RECT 10.6840 13.2165 10.7100 14.3100 ;
      RECT 10.5760 13.2165 10.6020 14.3100 ;
      RECT 10.4680 13.2165 10.4940 14.3100 ;
      RECT 10.3600 13.2165 10.3860 14.3100 ;
      RECT 10.2520 13.2165 10.2780 14.3100 ;
      RECT 10.1440 13.2165 10.1700 14.3100 ;
      RECT 10.0360 13.2165 10.0620 14.3100 ;
      RECT 9.9280 13.2165 9.9540 14.3100 ;
      RECT 9.8200 13.2165 9.8460 14.3100 ;
      RECT 9.7120 13.2165 9.7380 14.3100 ;
      RECT 9.6040 13.2165 9.6300 14.3100 ;
      RECT 9.4960 13.2165 9.5220 14.3100 ;
      RECT 9.3880 13.2165 9.4140 14.3100 ;
      RECT 9.1750 13.2165 9.2520 14.3100 ;
      RECT 7.2820 13.2165 7.3590 14.3100 ;
      RECT 7.1200 13.2165 7.1460 14.3100 ;
      RECT 7.0120 13.2165 7.0380 14.3100 ;
      RECT 6.9040 13.2165 6.9300 14.3100 ;
      RECT 6.7960 13.2165 6.8220 14.3100 ;
      RECT 6.6880 13.2165 6.7140 14.3100 ;
      RECT 6.5800 13.2165 6.6060 14.3100 ;
      RECT 6.4720 13.2165 6.4980 14.3100 ;
      RECT 6.3640 13.2165 6.3900 14.3100 ;
      RECT 6.2560 13.2165 6.2820 14.3100 ;
      RECT 6.1480 13.2165 6.1740 14.3100 ;
      RECT 6.0400 13.2165 6.0660 14.3100 ;
      RECT 5.9320 13.2165 5.9580 14.3100 ;
      RECT 5.8240 13.2165 5.8500 14.3100 ;
      RECT 5.7160 13.2165 5.7420 14.3100 ;
      RECT 5.6080 13.2165 5.6340 14.3100 ;
      RECT 5.5000 13.2165 5.5260 14.3100 ;
      RECT 5.3920 13.2165 5.4180 14.3100 ;
      RECT 5.2840 13.2165 5.3100 14.3100 ;
      RECT 5.1760 13.2165 5.2020 14.3100 ;
      RECT 5.0680 13.2165 5.0940 14.3100 ;
      RECT 4.9600 13.2165 4.9860 14.3100 ;
      RECT 4.8520 13.2165 4.8780 14.3100 ;
      RECT 4.7440 13.2165 4.7700 14.3100 ;
      RECT 4.6360 13.2165 4.6620 14.3100 ;
      RECT 4.5280 13.2165 4.5540 14.3100 ;
      RECT 4.4200 13.2165 4.4460 14.3100 ;
      RECT 4.3120 13.2165 4.3380 14.3100 ;
      RECT 4.2040 13.2165 4.2300 14.3100 ;
      RECT 4.0960 13.2165 4.1220 14.3100 ;
      RECT 3.9880 13.2165 4.0140 14.3100 ;
      RECT 3.8800 13.2165 3.9060 14.3100 ;
      RECT 3.7720 13.2165 3.7980 14.3100 ;
      RECT 3.6640 13.2165 3.6900 14.3100 ;
      RECT 3.5560 13.2165 3.5820 14.3100 ;
      RECT 3.4480 13.2165 3.4740 14.3100 ;
      RECT 3.3400 13.2165 3.3660 14.3100 ;
      RECT 3.2320 13.2165 3.2580 14.3100 ;
      RECT 3.1240 13.2165 3.1500 14.3100 ;
      RECT 3.0160 13.2165 3.0420 14.3100 ;
      RECT 2.9080 13.2165 2.9340 14.3100 ;
      RECT 2.8000 13.2165 2.8260 14.3100 ;
      RECT 2.6920 13.2165 2.7180 14.3100 ;
      RECT 2.5840 13.2165 2.6100 14.3100 ;
      RECT 2.4760 13.2165 2.5020 14.3100 ;
      RECT 2.3680 13.2165 2.3940 14.3100 ;
      RECT 2.2600 13.2165 2.2860 14.3100 ;
      RECT 2.1520 13.2165 2.1780 14.3100 ;
      RECT 2.0440 13.2165 2.0700 14.3100 ;
      RECT 1.9360 13.2165 1.9620 14.3100 ;
      RECT 1.8280 13.2165 1.8540 14.3100 ;
      RECT 1.7200 13.2165 1.7460 14.3100 ;
      RECT 1.6120 13.2165 1.6380 14.3100 ;
      RECT 1.5040 13.2165 1.5300 14.3100 ;
      RECT 1.3960 13.2165 1.4220 14.3100 ;
      RECT 1.2880 13.2165 1.3140 14.3100 ;
      RECT 1.1800 13.2165 1.2060 14.3100 ;
      RECT 1.0720 13.2165 1.0980 14.3100 ;
      RECT 0.9640 13.2165 0.9900 14.3100 ;
      RECT 0.8560 13.2165 0.8820 14.3100 ;
      RECT 0.7480 13.2165 0.7740 14.3100 ;
      RECT 0.6400 13.2165 0.6660 14.3100 ;
      RECT 0.5320 13.2165 0.5580 14.3100 ;
      RECT 0.4240 13.2165 0.4500 14.3100 ;
      RECT 0.3160 13.2165 0.3420 14.3100 ;
      RECT 0.2080 13.2165 0.2340 14.3100 ;
      RECT 0.0050 13.2165 0.0900 14.3100 ;
      RECT 8.6410 14.2965 8.7690 15.3900 ;
      RECT 8.6270 14.9620 8.7690 15.2845 ;
      RECT 8.4790 14.6890 8.5410 15.3900 ;
      RECT 8.4650 14.9985 8.5410 15.1520 ;
      RECT 8.4790 14.2965 8.5050 15.3900 ;
      RECT 8.4790 14.4175 8.5190 14.6570 ;
      RECT 8.4790 14.2965 8.5410 14.3855 ;
      RECT 8.1820 14.7470 8.3880 15.3900 ;
      RECT 8.3620 14.2965 8.3880 15.3900 ;
      RECT 8.1820 15.0240 8.4020 15.2820 ;
      RECT 8.1820 14.2965 8.2800 15.3900 ;
      RECT 7.7650 14.2965 7.8480 15.3900 ;
      RECT 7.7650 14.3850 7.8620 15.3205 ;
      RECT 16.4440 14.2965 16.5290 15.3900 ;
      RECT 16.3000 14.2965 16.3260 15.3900 ;
      RECT 16.1920 14.2965 16.2180 15.3900 ;
      RECT 16.0840 14.2965 16.1100 15.3900 ;
      RECT 15.9760 14.2965 16.0020 15.3900 ;
      RECT 15.8680 14.2965 15.8940 15.3900 ;
      RECT 15.7600 14.2965 15.7860 15.3900 ;
      RECT 15.6520 14.2965 15.6780 15.3900 ;
      RECT 15.5440 14.2965 15.5700 15.3900 ;
      RECT 15.4360 14.2965 15.4620 15.3900 ;
      RECT 15.3280 14.2965 15.3540 15.3900 ;
      RECT 15.2200 14.2965 15.2460 15.3900 ;
      RECT 15.1120 14.2965 15.1380 15.3900 ;
      RECT 15.0040 14.2965 15.0300 15.3900 ;
      RECT 14.8960 14.2965 14.9220 15.3900 ;
      RECT 14.7880 14.2965 14.8140 15.3900 ;
      RECT 14.6800 14.2965 14.7060 15.3900 ;
      RECT 14.5720 14.2965 14.5980 15.3900 ;
      RECT 14.4640 14.2965 14.4900 15.3900 ;
      RECT 14.3560 14.2965 14.3820 15.3900 ;
      RECT 14.2480 14.2965 14.2740 15.3900 ;
      RECT 14.1400 14.2965 14.1660 15.3900 ;
      RECT 14.0320 14.2965 14.0580 15.3900 ;
      RECT 13.9240 14.2965 13.9500 15.3900 ;
      RECT 13.8160 14.2965 13.8420 15.3900 ;
      RECT 13.7080 14.2965 13.7340 15.3900 ;
      RECT 13.6000 14.2965 13.6260 15.3900 ;
      RECT 13.4920 14.2965 13.5180 15.3900 ;
      RECT 13.3840 14.2965 13.4100 15.3900 ;
      RECT 13.2760 14.2965 13.3020 15.3900 ;
      RECT 13.1680 14.2965 13.1940 15.3900 ;
      RECT 13.0600 14.2965 13.0860 15.3900 ;
      RECT 12.9520 14.2965 12.9780 15.3900 ;
      RECT 12.8440 14.2965 12.8700 15.3900 ;
      RECT 12.7360 14.2965 12.7620 15.3900 ;
      RECT 12.6280 14.2965 12.6540 15.3900 ;
      RECT 12.5200 14.2965 12.5460 15.3900 ;
      RECT 12.4120 14.2965 12.4380 15.3900 ;
      RECT 12.3040 14.2965 12.3300 15.3900 ;
      RECT 12.1960 14.2965 12.2220 15.3900 ;
      RECT 12.0880 14.2965 12.1140 15.3900 ;
      RECT 11.9800 14.2965 12.0060 15.3900 ;
      RECT 11.8720 14.2965 11.8980 15.3900 ;
      RECT 11.7640 14.2965 11.7900 15.3900 ;
      RECT 11.6560 14.2965 11.6820 15.3900 ;
      RECT 11.5480 14.2965 11.5740 15.3900 ;
      RECT 11.4400 14.2965 11.4660 15.3900 ;
      RECT 11.3320 14.2965 11.3580 15.3900 ;
      RECT 11.2240 14.2965 11.2500 15.3900 ;
      RECT 11.1160 14.2965 11.1420 15.3900 ;
      RECT 11.0080 14.2965 11.0340 15.3900 ;
      RECT 10.9000 14.2965 10.9260 15.3900 ;
      RECT 10.7920 14.2965 10.8180 15.3900 ;
      RECT 10.6840 14.2965 10.7100 15.3900 ;
      RECT 10.5760 14.2965 10.6020 15.3900 ;
      RECT 10.4680 14.2965 10.4940 15.3900 ;
      RECT 10.3600 14.2965 10.3860 15.3900 ;
      RECT 10.2520 14.2965 10.2780 15.3900 ;
      RECT 10.1440 14.2965 10.1700 15.3900 ;
      RECT 10.0360 14.2965 10.0620 15.3900 ;
      RECT 9.9280 14.2965 9.9540 15.3900 ;
      RECT 9.8200 14.2965 9.8460 15.3900 ;
      RECT 9.7120 14.2965 9.7380 15.3900 ;
      RECT 9.6040 14.2965 9.6300 15.3900 ;
      RECT 9.4960 14.2965 9.5220 15.3900 ;
      RECT 9.3880 14.2965 9.4140 15.3900 ;
      RECT 9.1750 14.2965 9.2520 15.3900 ;
      RECT 7.2820 14.2965 7.3590 15.3900 ;
      RECT 7.1200 14.2965 7.1460 15.3900 ;
      RECT 7.0120 14.2965 7.0380 15.3900 ;
      RECT 6.9040 14.2965 6.9300 15.3900 ;
      RECT 6.7960 14.2965 6.8220 15.3900 ;
      RECT 6.6880 14.2965 6.7140 15.3900 ;
      RECT 6.5800 14.2965 6.6060 15.3900 ;
      RECT 6.4720 14.2965 6.4980 15.3900 ;
      RECT 6.3640 14.2965 6.3900 15.3900 ;
      RECT 6.2560 14.2965 6.2820 15.3900 ;
      RECT 6.1480 14.2965 6.1740 15.3900 ;
      RECT 6.0400 14.2965 6.0660 15.3900 ;
      RECT 5.9320 14.2965 5.9580 15.3900 ;
      RECT 5.8240 14.2965 5.8500 15.3900 ;
      RECT 5.7160 14.2965 5.7420 15.3900 ;
      RECT 5.6080 14.2965 5.6340 15.3900 ;
      RECT 5.5000 14.2965 5.5260 15.3900 ;
      RECT 5.3920 14.2965 5.4180 15.3900 ;
      RECT 5.2840 14.2965 5.3100 15.3900 ;
      RECT 5.1760 14.2965 5.2020 15.3900 ;
      RECT 5.0680 14.2965 5.0940 15.3900 ;
      RECT 4.9600 14.2965 4.9860 15.3900 ;
      RECT 4.8520 14.2965 4.8780 15.3900 ;
      RECT 4.7440 14.2965 4.7700 15.3900 ;
      RECT 4.6360 14.2965 4.6620 15.3900 ;
      RECT 4.5280 14.2965 4.5540 15.3900 ;
      RECT 4.4200 14.2965 4.4460 15.3900 ;
      RECT 4.3120 14.2965 4.3380 15.3900 ;
      RECT 4.2040 14.2965 4.2300 15.3900 ;
      RECT 4.0960 14.2965 4.1220 15.3900 ;
      RECT 3.9880 14.2965 4.0140 15.3900 ;
      RECT 3.8800 14.2965 3.9060 15.3900 ;
      RECT 3.7720 14.2965 3.7980 15.3900 ;
      RECT 3.6640 14.2965 3.6900 15.3900 ;
      RECT 3.5560 14.2965 3.5820 15.3900 ;
      RECT 3.4480 14.2965 3.4740 15.3900 ;
      RECT 3.3400 14.2965 3.3660 15.3900 ;
      RECT 3.2320 14.2965 3.2580 15.3900 ;
      RECT 3.1240 14.2965 3.1500 15.3900 ;
      RECT 3.0160 14.2965 3.0420 15.3900 ;
      RECT 2.9080 14.2965 2.9340 15.3900 ;
      RECT 2.8000 14.2965 2.8260 15.3900 ;
      RECT 2.6920 14.2965 2.7180 15.3900 ;
      RECT 2.5840 14.2965 2.6100 15.3900 ;
      RECT 2.4760 14.2965 2.5020 15.3900 ;
      RECT 2.3680 14.2965 2.3940 15.3900 ;
      RECT 2.2600 14.2965 2.2860 15.3900 ;
      RECT 2.1520 14.2965 2.1780 15.3900 ;
      RECT 2.0440 14.2965 2.0700 15.3900 ;
      RECT 1.9360 14.2965 1.9620 15.3900 ;
      RECT 1.8280 14.2965 1.8540 15.3900 ;
      RECT 1.7200 14.2965 1.7460 15.3900 ;
      RECT 1.6120 14.2965 1.6380 15.3900 ;
      RECT 1.5040 14.2965 1.5300 15.3900 ;
      RECT 1.3960 14.2965 1.4220 15.3900 ;
      RECT 1.2880 14.2965 1.3140 15.3900 ;
      RECT 1.1800 14.2965 1.2060 15.3900 ;
      RECT 1.0720 14.2965 1.0980 15.3900 ;
      RECT 0.9640 14.2965 0.9900 15.3900 ;
      RECT 0.8560 14.2965 0.8820 15.3900 ;
      RECT 0.7480 14.2965 0.7740 15.3900 ;
      RECT 0.6400 14.2965 0.6660 15.3900 ;
      RECT 0.5320 14.2965 0.5580 15.3900 ;
      RECT 0.4240 14.2965 0.4500 15.3900 ;
      RECT 0.3160 14.2965 0.3420 15.3900 ;
      RECT 0.2080 14.2965 0.2340 15.3900 ;
      RECT 0.0050 14.2965 0.0900 15.3900 ;
      RECT 8.6410 15.3765 8.7690 16.4700 ;
      RECT 8.6270 16.0420 8.7690 16.3645 ;
      RECT 8.4790 15.7690 8.5410 16.4700 ;
      RECT 8.4650 16.0785 8.5410 16.2320 ;
      RECT 8.4790 15.3765 8.5050 16.4700 ;
      RECT 8.4790 15.4975 8.5190 15.7370 ;
      RECT 8.4790 15.3765 8.5410 15.4655 ;
      RECT 8.1820 15.8270 8.3880 16.4700 ;
      RECT 8.3620 15.3765 8.3880 16.4700 ;
      RECT 8.1820 16.1040 8.4020 16.3620 ;
      RECT 8.1820 15.3765 8.2800 16.4700 ;
      RECT 7.7650 15.3765 7.8480 16.4700 ;
      RECT 7.7650 15.4650 7.8620 16.4005 ;
      RECT 16.4440 15.3765 16.5290 16.4700 ;
      RECT 16.3000 15.3765 16.3260 16.4700 ;
      RECT 16.1920 15.3765 16.2180 16.4700 ;
      RECT 16.0840 15.3765 16.1100 16.4700 ;
      RECT 15.9760 15.3765 16.0020 16.4700 ;
      RECT 15.8680 15.3765 15.8940 16.4700 ;
      RECT 15.7600 15.3765 15.7860 16.4700 ;
      RECT 15.6520 15.3765 15.6780 16.4700 ;
      RECT 15.5440 15.3765 15.5700 16.4700 ;
      RECT 15.4360 15.3765 15.4620 16.4700 ;
      RECT 15.3280 15.3765 15.3540 16.4700 ;
      RECT 15.2200 15.3765 15.2460 16.4700 ;
      RECT 15.1120 15.3765 15.1380 16.4700 ;
      RECT 15.0040 15.3765 15.0300 16.4700 ;
      RECT 14.8960 15.3765 14.9220 16.4700 ;
      RECT 14.7880 15.3765 14.8140 16.4700 ;
      RECT 14.6800 15.3765 14.7060 16.4700 ;
      RECT 14.5720 15.3765 14.5980 16.4700 ;
      RECT 14.4640 15.3765 14.4900 16.4700 ;
      RECT 14.3560 15.3765 14.3820 16.4700 ;
      RECT 14.2480 15.3765 14.2740 16.4700 ;
      RECT 14.1400 15.3765 14.1660 16.4700 ;
      RECT 14.0320 15.3765 14.0580 16.4700 ;
      RECT 13.9240 15.3765 13.9500 16.4700 ;
      RECT 13.8160 15.3765 13.8420 16.4700 ;
      RECT 13.7080 15.3765 13.7340 16.4700 ;
      RECT 13.6000 15.3765 13.6260 16.4700 ;
      RECT 13.4920 15.3765 13.5180 16.4700 ;
      RECT 13.3840 15.3765 13.4100 16.4700 ;
      RECT 13.2760 15.3765 13.3020 16.4700 ;
      RECT 13.1680 15.3765 13.1940 16.4700 ;
      RECT 13.0600 15.3765 13.0860 16.4700 ;
      RECT 12.9520 15.3765 12.9780 16.4700 ;
      RECT 12.8440 15.3765 12.8700 16.4700 ;
      RECT 12.7360 15.3765 12.7620 16.4700 ;
      RECT 12.6280 15.3765 12.6540 16.4700 ;
      RECT 12.5200 15.3765 12.5460 16.4700 ;
      RECT 12.4120 15.3765 12.4380 16.4700 ;
      RECT 12.3040 15.3765 12.3300 16.4700 ;
      RECT 12.1960 15.3765 12.2220 16.4700 ;
      RECT 12.0880 15.3765 12.1140 16.4700 ;
      RECT 11.9800 15.3765 12.0060 16.4700 ;
      RECT 11.8720 15.3765 11.8980 16.4700 ;
      RECT 11.7640 15.3765 11.7900 16.4700 ;
      RECT 11.6560 15.3765 11.6820 16.4700 ;
      RECT 11.5480 15.3765 11.5740 16.4700 ;
      RECT 11.4400 15.3765 11.4660 16.4700 ;
      RECT 11.3320 15.3765 11.3580 16.4700 ;
      RECT 11.2240 15.3765 11.2500 16.4700 ;
      RECT 11.1160 15.3765 11.1420 16.4700 ;
      RECT 11.0080 15.3765 11.0340 16.4700 ;
      RECT 10.9000 15.3765 10.9260 16.4700 ;
      RECT 10.7920 15.3765 10.8180 16.4700 ;
      RECT 10.6840 15.3765 10.7100 16.4700 ;
      RECT 10.5760 15.3765 10.6020 16.4700 ;
      RECT 10.4680 15.3765 10.4940 16.4700 ;
      RECT 10.3600 15.3765 10.3860 16.4700 ;
      RECT 10.2520 15.3765 10.2780 16.4700 ;
      RECT 10.1440 15.3765 10.1700 16.4700 ;
      RECT 10.0360 15.3765 10.0620 16.4700 ;
      RECT 9.9280 15.3765 9.9540 16.4700 ;
      RECT 9.8200 15.3765 9.8460 16.4700 ;
      RECT 9.7120 15.3765 9.7380 16.4700 ;
      RECT 9.6040 15.3765 9.6300 16.4700 ;
      RECT 9.4960 15.3765 9.5220 16.4700 ;
      RECT 9.3880 15.3765 9.4140 16.4700 ;
      RECT 9.1750 15.3765 9.2520 16.4700 ;
      RECT 7.2820 15.3765 7.3590 16.4700 ;
      RECT 7.1200 15.3765 7.1460 16.4700 ;
      RECT 7.0120 15.3765 7.0380 16.4700 ;
      RECT 6.9040 15.3765 6.9300 16.4700 ;
      RECT 6.7960 15.3765 6.8220 16.4700 ;
      RECT 6.6880 15.3765 6.7140 16.4700 ;
      RECT 6.5800 15.3765 6.6060 16.4700 ;
      RECT 6.4720 15.3765 6.4980 16.4700 ;
      RECT 6.3640 15.3765 6.3900 16.4700 ;
      RECT 6.2560 15.3765 6.2820 16.4700 ;
      RECT 6.1480 15.3765 6.1740 16.4700 ;
      RECT 6.0400 15.3765 6.0660 16.4700 ;
      RECT 5.9320 15.3765 5.9580 16.4700 ;
      RECT 5.8240 15.3765 5.8500 16.4700 ;
      RECT 5.7160 15.3765 5.7420 16.4700 ;
      RECT 5.6080 15.3765 5.6340 16.4700 ;
      RECT 5.5000 15.3765 5.5260 16.4700 ;
      RECT 5.3920 15.3765 5.4180 16.4700 ;
      RECT 5.2840 15.3765 5.3100 16.4700 ;
      RECT 5.1760 15.3765 5.2020 16.4700 ;
      RECT 5.0680 15.3765 5.0940 16.4700 ;
      RECT 4.9600 15.3765 4.9860 16.4700 ;
      RECT 4.8520 15.3765 4.8780 16.4700 ;
      RECT 4.7440 15.3765 4.7700 16.4700 ;
      RECT 4.6360 15.3765 4.6620 16.4700 ;
      RECT 4.5280 15.3765 4.5540 16.4700 ;
      RECT 4.4200 15.3765 4.4460 16.4700 ;
      RECT 4.3120 15.3765 4.3380 16.4700 ;
      RECT 4.2040 15.3765 4.2300 16.4700 ;
      RECT 4.0960 15.3765 4.1220 16.4700 ;
      RECT 3.9880 15.3765 4.0140 16.4700 ;
      RECT 3.8800 15.3765 3.9060 16.4700 ;
      RECT 3.7720 15.3765 3.7980 16.4700 ;
      RECT 3.6640 15.3765 3.6900 16.4700 ;
      RECT 3.5560 15.3765 3.5820 16.4700 ;
      RECT 3.4480 15.3765 3.4740 16.4700 ;
      RECT 3.3400 15.3765 3.3660 16.4700 ;
      RECT 3.2320 15.3765 3.2580 16.4700 ;
      RECT 3.1240 15.3765 3.1500 16.4700 ;
      RECT 3.0160 15.3765 3.0420 16.4700 ;
      RECT 2.9080 15.3765 2.9340 16.4700 ;
      RECT 2.8000 15.3765 2.8260 16.4700 ;
      RECT 2.6920 15.3765 2.7180 16.4700 ;
      RECT 2.5840 15.3765 2.6100 16.4700 ;
      RECT 2.4760 15.3765 2.5020 16.4700 ;
      RECT 2.3680 15.3765 2.3940 16.4700 ;
      RECT 2.2600 15.3765 2.2860 16.4700 ;
      RECT 2.1520 15.3765 2.1780 16.4700 ;
      RECT 2.0440 15.3765 2.0700 16.4700 ;
      RECT 1.9360 15.3765 1.9620 16.4700 ;
      RECT 1.8280 15.3765 1.8540 16.4700 ;
      RECT 1.7200 15.3765 1.7460 16.4700 ;
      RECT 1.6120 15.3765 1.6380 16.4700 ;
      RECT 1.5040 15.3765 1.5300 16.4700 ;
      RECT 1.3960 15.3765 1.4220 16.4700 ;
      RECT 1.2880 15.3765 1.3140 16.4700 ;
      RECT 1.1800 15.3765 1.2060 16.4700 ;
      RECT 1.0720 15.3765 1.0980 16.4700 ;
      RECT 0.9640 15.3765 0.9900 16.4700 ;
      RECT 0.8560 15.3765 0.8820 16.4700 ;
      RECT 0.7480 15.3765 0.7740 16.4700 ;
      RECT 0.6400 15.3765 0.6660 16.4700 ;
      RECT 0.5320 15.3765 0.5580 16.4700 ;
      RECT 0.4240 15.3765 0.4500 16.4700 ;
      RECT 0.3160 15.3765 0.3420 16.4700 ;
      RECT 0.2080 15.3765 0.2340 16.4700 ;
      RECT 0.0050 15.3765 0.0900 16.4700 ;
      RECT 8.6410 16.4565 8.7690 17.5500 ;
      RECT 8.6270 17.1220 8.7690 17.4445 ;
      RECT 8.4790 16.8490 8.5410 17.5500 ;
      RECT 8.4650 17.1585 8.5410 17.3120 ;
      RECT 8.4790 16.4565 8.5050 17.5500 ;
      RECT 8.4790 16.5775 8.5190 16.8170 ;
      RECT 8.4790 16.4565 8.5410 16.5455 ;
      RECT 8.1820 16.9070 8.3880 17.5500 ;
      RECT 8.3620 16.4565 8.3880 17.5500 ;
      RECT 8.1820 17.1840 8.4020 17.4420 ;
      RECT 8.1820 16.4565 8.2800 17.5500 ;
      RECT 7.7650 16.4565 7.8480 17.5500 ;
      RECT 7.7650 16.5450 7.8620 17.4805 ;
      RECT 16.4440 16.4565 16.5290 17.5500 ;
      RECT 16.3000 16.4565 16.3260 17.5500 ;
      RECT 16.1920 16.4565 16.2180 17.5500 ;
      RECT 16.0840 16.4565 16.1100 17.5500 ;
      RECT 15.9760 16.4565 16.0020 17.5500 ;
      RECT 15.8680 16.4565 15.8940 17.5500 ;
      RECT 15.7600 16.4565 15.7860 17.5500 ;
      RECT 15.6520 16.4565 15.6780 17.5500 ;
      RECT 15.5440 16.4565 15.5700 17.5500 ;
      RECT 15.4360 16.4565 15.4620 17.5500 ;
      RECT 15.3280 16.4565 15.3540 17.5500 ;
      RECT 15.2200 16.4565 15.2460 17.5500 ;
      RECT 15.1120 16.4565 15.1380 17.5500 ;
      RECT 15.0040 16.4565 15.0300 17.5500 ;
      RECT 14.8960 16.4565 14.9220 17.5500 ;
      RECT 14.7880 16.4565 14.8140 17.5500 ;
      RECT 14.6800 16.4565 14.7060 17.5500 ;
      RECT 14.5720 16.4565 14.5980 17.5500 ;
      RECT 14.4640 16.4565 14.4900 17.5500 ;
      RECT 14.3560 16.4565 14.3820 17.5500 ;
      RECT 14.2480 16.4565 14.2740 17.5500 ;
      RECT 14.1400 16.4565 14.1660 17.5500 ;
      RECT 14.0320 16.4565 14.0580 17.5500 ;
      RECT 13.9240 16.4565 13.9500 17.5500 ;
      RECT 13.8160 16.4565 13.8420 17.5500 ;
      RECT 13.7080 16.4565 13.7340 17.5500 ;
      RECT 13.6000 16.4565 13.6260 17.5500 ;
      RECT 13.4920 16.4565 13.5180 17.5500 ;
      RECT 13.3840 16.4565 13.4100 17.5500 ;
      RECT 13.2760 16.4565 13.3020 17.5500 ;
      RECT 13.1680 16.4565 13.1940 17.5500 ;
      RECT 13.0600 16.4565 13.0860 17.5500 ;
      RECT 12.9520 16.4565 12.9780 17.5500 ;
      RECT 12.8440 16.4565 12.8700 17.5500 ;
      RECT 12.7360 16.4565 12.7620 17.5500 ;
      RECT 12.6280 16.4565 12.6540 17.5500 ;
      RECT 12.5200 16.4565 12.5460 17.5500 ;
      RECT 12.4120 16.4565 12.4380 17.5500 ;
      RECT 12.3040 16.4565 12.3300 17.5500 ;
      RECT 12.1960 16.4565 12.2220 17.5500 ;
      RECT 12.0880 16.4565 12.1140 17.5500 ;
      RECT 11.9800 16.4565 12.0060 17.5500 ;
      RECT 11.8720 16.4565 11.8980 17.5500 ;
      RECT 11.7640 16.4565 11.7900 17.5500 ;
      RECT 11.6560 16.4565 11.6820 17.5500 ;
      RECT 11.5480 16.4565 11.5740 17.5500 ;
      RECT 11.4400 16.4565 11.4660 17.5500 ;
      RECT 11.3320 16.4565 11.3580 17.5500 ;
      RECT 11.2240 16.4565 11.2500 17.5500 ;
      RECT 11.1160 16.4565 11.1420 17.5500 ;
      RECT 11.0080 16.4565 11.0340 17.5500 ;
      RECT 10.9000 16.4565 10.9260 17.5500 ;
      RECT 10.7920 16.4565 10.8180 17.5500 ;
      RECT 10.6840 16.4565 10.7100 17.5500 ;
      RECT 10.5760 16.4565 10.6020 17.5500 ;
      RECT 10.4680 16.4565 10.4940 17.5500 ;
      RECT 10.3600 16.4565 10.3860 17.5500 ;
      RECT 10.2520 16.4565 10.2780 17.5500 ;
      RECT 10.1440 16.4565 10.1700 17.5500 ;
      RECT 10.0360 16.4565 10.0620 17.5500 ;
      RECT 9.9280 16.4565 9.9540 17.5500 ;
      RECT 9.8200 16.4565 9.8460 17.5500 ;
      RECT 9.7120 16.4565 9.7380 17.5500 ;
      RECT 9.6040 16.4565 9.6300 17.5500 ;
      RECT 9.4960 16.4565 9.5220 17.5500 ;
      RECT 9.3880 16.4565 9.4140 17.5500 ;
      RECT 9.1750 16.4565 9.2520 17.5500 ;
      RECT 7.2820 16.4565 7.3590 17.5500 ;
      RECT 7.1200 16.4565 7.1460 17.5500 ;
      RECT 7.0120 16.4565 7.0380 17.5500 ;
      RECT 6.9040 16.4565 6.9300 17.5500 ;
      RECT 6.7960 16.4565 6.8220 17.5500 ;
      RECT 6.6880 16.4565 6.7140 17.5500 ;
      RECT 6.5800 16.4565 6.6060 17.5500 ;
      RECT 6.4720 16.4565 6.4980 17.5500 ;
      RECT 6.3640 16.4565 6.3900 17.5500 ;
      RECT 6.2560 16.4565 6.2820 17.5500 ;
      RECT 6.1480 16.4565 6.1740 17.5500 ;
      RECT 6.0400 16.4565 6.0660 17.5500 ;
      RECT 5.9320 16.4565 5.9580 17.5500 ;
      RECT 5.8240 16.4565 5.8500 17.5500 ;
      RECT 5.7160 16.4565 5.7420 17.5500 ;
      RECT 5.6080 16.4565 5.6340 17.5500 ;
      RECT 5.5000 16.4565 5.5260 17.5500 ;
      RECT 5.3920 16.4565 5.4180 17.5500 ;
      RECT 5.2840 16.4565 5.3100 17.5500 ;
      RECT 5.1760 16.4565 5.2020 17.5500 ;
      RECT 5.0680 16.4565 5.0940 17.5500 ;
      RECT 4.9600 16.4565 4.9860 17.5500 ;
      RECT 4.8520 16.4565 4.8780 17.5500 ;
      RECT 4.7440 16.4565 4.7700 17.5500 ;
      RECT 4.6360 16.4565 4.6620 17.5500 ;
      RECT 4.5280 16.4565 4.5540 17.5500 ;
      RECT 4.4200 16.4565 4.4460 17.5500 ;
      RECT 4.3120 16.4565 4.3380 17.5500 ;
      RECT 4.2040 16.4565 4.2300 17.5500 ;
      RECT 4.0960 16.4565 4.1220 17.5500 ;
      RECT 3.9880 16.4565 4.0140 17.5500 ;
      RECT 3.8800 16.4565 3.9060 17.5500 ;
      RECT 3.7720 16.4565 3.7980 17.5500 ;
      RECT 3.6640 16.4565 3.6900 17.5500 ;
      RECT 3.5560 16.4565 3.5820 17.5500 ;
      RECT 3.4480 16.4565 3.4740 17.5500 ;
      RECT 3.3400 16.4565 3.3660 17.5500 ;
      RECT 3.2320 16.4565 3.2580 17.5500 ;
      RECT 3.1240 16.4565 3.1500 17.5500 ;
      RECT 3.0160 16.4565 3.0420 17.5500 ;
      RECT 2.9080 16.4565 2.9340 17.5500 ;
      RECT 2.8000 16.4565 2.8260 17.5500 ;
      RECT 2.6920 16.4565 2.7180 17.5500 ;
      RECT 2.5840 16.4565 2.6100 17.5500 ;
      RECT 2.4760 16.4565 2.5020 17.5500 ;
      RECT 2.3680 16.4565 2.3940 17.5500 ;
      RECT 2.2600 16.4565 2.2860 17.5500 ;
      RECT 2.1520 16.4565 2.1780 17.5500 ;
      RECT 2.0440 16.4565 2.0700 17.5500 ;
      RECT 1.9360 16.4565 1.9620 17.5500 ;
      RECT 1.8280 16.4565 1.8540 17.5500 ;
      RECT 1.7200 16.4565 1.7460 17.5500 ;
      RECT 1.6120 16.4565 1.6380 17.5500 ;
      RECT 1.5040 16.4565 1.5300 17.5500 ;
      RECT 1.3960 16.4565 1.4220 17.5500 ;
      RECT 1.2880 16.4565 1.3140 17.5500 ;
      RECT 1.1800 16.4565 1.2060 17.5500 ;
      RECT 1.0720 16.4565 1.0980 17.5500 ;
      RECT 0.9640 16.4565 0.9900 17.5500 ;
      RECT 0.8560 16.4565 0.8820 17.5500 ;
      RECT 0.7480 16.4565 0.7740 17.5500 ;
      RECT 0.6400 16.4565 0.6660 17.5500 ;
      RECT 0.5320 16.4565 0.5580 17.5500 ;
      RECT 0.4240 16.4565 0.4500 17.5500 ;
      RECT 0.3160 16.4565 0.3420 17.5500 ;
      RECT 0.2080 16.4565 0.2340 17.5500 ;
      RECT 0.0050 16.4565 0.0900 17.5500 ;
      RECT 8.6410 17.5365 8.7690 18.6300 ;
      RECT 8.6270 18.2020 8.7690 18.5245 ;
      RECT 8.4790 17.9290 8.5410 18.6300 ;
      RECT 8.4650 18.2385 8.5410 18.3920 ;
      RECT 8.4790 17.5365 8.5050 18.6300 ;
      RECT 8.4790 17.6575 8.5190 17.8970 ;
      RECT 8.4790 17.5365 8.5410 17.6255 ;
      RECT 8.1820 17.9870 8.3880 18.6300 ;
      RECT 8.3620 17.5365 8.3880 18.6300 ;
      RECT 8.1820 18.2640 8.4020 18.5220 ;
      RECT 8.1820 17.5365 8.2800 18.6300 ;
      RECT 7.7650 17.5365 7.8480 18.6300 ;
      RECT 7.7650 17.6250 7.8620 18.5605 ;
      RECT 16.4440 17.5365 16.5290 18.6300 ;
      RECT 16.3000 17.5365 16.3260 18.6300 ;
      RECT 16.1920 17.5365 16.2180 18.6300 ;
      RECT 16.0840 17.5365 16.1100 18.6300 ;
      RECT 15.9760 17.5365 16.0020 18.6300 ;
      RECT 15.8680 17.5365 15.8940 18.6300 ;
      RECT 15.7600 17.5365 15.7860 18.6300 ;
      RECT 15.6520 17.5365 15.6780 18.6300 ;
      RECT 15.5440 17.5365 15.5700 18.6300 ;
      RECT 15.4360 17.5365 15.4620 18.6300 ;
      RECT 15.3280 17.5365 15.3540 18.6300 ;
      RECT 15.2200 17.5365 15.2460 18.6300 ;
      RECT 15.1120 17.5365 15.1380 18.6300 ;
      RECT 15.0040 17.5365 15.0300 18.6300 ;
      RECT 14.8960 17.5365 14.9220 18.6300 ;
      RECT 14.7880 17.5365 14.8140 18.6300 ;
      RECT 14.6800 17.5365 14.7060 18.6300 ;
      RECT 14.5720 17.5365 14.5980 18.6300 ;
      RECT 14.4640 17.5365 14.4900 18.6300 ;
      RECT 14.3560 17.5365 14.3820 18.6300 ;
      RECT 14.2480 17.5365 14.2740 18.6300 ;
      RECT 14.1400 17.5365 14.1660 18.6300 ;
      RECT 14.0320 17.5365 14.0580 18.6300 ;
      RECT 13.9240 17.5365 13.9500 18.6300 ;
      RECT 13.8160 17.5365 13.8420 18.6300 ;
      RECT 13.7080 17.5365 13.7340 18.6300 ;
      RECT 13.6000 17.5365 13.6260 18.6300 ;
      RECT 13.4920 17.5365 13.5180 18.6300 ;
      RECT 13.3840 17.5365 13.4100 18.6300 ;
      RECT 13.2760 17.5365 13.3020 18.6300 ;
      RECT 13.1680 17.5365 13.1940 18.6300 ;
      RECT 13.0600 17.5365 13.0860 18.6300 ;
      RECT 12.9520 17.5365 12.9780 18.6300 ;
      RECT 12.8440 17.5365 12.8700 18.6300 ;
      RECT 12.7360 17.5365 12.7620 18.6300 ;
      RECT 12.6280 17.5365 12.6540 18.6300 ;
      RECT 12.5200 17.5365 12.5460 18.6300 ;
      RECT 12.4120 17.5365 12.4380 18.6300 ;
      RECT 12.3040 17.5365 12.3300 18.6300 ;
      RECT 12.1960 17.5365 12.2220 18.6300 ;
      RECT 12.0880 17.5365 12.1140 18.6300 ;
      RECT 11.9800 17.5365 12.0060 18.6300 ;
      RECT 11.8720 17.5365 11.8980 18.6300 ;
      RECT 11.7640 17.5365 11.7900 18.6300 ;
      RECT 11.6560 17.5365 11.6820 18.6300 ;
      RECT 11.5480 17.5365 11.5740 18.6300 ;
      RECT 11.4400 17.5365 11.4660 18.6300 ;
      RECT 11.3320 17.5365 11.3580 18.6300 ;
      RECT 11.2240 17.5365 11.2500 18.6300 ;
      RECT 11.1160 17.5365 11.1420 18.6300 ;
      RECT 11.0080 17.5365 11.0340 18.6300 ;
      RECT 10.9000 17.5365 10.9260 18.6300 ;
      RECT 10.7920 17.5365 10.8180 18.6300 ;
      RECT 10.6840 17.5365 10.7100 18.6300 ;
      RECT 10.5760 17.5365 10.6020 18.6300 ;
      RECT 10.4680 17.5365 10.4940 18.6300 ;
      RECT 10.3600 17.5365 10.3860 18.6300 ;
      RECT 10.2520 17.5365 10.2780 18.6300 ;
      RECT 10.1440 17.5365 10.1700 18.6300 ;
      RECT 10.0360 17.5365 10.0620 18.6300 ;
      RECT 9.9280 17.5365 9.9540 18.6300 ;
      RECT 9.8200 17.5365 9.8460 18.6300 ;
      RECT 9.7120 17.5365 9.7380 18.6300 ;
      RECT 9.6040 17.5365 9.6300 18.6300 ;
      RECT 9.4960 17.5365 9.5220 18.6300 ;
      RECT 9.3880 17.5365 9.4140 18.6300 ;
      RECT 9.1750 17.5365 9.2520 18.6300 ;
      RECT 7.2820 17.5365 7.3590 18.6300 ;
      RECT 7.1200 17.5365 7.1460 18.6300 ;
      RECT 7.0120 17.5365 7.0380 18.6300 ;
      RECT 6.9040 17.5365 6.9300 18.6300 ;
      RECT 6.7960 17.5365 6.8220 18.6300 ;
      RECT 6.6880 17.5365 6.7140 18.6300 ;
      RECT 6.5800 17.5365 6.6060 18.6300 ;
      RECT 6.4720 17.5365 6.4980 18.6300 ;
      RECT 6.3640 17.5365 6.3900 18.6300 ;
      RECT 6.2560 17.5365 6.2820 18.6300 ;
      RECT 6.1480 17.5365 6.1740 18.6300 ;
      RECT 6.0400 17.5365 6.0660 18.6300 ;
      RECT 5.9320 17.5365 5.9580 18.6300 ;
      RECT 5.8240 17.5365 5.8500 18.6300 ;
      RECT 5.7160 17.5365 5.7420 18.6300 ;
      RECT 5.6080 17.5365 5.6340 18.6300 ;
      RECT 5.5000 17.5365 5.5260 18.6300 ;
      RECT 5.3920 17.5365 5.4180 18.6300 ;
      RECT 5.2840 17.5365 5.3100 18.6300 ;
      RECT 5.1760 17.5365 5.2020 18.6300 ;
      RECT 5.0680 17.5365 5.0940 18.6300 ;
      RECT 4.9600 17.5365 4.9860 18.6300 ;
      RECT 4.8520 17.5365 4.8780 18.6300 ;
      RECT 4.7440 17.5365 4.7700 18.6300 ;
      RECT 4.6360 17.5365 4.6620 18.6300 ;
      RECT 4.5280 17.5365 4.5540 18.6300 ;
      RECT 4.4200 17.5365 4.4460 18.6300 ;
      RECT 4.3120 17.5365 4.3380 18.6300 ;
      RECT 4.2040 17.5365 4.2300 18.6300 ;
      RECT 4.0960 17.5365 4.1220 18.6300 ;
      RECT 3.9880 17.5365 4.0140 18.6300 ;
      RECT 3.8800 17.5365 3.9060 18.6300 ;
      RECT 3.7720 17.5365 3.7980 18.6300 ;
      RECT 3.6640 17.5365 3.6900 18.6300 ;
      RECT 3.5560 17.5365 3.5820 18.6300 ;
      RECT 3.4480 17.5365 3.4740 18.6300 ;
      RECT 3.3400 17.5365 3.3660 18.6300 ;
      RECT 3.2320 17.5365 3.2580 18.6300 ;
      RECT 3.1240 17.5365 3.1500 18.6300 ;
      RECT 3.0160 17.5365 3.0420 18.6300 ;
      RECT 2.9080 17.5365 2.9340 18.6300 ;
      RECT 2.8000 17.5365 2.8260 18.6300 ;
      RECT 2.6920 17.5365 2.7180 18.6300 ;
      RECT 2.5840 17.5365 2.6100 18.6300 ;
      RECT 2.4760 17.5365 2.5020 18.6300 ;
      RECT 2.3680 17.5365 2.3940 18.6300 ;
      RECT 2.2600 17.5365 2.2860 18.6300 ;
      RECT 2.1520 17.5365 2.1780 18.6300 ;
      RECT 2.0440 17.5365 2.0700 18.6300 ;
      RECT 1.9360 17.5365 1.9620 18.6300 ;
      RECT 1.8280 17.5365 1.8540 18.6300 ;
      RECT 1.7200 17.5365 1.7460 18.6300 ;
      RECT 1.6120 17.5365 1.6380 18.6300 ;
      RECT 1.5040 17.5365 1.5300 18.6300 ;
      RECT 1.3960 17.5365 1.4220 18.6300 ;
      RECT 1.2880 17.5365 1.3140 18.6300 ;
      RECT 1.1800 17.5365 1.2060 18.6300 ;
      RECT 1.0720 17.5365 1.0980 18.6300 ;
      RECT 0.9640 17.5365 0.9900 18.6300 ;
      RECT 0.8560 17.5365 0.8820 18.6300 ;
      RECT 0.7480 17.5365 0.7740 18.6300 ;
      RECT 0.6400 17.5365 0.6660 18.6300 ;
      RECT 0.5320 17.5365 0.5580 18.6300 ;
      RECT 0.4240 17.5365 0.4500 18.6300 ;
      RECT 0.3160 17.5365 0.3420 18.6300 ;
      RECT 0.2080 17.5365 0.2340 18.6300 ;
      RECT 0.0050 17.5365 0.0900 18.6300 ;
      RECT 8.6410 18.6165 8.7690 19.7100 ;
      RECT 8.6270 19.2820 8.7690 19.6045 ;
      RECT 8.4790 19.0090 8.5410 19.7100 ;
      RECT 8.4650 19.3185 8.5410 19.4720 ;
      RECT 8.4790 18.6165 8.5050 19.7100 ;
      RECT 8.4790 18.7375 8.5190 18.9770 ;
      RECT 8.4790 18.6165 8.5410 18.7055 ;
      RECT 8.1820 19.0670 8.3880 19.7100 ;
      RECT 8.3620 18.6165 8.3880 19.7100 ;
      RECT 8.1820 19.3440 8.4020 19.6020 ;
      RECT 8.1820 18.6165 8.2800 19.7100 ;
      RECT 7.7650 18.6165 7.8480 19.7100 ;
      RECT 7.7650 18.7050 7.8620 19.6405 ;
      RECT 16.4440 18.6165 16.5290 19.7100 ;
      RECT 16.3000 18.6165 16.3260 19.7100 ;
      RECT 16.1920 18.6165 16.2180 19.7100 ;
      RECT 16.0840 18.6165 16.1100 19.7100 ;
      RECT 15.9760 18.6165 16.0020 19.7100 ;
      RECT 15.8680 18.6165 15.8940 19.7100 ;
      RECT 15.7600 18.6165 15.7860 19.7100 ;
      RECT 15.6520 18.6165 15.6780 19.7100 ;
      RECT 15.5440 18.6165 15.5700 19.7100 ;
      RECT 15.4360 18.6165 15.4620 19.7100 ;
      RECT 15.3280 18.6165 15.3540 19.7100 ;
      RECT 15.2200 18.6165 15.2460 19.7100 ;
      RECT 15.1120 18.6165 15.1380 19.7100 ;
      RECT 15.0040 18.6165 15.0300 19.7100 ;
      RECT 14.8960 18.6165 14.9220 19.7100 ;
      RECT 14.7880 18.6165 14.8140 19.7100 ;
      RECT 14.6800 18.6165 14.7060 19.7100 ;
      RECT 14.5720 18.6165 14.5980 19.7100 ;
      RECT 14.4640 18.6165 14.4900 19.7100 ;
      RECT 14.3560 18.6165 14.3820 19.7100 ;
      RECT 14.2480 18.6165 14.2740 19.7100 ;
      RECT 14.1400 18.6165 14.1660 19.7100 ;
      RECT 14.0320 18.6165 14.0580 19.7100 ;
      RECT 13.9240 18.6165 13.9500 19.7100 ;
      RECT 13.8160 18.6165 13.8420 19.7100 ;
      RECT 13.7080 18.6165 13.7340 19.7100 ;
      RECT 13.6000 18.6165 13.6260 19.7100 ;
      RECT 13.4920 18.6165 13.5180 19.7100 ;
      RECT 13.3840 18.6165 13.4100 19.7100 ;
      RECT 13.2760 18.6165 13.3020 19.7100 ;
      RECT 13.1680 18.6165 13.1940 19.7100 ;
      RECT 13.0600 18.6165 13.0860 19.7100 ;
      RECT 12.9520 18.6165 12.9780 19.7100 ;
      RECT 12.8440 18.6165 12.8700 19.7100 ;
      RECT 12.7360 18.6165 12.7620 19.7100 ;
      RECT 12.6280 18.6165 12.6540 19.7100 ;
      RECT 12.5200 18.6165 12.5460 19.7100 ;
      RECT 12.4120 18.6165 12.4380 19.7100 ;
      RECT 12.3040 18.6165 12.3300 19.7100 ;
      RECT 12.1960 18.6165 12.2220 19.7100 ;
      RECT 12.0880 18.6165 12.1140 19.7100 ;
      RECT 11.9800 18.6165 12.0060 19.7100 ;
      RECT 11.8720 18.6165 11.8980 19.7100 ;
      RECT 11.7640 18.6165 11.7900 19.7100 ;
      RECT 11.6560 18.6165 11.6820 19.7100 ;
      RECT 11.5480 18.6165 11.5740 19.7100 ;
      RECT 11.4400 18.6165 11.4660 19.7100 ;
      RECT 11.3320 18.6165 11.3580 19.7100 ;
      RECT 11.2240 18.6165 11.2500 19.7100 ;
      RECT 11.1160 18.6165 11.1420 19.7100 ;
      RECT 11.0080 18.6165 11.0340 19.7100 ;
      RECT 10.9000 18.6165 10.9260 19.7100 ;
      RECT 10.7920 18.6165 10.8180 19.7100 ;
      RECT 10.6840 18.6165 10.7100 19.7100 ;
      RECT 10.5760 18.6165 10.6020 19.7100 ;
      RECT 10.4680 18.6165 10.4940 19.7100 ;
      RECT 10.3600 18.6165 10.3860 19.7100 ;
      RECT 10.2520 18.6165 10.2780 19.7100 ;
      RECT 10.1440 18.6165 10.1700 19.7100 ;
      RECT 10.0360 18.6165 10.0620 19.7100 ;
      RECT 9.9280 18.6165 9.9540 19.7100 ;
      RECT 9.8200 18.6165 9.8460 19.7100 ;
      RECT 9.7120 18.6165 9.7380 19.7100 ;
      RECT 9.6040 18.6165 9.6300 19.7100 ;
      RECT 9.4960 18.6165 9.5220 19.7100 ;
      RECT 9.3880 18.6165 9.4140 19.7100 ;
      RECT 9.1750 18.6165 9.2520 19.7100 ;
      RECT 7.2820 18.6165 7.3590 19.7100 ;
      RECT 7.1200 18.6165 7.1460 19.7100 ;
      RECT 7.0120 18.6165 7.0380 19.7100 ;
      RECT 6.9040 18.6165 6.9300 19.7100 ;
      RECT 6.7960 18.6165 6.8220 19.7100 ;
      RECT 6.6880 18.6165 6.7140 19.7100 ;
      RECT 6.5800 18.6165 6.6060 19.7100 ;
      RECT 6.4720 18.6165 6.4980 19.7100 ;
      RECT 6.3640 18.6165 6.3900 19.7100 ;
      RECT 6.2560 18.6165 6.2820 19.7100 ;
      RECT 6.1480 18.6165 6.1740 19.7100 ;
      RECT 6.0400 18.6165 6.0660 19.7100 ;
      RECT 5.9320 18.6165 5.9580 19.7100 ;
      RECT 5.8240 18.6165 5.8500 19.7100 ;
      RECT 5.7160 18.6165 5.7420 19.7100 ;
      RECT 5.6080 18.6165 5.6340 19.7100 ;
      RECT 5.5000 18.6165 5.5260 19.7100 ;
      RECT 5.3920 18.6165 5.4180 19.7100 ;
      RECT 5.2840 18.6165 5.3100 19.7100 ;
      RECT 5.1760 18.6165 5.2020 19.7100 ;
      RECT 5.0680 18.6165 5.0940 19.7100 ;
      RECT 4.9600 18.6165 4.9860 19.7100 ;
      RECT 4.8520 18.6165 4.8780 19.7100 ;
      RECT 4.7440 18.6165 4.7700 19.7100 ;
      RECT 4.6360 18.6165 4.6620 19.7100 ;
      RECT 4.5280 18.6165 4.5540 19.7100 ;
      RECT 4.4200 18.6165 4.4460 19.7100 ;
      RECT 4.3120 18.6165 4.3380 19.7100 ;
      RECT 4.2040 18.6165 4.2300 19.7100 ;
      RECT 4.0960 18.6165 4.1220 19.7100 ;
      RECT 3.9880 18.6165 4.0140 19.7100 ;
      RECT 3.8800 18.6165 3.9060 19.7100 ;
      RECT 3.7720 18.6165 3.7980 19.7100 ;
      RECT 3.6640 18.6165 3.6900 19.7100 ;
      RECT 3.5560 18.6165 3.5820 19.7100 ;
      RECT 3.4480 18.6165 3.4740 19.7100 ;
      RECT 3.3400 18.6165 3.3660 19.7100 ;
      RECT 3.2320 18.6165 3.2580 19.7100 ;
      RECT 3.1240 18.6165 3.1500 19.7100 ;
      RECT 3.0160 18.6165 3.0420 19.7100 ;
      RECT 2.9080 18.6165 2.9340 19.7100 ;
      RECT 2.8000 18.6165 2.8260 19.7100 ;
      RECT 2.6920 18.6165 2.7180 19.7100 ;
      RECT 2.5840 18.6165 2.6100 19.7100 ;
      RECT 2.4760 18.6165 2.5020 19.7100 ;
      RECT 2.3680 18.6165 2.3940 19.7100 ;
      RECT 2.2600 18.6165 2.2860 19.7100 ;
      RECT 2.1520 18.6165 2.1780 19.7100 ;
      RECT 2.0440 18.6165 2.0700 19.7100 ;
      RECT 1.9360 18.6165 1.9620 19.7100 ;
      RECT 1.8280 18.6165 1.8540 19.7100 ;
      RECT 1.7200 18.6165 1.7460 19.7100 ;
      RECT 1.6120 18.6165 1.6380 19.7100 ;
      RECT 1.5040 18.6165 1.5300 19.7100 ;
      RECT 1.3960 18.6165 1.4220 19.7100 ;
      RECT 1.2880 18.6165 1.3140 19.7100 ;
      RECT 1.1800 18.6165 1.2060 19.7100 ;
      RECT 1.0720 18.6165 1.0980 19.7100 ;
      RECT 0.9640 18.6165 0.9900 19.7100 ;
      RECT 0.8560 18.6165 0.8820 19.7100 ;
      RECT 0.7480 18.6165 0.7740 19.7100 ;
      RECT 0.6400 18.6165 0.6660 19.7100 ;
      RECT 0.5320 18.6165 0.5580 19.7100 ;
      RECT 0.4240 18.6165 0.4500 19.7100 ;
      RECT 0.3160 18.6165 0.3420 19.7100 ;
      RECT 0.2080 18.6165 0.2340 19.7100 ;
      RECT 0.0050 18.6165 0.0900 19.7100 ;
      RECT 8.6410 19.6965 8.7690 20.7900 ;
      RECT 8.6270 20.3620 8.7690 20.6845 ;
      RECT 8.4790 20.0890 8.5410 20.7900 ;
      RECT 8.4650 20.3985 8.5410 20.5520 ;
      RECT 8.4790 19.6965 8.5050 20.7900 ;
      RECT 8.4790 19.8175 8.5190 20.0570 ;
      RECT 8.4790 19.6965 8.5410 19.7855 ;
      RECT 8.1820 20.1470 8.3880 20.7900 ;
      RECT 8.3620 19.6965 8.3880 20.7900 ;
      RECT 8.1820 20.4240 8.4020 20.6820 ;
      RECT 8.1820 19.6965 8.2800 20.7900 ;
      RECT 7.7650 19.6965 7.8480 20.7900 ;
      RECT 7.7650 19.7850 7.8620 20.7205 ;
      RECT 16.4440 19.6965 16.5290 20.7900 ;
      RECT 16.3000 19.6965 16.3260 20.7900 ;
      RECT 16.1920 19.6965 16.2180 20.7900 ;
      RECT 16.0840 19.6965 16.1100 20.7900 ;
      RECT 15.9760 19.6965 16.0020 20.7900 ;
      RECT 15.8680 19.6965 15.8940 20.7900 ;
      RECT 15.7600 19.6965 15.7860 20.7900 ;
      RECT 15.6520 19.6965 15.6780 20.7900 ;
      RECT 15.5440 19.6965 15.5700 20.7900 ;
      RECT 15.4360 19.6965 15.4620 20.7900 ;
      RECT 15.3280 19.6965 15.3540 20.7900 ;
      RECT 15.2200 19.6965 15.2460 20.7900 ;
      RECT 15.1120 19.6965 15.1380 20.7900 ;
      RECT 15.0040 19.6965 15.0300 20.7900 ;
      RECT 14.8960 19.6965 14.9220 20.7900 ;
      RECT 14.7880 19.6965 14.8140 20.7900 ;
      RECT 14.6800 19.6965 14.7060 20.7900 ;
      RECT 14.5720 19.6965 14.5980 20.7900 ;
      RECT 14.4640 19.6965 14.4900 20.7900 ;
      RECT 14.3560 19.6965 14.3820 20.7900 ;
      RECT 14.2480 19.6965 14.2740 20.7900 ;
      RECT 14.1400 19.6965 14.1660 20.7900 ;
      RECT 14.0320 19.6965 14.0580 20.7900 ;
      RECT 13.9240 19.6965 13.9500 20.7900 ;
      RECT 13.8160 19.6965 13.8420 20.7900 ;
      RECT 13.7080 19.6965 13.7340 20.7900 ;
      RECT 13.6000 19.6965 13.6260 20.7900 ;
      RECT 13.4920 19.6965 13.5180 20.7900 ;
      RECT 13.3840 19.6965 13.4100 20.7900 ;
      RECT 13.2760 19.6965 13.3020 20.7900 ;
      RECT 13.1680 19.6965 13.1940 20.7900 ;
      RECT 13.0600 19.6965 13.0860 20.7900 ;
      RECT 12.9520 19.6965 12.9780 20.7900 ;
      RECT 12.8440 19.6965 12.8700 20.7900 ;
      RECT 12.7360 19.6965 12.7620 20.7900 ;
      RECT 12.6280 19.6965 12.6540 20.7900 ;
      RECT 12.5200 19.6965 12.5460 20.7900 ;
      RECT 12.4120 19.6965 12.4380 20.7900 ;
      RECT 12.3040 19.6965 12.3300 20.7900 ;
      RECT 12.1960 19.6965 12.2220 20.7900 ;
      RECT 12.0880 19.6965 12.1140 20.7900 ;
      RECT 11.9800 19.6965 12.0060 20.7900 ;
      RECT 11.8720 19.6965 11.8980 20.7900 ;
      RECT 11.7640 19.6965 11.7900 20.7900 ;
      RECT 11.6560 19.6965 11.6820 20.7900 ;
      RECT 11.5480 19.6965 11.5740 20.7900 ;
      RECT 11.4400 19.6965 11.4660 20.7900 ;
      RECT 11.3320 19.6965 11.3580 20.7900 ;
      RECT 11.2240 19.6965 11.2500 20.7900 ;
      RECT 11.1160 19.6965 11.1420 20.7900 ;
      RECT 11.0080 19.6965 11.0340 20.7900 ;
      RECT 10.9000 19.6965 10.9260 20.7900 ;
      RECT 10.7920 19.6965 10.8180 20.7900 ;
      RECT 10.6840 19.6965 10.7100 20.7900 ;
      RECT 10.5760 19.6965 10.6020 20.7900 ;
      RECT 10.4680 19.6965 10.4940 20.7900 ;
      RECT 10.3600 19.6965 10.3860 20.7900 ;
      RECT 10.2520 19.6965 10.2780 20.7900 ;
      RECT 10.1440 19.6965 10.1700 20.7900 ;
      RECT 10.0360 19.6965 10.0620 20.7900 ;
      RECT 9.9280 19.6965 9.9540 20.7900 ;
      RECT 9.8200 19.6965 9.8460 20.7900 ;
      RECT 9.7120 19.6965 9.7380 20.7900 ;
      RECT 9.6040 19.6965 9.6300 20.7900 ;
      RECT 9.4960 19.6965 9.5220 20.7900 ;
      RECT 9.3880 19.6965 9.4140 20.7900 ;
      RECT 9.1750 19.6965 9.2520 20.7900 ;
      RECT 7.2820 19.6965 7.3590 20.7900 ;
      RECT 7.1200 19.6965 7.1460 20.7900 ;
      RECT 7.0120 19.6965 7.0380 20.7900 ;
      RECT 6.9040 19.6965 6.9300 20.7900 ;
      RECT 6.7960 19.6965 6.8220 20.7900 ;
      RECT 6.6880 19.6965 6.7140 20.7900 ;
      RECT 6.5800 19.6965 6.6060 20.7900 ;
      RECT 6.4720 19.6965 6.4980 20.7900 ;
      RECT 6.3640 19.6965 6.3900 20.7900 ;
      RECT 6.2560 19.6965 6.2820 20.7900 ;
      RECT 6.1480 19.6965 6.1740 20.7900 ;
      RECT 6.0400 19.6965 6.0660 20.7900 ;
      RECT 5.9320 19.6965 5.9580 20.7900 ;
      RECT 5.8240 19.6965 5.8500 20.7900 ;
      RECT 5.7160 19.6965 5.7420 20.7900 ;
      RECT 5.6080 19.6965 5.6340 20.7900 ;
      RECT 5.5000 19.6965 5.5260 20.7900 ;
      RECT 5.3920 19.6965 5.4180 20.7900 ;
      RECT 5.2840 19.6965 5.3100 20.7900 ;
      RECT 5.1760 19.6965 5.2020 20.7900 ;
      RECT 5.0680 19.6965 5.0940 20.7900 ;
      RECT 4.9600 19.6965 4.9860 20.7900 ;
      RECT 4.8520 19.6965 4.8780 20.7900 ;
      RECT 4.7440 19.6965 4.7700 20.7900 ;
      RECT 4.6360 19.6965 4.6620 20.7900 ;
      RECT 4.5280 19.6965 4.5540 20.7900 ;
      RECT 4.4200 19.6965 4.4460 20.7900 ;
      RECT 4.3120 19.6965 4.3380 20.7900 ;
      RECT 4.2040 19.6965 4.2300 20.7900 ;
      RECT 4.0960 19.6965 4.1220 20.7900 ;
      RECT 3.9880 19.6965 4.0140 20.7900 ;
      RECT 3.8800 19.6965 3.9060 20.7900 ;
      RECT 3.7720 19.6965 3.7980 20.7900 ;
      RECT 3.6640 19.6965 3.6900 20.7900 ;
      RECT 3.5560 19.6965 3.5820 20.7900 ;
      RECT 3.4480 19.6965 3.4740 20.7900 ;
      RECT 3.3400 19.6965 3.3660 20.7900 ;
      RECT 3.2320 19.6965 3.2580 20.7900 ;
      RECT 3.1240 19.6965 3.1500 20.7900 ;
      RECT 3.0160 19.6965 3.0420 20.7900 ;
      RECT 2.9080 19.6965 2.9340 20.7900 ;
      RECT 2.8000 19.6965 2.8260 20.7900 ;
      RECT 2.6920 19.6965 2.7180 20.7900 ;
      RECT 2.5840 19.6965 2.6100 20.7900 ;
      RECT 2.4760 19.6965 2.5020 20.7900 ;
      RECT 2.3680 19.6965 2.3940 20.7900 ;
      RECT 2.2600 19.6965 2.2860 20.7900 ;
      RECT 2.1520 19.6965 2.1780 20.7900 ;
      RECT 2.0440 19.6965 2.0700 20.7900 ;
      RECT 1.9360 19.6965 1.9620 20.7900 ;
      RECT 1.8280 19.6965 1.8540 20.7900 ;
      RECT 1.7200 19.6965 1.7460 20.7900 ;
      RECT 1.6120 19.6965 1.6380 20.7900 ;
      RECT 1.5040 19.6965 1.5300 20.7900 ;
      RECT 1.3960 19.6965 1.4220 20.7900 ;
      RECT 1.2880 19.6965 1.3140 20.7900 ;
      RECT 1.1800 19.6965 1.2060 20.7900 ;
      RECT 1.0720 19.6965 1.0980 20.7900 ;
      RECT 0.9640 19.6965 0.9900 20.7900 ;
      RECT 0.8560 19.6965 0.8820 20.7900 ;
      RECT 0.7480 19.6965 0.7740 20.7900 ;
      RECT 0.6400 19.6965 0.6660 20.7900 ;
      RECT 0.5320 19.6965 0.5580 20.7900 ;
      RECT 0.4240 19.6965 0.4500 20.7900 ;
      RECT 0.3160 19.6965 0.3420 20.7900 ;
      RECT 0.2080 19.6965 0.2340 20.7900 ;
      RECT 0.0050 19.6965 0.0900 20.7900 ;
      RECT 8.6410 20.7765 8.7690 21.8700 ;
      RECT 8.6270 21.4420 8.7690 21.7645 ;
      RECT 8.4790 21.1690 8.5410 21.8700 ;
      RECT 8.4650 21.4785 8.5410 21.6320 ;
      RECT 8.4790 20.7765 8.5050 21.8700 ;
      RECT 8.4790 20.8975 8.5190 21.1370 ;
      RECT 8.4790 20.7765 8.5410 20.8655 ;
      RECT 8.1820 21.2270 8.3880 21.8700 ;
      RECT 8.3620 20.7765 8.3880 21.8700 ;
      RECT 8.1820 21.5040 8.4020 21.7620 ;
      RECT 8.1820 20.7765 8.2800 21.8700 ;
      RECT 7.7650 20.7765 7.8480 21.8700 ;
      RECT 7.7650 20.8650 7.8620 21.8005 ;
      RECT 16.4440 20.7765 16.5290 21.8700 ;
      RECT 16.3000 20.7765 16.3260 21.8700 ;
      RECT 16.1920 20.7765 16.2180 21.8700 ;
      RECT 16.0840 20.7765 16.1100 21.8700 ;
      RECT 15.9760 20.7765 16.0020 21.8700 ;
      RECT 15.8680 20.7765 15.8940 21.8700 ;
      RECT 15.7600 20.7765 15.7860 21.8700 ;
      RECT 15.6520 20.7765 15.6780 21.8700 ;
      RECT 15.5440 20.7765 15.5700 21.8700 ;
      RECT 15.4360 20.7765 15.4620 21.8700 ;
      RECT 15.3280 20.7765 15.3540 21.8700 ;
      RECT 15.2200 20.7765 15.2460 21.8700 ;
      RECT 15.1120 20.7765 15.1380 21.8700 ;
      RECT 15.0040 20.7765 15.0300 21.8700 ;
      RECT 14.8960 20.7765 14.9220 21.8700 ;
      RECT 14.7880 20.7765 14.8140 21.8700 ;
      RECT 14.6800 20.7765 14.7060 21.8700 ;
      RECT 14.5720 20.7765 14.5980 21.8700 ;
      RECT 14.4640 20.7765 14.4900 21.8700 ;
      RECT 14.3560 20.7765 14.3820 21.8700 ;
      RECT 14.2480 20.7765 14.2740 21.8700 ;
      RECT 14.1400 20.7765 14.1660 21.8700 ;
      RECT 14.0320 20.7765 14.0580 21.8700 ;
      RECT 13.9240 20.7765 13.9500 21.8700 ;
      RECT 13.8160 20.7765 13.8420 21.8700 ;
      RECT 13.7080 20.7765 13.7340 21.8700 ;
      RECT 13.6000 20.7765 13.6260 21.8700 ;
      RECT 13.4920 20.7765 13.5180 21.8700 ;
      RECT 13.3840 20.7765 13.4100 21.8700 ;
      RECT 13.2760 20.7765 13.3020 21.8700 ;
      RECT 13.1680 20.7765 13.1940 21.8700 ;
      RECT 13.0600 20.7765 13.0860 21.8700 ;
      RECT 12.9520 20.7765 12.9780 21.8700 ;
      RECT 12.8440 20.7765 12.8700 21.8700 ;
      RECT 12.7360 20.7765 12.7620 21.8700 ;
      RECT 12.6280 20.7765 12.6540 21.8700 ;
      RECT 12.5200 20.7765 12.5460 21.8700 ;
      RECT 12.4120 20.7765 12.4380 21.8700 ;
      RECT 12.3040 20.7765 12.3300 21.8700 ;
      RECT 12.1960 20.7765 12.2220 21.8700 ;
      RECT 12.0880 20.7765 12.1140 21.8700 ;
      RECT 11.9800 20.7765 12.0060 21.8700 ;
      RECT 11.8720 20.7765 11.8980 21.8700 ;
      RECT 11.7640 20.7765 11.7900 21.8700 ;
      RECT 11.6560 20.7765 11.6820 21.8700 ;
      RECT 11.5480 20.7765 11.5740 21.8700 ;
      RECT 11.4400 20.7765 11.4660 21.8700 ;
      RECT 11.3320 20.7765 11.3580 21.8700 ;
      RECT 11.2240 20.7765 11.2500 21.8700 ;
      RECT 11.1160 20.7765 11.1420 21.8700 ;
      RECT 11.0080 20.7765 11.0340 21.8700 ;
      RECT 10.9000 20.7765 10.9260 21.8700 ;
      RECT 10.7920 20.7765 10.8180 21.8700 ;
      RECT 10.6840 20.7765 10.7100 21.8700 ;
      RECT 10.5760 20.7765 10.6020 21.8700 ;
      RECT 10.4680 20.7765 10.4940 21.8700 ;
      RECT 10.3600 20.7765 10.3860 21.8700 ;
      RECT 10.2520 20.7765 10.2780 21.8700 ;
      RECT 10.1440 20.7765 10.1700 21.8700 ;
      RECT 10.0360 20.7765 10.0620 21.8700 ;
      RECT 9.9280 20.7765 9.9540 21.8700 ;
      RECT 9.8200 20.7765 9.8460 21.8700 ;
      RECT 9.7120 20.7765 9.7380 21.8700 ;
      RECT 9.6040 20.7765 9.6300 21.8700 ;
      RECT 9.4960 20.7765 9.5220 21.8700 ;
      RECT 9.3880 20.7765 9.4140 21.8700 ;
      RECT 9.1750 20.7765 9.2520 21.8700 ;
      RECT 7.2820 20.7765 7.3590 21.8700 ;
      RECT 7.1200 20.7765 7.1460 21.8700 ;
      RECT 7.0120 20.7765 7.0380 21.8700 ;
      RECT 6.9040 20.7765 6.9300 21.8700 ;
      RECT 6.7960 20.7765 6.8220 21.8700 ;
      RECT 6.6880 20.7765 6.7140 21.8700 ;
      RECT 6.5800 20.7765 6.6060 21.8700 ;
      RECT 6.4720 20.7765 6.4980 21.8700 ;
      RECT 6.3640 20.7765 6.3900 21.8700 ;
      RECT 6.2560 20.7765 6.2820 21.8700 ;
      RECT 6.1480 20.7765 6.1740 21.8700 ;
      RECT 6.0400 20.7765 6.0660 21.8700 ;
      RECT 5.9320 20.7765 5.9580 21.8700 ;
      RECT 5.8240 20.7765 5.8500 21.8700 ;
      RECT 5.7160 20.7765 5.7420 21.8700 ;
      RECT 5.6080 20.7765 5.6340 21.8700 ;
      RECT 5.5000 20.7765 5.5260 21.8700 ;
      RECT 5.3920 20.7765 5.4180 21.8700 ;
      RECT 5.2840 20.7765 5.3100 21.8700 ;
      RECT 5.1760 20.7765 5.2020 21.8700 ;
      RECT 5.0680 20.7765 5.0940 21.8700 ;
      RECT 4.9600 20.7765 4.9860 21.8700 ;
      RECT 4.8520 20.7765 4.8780 21.8700 ;
      RECT 4.7440 20.7765 4.7700 21.8700 ;
      RECT 4.6360 20.7765 4.6620 21.8700 ;
      RECT 4.5280 20.7765 4.5540 21.8700 ;
      RECT 4.4200 20.7765 4.4460 21.8700 ;
      RECT 4.3120 20.7765 4.3380 21.8700 ;
      RECT 4.2040 20.7765 4.2300 21.8700 ;
      RECT 4.0960 20.7765 4.1220 21.8700 ;
      RECT 3.9880 20.7765 4.0140 21.8700 ;
      RECT 3.8800 20.7765 3.9060 21.8700 ;
      RECT 3.7720 20.7765 3.7980 21.8700 ;
      RECT 3.6640 20.7765 3.6900 21.8700 ;
      RECT 3.5560 20.7765 3.5820 21.8700 ;
      RECT 3.4480 20.7765 3.4740 21.8700 ;
      RECT 3.3400 20.7765 3.3660 21.8700 ;
      RECT 3.2320 20.7765 3.2580 21.8700 ;
      RECT 3.1240 20.7765 3.1500 21.8700 ;
      RECT 3.0160 20.7765 3.0420 21.8700 ;
      RECT 2.9080 20.7765 2.9340 21.8700 ;
      RECT 2.8000 20.7765 2.8260 21.8700 ;
      RECT 2.6920 20.7765 2.7180 21.8700 ;
      RECT 2.5840 20.7765 2.6100 21.8700 ;
      RECT 2.4760 20.7765 2.5020 21.8700 ;
      RECT 2.3680 20.7765 2.3940 21.8700 ;
      RECT 2.2600 20.7765 2.2860 21.8700 ;
      RECT 2.1520 20.7765 2.1780 21.8700 ;
      RECT 2.0440 20.7765 2.0700 21.8700 ;
      RECT 1.9360 20.7765 1.9620 21.8700 ;
      RECT 1.8280 20.7765 1.8540 21.8700 ;
      RECT 1.7200 20.7765 1.7460 21.8700 ;
      RECT 1.6120 20.7765 1.6380 21.8700 ;
      RECT 1.5040 20.7765 1.5300 21.8700 ;
      RECT 1.3960 20.7765 1.4220 21.8700 ;
      RECT 1.2880 20.7765 1.3140 21.8700 ;
      RECT 1.1800 20.7765 1.2060 21.8700 ;
      RECT 1.0720 20.7765 1.0980 21.8700 ;
      RECT 0.9640 20.7765 0.9900 21.8700 ;
      RECT 0.8560 20.7765 0.8820 21.8700 ;
      RECT 0.7480 20.7765 0.7740 21.8700 ;
      RECT 0.6400 20.7765 0.6660 21.8700 ;
      RECT 0.5320 20.7765 0.5580 21.8700 ;
      RECT 0.4240 20.7765 0.4500 21.8700 ;
      RECT 0.3160 20.7765 0.3420 21.8700 ;
      RECT 0.2080 20.7765 0.2340 21.8700 ;
      RECT 0.0050 20.7765 0.0900 21.8700 ;
      RECT 8.6410 21.8565 8.7690 22.9500 ;
      RECT 8.6270 22.5220 8.7690 22.8445 ;
      RECT 8.4790 22.2490 8.5410 22.9500 ;
      RECT 8.4650 22.5585 8.5410 22.7120 ;
      RECT 8.4790 21.8565 8.5050 22.9500 ;
      RECT 8.4790 21.9775 8.5190 22.2170 ;
      RECT 8.4790 21.8565 8.5410 21.9455 ;
      RECT 8.1820 22.3070 8.3880 22.9500 ;
      RECT 8.3620 21.8565 8.3880 22.9500 ;
      RECT 8.1820 22.5840 8.4020 22.8420 ;
      RECT 8.1820 21.8565 8.2800 22.9500 ;
      RECT 7.7650 21.8565 7.8480 22.9500 ;
      RECT 7.7650 21.9450 7.8620 22.8805 ;
      RECT 16.4440 21.8565 16.5290 22.9500 ;
      RECT 16.3000 21.8565 16.3260 22.9500 ;
      RECT 16.1920 21.8565 16.2180 22.9500 ;
      RECT 16.0840 21.8565 16.1100 22.9500 ;
      RECT 15.9760 21.8565 16.0020 22.9500 ;
      RECT 15.8680 21.8565 15.8940 22.9500 ;
      RECT 15.7600 21.8565 15.7860 22.9500 ;
      RECT 15.6520 21.8565 15.6780 22.9500 ;
      RECT 15.5440 21.8565 15.5700 22.9500 ;
      RECT 15.4360 21.8565 15.4620 22.9500 ;
      RECT 15.3280 21.8565 15.3540 22.9500 ;
      RECT 15.2200 21.8565 15.2460 22.9500 ;
      RECT 15.1120 21.8565 15.1380 22.9500 ;
      RECT 15.0040 21.8565 15.0300 22.9500 ;
      RECT 14.8960 21.8565 14.9220 22.9500 ;
      RECT 14.7880 21.8565 14.8140 22.9500 ;
      RECT 14.6800 21.8565 14.7060 22.9500 ;
      RECT 14.5720 21.8565 14.5980 22.9500 ;
      RECT 14.4640 21.8565 14.4900 22.9500 ;
      RECT 14.3560 21.8565 14.3820 22.9500 ;
      RECT 14.2480 21.8565 14.2740 22.9500 ;
      RECT 14.1400 21.8565 14.1660 22.9500 ;
      RECT 14.0320 21.8565 14.0580 22.9500 ;
      RECT 13.9240 21.8565 13.9500 22.9500 ;
      RECT 13.8160 21.8565 13.8420 22.9500 ;
      RECT 13.7080 21.8565 13.7340 22.9500 ;
      RECT 13.6000 21.8565 13.6260 22.9500 ;
      RECT 13.4920 21.8565 13.5180 22.9500 ;
      RECT 13.3840 21.8565 13.4100 22.9500 ;
      RECT 13.2760 21.8565 13.3020 22.9500 ;
      RECT 13.1680 21.8565 13.1940 22.9500 ;
      RECT 13.0600 21.8565 13.0860 22.9500 ;
      RECT 12.9520 21.8565 12.9780 22.9500 ;
      RECT 12.8440 21.8565 12.8700 22.9500 ;
      RECT 12.7360 21.8565 12.7620 22.9500 ;
      RECT 12.6280 21.8565 12.6540 22.9500 ;
      RECT 12.5200 21.8565 12.5460 22.9500 ;
      RECT 12.4120 21.8565 12.4380 22.9500 ;
      RECT 12.3040 21.8565 12.3300 22.9500 ;
      RECT 12.1960 21.8565 12.2220 22.9500 ;
      RECT 12.0880 21.8565 12.1140 22.9500 ;
      RECT 11.9800 21.8565 12.0060 22.9500 ;
      RECT 11.8720 21.8565 11.8980 22.9500 ;
      RECT 11.7640 21.8565 11.7900 22.9500 ;
      RECT 11.6560 21.8565 11.6820 22.9500 ;
      RECT 11.5480 21.8565 11.5740 22.9500 ;
      RECT 11.4400 21.8565 11.4660 22.9500 ;
      RECT 11.3320 21.8565 11.3580 22.9500 ;
      RECT 11.2240 21.8565 11.2500 22.9500 ;
      RECT 11.1160 21.8565 11.1420 22.9500 ;
      RECT 11.0080 21.8565 11.0340 22.9500 ;
      RECT 10.9000 21.8565 10.9260 22.9500 ;
      RECT 10.7920 21.8565 10.8180 22.9500 ;
      RECT 10.6840 21.8565 10.7100 22.9500 ;
      RECT 10.5760 21.8565 10.6020 22.9500 ;
      RECT 10.4680 21.8565 10.4940 22.9500 ;
      RECT 10.3600 21.8565 10.3860 22.9500 ;
      RECT 10.2520 21.8565 10.2780 22.9500 ;
      RECT 10.1440 21.8565 10.1700 22.9500 ;
      RECT 10.0360 21.8565 10.0620 22.9500 ;
      RECT 9.9280 21.8565 9.9540 22.9500 ;
      RECT 9.8200 21.8565 9.8460 22.9500 ;
      RECT 9.7120 21.8565 9.7380 22.9500 ;
      RECT 9.6040 21.8565 9.6300 22.9500 ;
      RECT 9.4960 21.8565 9.5220 22.9500 ;
      RECT 9.3880 21.8565 9.4140 22.9500 ;
      RECT 9.1750 21.8565 9.2520 22.9500 ;
      RECT 7.2820 21.8565 7.3590 22.9500 ;
      RECT 7.1200 21.8565 7.1460 22.9500 ;
      RECT 7.0120 21.8565 7.0380 22.9500 ;
      RECT 6.9040 21.8565 6.9300 22.9500 ;
      RECT 6.7960 21.8565 6.8220 22.9500 ;
      RECT 6.6880 21.8565 6.7140 22.9500 ;
      RECT 6.5800 21.8565 6.6060 22.9500 ;
      RECT 6.4720 21.8565 6.4980 22.9500 ;
      RECT 6.3640 21.8565 6.3900 22.9500 ;
      RECT 6.2560 21.8565 6.2820 22.9500 ;
      RECT 6.1480 21.8565 6.1740 22.9500 ;
      RECT 6.0400 21.8565 6.0660 22.9500 ;
      RECT 5.9320 21.8565 5.9580 22.9500 ;
      RECT 5.8240 21.8565 5.8500 22.9500 ;
      RECT 5.7160 21.8565 5.7420 22.9500 ;
      RECT 5.6080 21.8565 5.6340 22.9500 ;
      RECT 5.5000 21.8565 5.5260 22.9500 ;
      RECT 5.3920 21.8565 5.4180 22.9500 ;
      RECT 5.2840 21.8565 5.3100 22.9500 ;
      RECT 5.1760 21.8565 5.2020 22.9500 ;
      RECT 5.0680 21.8565 5.0940 22.9500 ;
      RECT 4.9600 21.8565 4.9860 22.9500 ;
      RECT 4.8520 21.8565 4.8780 22.9500 ;
      RECT 4.7440 21.8565 4.7700 22.9500 ;
      RECT 4.6360 21.8565 4.6620 22.9500 ;
      RECT 4.5280 21.8565 4.5540 22.9500 ;
      RECT 4.4200 21.8565 4.4460 22.9500 ;
      RECT 4.3120 21.8565 4.3380 22.9500 ;
      RECT 4.2040 21.8565 4.2300 22.9500 ;
      RECT 4.0960 21.8565 4.1220 22.9500 ;
      RECT 3.9880 21.8565 4.0140 22.9500 ;
      RECT 3.8800 21.8565 3.9060 22.9500 ;
      RECT 3.7720 21.8565 3.7980 22.9500 ;
      RECT 3.6640 21.8565 3.6900 22.9500 ;
      RECT 3.5560 21.8565 3.5820 22.9500 ;
      RECT 3.4480 21.8565 3.4740 22.9500 ;
      RECT 3.3400 21.8565 3.3660 22.9500 ;
      RECT 3.2320 21.8565 3.2580 22.9500 ;
      RECT 3.1240 21.8565 3.1500 22.9500 ;
      RECT 3.0160 21.8565 3.0420 22.9500 ;
      RECT 2.9080 21.8565 2.9340 22.9500 ;
      RECT 2.8000 21.8565 2.8260 22.9500 ;
      RECT 2.6920 21.8565 2.7180 22.9500 ;
      RECT 2.5840 21.8565 2.6100 22.9500 ;
      RECT 2.4760 21.8565 2.5020 22.9500 ;
      RECT 2.3680 21.8565 2.3940 22.9500 ;
      RECT 2.2600 21.8565 2.2860 22.9500 ;
      RECT 2.1520 21.8565 2.1780 22.9500 ;
      RECT 2.0440 21.8565 2.0700 22.9500 ;
      RECT 1.9360 21.8565 1.9620 22.9500 ;
      RECT 1.8280 21.8565 1.8540 22.9500 ;
      RECT 1.7200 21.8565 1.7460 22.9500 ;
      RECT 1.6120 21.8565 1.6380 22.9500 ;
      RECT 1.5040 21.8565 1.5300 22.9500 ;
      RECT 1.3960 21.8565 1.4220 22.9500 ;
      RECT 1.2880 21.8565 1.3140 22.9500 ;
      RECT 1.1800 21.8565 1.2060 22.9500 ;
      RECT 1.0720 21.8565 1.0980 22.9500 ;
      RECT 0.9640 21.8565 0.9900 22.9500 ;
      RECT 0.8560 21.8565 0.8820 22.9500 ;
      RECT 0.7480 21.8565 0.7740 22.9500 ;
      RECT 0.6400 21.8565 0.6660 22.9500 ;
      RECT 0.5320 21.8565 0.5580 22.9500 ;
      RECT 0.4240 21.8565 0.4500 22.9500 ;
      RECT 0.3160 21.8565 0.3420 22.9500 ;
      RECT 0.2080 21.8565 0.2340 22.9500 ;
      RECT 0.0050 21.8565 0.0900 22.9500 ;
      RECT 8.6410 22.9365 8.7690 24.0300 ;
      RECT 8.6270 23.6020 8.7690 23.9245 ;
      RECT 8.4790 23.3290 8.5410 24.0300 ;
      RECT 8.4650 23.6385 8.5410 23.7920 ;
      RECT 8.4790 22.9365 8.5050 24.0300 ;
      RECT 8.4790 23.0575 8.5190 23.2970 ;
      RECT 8.4790 22.9365 8.5410 23.0255 ;
      RECT 8.1820 23.3870 8.3880 24.0300 ;
      RECT 8.3620 22.9365 8.3880 24.0300 ;
      RECT 8.1820 23.6640 8.4020 23.9220 ;
      RECT 8.1820 22.9365 8.2800 24.0300 ;
      RECT 7.7650 22.9365 7.8480 24.0300 ;
      RECT 7.7650 23.0250 7.8620 23.9605 ;
      RECT 16.4440 22.9365 16.5290 24.0300 ;
      RECT 16.3000 22.9365 16.3260 24.0300 ;
      RECT 16.1920 22.9365 16.2180 24.0300 ;
      RECT 16.0840 22.9365 16.1100 24.0300 ;
      RECT 15.9760 22.9365 16.0020 24.0300 ;
      RECT 15.8680 22.9365 15.8940 24.0300 ;
      RECT 15.7600 22.9365 15.7860 24.0300 ;
      RECT 15.6520 22.9365 15.6780 24.0300 ;
      RECT 15.5440 22.9365 15.5700 24.0300 ;
      RECT 15.4360 22.9365 15.4620 24.0300 ;
      RECT 15.3280 22.9365 15.3540 24.0300 ;
      RECT 15.2200 22.9365 15.2460 24.0300 ;
      RECT 15.1120 22.9365 15.1380 24.0300 ;
      RECT 15.0040 22.9365 15.0300 24.0300 ;
      RECT 14.8960 22.9365 14.9220 24.0300 ;
      RECT 14.7880 22.9365 14.8140 24.0300 ;
      RECT 14.6800 22.9365 14.7060 24.0300 ;
      RECT 14.5720 22.9365 14.5980 24.0300 ;
      RECT 14.4640 22.9365 14.4900 24.0300 ;
      RECT 14.3560 22.9365 14.3820 24.0300 ;
      RECT 14.2480 22.9365 14.2740 24.0300 ;
      RECT 14.1400 22.9365 14.1660 24.0300 ;
      RECT 14.0320 22.9365 14.0580 24.0300 ;
      RECT 13.9240 22.9365 13.9500 24.0300 ;
      RECT 13.8160 22.9365 13.8420 24.0300 ;
      RECT 13.7080 22.9365 13.7340 24.0300 ;
      RECT 13.6000 22.9365 13.6260 24.0300 ;
      RECT 13.4920 22.9365 13.5180 24.0300 ;
      RECT 13.3840 22.9365 13.4100 24.0300 ;
      RECT 13.2760 22.9365 13.3020 24.0300 ;
      RECT 13.1680 22.9365 13.1940 24.0300 ;
      RECT 13.0600 22.9365 13.0860 24.0300 ;
      RECT 12.9520 22.9365 12.9780 24.0300 ;
      RECT 12.8440 22.9365 12.8700 24.0300 ;
      RECT 12.7360 22.9365 12.7620 24.0300 ;
      RECT 12.6280 22.9365 12.6540 24.0300 ;
      RECT 12.5200 22.9365 12.5460 24.0300 ;
      RECT 12.4120 22.9365 12.4380 24.0300 ;
      RECT 12.3040 22.9365 12.3300 24.0300 ;
      RECT 12.1960 22.9365 12.2220 24.0300 ;
      RECT 12.0880 22.9365 12.1140 24.0300 ;
      RECT 11.9800 22.9365 12.0060 24.0300 ;
      RECT 11.8720 22.9365 11.8980 24.0300 ;
      RECT 11.7640 22.9365 11.7900 24.0300 ;
      RECT 11.6560 22.9365 11.6820 24.0300 ;
      RECT 11.5480 22.9365 11.5740 24.0300 ;
      RECT 11.4400 22.9365 11.4660 24.0300 ;
      RECT 11.3320 22.9365 11.3580 24.0300 ;
      RECT 11.2240 22.9365 11.2500 24.0300 ;
      RECT 11.1160 22.9365 11.1420 24.0300 ;
      RECT 11.0080 22.9365 11.0340 24.0300 ;
      RECT 10.9000 22.9365 10.9260 24.0300 ;
      RECT 10.7920 22.9365 10.8180 24.0300 ;
      RECT 10.6840 22.9365 10.7100 24.0300 ;
      RECT 10.5760 22.9365 10.6020 24.0300 ;
      RECT 10.4680 22.9365 10.4940 24.0300 ;
      RECT 10.3600 22.9365 10.3860 24.0300 ;
      RECT 10.2520 22.9365 10.2780 24.0300 ;
      RECT 10.1440 22.9365 10.1700 24.0300 ;
      RECT 10.0360 22.9365 10.0620 24.0300 ;
      RECT 9.9280 22.9365 9.9540 24.0300 ;
      RECT 9.8200 22.9365 9.8460 24.0300 ;
      RECT 9.7120 22.9365 9.7380 24.0300 ;
      RECT 9.6040 22.9365 9.6300 24.0300 ;
      RECT 9.4960 22.9365 9.5220 24.0300 ;
      RECT 9.3880 22.9365 9.4140 24.0300 ;
      RECT 9.1750 22.9365 9.2520 24.0300 ;
      RECT 7.2820 22.9365 7.3590 24.0300 ;
      RECT 7.1200 22.9365 7.1460 24.0300 ;
      RECT 7.0120 22.9365 7.0380 24.0300 ;
      RECT 6.9040 22.9365 6.9300 24.0300 ;
      RECT 6.7960 22.9365 6.8220 24.0300 ;
      RECT 6.6880 22.9365 6.7140 24.0300 ;
      RECT 6.5800 22.9365 6.6060 24.0300 ;
      RECT 6.4720 22.9365 6.4980 24.0300 ;
      RECT 6.3640 22.9365 6.3900 24.0300 ;
      RECT 6.2560 22.9365 6.2820 24.0300 ;
      RECT 6.1480 22.9365 6.1740 24.0300 ;
      RECT 6.0400 22.9365 6.0660 24.0300 ;
      RECT 5.9320 22.9365 5.9580 24.0300 ;
      RECT 5.8240 22.9365 5.8500 24.0300 ;
      RECT 5.7160 22.9365 5.7420 24.0300 ;
      RECT 5.6080 22.9365 5.6340 24.0300 ;
      RECT 5.5000 22.9365 5.5260 24.0300 ;
      RECT 5.3920 22.9365 5.4180 24.0300 ;
      RECT 5.2840 22.9365 5.3100 24.0300 ;
      RECT 5.1760 22.9365 5.2020 24.0300 ;
      RECT 5.0680 22.9365 5.0940 24.0300 ;
      RECT 4.9600 22.9365 4.9860 24.0300 ;
      RECT 4.8520 22.9365 4.8780 24.0300 ;
      RECT 4.7440 22.9365 4.7700 24.0300 ;
      RECT 4.6360 22.9365 4.6620 24.0300 ;
      RECT 4.5280 22.9365 4.5540 24.0300 ;
      RECT 4.4200 22.9365 4.4460 24.0300 ;
      RECT 4.3120 22.9365 4.3380 24.0300 ;
      RECT 4.2040 22.9365 4.2300 24.0300 ;
      RECT 4.0960 22.9365 4.1220 24.0300 ;
      RECT 3.9880 22.9365 4.0140 24.0300 ;
      RECT 3.8800 22.9365 3.9060 24.0300 ;
      RECT 3.7720 22.9365 3.7980 24.0300 ;
      RECT 3.6640 22.9365 3.6900 24.0300 ;
      RECT 3.5560 22.9365 3.5820 24.0300 ;
      RECT 3.4480 22.9365 3.4740 24.0300 ;
      RECT 3.3400 22.9365 3.3660 24.0300 ;
      RECT 3.2320 22.9365 3.2580 24.0300 ;
      RECT 3.1240 22.9365 3.1500 24.0300 ;
      RECT 3.0160 22.9365 3.0420 24.0300 ;
      RECT 2.9080 22.9365 2.9340 24.0300 ;
      RECT 2.8000 22.9365 2.8260 24.0300 ;
      RECT 2.6920 22.9365 2.7180 24.0300 ;
      RECT 2.5840 22.9365 2.6100 24.0300 ;
      RECT 2.4760 22.9365 2.5020 24.0300 ;
      RECT 2.3680 22.9365 2.3940 24.0300 ;
      RECT 2.2600 22.9365 2.2860 24.0300 ;
      RECT 2.1520 22.9365 2.1780 24.0300 ;
      RECT 2.0440 22.9365 2.0700 24.0300 ;
      RECT 1.9360 22.9365 1.9620 24.0300 ;
      RECT 1.8280 22.9365 1.8540 24.0300 ;
      RECT 1.7200 22.9365 1.7460 24.0300 ;
      RECT 1.6120 22.9365 1.6380 24.0300 ;
      RECT 1.5040 22.9365 1.5300 24.0300 ;
      RECT 1.3960 22.9365 1.4220 24.0300 ;
      RECT 1.2880 22.9365 1.3140 24.0300 ;
      RECT 1.1800 22.9365 1.2060 24.0300 ;
      RECT 1.0720 22.9365 1.0980 24.0300 ;
      RECT 0.9640 22.9365 0.9900 24.0300 ;
      RECT 0.8560 22.9365 0.8820 24.0300 ;
      RECT 0.7480 22.9365 0.7740 24.0300 ;
      RECT 0.6400 22.9365 0.6660 24.0300 ;
      RECT 0.5320 22.9365 0.5580 24.0300 ;
      RECT 0.4240 22.9365 0.4500 24.0300 ;
      RECT 0.3160 22.9365 0.3420 24.0300 ;
      RECT 0.2080 22.9365 0.2340 24.0300 ;
      RECT 0.0050 22.9365 0.0900 24.0300 ;
      RECT 8.6410 24.0165 8.7690 25.1100 ;
      RECT 8.6270 24.6820 8.7690 25.0045 ;
      RECT 8.4790 24.4090 8.5410 25.1100 ;
      RECT 8.4650 24.7185 8.5410 24.8720 ;
      RECT 8.4790 24.0165 8.5050 25.1100 ;
      RECT 8.4790 24.1375 8.5190 24.3770 ;
      RECT 8.4790 24.0165 8.5410 24.1055 ;
      RECT 8.1820 24.4670 8.3880 25.1100 ;
      RECT 8.3620 24.0165 8.3880 25.1100 ;
      RECT 8.1820 24.7440 8.4020 25.0020 ;
      RECT 8.1820 24.0165 8.2800 25.1100 ;
      RECT 7.7650 24.0165 7.8480 25.1100 ;
      RECT 7.7650 24.1050 7.8620 25.0405 ;
      RECT 16.4440 24.0165 16.5290 25.1100 ;
      RECT 16.3000 24.0165 16.3260 25.1100 ;
      RECT 16.1920 24.0165 16.2180 25.1100 ;
      RECT 16.0840 24.0165 16.1100 25.1100 ;
      RECT 15.9760 24.0165 16.0020 25.1100 ;
      RECT 15.8680 24.0165 15.8940 25.1100 ;
      RECT 15.7600 24.0165 15.7860 25.1100 ;
      RECT 15.6520 24.0165 15.6780 25.1100 ;
      RECT 15.5440 24.0165 15.5700 25.1100 ;
      RECT 15.4360 24.0165 15.4620 25.1100 ;
      RECT 15.3280 24.0165 15.3540 25.1100 ;
      RECT 15.2200 24.0165 15.2460 25.1100 ;
      RECT 15.1120 24.0165 15.1380 25.1100 ;
      RECT 15.0040 24.0165 15.0300 25.1100 ;
      RECT 14.8960 24.0165 14.9220 25.1100 ;
      RECT 14.7880 24.0165 14.8140 25.1100 ;
      RECT 14.6800 24.0165 14.7060 25.1100 ;
      RECT 14.5720 24.0165 14.5980 25.1100 ;
      RECT 14.4640 24.0165 14.4900 25.1100 ;
      RECT 14.3560 24.0165 14.3820 25.1100 ;
      RECT 14.2480 24.0165 14.2740 25.1100 ;
      RECT 14.1400 24.0165 14.1660 25.1100 ;
      RECT 14.0320 24.0165 14.0580 25.1100 ;
      RECT 13.9240 24.0165 13.9500 25.1100 ;
      RECT 13.8160 24.0165 13.8420 25.1100 ;
      RECT 13.7080 24.0165 13.7340 25.1100 ;
      RECT 13.6000 24.0165 13.6260 25.1100 ;
      RECT 13.4920 24.0165 13.5180 25.1100 ;
      RECT 13.3840 24.0165 13.4100 25.1100 ;
      RECT 13.2760 24.0165 13.3020 25.1100 ;
      RECT 13.1680 24.0165 13.1940 25.1100 ;
      RECT 13.0600 24.0165 13.0860 25.1100 ;
      RECT 12.9520 24.0165 12.9780 25.1100 ;
      RECT 12.8440 24.0165 12.8700 25.1100 ;
      RECT 12.7360 24.0165 12.7620 25.1100 ;
      RECT 12.6280 24.0165 12.6540 25.1100 ;
      RECT 12.5200 24.0165 12.5460 25.1100 ;
      RECT 12.4120 24.0165 12.4380 25.1100 ;
      RECT 12.3040 24.0165 12.3300 25.1100 ;
      RECT 12.1960 24.0165 12.2220 25.1100 ;
      RECT 12.0880 24.0165 12.1140 25.1100 ;
      RECT 11.9800 24.0165 12.0060 25.1100 ;
      RECT 11.8720 24.0165 11.8980 25.1100 ;
      RECT 11.7640 24.0165 11.7900 25.1100 ;
      RECT 11.6560 24.0165 11.6820 25.1100 ;
      RECT 11.5480 24.0165 11.5740 25.1100 ;
      RECT 11.4400 24.0165 11.4660 25.1100 ;
      RECT 11.3320 24.0165 11.3580 25.1100 ;
      RECT 11.2240 24.0165 11.2500 25.1100 ;
      RECT 11.1160 24.0165 11.1420 25.1100 ;
      RECT 11.0080 24.0165 11.0340 25.1100 ;
      RECT 10.9000 24.0165 10.9260 25.1100 ;
      RECT 10.7920 24.0165 10.8180 25.1100 ;
      RECT 10.6840 24.0165 10.7100 25.1100 ;
      RECT 10.5760 24.0165 10.6020 25.1100 ;
      RECT 10.4680 24.0165 10.4940 25.1100 ;
      RECT 10.3600 24.0165 10.3860 25.1100 ;
      RECT 10.2520 24.0165 10.2780 25.1100 ;
      RECT 10.1440 24.0165 10.1700 25.1100 ;
      RECT 10.0360 24.0165 10.0620 25.1100 ;
      RECT 9.9280 24.0165 9.9540 25.1100 ;
      RECT 9.8200 24.0165 9.8460 25.1100 ;
      RECT 9.7120 24.0165 9.7380 25.1100 ;
      RECT 9.6040 24.0165 9.6300 25.1100 ;
      RECT 9.4960 24.0165 9.5220 25.1100 ;
      RECT 9.3880 24.0165 9.4140 25.1100 ;
      RECT 9.1750 24.0165 9.2520 25.1100 ;
      RECT 7.2820 24.0165 7.3590 25.1100 ;
      RECT 7.1200 24.0165 7.1460 25.1100 ;
      RECT 7.0120 24.0165 7.0380 25.1100 ;
      RECT 6.9040 24.0165 6.9300 25.1100 ;
      RECT 6.7960 24.0165 6.8220 25.1100 ;
      RECT 6.6880 24.0165 6.7140 25.1100 ;
      RECT 6.5800 24.0165 6.6060 25.1100 ;
      RECT 6.4720 24.0165 6.4980 25.1100 ;
      RECT 6.3640 24.0165 6.3900 25.1100 ;
      RECT 6.2560 24.0165 6.2820 25.1100 ;
      RECT 6.1480 24.0165 6.1740 25.1100 ;
      RECT 6.0400 24.0165 6.0660 25.1100 ;
      RECT 5.9320 24.0165 5.9580 25.1100 ;
      RECT 5.8240 24.0165 5.8500 25.1100 ;
      RECT 5.7160 24.0165 5.7420 25.1100 ;
      RECT 5.6080 24.0165 5.6340 25.1100 ;
      RECT 5.5000 24.0165 5.5260 25.1100 ;
      RECT 5.3920 24.0165 5.4180 25.1100 ;
      RECT 5.2840 24.0165 5.3100 25.1100 ;
      RECT 5.1760 24.0165 5.2020 25.1100 ;
      RECT 5.0680 24.0165 5.0940 25.1100 ;
      RECT 4.9600 24.0165 4.9860 25.1100 ;
      RECT 4.8520 24.0165 4.8780 25.1100 ;
      RECT 4.7440 24.0165 4.7700 25.1100 ;
      RECT 4.6360 24.0165 4.6620 25.1100 ;
      RECT 4.5280 24.0165 4.5540 25.1100 ;
      RECT 4.4200 24.0165 4.4460 25.1100 ;
      RECT 4.3120 24.0165 4.3380 25.1100 ;
      RECT 4.2040 24.0165 4.2300 25.1100 ;
      RECT 4.0960 24.0165 4.1220 25.1100 ;
      RECT 3.9880 24.0165 4.0140 25.1100 ;
      RECT 3.8800 24.0165 3.9060 25.1100 ;
      RECT 3.7720 24.0165 3.7980 25.1100 ;
      RECT 3.6640 24.0165 3.6900 25.1100 ;
      RECT 3.5560 24.0165 3.5820 25.1100 ;
      RECT 3.4480 24.0165 3.4740 25.1100 ;
      RECT 3.3400 24.0165 3.3660 25.1100 ;
      RECT 3.2320 24.0165 3.2580 25.1100 ;
      RECT 3.1240 24.0165 3.1500 25.1100 ;
      RECT 3.0160 24.0165 3.0420 25.1100 ;
      RECT 2.9080 24.0165 2.9340 25.1100 ;
      RECT 2.8000 24.0165 2.8260 25.1100 ;
      RECT 2.6920 24.0165 2.7180 25.1100 ;
      RECT 2.5840 24.0165 2.6100 25.1100 ;
      RECT 2.4760 24.0165 2.5020 25.1100 ;
      RECT 2.3680 24.0165 2.3940 25.1100 ;
      RECT 2.2600 24.0165 2.2860 25.1100 ;
      RECT 2.1520 24.0165 2.1780 25.1100 ;
      RECT 2.0440 24.0165 2.0700 25.1100 ;
      RECT 1.9360 24.0165 1.9620 25.1100 ;
      RECT 1.8280 24.0165 1.8540 25.1100 ;
      RECT 1.7200 24.0165 1.7460 25.1100 ;
      RECT 1.6120 24.0165 1.6380 25.1100 ;
      RECT 1.5040 24.0165 1.5300 25.1100 ;
      RECT 1.3960 24.0165 1.4220 25.1100 ;
      RECT 1.2880 24.0165 1.3140 25.1100 ;
      RECT 1.1800 24.0165 1.2060 25.1100 ;
      RECT 1.0720 24.0165 1.0980 25.1100 ;
      RECT 0.9640 24.0165 0.9900 25.1100 ;
      RECT 0.8560 24.0165 0.8820 25.1100 ;
      RECT 0.7480 24.0165 0.7740 25.1100 ;
      RECT 0.6400 24.0165 0.6660 25.1100 ;
      RECT 0.5320 24.0165 0.5580 25.1100 ;
      RECT 0.4240 24.0165 0.4500 25.1100 ;
      RECT 0.3160 24.0165 0.3420 25.1100 ;
      RECT 0.2080 24.0165 0.2340 25.1100 ;
      RECT 0.0050 24.0165 0.0900 25.1100 ;
      RECT 8.6410 25.0965 8.7690 26.1900 ;
      RECT 8.6270 25.7620 8.7690 26.0845 ;
      RECT 8.4790 25.4890 8.5410 26.1900 ;
      RECT 8.4650 25.7985 8.5410 25.9520 ;
      RECT 8.4790 25.0965 8.5050 26.1900 ;
      RECT 8.4790 25.2175 8.5190 25.4570 ;
      RECT 8.4790 25.0965 8.5410 25.1855 ;
      RECT 8.1820 25.5470 8.3880 26.1900 ;
      RECT 8.3620 25.0965 8.3880 26.1900 ;
      RECT 8.1820 25.8240 8.4020 26.0820 ;
      RECT 8.1820 25.0965 8.2800 26.1900 ;
      RECT 7.7650 25.0965 7.8480 26.1900 ;
      RECT 7.7650 25.1850 7.8620 26.1205 ;
      RECT 16.4440 25.0965 16.5290 26.1900 ;
      RECT 16.3000 25.0965 16.3260 26.1900 ;
      RECT 16.1920 25.0965 16.2180 26.1900 ;
      RECT 16.0840 25.0965 16.1100 26.1900 ;
      RECT 15.9760 25.0965 16.0020 26.1900 ;
      RECT 15.8680 25.0965 15.8940 26.1900 ;
      RECT 15.7600 25.0965 15.7860 26.1900 ;
      RECT 15.6520 25.0965 15.6780 26.1900 ;
      RECT 15.5440 25.0965 15.5700 26.1900 ;
      RECT 15.4360 25.0965 15.4620 26.1900 ;
      RECT 15.3280 25.0965 15.3540 26.1900 ;
      RECT 15.2200 25.0965 15.2460 26.1900 ;
      RECT 15.1120 25.0965 15.1380 26.1900 ;
      RECT 15.0040 25.0965 15.0300 26.1900 ;
      RECT 14.8960 25.0965 14.9220 26.1900 ;
      RECT 14.7880 25.0965 14.8140 26.1900 ;
      RECT 14.6800 25.0965 14.7060 26.1900 ;
      RECT 14.5720 25.0965 14.5980 26.1900 ;
      RECT 14.4640 25.0965 14.4900 26.1900 ;
      RECT 14.3560 25.0965 14.3820 26.1900 ;
      RECT 14.2480 25.0965 14.2740 26.1900 ;
      RECT 14.1400 25.0965 14.1660 26.1900 ;
      RECT 14.0320 25.0965 14.0580 26.1900 ;
      RECT 13.9240 25.0965 13.9500 26.1900 ;
      RECT 13.8160 25.0965 13.8420 26.1900 ;
      RECT 13.7080 25.0965 13.7340 26.1900 ;
      RECT 13.6000 25.0965 13.6260 26.1900 ;
      RECT 13.4920 25.0965 13.5180 26.1900 ;
      RECT 13.3840 25.0965 13.4100 26.1900 ;
      RECT 13.2760 25.0965 13.3020 26.1900 ;
      RECT 13.1680 25.0965 13.1940 26.1900 ;
      RECT 13.0600 25.0965 13.0860 26.1900 ;
      RECT 12.9520 25.0965 12.9780 26.1900 ;
      RECT 12.8440 25.0965 12.8700 26.1900 ;
      RECT 12.7360 25.0965 12.7620 26.1900 ;
      RECT 12.6280 25.0965 12.6540 26.1900 ;
      RECT 12.5200 25.0965 12.5460 26.1900 ;
      RECT 12.4120 25.0965 12.4380 26.1900 ;
      RECT 12.3040 25.0965 12.3300 26.1900 ;
      RECT 12.1960 25.0965 12.2220 26.1900 ;
      RECT 12.0880 25.0965 12.1140 26.1900 ;
      RECT 11.9800 25.0965 12.0060 26.1900 ;
      RECT 11.8720 25.0965 11.8980 26.1900 ;
      RECT 11.7640 25.0965 11.7900 26.1900 ;
      RECT 11.6560 25.0965 11.6820 26.1900 ;
      RECT 11.5480 25.0965 11.5740 26.1900 ;
      RECT 11.4400 25.0965 11.4660 26.1900 ;
      RECT 11.3320 25.0965 11.3580 26.1900 ;
      RECT 11.2240 25.0965 11.2500 26.1900 ;
      RECT 11.1160 25.0965 11.1420 26.1900 ;
      RECT 11.0080 25.0965 11.0340 26.1900 ;
      RECT 10.9000 25.0965 10.9260 26.1900 ;
      RECT 10.7920 25.0965 10.8180 26.1900 ;
      RECT 10.6840 25.0965 10.7100 26.1900 ;
      RECT 10.5760 25.0965 10.6020 26.1900 ;
      RECT 10.4680 25.0965 10.4940 26.1900 ;
      RECT 10.3600 25.0965 10.3860 26.1900 ;
      RECT 10.2520 25.0965 10.2780 26.1900 ;
      RECT 10.1440 25.0965 10.1700 26.1900 ;
      RECT 10.0360 25.0965 10.0620 26.1900 ;
      RECT 9.9280 25.0965 9.9540 26.1900 ;
      RECT 9.8200 25.0965 9.8460 26.1900 ;
      RECT 9.7120 25.0965 9.7380 26.1900 ;
      RECT 9.6040 25.0965 9.6300 26.1900 ;
      RECT 9.4960 25.0965 9.5220 26.1900 ;
      RECT 9.3880 25.0965 9.4140 26.1900 ;
      RECT 9.1750 25.0965 9.2520 26.1900 ;
      RECT 7.2820 25.0965 7.3590 26.1900 ;
      RECT 7.1200 25.0965 7.1460 26.1900 ;
      RECT 7.0120 25.0965 7.0380 26.1900 ;
      RECT 6.9040 25.0965 6.9300 26.1900 ;
      RECT 6.7960 25.0965 6.8220 26.1900 ;
      RECT 6.6880 25.0965 6.7140 26.1900 ;
      RECT 6.5800 25.0965 6.6060 26.1900 ;
      RECT 6.4720 25.0965 6.4980 26.1900 ;
      RECT 6.3640 25.0965 6.3900 26.1900 ;
      RECT 6.2560 25.0965 6.2820 26.1900 ;
      RECT 6.1480 25.0965 6.1740 26.1900 ;
      RECT 6.0400 25.0965 6.0660 26.1900 ;
      RECT 5.9320 25.0965 5.9580 26.1900 ;
      RECT 5.8240 25.0965 5.8500 26.1900 ;
      RECT 5.7160 25.0965 5.7420 26.1900 ;
      RECT 5.6080 25.0965 5.6340 26.1900 ;
      RECT 5.5000 25.0965 5.5260 26.1900 ;
      RECT 5.3920 25.0965 5.4180 26.1900 ;
      RECT 5.2840 25.0965 5.3100 26.1900 ;
      RECT 5.1760 25.0965 5.2020 26.1900 ;
      RECT 5.0680 25.0965 5.0940 26.1900 ;
      RECT 4.9600 25.0965 4.9860 26.1900 ;
      RECT 4.8520 25.0965 4.8780 26.1900 ;
      RECT 4.7440 25.0965 4.7700 26.1900 ;
      RECT 4.6360 25.0965 4.6620 26.1900 ;
      RECT 4.5280 25.0965 4.5540 26.1900 ;
      RECT 4.4200 25.0965 4.4460 26.1900 ;
      RECT 4.3120 25.0965 4.3380 26.1900 ;
      RECT 4.2040 25.0965 4.2300 26.1900 ;
      RECT 4.0960 25.0965 4.1220 26.1900 ;
      RECT 3.9880 25.0965 4.0140 26.1900 ;
      RECT 3.8800 25.0965 3.9060 26.1900 ;
      RECT 3.7720 25.0965 3.7980 26.1900 ;
      RECT 3.6640 25.0965 3.6900 26.1900 ;
      RECT 3.5560 25.0965 3.5820 26.1900 ;
      RECT 3.4480 25.0965 3.4740 26.1900 ;
      RECT 3.3400 25.0965 3.3660 26.1900 ;
      RECT 3.2320 25.0965 3.2580 26.1900 ;
      RECT 3.1240 25.0965 3.1500 26.1900 ;
      RECT 3.0160 25.0965 3.0420 26.1900 ;
      RECT 2.9080 25.0965 2.9340 26.1900 ;
      RECT 2.8000 25.0965 2.8260 26.1900 ;
      RECT 2.6920 25.0965 2.7180 26.1900 ;
      RECT 2.5840 25.0965 2.6100 26.1900 ;
      RECT 2.4760 25.0965 2.5020 26.1900 ;
      RECT 2.3680 25.0965 2.3940 26.1900 ;
      RECT 2.2600 25.0965 2.2860 26.1900 ;
      RECT 2.1520 25.0965 2.1780 26.1900 ;
      RECT 2.0440 25.0965 2.0700 26.1900 ;
      RECT 1.9360 25.0965 1.9620 26.1900 ;
      RECT 1.8280 25.0965 1.8540 26.1900 ;
      RECT 1.7200 25.0965 1.7460 26.1900 ;
      RECT 1.6120 25.0965 1.6380 26.1900 ;
      RECT 1.5040 25.0965 1.5300 26.1900 ;
      RECT 1.3960 25.0965 1.4220 26.1900 ;
      RECT 1.2880 25.0965 1.3140 26.1900 ;
      RECT 1.1800 25.0965 1.2060 26.1900 ;
      RECT 1.0720 25.0965 1.0980 26.1900 ;
      RECT 0.9640 25.0965 0.9900 26.1900 ;
      RECT 0.8560 25.0965 0.8820 26.1900 ;
      RECT 0.7480 25.0965 0.7740 26.1900 ;
      RECT 0.6400 25.0965 0.6660 26.1900 ;
      RECT 0.5320 25.0965 0.5580 26.1900 ;
      RECT 0.4240 25.0965 0.4500 26.1900 ;
      RECT 0.3160 25.0965 0.3420 26.1900 ;
      RECT 0.2080 25.0965 0.2340 26.1900 ;
      RECT 0.0050 25.0965 0.0900 26.1900 ;
      RECT 8.6410 26.1765 8.7690 27.2700 ;
      RECT 8.6270 26.8420 8.7690 27.1645 ;
      RECT 8.4790 26.5690 8.5410 27.2700 ;
      RECT 8.4650 26.8785 8.5410 27.0320 ;
      RECT 8.4790 26.1765 8.5050 27.2700 ;
      RECT 8.4790 26.2975 8.5190 26.5370 ;
      RECT 8.4790 26.1765 8.5410 26.2655 ;
      RECT 8.1820 26.6270 8.3880 27.2700 ;
      RECT 8.3620 26.1765 8.3880 27.2700 ;
      RECT 8.1820 26.9040 8.4020 27.1620 ;
      RECT 8.1820 26.1765 8.2800 27.2700 ;
      RECT 7.7650 26.1765 7.8480 27.2700 ;
      RECT 7.7650 26.2650 7.8620 27.2005 ;
      RECT 16.4440 26.1765 16.5290 27.2700 ;
      RECT 16.3000 26.1765 16.3260 27.2700 ;
      RECT 16.1920 26.1765 16.2180 27.2700 ;
      RECT 16.0840 26.1765 16.1100 27.2700 ;
      RECT 15.9760 26.1765 16.0020 27.2700 ;
      RECT 15.8680 26.1765 15.8940 27.2700 ;
      RECT 15.7600 26.1765 15.7860 27.2700 ;
      RECT 15.6520 26.1765 15.6780 27.2700 ;
      RECT 15.5440 26.1765 15.5700 27.2700 ;
      RECT 15.4360 26.1765 15.4620 27.2700 ;
      RECT 15.3280 26.1765 15.3540 27.2700 ;
      RECT 15.2200 26.1765 15.2460 27.2700 ;
      RECT 15.1120 26.1765 15.1380 27.2700 ;
      RECT 15.0040 26.1765 15.0300 27.2700 ;
      RECT 14.8960 26.1765 14.9220 27.2700 ;
      RECT 14.7880 26.1765 14.8140 27.2700 ;
      RECT 14.6800 26.1765 14.7060 27.2700 ;
      RECT 14.5720 26.1765 14.5980 27.2700 ;
      RECT 14.4640 26.1765 14.4900 27.2700 ;
      RECT 14.3560 26.1765 14.3820 27.2700 ;
      RECT 14.2480 26.1765 14.2740 27.2700 ;
      RECT 14.1400 26.1765 14.1660 27.2700 ;
      RECT 14.0320 26.1765 14.0580 27.2700 ;
      RECT 13.9240 26.1765 13.9500 27.2700 ;
      RECT 13.8160 26.1765 13.8420 27.2700 ;
      RECT 13.7080 26.1765 13.7340 27.2700 ;
      RECT 13.6000 26.1765 13.6260 27.2700 ;
      RECT 13.4920 26.1765 13.5180 27.2700 ;
      RECT 13.3840 26.1765 13.4100 27.2700 ;
      RECT 13.2760 26.1765 13.3020 27.2700 ;
      RECT 13.1680 26.1765 13.1940 27.2700 ;
      RECT 13.0600 26.1765 13.0860 27.2700 ;
      RECT 12.9520 26.1765 12.9780 27.2700 ;
      RECT 12.8440 26.1765 12.8700 27.2700 ;
      RECT 12.7360 26.1765 12.7620 27.2700 ;
      RECT 12.6280 26.1765 12.6540 27.2700 ;
      RECT 12.5200 26.1765 12.5460 27.2700 ;
      RECT 12.4120 26.1765 12.4380 27.2700 ;
      RECT 12.3040 26.1765 12.3300 27.2700 ;
      RECT 12.1960 26.1765 12.2220 27.2700 ;
      RECT 12.0880 26.1765 12.1140 27.2700 ;
      RECT 11.9800 26.1765 12.0060 27.2700 ;
      RECT 11.8720 26.1765 11.8980 27.2700 ;
      RECT 11.7640 26.1765 11.7900 27.2700 ;
      RECT 11.6560 26.1765 11.6820 27.2700 ;
      RECT 11.5480 26.1765 11.5740 27.2700 ;
      RECT 11.4400 26.1765 11.4660 27.2700 ;
      RECT 11.3320 26.1765 11.3580 27.2700 ;
      RECT 11.2240 26.1765 11.2500 27.2700 ;
      RECT 11.1160 26.1765 11.1420 27.2700 ;
      RECT 11.0080 26.1765 11.0340 27.2700 ;
      RECT 10.9000 26.1765 10.9260 27.2700 ;
      RECT 10.7920 26.1765 10.8180 27.2700 ;
      RECT 10.6840 26.1765 10.7100 27.2700 ;
      RECT 10.5760 26.1765 10.6020 27.2700 ;
      RECT 10.4680 26.1765 10.4940 27.2700 ;
      RECT 10.3600 26.1765 10.3860 27.2700 ;
      RECT 10.2520 26.1765 10.2780 27.2700 ;
      RECT 10.1440 26.1765 10.1700 27.2700 ;
      RECT 10.0360 26.1765 10.0620 27.2700 ;
      RECT 9.9280 26.1765 9.9540 27.2700 ;
      RECT 9.8200 26.1765 9.8460 27.2700 ;
      RECT 9.7120 26.1765 9.7380 27.2700 ;
      RECT 9.6040 26.1765 9.6300 27.2700 ;
      RECT 9.4960 26.1765 9.5220 27.2700 ;
      RECT 9.3880 26.1765 9.4140 27.2700 ;
      RECT 9.1750 26.1765 9.2520 27.2700 ;
      RECT 7.2820 26.1765 7.3590 27.2700 ;
      RECT 7.1200 26.1765 7.1460 27.2700 ;
      RECT 7.0120 26.1765 7.0380 27.2700 ;
      RECT 6.9040 26.1765 6.9300 27.2700 ;
      RECT 6.7960 26.1765 6.8220 27.2700 ;
      RECT 6.6880 26.1765 6.7140 27.2700 ;
      RECT 6.5800 26.1765 6.6060 27.2700 ;
      RECT 6.4720 26.1765 6.4980 27.2700 ;
      RECT 6.3640 26.1765 6.3900 27.2700 ;
      RECT 6.2560 26.1765 6.2820 27.2700 ;
      RECT 6.1480 26.1765 6.1740 27.2700 ;
      RECT 6.0400 26.1765 6.0660 27.2700 ;
      RECT 5.9320 26.1765 5.9580 27.2700 ;
      RECT 5.8240 26.1765 5.8500 27.2700 ;
      RECT 5.7160 26.1765 5.7420 27.2700 ;
      RECT 5.6080 26.1765 5.6340 27.2700 ;
      RECT 5.5000 26.1765 5.5260 27.2700 ;
      RECT 5.3920 26.1765 5.4180 27.2700 ;
      RECT 5.2840 26.1765 5.3100 27.2700 ;
      RECT 5.1760 26.1765 5.2020 27.2700 ;
      RECT 5.0680 26.1765 5.0940 27.2700 ;
      RECT 4.9600 26.1765 4.9860 27.2700 ;
      RECT 4.8520 26.1765 4.8780 27.2700 ;
      RECT 4.7440 26.1765 4.7700 27.2700 ;
      RECT 4.6360 26.1765 4.6620 27.2700 ;
      RECT 4.5280 26.1765 4.5540 27.2700 ;
      RECT 4.4200 26.1765 4.4460 27.2700 ;
      RECT 4.3120 26.1765 4.3380 27.2700 ;
      RECT 4.2040 26.1765 4.2300 27.2700 ;
      RECT 4.0960 26.1765 4.1220 27.2700 ;
      RECT 3.9880 26.1765 4.0140 27.2700 ;
      RECT 3.8800 26.1765 3.9060 27.2700 ;
      RECT 3.7720 26.1765 3.7980 27.2700 ;
      RECT 3.6640 26.1765 3.6900 27.2700 ;
      RECT 3.5560 26.1765 3.5820 27.2700 ;
      RECT 3.4480 26.1765 3.4740 27.2700 ;
      RECT 3.3400 26.1765 3.3660 27.2700 ;
      RECT 3.2320 26.1765 3.2580 27.2700 ;
      RECT 3.1240 26.1765 3.1500 27.2700 ;
      RECT 3.0160 26.1765 3.0420 27.2700 ;
      RECT 2.9080 26.1765 2.9340 27.2700 ;
      RECT 2.8000 26.1765 2.8260 27.2700 ;
      RECT 2.6920 26.1765 2.7180 27.2700 ;
      RECT 2.5840 26.1765 2.6100 27.2700 ;
      RECT 2.4760 26.1765 2.5020 27.2700 ;
      RECT 2.3680 26.1765 2.3940 27.2700 ;
      RECT 2.2600 26.1765 2.2860 27.2700 ;
      RECT 2.1520 26.1765 2.1780 27.2700 ;
      RECT 2.0440 26.1765 2.0700 27.2700 ;
      RECT 1.9360 26.1765 1.9620 27.2700 ;
      RECT 1.8280 26.1765 1.8540 27.2700 ;
      RECT 1.7200 26.1765 1.7460 27.2700 ;
      RECT 1.6120 26.1765 1.6380 27.2700 ;
      RECT 1.5040 26.1765 1.5300 27.2700 ;
      RECT 1.3960 26.1765 1.4220 27.2700 ;
      RECT 1.2880 26.1765 1.3140 27.2700 ;
      RECT 1.1800 26.1765 1.2060 27.2700 ;
      RECT 1.0720 26.1765 1.0980 27.2700 ;
      RECT 0.9640 26.1765 0.9900 27.2700 ;
      RECT 0.8560 26.1765 0.8820 27.2700 ;
      RECT 0.7480 26.1765 0.7740 27.2700 ;
      RECT 0.6400 26.1765 0.6660 27.2700 ;
      RECT 0.5320 26.1765 0.5580 27.2700 ;
      RECT 0.4240 26.1765 0.4500 27.2700 ;
      RECT 0.3160 26.1765 0.3420 27.2700 ;
      RECT 0.2080 26.1765 0.2340 27.2700 ;
      RECT 0.0050 26.1765 0.0900 27.2700 ;
      RECT 8.6410 27.2565 8.7690 28.3500 ;
      RECT 8.6270 27.9220 8.7690 28.2445 ;
      RECT 8.4790 27.6490 8.5410 28.3500 ;
      RECT 8.4650 27.9585 8.5410 28.1120 ;
      RECT 8.4790 27.2565 8.5050 28.3500 ;
      RECT 8.4790 27.3775 8.5190 27.6170 ;
      RECT 8.4790 27.2565 8.5410 27.3455 ;
      RECT 8.1820 27.7070 8.3880 28.3500 ;
      RECT 8.3620 27.2565 8.3880 28.3500 ;
      RECT 8.1820 27.9840 8.4020 28.2420 ;
      RECT 8.1820 27.2565 8.2800 28.3500 ;
      RECT 7.7650 27.2565 7.8480 28.3500 ;
      RECT 7.7650 27.3450 7.8620 28.2805 ;
      RECT 16.4440 27.2565 16.5290 28.3500 ;
      RECT 16.3000 27.2565 16.3260 28.3500 ;
      RECT 16.1920 27.2565 16.2180 28.3500 ;
      RECT 16.0840 27.2565 16.1100 28.3500 ;
      RECT 15.9760 27.2565 16.0020 28.3500 ;
      RECT 15.8680 27.2565 15.8940 28.3500 ;
      RECT 15.7600 27.2565 15.7860 28.3500 ;
      RECT 15.6520 27.2565 15.6780 28.3500 ;
      RECT 15.5440 27.2565 15.5700 28.3500 ;
      RECT 15.4360 27.2565 15.4620 28.3500 ;
      RECT 15.3280 27.2565 15.3540 28.3500 ;
      RECT 15.2200 27.2565 15.2460 28.3500 ;
      RECT 15.1120 27.2565 15.1380 28.3500 ;
      RECT 15.0040 27.2565 15.0300 28.3500 ;
      RECT 14.8960 27.2565 14.9220 28.3500 ;
      RECT 14.7880 27.2565 14.8140 28.3500 ;
      RECT 14.6800 27.2565 14.7060 28.3500 ;
      RECT 14.5720 27.2565 14.5980 28.3500 ;
      RECT 14.4640 27.2565 14.4900 28.3500 ;
      RECT 14.3560 27.2565 14.3820 28.3500 ;
      RECT 14.2480 27.2565 14.2740 28.3500 ;
      RECT 14.1400 27.2565 14.1660 28.3500 ;
      RECT 14.0320 27.2565 14.0580 28.3500 ;
      RECT 13.9240 27.2565 13.9500 28.3500 ;
      RECT 13.8160 27.2565 13.8420 28.3500 ;
      RECT 13.7080 27.2565 13.7340 28.3500 ;
      RECT 13.6000 27.2565 13.6260 28.3500 ;
      RECT 13.4920 27.2565 13.5180 28.3500 ;
      RECT 13.3840 27.2565 13.4100 28.3500 ;
      RECT 13.2760 27.2565 13.3020 28.3500 ;
      RECT 13.1680 27.2565 13.1940 28.3500 ;
      RECT 13.0600 27.2565 13.0860 28.3500 ;
      RECT 12.9520 27.2565 12.9780 28.3500 ;
      RECT 12.8440 27.2565 12.8700 28.3500 ;
      RECT 12.7360 27.2565 12.7620 28.3500 ;
      RECT 12.6280 27.2565 12.6540 28.3500 ;
      RECT 12.5200 27.2565 12.5460 28.3500 ;
      RECT 12.4120 27.2565 12.4380 28.3500 ;
      RECT 12.3040 27.2565 12.3300 28.3500 ;
      RECT 12.1960 27.2565 12.2220 28.3500 ;
      RECT 12.0880 27.2565 12.1140 28.3500 ;
      RECT 11.9800 27.2565 12.0060 28.3500 ;
      RECT 11.8720 27.2565 11.8980 28.3500 ;
      RECT 11.7640 27.2565 11.7900 28.3500 ;
      RECT 11.6560 27.2565 11.6820 28.3500 ;
      RECT 11.5480 27.2565 11.5740 28.3500 ;
      RECT 11.4400 27.2565 11.4660 28.3500 ;
      RECT 11.3320 27.2565 11.3580 28.3500 ;
      RECT 11.2240 27.2565 11.2500 28.3500 ;
      RECT 11.1160 27.2565 11.1420 28.3500 ;
      RECT 11.0080 27.2565 11.0340 28.3500 ;
      RECT 10.9000 27.2565 10.9260 28.3500 ;
      RECT 10.7920 27.2565 10.8180 28.3500 ;
      RECT 10.6840 27.2565 10.7100 28.3500 ;
      RECT 10.5760 27.2565 10.6020 28.3500 ;
      RECT 10.4680 27.2565 10.4940 28.3500 ;
      RECT 10.3600 27.2565 10.3860 28.3500 ;
      RECT 10.2520 27.2565 10.2780 28.3500 ;
      RECT 10.1440 27.2565 10.1700 28.3500 ;
      RECT 10.0360 27.2565 10.0620 28.3500 ;
      RECT 9.9280 27.2565 9.9540 28.3500 ;
      RECT 9.8200 27.2565 9.8460 28.3500 ;
      RECT 9.7120 27.2565 9.7380 28.3500 ;
      RECT 9.6040 27.2565 9.6300 28.3500 ;
      RECT 9.4960 27.2565 9.5220 28.3500 ;
      RECT 9.3880 27.2565 9.4140 28.3500 ;
      RECT 9.1750 27.2565 9.2520 28.3500 ;
      RECT 7.2820 27.2565 7.3590 28.3500 ;
      RECT 7.1200 27.2565 7.1460 28.3500 ;
      RECT 7.0120 27.2565 7.0380 28.3500 ;
      RECT 6.9040 27.2565 6.9300 28.3500 ;
      RECT 6.7960 27.2565 6.8220 28.3500 ;
      RECT 6.6880 27.2565 6.7140 28.3500 ;
      RECT 6.5800 27.2565 6.6060 28.3500 ;
      RECT 6.4720 27.2565 6.4980 28.3500 ;
      RECT 6.3640 27.2565 6.3900 28.3500 ;
      RECT 6.2560 27.2565 6.2820 28.3500 ;
      RECT 6.1480 27.2565 6.1740 28.3500 ;
      RECT 6.0400 27.2565 6.0660 28.3500 ;
      RECT 5.9320 27.2565 5.9580 28.3500 ;
      RECT 5.8240 27.2565 5.8500 28.3500 ;
      RECT 5.7160 27.2565 5.7420 28.3500 ;
      RECT 5.6080 27.2565 5.6340 28.3500 ;
      RECT 5.5000 27.2565 5.5260 28.3500 ;
      RECT 5.3920 27.2565 5.4180 28.3500 ;
      RECT 5.2840 27.2565 5.3100 28.3500 ;
      RECT 5.1760 27.2565 5.2020 28.3500 ;
      RECT 5.0680 27.2565 5.0940 28.3500 ;
      RECT 4.9600 27.2565 4.9860 28.3500 ;
      RECT 4.8520 27.2565 4.8780 28.3500 ;
      RECT 4.7440 27.2565 4.7700 28.3500 ;
      RECT 4.6360 27.2565 4.6620 28.3500 ;
      RECT 4.5280 27.2565 4.5540 28.3500 ;
      RECT 4.4200 27.2565 4.4460 28.3500 ;
      RECT 4.3120 27.2565 4.3380 28.3500 ;
      RECT 4.2040 27.2565 4.2300 28.3500 ;
      RECT 4.0960 27.2565 4.1220 28.3500 ;
      RECT 3.9880 27.2565 4.0140 28.3500 ;
      RECT 3.8800 27.2565 3.9060 28.3500 ;
      RECT 3.7720 27.2565 3.7980 28.3500 ;
      RECT 3.6640 27.2565 3.6900 28.3500 ;
      RECT 3.5560 27.2565 3.5820 28.3500 ;
      RECT 3.4480 27.2565 3.4740 28.3500 ;
      RECT 3.3400 27.2565 3.3660 28.3500 ;
      RECT 3.2320 27.2565 3.2580 28.3500 ;
      RECT 3.1240 27.2565 3.1500 28.3500 ;
      RECT 3.0160 27.2565 3.0420 28.3500 ;
      RECT 2.9080 27.2565 2.9340 28.3500 ;
      RECT 2.8000 27.2565 2.8260 28.3500 ;
      RECT 2.6920 27.2565 2.7180 28.3500 ;
      RECT 2.5840 27.2565 2.6100 28.3500 ;
      RECT 2.4760 27.2565 2.5020 28.3500 ;
      RECT 2.3680 27.2565 2.3940 28.3500 ;
      RECT 2.2600 27.2565 2.2860 28.3500 ;
      RECT 2.1520 27.2565 2.1780 28.3500 ;
      RECT 2.0440 27.2565 2.0700 28.3500 ;
      RECT 1.9360 27.2565 1.9620 28.3500 ;
      RECT 1.8280 27.2565 1.8540 28.3500 ;
      RECT 1.7200 27.2565 1.7460 28.3500 ;
      RECT 1.6120 27.2565 1.6380 28.3500 ;
      RECT 1.5040 27.2565 1.5300 28.3500 ;
      RECT 1.3960 27.2565 1.4220 28.3500 ;
      RECT 1.2880 27.2565 1.3140 28.3500 ;
      RECT 1.1800 27.2565 1.2060 28.3500 ;
      RECT 1.0720 27.2565 1.0980 28.3500 ;
      RECT 0.9640 27.2565 0.9900 28.3500 ;
      RECT 0.8560 27.2565 0.8820 28.3500 ;
      RECT 0.7480 27.2565 0.7740 28.3500 ;
      RECT 0.6400 27.2565 0.6660 28.3500 ;
      RECT 0.5320 27.2565 0.5580 28.3500 ;
      RECT 0.4240 27.2565 0.4500 28.3500 ;
      RECT 0.3160 27.2565 0.3420 28.3500 ;
      RECT 0.2080 27.2565 0.2340 28.3500 ;
      RECT 0.0050 27.2565 0.0900 28.3500 ;
      RECT 8.6410 28.3365 8.7690 29.4300 ;
      RECT 8.6270 29.0020 8.7690 29.3245 ;
      RECT 8.4790 28.7290 8.5410 29.4300 ;
      RECT 8.4650 29.0385 8.5410 29.1920 ;
      RECT 8.4790 28.3365 8.5050 29.4300 ;
      RECT 8.4790 28.4575 8.5190 28.6970 ;
      RECT 8.4790 28.3365 8.5410 28.4255 ;
      RECT 8.1820 28.7870 8.3880 29.4300 ;
      RECT 8.3620 28.3365 8.3880 29.4300 ;
      RECT 8.1820 29.0640 8.4020 29.3220 ;
      RECT 8.1820 28.3365 8.2800 29.4300 ;
      RECT 7.7650 28.3365 7.8480 29.4300 ;
      RECT 7.7650 28.4250 7.8620 29.3605 ;
      RECT 16.4440 28.3365 16.5290 29.4300 ;
      RECT 16.3000 28.3365 16.3260 29.4300 ;
      RECT 16.1920 28.3365 16.2180 29.4300 ;
      RECT 16.0840 28.3365 16.1100 29.4300 ;
      RECT 15.9760 28.3365 16.0020 29.4300 ;
      RECT 15.8680 28.3365 15.8940 29.4300 ;
      RECT 15.7600 28.3365 15.7860 29.4300 ;
      RECT 15.6520 28.3365 15.6780 29.4300 ;
      RECT 15.5440 28.3365 15.5700 29.4300 ;
      RECT 15.4360 28.3365 15.4620 29.4300 ;
      RECT 15.3280 28.3365 15.3540 29.4300 ;
      RECT 15.2200 28.3365 15.2460 29.4300 ;
      RECT 15.1120 28.3365 15.1380 29.4300 ;
      RECT 15.0040 28.3365 15.0300 29.4300 ;
      RECT 14.8960 28.3365 14.9220 29.4300 ;
      RECT 14.7880 28.3365 14.8140 29.4300 ;
      RECT 14.6800 28.3365 14.7060 29.4300 ;
      RECT 14.5720 28.3365 14.5980 29.4300 ;
      RECT 14.4640 28.3365 14.4900 29.4300 ;
      RECT 14.3560 28.3365 14.3820 29.4300 ;
      RECT 14.2480 28.3365 14.2740 29.4300 ;
      RECT 14.1400 28.3365 14.1660 29.4300 ;
      RECT 14.0320 28.3365 14.0580 29.4300 ;
      RECT 13.9240 28.3365 13.9500 29.4300 ;
      RECT 13.8160 28.3365 13.8420 29.4300 ;
      RECT 13.7080 28.3365 13.7340 29.4300 ;
      RECT 13.6000 28.3365 13.6260 29.4300 ;
      RECT 13.4920 28.3365 13.5180 29.4300 ;
      RECT 13.3840 28.3365 13.4100 29.4300 ;
      RECT 13.2760 28.3365 13.3020 29.4300 ;
      RECT 13.1680 28.3365 13.1940 29.4300 ;
      RECT 13.0600 28.3365 13.0860 29.4300 ;
      RECT 12.9520 28.3365 12.9780 29.4300 ;
      RECT 12.8440 28.3365 12.8700 29.4300 ;
      RECT 12.7360 28.3365 12.7620 29.4300 ;
      RECT 12.6280 28.3365 12.6540 29.4300 ;
      RECT 12.5200 28.3365 12.5460 29.4300 ;
      RECT 12.4120 28.3365 12.4380 29.4300 ;
      RECT 12.3040 28.3365 12.3300 29.4300 ;
      RECT 12.1960 28.3365 12.2220 29.4300 ;
      RECT 12.0880 28.3365 12.1140 29.4300 ;
      RECT 11.9800 28.3365 12.0060 29.4300 ;
      RECT 11.8720 28.3365 11.8980 29.4300 ;
      RECT 11.7640 28.3365 11.7900 29.4300 ;
      RECT 11.6560 28.3365 11.6820 29.4300 ;
      RECT 11.5480 28.3365 11.5740 29.4300 ;
      RECT 11.4400 28.3365 11.4660 29.4300 ;
      RECT 11.3320 28.3365 11.3580 29.4300 ;
      RECT 11.2240 28.3365 11.2500 29.4300 ;
      RECT 11.1160 28.3365 11.1420 29.4300 ;
      RECT 11.0080 28.3365 11.0340 29.4300 ;
      RECT 10.9000 28.3365 10.9260 29.4300 ;
      RECT 10.7920 28.3365 10.8180 29.4300 ;
      RECT 10.6840 28.3365 10.7100 29.4300 ;
      RECT 10.5760 28.3365 10.6020 29.4300 ;
      RECT 10.4680 28.3365 10.4940 29.4300 ;
      RECT 10.3600 28.3365 10.3860 29.4300 ;
      RECT 10.2520 28.3365 10.2780 29.4300 ;
      RECT 10.1440 28.3365 10.1700 29.4300 ;
      RECT 10.0360 28.3365 10.0620 29.4300 ;
      RECT 9.9280 28.3365 9.9540 29.4300 ;
      RECT 9.8200 28.3365 9.8460 29.4300 ;
      RECT 9.7120 28.3365 9.7380 29.4300 ;
      RECT 9.6040 28.3365 9.6300 29.4300 ;
      RECT 9.4960 28.3365 9.5220 29.4300 ;
      RECT 9.3880 28.3365 9.4140 29.4300 ;
      RECT 9.1750 28.3365 9.2520 29.4300 ;
      RECT 7.2820 28.3365 7.3590 29.4300 ;
      RECT 7.1200 28.3365 7.1460 29.4300 ;
      RECT 7.0120 28.3365 7.0380 29.4300 ;
      RECT 6.9040 28.3365 6.9300 29.4300 ;
      RECT 6.7960 28.3365 6.8220 29.4300 ;
      RECT 6.6880 28.3365 6.7140 29.4300 ;
      RECT 6.5800 28.3365 6.6060 29.4300 ;
      RECT 6.4720 28.3365 6.4980 29.4300 ;
      RECT 6.3640 28.3365 6.3900 29.4300 ;
      RECT 6.2560 28.3365 6.2820 29.4300 ;
      RECT 6.1480 28.3365 6.1740 29.4300 ;
      RECT 6.0400 28.3365 6.0660 29.4300 ;
      RECT 5.9320 28.3365 5.9580 29.4300 ;
      RECT 5.8240 28.3365 5.8500 29.4300 ;
      RECT 5.7160 28.3365 5.7420 29.4300 ;
      RECT 5.6080 28.3365 5.6340 29.4300 ;
      RECT 5.5000 28.3365 5.5260 29.4300 ;
      RECT 5.3920 28.3365 5.4180 29.4300 ;
      RECT 5.2840 28.3365 5.3100 29.4300 ;
      RECT 5.1760 28.3365 5.2020 29.4300 ;
      RECT 5.0680 28.3365 5.0940 29.4300 ;
      RECT 4.9600 28.3365 4.9860 29.4300 ;
      RECT 4.8520 28.3365 4.8780 29.4300 ;
      RECT 4.7440 28.3365 4.7700 29.4300 ;
      RECT 4.6360 28.3365 4.6620 29.4300 ;
      RECT 4.5280 28.3365 4.5540 29.4300 ;
      RECT 4.4200 28.3365 4.4460 29.4300 ;
      RECT 4.3120 28.3365 4.3380 29.4300 ;
      RECT 4.2040 28.3365 4.2300 29.4300 ;
      RECT 4.0960 28.3365 4.1220 29.4300 ;
      RECT 3.9880 28.3365 4.0140 29.4300 ;
      RECT 3.8800 28.3365 3.9060 29.4300 ;
      RECT 3.7720 28.3365 3.7980 29.4300 ;
      RECT 3.6640 28.3365 3.6900 29.4300 ;
      RECT 3.5560 28.3365 3.5820 29.4300 ;
      RECT 3.4480 28.3365 3.4740 29.4300 ;
      RECT 3.3400 28.3365 3.3660 29.4300 ;
      RECT 3.2320 28.3365 3.2580 29.4300 ;
      RECT 3.1240 28.3365 3.1500 29.4300 ;
      RECT 3.0160 28.3365 3.0420 29.4300 ;
      RECT 2.9080 28.3365 2.9340 29.4300 ;
      RECT 2.8000 28.3365 2.8260 29.4300 ;
      RECT 2.6920 28.3365 2.7180 29.4300 ;
      RECT 2.5840 28.3365 2.6100 29.4300 ;
      RECT 2.4760 28.3365 2.5020 29.4300 ;
      RECT 2.3680 28.3365 2.3940 29.4300 ;
      RECT 2.2600 28.3365 2.2860 29.4300 ;
      RECT 2.1520 28.3365 2.1780 29.4300 ;
      RECT 2.0440 28.3365 2.0700 29.4300 ;
      RECT 1.9360 28.3365 1.9620 29.4300 ;
      RECT 1.8280 28.3365 1.8540 29.4300 ;
      RECT 1.7200 28.3365 1.7460 29.4300 ;
      RECT 1.6120 28.3365 1.6380 29.4300 ;
      RECT 1.5040 28.3365 1.5300 29.4300 ;
      RECT 1.3960 28.3365 1.4220 29.4300 ;
      RECT 1.2880 28.3365 1.3140 29.4300 ;
      RECT 1.1800 28.3365 1.2060 29.4300 ;
      RECT 1.0720 28.3365 1.0980 29.4300 ;
      RECT 0.9640 28.3365 0.9900 29.4300 ;
      RECT 0.8560 28.3365 0.8820 29.4300 ;
      RECT 0.7480 28.3365 0.7740 29.4300 ;
      RECT 0.6400 28.3365 0.6660 29.4300 ;
      RECT 0.5320 28.3365 0.5580 29.4300 ;
      RECT 0.4240 28.3365 0.4500 29.4300 ;
      RECT 0.3160 28.3365 0.3420 29.4300 ;
      RECT 0.2080 28.3365 0.2340 29.4300 ;
      RECT 0.0050 28.3365 0.0900 29.4300 ;
      RECT 8.6410 29.4165 8.7690 30.5100 ;
      RECT 8.6270 30.0820 8.7690 30.4045 ;
      RECT 8.4790 29.8090 8.5410 30.5100 ;
      RECT 8.4650 30.1185 8.5410 30.2720 ;
      RECT 8.4790 29.4165 8.5050 30.5100 ;
      RECT 8.4790 29.5375 8.5190 29.7770 ;
      RECT 8.4790 29.4165 8.5410 29.5055 ;
      RECT 8.1820 29.8670 8.3880 30.5100 ;
      RECT 8.3620 29.4165 8.3880 30.5100 ;
      RECT 8.1820 30.1440 8.4020 30.4020 ;
      RECT 8.1820 29.4165 8.2800 30.5100 ;
      RECT 7.7650 29.4165 7.8480 30.5100 ;
      RECT 7.7650 29.5050 7.8620 30.4405 ;
      RECT 16.4440 29.4165 16.5290 30.5100 ;
      RECT 16.3000 29.4165 16.3260 30.5100 ;
      RECT 16.1920 29.4165 16.2180 30.5100 ;
      RECT 16.0840 29.4165 16.1100 30.5100 ;
      RECT 15.9760 29.4165 16.0020 30.5100 ;
      RECT 15.8680 29.4165 15.8940 30.5100 ;
      RECT 15.7600 29.4165 15.7860 30.5100 ;
      RECT 15.6520 29.4165 15.6780 30.5100 ;
      RECT 15.5440 29.4165 15.5700 30.5100 ;
      RECT 15.4360 29.4165 15.4620 30.5100 ;
      RECT 15.3280 29.4165 15.3540 30.5100 ;
      RECT 15.2200 29.4165 15.2460 30.5100 ;
      RECT 15.1120 29.4165 15.1380 30.5100 ;
      RECT 15.0040 29.4165 15.0300 30.5100 ;
      RECT 14.8960 29.4165 14.9220 30.5100 ;
      RECT 14.7880 29.4165 14.8140 30.5100 ;
      RECT 14.6800 29.4165 14.7060 30.5100 ;
      RECT 14.5720 29.4165 14.5980 30.5100 ;
      RECT 14.4640 29.4165 14.4900 30.5100 ;
      RECT 14.3560 29.4165 14.3820 30.5100 ;
      RECT 14.2480 29.4165 14.2740 30.5100 ;
      RECT 14.1400 29.4165 14.1660 30.5100 ;
      RECT 14.0320 29.4165 14.0580 30.5100 ;
      RECT 13.9240 29.4165 13.9500 30.5100 ;
      RECT 13.8160 29.4165 13.8420 30.5100 ;
      RECT 13.7080 29.4165 13.7340 30.5100 ;
      RECT 13.6000 29.4165 13.6260 30.5100 ;
      RECT 13.4920 29.4165 13.5180 30.5100 ;
      RECT 13.3840 29.4165 13.4100 30.5100 ;
      RECT 13.2760 29.4165 13.3020 30.5100 ;
      RECT 13.1680 29.4165 13.1940 30.5100 ;
      RECT 13.0600 29.4165 13.0860 30.5100 ;
      RECT 12.9520 29.4165 12.9780 30.5100 ;
      RECT 12.8440 29.4165 12.8700 30.5100 ;
      RECT 12.7360 29.4165 12.7620 30.5100 ;
      RECT 12.6280 29.4165 12.6540 30.5100 ;
      RECT 12.5200 29.4165 12.5460 30.5100 ;
      RECT 12.4120 29.4165 12.4380 30.5100 ;
      RECT 12.3040 29.4165 12.3300 30.5100 ;
      RECT 12.1960 29.4165 12.2220 30.5100 ;
      RECT 12.0880 29.4165 12.1140 30.5100 ;
      RECT 11.9800 29.4165 12.0060 30.5100 ;
      RECT 11.8720 29.4165 11.8980 30.5100 ;
      RECT 11.7640 29.4165 11.7900 30.5100 ;
      RECT 11.6560 29.4165 11.6820 30.5100 ;
      RECT 11.5480 29.4165 11.5740 30.5100 ;
      RECT 11.4400 29.4165 11.4660 30.5100 ;
      RECT 11.3320 29.4165 11.3580 30.5100 ;
      RECT 11.2240 29.4165 11.2500 30.5100 ;
      RECT 11.1160 29.4165 11.1420 30.5100 ;
      RECT 11.0080 29.4165 11.0340 30.5100 ;
      RECT 10.9000 29.4165 10.9260 30.5100 ;
      RECT 10.7920 29.4165 10.8180 30.5100 ;
      RECT 10.6840 29.4165 10.7100 30.5100 ;
      RECT 10.5760 29.4165 10.6020 30.5100 ;
      RECT 10.4680 29.4165 10.4940 30.5100 ;
      RECT 10.3600 29.4165 10.3860 30.5100 ;
      RECT 10.2520 29.4165 10.2780 30.5100 ;
      RECT 10.1440 29.4165 10.1700 30.5100 ;
      RECT 10.0360 29.4165 10.0620 30.5100 ;
      RECT 9.9280 29.4165 9.9540 30.5100 ;
      RECT 9.8200 29.4165 9.8460 30.5100 ;
      RECT 9.7120 29.4165 9.7380 30.5100 ;
      RECT 9.6040 29.4165 9.6300 30.5100 ;
      RECT 9.4960 29.4165 9.5220 30.5100 ;
      RECT 9.3880 29.4165 9.4140 30.5100 ;
      RECT 9.1750 29.4165 9.2520 30.5100 ;
      RECT 7.2820 29.4165 7.3590 30.5100 ;
      RECT 7.1200 29.4165 7.1460 30.5100 ;
      RECT 7.0120 29.4165 7.0380 30.5100 ;
      RECT 6.9040 29.4165 6.9300 30.5100 ;
      RECT 6.7960 29.4165 6.8220 30.5100 ;
      RECT 6.6880 29.4165 6.7140 30.5100 ;
      RECT 6.5800 29.4165 6.6060 30.5100 ;
      RECT 6.4720 29.4165 6.4980 30.5100 ;
      RECT 6.3640 29.4165 6.3900 30.5100 ;
      RECT 6.2560 29.4165 6.2820 30.5100 ;
      RECT 6.1480 29.4165 6.1740 30.5100 ;
      RECT 6.0400 29.4165 6.0660 30.5100 ;
      RECT 5.9320 29.4165 5.9580 30.5100 ;
      RECT 5.8240 29.4165 5.8500 30.5100 ;
      RECT 5.7160 29.4165 5.7420 30.5100 ;
      RECT 5.6080 29.4165 5.6340 30.5100 ;
      RECT 5.5000 29.4165 5.5260 30.5100 ;
      RECT 5.3920 29.4165 5.4180 30.5100 ;
      RECT 5.2840 29.4165 5.3100 30.5100 ;
      RECT 5.1760 29.4165 5.2020 30.5100 ;
      RECT 5.0680 29.4165 5.0940 30.5100 ;
      RECT 4.9600 29.4165 4.9860 30.5100 ;
      RECT 4.8520 29.4165 4.8780 30.5100 ;
      RECT 4.7440 29.4165 4.7700 30.5100 ;
      RECT 4.6360 29.4165 4.6620 30.5100 ;
      RECT 4.5280 29.4165 4.5540 30.5100 ;
      RECT 4.4200 29.4165 4.4460 30.5100 ;
      RECT 4.3120 29.4165 4.3380 30.5100 ;
      RECT 4.2040 29.4165 4.2300 30.5100 ;
      RECT 4.0960 29.4165 4.1220 30.5100 ;
      RECT 3.9880 29.4165 4.0140 30.5100 ;
      RECT 3.8800 29.4165 3.9060 30.5100 ;
      RECT 3.7720 29.4165 3.7980 30.5100 ;
      RECT 3.6640 29.4165 3.6900 30.5100 ;
      RECT 3.5560 29.4165 3.5820 30.5100 ;
      RECT 3.4480 29.4165 3.4740 30.5100 ;
      RECT 3.3400 29.4165 3.3660 30.5100 ;
      RECT 3.2320 29.4165 3.2580 30.5100 ;
      RECT 3.1240 29.4165 3.1500 30.5100 ;
      RECT 3.0160 29.4165 3.0420 30.5100 ;
      RECT 2.9080 29.4165 2.9340 30.5100 ;
      RECT 2.8000 29.4165 2.8260 30.5100 ;
      RECT 2.6920 29.4165 2.7180 30.5100 ;
      RECT 2.5840 29.4165 2.6100 30.5100 ;
      RECT 2.4760 29.4165 2.5020 30.5100 ;
      RECT 2.3680 29.4165 2.3940 30.5100 ;
      RECT 2.2600 29.4165 2.2860 30.5100 ;
      RECT 2.1520 29.4165 2.1780 30.5100 ;
      RECT 2.0440 29.4165 2.0700 30.5100 ;
      RECT 1.9360 29.4165 1.9620 30.5100 ;
      RECT 1.8280 29.4165 1.8540 30.5100 ;
      RECT 1.7200 29.4165 1.7460 30.5100 ;
      RECT 1.6120 29.4165 1.6380 30.5100 ;
      RECT 1.5040 29.4165 1.5300 30.5100 ;
      RECT 1.3960 29.4165 1.4220 30.5100 ;
      RECT 1.2880 29.4165 1.3140 30.5100 ;
      RECT 1.1800 29.4165 1.2060 30.5100 ;
      RECT 1.0720 29.4165 1.0980 30.5100 ;
      RECT 0.9640 29.4165 0.9900 30.5100 ;
      RECT 0.8560 29.4165 0.8820 30.5100 ;
      RECT 0.7480 29.4165 0.7740 30.5100 ;
      RECT 0.6400 29.4165 0.6660 30.5100 ;
      RECT 0.5320 29.4165 0.5580 30.5100 ;
      RECT 0.4240 29.4165 0.4500 30.5100 ;
      RECT 0.3160 29.4165 0.3420 30.5100 ;
      RECT 0.2080 29.4165 0.2340 30.5100 ;
      RECT 0.0050 29.4165 0.0900 30.5100 ;
      RECT 8.6410 30.4965 8.7690 31.5900 ;
      RECT 8.6270 31.1620 8.7690 31.4845 ;
      RECT 8.4790 30.8890 8.5410 31.5900 ;
      RECT 8.4650 31.1985 8.5410 31.3520 ;
      RECT 8.4790 30.4965 8.5050 31.5900 ;
      RECT 8.4790 30.6175 8.5190 30.8570 ;
      RECT 8.4790 30.4965 8.5410 30.5855 ;
      RECT 8.1820 30.9470 8.3880 31.5900 ;
      RECT 8.3620 30.4965 8.3880 31.5900 ;
      RECT 8.1820 31.2240 8.4020 31.4820 ;
      RECT 8.1820 30.4965 8.2800 31.5900 ;
      RECT 7.7650 30.4965 7.8480 31.5900 ;
      RECT 7.7650 30.5850 7.8620 31.5205 ;
      RECT 16.4440 30.4965 16.5290 31.5900 ;
      RECT 16.3000 30.4965 16.3260 31.5900 ;
      RECT 16.1920 30.4965 16.2180 31.5900 ;
      RECT 16.0840 30.4965 16.1100 31.5900 ;
      RECT 15.9760 30.4965 16.0020 31.5900 ;
      RECT 15.8680 30.4965 15.8940 31.5900 ;
      RECT 15.7600 30.4965 15.7860 31.5900 ;
      RECT 15.6520 30.4965 15.6780 31.5900 ;
      RECT 15.5440 30.4965 15.5700 31.5900 ;
      RECT 15.4360 30.4965 15.4620 31.5900 ;
      RECT 15.3280 30.4965 15.3540 31.5900 ;
      RECT 15.2200 30.4965 15.2460 31.5900 ;
      RECT 15.1120 30.4965 15.1380 31.5900 ;
      RECT 15.0040 30.4965 15.0300 31.5900 ;
      RECT 14.8960 30.4965 14.9220 31.5900 ;
      RECT 14.7880 30.4965 14.8140 31.5900 ;
      RECT 14.6800 30.4965 14.7060 31.5900 ;
      RECT 14.5720 30.4965 14.5980 31.5900 ;
      RECT 14.4640 30.4965 14.4900 31.5900 ;
      RECT 14.3560 30.4965 14.3820 31.5900 ;
      RECT 14.2480 30.4965 14.2740 31.5900 ;
      RECT 14.1400 30.4965 14.1660 31.5900 ;
      RECT 14.0320 30.4965 14.0580 31.5900 ;
      RECT 13.9240 30.4965 13.9500 31.5900 ;
      RECT 13.8160 30.4965 13.8420 31.5900 ;
      RECT 13.7080 30.4965 13.7340 31.5900 ;
      RECT 13.6000 30.4965 13.6260 31.5900 ;
      RECT 13.4920 30.4965 13.5180 31.5900 ;
      RECT 13.3840 30.4965 13.4100 31.5900 ;
      RECT 13.2760 30.4965 13.3020 31.5900 ;
      RECT 13.1680 30.4965 13.1940 31.5900 ;
      RECT 13.0600 30.4965 13.0860 31.5900 ;
      RECT 12.9520 30.4965 12.9780 31.5900 ;
      RECT 12.8440 30.4965 12.8700 31.5900 ;
      RECT 12.7360 30.4965 12.7620 31.5900 ;
      RECT 12.6280 30.4965 12.6540 31.5900 ;
      RECT 12.5200 30.4965 12.5460 31.5900 ;
      RECT 12.4120 30.4965 12.4380 31.5900 ;
      RECT 12.3040 30.4965 12.3300 31.5900 ;
      RECT 12.1960 30.4965 12.2220 31.5900 ;
      RECT 12.0880 30.4965 12.1140 31.5900 ;
      RECT 11.9800 30.4965 12.0060 31.5900 ;
      RECT 11.8720 30.4965 11.8980 31.5900 ;
      RECT 11.7640 30.4965 11.7900 31.5900 ;
      RECT 11.6560 30.4965 11.6820 31.5900 ;
      RECT 11.5480 30.4965 11.5740 31.5900 ;
      RECT 11.4400 30.4965 11.4660 31.5900 ;
      RECT 11.3320 30.4965 11.3580 31.5900 ;
      RECT 11.2240 30.4965 11.2500 31.5900 ;
      RECT 11.1160 30.4965 11.1420 31.5900 ;
      RECT 11.0080 30.4965 11.0340 31.5900 ;
      RECT 10.9000 30.4965 10.9260 31.5900 ;
      RECT 10.7920 30.4965 10.8180 31.5900 ;
      RECT 10.6840 30.4965 10.7100 31.5900 ;
      RECT 10.5760 30.4965 10.6020 31.5900 ;
      RECT 10.4680 30.4965 10.4940 31.5900 ;
      RECT 10.3600 30.4965 10.3860 31.5900 ;
      RECT 10.2520 30.4965 10.2780 31.5900 ;
      RECT 10.1440 30.4965 10.1700 31.5900 ;
      RECT 10.0360 30.4965 10.0620 31.5900 ;
      RECT 9.9280 30.4965 9.9540 31.5900 ;
      RECT 9.8200 30.4965 9.8460 31.5900 ;
      RECT 9.7120 30.4965 9.7380 31.5900 ;
      RECT 9.6040 30.4965 9.6300 31.5900 ;
      RECT 9.4960 30.4965 9.5220 31.5900 ;
      RECT 9.3880 30.4965 9.4140 31.5900 ;
      RECT 9.1750 30.4965 9.2520 31.5900 ;
      RECT 7.2820 30.4965 7.3590 31.5900 ;
      RECT 7.1200 30.4965 7.1460 31.5900 ;
      RECT 7.0120 30.4965 7.0380 31.5900 ;
      RECT 6.9040 30.4965 6.9300 31.5900 ;
      RECT 6.7960 30.4965 6.8220 31.5900 ;
      RECT 6.6880 30.4965 6.7140 31.5900 ;
      RECT 6.5800 30.4965 6.6060 31.5900 ;
      RECT 6.4720 30.4965 6.4980 31.5900 ;
      RECT 6.3640 30.4965 6.3900 31.5900 ;
      RECT 6.2560 30.4965 6.2820 31.5900 ;
      RECT 6.1480 30.4965 6.1740 31.5900 ;
      RECT 6.0400 30.4965 6.0660 31.5900 ;
      RECT 5.9320 30.4965 5.9580 31.5900 ;
      RECT 5.8240 30.4965 5.8500 31.5900 ;
      RECT 5.7160 30.4965 5.7420 31.5900 ;
      RECT 5.6080 30.4965 5.6340 31.5900 ;
      RECT 5.5000 30.4965 5.5260 31.5900 ;
      RECT 5.3920 30.4965 5.4180 31.5900 ;
      RECT 5.2840 30.4965 5.3100 31.5900 ;
      RECT 5.1760 30.4965 5.2020 31.5900 ;
      RECT 5.0680 30.4965 5.0940 31.5900 ;
      RECT 4.9600 30.4965 4.9860 31.5900 ;
      RECT 4.8520 30.4965 4.8780 31.5900 ;
      RECT 4.7440 30.4965 4.7700 31.5900 ;
      RECT 4.6360 30.4965 4.6620 31.5900 ;
      RECT 4.5280 30.4965 4.5540 31.5900 ;
      RECT 4.4200 30.4965 4.4460 31.5900 ;
      RECT 4.3120 30.4965 4.3380 31.5900 ;
      RECT 4.2040 30.4965 4.2300 31.5900 ;
      RECT 4.0960 30.4965 4.1220 31.5900 ;
      RECT 3.9880 30.4965 4.0140 31.5900 ;
      RECT 3.8800 30.4965 3.9060 31.5900 ;
      RECT 3.7720 30.4965 3.7980 31.5900 ;
      RECT 3.6640 30.4965 3.6900 31.5900 ;
      RECT 3.5560 30.4965 3.5820 31.5900 ;
      RECT 3.4480 30.4965 3.4740 31.5900 ;
      RECT 3.3400 30.4965 3.3660 31.5900 ;
      RECT 3.2320 30.4965 3.2580 31.5900 ;
      RECT 3.1240 30.4965 3.1500 31.5900 ;
      RECT 3.0160 30.4965 3.0420 31.5900 ;
      RECT 2.9080 30.4965 2.9340 31.5900 ;
      RECT 2.8000 30.4965 2.8260 31.5900 ;
      RECT 2.6920 30.4965 2.7180 31.5900 ;
      RECT 2.5840 30.4965 2.6100 31.5900 ;
      RECT 2.4760 30.4965 2.5020 31.5900 ;
      RECT 2.3680 30.4965 2.3940 31.5900 ;
      RECT 2.2600 30.4965 2.2860 31.5900 ;
      RECT 2.1520 30.4965 2.1780 31.5900 ;
      RECT 2.0440 30.4965 2.0700 31.5900 ;
      RECT 1.9360 30.4965 1.9620 31.5900 ;
      RECT 1.8280 30.4965 1.8540 31.5900 ;
      RECT 1.7200 30.4965 1.7460 31.5900 ;
      RECT 1.6120 30.4965 1.6380 31.5900 ;
      RECT 1.5040 30.4965 1.5300 31.5900 ;
      RECT 1.3960 30.4965 1.4220 31.5900 ;
      RECT 1.2880 30.4965 1.3140 31.5900 ;
      RECT 1.1800 30.4965 1.2060 31.5900 ;
      RECT 1.0720 30.4965 1.0980 31.5900 ;
      RECT 0.9640 30.4965 0.9900 31.5900 ;
      RECT 0.8560 30.4965 0.8820 31.5900 ;
      RECT 0.7480 30.4965 0.7740 31.5900 ;
      RECT 0.6400 30.4965 0.6660 31.5900 ;
      RECT 0.5320 30.4965 0.5580 31.5900 ;
      RECT 0.4240 30.4965 0.4500 31.5900 ;
      RECT 0.3160 30.4965 0.3420 31.5900 ;
      RECT 0.2080 30.4965 0.2340 31.5900 ;
      RECT 0.0050 30.4965 0.0900 31.5900 ;
      RECT 8.6410 31.5765 8.7690 32.6700 ;
      RECT 8.6270 32.2420 8.7690 32.5645 ;
      RECT 8.4790 31.9690 8.5410 32.6700 ;
      RECT 8.4650 32.2785 8.5410 32.4320 ;
      RECT 8.4790 31.5765 8.5050 32.6700 ;
      RECT 8.4790 31.6975 8.5190 31.9370 ;
      RECT 8.4790 31.5765 8.5410 31.6655 ;
      RECT 8.1820 32.0270 8.3880 32.6700 ;
      RECT 8.3620 31.5765 8.3880 32.6700 ;
      RECT 8.1820 32.3040 8.4020 32.5620 ;
      RECT 8.1820 31.5765 8.2800 32.6700 ;
      RECT 7.7650 31.5765 7.8480 32.6700 ;
      RECT 7.7650 31.6650 7.8620 32.6005 ;
      RECT 16.4440 31.5765 16.5290 32.6700 ;
      RECT 16.3000 31.5765 16.3260 32.6700 ;
      RECT 16.1920 31.5765 16.2180 32.6700 ;
      RECT 16.0840 31.5765 16.1100 32.6700 ;
      RECT 15.9760 31.5765 16.0020 32.6700 ;
      RECT 15.8680 31.5765 15.8940 32.6700 ;
      RECT 15.7600 31.5765 15.7860 32.6700 ;
      RECT 15.6520 31.5765 15.6780 32.6700 ;
      RECT 15.5440 31.5765 15.5700 32.6700 ;
      RECT 15.4360 31.5765 15.4620 32.6700 ;
      RECT 15.3280 31.5765 15.3540 32.6700 ;
      RECT 15.2200 31.5765 15.2460 32.6700 ;
      RECT 15.1120 31.5765 15.1380 32.6700 ;
      RECT 15.0040 31.5765 15.0300 32.6700 ;
      RECT 14.8960 31.5765 14.9220 32.6700 ;
      RECT 14.7880 31.5765 14.8140 32.6700 ;
      RECT 14.6800 31.5765 14.7060 32.6700 ;
      RECT 14.5720 31.5765 14.5980 32.6700 ;
      RECT 14.4640 31.5765 14.4900 32.6700 ;
      RECT 14.3560 31.5765 14.3820 32.6700 ;
      RECT 14.2480 31.5765 14.2740 32.6700 ;
      RECT 14.1400 31.5765 14.1660 32.6700 ;
      RECT 14.0320 31.5765 14.0580 32.6700 ;
      RECT 13.9240 31.5765 13.9500 32.6700 ;
      RECT 13.8160 31.5765 13.8420 32.6700 ;
      RECT 13.7080 31.5765 13.7340 32.6700 ;
      RECT 13.6000 31.5765 13.6260 32.6700 ;
      RECT 13.4920 31.5765 13.5180 32.6700 ;
      RECT 13.3840 31.5765 13.4100 32.6700 ;
      RECT 13.2760 31.5765 13.3020 32.6700 ;
      RECT 13.1680 31.5765 13.1940 32.6700 ;
      RECT 13.0600 31.5765 13.0860 32.6700 ;
      RECT 12.9520 31.5765 12.9780 32.6700 ;
      RECT 12.8440 31.5765 12.8700 32.6700 ;
      RECT 12.7360 31.5765 12.7620 32.6700 ;
      RECT 12.6280 31.5765 12.6540 32.6700 ;
      RECT 12.5200 31.5765 12.5460 32.6700 ;
      RECT 12.4120 31.5765 12.4380 32.6700 ;
      RECT 12.3040 31.5765 12.3300 32.6700 ;
      RECT 12.1960 31.5765 12.2220 32.6700 ;
      RECT 12.0880 31.5765 12.1140 32.6700 ;
      RECT 11.9800 31.5765 12.0060 32.6700 ;
      RECT 11.8720 31.5765 11.8980 32.6700 ;
      RECT 11.7640 31.5765 11.7900 32.6700 ;
      RECT 11.6560 31.5765 11.6820 32.6700 ;
      RECT 11.5480 31.5765 11.5740 32.6700 ;
      RECT 11.4400 31.5765 11.4660 32.6700 ;
      RECT 11.3320 31.5765 11.3580 32.6700 ;
      RECT 11.2240 31.5765 11.2500 32.6700 ;
      RECT 11.1160 31.5765 11.1420 32.6700 ;
      RECT 11.0080 31.5765 11.0340 32.6700 ;
      RECT 10.9000 31.5765 10.9260 32.6700 ;
      RECT 10.7920 31.5765 10.8180 32.6700 ;
      RECT 10.6840 31.5765 10.7100 32.6700 ;
      RECT 10.5760 31.5765 10.6020 32.6700 ;
      RECT 10.4680 31.5765 10.4940 32.6700 ;
      RECT 10.3600 31.5765 10.3860 32.6700 ;
      RECT 10.2520 31.5765 10.2780 32.6700 ;
      RECT 10.1440 31.5765 10.1700 32.6700 ;
      RECT 10.0360 31.5765 10.0620 32.6700 ;
      RECT 9.9280 31.5765 9.9540 32.6700 ;
      RECT 9.8200 31.5765 9.8460 32.6700 ;
      RECT 9.7120 31.5765 9.7380 32.6700 ;
      RECT 9.6040 31.5765 9.6300 32.6700 ;
      RECT 9.4960 31.5765 9.5220 32.6700 ;
      RECT 9.3880 31.5765 9.4140 32.6700 ;
      RECT 9.1750 31.5765 9.2520 32.6700 ;
      RECT 7.2820 31.5765 7.3590 32.6700 ;
      RECT 7.1200 31.5765 7.1460 32.6700 ;
      RECT 7.0120 31.5765 7.0380 32.6700 ;
      RECT 6.9040 31.5765 6.9300 32.6700 ;
      RECT 6.7960 31.5765 6.8220 32.6700 ;
      RECT 6.6880 31.5765 6.7140 32.6700 ;
      RECT 6.5800 31.5765 6.6060 32.6700 ;
      RECT 6.4720 31.5765 6.4980 32.6700 ;
      RECT 6.3640 31.5765 6.3900 32.6700 ;
      RECT 6.2560 31.5765 6.2820 32.6700 ;
      RECT 6.1480 31.5765 6.1740 32.6700 ;
      RECT 6.0400 31.5765 6.0660 32.6700 ;
      RECT 5.9320 31.5765 5.9580 32.6700 ;
      RECT 5.8240 31.5765 5.8500 32.6700 ;
      RECT 5.7160 31.5765 5.7420 32.6700 ;
      RECT 5.6080 31.5765 5.6340 32.6700 ;
      RECT 5.5000 31.5765 5.5260 32.6700 ;
      RECT 5.3920 31.5765 5.4180 32.6700 ;
      RECT 5.2840 31.5765 5.3100 32.6700 ;
      RECT 5.1760 31.5765 5.2020 32.6700 ;
      RECT 5.0680 31.5765 5.0940 32.6700 ;
      RECT 4.9600 31.5765 4.9860 32.6700 ;
      RECT 4.8520 31.5765 4.8780 32.6700 ;
      RECT 4.7440 31.5765 4.7700 32.6700 ;
      RECT 4.6360 31.5765 4.6620 32.6700 ;
      RECT 4.5280 31.5765 4.5540 32.6700 ;
      RECT 4.4200 31.5765 4.4460 32.6700 ;
      RECT 4.3120 31.5765 4.3380 32.6700 ;
      RECT 4.2040 31.5765 4.2300 32.6700 ;
      RECT 4.0960 31.5765 4.1220 32.6700 ;
      RECT 3.9880 31.5765 4.0140 32.6700 ;
      RECT 3.8800 31.5765 3.9060 32.6700 ;
      RECT 3.7720 31.5765 3.7980 32.6700 ;
      RECT 3.6640 31.5765 3.6900 32.6700 ;
      RECT 3.5560 31.5765 3.5820 32.6700 ;
      RECT 3.4480 31.5765 3.4740 32.6700 ;
      RECT 3.3400 31.5765 3.3660 32.6700 ;
      RECT 3.2320 31.5765 3.2580 32.6700 ;
      RECT 3.1240 31.5765 3.1500 32.6700 ;
      RECT 3.0160 31.5765 3.0420 32.6700 ;
      RECT 2.9080 31.5765 2.9340 32.6700 ;
      RECT 2.8000 31.5765 2.8260 32.6700 ;
      RECT 2.6920 31.5765 2.7180 32.6700 ;
      RECT 2.5840 31.5765 2.6100 32.6700 ;
      RECT 2.4760 31.5765 2.5020 32.6700 ;
      RECT 2.3680 31.5765 2.3940 32.6700 ;
      RECT 2.2600 31.5765 2.2860 32.6700 ;
      RECT 2.1520 31.5765 2.1780 32.6700 ;
      RECT 2.0440 31.5765 2.0700 32.6700 ;
      RECT 1.9360 31.5765 1.9620 32.6700 ;
      RECT 1.8280 31.5765 1.8540 32.6700 ;
      RECT 1.7200 31.5765 1.7460 32.6700 ;
      RECT 1.6120 31.5765 1.6380 32.6700 ;
      RECT 1.5040 31.5765 1.5300 32.6700 ;
      RECT 1.3960 31.5765 1.4220 32.6700 ;
      RECT 1.2880 31.5765 1.3140 32.6700 ;
      RECT 1.1800 31.5765 1.2060 32.6700 ;
      RECT 1.0720 31.5765 1.0980 32.6700 ;
      RECT 0.9640 31.5765 0.9900 32.6700 ;
      RECT 0.8560 31.5765 0.8820 32.6700 ;
      RECT 0.7480 31.5765 0.7740 32.6700 ;
      RECT 0.6400 31.5765 0.6660 32.6700 ;
      RECT 0.5320 31.5765 0.5580 32.6700 ;
      RECT 0.4240 31.5765 0.4500 32.6700 ;
      RECT 0.3160 31.5765 0.3420 32.6700 ;
      RECT 0.2080 31.5765 0.2340 32.6700 ;
      RECT 0.0050 31.5765 0.0900 32.6700 ;
      RECT 8.6410 32.6565 8.7690 33.7500 ;
      RECT 8.6270 33.3220 8.7690 33.6445 ;
      RECT 8.4790 33.0490 8.5410 33.7500 ;
      RECT 8.4650 33.3585 8.5410 33.5120 ;
      RECT 8.4790 32.6565 8.5050 33.7500 ;
      RECT 8.4790 32.7775 8.5190 33.0170 ;
      RECT 8.4790 32.6565 8.5410 32.7455 ;
      RECT 8.1820 33.1070 8.3880 33.7500 ;
      RECT 8.3620 32.6565 8.3880 33.7500 ;
      RECT 8.1820 33.3840 8.4020 33.6420 ;
      RECT 8.1820 32.6565 8.2800 33.7500 ;
      RECT 7.7650 32.6565 7.8480 33.7500 ;
      RECT 7.7650 32.7450 7.8620 33.6805 ;
      RECT 16.4440 32.6565 16.5290 33.7500 ;
      RECT 16.3000 32.6565 16.3260 33.7500 ;
      RECT 16.1920 32.6565 16.2180 33.7500 ;
      RECT 16.0840 32.6565 16.1100 33.7500 ;
      RECT 15.9760 32.6565 16.0020 33.7500 ;
      RECT 15.8680 32.6565 15.8940 33.7500 ;
      RECT 15.7600 32.6565 15.7860 33.7500 ;
      RECT 15.6520 32.6565 15.6780 33.7500 ;
      RECT 15.5440 32.6565 15.5700 33.7500 ;
      RECT 15.4360 32.6565 15.4620 33.7500 ;
      RECT 15.3280 32.6565 15.3540 33.7500 ;
      RECT 15.2200 32.6565 15.2460 33.7500 ;
      RECT 15.1120 32.6565 15.1380 33.7500 ;
      RECT 15.0040 32.6565 15.0300 33.7500 ;
      RECT 14.8960 32.6565 14.9220 33.7500 ;
      RECT 14.7880 32.6565 14.8140 33.7500 ;
      RECT 14.6800 32.6565 14.7060 33.7500 ;
      RECT 14.5720 32.6565 14.5980 33.7500 ;
      RECT 14.4640 32.6565 14.4900 33.7500 ;
      RECT 14.3560 32.6565 14.3820 33.7500 ;
      RECT 14.2480 32.6565 14.2740 33.7500 ;
      RECT 14.1400 32.6565 14.1660 33.7500 ;
      RECT 14.0320 32.6565 14.0580 33.7500 ;
      RECT 13.9240 32.6565 13.9500 33.7500 ;
      RECT 13.8160 32.6565 13.8420 33.7500 ;
      RECT 13.7080 32.6565 13.7340 33.7500 ;
      RECT 13.6000 32.6565 13.6260 33.7500 ;
      RECT 13.4920 32.6565 13.5180 33.7500 ;
      RECT 13.3840 32.6565 13.4100 33.7500 ;
      RECT 13.2760 32.6565 13.3020 33.7500 ;
      RECT 13.1680 32.6565 13.1940 33.7500 ;
      RECT 13.0600 32.6565 13.0860 33.7500 ;
      RECT 12.9520 32.6565 12.9780 33.7500 ;
      RECT 12.8440 32.6565 12.8700 33.7500 ;
      RECT 12.7360 32.6565 12.7620 33.7500 ;
      RECT 12.6280 32.6565 12.6540 33.7500 ;
      RECT 12.5200 32.6565 12.5460 33.7500 ;
      RECT 12.4120 32.6565 12.4380 33.7500 ;
      RECT 12.3040 32.6565 12.3300 33.7500 ;
      RECT 12.1960 32.6565 12.2220 33.7500 ;
      RECT 12.0880 32.6565 12.1140 33.7500 ;
      RECT 11.9800 32.6565 12.0060 33.7500 ;
      RECT 11.8720 32.6565 11.8980 33.7500 ;
      RECT 11.7640 32.6565 11.7900 33.7500 ;
      RECT 11.6560 32.6565 11.6820 33.7500 ;
      RECT 11.5480 32.6565 11.5740 33.7500 ;
      RECT 11.4400 32.6565 11.4660 33.7500 ;
      RECT 11.3320 32.6565 11.3580 33.7500 ;
      RECT 11.2240 32.6565 11.2500 33.7500 ;
      RECT 11.1160 32.6565 11.1420 33.7500 ;
      RECT 11.0080 32.6565 11.0340 33.7500 ;
      RECT 10.9000 32.6565 10.9260 33.7500 ;
      RECT 10.7920 32.6565 10.8180 33.7500 ;
      RECT 10.6840 32.6565 10.7100 33.7500 ;
      RECT 10.5760 32.6565 10.6020 33.7500 ;
      RECT 10.4680 32.6565 10.4940 33.7500 ;
      RECT 10.3600 32.6565 10.3860 33.7500 ;
      RECT 10.2520 32.6565 10.2780 33.7500 ;
      RECT 10.1440 32.6565 10.1700 33.7500 ;
      RECT 10.0360 32.6565 10.0620 33.7500 ;
      RECT 9.9280 32.6565 9.9540 33.7500 ;
      RECT 9.8200 32.6565 9.8460 33.7500 ;
      RECT 9.7120 32.6565 9.7380 33.7500 ;
      RECT 9.6040 32.6565 9.6300 33.7500 ;
      RECT 9.4960 32.6565 9.5220 33.7500 ;
      RECT 9.3880 32.6565 9.4140 33.7500 ;
      RECT 9.1750 32.6565 9.2520 33.7500 ;
      RECT 7.2820 32.6565 7.3590 33.7500 ;
      RECT 7.1200 32.6565 7.1460 33.7500 ;
      RECT 7.0120 32.6565 7.0380 33.7500 ;
      RECT 6.9040 32.6565 6.9300 33.7500 ;
      RECT 6.7960 32.6565 6.8220 33.7500 ;
      RECT 6.6880 32.6565 6.7140 33.7500 ;
      RECT 6.5800 32.6565 6.6060 33.7500 ;
      RECT 6.4720 32.6565 6.4980 33.7500 ;
      RECT 6.3640 32.6565 6.3900 33.7500 ;
      RECT 6.2560 32.6565 6.2820 33.7500 ;
      RECT 6.1480 32.6565 6.1740 33.7500 ;
      RECT 6.0400 32.6565 6.0660 33.7500 ;
      RECT 5.9320 32.6565 5.9580 33.7500 ;
      RECT 5.8240 32.6565 5.8500 33.7500 ;
      RECT 5.7160 32.6565 5.7420 33.7500 ;
      RECT 5.6080 32.6565 5.6340 33.7500 ;
      RECT 5.5000 32.6565 5.5260 33.7500 ;
      RECT 5.3920 32.6565 5.4180 33.7500 ;
      RECT 5.2840 32.6565 5.3100 33.7500 ;
      RECT 5.1760 32.6565 5.2020 33.7500 ;
      RECT 5.0680 32.6565 5.0940 33.7500 ;
      RECT 4.9600 32.6565 4.9860 33.7500 ;
      RECT 4.8520 32.6565 4.8780 33.7500 ;
      RECT 4.7440 32.6565 4.7700 33.7500 ;
      RECT 4.6360 32.6565 4.6620 33.7500 ;
      RECT 4.5280 32.6565 4.5540 33.7500 ;
      RECT 4.4200 32.6565 4.4460 33.7500 ;
      RECT 4.3120 32.6565 4.3380 33.7500 ;
      RECT 4.2040 32.6565 4.2300 33.7500 ;
      RECT 4.0960 32.6565 4.1220 33.7500 ;
      RECT 3.9880 32.6565 4.0140 33.7500 ;
      RECT 3.8800 32.6565 3.9060 33.7500 ;
      RECT 3.7720 32.6565 3.7980 33.7500 ;
      RECT 3.6640 32.6565 3.6900 33.7500 ;
      RECT 3.5560 32.6565 3.5820 33.7500 ;
      RECT 3.4480 32.6565 3.4740 33.7500 ;
      RECT 3.3400 32.6565 3.3660 33.7500 ;
      RECT 3.2320 32.6565 3.2580 33.7500 ;
      RECT 3.1240 32.6565 3.1500 33.7500 ;
      RECT 3.0160 32.6565 3.0420 33.7500 ;
      RECT 2.9080 32.6565 2.9340 33.7500 ;
      RECT 2.8000 32.6565 2.8260 33.7500 ;
      RECT 2.6920 32.6565 2.7180 33.7500 ;
      RECT 2.5840 32.6565 2.6100 33.7500 ;
      RECT 2.4760 32.6565 2.5020 33.7500 ;
      RECT 2.3680 32.6565 2.3940 33.7500 ;
      RECT 2.2600 32.6565 2.2860 33.7500 ;
      RECT 2.1520 32.6565 2.1780 33.7500 ;
      RECT 2.0440 32.6565 2.0700 33.7500 ;
      RECT 1.9360 32.6565 1.9620 33.7500 ;
      RECT 1.8280 32.6565 1.8540 33.7500 ;
      RECT 1.7200 32.6565 1.7460 33.7500 ;
      RECT 1.6120 32.6565 1.6380 33.7500 ;
      RECT 1.5040 32.6565 1.5300 33.7500 ;
      RECT 1.3960 32.6565 1.4220 33.7500 ;
      RECT 1.2880 32.6565 1.3140 33.7500 ;
      RECT 1.1800 32.6565 1.2060 33.7500 ;
      RECT 1.0720 32.6565 1.0980 33.7500 ;
      RECT 0.9640 32.6565 0.9900 33.7500 ;
      RECT 0.8560 32.6565 0.8820 33.7500 ;
      RECT 0.7480 32.6565 0.7740 33.7500 ;
      RECT 0.6400 32.6565 0.6660 33.7500 ;
      RECT 0.5320 32.6565 0.5580 33.7500 ;
      RECT 0.4240 32.6565 0.4500 33.7500 ;
      RECT 0.3160 32.6565 0.3420 33.7500 ;
      RECT 0.2080 32.6565 0.2340 33.7500 ;
      RECT 0.0050 32.6565 0.0900 33.7500 ;
      RECT 8.6410 33.7365 8.7690 34.8300 ;
      RECT 8.6270 34.4020 8.7690 34.7245 ;
      RECT 8.4790 34.1290 8.5410 34.8300 ;
      RECT 8.4650 34.4385 8.5410 34.5920 ;
      RECT 8.4790 33.7365 8.5050 34.8300 ;
      RECT 8.4790 33.8575 8.5190 34.0970 ;
      RECT 8.4790 33.7365 8.5410 33.8255 ;
      RECT 8.1820 34.1870 8.3880 34.8300 ;
      RECT 8.3620 33.7365 8.3880 34.8300 ;
      RECT 8.1820 34.4640 8.4020 34.7220 ;
      RECT 8.1820 33.7365 8.2800 34.8300 ;
      RECT 7.7650 33.7365 7.8480 34.8300 ;
      RECT 7.7650 33.8250 7.8620 34.7605 ;
      RECT 16.4440 33.7365 16.5290 34.8300 ;
      RECT 16.3000 33.7365 16.3260 34.8300 ;
      RECT 16.1920 33.7365 16.2180 34.8300 ;
      RECT 16.0840 33.7365 16.1100 34.8300 ;
      RECT 15.9760 33.7365 16.0020 34.8300 ;
      RECT 15.8680 33.7365 15.8940 34.8300 ;
      RECT 15.7600 33.7365 15.7860 34.8300 ;
      RECT 15.6520 33.7365 15.6780 34.8300 ;
      RECT 15.5440 33.7365 15.5700 34.8300 ;
      RECT 15.4360 33.7365 15.4620 34.8300 ;
      RECT 15.3280 33.7365 15.3540 34.8300 ;
      RECT 15.2200 33.7365 15.2460 34.8300 ;
      RECT 15.1120 33.7365 15.1380 34.8300 ;
      RECT 15.0040 33.7365 15.0300 34.8300 ;
      RECT 14.8960 33.7365 14.9220 34.8300 ;
      RECT 14.7880 33.7365 14.8140 34.8300 ;
      RECT 14.6800 33.7365 14.7060 34.8300 ;
      RECT 14.5720 33.7365 14.5980 34.8300 ;
      RECT 14.4640 33.7365 14.4900 34.8300 ;
      RECT 14.3560 33.7365 14.3820 34.8300 ;
      RECT 14.2480 33.7365 14.2740 34.8300 ;
      RECT 14.1400 33.7365 14.1660 34.8300 ;
      RECT 14.0320 33.7365 14.0580 34.8300 ;
      RECT 13.9240 33.7365 13.9500 34.8300 ;
      RECT 13.8160 33.7365 13.8420 34.8300 ;
      RECT 13.7080 33.7365 13.7340 34.8300 ;
      RECT 13.6000 33.7365 13.6260 34.8300 ;
      RECT 13.4920 33.7365 13.5180 34.8300 ;
      RECT 13.3840 33.7365 13.4100 34.8300 ;
      RECT 13.2760 33.7365 13.3020 34.8300 ;
      RECT 13.1680 33.7365 13.1940 34.8300 ;
      RECT 13.0600 33.7365 13.0860 34.8300 ;
      RECT 12.9520 33.7365 12.9780 34.8300 ;
      RECT 12.8440 33.7365 12.8700 34.8300 ;
      RECT 12.7360 33.7365 12.7620 34.8300 ;
      RECT 12.6280 33.7365 12.6540 34.8300 ;
      RECT 12.5200 33.7365 12.5460 34.8300 ;
      RECT 12.4120 33.7365 12.4380 34.8300 ;
      RECT 12.3040 33.7365 12.3300 34.8300 ;
      RECT 12.1960 33.7365 12.2220 34.8300 ;
      RECT 12.0880 33.7365 12.1140 34.8300 ;
      RECT 11.9800 33.7365 12.0060 34.8300 ;
      RECT 11.8720 33.7365 11.8980 34.8300 ;
      RECT 11.7640 33.7365 11.7900 34.8300 ;
      RECT 11.6560 33.7365 11.6820 34.8300 ;
      RECT 11.5480 33.7365 11.5740 34.8300 ;
      RECT 11.4400 33.7365 11.4660 34.8300 ;
      RECT 11.3320 33.7365 11.3580 34.8300 ;
      RECT 11.2240 33.7365 11.2500 34.8300 ;
      RECT 11.1160 33.7365 11.1420 34.8300 ;
      RECT 11.0080 33.7365 11.0340 34.8300 ;
      RECT 10.9000 33.7365 10.9260 34.8300 ;
      RECT 10.7920 33.7365 10.8180 34.8300 ;
      RECT 10.6840 33.7365 10.7100 34.8300 ;
      RECT 10.5760 33.7365 10.6020 34.8300 ;
      RECT 10.4680 33.7365 10.4940 34.8300 ;
      RECT 10.3600 33.7365 10.3860 34.8300 ;
      RECT 10.2520 33.7365 10.2780 34.8300 ;
      RECT 10.1440 33.7365 10.1700 34.8300 ;
      RECT 10.0360 33.7365 10.0620 34.8300 ;
      RECT 9.9280 33.7365 9.9540 34.8300 ;
      RECT 9.8200 33.7365 9.8460 34.8300 ;
      RECT 9.7120 33.7365 9.7380 34.8300 ;
      RECT 9.6040 33.7365 9.6300 34.8300 ;
      RECT 9.4960 33.7365 9.5220 34.8300 ;
      RECT 9.3880 33.7365 9.4140 34.8300 ;
      RECT 9.1750 33.7365 9.2520 34.8300 ;
      RECT 7.2820 33.7365 7.3590 34.8300 ;
      RECT 7.1200 33.7365 7.1460 34.8300 ;
      RECT 7.0120 33.7365 7.0380 34.8300 ;
      RECT 6.9040 33.7365 6.9300 34.8300 ;
      RECT 6.7960 33.7365 6.8220 34.8300 ;
      RECT 6.6880 33.7365 6.7140 34.8300 ;
      RECT 6.5800 33.7365 6.6060 34.8300 ;
      RECT 6.4720 33.7365 6.4980 34.8300 ;
      RECT 6.3640 33.7365 6.3900 34.8300 ;
      RECT 6.2560 33.7365 6.2820 34.8300 ;
      RECT 6.1480 33.7365 6.1740 34.8300 ;
      RECT 6.0400 33.7365 6.0660 34.8300 ;
      RECT 5.9320 33.7365 5.9580 34.8300 ;
      RECT 5.8240 33.7365 5.8500 34.8300 ;
      RECT 5.7160 33.7365 5.7420 34.8300 ;
      RECT 5.6080 33.7365 5.6340 34.8300 ;
      RECT 5.5000 33.7365 5.5260 34.8300 ;
      RECT 5.3920 33.7365 5.4180 34.8300 ;
      RECT 5.2840 33.7365 5.3100 34.8300 ;
      RECT 5.1760 33.7365 5.2020 34.8300 ;
      RECT 5.0680 33.7365 5.0940 34.8300 ;
      RECT 4.9600 33.7365 4.9860 34.8300 ;
      RECT 4.8520 33.7365 4.8780 34.8300 ;
      RECT 4.7440 33.7365 4.7700 34.8300 ;
      RECT 4.6360 33.7365 4.6620 34.8300 ;
      RECT 4.5280 33.7365 4.5540 34.8300 ;
      RECT 4.4200 33.7365 4.4460 34.8300 ;
      RECT 4.3120 33.7365 4.3380 34.8300 ;
      RECT 4.2040 33.7365 4.2300 34.8300 ;
      RECT 4.0960 33.7365 4.1220 34.8300 ;
      RECT 3.9880 33.7365 4.0140 34.8300 ;
      RECT 3.8800 33.7365 3.9060 34.8300 ;
      RECT 3.7720 33.7365 3.7980 34.8300 ;
      RECT 3.6640 33.7365 3.6900 34.8300 ;
      RECT 3.5560 33.7365 3.5820 34.8300 ;
      RECT 3.4480 33.7365 3.4740 34.8300 ;
      RECT 3.3400 33.7365 3.3660 34.8300 ;
      RECT 3.2320 33.7365 3.2580 34.8300 ;
      RECT 3.1240 33.7365 3.1500 34.8300 ;
      RECT 3.0160 33.7365 3.0420 34.8300 ;
      RECT 2.9080 33.7365 2.9340 34.8300 ;
      RECT 2.8000 33.7365 2.8260 34.8300 ;
      RECT 2.6920 33.7365 2.7180 34.8300 ;
      RECT 2.5840 33.7365 2.6100 34.8300 ;
      RECT 2.4760 33.7365 2.5020 34.8300 ;
      RECT 2.3680 33.7365 2.3940 34.8300 ;
      RECT 2.2600 33.7365 2.2860 34.8300 ;
      RECT 2.1520 33.7365 2.1780 34.8300 ;
      RECT 2.0440 33.7365 2.0700 34.8300 ;
      RECT 1.9360 33.7365 1.9620 34.8300 ;
      RECT 1.8280 33.7365 1.8540 34.8300 ;
      RECT 1.7200 33.7365 1.7460 34.8300 ;
      RECT 1.6120 33.7365 1.6380 34.8300 ;
      RECT 1.5040 33.7365 1.5300 34.8300 ;
      RECT 1.3960 33.7365 1.4220 34.8300 ;
      RECT 1.2880 33.7365 1.3140 34.8300 ;
      RECT 1.1800 33.7365 1.2060 34.8300 ;
      RECT 1.0720 33.7365 1.0980 34.8300 ;
      RECT 0.9640 33.7365 0.9900 34.8300 ;
      RECT 0.8560 33.7365 0.8820 34.8300 ;
      RECT 0.7480 33.7365 0.7740 34.8300 ;
      RECT 0.6400 33.7365 0.6660 34.8300 ;
      RECT 0.5320 33.7365 0.5580 34.8300 ;
      RECT 0.4240 33.7365 0.4500 34.8300 ;
      RECT 0.3160 33.7365 0.3420 34.8300 ;
      RECT 0.2080 33.7365 0.2340 34.8300 ;
      RECT 0.0050 33.7365 0.0900 34.8300 ;
      RECT 8.6410 34.8165 8.7690 35.9100 ;
      RECT 8.6270 35.4820 8.7690 35.8045 ;
      RECT 8.4790 35.2090 8.5410 35.9100 ;
      RECT 8.4650 35.5185 8.5410 35.6720 ;
      RECT 8.4790 34.8165 8.5050 35.9100 ;
      RECT 8.4790 34.9375 8.5190 35.1770 ;
      RECT 8.4790 34.8165 8.5410 34.9055 ;
      RECT 8.1820 35.2670 8.3880 35.9100 ;
      RECT 8.3620 34.8165 8.3880 35.9100 ;
      RECT 8.1820 35.5440 8.4020 35.8020 ;
      RECT 8.1820 34.8165 8.2800 35.9100 ;
      RECT 7.7650 34.8165 7.8480 35.9100 ;
      RECT 7.7650 34.9050 7.8620 35.8405 ;
      RECT 16.4440 34.8165 16.5290 35.9100 ;
      RECT 16.3000 34.8165 16.3260 35.9100 ;
      RECT 16.1920 34.8165 16.2180 35.9100 ;
      RECT 16.0840 34.8165 16.1100 35.9100 ;
      RECT 15.9760 34.8165 16.0020 35.9100 ;
      RECT 15.8680 34.8165 15.8940 35.9100 ;
      RECT 15.7600 34.8165 15.7860 35.9100 ;
      RECT 15.6520 34.8165 15.6780 35.9100 ;
      RECT 15.5440 34.8165 15.5700 35.9100 ;
      RECT 15.4360 34.8165 15.4620 35.9100 ;
      RECT 15.3280 34.8165 15.3540 35.9100 ;
      RECT 15.2200 34.8165 15.2460 35.9100 ;
      RECT 15.1120 34.8165 15.1380 35.9100 ;
      RECT 15.0040 34.8165 15.0300 35.9100 ;
      RECT 14.8960 34.8165 14.9220 35.9100 ;
      RECT 14.7880 34.8165 14.8140 35.9100 ;
      RECT 14.6800 34.8165 14.7060 35.9100 ;
      RECT 14.5720 34.8165 14.5980 35.9100 ;
      RECT 14.4640 34.8165 14.4900 35.9100 ;
      RECT 14.3560 34.8165 14.3820 35.9100 ;
      RECT 14.2480 34.8165 14.2740 35.9100 ;
      RECT 14.1400 34.8165 14.1660 35.9100 ;
      RECT 14.0320 34.8165 14.0580 35.9100 ;
      RECT 13.9240 34.8165 13.9500 35.9100 ;
      RECT 13.8160 34.8165 13.8420 35.9100 ;
      RECT 13.7080 34.8165 13.7340 35.9100 ;
      RECT 13.6000 34.8165 13.6260 35.9100 ;
      RECT 13.4920 34.8165 13.5180 35.9100 ;
      RECT 13.3840 34.8165 13.4100 35.9100 ;
      RECT 13.2760 34.8165 13.3020 35.9100 ;
      RECT 13.1680 34.8165 13.1940 35.9100 ;
      RECT 13.0600 34.8165 13.0860 35.9100 ;
      RECT 12.9520 34.8165 12.9780 35.9100 ;
      RECT 12.8440 34.8165 12.8700 35.9100 ;
      RECT 12.7360 34.8165 12.7620 35.9100 ;
      RECT 12.6280 34.8165 12.6540 35.9100 ;
      RECT 12.5200 34.8165 12.5460 35.9100 ;
      RECT 12.4120 34.8165 12.4380 35.9100 ;
      RECT 12.3040 34.8165 12.3300 35.9100 ;
      RECT 12.1960 34.8165 12.2220 35.9100 ;
      RECT 12.0880 34.8165 12.1140 35.9100 ;
      RECT 11.9800 34.8165 12.0060 35.9100 ;
      RECT 11.8720 34.8165 11.8980 35.9100 ;
      RECT 11.7640 34.8165 11.7900 35.9100 ;
      RECT 11.6560 34.8165 11.6820 35.9100 ;
      RECT 11.5480 34.8165 11.5740 35.9100 ;
      RECT 11.4400 34.8165 11.4660 35.9100 ;
      RECT 11.3320 34.8165 11.3580 35.9100 ;
      RECT 11.2240 34.8165 11.2500 35.9100 ;
      RECT 11.1160 34.8165 11.1420 35.9100 ;
      RECT 11.0080 34.8165 11.0340 35.9100 ;
      RECT 10.9000 34.8165 10.9260 35.9100 ;
      RECT 10.7920 34.8165 10.8180 35.9100 ;
      RECT 10.6840 34.8165 10.7100 35.9100 ;
      RECT 10.5760 34.8165 10.6020 35.9100 ;
      RECT 10.4680 34.8165 10.4940 35.9100 ;
      RECT 10.3600 34.8165 10.3860 35.9100 ;
      RECT 10.2520 34.8165 10.2780 35.9100 ;
      RECT 10.1440 34.8165 10.1700 35.9100 ;
      RECT 10.0360 34.8165 10.0620 35.9100 ;
      RECT 9.9280 34.8165 9.9540 35.9100 ;
      RECT 9.8200 34.8165 9.8460 35.9100 ;
      RECT 9.7120 34.8165 9.7380 35.9100 ;
      RECT 9.6040 34.8165 9.6300 35.9100 ;
      RECT 9.4960 34.8165 9.5220 35.9100 ;
      RECT 9.3880 34.8165 9.4140 35.9100 ;
      RECT 9.1750 34.8165 9.2520 35.9100 ;
      RECT 7.2820 34.8165 7.3590 35.9100 ;
      RECT 7.1200 34.8165 7.1460 35.9100 ;
      RECT 7.0120 34.8165 7.0380 35.9100 ;
      RECT 6.9040 34.8165 6.9300 35.9100 ;
      RECT 6.7960 34.8165 6.8220 35.9100 ;
      RECT 6.6880 34.8165 6.7140 35.9100 ;
      RECT 6.5800 34.8165 6.6060 35.9100 ;
      RECT 6.4720 34.8165 6.4980 35.9100 ;
      RECT 6.3640 34.8165 6.3900 35.9100 ;
      RECT 6.2560 34.8165 6.2820 35.9100 ;
      RECT 6.1480 34.8165 6.1740 35.9100 ;
      RECT 6.0400 34.8165 6.0660 35.9100 ;
      RECT 5.9320 34.8165 5.9580 35.9100 ;
      RECT 5.8240 34.8165 5.8500 35.9100 ;
      RECT 5.7160 34.8165 5.7420 35.9100 ;
      RECT 5.6080 34.8165 5.6340 35.9100 ;
      RECT 5.5000 34.8165 5.5260 35.9100 ;
      RECT 5.3920 34.8165 5.4180 35.9100 ;
      RECT 5.2840 34.8165 5.3100 35.9100 ;
      RECT 5.1760 34.8165 5.2020 35.9100 ;
      RECT 5.0680 34.8165 5.0940 35.9100 ;
      RECT 4.9600 34.8165 4.9860 35.9100 ;
      RECT 4.8520 34.8165 4.8780 35.9100 ;
      RECT 4.7440 34.8165 4.7700 35.9100 ;
      RECT 4.6360 34.8165 4.6620 35.9100 ;
      RECT 4.5280 34.8165 4.5540 35.9100 ;
      RECT 4.4200 34.8165 4.4460 35.9100 ;
      RECT 4.3120 34.8165 4.3380 35.9100 ;
      RECT 4.2040 34.8165 4.2300 35.9100 ;
      RECT 4.0960 34.8165 4.1220 35.9100 ;
      RECT 3.9880 34.8165 4.0140 35.9100 ;
      RECT 3.8800 34.8165 3.9060 35.9100 ;
      RECT 3.7720 34.8165 3.7980 35.9100 ;
      RECT 3.6640 34.8165 3.6900 35.9100 ;
      RECT 3.5560 34.8165 3.5820 35.9100 ;
      RECT 3.4480 34.8165 3.4740 35.9100 ;
      RECT 3.3400 34.8165 3.3660 35.9100 ;
      RECT 3.2320 34.8165 3.2580 35.9100 ;
      RECT 3.1240 34.8165 3.1500 35.9100 ;
      RECT 3.0160 34.8165 3.0420 35.9100 ;
      RECT 2.9080 34.8165 2.9340 35.9100 ;
      RECT 2.8000 34.8165 2.8260 35.9100 ;
      RECT 2.6920 34.8165 2.7180 35.9100 ;
      RECT 2.5840 34.8165 2.6100 35.9100 ;
      RECT 2.4760 34.8165 2.5020 35.9100 ;
      RECT 2.3680 34.8165 2.3940 35.9100 ;
      RECT 2.2600 34.8165 2.2860 35.9100 ;
      RECT 2.1520 34.8165 2.1780 35.9100 ;
      RECT 2.0440 34.8165 2.0700 35.9100 ;
      RECT 1.9360 34.8165 1.9620 35.9100 ;
      RECT 1.8280 34.8165 1.8540 35.9100 ;
      RECT 1.7200 34.8165 1.7460 35.9100 ;
      RECT 1.6120 34.8165 1.6380 35.9100 ;
      RECT 1.5040 34.8165 1.5300 35.9100 ;
      RECT 1.3960 34.8165 1.4220 35.9100 ;
      RECT 1.2880 34.8165 1.3140 35.9100 ;
      RECT 1.1800 34.8165 1.2060 35.9100 ;
      RECT 1.0720 34.8165 1.0980 35.9100 ;
      RECT 0.9640 34.8165 0.9900 35.9100 ;
      RECT 0.8560 34.8165 0.8820 35.9100 ;
      RECT 0.7480 34.8165 0.7740 35.9100 ;
      RECT 0.6400 34.8165 0.6660 35.9100 ;
      RECT 0.5320 34.8165 0.5580 35.9100 ;
      RECT 0.4240 34.8165 0.4500 35.9100 ;
      RECT 0.3160 34.8165 0.3420 35.9100 ;
      RECT 0.2080 34.8165 0.2340 35.9100 ;
      RECT 0.0050 34.8165 0.0900 35.9100 ;
      RECT 8.6410 35.8965 8.7690 36.9900 ;
      RECT 8.6270 36.5620 8.7690 36.8845 ;
      RECT 8.4790 36.2890 8.5410 36.9900 ;
      RECT 8.4650 36.5985 8.5410 36.7520 ;
      RECT 8.4790 35.8965 8.5050 36.9900 ;
      RECT 8.4790 36.0175 8.5190 36.2570 ;
      RECT 8.4790 35.8965 8.5410 35.9855 ;
      RECT 8.1820 36.3470 8.3880 36.9900 ;
      RECT 8.3620 35.8965 8.3880 36.9900 ;
      RECT 8.1820 36.6240 8.4020 36.8820 ;
      RECT 8.1820 35.8965 8.2800 36.9900 ;
      RECT 7.7650 35.8965 7.8480 36.9900 ;
      RECT 7.7650 35.9850 7.8620 36.9205 ;
      RECT 16.4440 35.8965 16.5290 36.9900 ;
      RECT 16.3000 35.8965 16.3260 36.9900 ;
      RECT 16.1920 35.8965 16.2180 36.9900 ;
      RECT 16.0840 35.8965 16.1100 36.9900 ;
      RECT 15.9760 35.8965 16.0020 36.9900 ;
      RECT 15.8680 35.8965 15.8940 36.9900 ;
      RECT 15.7600 35.8965 15.7860 36.9900 ;
      RECT 15.6520 35.8965 15.6780 36.9900 ;
      RECT 15.5440 35.8965 15.5700 36.9900 ;
      RECT 15.4360 35.8965 15.4620 36.9900 ;
      RECT 15.3280 35.8965 15.3540 36.9900 ;
      RECT 15.2200 35.8965 15.2460 36.9900 ;
      RECT 15.1120 35.8965 15.1380 36.9900 ;
      RECT 15.0040 35.8965 15.0300 36.9900 ;
      RECT 14.8960 35.8965 14.9220 36.9900 ;
      RECT 14.7880 35.8965 14.8140 36.9900 ;
      RECT 14.6800 35.8965 14.7060 36.9900 ;
      RECT 14.5720 35.8965 14.5980 36.9900 ;
      RECT 14.4640 35.8965 14.4900 36.9900 ;
      RECT 14.3560 35.8965 14.3820 36.9900 ;
      RECT 14.2480 35.8965 14.2740 36.9900 ;
      RECT 14.1400 35.8965 14.1660 36.9900 ;
      RECT 14.0320 35.8965 14.0580 36.9900 ;
      RECT 13.9240 35.8965 13.9500 36.9900 ;
      RECT 13.8160 35.8965 13.8420 36.9900 ;
      RECT 13.7080 35.8965 13.7340 36.9900 ;
      RECT 13.6000 35.8965 13.6260 36.9900 ;
      RECT 13.4920 35.8965 13.5180 36.9900 ;
      RECT 13.3840 35.8965 13.4100 36.9900 ;
      RECT 13.2760 35.8965 13.3020 36.9900 ;
      RECT 13.1680 35.8965 13.1940 36.9900 ;
      RECT 13.0600 35.8965 13.0860 36.9900 ;
      RECT 12.9520 35.8965 12.9780 36.9900 ;
      RECT 12.8440 35.8965 12.8700 36.9900 ;
      RECT 12.7360 35.8965 12.7620 36.9900 ;
      RECT 12.6280 35.8965 12.6540 36.9900 ;
      RECT 12.5200 35.8965 12.5460 36.9900 ;
      RECT 12.4120 35.8965 12.4380 36.9900 ;
      RECT 12.3040 35.8965 12.3300 36.9900 ;
      RECT 12.1960 35.8965 12.2220 36.9900 ;
      RECT 12.0880 35.8965 12.1140 36.9900 ;
      RECT 11.9800 35.8965 12.0060 36.9900 ;
      RECT 11.8720 35.8965 11.8980 36.9900 ;
      RECT 11.7640 35.8965 11.7900 36.9900 ;
      RECT 11.6560 35.8965 11.6820 36.9900 ;
      RECT 11.5480 35.8965 11.5740 36.9900 ;
      RECT 11.4400 35.8965 11.4660 36.9900 ;
      RECT 11.3320 35.8965 11.3580 36.9900 ;
      RECT 11.2240 35.8965 11.2500 36.9900 ;
      RECT 11.1160 35.8965 11.1420 36.9900 ;
      RECT 11.0080 35.8965 11.0340 36.9900 ;
      RECT 10.9000 35.8965 10.9260 36.9900 ;
      RECT 10.7920 35.8965 10.8180 36.9900 ;
      RECT 10.6840 35.8965 10.7100 36.9900 ;
      RECT 10.5760 35.8965 10.6020 36.9900 ;
      RECT 10.4680 35.8965 10.4940 36.9900 ;
      RECT 10.3600 35.8965 10.3860 36.9900 ;
      RECT 10.2520 35.8965 10.2780 36.9900 ;
      RECT 10.1440 35.8965 10.1700 36.9900 ;
      RECT 10.0360 35.8965 10.0620 36.9900 ;
      RECT 9.9280 35.8965 9.9540 36.9900 ;
      RECT 9.8200 35.8965 9.8460 36.9900 ;
      RECT 9.7120 35.8965 9.7380 36.9900 ;
      RECT 9.6040 35.8965 9.6300 36.9900 ;
      RECT 9.4960 35.8965 9.5220 36.9900 ;
      RECT 9.3880 35.8965 9.4140 36.9900 ;
      RECT 9.1750 35.8965 9.2520 36.9900 ;
      RECT 7.2820 35.8965 7.3590 36.9900 ;
      RECT 7.1200 35.8965 7.1460 36.9900 ;
      RECT 7.0120 35.8965 7.0380 36.9900 ;
      RECT 6.9040 35.8965 6.9300 36.9900 ;
      RECT 6.7960 35.8965 6.8220 36.9900 ;
      RECT 6.6880 35.8965 6.7140 36.9900 ;
      RECT 6.5800 35.8965 6.6060 36.9900 ;
      RECT 6.4720 35.8965 6.4980 36.9900 ;
      RECT 6.3640 35.8965 6.3900 36.9900 ;
      RECT 6.2560 35.8965 6.2820 36.9900 ;
      RECT 6.1480 35.8965 6.1740 36.9900 ;
      RECT 6.0400 35.8965 6.0660 36.9900 ;
      RECT 5.9320 35.8965 5.9580 36.9900 ;
      RECT 5.8240 35.8965 5.8500 36.9900 ;
      RECT 5.7160 35.8965 5.7420 36.9900 ;
      RECT 5.6080 35.8965 5.6340 36.9900 ;
      RECT 5.5000 35.8965 5.5260 36.9900 ;
      RECT 5.3920 35.8965 5.4180 36.9900 ;
      RECT 5.2840 35.8965 5.3100 36.9900 ;
      RECT 5.1760 35.8965 5.2020 36.9900 ;
      RECT 5.0680 35.8965 5.0940 36.9900 ;
      RECT 4.9600 35.8965 4.9860 36.9900 ;
      RECT 4.8520 35.8965 4.8780 36.9900 ;
      RECT 4.7440 35.8965 4.7700 36.9900 ;
      RECT 4.6360 35.8965 4.6620 36.9900 ;
      RECT 4.5280 35.8965 4.5540 36.9900 ;
      RECT 4.4200 35.8965 4.4460 36.9900 ;
      RECT 4.3120 35.8965 4.3380 36.9900 ;
      RECT 4.2040 35.8965 4.2300 36.9900 ;
      RECT 4.0960 35.8965 4.1220 36.9900 ;
      RECT 3.9880 35.8965 4.0140 36.9900 ;
      RECT 3.8800 35.8965 3.9060 36.9900 ;
      RECT 3.7720 35.8965 3.7980 36.9900 ;
      RECT 3.6640 35.8965 3.6900 36.9900 ;
      RECT 3.5560 35.8965 3.5820 36.9900 ;
      RECT 3.4480 35.8965 3.4740 36.9900 ;
      RECT 3.3400 35.8965 3.3660 36.9900 ;
      RECT 3.2320 35.8965 3.2580 36.9900 ;
      RECT 3.1240 35.8965 3.1500 36.9900 ;
      RECT 3.0160 35.8965 3.0420 36.9900 ;
      RECT 2.9080 35.8965 2.9340 36.9900 ;
      RECT 2.8000 35.8965 2.8260 36.9900 ;
      RECT 2.6920 35.8965 2.7180 36.9900 ;
      RECT 2.5840 35.8965 2.6100 36.9900 ;
      RECT 2.4760 35.8965 2.5020 36.9900 ;
      RECT 2.3680 35.8965 2.3940 36.9900 ;
      RECT 2.2600 35.8965 2.2860 36.9900 ;
      RECT 2.1520 35.8965 2.1780 36.9900 ;
      RECT 2.0440 35.8965 2.0700 36.9900 ;
      RECT 1.9360 35.8965 1.9620 36.9900 ;
      RECT 1.8280 35.8965 1.8540 36.9900 ;
      RECT 1.7200 35.8965 1.7460 36.9900 ;
      RECT 1.6120 35.8965 1.6380 36.9900 ;
      RECT 1.5040 35.8965 1.5300 36.9900 ;
      RECT 1.3960 35.8965 1.4220 36.9900 ;
      RECT 1.2880 35.8965 1.3140 36.9900 ;
      RECT 1.1800 35.8965 1.2060 36.9900 ;
      RECT 1.0720 35.8965 1.0980 36.9900 ;
      RECT 0.9640 35.8965 0.9900 36.9900 ;
      RECT 0.8560 35.8965 0.8820 36.9900 ;
      RECT 0.7480 35.8965 0.7740 36.9900 ;
      RECT 0.6400 35.8965 0.6660 36.9900 ;
      RECT 0.5320 35.8965 0.5580 36.9900 ;
      RECT 0.4240 35.8965 0.4500 36.9900 ;
      RECT 0.3160 35.8965 0.3420 36.9900 ;
      RECT 0.2080 35.8965 0.2340 36.9900 ;
      RECT 0.0050 35.8965 0.0900 36.9900 ;
      RECT 8.6410 36.9765 8.7690 38.0700 ;
      RECT 8.6270 37.6420 8.7690 37.9645 ;
      RECT 8.4790 37.3690 8.5410 38.0700 ;
      RECT 8.4650 37.6785 8.5410 37.8320 ;
      RECT 8.4790 36.9765 8.5050 38.0700 ;
      RECT 8.4790 37.0975 8.5190 37.3370 ;
      RECT 8.4790 36.9765 8.5410 37.0655 ;
      RECT 8.1820 37.4270 8.3880 38.0700 ;
      RECT 8.3620 36.9765 8.3880 38.0700 ;
      RECT 8.1820 37.7040 8.4020 37.9620 ;
      RECT 8.1820 36.9765 8.2800 38.0700 ;
      RECT 7.7650 36.9765 7.8480 38.0700 ;
      RECT 7.7650 37.0650 7.8620 38.0005 ;
      RECT 16.4440 36.9765 16.5290 38.0700 ;
      RECT 16.3000 36.9765 16.3260 38.0700 ;
      RECT 16.1920 36.9765 16.2180 38.0700 ;
      RECT 16.0840 36.9765 16.1100 38.0700 ;
      RECT 15.9760 36.9765 16.0020 38.0700 ;
      RECT 15.8680 36.9765 15.8940 38.0700 ;
      RECT 15.7600 36.9765 15.7860 38.0700 ;
      RECT 15.6520 36.9765 15.6780 38.0700 ;
      RECT 15.5440 36.9765 15.5700 38.0700 ;
      RECT 15.4360 36.9765 15.4620 38.0700 ;
      RECT 15.3280 36.9765 15.3540 38.0700 ;
      RECT 15.2200 36.9765 15.2460 38.0700 ;
      RECT 15.1120 36.9765 15.1380 38.0700 ;
      RECT 15.0040 36.9765 15.0300 38.0700 ;
      RECT 14.8960 36.9765 14.9220 38.0700 ;
      RECT 14.7880 36.9765 14.8140 38.0700 ;
      RECT 14.6800 36.9765 14.7060 38.0700 ;
      RECT 14.5720 36.9765 14.5980 38.0700 ;
      RECT 14.4640 36.9765 14.4900 38.0700 ;
      RECT 14.3560 36.9765 14.3820 38.0700 ;
      RECT 14.2480 36.9765 14.2740 38.0700 ;
      RECT 14.1400 36.9765 14.1660 38.0700 ;
      RECT 14.0320 36.9765 14.0580 38.0700 ;
      RECT 13.9240 36.9765 13.9500 38.0700 ;
      RECT 13.8160 36.9765 13.8420 38.0700 ;
      RECT 13.7080 36.9765 13.7340 38.0700 ;
      RECT 13.6000 36.9765 13.6260 38.0700 ;
      RECT 13.4920 36.9765 13.5180 38.0700 ;
      RECT 13.3840 36.9765 13.4100 38.0700 ;
      RECT 13.2760 36.9765 13.3020 38.0700 ;
      RECT 13.1680 36.9765 13.1940 38.0700 ;
      RECT 13.0600 36.9765 13.0860 38.0700 ;
      RECT 12.9520 36.9765 12.9780 38.0700 ;
      RECT 12.8440 36.9765 12.8700 38.0700 ;
      RECT 12.7360 36.9765 12.7620 38.0700 ;
      RECT 12.6280 36.9765 12.6540 38.0700 ;
      RECT 12.5200 36.9765 12.5460 38.0700 ;
      RECT 12.4120 36.9765 12.4380 38.0700 ;
      RECT 12.3040 36.9765 12.3300 38.0700 ;
      RECT 12.1960 36.9765 12.2220 38.0700 ;
      RECT 12.0880 36.9765 12.1140 38.0700 ;
      RECT 11.9800 36.9765 12.0060 38.0700 ;
      RECT 11.8720 36.9765 11.8980 38.0700 ;
      RECT 11.7640 36.9765 11.7900 38.0700 ;
      RECT 11.6560 36.9765 11.6820 38.0700 ;
      RECT 11.5480 36.9765 11.5740 38.0700 ;
      RECT 11.4400 36.9765 11.4660 38.0700 ;
      RECT 11.3320 36.9765 11.3580 38.0700 ;
      RECT 11.2240 36.9765 11.2500 38.0700 ;
      RECT 11.1160 36.9765 11.1420 38.0700 ;
      RECT 11.0080 36.9765 11.0340 38.0700 ;
      RECT 10.9000 36.9765 10.9260 38.0700 ;
      RECT 10.7920 36.9765 10.8180 38.0700 ;
      RECT 10.6840 36.9765 10.7100 38.0700 ;
      RECT 10.5760 36.9765 10.6020 38.0700 ;
      RECT 10.4680 36.9765 10.4940 38.0700 ;
      RECT 10.3600 36.9765 10.3860 38.0700 ;
      RECT 10.2520 36.9765 10.2780 38.0700 ;
      RECT 10.1440 36.9765 10.1700 38.0700 ;
      RECT 10.0360 36.9765 10.0620 38.0700 ;
      RECT 9.9280 36.9765 9.9540 38.0700 ;
      RECT 9.8200 36.9765 9.8460 38.0700 ;
      RECT 9.7120 36.9765 9.7380 38.0700 ;
      RECT 9.6040 36.9765 9.6300 38.0700 ;
      RECT 9.4960 36.9765 9.5220 38.0700 ;
      RECT 9.3880 36.9765 9.4140 38.0700 ;
      RECT 9.1750 36.9765 9.2520 38.0700 ;
      RECT 7.2820 36.9765 7.3590 38.0700 ;
      RECT 7.1200 36.9765 7.1460 38.0700 ;
      RECT 7.0120 36.9765 7.0380 38.0700 ;
      RECT 6.9040 36.9765 6.9300 38.0700 ;
      RECT 6.7960 36.9765 6.8220 38.0700 ;
      RECT 6.6880 36.9765 6.7140 38.0700 ;
      RECT 6.5800 36.9765 6.6060 38.0700 ;
      RECT 6.4720 36.9765 6.4980 38.0700 ;
      RECT 6.3640 36.9765 6.3900 38.0700 ;
      RECT 6.2560 36.9765 6.2820 38.0700 ;
      RECT 6.1480 36.9765 6.1740 38.0700 ;
      RECT 6.0400 36.9765 6.0660 38.0700 ;
      RECT 5.9320 36.9765 5.9580 38.0700 ;
      RECT 5.8240 36.9765 5.8500 38.0700 ;
      RECT 5.7160 36.9765 5.7420 38.0700 ;
      RECT 5.6080 36.9765 5.6340 38.0700 ;
      RECT 5.5000 36.9765 5.5260 38.0700 ;
      RECT 5.3920 36.9765 5.4180 38.0700 ;
      RECT 5.2840 36.9765 5.3100 38.0700 ;
      RECT 5.1760 36.9765 5.2020 38.0700 ;
      RECT 5.0680 36.9765 5.0940 38.0700 ;
      RECT 4.9600 36.9765 4.9860 38.0700 ;
      RECT 4.8520 36.9765 4.8780 38.0700 ;
      RECT 4.7440 36.9765 4.7700 38.0700 ;
      RECT 4.6360 36.9765 4.6620 38.0700 ;
      RECT 4.5280 36.9765 4.5540 38.0700 ;
      RECT 4.4200 36.9765 4.4460 38.0700 ;
      RECT 4.3120 36.9765 4.3380 38.0700 ;
      RECT 4.2040 36.9765 4.2300 38.0700 ;
      RECT 4.0960 36.9765 4.1220 38.0700 ;
      RECT 3.9880 36.9765 4.0140 38.0700 ;
      RECT 3.8800 36.9765 3.9060 38.0700 ;
      RECT 3.7720 36.9765 3.7980 38.0700 ;
      RECT 3.6640 36.9765 3.6900 38.0700 ;
      RECT 3.5560 36.9765 3.5820 38.0700 ;
      RECT 3.4480 36.9765 3.4740 38.0700 ;
      RECT 3.3400 36.9765 3.3660 38.0700 ;
      RECT 3.2320 36.9765 3.2580 38.0700 ;
      RECT 3.1240 36.9765 3.1500 38.0700 ;
      RECT 3.0160 36.9765 3.0420 38.0700 ;
      RECT 2.9080 36.9765 2.9340 38.0700 ;
      RECT 2.8000 36.9765 2.8260 38.0700 ;
      RECT 2.6920 36.9765 2.7180 38.0700 ;
      RECT 2.5840 36.9765 2.6100 38.0700 ;
      RECT 2.4760 36.9765 2.5020 38.0700 ;
      RECT 2.3680 36.9765 2.3940 38.0700 ;
      RECT 2.2600 36.9765 2.2860 38.0700 ;
      RECT 2.1520 36.9765 2.1780 38.0700 ;
      RECT 2.0440 36.9765 2.0700 38.0700 ;
      RECT 1.9360 36.9765 1.9620 38.0700 ;
      RECT 1.8280 36.9765 1.8540 38.0700 ;
      RECT 1.7200 36.9765 1.7460 38.0700 ;
      RECT 1.6120 36.9765 1.6380 38.0700 ;
      RECT 1.5040 36.9765 1.5300 38.0700 ;
      RECT 1.3960 36.9765 1.4220 38.0700 ;
      RECT 1.2880 36.9765 1.3140 38.0700 ;
      RECT 1.1800 36.9765 1.2060 38.0700 ;
      RECT 1.0720 36.9765 1.0980 38.0700 ;
      RECT 0.9640 36.9765 0.9900 38.0700 ;
      RECT 0.8560 36.9765 0.8820 38.0700 ;
      RECT 0.7480 36.9765 0.7740 38.0700 ;
      RECT 0.6400 36.9765 0.6660 38.0700 ;
      RECT 0.5320 36.9765 0.5580 38.0700 ;
      RECT 0.4240 36.9765 0.4500 38.0700 ;
      RECT 0.3160 36.9765 0.3420 38.0700 ;
      RECT 0.2080 36.9765 0.2340 38.0700 ;
      RECT 0.0050 36.9765 0.0900 38.0700 ;
      RECT 8.6410 38.0565 8.7690 39.1500 ;
      RECT 8.6270 38.7220 8.7690 39.0445 ;
      RECT 8.4790 38.4490 8.5410 39.1500 ;
      RECT 8.4650 38.7585 8.5410 38.9120 ;
      RECT 8.4790 38.0565 8.5050 39.1500 ;
      RECT 8.4790 38.1775 8.5190 38.4170 ;
      RECT 8.4790 38.0565 8.5410 38.1455 ;
      RECT 8.1820 38.5070 8.3880 39.1500 ;
      RECT 8.3620 38.0565 8.3880 39.1500 ;
      RECT 8.1820 38.7840 8.4020 39.0420 ;
      RECT 8.1820 38.0565 8.2800 39.1500 ;
      RECT 7.7650 38.0565 7.8480 39.1500 ;
      RECT 7.7650 38.1450 7.8620 39.0805 ;
      RECT 16.4440 38.0565 16.5290 39.1500 ;
      RECT 16.3000 38.0565 16.3260 39.1500 ;
      RECT 16.1920 38.0565 16.2180 39.1500 ;
      RECT 16.0840 38.0565 16.1100 39.1500 ;
      RECT 15.9760 38.0565 16.0020 39.1500 ;
      RECT 15.8680 38.0565 15.8940 39.1500 ;
      RECT 15.7600 38.0565 15.7860 39.1500 ;
      RECT 15.6520 38.0565 15.6780 39.1500 ;
      RECT 15.5440 38.0565 15.5700 39.1500 ;
      RECT 15.4360 38.0565 15.4620 39.1500 ;
      RECT 15.3280 38.0565 15.3540 39.1500 ;
      RECT 15.2200 38.0565 15.2460 39.1500 ;
      RECT 15.1120 38.0565 15.1380 39.1500 ;
      RECT 15.0040 38.0565 15.0300 39.1500 ;
      RECT 14.8960 38.0565 14.9220 39.1500 ;
      RECT 14.7880 38.0565 14.8140 39.1500 ;
      RECT 14.6800 38.0565 14.7060 39.1500 ;
      RECT 14.5720 38.0565 14.5980 39.1500 ;
      RECT 14.4640 38.0565 14.4900 39.1500 ;
      RECT 14.3560 38.0565 14.3820 39.1500 ;
      RECT 14.2480 38.0565 14.2740 39.1500 ;
      RECT 14.1400 38.0565 14.1660 39.1500 ;
      RECT 14.0320 38.0565 14.0580 39.1500 ;
      RECT 13.9240 38.0565 13.9500 39.1500 ;
      RECT 13.8160 38.0565 13.8420 39.1500 ;
      RECT 13.7080 38.0565 13.7340 39.1500 ;
      RECT 13.6000 38.0565 13.6260 39.1500 ;
      RECT 13.4920 38.0565 13.5180 39.1500 ;
      RECT 13.3840 38.0565 13.4100 39.1500 ;
      RECT 13.2760 38.0565 13.3020 39.1500 ;
      RECT 13.1680 38.0565 13.1940 39.1500 ;
      RECT 13.0600 38.0565 13.0860 39.1500 ;
      RECT 12.9520 38.0565 12.9780 39.1500 ;
      RECT 12.8440 38.0565 12.8700 39.1500 ;
      RECT 12.7360 38.0565 12.7620 39.1500 ;
      RECT 12.6280 38.0565 12.6540 39.1500 ;
      RECT 12.5200 38.0565 12.5460 39.1500 ;
      RECT 12.4120 38.0565 12.4380 39.1500 ;
      RECT 12.3040 38.0565 12.3300 39.1500 ;
      RECT 12.1960 38.0565 12.2220 39.1500 ;
      RECT 12.0880 38.0565 12.1140 39.1500 ;
      RECT 11.9800 38.0565 12.0060 39.1500 ;
      RECT 11.8720 38.0565 11.8980 39.1500 ;
      RECT 11.7640 38.0565 11.7900 39.1500 ;
      RECT 11.6560 38.0565 11.6820 39.1500 ;
      RECT 11.5480 38.0565 11.5740 39.1500 ;
      RECT 11.4400 38.0565 11.4660 39.1500 ;
      RECT 11.3320 38.0565 11.3580 39.1500 ;
      RECT 11.2240 38.0565 11.2500 39.1500 ;
      RECT 11.1160 38.0565 11.1420 39.1500 ;
      RECT 11.0080 38.0565 11.0340 39.1500 ;
      RECT 10.9000 38.0565 10.9260 39.1500 ;
      RECT 10.7920 38.0565 10.8180 39.1500 ;
      RECT 10.6840 38.0565 10.7100 39.1500 ;
      RECT 10.5760 38.0565 10.6020 39.1500 ;
      RECT 10.4680 38.0565 10.4940 39.1500 ;
      RECT 10.3600 38.0565 10.3860 39.1500 ;
      RECT 10.2520 38.0565 10.2780 39.1500 ;
      RECT 10.1440 38.0565 10.1700 39.1500 ;
      RECT 10.0360 38.0565 10.0620 39.1500 ;
      RECT 9.9280 38.0565 9.9540 39.1500 ;
      RECT 9.8200 38.0565 9.8460 39.1500 ;
      RECT 9.7120 38.0565 9.7380 39.1500 ;
      RECT 9.6040 38.0565 9.6300 39.1500 ;
      RECT 9.4960 38.0565 9.5220 39.1500 ;
      RECT 9.3880 38.0565 9.4140 39.1500 ;
      RECT 9.1750 38.0565 9.2520 39.1500 ;
      RECT 7.2820 38.0565 7.3590 39.1500 ;
      RECT 7.1200 38.0565 7.1460 39.1500 ;
      RECT 7.0120 38.0565 7.0380 39.1500 ;
      RECT 6.9040 38.0565 6.9300 39.1500 ;
      RECT 6.7960 38.0565 6.8220 39.1500 ;
      RECT 6.6880 38.0565 6.7140 39.1500 ;
      RECT 6.5800 38.0565 6.6060 39.1500 ;
      RECT 6.4720 38.0565 6.4980 39.1500 ;
      RECT 6.3640 38.0565 6.3900 39.1500 ;
      RECT 6.2560 38.0565 6.2820 39.1500 ;
      RECT 6.1480 38.0565 6.1740 39.1500 ;
      RECT 6.0400 38.0565 6.0660 39.1500 ;
      RECT 5.9320 38.0565 5.9580 39.1500 ;
      RECT 5.8240 38.0565 5.8500 39.1500 ;
      RECT 5.7160 38.0565 5.7420 39.1500 ;
      RECT 5.6080 38.0565 5.6340 39.1500 ;
      RECT 5.5000 38.0565 5.5260 39.1500 ;
      RECT 5.3920 38.0565 5.4180 39.1500 ;
      RECT 5.2840 38.0565 5.3100 39.1500 ;
      RECT 5.1760 38.0565 5.2020 39.1500 ;
      RECT 5.0680 38.0565 5.0940 39.1500 ;
      RECT 4.9600 38.0565 4.9860 39.1500 ;
      RECT 4.8520 38.0565 4.8780 39.1500 ;
      RECT 4.7440 38.0565 4.7700 39.1500 ;
      RECT 4.6360 38.0565 4.6620 39.1500 ;
      RECT 4.5280 38.0565 4.5540 39.1500 ;
      RECT 4.4200 38.0565 4.4460 39.1500 ;
      RECT 4.3120 38.0565 4.3380 39.1500 ;
      RECT 4.2040 38.0565 4.2300 39.1500 ;
      RECT 4.0960 38.0565 4.1220 39.1500 ;
      RECT 3.9880 38.0565 4.0140 39.1500 ;
      RECT 3.8800 38.0565 3.9060 39.1500 ;
      RECT 3.7720 38.0565 3.7980 39.1500 ;
      RECT 3.6640 38.0565 3.6900 39.1500 ;
      RECT 3.5560 38.0565 3.5820 39.1500 ;
      RECT 3.4480 38.0565 3.4740 39.1500 ;
      RECT 3.3400 38.0565 3.3660 39.1500 ;
      RECT 3.2320 38.0565 3.2580 39.1500 ;
      RECT 3.1240 38.0565 3.1500 39.1500 ;
      RECT 3.0160 38.0565 3.0420 39.1500 ;
      RECT 2.9080 38.0565 2.9340 39.1500 ;
      RECT 2.8000 38.0565 2.8260 39.1500 ;
      RECT 2.6920 38.0565 2.7180 39.1500 ;
      RECT 2.5840 38.0565 2.6100 39.1500 ;
      RECT 2.4760 38.0565 2.5020 39.1500 ;
      RECT 2.3680 38.0565 2.3940 39.1500 ;
      RECT 2.2600 38.0565 2.2860 39.1500 ;
      RECT 2.1520 38.0565 2.1780 39.1500 ;
      RECT 2.0440 38.0565 2.0700 39.1500 ;
      RECT 1.9360 38.0565 1.9620 39.1500 ;
      RECT 1.8280 38.0565 1.8540 39.1500 ;
      RECT 1.7200 38.0565 1.7460 39.1500 ;
      RECT 1.6120 38.0565 1.6380 39.1500 ;
      RECT 1.5040 38.0565 1.5300 39.1500 ;
      RECT 1.3960 38.0565 1.4220 39.1500 ;
      RECT 1.2880 38.0565 1.3140 39.1500 ;
      RECT 1.1800 38.0565 1.2060 39.1500 ;
      RECT 1.0720 38.0565 1.0980 39.1500 ;
      RECT 0.9640 38.0565 0.9900 39.1500 ;
      RECT 0.8560 38.0565 0.8820 39.1500 ;
      RECT 0.7480 38.0565 0.7740 39.1500 ;
      RECT 0.6400 38.0565 0.6660 39.1500 ;
      RECT 0.5320 38.0565 0.5580 39.1500 ;
      RECT 0.4240 38.0565 0.4500 39.1500 ;
      RECT 0.3160 38.0565 0.3420 39.1500 ;
      RECT 0.2080 38.0565 0.2340 39.1500 ;
      RECT 0.0050 38.0565 0.0900 39.1500 ;
      RECT 8.6410 39.1365 8.7690 40.2300 ;
      RECT 8.6270 39.8020 8.7690 40.1245 ;
      RECT 8.4790 39.5290 8.5410 40.2300 ;
      RECT 8.4650 39.8385 8.5410 39.9920 ;
      RECT 8.4790 39.1365 8.5050 40.2300 ;
      RECT 8.4790 39.2575 8.5190 39.4970 ;
      RECT 8.4790 39.1365 8.5410 39.2255 ;
      RECT 8.1820 39.5870 8.3880 40.2300 ;
      RECT 8.3620 39.1365 8.3880 40.2300 ;
      RECT 8.1820 39.8640 8.4020 40.1220 ;
      RECT 8.1820 39.1365 8.2800 40.2300 ;
      RECT 7.7650 39.1365 7.8480 40.2300 ;
      RECT 7.7650 39.2250 7.8620 40.1605 ;
      RECT 16.4440 39.1365 16.5290 40.2300 ;
      RECT 16.3000 39.1365 16.3260 40.2300 ;
      RECT 16.1920 39.1365 16.2180 40.2300 ;
      RECT 16.0840 39.1365 16.1100 40.2300 ;
      RECT 15.9760 39.1365 16.0020 40.2300 ;
      RECT 15.8680 39.1365 15.8940 40.2300 ;
      RECT 15.7600 39.1365 15.7860 40.2300 ;
      RECT 15.6520 39.1365 15.6780 40.2300 ;
      RECT 15.5440 39.1365 15.5700 40.2300 ;
      RECT 15.4360 39.1365 15.4620 40.2300 ;
      RECT 15.3280 39.1365 15.3540 40.2300 ;
      RECT 15.2200 39.1365 15.2460 40.2300 ;
      RECT 15.1120 39.1365 15.1380 40.2300 ;
      RECT 15.0040 39.1365 15.0300 40.2300 ;
      RECT 14.8960 39.1365 14.9220 40.2300 ;
      RECT 14.7880 39.1365 14.8140 40.2300 ;
      RECT 14.6800 39.1365 14.7060 40.2300 ;
      RECT 14.5720 39.1365 14.5980 40.2300 ;
      RECT 14.4640 39.1365 14.4900 40.2300 ;
      RECT 14.3560 39.1365 14.3820 40.2300 ;
      RECT 14.2480 39.1365 14.2740 40.2300 ;
      RECT 14.1400 39.1365 14.1660 40.2300 ;
      RECT 14.0320 39.1365 14.0580 40.2300 ;
      RECT 13.9240 39.1365 13.9500 40.2300 ;
      RECT 13.8160 39.1365 13.8420 40.2300 ;
      RECT 13.7080 39.1365 13.7340 40.2300 ;
      RECT 13.6000 39.1365 13.6260 40.2300 ;
      RECT 13.4920 39.1365 13.5180 40.2300 ;
      RECT 13.3840 39.1365 13.4100 40.2300 ;
      RECT 13.2760 39.1365 13.3020 40.2300 ;
      RECT 13.1680 39.1365 13.1940 40.2300 ;
      RECT 13.0600 39.1365 13.0860 40.2300 ;
      RECT 12.9520 39.1365 12.9780 40.2300 ;
      RECT 12.8440 39.1365 12.8700 40.2300 ;
      RECT 12.7360 39.1365 12.7620 40.2300 ;
      RECT 12.6280 39.1365 12.6540 40.2300 ;
      RECT 12.5200 39.1365 12.5460 40.2300 ;
      RECT 12.4120 39.1365 12.4380 40.2300 ;
      RECT 12.3040 39.1365 12.3300 40.2300 ;
      RECT 12.1960 39.1365 12.2220 40.2300 ;
      RECT 12.0880 39.1365 12.1140 40.2300 ;
      RECT 11.9800 39.1365 12.0060 40.2300 ;
      RECT 11.8720 39.1365 11.8980 40.2300 ;
      RECT 11.7640 39.1365 11.7900 40.2300 ;
      RECT 11.6560 39.1365 11.6820 40.2300 ;
      RECT 11.5480 39.1365 11.5740 40.2300 ;
      RECT 11.4400 39.1365 11.4660 40.2300 ;
      RECT 11.3320 39.1365 11.3580 40.2300 ;
      RECT 11.2240 39.1365 11.2500 40.2300 ;
      RECT 11.1160 39.1365 11.1420 40.2300 ;
      RECT 11.0080 39.1365 11.0340 40.2300 ;
      RECT 10.9000 39.1365 10.9260 40.2300 ;
      RECT 10.7920 39.1365 10.8180 40.2300 ;
      RECT 10.6840 39.1365 10.7100 40.2300 ;
      RECT 10.5760 39.1365 10.6020 40.2300 ;
      RECT 10.4680 39.1365 10.4940 40.2300 ;
      RECT 10.3600 39.1365 10.3860 40.2300 ;
      RECT 10.2520 39.1365 10.2780 40.2300 ;
      RECT 10.1440 39.1365 10.1700 40.2300 ;
      RECT 10.0360 39.1365 10.0620 40.2300 ;
      RECT 9.9280 39.1365 9.9540 40.2300 ;
      RECT 9.8200 39.1365 9.8460 40.2300 ;
      RECT 9.7120 39.1365 9.7380 40.2300 ;
      RECT 9.6040 39.1365 9.6300 40.2300 ;
      RECT 9.4960 39.1365 9.5220 40.2300 ;
      RECT 9.3880 39.1365 9.4140 40.2300 ;
      RECT 9.1750 39.1365 9.2520 40.2300 ;
      RECT 7.2820 39.1365 7.3590 40.2300 ;
      RECT 7.1200 39.1365 7.1460 40.2300 ;
      RECT 7.0120 39.1365 7.0380 40.2300 ;
      RECT 6.9040 39.1365 6.9300 40.2300 ;
      RECT 6.7960 39.1365 6.8220 40.2300 ;
      RECT 6.6880 39.1365 6.7140 40.2300 ;
      RECT 6.5800 39.1365 6.6060 40.2300 ;
      RECT 6.4720 39.1365 6.4980 40.2300 ;
      RECT 6.3640 39.1365 6.3900 40.2300 ;
      RECT 6.2560 39.1365 6.2820 40.2300 ;
      RECT 6.1480 39.1365 6.1740 40.2300 ;
      RECT 6.0400 39.1365 6.0660 40.2300 ;
      RECT 5.9320 39.1365 5.9580 40.2300 ;
      RECT 5.8240 39.1365 5.8500 40.2300 ;
      RECT 5.7160 39.1365 5.7420 40.2300 ;
      RECT 5.6080 39.1365 5.6340 40.2300 ;
      RECT 5.5000 39.1365 5.5260 40.2300 ;
      RECT 5.3920 39.1365 5.4180 40.2300 ;
      RECT 5.2840 39.1365 5.3100 40.2300 ;
      RECT 5.1760 39.1365 5.2020 40.2300 ;
      RECT 5.0680 39.1365 5.0940 40.2300 ;
      RECT 4.9600 39.1365 4.9860 40.2300 ;
      RECT 4.8520 39.1365 4.8780 40.2300 ;
      RECT 4.7440 39.1365 4.7700 40.2300 ;
      RECT 4.6360 39.1365 4.6620 40.2300 ;
      RECT 4.5280 39.1365 4.5540 40.2300 ;
      RECT 4.4200 39.1365 4.4460 40.2300 ;
      RECT 4.3120 39.1365 4.3380 40.2300 ;
      RECT 4.2040 39.1365 4.2300 40.2300 ;
      RECT 4.0960 39.1365 4.1220 40.2300 ;
      RECT 3.9880 39.1365 4.0140 40.2300 ;
      RECT 3.8800 39.1365 3.9060 40.2300 ;
      RECT 3.7720 39.1365 3.7980 40.2300 ;
      RECT 3.6640 39.1365 3.6900 40.2300 ;
      RECT 3.5560 39.1365 3.5820 40.2300 ;
      RECT 3.4480 39.1365 3.4740 40.2300 ;
      RECT 3.3400 39.1365 3.3660 40.2300 ;
      RECT 3.2320 39.1365 3.2580 40.2300 ;
      RECT 3.1240 39.1365 3.1500 40.2300 ;
      RECT 3.0160 39.1365 3.0420 40.2300 ;
      RECT 2.9080 39.1365 2.9340 40.2300 ;
      RECT 2.8000 39.1365 2.8260 40.2300 ;
      RECT 2.6920 39.1365 2.7180 40.2300 ;
      RECT 2.5840 39.1365 2.6100 40.2300 ;
      RECT 2.4760 39.1365 2.5020 40.2300 ;
      RECT 2.3680 39.1365 2.3940 40.2300 ;
      RECT 2.2600 39.1365 2.2860 40.2300 ;
      RECT 2.1520 39.1365 2.1780 40.2300 ;
      RECT 2.0440 39.1365 2.0700 40.2300 ;
      RECT 1.9360 39.1365 1.9620 40.2300 ;
      RECT 1.8280 39.1365 1.8540 40.2300 ;
      RECT 1.7200 39.1365 1.7460 40.2300 ;
      RECT 1.6120 39.1365 1.6380 40.2300 ;
      RECT 1.5040 39.1365 1.5300 40.2300 ;
      RECT 1.3960 39.1365 1.4220 40.2300 ;
      RECT 1.2880 39.1365 1.3140 40.2300 ;
      RECT 1.1800 39.1365 1.2060 40.2300 ;
      RECT 1.0720 39.1365 1.0980 40.2300 ;
      RECT 0.9640 39.1365 0.9900 40.2300 ;
      RECT 0.8560 39.1365 0.8820 40.2300 ;
      RECT 0.7480 39.1365 0.7740 40.2300 ;
      RECT 0.6400 39.1365 0.6660 40.2300 ;
      RECT 0.5320 39.1365 0.5580 40.2300 ;
      RECT 0.4240 39.1365 0.4500 40.2300 ;
      RECT 0.3160 39.1365 0.3420 40.2300 ;
      RECT 0.2080 39.1365 0.2340 40.2300 ;
      RECT 0.0050 39.1365 0.0900 40.2300 ;
      RECT 0.0000 48.4095 16.5240 48.8505 ;
      RECT 16.4390 40.1970 16.5240 48.8505 ;
      RECT 9.3830 41.7010 16.3210 48.8505 ;
      RECT 10.8410 40.1970 16.3210 48.8505 ;
      RECT 7.2230 48.4020 9.3010 48.8505 ;
      RECT 7.9970 48.3705 9.3010 48.8505 ;
      RECT 0.2030 41.5060 7.1410 48.8505 ;
      RECT 6.8450 40.1970 7.1410 48.8505 ;
      RECT 0.0000 40.1970 0.0850 48.8505 ;
      RECT 7.2230 41.8090 7.8430 48.8505 ;
      RECT 7.9970 48.3660 9.2650 48.8505 ;
      RECT 8.6450 41.6020 9.2650 48.8505 ;
      RECT 8.6360 48.1090 9.2650 48.8505 ;
      RECT 8.4740 48.1090 8.5360 48.8505 ;
      RECT 7.9970 48.1090 8.3830 48.8505 ;
      RECT 9.3830 43.9900 16.3350 48.3440 ;
      RECT 0.1890 43.9900 7.1410 48.3440 ;
      RECT 9.3690 43.9900 16.3350 48.3395 ;
      RECT 0.1890 43.9900 7.1550 48.3395 ;
      RECT 7.2090 43.9900 7.8430 48.3385 ;
      RECT 8.1770 40.8820 8.3470 48.8505 ;
      RECT 8.2850 40.1970 8.3470 48.8505 ;
      RECT 7.4930 40.6180 7.8790 47.9620 ;
      RECT 7.2090 47.9170 7.8930 47.9540 ;
      RECT 8.6310 46.8430 9.2650 47.9510 ;
      RECT 8.1630 47.6530 8.3470 47.8790 ;
      RECT 8.1770 47.0770 8.3610 47.3390 ;
      RECT 7.2090 46.8790 7.8930 47.3390 ;
      RECT 8.1630 46.3390 8.3470 46.7990 ;
      RECT 8.6310 44.3050 9.2650 46.6370 ;
      RECT 7.2090 44.9530 7.8930 46.0970 ;
      RECT 8.1770 44.6830 8.3610 45.9890 ;
      RECT 8.1630 45.2590 8.3610 45.7190 ;
      RECT 8.1630 42.0190 8.3470 45.1790 ;
      RECT 8.1630 42.0190 8.3610 44.6390 ;
      RECT 7.2090 44.4130 7.8930 44.6390 ;
      RECT 8.6450 41.6020 9.3010 43.9580 ;
      RECT 8.6310 41.4790 9.2470 43.2650 ;
      RECT 7.2230 42.4510 7.8930 42.8210 ;
      RECT 8.1770 41.7490 8.3610 41.9390 ;
      RECT 7.2770 41.7130 7.8930 41.9030 ;
      RECT 8.1630 41.6050 8.3470 41.7410 ;
      RECT 7.2770 40.9630 7.8790 47.9620 ;
      RECT 8.1770 41.4790 8.3610 41.7050 ;
      RECT 9.5450 41.5090 16.3210 48.8505 ;
      RECT 10.6250 41.5060 16.3210 48.8505 ;
      RECT 9.3830 40.1970 9.4630 48.8505 ;
      RECT 7.2230 40.8820 7.4110 41.6960 ;
      RECT 9.3830 40.1970 9.6790 41.6000 ;
      RECT 9.3830 41.3140 10.5430 41.6000 ;
      RECT 10.6250 40.1970 10.7590 48.8505 ;
      RECT 5.9810 41.1250 6.7630 48.8505 ;
      RECT 0.2030 40.1970 5.8990 48.8505 ;
      RECT 8.6450 40.9630 9.2470 48.8505 ;
      RECT 8.6810 40.3735 9.3010 41.4470 ;
      RECT 9.3830 41.3140 10.7590 41.4080 ;
      RECT 10.4090 40.1970 16.3210 41.4050 ;
      RECT 6.6290 40.1970 7.1410 41.4050 ;
      RECT 8.1630 41.3350 8.3610 41.3990 ;
      RECT 8.1630 41.2090 8.3470 41.3990 ;
      RECT 10.1930 40.9300 16.3210 41.4050 ;
      RECT 9.3830 40.9630 10.1110 41.6000 ;
      RECT 8.1770 40.9390 8.3610 41.2010 ;
      RECT 0.2030 40.9300 6.5470 41.4050 ;
      RECT 6.4130 40.1970 6.5470 48.8505 ;
      RECT 9.9770 40.1970 10.3270 41.0690 ;
      RECT 9.3830 40.8820 9.8950 41.6000 ;
      RECT 9.7610 40.1970 9.8950 48.8505 ;
      RECT 6.1970 40.8820 6.5470 48.8505 ;
      RECT 0.2030 40.1970 6.1150 41.4050 ;
      RECT 8.1770 40.1970 8.2030 48.8505 ;
      RECT 7.3130 40.1970 7.4110 48.8505 ;
      RECT 6.1970 40.1970 6.3310 48.8505 ;
      RECT 9.7610 40.1970 10.3270 40.8320 ;
      RECT 8.6450 40.1970 9.2470 40.8320 ;
      RECT 7.3130 40.1970 7.8430 40.8320 ;
      RECT 6.4130 40.1970 7.1410 40.8320 ;
      RECT 9.7610 40.1970 16.3210 40.8290 ;
      RECT 0.2030 40.1970 6.3310 40.8290 ;
      RECT 8.6310 40.6690 9.3010 40.8230 ;
      RECT 9.3830 40.1970 16.3210 40.5650 ;
      RECT 8.1770 40.1970 8.3470 40.5650 ;
      RECT 7.2230 40.1970 7.8430 40.5650 ;
      RECT 0.2030 40.1970 7.1410 40.5650 ;
      RECT 7.9970 40.1970 8.3470 40.4620 ;
      RECT 8.6360 40.1970 9.2470 40.3620 ;
      RECT 7.9970 40.1970 8.3830 40.3620 ;
      RECT 9.7650 40.1705 9.7830 48.8505 ;
      RECT 9.6570 40.1705 9.6750 48.8505 ;
      RECT 6.8490 40.1830 6.8670 48.8505 ;
      RECT 6.7410 40.1830 6.7590 48.8505 ;
      RECT 6.6330 40.1830 6.6510 48.8505 ;
      RECT 6.5250 40.1830 6.5430 48.8505 ;
      RECT 6.4170 40.1705 6.4350 48.8505 ;
      RECT 6.3090 40.1705 6.3270 48.8505 ;
      RECT 6.2010 40.1830 6.2190 48.8505 ;
      RECT 6.0930 40.1830 6.1110 48.8505 ;
      RECT 5.9850 40.1830 6.0030 48.8505 ;
      RECT 5.8770 40.1830 5.8950 48.8505 ;
      RECT 8.4740 40.1970 8.5360 40.3620 ;
        RECT 8.6410 48.3435 8.7690 49.4370 ;
        RECT 8.6270 49.0090 8.7690 49.3315 ;
        RECT 8.4790 48.7360 8.5410 49.4370 ;
        RECT 8.4650 49.0455 8.5410 49.1990 ;
        RECT 8.4790 48.3435 8.5050 49.4370 ;
        RECT 8.4790 48.4645 8.5190 48.7040 ;
        RECT 8.4790 48.3435 8.5410 48.4325 ;
        RECT 8.1820 48.7940 8.3880 49.4370 ;
        RECT 8.3620 48.3435 8.3880 49.4370 ;
        RECT 8.1820 49.0710 8.4020 49.3290 ;
        RECT 8.1820 48.3435 8.2800 49.4370 ;
        RECT 7.7650 48.3435 7.8480 49.4370 ;
        RECT 7.7650 48.4320 7.8620 49.3675 ;
        RECT 16.4440 48.3435 16.5290 49.4370 ;
        RECT 16.3000 48.3435 16.3260 49.4370 ;
        RECT 16.1920 48.3435 16.2180 49.4370 ;
        RECT 16.0840 48.3435 16.1100 49.4370 ;
        RECT 15.9760 48.3435 16.0020 49.4370 ;
        RECT 15.8680 48.3435 15.8940 49.4370 ;
        RECT 15.7600 48.3435 15.7860 49.4370 ;
        RECT 15.6520 48.3435 15.6780 49.4370 ;
        RECT 15.5440 48.3435 15.5700 49.4370 ;
        RECT 15.4360 48.3435 15.4620 49.4370 ;
        RECT 15.3280 48.3435 15.3540 49.4370 ;
        RECT 15.2200 48.3435 15.2460 49.4370 ;
        RECT 15.1120 48.3435 15.1380 49.4370 ;
        RECT 15.0040 48.3435 15.0300 49.4370 ;
        RECT 14.8960 48.3435 14.9220 49.4370 ;
        RECT 14.7880 48.3435 14.8140 49.4370 ;
        RECT 14.6800 48.3435 14.7060 49.4370 ;
        RECT 14.5720 48.3435 14.5980 49.4370 ;
        RECT 14.4640 48.3435 14.4900 49.4370 ;
        RECT 14.3560 48.3435 14.3820 49.4370 ;
        RECT 14.2480 48.3435 14.2740 49.4370 ;
        RECT 14.1400 48.3435 14.1660 49.4370 ;
        RECT 14.0320 48.3435 14.0580 49.4370 ;
        RECT 13.9240 48.3435 13.9500 49.4370 ;
        RECT 13.8160 48.3435 13.8420 49.4370 ;
        RECT 13.7080 48.3435 13.7340 49.4370 ;
        RECT 13.6000 48.3435 13.6260 49.4370 ;
        RECT 13.4920 48.3435 13.5180 49.4370 ;
        RECT 13.3840 48.3435 13.4100 49.4370 ;
        RECT 13.2760 48.3435 13.3020 49.4370 ;
        RECT 13.1680 48.3435 13.1940 49.4370 ;
        RECT 13.0600 48.3435 13.0860 49.4370 ;
        RECT 12.9520 48.3435 12.9780 49.4370 ;
        RECT 12.8440 48.3435 12.8700 49.4370 ;
        RECT 12.7360 48.3435 12.7620 49.4370 ;
        RECT 12.6280 48.3435 12.6540 49.4370 ;
        RECT 12.5200 48.3435 12.5460 49.4370 ;
        RECT 12.4120 48.3435 12.4380 49.4370 ;
        RECT 12.3040 48.3435 12.3300 49.4370 ;
        RECT 12.1960 48.3435 12.2220 49.4370 ;
        RECT 12.0880 48.3435 12.1140 49.4370 ;
        RECT 11.9800 48.3435 12.0060 49.4370 ;
        RECT 11.8720 48.3435 11.8980 49.4370 ;
        RECT 11.7640 48.3435 11.7900 49.4370 ;
        RECT 11.6560 48.3435 11.6820 49.4370 ;
        RECT 11.5480 48.3435 11.5740 49.4370 ;
        RECT 11.4400 48.3435 11.4660 49.4370 ;
        RECT 11.3320 48.3435 11.3580 49.4370 ;
        RECT 11.2240 48.3435 11.2500 49.4370 ;
        RECT 11.1160 48.3435 11.1420 49.4370 ;
        RECT 11.0080 48.3435 11.0340 49.4370 ;
        RECT 10.9000 48.3435 10.9260 49.4370 ;
        RECT 10.7920 48.3435 10.8180 49.4370 ;
        RECT 10.6840 48.3435 10.7100 49.4370 ;
        RECT 10.5760 48.3435 10.6020 49.4370 ;
        RECT 10.4680 48.3435 10.4940 49.4370 ;
        RECT 10.3600 48.3435 10.3860 49.4370 ;
        RECT 10.2520 48.3435 10.2780 49.4370 ;
        RECT 10.1440 48.3435 10.1700 49.4370 ;
        RECT 10.0360 48.3435 10.0620 49.4370 ;
        RECT 9.9280 48.3435 9.9540 49.4370 ;
        RECT 9.8200 48.3435 9.8460 49.4370 ;
        RECT 9.7120 48.3435 9.7380 49.4370 ;
        RECT 9.6040 48.3435 9.6300 49.4370 ;
        RECT 9.4960 48.3435 9.5220 49.4370 ;
        RECT 9.3880 48.3435 9.4140 49.4370 ;
        RECT 9.1750 48.3435 9.2520 49.4370 ;
        RECT 7.2820 48.3435 7.3590 49.4370 ;
        RECT 7.1200 48.3435 7.1460 49.4370 ;
        RECT 7.0120 48.3435 7.0380 49.4370 ;
        RECT 6.9040 48.3435 6.9300 49.4370 ;
        RECT 6.7960 48.3435 6.8220 49.4370 ;
        RECT 6.6880 48.3435 6.7140 49.4370 ;
        RECT 6.5800 48.3435 6.6060 49.4370 ;
        RECT 6.4720 48.3435 6.4980 49.4370 ;
        RECT 6.3640 48.3435 6.3900 49.4370 ;
        RECT 6.2560 48.3435 6.2820 49.4370 ;
        RECT 6.1480 48.3435 6.1740 49.4370 ;
        RECT 6.0400 48.3435 6.0660 49.4370 ;
        RECT 5.9320 48.3435 5.9580 49.4370 ;
        RECT 5.8240 48.3435 5.8500 49.4370 ;
        RECT 5.7160 48.3435 5.7420 49.4370 ;
        RECT 5.6080 48.3435 5.6340 49.4370 ;
        RECT 5.5000 48.3435 5.5260 49.4370 ;
        RECT 5.3920 48.3435 5.4180 49.4370 ;
        RECT 5.2840 48.3435 5.3100 49.4370 ;
        RECT 5.1760 48.3435 5.2020 49.4370 ;
        RECT 5.0680 48.3435 5.0940 49.4370 ;
        RECT 4.9600 48.3435 4.9860 49.4370 ;
        RECT 4.8520 48.3435 4.8780 49.4370 ;
        RECT 4.7440 48.3435 4.7700 49.4370 ;
        RECT 4.6360 48.3435 4.6620 49.4370 ;
        RECT 4.5280 48.3435 4.5540 49.4370 ;
        RECT 4.4200 48.3435 4.4460 49.4370 ;
        RECT 4.3120 48.3435 4.3380 49.4370 ;
        RECT 4.2040 48.3435 4.2300 49.4370 ;
        RECT 4.0960 48.3435 4.1220 49.4370 ;
        RECT 3.9880 48.3435 4.0140 49.4370 ;
        RECT 3.8800 48.3435 3.9060 49.4370 ;
        RECT 3.7720 48.3435 3.7980 49.4370 ;
        RECT 3.6640 48.3435 3.6900 49.4370 ;
        RECT 3.5560 48.3435 3.5820 49.4370 ;
        RECT 3.4480 48.3435 3.4740 49.4370 ;
        RECT 3.3400 48.3435 3.3660 49.4370 ;
        RECT 3.2320 48.3435 3.2580 49.4370 ;
        RECT 3.1240 48.3435 3.1500 49.4370 ;
        RECT 3.0160 48.3435 3.0420 49.4370 ;
        RECT 2.9080 48.3435 2.9340 49.4370 ;
        RECT 2.8000 48.3435 2.8260 49.4370 ;
        RECT 2.6920 48.3435 2.7180 49.4370 ;
        RECT 2.5840 48.3435 2.6100 49.4370 ;
        RECT 2.4760 48.3435 2.5020 49.4370 ;
        RECT 2.3680 48.3435 2.3940 49.4370 ;
        RECT 2.2600 48.3435 2.2860 49.4370 ;
        RECT 2.1520 48.3435 2.1780 49.4370 ;
        RECT 2.0440 48.3435 2.0700 49.4370 ;
        RECT 1.9360 48.3435 1.9620 49.4370 ;
        RECT 1.8280 48.3435 1.8540 49.4370 ;
        RECT 1.7200 48.3435 1.7460 49.4370 ;
        RECT 1.6120 48.3435 1.6380 49.4370 ;
        RECT 1.5040 48.3435 1.5300 49.4370 ;
        RECT 1.3960 48.3435 1.4220 49.4370 ;
        RECT 1.2880 48.3435 1.3140 49.4370 ;
        RECT 1.1800 48.3435 1.2060 49.4370 ;
        RECT 1.0720 48.3435 1.0980 49.4370 ;
        RECT 0.9640 48.3435 0.9900 49.4370 ;
        RECT 0.8560 48.3435 0.8820 49.4370 ;
        RECT 0.7480 48.3435 0.7740 49.4370 ;
        RECT 0.6400 48.3435 0.6660 49.4370 ;
        RECT 0.5320 48.3435 0.5580 49.4370 ;
        RECT 0.4240 48.3435 0.4500 49.4370 ;
        RECT 0.3160 48.3435 0.3420 49.4370 ;
        RECT 0.2080 48.3435 0.2340 49.4370 ;
        RECT 0.0050 48.3435 0.0900 49.4370 ;
        RECT 8.6410 49.4235 8.7690 50.5170 ;
        RECT 8.6270 50.0890 8.7690 50.4115 ;
        RECT 8.4790 49.8160 8.5410 50.5170 ;
        RECT 8.4650 50.1255 8.5410 50.2790 ;
        RECT 8.4790 49.4235 8.5050 50.5170 ;
        RECT 8.4790 49.5445 8.5190 49.7840 ;
        RECT 8.4790 49.4235 8.5410 49.5125 ;
        RECT 8.1820 49.8740 8.3880 50.5170 ;
        RECT 8.3620 49.4235 8.3880 50.5170 ;
        RECT 8.1820 50.1510 8.4020 50.4090 ;
        RECT 8.1820 49.4235 8.2800 50.5170 ;
        RECT 7.7650 49.4235 7.8480 50.5170 ;
        RECT 7.7650 49.5120 7.8620 50.4475 ;
        RECT 16.4440 49.4235 16.5290 50.5170 ;
        RECT 16.3000 49.4235 16.3260 50.5170 ;
        RECT 16.1920 49.4235 16.2180 50.5170 ;
        RECT 16.0840 49.4235 16.1100 50.5170 ;
        RECT 15.9760 49.4235 16.0020 50.5170 ;
        RECT 15.8680 49.4235 15.8940 50.5170 ;
        RECT 15.7600 49.4235 15.7860 50.5170 ;
        RECT 15.6520 49.4235 15.6780 50.5170 ;
        RECT 15.5440 49.4235 15.5700 50.5170 ;
        RECT 15.4360 49.4235 15.4620 50.5170 ;
        RECT 15.3280 49.4235 15.3540 50.5170 ;
        RECT 15.2200 49.4235 15.2460 50.5170 ;
        RECT 15.1120 49.4235 15.1380 50.5170 ;
        RECT 15.0040 49.4235 15.0300 50.5170 ;
        RECT 14.8960 49.4235 14.9220 50.5170 ;
        RECT 14.7880 49.4235 14.8140 50.5170 ;
        RECT 14.6800 49.4235 14.7060 50.5170 ;
        RECT 14.5720 49.4235 14.5980 50.5170 ;
        RECT 14.4640 49.4235 14.4900 50.5170 ;
        RECT 14.3560 49.4235 14.3820 50.5170 ;
        RECT 14.2480 49.4235 14.2740 50.5170 ;
        RECT 14.1400 49.4235 14.1660 50.5170 ;
        RECT 14.0320 49.4235 14.0580 50.5170 ;
        RECT 13.9240 49.4235 13.9500 50.5170 ;
        RECT 13.8160 49.4235 13.8420 50.5170 ;
        RECT 13.7080 49.4235 13.7340 50.5170 ;
        RECT 13.6000 49.4235 13.6260 50.5170 ;
        RECT 13.4920 49.4235 13.5180 50.5170 ;
        RECT 13.3840 49.4235 13.4100 50.5170 ;
        RECT 13.2760 49.4235 13.3020 50.5170 ;
        RECT 13.1680 49.4235 13.1940 50.5170 ;
        RECT 13.0600 49.4235 13.0860 50.5170 ;
        RECT 12.9520 49.4235 12.9780 50.5170 ;
        RECT 12.8440 49.4235 12.8700 50.5170 ;
        RECT 12.7360 49.4235 12.7620 50.5170 ;
        RECT 12.6280 49.4235 12.6540 50.5170 ;
        RECT 12.5200 49.4235 12.5460 50.5170 ;
        RECT 12.4120 49.4235 12.4380 50.5170 ;
        RECT 12.3040 49.4235 12.3300 50.5170 ;
        RECT 12.1960 49.4235 12.2220 50.5170 ;
        RECT 12.0880 49.4235 12.1140 50.5170 ;
        RECT 11.9800 49.4235 12.0060 50.5170 ;
        RECT 11.8720 49.4235 11.8980 50.5170 ;
        RECT 11.7640 49.4235 11.7900 50.5170 ;
        RECT 11.6560 49.4235 11.6820 50.5170 ;
        RECT 11.5480 49.4235 11.5740 50.5170 ;
        RECT 11.4400 49.4235 11.4660 50.5170 ;
        RECT 11.3320 49.4235 11.3580 50.5170 ;
        RECT 11.2240 49.4235 11.2500 50.5170 ;
        RECT 11.1160 49.4235 11.1420 50.5170 ;
        RECT 11.0080 49.4235 11.0340 50.5170 ;
        RECT 10.9000 49.4235 10.9260 50.5170 ;
        RECT 10.7920 49.4235 10.8180 50.5170 ;
        RECT 10.6840 49.4235 10.7100 50.5170 ;
        RECT 10.5760 49.4235 10.6020 50.5170 ;
        RECT 10.4680 49.4235 10.4940 50.5170 ;
        RECT 10.3600 49.4235 10.3860 50.5170 ;
        RECT 10.2520 49.4235 10.2780 50.5170 ;
        RECT 10.1440 49.4235 10.1700 50.5170 ;
        RECT 10.0360 49.4235 10.0620 50.5170 ;
        RECT 9.9280 49.4235 9.9540 50.5170 ;
        RECT 9.8200 49.4235 9.8460 50.5170 ;
        RECT 9.7120 49.4235 9.7380 50.5170 ;
        RECT 9.6040 49.4235 9.6300 50.5170 ;
        RECT 9.4960 49.4235 9.5220 50.5170 ;
        RECT 9.3880 49.4235 9.4140 50.5170 ;
        RECT 9.1750 49.4235 9.2520 50.5170 ;
        RECT 7.2820 49.4235 7.3590 50.5170 ;
        RECT 7.1200 49.4235 7.1460 50.5170 ;
        RECT 7.0120 49.4235 7.0380 50.5170 ;
        RECT 6.9040 49.4235 6.9300 50.5170 ;
        RECT 6.7960 49.4235 6.8220 50.5170 ;
        RECT 6.6880 49.4235 6.7140 50.5170 ;
        RECT 6.5800 49.4235 6.6060 50.5170 ;
        RECT 6.4720 49.4235 6.4980 50.5170 ;
        RECT 6.3640 49.4235 6.3900 50.5170 ;
        RECT 6.2560 49.4235 6.2820 50.5170 ;
        RECT 6.1480 49.4235 6.1740 50.5170 ;
        RECT 6.0400 49.4235 6.0660 50.5170 ;
        RECT 5.9320 49.4235 5.9580 50.5170 ;
        RECT 5.8240 49.4235 5.8500 50.5170 ;
        RECT 5.7160 49.4235 5.7420 50.5170 ;
        RECT 5.6080 49.4235 5.6340 50.5170 ;
        RECT 5.5000 49.4235 5.5260 50.5170 ;
        RECT 5.3920 49.4235 5.4180 50.5170 ;
        RECT 5.2840 49.4235 5.3100 50.5170 ;
        RECT 5.1760 49.4235 5.2020 50.5170 ;
        RECT 5.0680 49.4235 5.0940 50.5170 ;
        RECT 4.9600 49.4235 4.9860 50.5170 ;
        RECT 4.8520 49.4235 4.8780 50.5170 ;
        RECT 4.7440 49.4235 4.7700 50.5170 ;
        RECT 4.6360 49.4235 4.6620 50.5170 ;
        RECT 4.5280 49.4235 4.5540 50.5170 ;
        RECT 4.4200 49.4235 4.4460 50.5170 ;
        RECT 4.3120 49.4235 4.3380 50.5170 ;
        RECT 4.2040 49.4235 4.2300 50.5170 ;
        RECT 4.0960 49.4235 4.1220 50.5170 ;
        RECT 3.9880 49.4235 4.0140 50.5170 ;
        RECT 3.8800 49.4235 3.9060 50.5170 ;
        RECT 3.7720 49.4235 3.7980 50.5170 ;
        RECT 3.6640 49.4235 3.6900 50.5170 ;
        RECT 3.5560 49.4235 3.5820 50.5170 ;
        RECT 3.4480 49.4235 3.4740 50.5170 ;
        RECT 3.3400 49.4235 3.3660 50.5170 ;
        RECT 3.2320 49.4235 3.2580 50.5170 ;
        RECT 3.1240 49.4235 3.1500 50.5170 ;
        RECT 3.0160 49.4235 3.0420 50.5170 ;
        RECT 2.9080 49.4235 2.9340 50.5170 ;
        RECT 2.8000 49.4235 2.8260 50.5170 ;
        RECT 2.6920 49.4235 2.7180 50.5170 ;
        RECT 2.5840 49.4235 2.6100 50.5170 ;
        RECT 2.4760 49.4235 2.5020 50.5170 ;
        RECT 2.3680 49.4235 2.3940 50.5170 ;
        RECT 2.2600 49.4235 2.2860 50.5170 ;
        RECT 2.1520 49.4235 2.1780 50.5170 ;
        RECT 2.0440 49.4235 2.0700 50.5170 ;
        RECT 1.9360 49.4235 1.9620 50.5170 ;
        RECT 1.8280 49.4235 1.8540 50.5170 ;
        RECT 1.7200 49.4235 1.7460 50.5170 ;
        RECT 1.6120 49.4235 1.6380 50.5170 ;
        RECT 1.5040 49.4235 1.5300 50.5170 ;
        RECT 1.3960 49.4235 1.4220 50.5170 ;
        RECT 1.2880 49.4235 1.3140 50.5170 ;
        RECT 1.1800 49.4235 1.2060 50.5170 ;
        RECT 1.0720 49.4235 1.0980 50.5170 ;
        RECT 0.9640 49.4235 0.9900 50.5170 ;
        RECT 0.8560 49.4235 0.8820 50.5170 ;
        RECT 0.7480 49.4235 0.7740 50.5170 ;
        RECT 0.6400 49.4235 0.6660 50.5170 ;
        RECT 0.5320 49.4235 0.5580 50.5170 ;
        RECT 0.4240 49.4235 0.4500 50.5170 ;
        RECT 0.3160 49.4235 0.3420 50.5170 ;
        RECT 0.2080 49.4235 0.2340 50.5170 ;
        RECT 0.0050 49.4235 0.0900 50.5170 ;
        RECT 8.6410 50.5035 8.7690 51.5970 ;
        RECT 8.6270 51.1690 8.7690 51.4915 ;
        RECT 8.4790 50.8960 8.5410 51.5970 ;
        RECT 8.4650 51.2055 8.5410 51.3590 ;
        RECT 8.4790 50.5035 8.5050 51.5970 ;
        RECT 8.4790 50.6245 8.5190 50.8640 ;
        RECT 8.4790 50.5035 8.5410 50.5925 ;
        RECT 8.1820 50.9540 8.3880 51.5970 ;
        RECT 8.3620 50.5035 8.3880 51.5970 ;
        RECT 8.1820 51.2310 8.4020 51.4890 ;
        RECT 8.1820 50.5035 8.2800 51.5970 ;
        RECT 7.7650 50.5035 7.8480 51.5970 ;
        RECT 7.7650 50.5920 7.8620 51.5275 ;
        RECT 16.4440 50.5035 16.5290 51.5970 ;
        RECT 16.3000 50.5035 16.3260 51.5970 ;
        RECT 16.1920 50.5035 16.2180 51.5970 ;
        RECT 16.0840 50.5035 16.1100 51.5970 ;
        RECT 15.9760 50.5035 16.0020 51.5970 ;
        RECT 15.8680 50.5035 15.8940 51.5970 ;
        RECT 15.7600 50.5035 15.7860 51.5970 ;
        RECT 15.6520 50.5035 15.6780 51.5970 ;
        RECT 15.5440 50.5035 15.5700 51.5970 ;
        RECT 15.4360 50.5035 15.4620 51.5970 ;
        RECT 15.3280 50.5035 15.3540 51.5970 ;
        RECT 15.2200 50.5035 15.2460 51.5970 ;
        RECT 15.1120 50.5035 15.1380 51.5970 ;
        RECT 15.0040 50.5035 15.0300 51.5970 ;
        RECT 14.8960 50.5035 14.9220 51.5970 ;
        RECT 14.7880 50.5035 14.8140 51.5970 ;
        RECT 14.6800 50.5035 14.7060 51.5970 ;
        RECT 14.5720 50.5035 14.5980 51.5970 ;
        RECT 14.4640 50.5035 14.4900 51.5970 ;
        RECT 14.3560 50.5035 14.3820 51.5970 ;
        RECT 14.2480 50.5035 14.2740 51.5970 ;
        RECT 14.1400 50.5035 14.1660 51.5970 ;
        RECT 14.0320 50.5035 14.0580 51.5970 ;
        RECT 13.9240 50.5035 13.9500 51.5970 ;
        RECT 13.8160 50.5035 13.8420 51.5970 ;
        RECT 13.7080 50.5035 13.7340 51.5970 ;
        RECT 13.6000 50.5035 13.6260 51.5970 ;
        RECT 13.4920 50.5035 13.5180 51.5970 ;
        RECT 13.3840 50.5035 13.4100 51.5970 ;
        RECT 13.2760 50.5035 13.3020 51.5970 ;
        RECT 13.1680 50.5035 13.1940 51.5970 ;
        RECT 13.0600 50.5035 13.0860 51.5970 ;
        RECT 12.9520 50.5035 12.9780 51.5970 ;
        RECT 12.8440 50.5035 12.8700 51.5970 ;
        RECT 12.7360 50.5035 12.7620 51.5970 ;
        RECT 12.6280 50.5035 12.6540 51.5970 ;
        RECT 12.5200 50.5035 12.5460 51.5970 ;
        RECT 12.4120 50.5035 12.4380 51.5970 ;
        RECT 12.3040 50.5035 12.3300 51.5970 ;
        RECT 12.1960 50.5035 12.2220 51.5970 ;
        RECT 12.0880 50.5035 12.1140 51.5970 ;
        RECT 11.9800 50.5035 12.0060 51.5970 ;
        RECT 11.8720 50.5035 11.8980 51.5970 ;
        RECT 11.7640 50.5035 11.7900 51.5970 ;
        RECT 11.6560 50.5035 11.6820 51.5970 ;
        RECT 11.5480 50.5035 11.5740 51.5970 ;
        RECT 11.4400 50.5035 11.4660 51.5970 ;
        RECT 11.3320 50.5035 11.3580 51.5970 ;
        RECT 11.2240 50.5035 11.2500 51.5970 ;
        RECT 11.1160 50.5035 11.1420 51.5970 ;
        RECT 11.0080 50.5035 11.0340 51.5970 ;
        RECT 10.9000 50.5035 10.9260 51.5970 ;
        RECT 10.7920 50.5035 10.8180 51.5970 ;
        RECT 10.6840 50.5035 10.7100 51.5970 ;
        RECT 10.5760 50.5035 10.6020 51.5970 ;
        RECT 10.4680 50.5035 10.4940 51.5970 ;
        RECT 10.3600 50.5035 10.3860 51.5970 ;
        RECT 10.2520 50.5035 10.2780 51.5970 ;
        RECT 10.1440 50.5035 10.1700 51.5970 ;
        RECT 10.0360 50.5035 10.0620 51.5970 ;
        RECT 9.9280 50.5035 9.9540 51.5970 ;
        RECT 9.8200 50.5035 9.8460 51.5970 ;
        RECT 9.7120 50.5035 9.7380 51.5970 ;
        RECT 9.6040 50.5035 9.6300 51.5970 ;
        RECT 9.4960 50.5035 9.5220 51.5970 ;
        RECT 9.3880 50.5035 9.4140 51.5970 ;
        RECT 9.1750 50.5035 9.2520 51.5970 ;
        RECT 7.2820 50.5035 7.3590 51.5970 ;
        RECT 7.1200 50.5035 7.1460 51.5970 ;
        RECT 7.0120 50.5035 7.0380 51.5970 ;
        RECT 6.9040 50.5035 6.9300 51.5970 ;
        RECT 6.7960 50.5035 6.8220 51.5970 ;
        RECT 6.6880 50.5035 6.7140 51.5970 ;
        RECT 6.5800 50.5035 6.6060 51.5970 ;
        RECT 6.4720 50.5035 6.4980 51.5970 ;
        RECT 6.3640 50.5035 6.3900 51.5970 ;
        RECT 6.2560 50.5035 6.2820 51.5970 ;
        RECT 6.1480 50.5035 6.1740 51.5970 ;
        RECT 6.0400 50.5035 6.0660 51.5970 ;
        RECT 5.9320 50.5035 5.9580 51.5970 ;
        RECT 5.8240 50.5035 5.8500 51.5970 ;
        RECT 5.7160 50.5035 5.7420 51.5970 ;
        RECT 5.6080 50.5035 5.6340 51.5970 ;
        RECT 5.5000 50.5035 5.5260 51.5970 ;
        RECT 5.3920 50.5035 5.4180 51.5970 ;
        RECT 5.2840 50.5035 5.3100 51.5970 ;
        RECT 5.1760 50.5035 5.2020 51.5970 ;
        RECT 5.0680 50.5035 5.0940 51.5970 ;
        RECT 4.9600 50.5035 4.9860 51.5970 ;
        RECT 4.8520 50.5035 4.8780 51.5970 ;
        RECT 4.7440 50.5035 4.7700 51.5970 ;
        RECT 4.6360 50.5035 4.6620 51.5970 ;
        RECT 4.5280 50.5035 4.5540 51.5970 ;
        RECT 4.4200 50.5035 4.4460 51.5970 ;
        RECT 4.3120 50.5035 4.3380 51.5970 ;
        RECT 4.2040 50.5035 4.2300 51.5970 ;
        RECT 4.0960 50.5035 4.1220 51.5970 ;
        RECT 3.9880 50.5035 4.0140 51.5970 ;
        RECT 3.8800 50.5035 3.9060 51.5970 ;
        RECT 3.7720 50.5035 3.7980 51.5970 ;
        RECT 3.6640 50.5035 3.6900 51.5970 ;
        RECT 3.5560 50.5035 3.5820 51.5970 ;
        RECT 3.4480 50.5035 3.4740 51.5970 ;
        RECT 3.3400 50.5035 3.3660 51.5970 ;
        RECT 3.2320 50.5035 3.2580 51.5970 ;
        RECT 3.1240 50.5035 3.1500 51.5970 ;
        RECT 3.0160 50.5035 3.0420 51.5970 ;
        RECT 2.9080 50.5035 2.9340 51.5970 ;
        RECT 2.8000 50.5035 2.8260 51.5970 ;
        RECT 2.6920 50.5035 2.7180 51.5970 ;
        RECT 2.5840 50.5035 2.6100 51.5970 ;
        RECT 2.4760 50.5035 2.5020 51.5970 ;
        RECT 2.3680 50.5035 2.3940 51.5970 ;
        RECT 2.2600 50.5035 2.2860 51.5970 ;
        RECT 2.1520 50.5035 2.1780 51.5970 ;
        RECT 2.0440 50.5035 2.0700 51.5970 ;
        RECT 1.9360 50.5035 1.9620 51.5970 ;
        RECT 1.8280 50.5035 1.8540 51.5970 ;
        RECT 1.7200 50.5035 1.7460 51.5970 ;
        RECT 1.6120 50.5035 1.6380 51.5970 ;
        RECT 1.5040 50.5035 1.5300 51.5970 ;
        RECT 1.3960 50.5035 1.4220 51.5970 ;
        RECT 1.2880 50.5035 1.3140 51.5970 ;
        RECT 1.1800 50.5035 1.2060 51.5970 ;
        RECT 1.0720 50.5035 1.0980 51.5970 ;
        RECT 0.9640 50.5035 0.9900 51.5970 ;
        RECT 0.8560 50.5035 0.8820 51.5970 ;
        RECT 0.7480 50.5035 0.7740 51.5970 ;
        RECT 0.6400 50.5035 0.6660 51.5970 ;
        RECT 0.5320 50.5035 0.5580 51.5970 ;
        RECT 0.4240 50.5035 0.4500 51.5970 ;
        RECT 0.3160 50.5035 0.3420 51.5970 ;
        RECT 0.2080 50.5035 0.2340 51.5970 ;
        RECT 0.0050 50.5035 0.0900 51.5970 ;
        RECT 8.6410 51.5835 8.7690 52.6770 ;
        RECT 8.6270 52.2490 8.7690 52.5715 ;
        RECT 8.4790 51.9760 8.5410 52.6770 ;
        RECT 8.4650 52.2855 8.5410 52.4390 ;
        RECT 8.4790 51.5835 8.5050 52.6770 ;
        RECT 8.4790 51.7045 8.5190 51.9440 ;
        RECT 8.4790 51.5835 8.5410 51.6725 ;
        RECT 8.1820 52.0340 8.3880 52.6770 ;
        RECT 8.3620 51.5835 8.3880 52.6770 ;
        RECT 8.1820 52.3110 8.4020 52.5690 ;
        RECT 8.1820 51.5835 8.2800 52.6770 ;
        RECT 7.7650 51.5835 7.8480 52.6770 ;
        RECT 7.7650 51.6720 7.8620 52.6075 ;
        RECT 16.4440 51.5835 16.5290 52.6770 ;
        RECT 16.3000 51.5835 16.3260 52.6770 ;
        RECT 16.1920 51.5835 16.2180 52.6770 ;
        RECT 16.0840 51.5835 16.1100 52.6770 ;
        RECT 15.9760 51.5835 16.0020 52.6770 ;
        RECT 15.8680 51.5835 15.8940 52.6770 ;
        RECT 15.7600 51.5835 15.7860 52.6770 ;
        RECT 15.6520 51.5835 15.6780 52.6770 ;
        RECT 15.5440 51.5835 15.5700 52.6770 ;
        RECT 15.4360 51.5835 15.4620 52.6770 ;
        RECT 15.3280 51.5835 15.3540 52.6770 ;
        RECT 15.2200 51.5835 15.2460 52.6770 ;
        RECT 15.1120 51.5835 15.1380 52.6770 ;
        RECT 15.0040 51.5835 15.0300 52.6770 ;
        RECT 14.8960 51.5835 14.9220 52.6770 ;
        RECT 14.7880 51.5835 14.8140 52.6770 ;
        RECT 14.6800 51.5835 14.7060 52.6770 ;
        RECT 14.5720 51.5835 14.5980 52.6770 ;
        RECT 14.4640 51.5835 14.4900 52.6770 ;
        RECT 14.3560 51.5835 14.3820 52.6770 ;
        RECT 14.2480 51.5835 14.2740 52.6770 ;
        RECT 14.1400 51.5835 14.1660 52.6770 ;
        RECT 14.0320 51.5835 14.0580 52.6770 ;
        RECT 13.9240 51.5835 13.9500 52.6770 ;
        RECT 13.8160 51.5835 13.8420 52.6770 ;
        RECT 13.7080 51.5835 13.7340 52.6770 ;
        RECT 13.6000 51.5835 13.6260 52.6770 ;
        RECT 13.4920 51.5835 13.5180 52.6770 ;
        RECT 13.3840 51.5835 13.4100 52.6770 ;
        RECT 13.2760 51.5835 13.3020 52.6770 ;
        RECT 13.1680 51.5835 13.1940 52.6770 ;
        RECT 13.0600 51.5835 13.0860 52.6770 ;
        RECT 12.9520 51.5835 12.9780 52.6770 ;
        RECT 12.8440 51.5835 12.8700 52.6770 ;
        RECT 12.7360 51.5835 12.7620 52.6770 ;
        RECT 12.6280 51.5835 12.6540 52.6770 ;
        RECT 12.5200 51.5835 12.5460 52.6770 ;
        RECT 12.4120 51.5835 12.4380 52.6770 ;
        RECT 12.3040 51.5835 12.3300 52.6770 ;
        RECT 12.1960 51.5835 12.2220 52.6770 ;
        RECT 12.0880 51.5835 12.1140 52.6770 ;
        RECT 11.9800 51.5835 12.0060 52.6770 ;
        RECT 11.8720 51.5835 11.8980 52.6770 ;
        RECT 11.7640 51.5835 11.7900 52.6770 ;
        RECT 11.6560 51.5835 11.6820 52.6770 ;
        RECT 11.5480 51.5835 11.5740 52.6770 ;
        RECT 11.4400 51.5835 11.4660 52.6770 ;
        RECT 11.3320 51.5835 11.3580 52.6770 ;
        RECT 11.2240 51.5835 11.2500 52.6770 ;
        RECT 11.1160 51.5835 11.1420 52.6770 ;
        RECT 11.0080 51.5835 11.0340 52.6770 ;
        RECT 10.9000 51.5835 10.9260 52.6770 ;
        RECT 10.7920 51.5835 10.8180 52.6770 ;
        RECT 10.6840 51.5835 10.7100 52.6770 ;
        RECT 10.5760 51.5835 10.6020 52.6770 ;
        RECT 10.4680 51.5835 10.4940 52.6770 ;
        RECT 10.3600 51.5835 10.3860 52.6770 ;
        RECT 10.2520 51.5835 10.2780 52.6770 ;
        RECT 10.1440 51.5835 10.1700 52.6770 ;
        RECT 10.0360 51.5835 10.0620 52.6770 ;
        RECT 9.9280 51.5835 9.9540 52.6770 ;
        RECT 9.8200 51.5835 9.8460 52.6770 ;
        RECT 9.7120 51.5835 9.7380 52.6770 ;
        RECT 9.6040 51.5835 9.6300 52.6770 ;
        RECT 9.4960 51.5835 9.5220 52.6770 ;
        RECT 9.3880 51.5835 9.4140 52.6770 ;
        RECT 9.1750 51.5835 9.2520 52.6770 ;
        RECT 7.2820 51.5835 7.3590 52.6770 ;
        RECT 7.1200 51.5835 7.1460 52.6770 ;
        RECT 7.0120 51.5835 7.0380 52.6770 ;
        RECT 6.9040 51.5835 6.9300 52.6770 ;
        RECT 6.7960 51.5835 6.8220 52.6770 ;
        RECT 6.6880 51.5835 6.7140 52.6770 ;
        RECT 6.5800 51.5835 6.6060 52.6770 ;
        RECT 6.4720 51.5835 6.4980 52.6770 ;
        RECT 6.3640 51.5835 6.3900 52.6770 ;
        RECT 6.2560 51.5835 6.2820 52.6770 ;
        RECT 6.1480 51.5835 6.1740 52.6770 ;
        RECT 6.0400 51.5835 6.0660 52.6770 ;
        RECT 5.9320 51.5835 5.9580 52.6770 ;
        RECT 5.8240 51.5835 5.8500 52.6770 ;
        RECT 5.7160 51.5835 5.7420 52.6770 ;
        RECT 5.6080 51.5835 5.6340 52.6770 ;
        RECT 5.5000 51.5835 5.5260 52.6770 ;
        RECT 5.3920 51.5835 5.4180 52.6770 ;
        RECT 5.2840 51.5835 5.3100 52.6770 ;
        RECT 5.1760 51.5835 5.2020 52.6770 ;
        RECT 5.0680 51.5835 5.0940 52.6770 ;
        RECT 4.9600 51.5835 4.9860 52.6770 ;
        RECT 4.8520 51.5835 4.8780 52.6770 ;
        RECT 4.7440 51.5835 4.7700 52.6770 ;
        RECT 4.6360 51.5835 4.6620 52.6770 ;
        RECT 4.5280 51.5835 4.5540 52.6770 ;
        RECT 4.4200 51.5835 4.4460 52.6770 ;
        RECT 4.3120 51.5835 4.3380 52.6770 ;
        RECT 4.2040 51.5835 4.2300 52.6770 ;
        RECT 4.0960 51.5835 4.1220 52.6770 ;
        RECT 3.9880 51.5835 4.0140 52.6770 ;
        RECT 3.8800 51.5835 3.9060 52.6770 ;
        RECT 3.7720 51.5835 3.7980 52.6770 ;
        RECT 3.6640 51.5835 3.6900 52.6770 ;
        RECT 3.5560 51.5835 3.5820 52.6770 ;
        RECT 3.4480 51.5835 3.4740 52.6770 ;
        RECT 3.3400 51.5835 3.3660 52.6770 ;
        RECT 3.2320 51.5835 3.2580 52.6770 ;
        RECT 3.1240 51.5835 3.1500 52.6770 ;
        RECT 3.0160 51.5835 3.0420 52.6770 ;
        RECT 2.9080 51.5835 2.9340 52.6770 ;
        RECT 2.8000 51.5835 2.8260 52.6770 ;
        RECT 2.6920 51.5835 2.7180 52.6770 ;
        RECT 2.5840 51.5835 2.6100 52.6770 ;
        RECT 2.4760 51.5835 2.5020 52.6770 ;
        RECT 2.3680 51.5835 2.3940 52.6770 ;
        RECT 2.2600 51.5835 2.2860 52.6770 ;
        RECT 2.1520 51.5835 2.1780 52.6770 ;
        RECT 2.0440 51.5835 2.0700 52.6770 ;
        RECT 1.9360 51.5835 1.9620 52.6770 ;
        RECT 1.8280 51.5835 1.8540 52.6770 ;
        RECT 1.7200 51.5835 1.7460 52.6770 ;
        RECT 1.6120 51.5835 1.6380 52.6770 ;
        RECT 1.5040 51.5835 1.5300 52.6770 ;
        RECT 1.3960 51.5835 1.4220 52.6770 ;
        RECT 1.2880 51.5835 1.3140 52.6770 ;
        RECT 1.1800 51.5835 1.2060 52.6770 ;
        RECT 1.0720 51.5835 1.0980 52.6770 ;
        RECT 0.9640 51.5835 0.9900 52.6770 ;
        RECT 0.8560 51.5835 0.8820 52.6770 ;
        RECT 0.7480 51.5835 0.7740 52.6770 ;
        RECT 0.6400 51.5835 0.6660 52.6770 ;
        RECT 0.5320 51.5835 0.5580 52.6770 ;
        RECT 0.4240 51.5835 0.4500 52.6770 ;
        RECT 0.3160 51.5835 0.3420 52.6770 ;
        RECT 0.2080 51.5835 0.2340 52.6770 ;
        RECT 0.0050 51.5835 0.0900 52.6770 ;
        RECT 8.6410 52.6635 8.7690 53.7570 ;
        RECT 8.6270 53.3290 8.7690 53.6515 ;
        RECT 8.4790 53.0560 8.5410 53.7570 ;
        RECT 8.4650 53.3655 8.5410 53.5190 ;
        RECT 8.4790 52.6635 8.5050 53.7570 ;
        RECT 8.4790 52.7845 8.5190 53.0240 ;
        RECT 8.4790 52.6635 8.5410 52.7525 ;
        RECT 8.1820 53.1140 8.3880 53.7570 ;
        RECT 8.3620 52.6635 8.3880 53.7570 ;
        RECT 8.1820 53.3910 8.4020 53.6490 ;
        RECT 8.1820 52.6635 8.2800 53.7570 ;
        RECT 7.7650 52.6635 7.8480 53.7570 ;
        RECT 7.7650 52.7520 7.8620 53.6875 ;
        RECT 16.4440 52.6635 16.5290 53.7570 ;
        RECT 16.3000 52.6635 16.3260 53.7570 ;
        RECT 16.1920 52.6635 16.2180 53.7570 ;
        RECT 16.0840 52.6635 16.1100 53.7570 ;
        RECT 15.9760 52.6635 16.0020 53.7570 ;
        RECT 15.8680 52.6635 15.8940 53.7570 ;
        RECT 15.7600 52.6635 15.7860 53.7570 ;
        RECT 15.6520 52.6635 15.6780 53.7570 ;
        RECT 15.5440 52.6635 15.5700 53.7570 ;
        RECT 15.4360 52.6635 15.4620 53.7570 ;
        RECT 15.3280 52.6635 15.3540 53.7570 ;
        RECT 15.2200 52.6635 15.2460 53.7570 ;
        RECT 15.1120 52.6635 15.1380 53.7570 ;
        RECT 15.0040 52.6635 15.0300 53.7570 ;
        RECT 14.8960 52.6635 14.9220 53.7570 ;
        RECT 14.7880 52.6635 14.8140 53.7570 ;
        RECT 14.6800 52.6635 14.7060 53.7570 ;
        RECT 14.5720 52.6635 14.5980 53.7570 ;
        RECT 14.4640 52.6635 14.4900 53.7570 ;
        RECT 14.3560 52.6635 14.3820 53.7570 ;
        RECT 14.2480 52.6635 14.2740 53.7570 ;
        RECT 14.1400 52.6635 14.1660 53.7570 ;
        RECT 14.0320 52.6635 14.0580 53.7570 ;
        RECT 13.9240 52.6635 13.9500 53.7570 ;
        RECT 13.8160 52.6635 13.8420 53.7570 ;
        RECT 13.7080 52.6635 13.7340 53.7570 ;
        RECT 13.6000 52.6635 13.6260 53.7570 ;
        RECT 13.4920 52.6635 13.5180 53.7570 ;
        RECT 13.3840 52.6635 13.4100 53.7570 ;
        RECT 13.2760 52.6635 13.3020 53.7570 ;
        RECT 13.1680 52.6635 13.1940 53.7570 ;
        RECT 13.0600 52.6635 13.0860 53.7570 ;
        RECT 12.9520 52.6635 12.9780 53.7570 ;
        RECT 12.8440 52.6635 12.8700 53.7570 ;
        RECT 12.7360 52.6635 12.7620 53.7570 ;
        RECT 12.6280 52.6635 12.6540 53.7570 ;
        RECT 12.5200 52.6635 12.5460 53.7570 ;
        RECT 12.4120 52.6635 12.4380 53.7570 ;
        RECT 12.3040 52.6635 12.3300 53.7570 ;
        RECT 12.1960 52.6635 12.2220 53.7570 ;
        RECT 12.0880 52.6635 12.1140 53.7570 ;
        RECT 11.9800 52.6635 12.0060 53.7570 ;
        RECT 11.8720 52.6635 11.8980 53.7570 ;
        RECT 11.7640 52.6635 11.7900 53.7570 ;
        RECT 11.6560 52.6635 11.6820 53.7570 ;
        RECT 11.5480 52.6635 11.5740 53.7570 ;
        RECT 11.4400 52.6635 11.4660 53.7570 ;
        RECT 11.3320 52.6635 11.3580 53.7570 ;
        RECT 11.2240 52.6635 11.2500 53.7570 ;
        RECT 11.1160 52.6635 11.1420 53.7570 ;
        RECT 11.0080 52.6635 11.0340 53.7570 ;
        RECT 10.9000 52.6635 10.9260 53.7570 ;
        RECT 10.7920 52.6635 10.8180 53.7570 ;
        RECT 10.6840 52.6635 10.7100 53.7570 ;
        RECT 10.5760 52.6635 10.6020 53.7570 ;
        RECT 10.4680 52.6635 10.4940 53.7570 ;
        RECT 10.3600 52.6635 10.3860 53.7570 ;
        RECT 10.2520 52.6635 10.2780 53.7570 ;
        RECT 10.1440 52.6635 10.1700 53.7570 ;
        RECT 10.0360 52.6635 10.0620 53.7570 ;
        RECT 9.9280 52.6635 9.9540 53.7570 ;
        RECT 9.8200 52.6635 9.8460 53.7570 ;
        RECT 9.7120 52.6635 9.7380 53.7570 ;
        RECT 9.6040 52.6635 9.6300 53.7570 ;
        RECT 9.4960 52.6635 9.5220 53.7570 ;
        RECT 9.3880 52.6635 9.4140 53.7570 ;
        RECT 9.1750 52.6635 9.2520 53.7570 ;
        RECT 7.2820 52.6635 7.3590 53.7570 ;
        RECT 7.1200 52.6635 7.1460 53.7570 ;
        RECT 7.0120 52.6635 7.0380 53.7570 ;
        RECT 6.9040 52.6635 6.9300 53.7570 ;
        RECT 6.7960 52.6635 6.8220 53.7570 ;
        RECT 6.6880 52.6635 6.7140 53.7570 ;
        RECT 6.5800 52.6635 6.6060 53.7570 ;
        RECT 6.4720 52.6635 6.4980 53.7570 ;
        RECT 6.3640 52.6635 6.3900 53.7570 ;
        RECT 6.2560 52.6635 6.2820 53.7570 ;
        RECT 6.1480 52.6635 6.1740 53.7570 ;
        RECT 6.0400 52.6635 6.0660 53.7570 ;
        RECT 5.9320 52.6635 5.9580 53.7570 ;
        RECT 5.8240 52.6635 5.8500 53.7570 ;
        RECT 5.7160 52.6635 5.7420 53.7570 ;
        RECT 5.6080 52.6635 5.6340 53.7570 ;
        RECT 5.5000 52.6635 5.5260 53.7570 ;
        RECT 5.3920 52.6635 5.4180 53.7570 ;
        RECT 5.2840 52.6635 5.3100 53.7570 ;
        RECT 5.1760 52.6635 5.2020 53.7570 ;
        RECT 5.0680 52.6635 5.0940 53.7570 ;
        RECT 4.9600 52.6635 4.9860 53.7570 ;
        RECT 4.8520 52.6635 4.8780 53.7570 ;
        RECT 4.7440 52.6635 4.7700 53.7570 ;
        RECT 4.6360 52.6635 4.6620 53.7570 ;
        RECT 4.5280 52.6635 4.5540 53.7570 ;
        RECT 4.4200 52.6635 4.4460 53.7570 ;
        RECT 4.3120 52.6635 4.3380 53.7570 ;
        RECT 4.2040 52.6635 4.2300 53.7570 ;
        RECT 4.0960 52.6635 4.1220 53.7570 ;
        RECT 3.9880 52.6635 4.0140 53.7570 ;
        RECT 3.8800 52.6635 3.9060 53.7570 ;
        RECT 3.7720 52.6635 3.7980 53.7570 ;
        RECT 3.6640 52.6635 3.6900 53.7570 ;
        RECT 3.5560 52.6635 3.5820 53.7570 ;
        RECT 3.4480 52.6635 3.4740 53.7570 ;
        RECT 3.3400 52.6635 3.3660 53.7570 ;
        RECT 3.2320 52.6635 3.2580 53.7570 ;
        RECT 3.1240 52.6635 3.1500 53.7570 ;
        RECT 3.0160 52.6635 3.0420 53.7570 ;
        RECT 2.9080 52.6635 2.9340 53.7570 ;
        RECT 2.8000 52.6635 2.8260 53.7570 ;
        RECT 2.6920 52.6635 2.7180 53.7570 ;
        RECT 2.5840 52.6635 2.6100 53.7570 ;
        RECT 2.4760 52.6635 2.5020 53.7570 ;
        RECT 2.3680 52.6635 2.3940 53.7570 ;
        RECT 2.2600 52.6635 2.2860 53.7570 ;
        RECT 2.1520 52.6635 2.1780 53.7570 ;
        RECT 2.0440 52.6635 2.0700 53.7570 ;
        RECT 1.9360 52.6635 1.9620 53.7570 ;
        RECT 1.8280 52.6635 1.8540 53.7570 ;
        RECT 1.7200 52.6635 1.7460 53.7570 ;
        RECT 1.6120 52.6635 1.6380 53.7570 ;
        RECT 1.5040 52.6635 1.5300 53.7570 ;
        RECT 1.3960 52.6635 1.4220 53.7570 ;
        RECT 1.2880 52.6635 1.3140 53.7570 ;
        RECT 1.1800 52.6635 1.2060 53.7570 ;
        RECT 1.0720 52.6635 1.0980 53.7570 ;
        RECT 0.9640 52.6635 0.9900 53.7570 ;
        RECT 0.8560 52.6635 0.8820 53.7570 ;
        RECT 0.7480 52.6635 0.7740 53.7570 ;
        RECT 0.6400 52.6635 0.6660 53.7570 ;
        RECT 0.5320 52.6635 0.5580 53.7570 ;
        RECT 0.4240 52.6635 0.4500 53.7570 ;
        RECT 0.3160 52.6635 0.3420 53.7570 ;
        RECT 0.2080 52.6635 0.2340 53.7570 ;
        RECT 0.0050 52.6635 0.0900 53.7570 ;
        RECT 8.6410 53.7435 8.7690 54.8370 ;
        RECT 8.6270 54.4090 8.7690 54.7315 ;
        RECT 8.4790 54.1360 8.5410 54.8370 ;
        RECT 8.4650 54.4455 8.5410 54.5990 ;
        RECT 8.4790 53.7435 8.5050 54.8370 ;
        RECT 8.4790 53.8645 8.5190 54.1040 ;
        RECT 8.4790 53.7435 8.5410 53.8325 ;
        RECT 8.1820 54.1940 8.3880 54.8370 ;
        RECT 8.3620 53.7435 8.3880 54.8370 ;
        RECT 8.1820 54.4710 8.4020 54.7290 ;
        RECT 8.1820 53.7435 8.2800 54.8370 ;
        RECT 7.7650 53.7435 7.8480 54.8370 ;
        RECT 7.7650 53.8320 7.8620 54.7675 ;
        RECT 16.4440 53.7435 16.5290 54.8370 ;
        RECT 16.3000 53.7435 16.3260 54.8370 ;
        RECT 16.1920 53.7435 16.2180 54.8370 ;
        RECT 16.0840 53.7435 16.1100 54.8370 ;
        RECT 15.9760 53.7435 16.0020 54.8370 ;
        RECT 15.8680 53.7435 15.8940 54.8370 ;
        RECT 15.7600 53.7435 15.7860 54.8370 ;
        RECT 15.6520 53.7435 15.6780 54.8370 ;
        RECT 15.5440 53.7435 15.5700 54.8370 ;
        RECT 15.4360 53.7435 15.4620 54.8370 ;
        RECT 15.3280 53.7435 15.3540 54.8370 ;
        RECT 15.2200 53.7435 15.2460 54.8370 ;
        RECT 15.1120 53.7435 15.1380 54.8370 ;
        RECT 15.0040 53.7435 15.0300 54.8370 ;
        RECT 14.8960 53.7435 14.9220 54.8370 ;
        RECT 14.7880 53.7435 14.8140 54.8370 ;
        RECT 14.6800 53.7435 14.7060 54.8370 ;
        RECT 14.5720 53.7435 14.5980 54.8370 ;
        RECT 14.4640 53.7435 14.4900 54.8370 ;
        RECT 14.3560 53.7435 14.3820 54.8370 ;
        RECT 14.2480 53.7435 14.2740 54.8370 ;
        RECT 14.1400 53.7435 14.1660 54.8370 ;
        RECT 14.0320 53.7435 14.0580 54.8370 ;
        RECT 13.9240 53.7435 13.9500 54.8370 ;
        RECT 13.8160 53.7435 13.8420 54.8370 ;
        RECT 13.7080 53.7435 13.7340 54.8370 ;
        RECT 13.6000 53.7435 13.6260 54.8370 ;
        RECT 13.4920 53.7435 13.5180 54.8370 ;
        RECT 13.3840 53.7435 13.4100 54.8370 ;
        RECT 13.2760 53.7435 13.3020 54.8370 ;
        RECT 13.1680 53.7435 13.1940 54.8370 ;
        RECT 13.0600 53.7435 13.0860 54.8370 ;
        RECT 12.9520 53.7435 12.9780 54.8370 ;
        RECT 12.8440 53.7435 12.8700 54.8370 ;
        RECT 12.7360 53.7435 12.7620 54.8370 ;
        RECT 12.6280 53.7435 12.6540 54.8370 ;
        RECT 12.5200 53.7435 12.5460 54.8370 ;
        RECT 12.4120 53.7435 12.4380 54.8370 ;
        RECT 12.3040 53.7435 12.3300 54.8370 ;
        RECT 12.1960 53.7435 12.2220 54.8370 ;
        RECT 12.0880 53.7435 12.1140 54.8370 ;
        RECT 11.9800 53.7435 12.0060 54.8370 ;
        RECT 11.8720 53.7435 11.8980 54.8370 ;
        RECT 11.7640 53.7435 11.7900 54.8370 ;
        RECT 11.6560 53.7435 11.6820 54.8370 ;
        RECT 11.5480 53.7435 11.5740 54.8370 ;
        RECT 11.4400 53.7435 11.4660 54.8370 ;
        RECT 11.3320 53.7435 11.3580 54.8370 ;
        RECT 11.2240 53.7435 11.2500 54.8370 ;
        RECT 11.1160 53.7435 11.1420 54.8370 ;
        RECT 11.0080 53.7435 11.0340 54.8370 ;
        RECT 10.9000 53.7435 10.9260 54.8370 ;
        RECT 10.7920 53.7435 10.8180 54.8370 ;
        RECT 10.6840 53.7435 10.7100 54.8370 ;
        RECT 10.5760 53.7435 10.6020 54.8370 ;
        RECT 10.4680 53.7435 10.4940 54.8370 ;
        RECT 10.3600 53.7435 10.3860 54.8370 ;
        RECT 10.2520 53.7435 10.2780 54.8370 ;
        RECT 10.1440 53.7435 10.1700 54.8370 ;
        RECT 10.0360 53.7435 10.0620 54.8370 ;
        RECT 9.9280 53.7435 9.9540 54.8370 ;
        RECT 9.8200 53.7435 9.8460 54.8370 ;
        RECT 9.7120 53.7435 9.7380 54.8370 ;
        RECT 9.6040 53.7435 9.6300 54.8370 ;
        RECT 9.4960 53.7435 9.5220 54.8370 ;
        RECT 9.3880 53.7435 9.4140 54.8370 ;
        RECT 9.1750 53.7435 9.2520 54.8370 ;
        RECT 7.2820 53.7435 7.3590 54.8370 ;
        RECT 7.1200 53.7435 7.1460 54.8370 ;
        RECT 7.0120 53.7435 7.0380 54.8370 ;
        RECT 6.9040 53.7435 6.9300 54.8370 ;
        RECT 6.7960 53.7435 6.8220 54.8370 ;
        RECT 6.6880 53.7435 6.7140 54.8370 ;
        RECT 6.5800 53.7435 6.6060 54.8370 ;
        RECT 6.4720 53.7435 6.4980 54.8370 ;
        RECT 6.3640 53.7435 6.3900 54.8370 ;
        RECT 6.2560 53.7435 6.2820 54.8370 ;
        RECT 6.1480 53.7435 6.1740 54.8370 ;
        RECT 6.0400 53.7435 6.0660 54.8370 ;
        RECT 5.9320 53.7435 5.9580 54.8370 ;
        RECT 5.8240 53.7435 5.8500 54.8370 ;
        RECT 5.7160 53.7435 5.7420 54.8370 ;
        RECT 5.6080 53.7435 5.6340 54.8370 ;
        RECT 5.5000 53.7435 5.5260 54.8370 ;
        RECT 5.3920 53.7435 5.4180 54.8370 ;
        RECT 5.2840 53.7435 5.3100 54.8370 ;
        RECT 5.1760 53.7435 5.2020 54.8370 ;
        RECT 5.0680 53.7435 5.0940 54.8370 ;
        RECT 4.9600 53.7435 4.9860 54.8370 ;
        RECT 4.8520 53.7435 4.8780 54.8370 ;
        RECT 4.7440 53.7435 4.7700 54.8370 ;
        RECT 4.6360 53.7435 4.6620 54.8370 ;
        RECT 4.5280 53.7435 4.5540 54.8370 ;
        RECT 4.4200 53.7435 4.4460 54.8370 ;
        RECT 4.3120 53.7435 4.3380 54.8370 ;
        RECT 4.2040 53.7435 4.2300 54.8370 ;
        RECT 4.0960 53.7435 4.1220 54.8370 ;
        RECT 3.9880 53.7435 4.0140 54.8370 ;
        RECT 3.8800 53.7435 3.9060 54.8370 ;
        RECT 3.7720 53.7435 3.7980 54.8370 ;
        RECT 3.6640 53.7435 3.6900 54.8370 ;
        RECT 3.5560 53.7435 3.5820 54.8370 ;
        RECT 3.4480 53.7435 3.4740 54.8370 ;
        RECT 3.3400 53.7435 3.3660 54.8370 ;
        RECT 3.2320 53.7435 3.2580 54.8370 ;
        RECT 3.1240 53.7435 3.1500 54.8370 ;
        RECT 3.0160 53.7435 3.0420 54.8370 ;
        RECT 2.9080 53.7435 2.9340 54.8370 ;
        RECT 2.8000 53.7435 2.8260 54.8370 ;
        RECT 2.6920 53.7435 2.7180 54.8370 ;
        RECT 2.5840 53.7435 2.6100 54.8370 ;
        RECT 2.4760 53.7435 2.5020 54.8370 ;
        RECT 2.3680 53.7435 2.3940 54.8370 ;
        RECT 2.2600 53.7435 2.2860 54.8370 ;
        RECT 2.1520 53.7435 2.1780 54.8370 ;
        RECT 2.0440 53.7435 2.0700 54.8370 ;
        RECT 1.9360 53.7435 1.9620 54.8370 ;
        RECT 1.8280 53.7435 1.8540 54.8370 ;
        RECT 1.7200 53.7435 1.7460 54.8370 ;
        RECT 1.6120 53.7435 1.6380 54.8370 ;
        RECT 1.5040 53.7435 1.5300 54.8370 ;
        RECT 1.3960 53.7435 1.4220 54.8370 ;
        RECT 1.2880 53.7435 1.3140 54.8370 ;
        RECT 1.1800 53.7435 1.2060 54.8370 ;
        RECT 1.0720 53.7435 1.0980 54.8370 ;
        RECT 0.9640 53.7435 0.9900 54.8370 ;
        RECT 0.8560 53.7435 0.8820 54.8370 ;
        RECT 0.7480 53.7435 0.7740 54.8370 ;
        RECT 0.6400 53.7435 0.6660 54.8370 ;
        RECT 0.5320 53.7435 0.5580 54.8370 ;
        RECT 0.4240 53.7435 0.4500 54.8370 ;
        RECT 0.3160 53.7435 0.3420 54.8370 ;
        RECT 0.2080 53.7435 0.2340 54.8370 ;
        RECT 0.0050 53.7435 0.0900 54.8370 ;
        RECT 8.6410 54.8235 8.7690 55.9170 ;
        RECT 8.6270 55.4890 8.7690 55.8115 ;
        RECT 8.4790 55.2160 8.5410 55.9170 ;
        RECT 8.4650 55.5255 8.5410 55.6790 ;
        RECT 8.4790 54.8235 8.5050 55.9170 ;
        RECT 8.4790 54.9445 8.5190 55.1840 ;
        RECT 8.4790 54.8235 8.5410 54.9125 ;
        RECT 8.1820 55.2740 8.3880 55.9170 ;
        RECT 8.3620 54.8235 8.3880 55.9170 ;
        RECT 8.1820 55.5510 8.4020 55.8090 ;
        RECT 8.1820 54.8235 8.2800 55.9170 ;
        RECT 7.7650 54.8235 7.8480 55.9170 ;
        RECT 7.7650 54.9120 7.8620 55.8475 ;
        RECT 16.4440 54.8235 16.5290 55.9170 ;
        RECT 16.3000 54.8235 16.3260 55.9170 ;
        RECT 16.1920 54.8235 16.2180 55.9170 ;
        RECT 16.0840 54.8235 16.1100 55.9170 ;
        RECT 15.9760 54.8235 16.0020 55.9170 ;
        RECT 15.8680 54.8235 15.8940 55.9170 ;
        RECT 15.7600 54.8235 15.7860 55.9170 ;
        RECT 15.6520 54.8235 15.6780 55.9170 ;
        RECT 15.5440 54.8235 15.5700 55.9170 ;
        RECT 15.4360 54.8235 15.4620 55.9170 ;
        RECT 15.3280 54.8235 15.3540 55.9170 ;
        RECT 15.2200 54.8235 15.2460 55.9170 ;
        RECT 15.1120 54.8235 15.1380 55.9170 ;
        RECT 15.0040 54.8235 15.0300 55.9170 ;
        RECT 14.8960 54.8235 14.9220 55.9170 ;
        RECT 14.7880 54.8235 14.8140 55.9170 ;
        RECT 14.6800 54.8235 14.7060 55.9170 ;
        RECT 14.5720 54.8235 14.5980 55.9170 ;
        RECT 14.4640 54.8235 14.4900 55.9170 ;
        RECT 14.3560 54.8235 14.3820 55.9170 ;
        RECT 14.2480 54.8235 14.2740 55.9170 ;
        RECT 14.1400 54.8235 14.1660 55.9170 ;
        RECT 14.0320 54.8235 14.0580 55.9170 ;
        RECT 13.9240 54.8235 13.9500 55.9170 ;
        RECT 13.8160 54.8235 13.8420 55.9170 ;
        RECT 13.7080 54.8235 13.7340 55.9170 ;
        RECT 13.6000 54.8235 13.6260 55.9170 ;
        RECT 13.4920 54.8235 13.5180 55.9170 ;
        RECT 13.3840 54.8235 13.4100 55.9170 ;
        RECT 13.2760 54.8235 13.3020 55.9170 ;
        RECT 13.1680 54.8235 13.1940 55.9170 ;
        RECT 13.0600 54.8235 13.0860 55.9170 ;
        RECT 12.9520 54.8235 12.9780 55.9170 ;
        RECT 12.8440 54.8235 12.8700 55.9170 ;
        RECT 12.7360 54.8235 12.7620 55.9170 ;
        RECT 12.6280 54.8235 12.6540 55.9170 ;
        RECT 12.5200 54.8235 12.5460 55.9170 ;
        RECT 12.4120 54.8235 12.4380 55.9170 ;
        RECT 12.3040 54.8235 12.3300 55.9170 ;
        RECT 12.1960 54.8235 12.2220 55.9170 ;
        RECT 12.0880 54.8235 12.1140 55.9170 ;
        RECT 11.9800 54.8235 12.0060 55.9170 ;
        RECT 11.8720 54.8235 11.8980 55.9170 ;
        RECT 11.7640 54.8235 11.7900 55.9170 ;
        RECT 11.6560 54.8235 11.6820 55.9170 ;
        RECT 11.5480 54.8235 11.5740 55.9170 ;
        RECT 11.4400 54.8235 11.4660 55.9170 ;
        RECT 11.3320 54.8235 11.3580 55.9170 ;
        RECT 11.2240 54.8235 11.2500 55.9170 ;
        RECT 11.1160 54.8235 11.1420 55.9170 ;
        RECT 11.0080 54.8235 11.0340 55.9170 ;
        RECT 10.9000 54.8235 10.9260 55.9170 ;
        RECT 10.7920 54.8235 10.8180 55.9170 ;
        RECT 10.6840 54.8235 10.7100 55.9170 ;
        RECT 10.5760 54.8235 10.6020 55.9170 ;
        RECT 10.4680 54.8235 10.4940 55.9170 ;
        RECT 10.3600 54.8235 10.3860 55.9170 ;
        RECT 10.2520 54.8235 10.2780 55.9170 ;
        RECT 10.1440 54.8235 10.1700 55.9170 ;
        RECT 10.0360 54.8235 10.0620 55.9170 ;
        RECT 9.9280 54.8235 9.9540 55.9170 ;
        RECT 9.8200 54.8235 9.8460 55.9170 ;
        RECT 9.7120 54.8235 9.7380 55.9170 ;
        RECT 9.6040 54.8235 9.6300 55.9170 ;
        RECT 9.4960 54.8235 9.5220 55.9170 ;
        RECT 9.3880 54.8235 9.4140 55.9170 ;
        RECT 9.1750 54.8235 9.2520 55.9170 ;
        RECT 7.2820 54.8235 7.3590 55.9170 ;
        RECT 7.1200 54.8235 7.1460 55.9170 ;
        RECT 7.0120 54.8235 7.0380 55.9170 ;
        RECT 6.9040 54.8235 6.9300 55.9170 ;
        RECT 6.7960 54.8235 6.8220 55.9170 ;
        RECT 6.6880 54.8235 6.7140 55.9170 ;
        RECT 6.5800 54.8235 6.6060 55.9170 ;
        RECT 6.4720 54.8235 6.4980 55.9170 ;
        RECT 6.3640 54.8235 6.3900 55.9170 ;
        RECT 6.2560 54.8235 6.2820 55.9170 ;
        RECT 6.1480 54.8235 6.1740 55.9170 ;
        RECT 6.0400 54.8235 6.0660 55.9170 ;
        RECT 5.9320 54.8235 5.9580 55.9170 ;
        RECT 5.8240 54.8235 5.8500 55.9170 ;
        RECT 5.7160 54.8235 5.7420 55.9170 ;
        RECT 5.6080 54.8235 5.6340 55.9170 ;
        RECT 5.5000 54.8235 5.5260 55.9170 ;
        RECT 5.3920 54.8235 5.4180 55.9170 ;
        RECT 5.2840 54.8235 5.3100 55.9170 ;
        RECT 5.1760 54.8235 5.2020 55.9170 ;
        RECT 5.0680 54.8235 5.0940 55.9170 ;
        RECT 4.9600 54.8235 4.9860 55.9170 ;
        RECT 4.8520 54.8235 4.8780 55.9170 ;
        RECT 4.7440 54.8235 4.7700 55.9170 ;
        RECT 4.6360 54.8235 4.6620 55.9170 ;
        RECT 4.5280 54.8235 4.5540 55.9170 ;
        RECT 4.4200 54.8235 4.4460 55.9170 ;
        RECT 4.3120 54.8235 4.3380 55.9170 ;
        RECT 4.2040 54.8235 4.2300 55.9170 ;
        RECT 4.0960 54.8235 4.1220 55.9170 ;
        RECT 3.9880 54.8235 4.0140 55.9170 ;
        RECT 3.8800 54.8235 3.9060 55.9170 ;
        RECT 3.7720 54.8235 3.7980 55.9170 ;
        RECT 3.6640 54.8235 3.6900 55.9170 ;
        RECT 3.5560 54.8235 3.5820 55.9170 ;
        RECT 3.4480 54.8235 3.4740 55.9170 ;
        RECT 3.3400 54.8235 3.3660 55.9170 ;
        RECT 3.2320 54.8235 3.2580 55.9170 ;
        RECT 3.1240 54.8235 3.1500 55.9170 ;
        RECT 3.0160 54.8235 3.0420 55.9170 ;
        RECT 2.9080 54.8235 2.9340 55.9170 ;
        RECT 2.8000 54.8235 2.8260 55.9170 ;
        RECT 2.6920 54.8235 2.7180 55.9170 ;
        RECT 2.5840 54.8235 2.6100 55.9170 ;
        RECT 2.4760 54.8235 2.5020 55.9170 ;
        RECT 2.3680 54.8235 2.3940 55.9170 ;
        RECT 2.2600 54.8235 2.2860 55.9170 ;
        RECT 2.1520 54.8235 2.1780 55.9170 ;
        RECT 2.0440 54.8235 2.0700 55.9170 ;
        RECT 1.9360 54.8235 1.9620 55.9170 ;
        RECT 1.8280 54.8235 1.8540 55.9170 ;
        RECT 1.7200 54.8235 1.7460 55.9170 ;
        RECT 1.6120 54.8235 1.6380 55.9170 ;
        RECT 1.5040 54.8235 1.5300 55.9170 ;
        RECT 1.3960 54.8235 1.4220 55.9170 ;
        RECT 1.2880 54.8235 1.3140 55.9170 ;
        RECT 1.1800 54.8235 1.2060 55.9170 ;
        RECT 1.0720 54.8235 1.0980 55.9170 ;
        RECT 0.9640 54.8235 0.9900 55.9170 ;
        RECT 0.8560 54.8235 0.8820 55.9170 ;
        RECT 0.7480 54.8235 0.7740 55.9170 ;
        RECT 0.6400 54.8235 0.6660 55.9170 ;
        RECT 0.5320 54.8235 0.5580 55.9170 ;
        RECT 0.4240 54.8235 0.4500 55.9170 ;
        RECT 0.3160 54.8235 0.3420 55.9170 ;
        RECT 0.2080 54.8235 0.2340 55.9170 ;
        RECT 0.0050 54.8235 0.0900 55.9170 ;
        RECT 8.6410 55.9035 8.7690 56.9970 ;
        RECT 8.6270 56.5690 8.7690 56.8915 ;
        RECT 8.4790 56.2960 8.5410 56.9970 ;
        RECT 8.4650 56.6055 8.5410 56.7590 ;
        RECT 8.4790 55.9035 8.5050 56.9970 ;
        RECT 8.4790 56.0245 8.5190 56.2640 ;
        RECT 8.4790 55.9035 8.5410 55.9925 ;
        RECT 8.1820 56.3540 8.3880 56.9970 ;
        RECT 8.3620 55.9035 8.3880 56.9970 ;
        RECT 8.1820 56.6310 8.4020 56.8890 ;
        RECT 8.1820 55.9035 8.2800 56.9970 ;
        RECT 7.7650 55.9035 7.8480 56.9970 ;
        RECT 7.7650 55.9920 7.8620 56.9275 ;
        RECT 16.4440 55.9035 16.5290 56.9970 ;
        RECT 16.3000 55.9035 16.3260 56.9970 ;
        RECT 16.1920 55.9035 16.2180 56.9970 ;
        RECT 16.0840 55.9035 16.1100 56.9970 ;
        RECT 15.9760 55.9035 16.0020 56.9970 ;
        RECT 15.8680 55.9035 15.8940 56.9970 ;
        RECT 15.7600 55.9035 15.7860 56.9970 ;
        RECT 15.6520 55.9035 15.6780 56.9970 ;
        RECT 15.5440 55.9035 15.5700 56.9970 ;
        RECT 15.4360 55.9035 15.4620 56.9970 ;
        RECT 15.3280 55.9035 15.3540 56.9970 ;
        RECT 15.2200 55.9035 15.2460 56.9970 ;
        RECT 15.1120 55.9035 15.1380 56.9970 ;
        RECT 15.0040 55.9035 15.0300 56.9970 ;
        RECT 14.8960 55.9035 14.9220 56.9970 ;
        RECT 14.7880 55.9035 14.8140 56.9970 ;
        RECT 14.6800 55.9035 14.7060 56.9970 ;
        RECT 14.5720 55.9035 14.5980 56.9970 ;
        RECT 14.4640 55.9035 14.4900 56.9970 ;
        RECT 14.3560 55.9035 14.3820 56.9970 ;
        RECT 14.2480 55.9035 14.2740 56.9970 ;
        RECT 14.1400 55.9035 14.1660 56.9970 ;
        RECT 14.0320 55.9035 14.0580 56.9970 ;
        RECT 13.9240 55.9035 13.9500 56.9970 ;
        RECT 13.8160 55.9035 13.8420 56.9970 ;
        RECT 13.7080 55.9035 13.7340 56.9970 ;
        RECT 13.6000 55.9035 13.6260 56.9970 ;
        RECT 13.4920 55.9035 13.5180 56.9970 ;
        RECT 13.3840 55.9035 13.4100 56.9970 ;
        RECT 13.2760 55.9035 13.3020 56.9970 ;
        RECT 13.1680 55.9035 13.1940 56.9970 ;
        RECT 13.0600 55.9035 13.0860 56.9970 ;
        RECT 12.9520 55.9035 12.9780 56.9970 ;
        RECT 12.8440 55.9035 12.8700 56.9970 ;
        RECT 12.7360 55.9035 12.7620 56.9970 ;
        RECT 12.6280 55.9035 12.6540 56.9970 ;
        RECT 12.5200 55.9035 12.5460 56.9970 ;
        RECT 12.4120 55.9035 12.4380 56.9970 ;
        RECT 12.3040 55.9035 12.3300 56.9970 ;
        RECT 12.1960 55.9035 12.2220 56.9970 ;
        RECT 12.0880 55.9035 12.1140 56.9970 ;
        RECT 11.9800 55.9035 12.0060 56.9970 ;
        RECT 11.8720 55.9035 11.8980 56.9970 ;
        RECT 11.7640 55.9035 11.7900 56.9970 ;
        RECT 11.6560 55.9035 11.6820 56.9970 ;
        RECT 11.5480 55.9035 11.5740 56.9970 ;
        RECT 11.4400 55.9035 11.4660 56.9970 ;
        RECT 11.3320 55.9035 11.3580 56.9970 ;
        RECT 11.2240 55.9035 11.2500 56.9970 ;
        RECT 11.1160 55.9035 11.1420 56.9970 ;
        RECT 11.0080 55.9035 11.0340 56.9970 ;
        RECT 10.9000 55.9035 10.9260 56.9970 ;
        RECT 10.7920 55.9035 10.8180 56.9970 ;
        RECT 10.6840 55.9035 10.7100 56.9970 ;
        RECT 10.5760 55.9035 10.6020 56.9970 ;
        RECT 10.4680 55.9035 10.4940 56.9970 ;
        RECT 10.3600 55.9035 10.3860 56.9970 ;
        RECT 10.2520 55.9035 10.2780 56.9970 ;
        RECT 10.1440 55.9035 10.1700 56.9970 ;
        RECT 10.0360 55.9035 10.0620 56.9970 ;
        RECT 9.9280 55.9035 9.9540 56.9970 ;
        RECT 9.8200 55.9035 9.8460 56.9970 ;
        RECT 9.7120 55.9035 9.7380 56.9970 ;
        RECT 9.6040 55.9035 9.6300 56.9970 ;
        RECT 9.4960 55.9035 9.5220 56.9970 ;
        RECT 9.3880 55.9035 9.4140 56.9970 ;
        RECT 9.1750 55.9035 9.2520 56.9970 ;
        RECT 7.2820 55.9035 7.3590 56.9970 ;
        RECT 7.1200 55.9035 7.1460 56.9970 ;
        RECT 7.0120 55.9035 7.0380 56.9970 ;
        RECT 6.9040 55.9035 6.9300 56.9970 ;
        RECT 6.7960 55.9035 6.8220 56.9970 ;
        RECT 6.6880 55.9035 6.7140 56.9970 ;
        RECT 6.5800 55.9035 6.6060 56.9970 ;
        RECT 6.4720 55.9035 6.4980 56.9970 ;
        RECT 6.3640 55.9035 6.3900 56.9970 ;
        RECT 6.2560 55.9035 6.2820 56.9970 ;
        RECT 6.1480 55.9035 6.1740 56.9970 ;
        RECT 6.0400 55.9035 6.0660 56.9970 ;
        RECT 5.9320 55.9035 5.9580 56.9970 ;
        RECT 5.8240 55.9035 5.8500 56.9970 ;
        RECT 5.7160 55.9035 5.7420 56.9970 ;
        RECT 5.6080 55.9035 5.6340 56.9970 ;
        RECT 5.5000 55.9035 5.5260 56.9970 ;
        RECT 5.3920 55.9035 5.4180 56.9970 ;
        RECT 5.2840 55.9035 5.3100 56.9970 ;
        RECT 5.1760 55.9035 5.2020 56.9970 ;
        RECT 5.0680 55.9035 5.0940 56.9970 ;
        RECT 4.9600 55.9035 4.9860 56.9970 ;
        RECT 4.8520 55.9035 4.8780 56.9970 ;
        RECT 4.7440 55.9035 4.7700 56.9970 ;
        RECT 4.6360 55.9035 4.6620 56.9970 ;
        RECT 4.5280 55.9035 4.5540 56.9970 ;
        RECT 4.4200 55.9035 4.4460 56.9970 ;
        RECT 4.3120 55.9035 4.3380 56.9970 ;
        RECT 4.2040 55.9035 4.2300 56.9970 ;
        RECT 4.0960 55.9035 4.1220 56.9970 ;
        RECT 3.9880 55.9035 4.0140 56.9970 ;
        RECT 3.8800 55.9035 3.9060 56.9970 ;
        RECT 3.7720 55.9035 3.7980 56.9970 ;
        RECT 3.6640 55.9035 3.6900 56.9970 ;
        RECT 3.5560 55.9035 3.5820 56.9970 ;
        RECT 3.4480 55.9035 3.4740 56.9970 ;
        RECT 3.3400 55.9035 3.3660 56.9970 ;
        RECT 3.2320 55.9035 3.2580 56.9970 ;
        RECT 3.1240 55.9035 3.1500 56.9970 ;
        RECT 3.0160 55.9035 3.0420 56.9970 ;
        RECT 2.9080 55.9035 2.9340 56.9970 ;
        RECT 2.8000 55.9035 2.8260 56.9970 ;
        RECT 2.6920 55.9035 2.7180 56.9970 ;
        RECT 2.5840 55.9035 2.6100 56.9970 ;
        RECT 2.4760 55.9035 2.5020 56.9970 ;
        RECT 2.3680 55.9035 2.3940 56.9970 ;
        RECT 2.2600 55.9035 2.2860 56.9970 ;
        RECT 2.1520 55.9035 2.1780 56.9970 ;
        RECT 2.0440 55.9035 2.0700 56.9970 ;
        RECT 1.9360 55.9035 1.9620 56.9970 ;
        RECT 1.8280 55.9035 1.8540 56.9970 ;
        RECT 1.7200 55.9035 1.7460 56.9970 ;
        RECT 1.6120 55.9035 1.6380 56.9970 ;
        RECT 1.5040 55.9035 1.5300 56.9970 ;
        RECT 1.3960 55.9035 1.4220 56.9970 ;
        RECT 1.2880 55.9035 1.3140 56.9970 ;
        RECT 1.1800 55.9035 1.2060 56.9970 ;
        RECT 1.0720 55.9035 1.0980 56.9970 ;
        RECT 0.9640 55.9035 0.9900 56.9970 ;
        RECT 0.8560 55.9035 0.8820 56.9970 ;
        RECT 0.7480 55.9035 0.7740 56.9970 ;
        RECT 0.6400 55.9035 0.6660 56.9970 ;
        RECT 0.5320 55.9035 0.5580 56.9970 ;
        RECT 0.4240 55.9035 0.4500 56.9970 ;
        RECT 0.3160 55.9035 0.3420 56.9970 ;
        RECT 0.2080 55.9035 0.2340 56.9970 ;
        RECT 0.0050 55.9035 0.0900 56.9970 ;
        RECT 8.6410 56.9835 8.7690 58.0770 ;
        RECT 8.6270 57.6490 8.7690 57.9715 ;
        RECT 8.4790 57.3760 8.5410 58.0770 ;
        RECT 8.4650 57.6855 8.5410 57.8390 ;
        RECT 8.4790 56.9835 8.5050 58.0770 ;
        RECT 8.4790 57.1045 8.5190 57.3440 ;
        RECT 8.4790 56.9835 8.5410 57.0725 ;
        RECT 8.1820 57.4340 8.3880 58.0770 ;
        RECT 8.3620 56.9835 8.3880 58.0770 ;
        RECT 8.1820 57.7110 8.4020 57.9690 ;
        RECT 8.1820 56.9835 8.2800 58.0770 ;
        RECT 7.7650 56.9835 7.8480 58.0770 ;
        RECT 7.7650 57.0720 7.8620 58.0075 ;
        RECT 16.4440 56.9835 16.5290 58.0770 ;
        RECT 16.3000 56.9835 16.3260 58.0770 ;
        RECT 16.1920 56.9835 16.2180 58.0770 ;
        RECT 16.0840 56.9835 16.1100 58.0770 ;
        RECT 15.9760 56.9835 16.0020 58.0770 ;
        RECT 15.8680 56.9835 15.8940 58.0770 ;
        RECT 15.7600 56.9835 15.7860 58.0770 ;
        RECT 15.6520 56.9835 15.6780 58.0770 ;
        RECT 15.5440 56.9835 15.5700 58.0770 ;
        RECT 15.4360 56.9835 15.4620 58.0770 ;
        RECT 15.3280 56.9835 15.3540 58.0770 ;
        RECT 15.2200 56.9835 15.2460 58.0770 ;
        RECT 15.1120 56.9835 15.1380 58.0770 ;
        RECT 15.0040 56.9835 15.0300 58.0770 ;
        RECT 14.8960 56.9835 14.9220 58.0770 ;
        RECT 14.7880 56.9835 14.8140 58.0770 ;
        RECT 14.6800 56.9835 14.7060 58.0770 ;
        RECT 14.5720 56.9835 14.5980 58.0770 ;
        RECT 14.4640 56.9835 14.4900 58.0770 ;
        RECT 14.3560 56.9835 14.3820 58.0770 ;
        RECT 14.2480 56.9835 14.2740 58.0770 ;
        RECT 14.1400 56.9835 14.1660 58.0770 ;
        RECT 14.0320 56.9835 14.0580 58.0770 ;
        RECT 13.9240 56.9835 13.9500 58.0770 ;
        RECT 13.8160 56.9835 13.8420 58.0770 ;
        RECT 13.7080 56.9835 13.7340 58.0770 ;
        RECT 13.6000 56.9835 13.6260 58.0770 ;
        RECT 13.4920 56.9835 13.5180 58.0770 ;
        RECT 13.3840 56.9835 13.4100 58.0770 ;
        RECT 13.2760 56.9835 13.3020 58.0770 ;
        RECT 13.1680 56.9835 13.1940 58.0770 ;
        RECT 13.0600 56.9835 13.0860 58.0770 ;
        RECT 12.9520 56.9835 12.9780 58.0770 ;
        RECT 12.8440 56.9835 12.8700 58.0770 ;
        RECT 12.7360 56.9835 12.7620 58.0770 ;
        RECT 12.6280 56.9835 12.6540 58.0770 ;
        RECT 12.5200 56.9835 12.5460 58.0770 ;
        RECT 12.4120 56.9835 12.4380 58.0770 ;
        RECT 12.3040 56.9835 12.3300 58.0770 ;
        RECT 12.1960 56.9835 12.2220 58.0770 ;
        RECT 12.0880 56.9835 12.1140 58.0770 ;
        RECT 11.9800 56.9835 12.0060 58.0770 ;
        RECT 11.8720 56.9835 11.8980 58.0770 ;
        RECT 11.7640 56.9835 11.7900 58.0770 ;
        RECT 11.6560 56.9835 11.6820 58.0770 ;
        RECT 11.5480 56.9835 11.5740 58.0770 ;
        RECT 11.4400 56.9835 11.4660 58.0770 ;
        RECT 11.3320 56.9835 11.3580 58.0770 ;
        RECT 11.2240 56.9835 11.2500 58.0770 ;
        RECT 11.1160 56.9835 11.1420 58.0770 ;
        RECT 11.0080 56.9835 11.0340 58.0770 ;
        RECT 10.9000 56.9835 10.9260 58.0770 ;
        RECT 10.7920 56.9835 10.8180 58.0770 ;
        RECT 10.6840 56.9835 10.7100 58.0770 ;
        RECT 10.5760 56.9835 10.6020 58.0770 ;
        RECT 10.4680 56.9835 10.4940 58.0770 ;
        RECT 10.3600 56.9835 10.3860 58.0770 ;
        RECT 10.2520 56.9835 10.2780 58.0770 ;
        RECT 10.1440 56.9835 10.1700 58.0770 ;
        RECT 10.0360 56.9835 10.0620 58.0770 ;
        RECT 9.9280 56.9835 9.9540 58.0770 ;
        RECT 9.8200 56.9835 9.8460 58.0770 ;
        RECT 9.7120 56.9835 9.7380 58.0770 ;
        RECT 9.6040 56.9835 9.6300 58.0770 ;
        RECT 9.4960 56.9835 9.5220 58.0770 ;
        RECT 9.3880 56.9835 9.4140 58.0770 ;
        RECT 9.1750 56.9835 9.2520 58.0770 ;
        RECT 7.2820 56.9835 7.3590 58.0770 ;
        RECT 7.1200 56.9835 7.1460 58.0770 ;
        RECT 7.0120 56.9835 7.0380 58.0770 ;
        RECT 6.9040 56.9835 6.9300 58.0770 ;
        RECT 6.7960 56.9835 6.8220 58.0770 ;
        RECT 6.6880 56.9835 6.7140 58.0770 ;
        RECT 6.5800 56.9835 6.6060 58.0770 ;
        RECT 6.4720 56.9835 6.4980 58.0770 ;
        RECT 6.3640 56.9835 6.3900 58.0770 ;
        RECT 6.2560 56.9835 6.2820 58.0770 ;
        RECT 6.1480 56.9835 6.1740 58.0770 ;
        RECT 6.0400 56.9835 6.0660 58.0770 ;
        RECT 5.9320 56.9835 5.9580 58.0770 ;
        RECT 5.8240 56.9835 5.8500 58.0770 ;
        RECT 5.7160 56.9835 5.7420 58.0770 ;
        RECT 5.6080 56.9835 5.6340 58.0770 ;
        RECT 5.5000 56.9835 5.5260 58.0770 ;
        RECT 5.3920 56.9835 5.4180 58.0770 ;
        RECT 5.2840 56.9835 5.3100 58.0770 ;
        RECT 5.1760 56.9835 5.2020 58.0770 ;
        RECT 5.0680 56.9835 5.0940 58.0770 ;
        RECT 4.9600 56.9835 4.9860 58.0770 ;
        RECT 4.8520 56.9835 4.8780 58.0770 ;
        RECT 4.7440 56.9835 4.7700 58.0770 ;
        RECT 4.6360 56.9835 4.6620 58.0770 ;
        RECT 4.5280 56.9835 4.5540 58.0770 ;
        RECT 4.4200 56.9835 4.4460 58.0770 ;
        RECT 4.3120 56.9835 4.3380 58.0770 ;
        RECT 4.2040 56.9835 4.2300 58.0770 ;
        RECT 4.0960 56.9835 4.1220 58.0770 ;
        RECT 3.9880 56.9835 4.0140 58.0770 ;
        RECT 3.8800 56.9835 3.9060 58.0770 ;
        RECT 3.7720 56.9835 3.7980 58.0770 ;
        RECT 3.6640 56.9835 3.6900 58.0770 ;
        RECT 3.5560 56.9835 3.5820 58.0770 ;
        RECT 3.4480 56.9835 3.4740 58.0770 ;
        RECT 3.3400 56.9835 3.3660 58.0770 ;
        RECT 3.2320 56.9835 3.2580 58.0770 ;
        RECT 3.1240 56.9835 3.1500 58.0770 ;
        RECT 3.0160 56.9835 3.0420 58.0770 ;
        RECT 2.9080 56.9835 2.9340 58.0770 ;
        RECT 2.8000 56.9835 2.8260 58.0770 ;
        RECT 2.6920 56.9835 2.7180 58.0770 ;
        RECT 2.5840 56.9835 2.6100 58.0770 ;
        RECT 2.4760 56.9835 2.5020 58.0770 ;
        RECT 2.3680 56.9835 2.3940 58.0770 ;
        RECT 2.2600 56.9835 2.2860 58.0770 ;
        RECT 2.1520 56.9835 2.1780 58.0770 ;
        RECT 2.0440 56.9835 2.0700 58.0770 ;
        RECT 1.9360 56.9835 1.9620 58.0770 ;
        RECT 1.8280 56.9835 1.8540 58.0770 ;
        RECT 1.7200 56.9835 1.7460 58.0770 ;
        RECT 1.6120 56.9835 1.6380 58.0770 ;
        RECT 1.5040 56.9835 1.5300 58.0770 ;
        RECT 1.3960 56.9835 1.4220 58.0770 ;
        RECT 1.2880 56.9835 1.3140 58.0770 ;
        RECT 1.1800 56.9835 1.2060 58.0770 ;
        RECT 1.0720 56.9835 1.0980 58.0770 ;
        RECT 0.9640 56.9835 0.9900 58.0770 ;
        RECT 0.8560 56.9835 0.8820 58.0770 ;
        RECT 0.7480 56.9835 0.7740 58.0770 ;
        RECT 0.6400 56.9835 0.6660 58.0770 ;
        RECT 0.5320 56.9835 0.5580 58.0770 ;
        RECT 0.4240 56.9835 0.4500 58.0770 ;
        RECT 0.3160 56.9835 0.3420 58.0770 ;
        RECT 0.2080 56.9835 0.2340 58.0770 ;
        RECT 0.0050 56.9835 0.0900 58.0770 ;
        RECT 8.6410 58.0635 8.7690 59.1570 ;
        RECT 8.6270 58.7290 8.7690 59.0515 ;
        RECT 8.4790 58.4560 8.5410 59.1570 ;
        RECT 8.4650 58.7655 8.5410 58.9190 ;
        RECT 8.4790 58.0635 8.5050 59.1570 ;
        RECT 8.4790 58.1845 8.5190 58.4240 ;
        RECT 8.4790 58.0635 8.5410 58.1525 ;
        RECT 8.1820 58.5140 8.3880 59.1570 ;
        RECT 8.3620 58.0635 8.3880 59.1570 ;
        RECT 8.1820 58.7910 8.4020 59.0490 ;
        RECT 8.1820 58.0635 8.2800 59.1570 ;
        RECT 7.7650 58.0635 7.8480 59.1570 ;
        RECT 7.7650 58.1520 7.8620 59.0875 ;
        RECT 16.4440 58.0635 16.5290 59.1570 ;
        RECT 16.3000 58.0635 16.3260 59.1570 ;
        RECT 16.1920 58.0635 16.2180 59.1570 ;
        RECT 16.0840 58.0635 16.1100 59.1570 ;
        RECT 15.9760 58.0635 16.0020 59.1570 ;
        RECT 15.8680 58.0635 15.8940 59.1570 ;
        RECT 15.7600 58.0635 15.7860 59.1570 ;
        RECT 15.6520 58.0635 15.6780 59.1570 ;
        RECT 15.5440 58.0635 15.5700 59.1570 ;
        RECT 15.4360 58.0635 15.4620 59.1570 ;
        RECT 15.3280 58.0635 15.3540 59.1570 ;
        RECT 15.2200 58.0635 15.2460 59.1570 ;
        RECT 15.1120 58.0635 15.1380 59.1570 ;
        RECT 15.0040 58.0635 15.0300 59.1570 ;
        RECT 14.8960 58.0635 14.9220 59.1570 ;
        RECT 14.7880 58.0635 14.8140 59.1570 ;
        RECT 14.6800 58.0635 14.7060 59.1570 ;
        RECT 14.5720 58.0635 14.5980 59.1570 ;
        RECT 14.4640 58.0635 14.4900 59.1570 ;
        RECT 14.3560 58.0635 14.3820 59.1570 ;
        RECT 14.2480 58.0635 14.2740 59.1570 ;
        RECT 14.1400 58.0635 14.1660 59.1570 ;
        RECT 14.0320 58.0635 14.0580 59.1570 ;
        RECT 13.9240 58.0635 13.9500 59.1570 ;
        RECT 13.8160 58.0635 13.8420 59.1570 ;
        RECT 13.7080 58.0635 13.7340 59.1570 ;
        RECT 13.6000 58.0635 13.6260 59.1570 ;
        RECT 13.4920 58.0635 13.5180 59.1570 ;
        RECT 13.3840 58.0635 13.4100 59.1570 ;
        RECT 13.2760 58.0635 13.3020 59.1570 ;
        RECT 13.1680 58.0635 13.1940 59.1570 ;
        RECT 13.0600 58.0635 13.0860 59.1570 ;
        RECT 12.9520 58.0635 12.9780 59.1570 ;
        RECT 12.8440 58.0635 12.8700 59.1570 ;
        RECT 12.7360 58.0635 12.7620 59.1570 ;
        RECT 12.6280 58.0635 12.6540 59.1570 ;
        RECT 12.5200 58.0635 12.5460 59.1570 ;
        RECT 12.4120 58.0635 12.4380 59.1570 ;
        RECT 12.3040 58.0635 12.3300 59.1570 ;
        RECT 12.1960 58.0635 12.2220 59.1570 ;
        RECT 12.0880 58.0635 12.1140 59.1570 ;
        RECT 11.9800 58.0635 12.0060 59.1570 ;
        RECT 11.8720 58.0635 11.8980 59.1570 ;
        RECT 11.7640 58.0635 11.7900 59.1570 ;
        RECT 11.6560 58.0635 11.6820 59.1570 ;
        RECT 11.5480 58.0635 11.5740 59.1570 ;
        RECT 11.4400 58.0635 11.4660 59.1570 ;
        RECT 11.3320 58.0635 11.3580 59.1570 ;
        RECT 11.2240 58.0635 11.2500 59.1570 ;
        RECT 11.1160 58.0635 11.1420 59.1570 ;
        RECT 11.0080 58.0635 11.0340 59.1570 ;
        RECT 10.9000 58.0635 10.9260 59.1570 ;
        RECT 10.7920 58.0635 10.8180 59.1570 ;
        RECT 10.6840 58.0635 10.7100 59.1570 ;
        RECT 10.5760 58.0635 10.6020 59.1570 ;
        RECT 10.4680 58.0635 10.4940 59.1570 ;
        RECT 10.3600 58.0635 10.3860 59.1570 ;
        RECT 10.2520 58.0635 10.2780 59.1570 ;
        RECT 10.1440 58.0635 10.1700 59.1570 ;
        RECT 10.0360 58.0635 10.0620 59.1570 ;
        RECT 9.9280 58.0635 9.9540 59.1570 ;
        RECT 9.8200 58.0635 9.8460 59.1570 ;
        RECT 9.7120 58.0635 9.7380 59.1570 ;
        RECT 9.6040 58.0635 9.6300 59.1570 ;
        RECT 9.4960 58.0635 9.5220 59.1570 ;
        RECT 9.3880 58.0635 9.4140 59.1570 ;
        RECT 9.1750 58.0635 9.2520 59.1570 ;
        RECT 7.2820 58.0635 7.3590 59.1570 ;
        RECT 7.1200 58.0635 7.1460 59.1570 ;
        RECT 7.0120 58.0635 7.0380 59.1570 ;
        RECT 6.9040 58.0635 6.9300 59.1570 ;
        RECT 6.7960 58.0635 6.8220 59.1570 ;
        RECT 6.6880 58.0635 6.7140 59.1570 ;
        RECT 6.5800 58.0635 6.6060 59.1570 ;
        RECT 6.4720 58.0635 6.4980 59.1570 ;
        RECT 6.3640 58.0635 6.3900 59.1570 ;
        RECT 6.2560 58.0635 6.2820 59.1570 ;
        RECT 6.1480 58.0635 6.1740 59.1570 ;
        RECT 6.0400 58.0635 6.0660 59.1570 ;
        RECT 5.9320 58.0635 5.9580 59.1570 ;
        RECT 5.8240 58.0635 5.8500 59.1570 ;
        RECT 5.7160 58.0635 5.7420 59.1570 ;
        RECT 5.6080 58.0635 5.6340 59.1570 ;
        RECT 5.5000 58.0635 5.5260 59.1570 ;
        RECT 5.3920 58.0635 5.4180 59.1570 ;
        RECT 5.2840 58.0635 5.3100 59.1570 ;
        RECT 5.1760 58.0635 5.2020 59.1570 ;
        RECT 5.0680 58.0635 5.0940 59.1570 ;
        RECT 4.9600 58.0635 4.9860 59.1570 ;
        RECT 4.8520 58.0635 4.8780 59.1570 ;
        RECT 4.7440 58.0635 4.7700 59.1570 ;
        RECT 4.6360 58.0635 4.6620 59.1570 ;
        RECT 4.5280 58.0635 4.5540 59.1570 ;
        RECT 4.4200 58.0635 4.4460 59.1570 ;
        RECT 4.3120 58.0635 4.3380 59.1570 ;
        RECT 4.2040 58.0635 4.2300 59.1570 ;
        RECT 4.0960 58.0635 4.1220 59.1570 ;
        RECT 3.9880 58.0635 4.0140 59.1570 ;
        RECT 3.8800 58.0635 3.9060 59.1570 ;
        RECT 3.7720 58.0635 3.7980 59.1570 ;
        RECT 3.6640 58.0635 3.6900 59.1570 ;
        RECT 3.5560 58.0635 3.5820 59.1570 ;
        RECT 3.4480 58.0635 3.4740 59.1570 ;
        RECT 3.3400 58.0635 3.3660 59.1570 ;
        RECT 3.2320 58.0635 3.2580 59.1570 ;
        RECT 3.1240 58.0635 3.1500 59.1570 ;
        RECT 3.0160 58.0635 3.0420 59.1570 ;
        RECT 2.9080 58.0635 2.9340 59.1570 ;
        RECT 2.8000 58.0635 2.8260 59.1570 ;
        RECT 2.6920 58.0635 2.7180 59.1570 ;
        RECT 2.5840 58.0635 2.6100 59.1570 ;
        RECT 2.4760 58.0635 2.5020 59.1570 ;
        RECT 2.3680 58.0635 2.3940 59.1570 ;
        RECT 2.2600 58.0635 2.2860 59.1570 ;
        RECT 2.1520 58.0635 2.1780 59.1570 ;
        RECT 2.0440 58.0635 2.0700 59.1570 ;
        RECT 1.9360 58.0635 1.9620 59.1570 ;
        RECT 1.8280 58.0635 1.8540 59.1570 ;
        RECT 1.7200 58.0635 1.7460 59.1570 ;
        RECT 1.6120 58.0635 1.6380 59.1570 ;
        RECT 1.5040 58.0635 1.5300 59.1570 ;
        RECT 1.3960 58.0635 1.4220 59.1570 ;
        RECT 1.2880 58.0635 1.3140 59.1570 ;
        RECT 1.1800 58.0635 1.2060 59.1570 ;
        RECT 1.0720 58.0635 1.0980 59.1570 ;
        RECT 0.9640 58.0635 0.9900 59.1570 ;
        RECT 0.8560 58.0635 0.8820 59.1570 ;
        RECT 0.7480 58.0635 0.7740 59.1570 ;
        RECT 0.6400 58.0635 0.6660 59.1570 ;
        RECT 0.5320 58.0635 0.5580 59.1570 ;
        RECT 0.4240 58.0635 0.4500 59.1570 ;
        RECT 0.3160 58.0635 0.3420 59.1570 ;
        RECT 0.2080 58.0635 0.2340 59.1570 ;
        RECT 0.0050 58.0635 0.0900 59.1570 ;
        RECT 8.6410 59.1435 8.7690 60.2370 ;
        RECT 8.6270 59.8090 8.7690 60.1315 ;
        RECT 8.4790 59.5360 8.5410 60.2370 ;
        RECT 8.4650 59.8455 8.5410 59.9990 ;
        RECT 8.4790 59.1435 8.5050 60.2370 ;
        RECT 8.4790 59.2645 8.5190 59.5040 ;
        RECT 8.4790 59.1435 8.5410 59.2325 ;
        RECT 8.1820 59.5940 8.3880 60.2370 ;
        RECT 8.3620 59.1435 8.3880 60.2370 ;
        RECT 8.1820 59.8710 8.4020 60.1290 ;
        RECT 8.1820 59.1435 8.2800 60.2370 ;
        RECT 7.7650 59.1435 7.8480 60.2370 ;
        RECT 7.7650 59.2320 7.8620 60.1675 ;
        RECT 16.4440 59.1435 16.5290 60.2370 ;
        RECT 16.3000 59.1435 16.3260 60.2370 ;
        RECT 16.1920 59.1435 16.2180 60.2370 ;
        RECT 16.0840 59.1435 16.1100 60.2370 ;
        RECT 15.9760 59.1435 16.0020 60.2370 ;
        RECT 15.8680 59.1435 15.8940 60.2370 ;
        RECT 15.7600 59.1435 15.7860 60.2370 ;
        RECT 15.6520 59.1435 15.6780 60.2370 ;
        RECT 15.5440 59.1435 15.5700 60.2370 ;
        RECT 15.4360 59.1435 15.4620 60.2370 ;
        RECT 15.3280 59.1435 15.3540 60.2370 ;
        RECT 15.2200 59.1435 15.2460 60.2370 ;
        RECT 15.1120 59.1435 15.1380 60.2370 ;
        RECT 15.0040 59.1435 15.0300 60.2370 ;
        RECT 14.8960 59.1435 14.9220 60.2370 ;
        RECT 14.7880 59.1435 14.8140 60.2370 ;
        RECT 14.6800 59.1435 14.7060 60.2370 ;
        RECT 14.5720 59.1435 14.5980 60.2370 ;
        RECT 14.4640 59.1435 14.4900 60.2370 ;
        RECT 14.3560 59.1435 14.3820 60.2370 ;
        RECT 14.2480 59.1435 14.2740 60.2370 ;
        RECT 14.1400 59.1435 14.1660 60.2370 ;
        RECT 14.0320 59.1435 14.0580 60.2370 ;
        RECT 13.9240 59.1435 13.9500 60.2370 ;
        RECT 13.8160 59.1435 13.8420 60.2370 ;
        RECT 13.7080 59.1435 13.7340 60.2370 ;
        RECT 13.6000 59.1435 13.6260 60.2370 ;
        RECT 13.4920 59.1435 13.5180 60.2370 ;
        RECT 13.3840 59.1435 13.4100 60.2370 ;
        RECT 13.2760 59.1435 13.3020 60.2370 ;
        RECT 13.1680 59.1435 13.1940 60.2370 ;
        RECT 13.0600 59.1435 13.0860 60.2370 ;
        RECT 12.9520 59.1435 12.9780 60.2370 ;
        RECT 12.8440 59.1435 12.8700 60.2370 ;
        RECT 12.7360 59.1435 12.7620 60.2370 ;
        RECT 12.6280 59.1435 12.6540 60.2370 ;
        RECT 12.5200 59.1435 12.5460 60.2370 ;
        RECT 12.4120 59.1435 12.4380 60.2370 ;
        RECT 12.3040 59.1435 12.3300 60.2370 ;
        RECT 12.1960 59.1435 12.2220 60.2370 ;
        RECT 12.0880 59.1435 12.1140 60.2370 ;
        RECT 11.9800 59.1435 12.0060 60.2370 ;
        RECT 11.8720 59.1435 11.8980 60.2370 ;
        RECT 11.7640 59.1435 11.7900 60.2370 ;
        RECT 11.6560 59.1435 11.6820 60.2370 ;
        RECT 11.5480 59.1435 11.5740 60.2370 ;
        RECT 11.4400 59.1435 11.4660 60.2370 ;
        RECT 11.3320 59.1435 11.3580 60.2370 ;
        RECT 11.2240 59.1435 11.2500 60.2370 ;
        RECT 11.1160 59.1435 11.1420 60.2370 ;
        RECT 11.0080 59.1435 11.0340 60.2370 ;
        RECT 10.9000 59.1435 10.9260 60.2370 ;
        RECT 10.7920 59.1435 10.8180 60.2370 ;
        RECT 10.6840 59.1435 10.7100 60.2370 ;
        RECT 10.5760 59.1435 10.6020 60.2370 ;
        RECT 10.4680 59.1435 10.4940 60.2370 ;
        RECT 10.3600 59.1435 10.3860 60.2370 ;
        RECT 10.2520 59.1435 10.2780 60.2370 ;
        RECT 10.1440 59.1435 10.1700 60.2370 ;
        RECT 10.0360 59.1435 10.0620 60.2370 ;
        RECT 9.9280 59.1435 9.9540 60.2370 ;
        RECT 9.8200 59.1435 9.8460 60.2370 ;
        RECT 9.7120 59.1435 9.7380 60.2370 ;
        RECT 9.6040 59.1435 9.6300 60.2370 ;
        RECT 9.4960 59.1435 9.5220 60.2370 ;
        RECT 9.3880 59.1435 9.4140 60.2370 ;
        RECT 9.1750 59.1435 9.2520 60.2370 ;
        RECT 7.2820 59.1435 7.3590 60.2370 ;
        RECT 7.1200 59.1435 7.1460 60.2370 ;
        RECT 7.0120 59.1435 7.0380 60.2370 ;
        RECT 6.9040 59.1435 6.9300 60.2370 ;
        RECT 6.7960 59.1435 6.8220 60.2370 ;
        RECT 6.6880 59.1435 6.7140 60.2370 ;
        RECT 6.5800 59.1435 6.6060 60.2370 ;
        RECT 6.4720 59.1435 6.4980 60.2370 ;
        RECT 6.3640 59.1435 6.3900 60.2370 ;
        RECT 6.2560 59.1435 6.2820 60.2370 ;
        RECT 6.1480 59.1435 6.1740 60.2370 ;
        RECT 6.0400 59.1435 6.0660 60.2370 ;
        RECT 5.9320 59.1435 5.9580 60.2370 ;
        RECT 5.8240 59.1435 5.8500 60.2370 ;
        RECT 5.7160 59.1435 5.7420 60.2370 ;
        RECT 5.6080 59.1435 5.6340 60.2370 ;
        RECT 5.5000 59.1435 5.5260 60.2370 ;
        RECT 5.3920 59.1435 5.4180 60.2370 ;
        RECT 5.2840 59.1435 5.3100 60.2370 ;
        RECT 5.1760 59.1435 5.2020 60.2370 ;
        RECT 5.0680 59.1435 5.0940 60.2370 ;
        RECT 4.9600 59.1435 4.9860 60.2370 ;
        RECT 4.8520 59.1435 4.8780 60.2370 ;
        RECT 4.7440 59.1435 4.7700 60.2370 ;
        RECT 4.6360 59.1435 4.6620 60.2370 ;
        RECT 4.5280 59.1435 4.5540 60.2370 ;
        RECT 4.4200 59.1435 4.4460 60.2370 ;
        RECT 4.3120 59.1435 4.3380 60.2370 ;
        RECT 4.2040 59.1435 4.2300 60.2370 ;
        RECT 4.0960 59.1435 4.1220 60.2370 ;
        RECT 3.9880 59.1435 4.0140 60.2370 ;
        RECT 3.8800 59.1435 3.9060 60.2370 ;
        RECT 3.7720 59.1435 3.7980 60.2370 ;
        RECT 3.6640 59.1435 3.6900 60.2370 ;
        RECT 3.5560 59.1435 3.5820 60.2370 ;
        RECT 3.4480 59.1435 3.4740 60.2370 ;
        RECT 3.3400 59.1435 3.3660 60.2370 ;
        RECT 3.2320 59.1435 3.2580 60.2370 ;
        RECT 3.1240 59.1435 3.1500 60.2370 ;
        RECT 3.0160 59.1435 3.0420 60.2370 ;
        RECT 2.9080 59.1435 2.9340 60.2370 ;
        RECT 2.8000 59.1435 2.8260 60.2370 ;
        RECT 2.6920 59.1435 2.7180 60.2370 ;
        RECT 2.5840 59.1435 2.6100 60.2370 ;
        RECT 2.4760 59.1435 2.5020 60.2370 ;
        RECT 2.3680 59.1435 2.3940 60.2370 ;
        RECT 2.2600 59.1435 2.2860 60.2370 ;
        RECT 2.1520 59.1435 2.1780 60.2370 ;
        RECT 2.0440 59.1435 2.0700 60.2370 ;
        RECT 1.9360 59.1435 1.9620 60.2370 ;
        RECT 1.8280 59.1435 1.8540 60.2370 ;
        RECT 1.7200 59.1435 1.7460 60.2370 ;
        RECT 1.6120 59.1435 1.6380 60.2370 ;
        RECT 1.5040 59.1435 1.5300 60.2370 ;
        RECT 1.3960 59.1435 1.4220 60.2370 ;
        RECT 1.2880 59.1435 1.3140 60.2370 ;
        RECT 1.1800 59.1435 1.2060 60.2370 ;
        RECT 1.0720 59.1435 1.0980 60.2370 ;
        RECT 0.9640 59.1435 0.9900 60.2370 ;
        RECT 0.8560 59.1435 0.8820 60.2370 ;
        RECT 0.7480 59.1435 0.7740 60.2370 ;
        RECT 0.6400 59.1435 0.6660 60.2370 ;
        RECT 0.5320 59.1435 0.5580 60.2370 ;
        RECT 0.4240 59.1435 0.4500 60.2370 ;
        RECT 0.3160 59.1435 0.3420 60.2370 ;
        RECT 0.2080 59.1435 0.2340 60.2370 ;
        RECT 0.0050 59.1435 0.0900 60.2370 ;
        RECT 8.6410 60.2235 8.7690 61.3170 ;
        RECT 8.6270 60.8890 8.7690 61.2115 ;
        RECT 8.4790 60.6160 8.5410 61.3170 ;
        RECT 8.4650 60.9255 8.5410 61.0790 ;
        RECT 8.4790 60.2235 8.5050 61.3170 ;
        RECT 8.4790 60.3445 8.5190 60.5840 ;
        RECT 8.4790 60.2235 8.5410 60.3125 ;
        RECT 8.1820 60.6740 8.3880 61.3170 ;
        RECT 8.3620 60.2235 8.3880 61.3170 ;
        RECT 8.1820 60.9510 8.4020 61.2090 ;
        RECT 8.1820 60.2235 8.2800 61.3170 ;
        RECT 7.7650 60.2235 7.8480 61.3170 ;
        RECT 7.7650 60.3120 7.8620 61.2475 ;
        RECT 16.4440 60.2235 16.5290 61.3170 ;
        RECT 16.3000 60.2235 16.3260 61.3170 ;
        RECT 16.1920 60.2235 16.2180 61.3170 ;
        RECT 16.0840 60.2235 16.1100 61.3170 ;
        RECT 15.9760 60.2235 16.0020 61.3170 ;
        RECT 15.8680 60.2235 15.8940 61.3170 ;
        RECT 15.7600 60.2235 15.7860 61.3170 ;
        RECT 15.6520 60.2235 15.6780 61.3170 ;
        RECT 15.5440 60.2235 15.5700 61.3170 ;
        RECT 15.4360 60.2235 15.4620 61.3170 ;
        RECT 15.3280 60.2235 15.3540 61.3170 ;
        RECT 15.2200 60.2235 15.2460 61.3170 ;
        RECT 15.1120 60.2235 15.1380 61.3170 ;
        RECT 15.0040 60.2235 15.0300 61.3170 ;
        RECT 14.8960 60.2235 14.9220 61.3170 ;
        RECT 14.7880 60.2235 14.8140 61.3170 ;
        RECT 14.6800 60.2235 14.7060 61.3170 ;
        RECT 14.5720 60.2235 14.5980 61.3170 ;
        RECT 14.4640 60.2235 14.4900 61.3170 ;
        RECT 14.3560 60.2235 14.3820 61.3170 ;
        RECT 14.2480 60.2235 14.2740 61.3170 ;
        RECT 14.1400 60.2235 14.1660 61.3170 ;
        RECT 14.0320 60.2235 14.0580 61.3170 ;
        RECT 13.9240 60.2235 13.9500 61.3170 ;
        RECT 13.8160 60.2235 13.8420 61.3170 ;
        RECT 13.7080 60.2235 13.7340 61.3170 ;
        RECT 13.6000 60.2235 13.6260 61.3170 ;
        RECT 13.4920 60.2235 13.5180 61.3170 ;
        RECT 13.3840 60.2235 13.4100 61.3170 ;
        RECT 13.2760 60.2235 13.3020 61.3170 ;
        RECT 13.1680 60.2235 13.1940 61.3170 ;
        RECT 13.0600 60.2235 13.0860 61.3170 ;
        RECT 12.9520 60.2235 12.9780 61.3170 ;
        RECT 12.8440 60.2235 12.8700 61.3170 ;
        RECT 12.7360 60.2235 12.7620 61.3170 ;
        RECT 12.6280 60.2235 12.6540 61.3170 ;
        RECT 12.5200 60.2235 12.5460 61.3170 ;
        RECT 12.4120 60.2235 12.4380 61.3170 ;
        RECT 12.3040 60.2235 12.3300 61.3170 ;
        RECT 12.1960 60.2235 12.2220 61.3170 ;
        RECT 12.0880 60.2235 12.1140 61.3170 ;
        RECT 11.9800 60.2235 12.0060 61.3170 ;
        RECT 11.8720 60.2235 11.8980 61.3170 ;
        RECT 11.7640 60.2235 11.7900 61.3170 ;
        RECT 11.6560 60.2235 11.6820 61.3170 ;
        RECT 11.5480 60.2235 11.5740 61.3170 ;
        RECT 11.4400 60.2235 11.4660 61.3170 ;
        RECT 11.3320 60.2235 11.3580 61.3170 ;
        RECT 11.2240 60.2235 11.2500 61.3170 ;
        RECT 11.1160 60.2235 11.1420 61.3170 ;
        RECT 11.0080 60.2235 11.0340 61.3170 ;
        RECT 10.9000 60.2235 10.9260 61.3170 ;
        RECT 10.7920 60.2235 10.8180 61.3170 ;
        RECT 10.6840 60.2235 10.7100 61.3170 ;
        RECT 10.5760 60.2235 10.6020 61.3170 ;
        RECT 10.4680 60.2235 10.4940 61.3170 ;
        RECT 10.3600 60.2235 10.3860 61.3170 ;
        RECT 10.2520 60.2235 10.2780 61.3170 ;
        RECT 10.1440 60.2235 10.1700 61.3170 ;
        RECT 10.0360 60.2235 10.0620 61.3170 ;
        RECT 9.9280 60.2235 9.9540 61.3170 ;
        RECT 9.8200 60.2235 9.8460 61.3170 ;
        RECT 9.7120 60.2235 9.7380 61.3170 ;
        RECT 9.6040 60.2235 9.6300 61.3170 ;
        RECT 9.4960 60.2235 9.5220 61.3170 ;
        RECT 9.3880 60.2235 9.4140 61.3170 ;
        RECT 9.1750 60.2235 9.2520 61.3170 ;
        RECT 7.2820 60.2235 7.3590 61.3170 ;
        RECT 7.1200 60.2235 7.1460 61.3170 ;
        RECT 7.0120 60.2235 7.0380 61.3170 ;
        RECT 6.9040 60.2235 6.9300 61.3170 ;
        RECT 6.7960 60.2235 6.8220 61.3170 ;
        RECT 6.6880 60.2235 6.7140 61.3170 ;
        RECT 6.5800 60.2235 6.6060 61.3170 ;
        RECT 6.4720 60.2235 6.4980 61.3170 ;
        RECT 6.3640 60.2235 6.3900 61.3170 ;
        RECT 6.2560 60.2235 6.2820 61.3170 ;
        RECT 6.1480 60.2235 6.1740 61.3170 ;
        RECT 6.0400 60.2235 6.0660 61.3170 ;
        RECT 5.9320 60.2235 5.9580 61.3170 ;
        RECT 5.8240 60.2235 5.8500 61.3170 ;
        RECT 5.7160 60.2235 5.7420 61.3170 ;
        RECT 5.6080 60.2235 5.6340 61.3170 ;
        RECT 5.5000 60.2235 5.5260 61.3170 ;
        RECT 5.3920 60.2235 5.4180 61.3170 ;
        RECT 5.2840 60.2235 5.3100 61.3170 ;
        RECT 5.1760 60.2235 5.2020 61.3170 ;
        RECT 5.0680 60.2235 5.0940 61.3170 ;
        RECT 4.9600 60.2235 4.9860 61.3170 ;
        RECT 4.8520 60.2235 4.8780 61.3170 ;
        RECT 4.7440 60.2235 4.7700 61.3170 ;
        RECT 4.6360 60.2235 4.6620 61.3170 ;
        RECT 4.5280 60.2235 4.5540 61.3170 ;
        RECT 4.4200 60.2235 4.4460 61.3170 ;
        RECT 4.3120 60.2235 4.3380 61.3170 ;
        RECT 4.2040 60.2235 4.2300 61.3170 ;
        RECT 4.0960 60.2235 4.1220 61.3170 ;
        RECT 3.9880 60.2235 4.0140 61.3170 ;
        RECT 3.8800 60.2235 3.9060 61.3170 ;
        RECT 3.7720 60.2235 3.7980 61.3170 ;
        RECT 3.6640 60.2235 3.6900 61.3170 ;
        RECT 3.5560 60.2235 3.5820 61.3170 ;
        RECT 3.4480 60.2235 3.4740 61.3170 ;
        RECT 3.3400 60.2235 3.3660 61.3170 ;
        RECT 3.2320 60.2235 3.2580 61.3170 ;
        RECT 3.1240 60.2235 3.1500 61.3170 ;
        RECT 3.0160 60.2235 3.0420 61.3170 ;
        RECT 2.9080 60.2235 2.9340 61.3170 ;
        RECT 2.8000 60.2235 2.8260 61.3170 ;
        RECT 2.6920 60.2235 2.7180 61.3170 ;
        RECT 2.5840 60.2235 2.6100 61.3170 ;
        RECT 2.4760 60.2235 2.5020 61.3170 ;
        RECT 2.3680 60.2235 2.3940 61.3170 ;
        RECT 2.2600 60.2235 2.2860 61.3170 ;
        RECT 2.1520 60.2235 2.1780 61.3170 ;
        RECT 2.0440 60.2235 2.0700 61.3170 ;
        RECT 1.9360 60.2235 1.9620 61.3170 ;
        RECT 1.8280 60.2235 1.8540 61.3170 ;
        RECT 1.7200 60.2235 1.7460 61.3170 ;
        RECT 1.6120 60.2235 1.6380 61.3170 ;
        RECT 1.5040 60.2235 1.5300 61.3170 ;
        RECT 1.3960 60.2235 1.4220 61.3170 ;
        RECT 1.2880 60.2235 1.3140 61.3170 ;
        RECT 1.1800 60.2235 1.2060 61.3170 ;
        RECT 1.0720 60.2235 1.0980 61.3170 ;
        RECT 0.9640 60.2235 0.9900 61.3170 ;
        RECT 0.8560 60.2235 0.8820 61.3170 ;
        RECT 0.7480 60.2235 0.7740 61.3170 ;
        RECT 0.6400 60.2235 0.6660 61.3170 ;
        RECT 0.5320 60.2235 0.5580 61.3170 ;
        RECT 0.4240 60.2235 0.4500 61.3170 ;
        RECT 0.3160 60.2235 0.3420 61.3170 ;
        RECT 0.2080 60.2235 0.2340 61.3170 ;
        RECT 0.0050 60.2235 0.0900 61.3170 ;
        RECT 8.6410 61.3035 8.7690 62.3970 ;
        RECT 8.6270 61.9690 8.7690 62.2915 ;
        RECT 8.4790 61.6960 8.5410 62.3970 ;
        RECT 8.4650 62.0055 8.5410 62.1590 ;
        RECT 8.4790 61.3035 8.5050 62.3970 ;
        RECT 8.4790 61.4245 8.5190 61.6640 ;
        RECT 8.4790 61.3035 8.5410 61.3925 ;
        RECT 8.1820 61.7540 8.3880 62.3970 ;
        RECT 8.3620 61.3035 8.3880 62.3970 ;
        RECT 8.1820 62.0310 8.4020 62.2890 ;
        RECT 8.1820 61.3035 8.2800 62.3970 ;
        RECT 7.7650 61.3035 7.8480 62.3970 ;
        RECT 7.7650 61.3920 7.8620 62.3275 ;
        RECT 16.4440 61.3035 16.5290 62.3970 ;
        RECT 16.3000 61.3035 16.3260 62.3970 ;
        RECT 16.1920 61.3035 16.2180 62.3970 ;
        RECT 16.0840 61.3035 16.1100 62.3970 ;
        RECT 15.9760 61.3035 16.0020 62.3970 ;
        RECT 15.8680 61.3035 15.8940 62.3970 ;
        RECT 15.7600 61.3035 15.7860 62.3970 ;
        RECT 15.6520 61.3035 15.6780 62.3970 ;
        RECT 15.5440 61.3035 15.5700 62.3970 ;
        RECT 15.4360 61.3035 15.4620 62.3970 ;
        RECT 15.3280 61.3035 15.3540 62.3970 ;
        RECT 15.2200 61.3035 15.2460 62.3970 ;
        RECT 15.1120 61.3035 15.1380 62.3970 ;
        RECT 15.0040 61.3035 15.0300 62.3970 ;
        RECT 14.8960 61.3035 14.9220 62.3970 ;
        RECT 14.7880 61.3035 14.8140 62.3970 ;
        RECT 14.6800 61.3035 14.7060 62.3970 ;
        RECT 14.5720 61.3035 14.5980 62.3970 ;
        RECT 14.4640 61.3035 14.4900 62.3970 ;
        RECT 14.3560 61.3035 14.3820 62.3970 ;
        RECT 14.2480 61.3035 14.2740 62.3970 ;
        RECT 14.1400 61.3035 14.1660 62.3970 ;
        RECT 14.0320 61.3035 14.0580 62.3970 ;
        RECT 13.9240 61.3035 13.9500 62.3970 ;
        RECT 13.8160 61.3035 13.8420 62.3970 ;
        RECT 13.7080 61.3035 13.7340 62.3970 ;
        RECT 13.6000 61.3035 13.6260 62.3970 ;
        RECT 13.4920 61.3035 13.5180 62.3970 ;
        RECT 13.3840 61.3035 13.4100 62.3970 ;
        RECT 13.2760 61.3035 13.3020 62.3970 ;
        RECT 13.1680 61.3035 13.1940 62.3970 ;
        RECT 13.0600 61.3035 13.0860 62.3970 ;
        RECT 12.9520 61.3035 12.9780 62.3970 ;
        RECT 12.8440 61.3035 12.8700 62.3970 ;
        RECT 12.7360 61.3035 12.7620 62.3970 ;
        RECT 12.6280 61.3035 12.6540 62.3970 ;
        RECT 12.5200 61.3035 12.5460 62.3970 ;
        RECT 12.4120 61.3035 12.4380 62.3970 ;
        RECT 12.3040 61.3035 12.3300 62.3970 ;
        RECT 12.1960 61.3035 12.2220 62.3970 ;
        RECT 12.0880 61.3035 12.1140 62.3970 ;
        RECT 11.9800 61.3035 12.0060 62.3970 ;
        RECT 11.8720 61.3035 11.8980 62.3970 ;
        RECT 11.7640 61.3035 11.7900 62.3970 ;
        RECT 11.6560 61.3035 11.6820 62.3970 ;
        RECT 11.5480 61.3035 11.5740 62.3970 ;
        RECT 11.4400 61.3035 11.4660 62.3970 ;
        RECT 11.3320 61.3035 11.3580 62.3970 ;
        RECT 11.2240 61.3035 11.2500 62.3970 ;
        RECT 11.1160 61.3035 11.1420 62.3970 ;
        RECT 11.0080 61.3035 11.0340 62.3970 ;
        RECT 10.9000 61.3035 10.9260 62.3970 ;
        RECT 10.7920 61.3035 10.8180 62.3970 ;
        RECT 10.6840 61.3035 10.7100 62.3970 ;
        RECT 10.5760 61.3035 10.6020 62.3970 ;
        RECT 10.4680 61.3035 10.4940 62.3970 ;
        RECT 10.3600 61.3035 10.3860 62.3970 ;
        RECT 10.2520 61.3035 10.2780 62.3970 ;
        RECT 10.1440 61.3035 10.1700 62.3970 ;
        RECT 10.0360 61.3035 10.0620 62.3970 ;
        RECT 9.9280 61.3035 9.9540 62.3970 ;
        RECT 9.8200 61.3035 9.8460 62.3970 ;
        RECT 9.7120 61.3035 9.7380 62.3970 ;
        RECT 9.6040 61.3035 9.6300 62.3970 ;
        RECT 9.4960 61.3035 9.5220 62.3970 ;
        RECT 9.3880 61.3035 9.4140 62.3970 ;
        RECT 9.1750 61.3035 9.2520 62.3970 ;
        RECT 7.2820 61.3035 7.3590 62.3970 ;
        RECT 7.1200 61.3035 7.1460 62.3970 ;
        RECT 7.0120 61.3035 7.0380 62.3970 ;
        RECT 6.9040 61.3035 6.9300 62.3970 ;
        RECT 6.7960 61.3035 6.8220 62.3970 ;
        RECT 6.6880 61.3035 6.7140 62.3970 ;
        RECT 6.5800 61.3035 6.6060 62.3970 ;
        RECT 6.4720 61.3035 6.4980 62.3970 ;
        RECT 6.3640 61.3035 6.3900 62.3970 ;
        RECT 6.2560 61.3035 6.2820 62.3970 ;
        RECT 6.1480 61.3035 6.1740 62.3970 ;
        RECT 6.0400 61.3035 6.0660 62.3970 ;
        RECT 5.9320 61.3035 5.9580 62.3970 ;
        RECT 5.8240 61.3035 5.8500 62.3970 ;
        RECT 5.7160 61.3035 5.7420 62.3970 ;
        RECT 5.6080 61.3035 5.6340 62.3970 ;
        RECT 5.5000 61.3035 5.5260 62.3970 ;
        RECT 5.3920 61.3035 5.4180 62.3970 ;
        RECT 5.2840 61.3035 5.3100 62.3970 ;
        RECT 5.1760 61.3035 5.2020 62.3970 ;
        RECT 5.0680 61.3035 5.0940 62.3970 ;
        RECT 4.9600 61.3035 4.9860 62.3970 ;
        RECT 4.8520 61.3035 4.8780 62.3970 ;
        RECT 4.7440 61.3035 4.7700 62.3970 ;
        RECT 4.6360 61.3035 4.6620 62.3970 ;
        RECT 4.5280 61.3035 4.5540 62.3970 ;
        RECT 4.4200 61.3035 4.4460 62.3970 ;
        RECT 4.3120 61.3035 4.3380 62.3970 ;
        RECT 4.2040 61.3035 4.2300 62.3970 ;
        RECT 4.0960 61.3035 4.1220 62.3970 ;
        RECT 3.9880 61.3035 4.0140 62.3970 ;
        RECT 3.8800 61.3035 3.9060 62.3970 ;
        RECT 3.7720 61.3035 3.7980 62.3970 ;
        RECT 3.6640 61.3035 3.6900 62.3970 ;
        RECT 3.5560 61.3035 3.5820 62.3970 ;
        RECT 3.4480 61.3035 3.4740 62.3970 ;
        RECT 3.3400 61.3035 3.3660 62.3970 ;
        RECT 3.2320 61.3035 3.2580 62.3970 ;
        RECT 3.1240 61.3035 3.1500 62.3970 ;
        RECT 3.0160 61.3035 3.0420 62.3970 ;
        RECT 2.9080 61.3035 2.9340 62.3970 ;
        RECT 2.8000 61.3035 2.8260 62.3970 ;
        RECT 2.6920 61.3035 2.7180 62.3970 ;
        RECT 2.5840 61.3035 2.6100 62.3970 ;
        RECT 2.4760 61.3035 2.5020 62.3970 ;
        RECT 2.3680 61.3035 2.3940 62.3970 ;
        RECT 2.2600 61.3035 2.2860 62.3970 ;
        RECT 2.1520 61.3035 2.1780 62.3970 ;
        RECT 2.0440 61.3035 2.0700 62.3970 ;
        RECT 1.9360 61.3035 1.9620 62.3970 ;
        RECT 1.8280 61.3035 1.8540 62.3970 ;
        RECT 1.7200 61.3035 1.7460 62.3970 ;
        RECT 1.6120 61.3035 1.6380 62.3970 ;
        RECT 1.5040 61.3035 1.5300 62.3970 ;
        RECT 1.3960 61.3035 1.4220 62.3970 ;
        RECT 1.2880 61.3035 1.3140 62.3970 ;
        RECT 1.1800 61.3035 1.2060 62.3970 ;
        RECT 1.0720 61.3035 1.0980 62.3970 ;
        RECT 0.9640 61.3035 0.9900 62.3970 ;
        RECT 0.8560 61.3035 0.8820 62.3970 ;
        RECT 0.7480 61.3035 0.7740 62.3970 ;
        RECT 0.6400 61.3035 0.6660 62.3970 ;
        RECT 0.5320 61.3035 0.5580 62.3970 ;
        RECT 0.4240 61.3035 0.4500 62.3970 ;
        RECT 0.3160 61.3035 0.3420 62.3970 ;
        RECT 0.2080 61.3035 0.2340 62.3970 ;
        RECT 0.0050 61.3035 0.0900 62.3970 ;
        RECT 8.6410 62.3835 8.7690 63.4770 ;
        RECT 8.6270 63.0490 8.7690 63.3715 ;
        RECT 8.4790 62.7760 8.5410 63.4770 ;
        RECT 8.4650 63.0855 8.5410 63.2390 ;
        RECT 8.4790 62.3835 8.5050 63.4770 ;
        RECT 8.4790 62.5045 8.5190 62.7440 ;
        RECT 8.4790 62.3835 8.5410 62.4725 ;
        RECT 8.1820 62.8340 8.3880 63.4770 ;
        RECT 8.3620 62.3835 8.3880 63.4770 ;
        RECT 8.1820 63.1110 8.4020 63.3690 ;
        RECT 8.1820 62.3835 8.2800 63.4770 ;
        RECT 7.7650 62.3835 7.8480 63.4770 ;
        RECT 7.7650 62.4720 7.8620 63.4075 ;
        RECT 16.4440 62.3835 16.5290 63.4770 ;
        RECT 16.3000 62.3835 16.3260 63.4770 ;
        RECT 16.1920 62.3835 16.2180 63.4770 ;
        RECT 16.0840 62.3835 16.1100 63.4770 ;
        RECT 15.9760 62.3835 16.0020 63.4770 ;
        RECT 15.8680 62.3835 15.8940 63.4770 ;
        RECT 15.7600 62.3835 15.7860 63.4770 ;
        RECT 15.6520 62.3835 15.6780 63.4770 ;
        RECT 15.5440 62.3835 15.5700 63.4770 ;
        RECT 15.4360 62.3835 15.4620 63.4770 ;
        RECT 15.3280 62.3835 15.3540 63.4770 ;
        RECT 15.2200 62.3835 15.2460 63.4770 ;
        RECT 15.1120 62.3835 15.1380 63.4770 ;
        RECT 15.0040 62.3835 15.0300 63.4770 ;
        RECT 14.8960 62.3835 14.9220 63.4770 ;
        RECT 14.7880 62.3835 14.8140 63.4770 ;
        RECT 14.6800 62.3835 14.7060 63.4770 ;
        RECT 14.5720 62.3835 14.5980 63.4770 ;
        RECT 14.4640 62.3835 14.4900 63.4770 ;
        RECT 14.3560 62.3835 14.3820 63.4770 ;
        RECT 14.2480 62.3835 14.2740 63.4770 ;
        RECT 14.1400 62.3835 14.1660 63.4770 ;
        RECT 14.0320 62.3835 14.0580 63.4770 ;
        RECT 13.9240 62.3835 13.9500 63.4770 ;
        RECT 13.8160 62.3835 13.8420 63.4770 ;
        RECT 13.7080 62.3835 13.7340 63.4770 ;
        RECT 13.6000 62.3835 13.6260 63.4770 ;
        RECT 13.4920 62.3835 13.5180 63.4770 ;
        RECT 13.3840 62.3835 13.4100 63.4770 ;
        RECT 13.2760 62.3835 13.3020 63.4770 ;
        RECT 13.1680 62.3835 13.1940 63.4770 ;
        RECT 13.0600 62.3835 13.0860 63.4770 ;
        RECT 12.9520 62.3835 12.9780 63.4770 ;
        RECT 12.8440 62.3835 12.8700 63.4770 ;
        RECT 12.7360 62.3835 12.7620 63.4770 ;
        RECT 12.6280 62.3835 12.6540 63.4770 ;
        RECT 12.5200 62.3835 12.5460 63.4770 ;
        RECT 12.4120 62.3835 12.4380 63.4770 ;
        RECT 12.3040 62.3835 12.3300 63.4770 ;
        RECT 12.1960 62.3835 12.2220 63.4770 ;
        RECT 12.0880 62.3835 12.1140 63.4770 ;
        RECT 11.9800 62.3835 12.0060 63.4770 ;
        RECT 11.8720 62.3835 11.8980 63.4770 ;
        RECT 11.7640 62.3835 11.7900 63.4770 ;
        RECT 11.6560 62.3835 11.6820 63.4770 ;
        RECT 11.5480 62.3835 11.5740 63.4770 ;
        RECT 11.4400 62.3835 11.4660 63.4770 ;
        RECT 11.3320 62.3835 11.3580 63.4770 ;
        RECT 11.2240 62.3835 11.2500 63.4770 ;
        RECT 11.1160 62.3835 11.1420 63.4770 ;
        RECT 11.0080 62.3835 11.0340 63.4770 ;
        RECT 10.9000 62.3835 10.9260 63.4770 ;
        RECT 10.7920 62.3835 10.8180 63.4770 ;
        RECT 10.6840 62.3835 10.7100 63.4770 ;
        RECT 10.5760 62.3835 10.6020 63.4770 ;
        RECT 10.4680 62.3835 10.4940 63.4770 ;
        RECT 10.3600 62.3835 10.3860 63.4770 ;
        RECT 10.2520 62.3835 10.2780 63.4770 ;
        RECT 10.1440 62.3835 10.1700 63.4770 ;
        RECT 10.0360 62.3835 10.0620 63.4770 ;
        RECT 9.9280 62.3835 9.9540 63.4770 ;
        RECT 9.8200 62.3835 9.8460 63.4770 ;
        RECT 9.7120 62.3835 9.7380 63.4770 ;
        RECT 9.6040 62.3835 9.6300 63.4770 ;
        RECT 9.4960 62.3835 9.5220 63.4770 ;
        RECT 9.3880 62.3835 9.4140 63.4770 ;
        RECT 9.1750 62.3835 9.2520 63.4770 ;
        RECT 7.2820 62.3835 7.3590 63.4770 ;
        RECT 7.1200 62.3835 7.1460 63.4770 ;
        RECT 7.0120 62.3835 7.0380 63.4770 ;
        RECT 6.9040 62.3835 6.9300 63.4770 ;
        RECT 6.7960 62.3835 6.8220 63.4770 ;
        RECT 6.6880 62.3835 6.7140 63.4770 ;
        RECT 6.5800 62.3835 6.6060 63.4770 ;
        RECT 6.4720 62.3835 6.4980 63.4770 ;
        RECT 6.3640 62.3835 6.3900 63.4770 ;
        RECT 6.2560 62.3835 6.2820 63.4770 ;
        RECT 6.1480 62.3835 6.1740 63.4770 ;
        RECT 6.0400 62.3835 6.0660 63.4770 ;
        RECT 5.9320 62.3835 5.9580 63.4770 ;
        RECT 5.8240 62.3835 5.8500 63.4770 ;
        RECT 5.7160 62.3835 5.7420 63.4770 ;
        RECT 5.6080 62.3835 5.6340 63.4770 ;
        RECT 5.5000 62.3835 5.5260 63.4770 ;
        RECT 5.3920 62.3835 5.4180 63.4770 ;
        RECT 5.2840 62.3835 5.3100 63.4770 ;
        RECT 5.1760 62.3835 5.2020 63.4770 ;
        RECT 5.0680 62.3835 5.0940 63.4770 ;
        RECT 4.9600 62.3835 4.9860 63.4770 ;
        RECT 4.8520 62.3835 4.8780 63.4770 ;
        RECT 4.7440 62.3835 4.7700 63.4770 ;
        RECT 4.6360 62.3835 4.6620 63.4770 ;
        RECT 4.5280 62.3835 4.5540 63.4770 ;
        RECT 4.4200 62.3835 4.4460 63.4770 ;
        RECT 4.3120 62.3835 4.3380 63.4770 ;
        RECT 4.2040 62.3835 4.2300 63.4770 ;
        RECT 4.0960 62.3835 4.1220 63.4770 ;
        RECT 3.9880 62.3835 4.0140 63.4770 ;
        RECT 3.8800 62.3835 3.9060 63.4770 ;
        RECT 3.7720 62.3835 3.7980 63.4770 ;
        RECT 3.6640 62.3835 3.6900 63.4770 ;
        RECT 3.5560 62.3835 3.5820 63.4770 ;
        RECT 3.4480 62.3835 3.4740 63.4770 ;
        RECT 3.3400 62.3835 3.3660 63.4770 ;
        RECT 3.2320 62.3835 3.2580 63.4770 ;
        RECT 3.1240 62.3835 3.1500 63.4770 ;
        RECT 3.0160 62.3835 3.0420 63.4770 ;
        RECT 2.9080 62.3835 2.9340 63.4770 ;
        RECT 2.8000 62.3835 2.8260 63.4770 ;
        RECT 2.6920 62.3835 2.7180 63.4770 ;
        RECT 2.5840 62.3835 2.6100 63.4770 ;
        RECT 2.4760 62.3835 2.5020 63.4770 ;
        RECT 2.3680 62.3835 2.3940 63.4770 ;
        RECT 2.2600 62.3835 2.2860 63.4770 ;
        RECT 2.1520 62.3835 2.1780 63.4770 ;
        RECT 2.0440 62.3835 2.0700 63.4770 ;
        RECT 1.9360 62.3835 1.9620 63.4770 ;
        RECT 1.8280 62.3835 1.8540 63.4770 ;
        RECT 1.7200 62.3835 1.7460 63.4770 ;
        RECT 1.6120 62.3835 1.6380 63.4770 ;
        RECT 1.5040 62.3835 1.5300 63.4770 ;
        RECT 1.3960 62.3835 1.4220 63.4770 ;
        RECT 1.2880 62.3835 1.3140 63.4770 ;
        RECT 1.1800 62.3835 1.2060 63.4770 ;
        RECT 1.0720 62.3835 1.0980 63.4770 ;
        RECT 0.9640 62.3835 0.9900 63.4770 ;
        RECT 0.8560 62.3835 0.8820 63.4770 ;
        RECT 0.7480 62.3835 0.7740 63.4770 ;
        RECT 0.6400 62.3835 0.6660 63.4770 ;
        RECT 0.5320 62.3835 0.5580 63.4770 ;
        RECT 0.4240 62.3835 0.4500 63.4770 ;
        RECT 0.3160 62.3835 0.3420 63.4770 ;
        RECT 0.2080 62.3835 0.2340 63.4770 ;
        RECT 0.0050 62.3835 0.0900 63.4770 ;
        RECT 8.6410 63.4635 8.7690 64.5570 ;
        RECT 8.6270 64.1290 8.7690 64.4515 ;
        RECT 8.4790 63.8560 8.5410 64.5570 ;
        RECT 8.4650 64.1655 8.5410 64.3190 ;
        RECT 8.4790 63.4635 8.5050 64.5570 ;
        RECT 8.4790 63.5845 8.5190 63.8240 ;
        RECT 8.4790 63.4635 8.5410 63.5525 ;
        RECT 8.1820 63.9140 8.3880 64.5570 ;
        RECT 8.3620 63.4635 8.3880 64.5570 ;
        RECT 8.1820 64.1910 8.4020 64.4490 ;
        RECT 8.1820 63.4635 8.2800 64.5570 ;
        RECT 7.7650 63.4635 7.8480 64.5570 ;
        RECT 7.7650 63.5520 7.8620 64.4875 ;
        RECT 16.4440 63.4635 16.5290 64.5570 ;
        RECT 16.3000 63.4635 16.3260 64.5570 ;
        RECT 16.1920 63.4635 16.2180 64.5570 ;
        RECT 16.0840 63.4635 16.1100 64.5570 ;
        RECT 15.9760 63.4635 16.0020 64.5570 ;
        RECT 15.8680 63.4635 15.8940 64.5570 ;
        RECT 15.7600 63.4635 15.7860 64.5570 ;
        RECT 15.6520 63.4635 15.6780 64.5570 ;
        RECT 15.5440 63.4635 15.5700 64.5570 ;
        RECT 15.4360 63.4635 15.4620 64.5570 ;
        RECT 15.3280 63.4635 15.3540 64.5570 ;
        RECT 15.2200 63.4635 15.2460 64.5570 ;
        RECT 15.1120 63.4635 15.1380 64.5570 ;
        RECT 15.0040 63.4635 15.0300 64.5570 ;
        RECT 14.8960 63.4635 14.9220 64.5570 ;
        RECT 14.7880 63.4635 14.8140 64.5570 ;
        RECT 14.6800 63.4635 14.7060 64.5570 ;
        RECT 14.5720 63.4635 14.5980 64.5570 ;
        RECT 14.4640 63.4635 14.4900 64.5570 ;
        RECT 14.3560 63.4635 14.3820 64.5570 ;
        RECT 14.2480 63.4635 14.2740 64.5570 ;
        RECT 14.1400 63.4635 14.1660 64.5570 ;
        RECT 14.0320 63.4635 14.0580 64.5570 ;
        RECT 13.9240 63.4635 13.9500 64.5570 ;
        RECT 13.8160 63.4635 13.8420 64.5570 ;
        RECT 13.7080 63.4635 13.7340 64.5570 ;
        RECT 13.6000 63.4635 13.6260 64.5570 ;
        RECT 13.4920 63.4635 13.5180 64.5570 ;
        RECT 13.3840 63.4635 13.4100 64.5570 ;
        RECT 13.2760 63.4635 13.3020 64.5570 ;
        RECT 13.1680 63.4635 13.1940 64.5570 ;
        RECT 13.0600 63.4635 13.0860 64.5570 ;
        RECT 12.9520 63.4635 12.9780 64.5570 ;
        RECT 12.8440 63.4635 12.8700 64.5570 ;
        RECT 12.7360 63.4635 12.7620 64.5570 ;
        RECT 12.6280 63.4635 12.6540 64.5570 ;
        RECT 12.5200 63.4635 12.5460 64.5570 ;
        RECT 12.4120 63.4635 12.4380 64.5570 ;
        RECT 12.3040 63.4635 12.3300 64.5570 ;
        RECT 12.1960 63.4635 12.2220 64.5570 ;
        RECT 12.0880 63.4635 12.1140 64.5570 ;
        RECT 11.9800 63.4635 12.0060 64.5570 ;
        RECT 11.8720 63.4635 11.8980 64.5570 ;
        RECT 11.7640 63.4635 11.7900 64.5570 ;
        RECT 11.6560 63.4635 11.6820 64.5570 ;
        RECT 11.5480 63.4635 11.5740 64.5570 ;
        RECT 11.4400 63.4635 11.4660 64.5570 ;
        RECT 11.3320 63.4635 11.3580 64.5570 ;
        RECT 11.2240 63.4635 11.2500 64.5570 ;
        RECT 11.1160 63.4635 11.1420 64.5570 ;
        RECT 11.0080 63.4635 11.0340 64.5570 ;
        RECT 10.9000 63.4635 10.9260 64.5570 ;
        RECT 10.7920 63.4635 10.8180 64.5570 ;
        RECT 10.6840 63.4635 10.7100 64.5570 ;
        RECT 10.5760 63.4635 10.6020 64.5570 ;
        RECT 10.4680 63.4635 10.4940 64.5570 ;
        RECT 10.3600 63.4635 10.3860 64.5570 ;
        RECT 10.2520 63.4635 10.2780 64.5570 ;
        RECT 10.1440 63.4635 10.1700 64.5570 ;
        RECT 10.0360 63.4635 10.0620 64.5570 ;
        RECT 9.9280 63.4635 9.9540 64.5570 ;
        RECT 9.8200 63.4635 9.8460 64.5570 ;
        RECT 9.7120 63.4635 9.7380 64.5570 ;
        RECT 9.6040 63.4635 9.6300 64.5570 ;
        RECT 9.4960 63.4635 9.5220 64.5570 ;
        RECT 9.3880 63.4635 9.4140 64.5570 ;
        RECT 9.1750 63.4635 9.2520 64.5570 ;
        RECT 7.2820 63.4635 7.3590 64.5570 ;
        RECT 7.1200 63.4635 7.1460 64.5570 ;
        RECT 7.0120 63.4635 7.0380 64.5570 ;
        RECT 6.9040 63.4635 6.9300 64.5570 ;
        RECT 6.7960 63.4635 6.8220 64.5570 ;
        RECT 6.6880 63.4635 6.7140 64.5570 ;
        RECT 6.5800 63.4635 6.6060 64.5570 ;
        RECT 6.4720 63.4635 6.4980 64.5570 ;
        RECT 6.3640 63.4635 6.3900 64.5570 ;
        RECT 6.2560 63.4635 6.2820 64.5570 ;
        RECT 6.1480 63.4635 6.1740 64.5570 ;
        RECT 6.0400 63.4635 6.0660 64.5570 ;
        RECT 5.9320 63.4635 5.9580 64.5570 ;
        RECT 5.8240 63.4635 5.8500 64.5570 ;
        RECT 5.7160 63.4635 5.7420 64.5570 ;
        RECT 5.6080 63.4635 5.6340 64.5570 ;
        RECT 5.5000 63.4635 5.5260 64.5570 ;
        RECT 5.3920 63.4635 5.4180 64.5570 ;
        RECT 5.2840 63.4635 5.3100 64.5570 ;
        RECT 5.1760 63.4635 5.2020 64.5570 ;
        RECT 5.0680 63.4635 5.0940 64.5570 ;
        RECT 4.9600 63.4635 4.9860 64.5570 ;
        RECT 4.8520 63.4635 4.8780 64.5570 ;
        RECT 4.7440 63.4635 4.7700 64.5570 ;
        RECT 4.6360 63.4635 4.6620 64.5570 ;
        RECT 4.5280 63.4635 4.5540 64.5570 ;
        RECT 4.4200 63.4635 4.4460 64.5570 ;
        RECT 4.3120 63.4635 4.3380 64.5570 ;
        RECT 4.2040 63.4635 4.2300 64.5570 ;
        RECT 4.0960 63.4635 4.1220 64.5570 ;
        RECT 3.9880 63.4635 4.0140 64.5570 ;
        RECT 3.8800 63.4635 3.9060 64.5570 ;
        RECT 3.7720 63.4635 3.7980 64.5570 ;
        RECT 3.6640 63.4635 3.6900 64.5570 ;
        RECT 3.5560 63.4635 3.5820 64.5570 ;
        RECT 3.4480 63.4635 3.4740 64.5570 ;
        RECT 3.3400 63.4635 3.3660 64.5570 ;
        RECT 3.2320 63.4635 3.2580 64.5570 ;
        RECT 3.1240 63.4635 3.1500 64.5570 ;
        RECT 3.0160 63.4635 3.0420 64.5570 ;
        RECT 2.9080 63.4635 2.9340 64.5570 ;
        RECT 2.8000 63.4635 2.8260 64.5570 ;
        RECT 2.6920 63.4635 2.7180 64.5570 ;
        RECT 2.5840 63.4635 2.6100 64.5570 ;
        RECT 2.4760 63.4635 2.5020 64.5570 ;
        RECT 2.3680 63.4635 2.3940 64.5570 ;
        RECT 2.2600 63.4635 2.2860 64.5570 ;
        RECT 2.1520 63.4635 2.1780 64.5570 ;
        RECT 2.0440 63.4635 2.0700 64.5570 ;
        RECT 1.9360 63.4635 1.9620 64.5570 ;
        RECT 1.8280 63.4635 1.8540 64.5570 ;
        RECT 1.7200 63.4635 1.7460 64.5570 ;
        RECT 1.6120 63.4635 1.6380 64.5570 ;
        RECT 1.5040 63.4635 1.5300 64.5570 ;
        RECT 1.3960 63.4635 1.4220 64.5570 ;
        RECT 1.2880 63.4635 1.3140 64.5570 ;
        RECT 1.1800 63.4635 1.2060 64.5570 ;
        RECT 1.0720 63.4635 1.0980 64.5570 ;
        RECT 0.9640 63.4635 0.9900 64.5570 ;
        RECT 0.8560 63.4635 0.8820 64.5570 ;
        RECT 0.7480 63.4635 0.7740 64.5570 ;
        RECT 0.6400 63.4635 0.6660 64.5570 ;
        RECT 0.5320 63.4635 0.5580 64.5570 ;
        RECT 0.4240 63.4635 0.4500 64.5570 ;
        RECT 0.3160 63.4635 0.3420 64.5570 ;
        RECT 0.2080 63.4635 0.2340 64.5570 ;
        RECT 0.0050 63.4635 0.0900 64.5570 ;
        RECT 8.6410 64.5435 8.7690 65.6370 ;
        RECT 8.6270 65.2090 8.7690 65.5315 ;
        RECT 8.4790 64.9360 8.5410 65.6370 ;
        RECT 8.4650 65.2455 8.5410 65.3990 ;
        RECT 8.4790 64.5435 8.5050 65.6370 ;
        RECT 8.4790 64.6645 8.5190 64.9040 ;
        RECT 8.4790 64.5435 8.5410 64.6325 ;
        RECT 8.1820 64.9940 8.3880 65.6370 ;
        RECT 8.3620 64.5435 8.3880 65.6370 ;
        RECT 8.1820 65.2710 8.4020 65.5290 ;
        RECT 8.1820 64.5435 8.2800 65.6370 ;
        RECT 7.7650 64.5435 7.8480 65.6370 ;
        RECT 7.7650 64.6320 7.8620 65.5675 ;
        RECT 16.4440 64.5435 16.5290 65.6370 ;
        RECT 16.3000 64.5435 16.3260 65.6370 ;
        RECT 16.1920 64.5435 16.2180 65.6370 ;
        RECT 16.0840 64.5435 16.1100 65.6370 ;
        RECT 15.9760 64.5435 16.0020 65.6370 ;
        RECT 15.8680 64.5435 15.8940 65.6370 ;
        RECT 15.7600 64.5435 15.7860 65.6370 ;
        RECT 15.6520 64.5435 15.6780 65.6370 ;
        RECT 15.5440 64.5435 15.5700 65.6370 ;
        RECT 15.4360 64.5435 15.4620 65.6370 ;
        RECT 15.3280 64.5435 15.3540 65.6370 ;
        RECT 15.2200 64.5435 15.2460 65.6370 ;
        RECT 15.1120 64.5435 15.1380 65.6370 ;
        RECT 15.0040 64.5435 15.0300 65.6370 ;
        RECT 14.8960 64.5435 14.9220 65.6370 ;
        RECT 14.7880 64.5435 14.8140 65.6370 ;
        RECT 14.6800 64.5435 14.7060 65.6370 ;
        RECT 14.5720 64.5435 14.5980 65.6370 ;
        RECT 14.4640 64.5435 14.4900 65.6370 ;
        RECT 14.3560 64.5435 14.3820 65.6370 ;
        RECT 14.2480 64.5435 14.2740 65.6370 ;
        RECT 14.1400 64.5435 14.1660 65.6370 ;
        RECT 14.0320 64.5435 14.0580 65.6370 ;
        RECT 13.9240 64.5435 13.9500 65.6370 ;
        RECT 13.8160 64.5435 13.8420 65.6370 ;
        RECT 13.7080 64.5435 13.7340 65.6370 ;
        RECT 13.6000 64.5435 13.6260 65.6370 ;
        RECT 13.4920 64.5435 13.5180 65.6370 ;
        RECT 13.3840 64.5435 13.4100 65.6370 ;
        RECT 13.2760 64.5435 13.3020 65.6370 ;
        RECT 13.1680 64.5435 13.1940 65.6370 ;
        RECT 13.0600 64.5435 13.0860 65.6370 ;
        RECT 12.9520 64.5435 12.9780 65.6370 ;
        RECT 12.8440 64.5435 12.8700 65.6370 ;
        RECT 12.7360 64.5435 12.7620 65.6370 ;
        RECT 12.6280 64.5435 12.6540 65.6370 ;
        RECT 12.5200 64.5435 12.5460 65.6370 ;
        RECT 12.4120 64.5435 12.4380 65.6370 ;
        RECT 12.3040 64.5435 12.3300 65.6370 ;
        RECT 12.1960 64.5435 12.2220 65.6370 ;
        RECT 12.0880 64.5435 12.1140 65.6370 ;
        RECT 11.9800 64.5435 12.0060 65.6370 ;
        RECT 11.8720 64.5435 11.8980 65.6370 ;
        RECT 11.7640 64.5435 11.7900 65.6370 ;
        RECT 11.6560 64.5435 11.6820 65.6370 ;
        RECT 11.5480 64.5435 11.5740 65.6370 ;
        RECT 11.4400 64.5435 11.4660 65.6370 ;
        RECT 11.3320 64.5435 11.3580 65.6370 ;
        RECT 11.2240 64.5435 11.2500 65.6370 ;
        RECT 11.1160 64.5435 11.1420 65.6370 ;
        RECT 11.0080 64.5435 11.0340 65.6370 ;
        RECT 10.9000 64.5435 10.9260 65.6370 ;
        RECT 10.7920 64.5435 10.8180 65.6370 ;
        RECT 10.6840 64.5435 10.7100 65.6370 ;
        RECT 10.5760 64.5435 10.6020 65.6370 ;
        RECT 10.4680 64.5435 10.4940 65.6370 ;
        RECT 10.3600 64.5435 10.3860 65.6370 ;
        RECT 10.2520 64.5435 10.2780 65.6370 ;
        RECT 10.1440 64.5435 10.1700 65.6370 ;
        RECT 10.0360 64.5435 10.0620 65.6370 ;
        RECT 9.9280 64.5435 9.9540 65.6370 ;
        RECT 9.8200 64.5435 9.8460 65.6370 ;
        RECT 9.7120 64.5435 9.7380 65.6370 ;
        RECT 9.6040 64.5435 9.6300 65.6370 ;
        RECT 9.4960 64.5435 9.5220 65.6370 ;
        RECT 9.3880 64.5435 9.4140 65.6370 ;
        RECT 9.1750 64.5435 9.2520 65.6370 ;
        RECT 7.2820 64.5435 7.3590 65.6370 ;
        RECT 7.1200 64.5435 7.1460 65.6370 ;
        RECT 7.0120 64.5435 7.0380 65.6370 ;
        RECT 6.9040 64.5435 6.9300 65.6370 ;
        RECT 6.7960 64.5435 6.8220 65.6370 ;
        RECT 6.6880 64.5435 6.7140 65.6370 ;
        RECT 6.5800 64.5435 6.6060 65.6370 ;
        RECT 6.4720 64.5435 6.4980 65.6370 ;
        RECT 6.3640 64.5435 6.3900 65.6370 ;
        RECT 6.2560 64.5435 6.2820 65.6370 ;
        RECT 6.1480 64.5435 6.1740 65.6370 ;
        RECT 6.0400 64.5435 6.0660 65.6370 ;
        RECT 5.9320 64.5435 5.9580 65.6370 ;
        RECT 5.8240 64.5435 5.8500 65.6370 ;
        RECT 5.7160 64.5435 5.7420 65.6370 ;
        RECT 5.6080 64.5435 5.6340 65.6370 ;
        RECT 5.5000 64.5435 5.5260 65.6370 ;
        RECT 5.3920 64.5435 5.4180 65.6370 ;
        RECT 5.2840 64.5435 5.3100 65.6370 ;
        RECT 5.1760 64.5435 5.2020 65.6370 ;
        RECT 5.0680 64.5435 5.0940 65.6370 ;
        RECT 4.9600 64.5435 4.9860 65.6370 ;
        RECT 4.8520 64.5435 4.8780 65.6370 ;
        RECT 4.7440 64.5435 4.7700 65.6370 ;
        RECT 4.6360 64.5435 4.6620 65.6370 ;
        RECT 4.5280 64.5435 4.5540 65.6370 ;
        RECT 4.4200 64.5435 4.4460 65.6370 ;
        RECT 4.3120 64.5435 4.3380 65.6370 ;
        RECT 4.2040 64.5435 4.2300 65.6370 ;
        RECT 4.0960 64.5435 4.1220 65.6370 ;
        RECT 3.9880 64.5435 4.0140 65.6370 ;
        RECT 3.8800 64.5435 3.9060 65.6370 ;
        RECT 3.7720 64.5435 3.7980 65.6370 ;
        RECT 3.6640 64.5435 3.6900 65.6370 ;
        RECT 3.5560 64.5435 3.5820 65.6370 ;
        RECT 3.4480 64.5435 3.4740 65.6370 ;
        RECT 3.3400 64.5435 3.3660 65.6370 ;
        RECT 3.2320 64.5435 3.2580 65.6370 ;
        RECT 3.1240 64.5435 3.1500 65.6370 ;
        RECT 3.0160 64.5435 3.0420 65.6370 ;
        RECT 2.9080 64.5435 2.9340 65.6370 ;
        RECT 2.8000 64.5435 2.8260 65.6370 ;
        RECT 2.6920 64.5435 2.7180 65.6370 ;
        RECT 2.5840 64.5435 2.6100 65.6370 ;
        RECT 2.4760 64.5435 2.5020 65.6370 ;
        RECT 2.3680 64.5435 2.3940 65.6370 ;
        RECT 2.2600 64.5435 2.2860 65.6370 ;
        RECT 2.1520 64.5435 2.1780 65.6370 ;
        RECT 2.0440 64.5435 2.0700 65.6370 ;
        RECT 1.9360 64.5435 1.9620 65.6370 ;
        RECT 1.8280 64.5435 1.8540 65.6370 ;
        RECT 1.7200 64.5435 1.7460 65.6370 ;
        RECT 1.6120 64.5435 1.6380 65.6370 ;
        RECT 1.5040 64.5435 1.5300 65.6370 ;
        RECT 1.3960 64.5435 1.4220 65.6370 ;
        RECT 1.2880 64.5435 1.3140 65.6370 ;
        RECT 1.1800 64.5435 1.2060 65.6370 ;
        RECT 1.0720 64.5435 1.0980 65.6370 ;
        RECT 0.9640 64.5435 0.9900 65.6370 ;
        RECT 0.8560 64.5435 0.8820 65.6370 ;
        RECT 0.7480 64.5435 0.7740 65.6370 ;
        RECT 0.6400 64.5435 0.6660 65.6370 ;
        RECT 0.5320 64.5435 0.5580 65.6370 ;
        RECT 0.4240 64.5435 0.4500 65.6370 ;
        RECT 0.3160 64.5435 0.3420 65.6370 ;
        RECT 0.2080 64.5435 0.2340 65.6370 ;
        RECT 0.0050 64.5435 0.0900 65.6370 ;
        RECT 8.6410 65.6235 8.7690 66.7170 ;
        RECT 8.6270 66.2890 8.7690 66.6115 ;
        RECT 8.4790 66.0160 8.5410 66.7170 ;
        RECT 8.4650 66.3255 8.5410 66.4790 ;
        RECT 8.4790 65.6235 8.5050 66.7170 ;
        RECT 8.4790 65.7445 8.5190 65.9840 ;
        RECT 8.4790 65.6235 8.5410 65.7125 ;
        RECT 8.1820 66.0740 8.3880 66.7170 ;
        RECT 8.3620 65.6235 8.3880 66.7170 ;
        RECT 8.1820 66.3510 8.4020 66.6090 ;
        RECT 8.1820 65.6235 8.2800 66.7170 ;
        RECT 7.7650 65.6235 7.8480 66.7170 ;
        RECT 7.7650 65.7120 7.8620 66.6475 ;
        RECT 16.4440 65.6235 16.5290 66.7170 ;
        RECT 16.3000 65.6235 16.3260 66.7170 ;
        RECT 16.1920 65.6235 16.2180 66.7170 ;
        RECT 16.0840 65.6235 16.1100 66.7170 ;
        RECT 15.9760 65.6235 16.0020 66.7170 ;
        RECT 15.8680 65.6235 15.8940 66.7170 ;
        RECT 15.7600 65.6235 15.7860 66.7170 ;
        RECT 15.6520 65.6235 15.6780 66.7170 ;
        RECT 15.5440 65.6235 15.5700 66.7170 ;
        RECT 15.4360 65.6235 15.4620 66.7170 ;
        RECT 15.3280 65.6235 15.3540 66.7170 ;
        RECT 15.2200 65.6235 15.2460 66.7170 ;
        RECT 15.1120 65.6235 15.1380 66.7170 ;
        RECT 15.0040 65.6235 15.0300 66.7170 ;
        RECT 14.8960 65.6235 14.9220 66.7170 ;
        RECT 14.7880 65.6235 14.8140 66.7170 ;
        RECT 14.6800 65.6235 14.7060 66.7170 ;
        RECT 14.5720 65.6235 14.5980 66.7170 ;
        RECT 14.4640 65.6235 14.4900 66.7170 ;
        RECT 14.3560 65.6235 14.3820 66.7170 ;
        RECT 14.2480 65.6235 14.2740 66.7170 ;
        RECT 14.1400 65.6235 14.1660 66.7170 ;
        RECT 14.0320 65.6235 14.0580 66.7170 ;
        RECT 13.9240 65.6235 13.9500 66.7170 ;
        RECT 13.8160 65.6235 13.8420 66.7170 ;
        RECT 13.7080 65.6235 13.7340 66.7170 ;
        RECT 13.6000 65.6235 13.6260 66.7170 ;
        RECT 13.4920 65.6235 13.5180 66.7170 ;
        RECT 13.3840 65.6235 13.4100 66.7170 ;
        RECT 13.2760 65.6235 13.3020 66.7170 ;
        RECT 13.1680 65.6235 13.1940 66.7170 ;
        RECT 13.0600 65.6235 13.0860 66.7170 ;
        RECT 12.9520 65.6235 12.9780 66.7170 ;
        RECT 12.8440 65.6235 12.8700 66.7170 ;
        RECT 12.7360 65.6235 12.7620 66.7170 ;
        RECT 12.6280 65.6235 12.6540 66.7170 ;
        RECT 12.5200 65.6235 12.5460 66.7170 ;
        RECT 12.4120 65.6235 12.4380 66.7170 ;
        RECT 12.3040 65.6235 12.3300 66.7170 ;
        RECT 12.1960 65.6235 12.2220 66.7170 ;
        RECT 12.0880 65.6235 12.1140 66.7170 ;
        RECT 11.9800 65.6235 12.0060 66.7170 ;
        RECT 11.8720 65.6235 11.8980 66.7170 ;
        RECT 11.7640 65.6235 11.7900 66.7170 ;
        RECT 11.6560 65.6235 11.6820 66.7170 ;
        RECT 11.5480 65.6235 11.5740 66.7170 ;
        RECT 11.4400 65.6235 11.4660 66.7170 ;
        RECT 11.3320 65.6235 11.3580 66.7170 ;
        RECT 11.2240 65.6235 11.2500 66.7170 ;
        RECT 11.1160 65.6235 11.1420 66.7170 ;
        RECT 11.0080 65.6235 11.0340 66.7170 ;
        RECT 10.9000 65.6235 10.9260 66.7170 ;
        RECT 10.7920 65.6235 10.8180 66.7170 ;
        RECT 10.6840 65.6235 10.7100 66.7170 ;
        RECT 10.5760 65.6235 10.6020 66.7170 ;
        RECT 10.4680 65.6235 10.4940 66.7170 ;
        RECT 10.3600 65.6235 10.3860 66.7170 ;
        RECT 10.2520 65.6235 10.2780 66.7170 ;
        RECT 10.1440 65.6235 10.1700 66.7170 ;
        RECT 10.0360 65.6235 10.0620 66.7170 ;
        RECT 9.9280 65.6235 9.9540 66.7170 ;
        RECT 9.8200 65.6235 9.8460 66.7170 ;
        RECT 9.7120 65.6235 9.7380 66.7170 ;
        RECT 9.6040 65.6235 9.6300 66.7170 ;
        RECT 9.4960 65.6235 9.5220 66.7170 ;
        RECT 9.3880 65.6235 9.4140 66.7170 ;
        RECT 9.1750 65.6235 9.2520 66.7170 ;
        RECT 7.2820 65.6235 7.3590 66.7170 ;
        RECT 7.1200 65.6235 7.1460 66.7170 ;
        RECT 7.0120 65.6235 7.0380 66.7170 ;
        RECT 6.9040 65.6235 6.9300 66.7170 ;
        RECT 6.7960 65.6235 6.8220 66.7170 ;
        RECT 6.6880 65.6235 6.7140 66.7170 ;
        RECT 6.5800 65.6235 6.6060 66.7170 ;
        RECT 6.4720 65.6235 6.4980 66.7170 ;
        RECT 6.3640 65.6235 6.3900 66.7170 ;
        RECT 6.2560 65.6235 6.2820 66.7170 ;
        RECT 6.1480 65.6235 6.1740 66.7170 ;
        RECT 6.0400 65.6235 6.0660 66.7170 ;
        RECT 5.9320 65.6235 5.9580 66.7170 ;
        RECT 5.8240 65.6235 5.8500 66.7170 ;
        RECT 5.7160 65.6235 5.7420 66.7170 ;
        RECT 5.6080 65.6235 5.6340 66.7170 ;
        RECT 5.5000 65.6235 5.5260 66.7170 ;
        RECT 5.3920 65.6235 5.4180 66.7170 ;
        RECT 5.2840 65.6235 5.3100 66.7170 ;
        RECT 5.1760 65.6235 5.2020 66.7170 ;
        RECT 5.0680 65.6235 5.0940 66.7170 ;
        RECT 4.9600 65.6235 4.9860 66.7170 ;
        RECT 4.8520 65.6235 4.8780 66.7170 ;
        RECT 4.7440 65.6235 4.7700 66.7170 ;
        RECT 4.6360 65.6235 4.6620 66.7170 ;
        RECT 4.5280 65.6235 4.5540 66.7170 ;
        RECT 4.4200 65.6235 4.4460 66.7170 ;
        RECT 4.3120 65.6235 4.3380 66.7170 ;
        RECT 4.2040 65.6235 4.2300 66.7170 ;
        RECT 4.0960 65.6235 4.1220 66.7170 ;
        RECT 3.9880 65.6235 4.0140 66.7170 ;
        RECT 3.8800 65.6235 3.9060 66.7170 ;
        RECT 3.7720 65.6235 3.7980 66.7170 ;
        RECT 3.6640 65.6235 3.6900 66.7170 ;
        RECT 3.5560 65.6235 3.5820 66.7170 ;
        RECT 3.4480 65.6235 3.4740 66.7170 ;
        RECT 3.3400 65.6235 3.3660 66.7170 ;
        RECT 3.2320 65.6235 3.2580 66.7170 ;
        RECT 3.1240 65.6235 3.1500 66.7170 ;
        RECT 3.0160 65.6235 3.0420 66.7170 ;
        RECT 2.9080 65.6235 2.9340 66.7170 ;
        RECT 2.8000 65.6235 2.8260 66.7170 ;
        RECT 2.6920 65.6235 2.7180 66.7170 ;
        RECT 2.5840 65.6235 2.6100 66.7170 ;
        RECT 2.4760 65.6235 2.5020 66.7170 ;
        RECT 2.3680 65.6235 2.3940 66.7170 ;
        RECT 2.2600 65.6235 2.2860 66.7170 ;
        RECT 2.1520 65.6235 2.1780 66.7170 ;
        RECT 2.0440 65.6235 2.0700 66.7170 ;
        RECT 1.9360 65.6235 1.9620 66.7170 ;
        RECT 1.8280 65.6235 1.8540 66.7170 ;
        RECT 1.7200 65.6235 1.7460 66.7170 ;
        RECT 1.6120 65.6235 1.6380 66.7170 ;
        RECT 1.5040 65.6235 1.5300 66.7170 ;
        RECT 1.3960 65.6235 1.4220 66.7170 ;
        RECT 1.2880 65.6235 1.3140 66.7170 ;
        RECT 1.1800 65.6235 1.2060 66.7170 ;
        RECT 1.0720 65.6235 1.0980 66.7170 ;
        RECT 0.9640 65.6235 0.9900 66.7170 ;
        RECT 0.8560 65.6235 0.8820 66.7170 ;
        RECT 0.7480 65.6235 0.7740 66.7170 ;
        RECT 0.6400 65.6235 0.6660 66.7170 ;
        RECT 0.5320 65.6235 0.5580 66.7170 ;
        RECT 0.4240 65.6235 0.4500 66.7170 ;
        RECT 0.3160 65.6235 0.3420 66.7170 ;
        RECT 0.2080 65.6235 0.2340 66.7170 ;
        RECT 0.0050 65.6235 0.0900 66.7170 ;
        RECT 8.6410 66.7035 8.7690 67.7970 ;
        RECT 8.6270 67.3690 8.7690 67.6915 ;
        RECT 8.4790 67.0960 8.5410 67.7970 ;
        RECT 8.4650 67.4055 8.5410 67.5590 ;
        RECT 8.4790 66.7035 8.5050 67.7970 ;
        RECT 8.4790 66.8245 8.5190 67.0640 ;
        RECT 8.4790 66.7035 8.5410 66.7925 ;
        RECT 8.1820 67.1540 8.3880 67.7970 ;
        RECT 8.3620 66.7035 8.3880 67.7970 ;
        RECT 8.1820 67.4310 8.4020 67.6890 ;
        RECT 8.1820 66.7035 8.2800 67.7970 ;
        RECT 7.7650 66.7035 7.8480 67.7970 ;
        RECT 7.7650 66.7920 7.8620 67.7275 ;
        RECT 16.4440 66.7035 16.5290 67.7970 ;
        RECT 16.3000 66.7035 16.3260 67.7970 ;
        RECT 16.1920 66.7035 16.2180 67.7970 ;
        RECT 16.0840 66.7035 16.1100 67.7970 ;
        RECT 15.9760 66.7035 16.0020 67.7970 ;
        RECT 15.8680 66.7035 15.8940 67.7970 ;
        RECT 15.7600 66.7035 15.7860 67.7970 ;
        RECT 15.6520 66.7035 15.6780 67.7970 ;
        RECT 15.5440 66.7035 15.5700 67.7970 ;
        RECT 15.4360 66.7035 15.4620 67.7970 ;
        RECT 15.3280 66.7035 15.3540 67.7970 ;
        RECT 15.2200 66.7035 15.2460 67.7970 ;
        RECT 15.1120 66.7035 15.1380 67.7970 ;
        RECT 15.0040 66.7035 15.0300 67.7970 ;
        RECT 14.8960 66.7035 14.9220 67.7970 ;
        RECT 14.7880 66.7035 14.8140 67.7970 ;
        RECT 14.6800 66.7035 14.7060 67.7970 ;
        RECT 14.5720 66.7035 14.5980 67.7970 ;
        RECT 14.4640 66.7035 14.4900 67.7970 ;
        RECT 14.3560 66.7035 14.3820 67.7970 ;
        RECT 14.2480 66.7035 14.2740 67.7970 ;
        RECT 14.1400 66.7035 14.1660 67.7970 ;
        RECT 14.0320 66.7035 14.0580 67.7970 ;
        RECT 13.9240 66.7035 13.9500 67.7970 ;
        RECT 13.8160 66.7035 13.8420 67.7970 ;
        RECT 13.7080 66.7035 13.7340 67.7970 ;
        RECT 13.6000 66.7035 13.6260 67.7970 ;
        RECT 13.4920 66.7035 13.5180 67.7970 ;
        RECT 13.3840 66.7035 13.4100 67.7970 ;
        RECT 13.2760 66.7035 13.3020 67.7970 ;
        RECT 13.1680 66.7035 13.1940 67.7970 ;
        RECT 13.0600 66.7035 13.0860 67.7970 ;
        RECT 12.9520 66.7035 12.9780 67.7970 ;
        RECT 12.8440 66.7035 12.8700 67.7970 ;
        RECT 12.7360 66.7035 12.7620 67.7970 ;
        RECT 12.6280 66.7035 12.6540 67.7970 ;
        RECT 12.5200 66.7035 12.5460 67.7970 ;
        RECT 12.4120 66.7035 12.4380 67.7970 ;
        RECT 12.3040 66.7035 12.3300 67.7970 ;
        RECT 12.1960 66.7035 12.2220 67.7970 ;
        RECT 12.0880 66.7035 12.1140 67.7970 ;
        RECT 11.9800 66.7035 12.0060 67.7970 ;
        RECT 11.8720 66.7035 11.8980 67.7970 ;
        RECT 11.7640 66.7035 11.7900 67.7970 ;
        RECT 11.6560 66.7035 11.6820 67.7970 ;
        RECT 11.5480 66.7035 11.5740 67.7970 ;
        RECT 11.4400 66.7035 11.4660 67.7970 ;
        RECT 11.3320 66.7035 11.3580 67.7970 ;
        RECT 11.2240 66.7035 11.2500 67.7970 ;
        RECT 11.1160 66.7035 11.1420 67.7970 ;
        RECT 11.0080 66.7035 11.0340 67.7970 ;
        RECT 10.9000 66.7035 10.9260 67.7970 ;
        RECT 10.7920 66.7035 10.8180 67.7970 ;
        RECT 10.6840 66.7035 10.7100 67.7970 ;
        RECT 10.5760 66.7035 10.6020 67.7970 ;
        RECT 10.4680 66.7035 10.4940 67.7970 ;
        RECT 10.3600 66.7035 10.3860 67.7970 ;
        RECT 10.2520 66.7035 10.2780 67.7970 ;
        RECT 10.1440 66.7035 10.1700 67.7970 ;
        RECT 10.0360 66.7035 10.0620 67.7970 ;
        RECT 9.9280 66.7035 9.9540 67.7970 ;
        RECT 9.8200 66.7035 9.8460 67.7970 ;
        RECT 9.7120 66.7035 9.7380 67.7970 ;
        RECT 9.6040 66.7035 9.6300 67.7970 ;
        RECT 9.4960 66.7035 9.5220 67.7970 ;
        RECT 9.3880 66.7035 9.4140 67.7970 ;
        RECT 9.1750 66.7035 9.2520 67.7970 ;
        RECT 7.2820 66.7035 7.3590 67.7970 ;
        RECT 7.1200 66.7035 7.1460 67.7970 ;
        RECT 7.0120 66.7035 7.0380 67.7970 ;
        RECT 6.9040 66.7035 6.9300 67.7970 ;
        RECT 6.7960 66.7035 6.8220 67.7970 ;
        RECT 6.6880 66.7035 6.7140 67.7970 ;
        RECT 6.5800 66.7035 6.6060 67.7970 ;
        RECT 6.4720 66.7035 6.4980 67.7970 ;
        RECT 6.3640 66.7035 6.3900 67.7970 ;
        RECT 6.2560 66.7035 6.2820 67.7970 ;
        RECT 6.1480 66.7035 6.1740 67.7970 ;
        RECT 6.0400 66.7035 6.0660 67.7970 ;
        RECT 5.9320 66.7035 5.9580 67.7970 ;
        RECT 5.8240 66.7035 5.8500 67.7970 ;
        RECT 5.7160 66.7035 5.7420 67.7970 ;
        RECT 5.6080 66.7035 5.6340 67.7970 ;
        RECT 5.5000 66.7035 5.5260 67.7970 ;
        RECT 5.3920 66.7035 5.4180 67.7970 ;
        RECT 5.2840 66.7035 5.3100 67.7970 ;
        RECT 5.1760 66.7035 5.2020 67.7970 ;
        RECT 5.0680 66.7035 5.0940 67.7970 ;
        RECT 4.9600 66.7035 4.9860 67.7970 ;
        RECT 4.8520 66.7035 4.8780 67.7970 ;
        RECT 4.7440 66.7035 4.7700 67.7970 ;
        RECT 4.6360 66.7035 4.6620 67.7970 ;
        RECT 4.5280 66.7035 4.5540 67.7970 ;
        RECT 4.4200 66.7035 4.4460 67.7970 ;
        RECT 4.3120 66.7035 4.3380 67.7970 ;
        RECT 4.2040 66.7035 4.2300 67.7970 ;
        RECT 4.0960 66.7035 4.1220 67.7970 ;
        RECT 3.9880 66.7035 4.0140 67.7970 ;
        RECT 3.8800 66.7035 3.9060 67.7970 ;
        RECT 3.7720 66.7035 3.7980 67.7970 ;
        RECT 3.6640 66.7035 3.6900 67.7970 ;
        RECT 3.5560 66.7035 3.5820 67.7970 ;
        RECT 3.4480 66.7035 3.4740 67.7970 ;
        RECT 3.3400 66.7035 3.3660 67.7970 ;
        RECT 3.2320 66.7035 3.2580 67.7970 ;
        RECT 3.1240 66.7035 3.1500 67.7970 ;
        RECT 3.0160 66.7035 3.0420 67.7970 ;
        RECT 2.9080 66.7035 2.9340 67.7970 ;
        RECT 2.8000 66.7035 2.8260 67.7970 ;
        RECT 2.6920 66.7035 2.7180 67.7970 ;
        RECT 2.5840 66.7035 2.6100 67.7970 ;
        RECT 2.4760 66.7035 2.5020 67.7970 ;
        RECT 2.3680 66.7035 2.3940 67.7970 ;
        RECT 2.2600 66.7035 2.2860 67.7970 ;
        RECT 2.1520 66.7035 2.1780 67.7970 ;
        RECT 2.0440 66.7035 2.0700 67.7970 ;
        RECT 1.9360 66.7035 1.9620 67.7970 ;
        RECT 1.8280 66.7035 1.8540 67.7970 ;
        RECT 1.7200 66.7035 1.7460 67.7970 ;
        RECT 1.6120 66.7035 1.6380 67.7970 ;
        RECT 1.5040 66.7035 1.5300 67.7970 ;
        RECT 1.3960 66.7035 1.4220 67.7970 ;
        RECT 1.2880 66.7035 1.3140 67.7970 ;
        RECT 1.1800 66.7035 1.2060 67.7970 ;
        RECT 1.0720 66.7035 1.0980 67.7970 ;
        RECT 0.9640 66.7035 0.9900 67.7970 ;
        RECT 0.8560 66.7035 0.8820 67.7970 ;
        RECT 0.7480 66.7035 0.7740 67.7970 ;
        RECT 0.6400 66.7035 0.6660 67.7970 ;
        RECT 0.5320 66.7035 0.5580 67.7970 ;
        RECT 0.4240 66.7035 0.4500 67.7970 ;
        RECT 0.3160 66.7035 0.3420 67.7970 ;
        RECT 0.2080 66.7035 0.2340 67.7970 ;
        RECT 0.0050 66.7035 0.0900 67.7970 ;
        RECT 8.6410 67.7835 8.7690 68.8770 ;
        RECT 8.6270 68.4490 8.7690 68.7715 ;
        RECT 8.4790 68.1760 8.5410 68.8770 ;
        RECT 8.4650 68.4855 8.5410 68.6390 ;
        RECT 8.4790 67.7835 8.5050 68.8770 ;
        RECT 8.4790 67.9045 8.5190 68.1440 ;
        RECT 8.4790 67.7835 8.5410 67.8725 ;
        RECT 8.1820 68.2340 8.3880 68.8770 ;
        RECT 8.3620 67.7835 8.3880 68.8770 ;
        RECT 8.1820 68.5110 8.4020 68.7690 ;
        RECT 8.1820 67.7835 8.2800 68.8770 ;
        RECT 7.7650 67.7835 7.8480 68.8770 ;
        RECT 7.7650 67.8720 7.8620 68.8075 ;
        RECT 16.4440 67.7835 16.5290 68.8770 ;
        RECT 16.3000 67.7835 16.3260 68.8770 ;
        RECT 16.1920 67.7835 16.2180 68.8770 ;
        RECT 16.0840 67.7835 16.1100 68.8770 ;
        RECT 15.9760 67.7835 16.0020 68.8770 ;
        RECT 15.8680 67.7835 15.8940 68.8770 ;
        RECT 15.7600 67.7835 15.7860 68.8770 ;
        RECT 15.6520 67.7835 15.6780 68.8770 ;
        RECT 15.5440 67.7835 15.5700 68.8770 ;
        RECT 15.4360 67.7835 15.4620 68.8770 ;
        RECT 15.3280 67.7835 15.3540 68.8770 ;
        RECT 15.2200 67.7835 15.2460 68.8770 ;
        RECT 15.1120 67.7835 15.1380 68.8770 ;
        RECT 15.0040 67.7835 15.0300 68.8770 ;
        RECT 14.8960 67.7835 14.9220 68.8770 ;
        RECT 14.7880 67.7835 14.8140 68.8770 ;
        RECT 14.6800 67.7835 14.7060 68.8770 ;
        RECT 14.5720 67.7835 14.5980 68.8770 ;
        RECT 14.4640 67.7835 14.4900 68.8770 ;
        RECT 14.3560 67.7835 14.3820 68.8770 ;
        RECT 14.2480 67.7835 14.2740 68.8770 ;
        RECT 14.1400 67.7835 14.1660 68.8770 ;
        RECT 14.0320 67.7835 14.0580 68.8770 ;
        RECT 13.9240 67.7835 13.9500 68.8770 ;
        RECT 13.8160 67.7835 13.8420 68.8770 ;
        RECT 13.7080 67.7835 13.7340 68.8770 ;
        RECT 13.6000 67.7835 13.6260 68.8770 ;
        RECT 13.4920 67.7835 13.5180 68.8770 ;
        RECT 13.3840 67.7835 13.4100 68.8770 ;
        RECT 13.2760 67.7835 13.3020 68.8770 ;
        RECT 13.1680 67.7835 13.1940 68.8770 ;
        RECT 13.0600 67.7835 13.0860 68.8770 ;
        RECT 12.9520 67.7835 12.9780 68.8770 ;
        RECT 12.8440 67.7835 12.8700 68.8770 ;
        RECT 12.7360 67.7835 12.7620 68.8770 ;
        RECT 12.6280 67.7835 12.6540 68.8770 ;
        RECT 12.5200 67.7835 12.5460 68.8770 ;
        RECT 12.4120 67.7835 12.4380 68.8770 ;
        RECT 12.3040 67.7835 12.3300 68.8770 ;
        RECT 12.1960 67.7835 12.2220 68.8770 ;
        RECT 12.0880 67.7835 12.1140 68.8770 ;
        RECT 11.9800 67.7835 12.0060 68.8770 ;
        RECT 11.8720 67.7835 11.8980 68.8770 ;
        RECT 11.7640 67.7835 11.7900 68.8770 ;
        RECT 11.6560 67.7835 11.6820 68.8770 ;
        RECT 11.5480 67.7835 11.5740 68.8770 ;
        RECT 11.4400 67.7835 11.4660 68.8770 ;
        RECT 11.3320 67.7835 11.3580 68.8770 ;
        RECT 11.2240 67.7835 11.2500 68.8770 ;
        RECT 11.1160 67.7835 11.1420 68.8770 ;
        RECT 11.0080 67.7835 11.0340 68.8770 ;
        RECT 10.9000 67.7835 10.9260 68.8770 ;
        RECT 10.7920 67.7835 10.8180 68.8770 ;
        RECT 10.6840 67.7835 10.7100 68.8770 ;
        RECT 10.5760 67.7835 10.6020 68.8770 ;
        RECT 10.4680 67.7835 10.4940 68.8770 ;
        RECT 10.3600 67.7835 10.3860 68.8770 ;
        RECT 10.2520 67.7835 10.2780 68.8770 ;
        RECT 10.1440 67.7835 10.1700 68.8770 ;
        RECT 10.0360 67.7835 10.0620 68.8770 ;
        RECT 9.9280 67.7835 9.9540 68.8770 ;
        RECT 9.8200 67.7835 9.8460 68.8770 ;
        RECT 9.7120 67.7835 9.7380 68.8770 ;
        RECT 9.6040 67.7835 9.6300 68.8770 ;
        RECT 9.4960 67.7835 9.5220 68.8770 ;
        RECT 9.3880 67.7835 9.4140 68.8770 ;
        RECT 9.1750 67.7835 9.2520 68.8770 ;
        RECT 7.2820 67.7835 7.3590 68.8770 ;
        RECT 7.1200 67.7835 7.1460 68.8770 ;
        RECT 7.0120 67.7835 7.0380 68.8770 ;
        RECT 6.9040 67.7835 6.9300 68.8770 ;
        RECT 6.7960 67.7835 6.8220 68.8770 ;
        RECT 6.6880 67.7835 6.7140 68.8770 ;
        RECT 6.5800 67.7835 6.6060 68.8770 ;
        RECT 6.4720 67.7835 6.4980 68.8770 ;
        RECT 6.3640 67.7835 6.3900 68.8770 ;
        RECT 6.2560 67.7835 6.2820 68.8770 ;
        RECT 6.1480 67.7835 6.1740 68.8770 ;
        RECT 6.0400 67.7835 6.0660 68.8770 ;
        RECT 5.9320 67.7835 5.9580 68.8770 ;
        RECT 5.8240 67.7835 5.8500 68.8770 ;
        RECT 5.7160 67.7835 5.7420 68.8770 ;
        RECT 5.6080 67.7835 5.6340 68.8770 ;
        RECT 5.5000 67.7835 5.5260 68.8770 ;
        RECT 5.3920 67.7835 5.4180 68.8770 ;
        RECT 5.2840 67.7835 5.3100 68.8770 ;
        RECT 5.1760 67.7835 5.2020 68.8770 ;
        RECT 5.0680 67.7835 5.0940 68.8770 ;
        RECT 4.9600 67.7835 4.9860 68.8770 ;
        RECT 4.8520 67.7835 4.8780 68.8770 ;
        RECT 4.7440 67.7835 4.7700 68.8770 ;
        RECT 4.6360 67.7835 4.6620 68.8770 ;
        RECT 4.5280 67.7835 4.5540 68.8770 ;
        RECT 4.4200 67.7835 4.4460 68.8770 ;
        RECT 4.3120 67.7835 4.3380 68.8770 ;
        RECT 4.2040 67.7835 4.2300 68.8770 ;
        RECT 4.0960 67.7835 4.1220 68.8770 ;
        RECT 3.9880 67.7835 4.0140 68.8770 ;
        RECT 3.8800 67.7835 3.9060 68.8770 ;
        RECT 3.7720 67.7835 3.7980 68.8770 ;
        RECT 3.6640 67.7835 3.6900 68.8770 ;
        RECT 3.5560 67.7835 3.5820 68.8770 ;
        RECT 3.4480 67.7835 3.4740 68.8770 ;
        RECT 3.3400 67.7835 3.3660 68.8770 ;
        RECT 3.2320 67.7835 3.2580 68.8770 ;
        RECT 3.1240 67.7835 3.1500 68.8770 ;
        RECT 3.0160 67.7835 3.0420 68.8770 ;
        RECT 2.9080 67.7835 2.9340 68.8770 ;
        RECT 2.8000 67.7835 2.8260 68.8770 ;
        RECT 2.6920 67.7835 2.7180 68.8770 ;
        RECT 2.5840 67.7835 2.6100 68.8770 ;
        RECT 2.4760 67.7835 2.5020 68.8770 ;
        RECT 2.3680 67.7835 2.3940 68.8770 ;
        RECT 2.2600 67.7835 2.2860 68.8770 ;
        RECT 2.1520 67.7835 2.1780 68.8770 ;
        RECT 2.0440 67.7835 2.0700 68.8770 ;
        RECT 1.9360 67.7835 1.9620 68.8770 ;
        RECT 1.8280 67.7835 1.8540 68.8770 ;
        RECT 1.7200 67.7835 1.7460 68.8770 ;
        RECT 1.6120 67.7835 1.6380 68.8770 ;
        RECT 1.5040 67.7835 1.5300 68.8770 ;
        RECT 1.3960 67.7835 1.4220 68.8770 ;
        RECT 1.2880 67.7835 1.3140 68.8770 ;
        RECT 1.1800 67.7835 1.2060 68.8770 ;
        RECT 1.0720 67.7835 1.0980 68.8770 ;
        RECT 0.9640 67.7835 0.9900 68.8770 ;
        RECT 0.8560 67.7835 0.8820 68.8770 ;
        RECT 0.7480 67.7835 0.7740 68.8770 ;
        RECT 0.6400 67.7835 0.6660 68.8770 ;
        RECT 0.5320 67.7835 0.5580 68.8770 ;
        RECT 0.4240 67.7835 0.4500 68.8770 ;
        RECT 0.3160 67.7835 0.3420 68.8770 ;
        RECT 0.2080 67.7835 0.2340 68.8770 ;
        RECT 0.0050 67.7835 0.0900 68.8770 ;
        RECT 8.6410 68.8635 8.7690 69.9570 ;
        RECT 8.6270 69.5290 8.7690 69.8515 ;
        RECT 8.4790 69.2560 8.5410 69.9570 ;
        RECT 8.4650 69.5655 8.5410 69.7190 ;
        RECT 8.4790 68.8635 8.5050 69.9570 ;
        RECT 8.4790 68.9845 8.5190 69.2240 ;
        RECT 8.4790 68.8635 8.5410 68.9525 ;
        RECT 8.1820 69.3140 8.3880 69.9570 ;
        RECT 8.3620 68.8635 8.3880 69.9570 ;
        RECT 8.1820 69.5910 8.4020 69.8490 ;
        RECT 8.1820 68.8635 8.2800 69.9570 ;
        RECT 7.7650 68.8635 7.8480 69.9570 ;
        RECT 7.7650 68.9520 7.8620 69.8875 ;
        RECT 16.4440 68.8635 16.5290 69.9570 ;
        RECT 16.3000 68.8635 16.3260 69.9570 ;
        RECT 16.1920 68.8635 16.2180 69.9570 ;
        RECT 16.0840 68.8635 16.1100 69.9570 ;
        RECT 15.9760 68.8635 16.0020 69.9570 ;
        RECT 15.8680 68.8635 15.8940 69.9570 ;
        RECT 15.7600 68.8635 15.7860 69.9570 ;
        RECT 15.6520 68.8635 15.6780 69.9570 ;
        RECT 15.5440 68.8635 15.5700 69.9570 ;
        RECT 15.4360 68.8635 15.4620 69.9570 ;
        RECT 15.3280 68.8635 15.3540 69.9570 ;
        RECT 15.2200 68.8635 15.2460 69.9570 ;
        RECT 15.1120 68.8635 15.1380 69.9570 ;
        RECT 15.0040 68.8635 15.0300 69.9570 ;
        RECT 14.8960 68.8635 14.9220 69.9570 ;
        RECT 14.7880 68.8635 14.8140 69.9570 ;
        RECT 14.6800 68.8635 14.7060 69.9570 ;
        RECT 14.5720 68.8635 14.5980 69.9570 ;
        RECT 14.4640 68.8635 14.4900 69.9570 ;
        RECT 14.3560 68.8635 14.3820 69.9570 ;
        RECT 14.2480 68.8635 14.2740 69.9570 ;
        RECT 14.1400 68.8635 14.1660 69.9570 ;
        RECT 14.0320 68.8635 14.0580 69.9570 ;
        RECT 13.9240 68.8635 13.9500 69.9570 ;
        RECT 13.8160 68.8635 13.8420 69.9570 ;
        RECT 13.7080 68.8635 13.7340 69.9570 ;
        RECT 13.6000 68.8635 13.6260 69.9570 ;
        RECT 13.4920 68.8635 13.5180 69.9570 ;
        RECT 13.3840 68.8635 13.4100 69.9570 ;
        RECT 13.2760 68.8635 13.3020 69.9570 ;
        RECT 13.1680 68.8635 13.1940 69.9570 ;
        RECT 13.0600 68.8635 13.0860 69.9570 ;
        RECT 12.9520 68.8635 12.9780 69.9570 ;
        RECT 12.8440 68.8635 12.8700 69.9570 ;
        RECT 12.7360 68.8635 12.7620 69.9570 ;
        RECT 12.6280 68.8635 12.6540 69.9570 ;
        RECT 12.5200 68.8635 12.5460 69.9570 ;
        RECT 12.4120 68.8635 12.4380 69.9570 ;
        RECT 12.3040 68.8635 12.3300 69.9570 ;
        RECT 12.1960 68.8635 12.2220 69.9570 ;
        RECT 12.0880 68.8635 12.1140 69.9570 ;
        RECT 11.9800 68.8635 12.0060 69.9570 ;
        RECT 11.8720 68.8635 11.8980 69.9570 ;
        RECT 11.7640 68.8635 11.7900 69.9570 ;
        RECT 11.6560 68.8635 11.6820 69.9570 ;
        RECT 11.5480 68.8635 11.5740 69.9570 ;
        RECT 11.4400 68.8635 11.4660 69.9570 ;
        RECT 11.3320 68.8635 11.3580 69.9570 ;
        RECT 11.2240 68.8635 11.2500 69.9570 ;
        RECT 11.1160 68.8635 11.1420 69.9570 ;
        RECT 11.0080 68.8635 11.0340 69.9570 ;
        RECT 10.9000 68.8635 10.9260 69.9570 ;
        RECT 10.7920 68.8635 10.8180 69.9570 ;
        RECT 10.6840 68.8635 10.7100 69.9570 ;
        RECT 10.5760 68.8635 10.6020 69.9570 ;
        RECT 10.4680 68.8635 10.4940 69.9570 ;
        RECT 10.3600 68.8635 10.3860 69.9570 ;
        RECT 10.2520 68.8635 10.2780 69.9570 ;
        RECT 10.1440 68.8635 10.1700 69.9570 ;
        RECT 10.0360 68.8635 10.0620 69.9570 ;
        RECT 9.9280 68.8635 9.9540 69.9570 ;
        RECT 9.8200 68.8635 9.8460 69.9570 ;
        RECT 9.7120 68.8635 9.7380 69.9570 ;
        RECT 9.6040 68.8635 9.6300 69.9570 ;
        RECT 9.4960 68.8635 9.5220 69.9570 ;
        RECT 9.3880 68.8635 9.4140 69.9570 ;
        RECT 9.1750 68.8635 9.2520 69.9570 ;
        RECT 7.2820 68.8635 7.3590 69.9570 ;
        RECT 7.1200 68.8635 7.1460 69.9570 ;
        RECT 7.0120 68.8635 7.0380 69.9570 ;
        RECT 6.9040 68.8635 6.9300 69.9570 ;
        RECT 6.7960 68.8635 6.8220 69.9570 ;
        RECT 6.6880 68.8635 6.7140 69.9570 ;
        RECT 6.5800 68.8635 6.6060 69.9570 ;
        RECT 6.4720 68.8635 6.4980 69.9570 ;
        RECT 6.3640 68.8635 6.3900 69.9570 ;
        RECT 6.2560 68.8635 6.2820 69.9570 ;
        RECT 6.1480 68.8635 6.1740 69.9570 ;
        RECT 6.0400 68.8635 6.0660 69.9570 ;
        RECT 5.9320 68.8635 5.9580 69.9570 ;
        RECT 5.8240 68.8635 5.8500 69.9570 ;
        RECT 5.7160 68.8635 5.7420 69.9570 ;
        RECT 5.6080 68.8635 5.6340 69.9570 ;
        RECT 5.5000 68.8635 5.5260 69.9570 ;
        RECT 5.3920 68.8635 5.4180 69.9570 ;
        RECT 5.2840 68.8635 5.3100 69.9570 ;
        RECT 5.1760 68.8635 5.2020 69.9570 ;
        RECT 5.0680 68.8635 5.0940 69.9570 ;
        RECT 4.9600 68.8635 4.9860 69.9570 ;
        RECT 4.8520 68.8635 4.8780 69.9570 ;
        RECT 4.7440 68.8635 4.7700 69.9570 ;
        RECT 4.6360 68.8635 4.6620 69.9570 ;
        RECT 4.5280 68.8635 4.5540 69.9570 ;
        RECT 4.4200 68.8635 4.4460 69.9570 ;
        RECT 4.3120 68.8635 4.3380 69.9570 ;
        RECT 4.2040 68.8635 4.2300 69.9570 ;
        RECT 4.0960 68.8635 4.1220 69.9570 ;
        RECT 3.9880 68.8635 4.0140 69.9570 ;
        RECT 3.8800 68.8635 3.9060 69.9570 ;
        RECT 3.7720 68.8635 3.7980 69.9570 ;
        RECT 3.6640 68.8635 3.6900 69.9570 ;
        RECT 3.5560 68.8635 3.5820 69.9570 ;
        RECT 3.4480 68.8635 3.4740 69.9570 ;
        RECT 3.3400 68.8635 3.3660 69.9570 ;
        RECT 3.2320 68.8635 3.2580 69.9570 ;
        RECT 3.1240 68.8635 3.1500 69.9570 ;
        RECT 3.0160 68.8635 3.0420 69.9570 ;
        RECT 2.9080 68.8635 2.9340 69.9570 ;
        RECT 2.8000 68.8635 2.8260 69.9570 ;
        RECT 2.6920 68.8635 2.7180 69.9570 ;
        RECT 2.5840 68.8635 2.6100 69.9570 ;
        RECT 2.4760 68.8635 2.5020 69.9570 ;
        RECT 2.3680 68.8635 2.3940 69.9570 ;
        RECT 2.2600 68.8635 2.2860 69.9570 ;
        RECT 2.1520 68.8635 2.1780 69.9570 ;
        RECT 2.0440 68.8635 2.0700 69.9570 ;
        RECT 1.9360 68.8635 1.9620 69.9570 ;
        RECT 1.8280 68.8635 1.8540 69.9570 ;
        RECT 1.7200 68.8635 1.7460 69.9570 ;
        RECT 1.6120 68.8635 1.6380 69.9570 ;
        RECT 1.5040 68.8635 1.5300 69.9570 ;
        RECT 1.3960 68.8635 1.4220 69.9570 ;
        RECT 1.2880 68.8635 1.3140 69.9570 ;
        RECT 1.1800 68.8635 1.2060 69.9570 ;
        RECT 1.0720 68.8635 1.0980 69.9570 ;
        RECT 0.9640 68.8635 0.9900 69.9570 ;
        RECT 0.8560 68.8635 0.8820 69.9570 ;
        RECT 0.7480 68.8635 0.7740 69.9570 ;
        RECT 0.6400 68.8635 0.6660 69.9570 ;
        RECT 0.5320 68.8635 0.5580 69.9570 ;
        RECT 0.4240 68.8635 0.4500 69.9570 ;
        RECT 0.3160 68.8635 0.3420 69.9570 ;
        RECT 0.2080 68.8635 0.2340 69.9570 ;
        RECT 0.0050 68.8635 0.0900 69.9570 ;
        RECT 8.6410 69.9435 8.7690 71.0370 ;
        RECT 8.6270 70.6090 8.7690 70.9315 ;
        RECT 8.4790 70.3360 8.5410 71.0370 ;
        RECT 8.4650 70.6455 8.5410 70.7990 ;
        RECT 8.4790 69.9435 8.5050 71.0370 ;
        RECT 8.4790 70.0645 8.5190 70.3040 ;
        RECT 8.4790 69.9435 8.5410 70.0325 ;
        RECT 8.1820 70.3940 8.3880 71.0370 ;
        RECT 8.3620 69.9435 8.3880 71.0370 ;
        RECT 8.1820 70.6710 8.4020 70.9290 ;
        RECT 8.1820 69.9435 8.2800 71.0370 ;
        RECT 7.7650 69.9435 7.8480 71.0370 ;
        RECT 7.7650 70.0320 7.8620 70.9675 ;
        RECT 16.4440 69.9435 16.5290 71.0370 ;
        RECT 16.3000 69.9435 16.3260 71.0370 ;
        RECT 16.1920 69.9435 16.2180 71.0370 ;
        RECT 16.0840 69.9435 16.1100 71.0370 ;
        RECT 15.9760 69.9435 16.0020 71.0370 ;
        RECT 15.8680 69.9435 15.8940 71.0370 ;
        RECT 15.7600 69.9435 15.7860 71.0370 ;
        RECT 15.6520 69.9435 15.6780 71.0370 ;
        RECT 15.5440 69.9435 15.5700 71.0370 ;
        RECT 15.4360 69.9435 15.4620 71.0370 ;
        RECT 15.3280 69.9435 15.3540 71.0370 ;
        RECT 15.2200 69.9435 15.2460 71.0370 ;
        RECT 15.1120 69.9435 15.1380 71.0370 ;
        RECT 15.0040 69.9435 15.0300 71.0370 ;
        RECT 14.8960 69.9435 14.9220 71.0370 ;
        RECT 14.7880 69.9435 14.8140 71.0370 ;
        RECT 14.6800 69.9435 14.7060 71.0370 ;
        RECT 14.5720 69.9435 14.5980 71.0370 ;
        RECT 14.4640 69.9435 14.4900 71.0370 ;
        RECT 14.3560 69.9435 14.3820 71.0370 ;
        RECT 14.2480 69.9435 14.2740 71.0370 ;
        RECT 14.1400 69.9435 14.1660 71.0370 ;
        RECT 14.0320 69.9435 14.0580 71.0370 ;
        RECT 13.9240 69.9435 13.9500 71.0370 ;
        RECT 13.8160 69.9435 13.8420 71.0370 ;
        RECT 13.7080 69.9435 13.7340 71.0370 ;
        RECT 13.6000 69.9435 13.6260 71.0370 ;
        RECT 13.4920 69.9435 13.5180 71.0370 ;
        RECT 13.3840 69.9435 13.4100 71.0370 ;
        RECT 13.2760 69.9435 13.3020 71.0370 ;
        RECT 13.1680 69.9435 13.1940 71.0370 ;
        RECT 13.0600 69.9435 13.0860 71.0370 ;
        RECT 12.9520 69.9435 12.9780 71.0370 ;
        RECT 12.8440 69.9435 12.8700 71.0370 ;
        RECT 12.7360 69.9435 12.7620 71.0370 ;
        RECT 12.6280 69.9435 12.6540 71.0370 ;
        RECT 12.5200 69.9435 12.5460 71.0370 ;
        RECT 12.4120 69.9435 12.4380 71.0370 ;
        RECT 12.3040 69.9435 12.3300 71.0370 ;
        RECT 12.1960 69.9435 12.2220 71.0370 ;
        RECT 12.0880 69.9435 12.1140 71.0370 ;
        RECT 11.9800 69.9435 12.0060 71.0370 ;
        RECT 11.8720 69.9435 11.8980 71.0370 ;
        RECT 11.7640 69.9435 11.7900 71.0370 ;
        RECT 11.6560 69.9435 11.6820 71.0370 ;
        RECT 11.5480 69.9435 11.5740 71.0370 ;
        RECT 11.4400 69.9435 11.4660 71.0370 ;
        RECT 11.3320 69.9435 11.3580 71.0370 ;
        RECT 11.2240 69.9435 11.2500 71.0370 ;
        RECT 11.1160 69.9435 11.1420 71.0370 ;
        RECT 11.0080 69.9435 11.0340 71.0370 ;
        RECT 10.9000 69.9435 10.9260 71.0370 ;
        RECT 10.7920 69.9435 10.8180 71.0370 ;
        RECT 10.6840 69.9435 10.7100 71.0370 ;
        RECT 10.5760 69.9435 10.6020 71.0370 ;
        RECT 10.4680 69.9435 10.4940 71.0370 ;
        RECT 10.3600 69.9435 10.3860 71.0370 ;
        RECT 10.2520 69.9435 10.2780 71.0370 ;
        RECT 10.1440 69.9435 10.1700 71.0370 ;
        RECT 10.0360 69.9435 10.0620 71.0370 ;
        RECT 9.9280 69.9435 9.9540 71.0370 ;
        RECT 9.8200 69.9435 9.8460 71.0370 ;
        RECT 9.7120 69.9435 9.7380 71.0370 ;
        RECT 9.6040 69.9435 9.6300 71.0370 ;
        RECT 9.4960 69.9435 9.5220 71.0370 ;
        RECT 9.3880 69.9435 9.4140 71.0370 ;
        RECT 9.1750 69.9435 9.2520 71.0370 ;
        RECT 7.2820 69.9435 7.3590 71.0370 ;
        RECT 7.1200 69.9435 7.1460 71.0370 ;
        RECT 7.0120 69.9435 7.0380 71.0370 ;
        RECT 6.9040 69.9435 6.9300 71.0370 ;
        RECT 6.7960 69.9435 6.8220 71.0370 ;
        RECT 6.6880 69.9435 6.7140 71.0370 ;
        RECT 6.5800 69.9435 6.6060 71.0370 ;
        RECT 6.4720 69.9435 6.4980 71.0370 ;
        RECT 6.3640 69.9435 6.3900 71.0370 ;
        RECT 6.2560 69.9435 6.2820 71.0370 ;
        RECT 6.1480 69.9435 6.1740 71.0370 ;
        RECT 6.0400 69.9435 6.0660 71.0370 ;
        RECT 5.9320 69.9435 5.9580 71.0370 ;
        RECT 5.8240 69.9435 5.8500 71.0370 ;
        RECT 5.7160 69.9435 5.7420 71.0370 ;
        RECT 5.6080 69.9435 5.6340 71.0370 ;
        RECT 5.5000 69.9435 5.5260 71.0370 ;
        RECT 5.3920 69.9435 5.4180 71.0370 ;
        RECT 5.2840 69.9435 5.3100 71.0370 ;
        RECT 5.1760 69.9435 5.2020 71.0370 ;
        RECT 5.0680 69.9435 5.0940 71.0370 ;
        RECT 4.9600 69.9435 4.9860 71.0370 ;
        RECT 4.8520 69.9435 4.8780 71.0370 ;
        RECT 4.7440 69.9435 4.7700 71.0370 ;
        RECT 4.6360 69.9435 4.6620 71.0370 ;
        RECT 4.5280 69.9435 4.5540 71.0370 ;
        RECT 4.4200 69.9435 4.4460 71.0370 ;
        RECT 4.3120 69.9435 4.3380 71.0370 ;
        RECT 4.2040 69.9435 4.2300 71.0370 ;
        RECT 4.0960 69.9435 4.1220 71.0370 ;
        RECT 3.9880 69.9435 4.0140 71.0370 ;
        RECT 3.8800 69.9435 3.9060 71.0370 ;
        RECT 3.7720 69.9435 3.7980 71.0370 ;
        RECT 3.6640 69.9435 3.6900 71.0370 ;
        RECT 3.5560 69.9435 3.5820 71.0370 ;
        RECT 3.4480 69.9435 3.4740 71.0370 ;
        RECT 3.3400 69.9435 3.3660 71.0370 ;
        RECT 3.2320 69.9435 3.2580 71.0370 ;
        RECT 3.1240 69.9435 3.1500 71.0370 ;
        RECT 3.0160 69.9435 3.0420 71.0370 ;
        RECT 2.9080 69.9435 2.9340 71.0370 ;
        RECT 2.8000 69.9435 2.8260 71.0370 ;
        RECT 2.6920 69.9435 2.7180 71.0370 ;
        RECT 2.5840 69.9435 2.6100 71.0370 ;
        RECT 2.4760 69.9435 2.5020 71.0370 ;
        RECT 2.3680 69.9435 2.3940 71.0370 ;
        RECT 2.2600 69.9435 2.2860 71.0370 ;
        RECT 2.1520 69.9435 2.1780 71.0370 ;
        RECT 2.0440 69.9435 2.0700 71.0370 ;
        RECT 1.9360 69.9435 1.9620 71.0370 ;
        RECT 1.8280 69.9435 1.8540 71.0370 ;
        RECT 1.7200 69.9435 1.7460 71.0370 ;
        RECT 1.6120 69.9435 1.6380 71.0370 ;
        RECT 1.5040 69.9435 1.5300 71.0370 ;
        RECT 1.3960 69.9435 1.4220 71.0370 ;
        RECT 1.2880 69.9435 1.3140 71.0370 ;
        RECT 1.1800 69.9435 1.2060 71.0370 ;
        RECT 1.0720 69.9435 1.0980 71.0370 ;
        RECT 0.9640 69.9435 0.9900 71.0370 ;
        RECT 0.8560 69.9435 0.8820 71.0370 ;
        RECT 0.7480 69.9435 0.7740 71.0370 ;
        RECT 0.6400 69.9435 0.6660 71.0370 ;
        RECT 0.5320 69.9435 0.5580 71.0370 ;
        RECT 0.4240 69.9435 0.4500 71.0370 ;
        RECT 0.3160 69.9435 0.3420 71.0370 ;
        RECT 0.2080 69.9435 0.2340 71.0370 ;
        RECT 0.0050 69.9435 0.0900 71.0370 ;
        RECT 8.6410 71.0235 8.7690 72.1170 ;
        RECT 8.6270 71.6890 8.7690 72.0115 ;
        RECT 8.4790 71.4160 8.5410 72.1170 ;
        RECT 8.4650 71.7255 8.5410 71.8790 ;
        RECT 8.4790 71.0235 8.5050 72.1170 ;
        RECT 8.4790 71.1445 8.5190 71.3840 ;
        RECT 8.4790 71.0235 8.5410 71.1125 ;
        RECT 8.1820 71.4740 8.3880 72.1170 ;
        RECT 8.3620 71.0235 8.3880 72.1170 ;
        RECT 8.1820 71.7510 8.4020 72.0090 ;
        RECT 8.1820 71.0235 8.2800 72.1170 ;
        RECT 7.7650 71.0235 7.8480 72.1170 ;
        RECT 7.7650 71.1120 7.8620 72.0475 ;
        RECT 16.4440 71.0235 16.5290 72.1170 ;
        RECT 16.3000 71.0235 16.3260 72.1170 ;
        RECT 16.1920 71.0235 16.2180 72.1170 ;
        RECT 16.0840 71.0235 16.1100 72.1170 ;
        RECT 15.9760 71.0235 16.0020 72.1170 ;
        RECT 15.8680 71.0235 15.8940 72.1170 ;
        RECT 15.7600 71.0235 15.7860 72.1170 ;
        RECT 15.6520 71.0235 15.6780 72.1170 ;
        RECT 15.5440 71.0235 15.5700 72.1170 ;
        RECT 15.4360 71.0235 15.4620 72.1170 ;
        RECT 15.3280 71.0235 15.3540 72.1170 ;
        RECT 15.2200 71.0235 15.2460 72.1170 ;
        RECT 15.1120 71.0235 15.1380 72.1170 ;
        RECT 15.0040 71.0235 15.0300 72.1170 ;
        RECT 14.8960 71.0235 14.9220 72.1170 ;
        RECT 14.7880 71.0235 14.8140 72.1170 ;
        RECT 14.6800 71.0235 14.7060 72.1170 ;
        RECT 14.5720 71.0235 14.5980 72.1170 ;
        RECT 14.4640 71.0235 14.4900 72.1170 ;
        RECT 14.3560 71.0235 14.3820 72.1170 ;
        RECT 14.2480 71.0235 14.2740 72.1170 ;
        RECT 14.1400 71.0235 14.1660 72.1170 ;
        RECT 14.0320 71.0235 14.0580 72.1170 ;
        RECT 13.9240 71.0235 13.9500 72.1170 ;
        RECT 13.8160 71.0235 13.8420 72.1170 ;
        RECT 13.7080 71.0235 13.7340 72.1170 ;
        RECT 13.6000 71.0235 13.6260 72.1170 ;
        RECT 13.4920 71.0235 13.5180 72.1170 ;
        RECT 13.3840 71.0235 13.4100 72.1170 ;
        RECT 13.2760 71.0235 13.3020 72.1170 ;
        RECT 13.1680 71.0235 13.1940 72.1170 ;
        RECT 13.0600 71.0235 13.0860 72.1170 ;
        RECT 12.9520 71.0235 12.9780 72.1170 ;
        RECT 12.8440 71.0235 12.8700 72.1170 ;
        RECT 12.7360 71.0235 12.7620 72.1170 ;
        RECT 12.6280 71.0235 12.6540 72.1170 ;
        RECT 12.5200 71.0235 12.5460 72.1170 ;
        RECT 12.4120 71.0235 12.4380 72.1170 ;
        RECT 12.3040 71.0235 12.3300 72.1170 ;
        RECT 12.1960 71.0235 12.2220 72.1170 ;
        RECT 12.0880 71.0235 12.1140 72.1170 ;
        RECT 11.9800 71.0235 12.0060 72.1170 ;
        RECT 11.8720 71.0235 11.8980 72.1170 ;
        RECT 11.7640 71.0235 11.7900 72.1170 ;
        RECT 11.6560 71.0235 11.6820 72.1170 ;
        RECT 11.5480 71.0235 11.5740 72.1170 ;
        RECT 11.4400 71.0235 11.4660 72.1170 ;
        RECT 11.3320 71.0235 11.3580 72.1170 ;
        RECT 11.2240 71.0235 11.2500 72.1170 ;
        RECT 11.1160 71.0235 11.1420 72.1170 ;
        RECT 11.0080 71.0235 11.0340 72.1170 ;
        RECT 10.9000 71.0235 10.9260 72.1170 ;
        RECT 10.7920 71.0235 10.8180 72.1170 ;
        RECT 10.6840 71.0235 10.7100 72.1170 ;
        RECT 10.5760 71.0235 10.6020 72.1170 ;
        RECT 10.4680 71.0235 10.4940 72.1170 ;
        RECT 10.3600 71.0235 10.3860 72.1170 ;
        RECT 10.2520 71.0235 10.2780 72.1170 ;
        RECT 10.1440 71.0235 10.1700 72.1170 ;
        RECT 10.0360 71.0235 10.0620 72.1170 ;
        RECT 9.9280 71.0235 9.9540 72.1170 ;
        RECT 9.8200 71.0235 9.8460 72.1170 ;
        RECT 9.7120 71.0235 9.7380 72.1170 ;
        RECT 9.6040 71.0235 9.6300 72.1170 ;
        RECT 9.4960 71.0235 9.5220 72.1170 ;
        RECT 9.3880 71.0235 9.4140 72.1170 ;
        RECT 9.1750 71.0235 9.2520 72.1170 ;
        RECT 7.2820 71.0235 7.3590 72.1170 ;
        RECT 7.1200 71.0235 7.1460 72.1170 ;
        RECT 7.0120 71.0235 7.0380 72.1170 ;
        RECT 6.9040 71.0235 6.9300 72.1170 ;
        RECT 6.7960 71.0235 6.8220 72.1170 ;
        RECT 6.6880 71.0235 6.7140 72.1170 ;
        RECT 6.5800 71.0235 6.6060 72.1170 ;
        RECT 6.4720 71.0235 6.4980 72.1170 ;
        RECT 6.3640 71.0235 6.3900 72.1170 ;
        RECT 6.2560 71.0235 6.2820 72.1170 ;
        RECT 6.1480 71.0235 6.1740 72.1170 ;
        RECT 6.0400 71.0235 6.0660 72.1170 ;
        RECT 5.9320 71.0235 5.9580 72.1170 ;
        RECT 5.8240 71.0235 5.8500 72.1170 ;
        RECT 5.7160 71.0235 5.7420 72.1170 ;
        RECT 5.6080 71.0235 5.6340 72.1170 ;
        RECT 5.5000 71.0235 5.5260 72.1170 ;
        RECT 5.3920 71.0235 5.4180 72.1170 ;
        RECT 5.2840 71.0235 5.3100 72.1170 ;
        RECT 5.1760 71.0235 5.2020 72.1170 ;
        RECT 5.0680 71.0235 5.0940 72.1170 ;
        RECT 4.9600 71.0235 4.9860 72.1170 ;
        RECT 4.8520 71.0235 4.8780 72.1170 ;
        RECT 4.7440 71.0235 4.7700 72.1170 ;
        RECT 4.6360 71.0235 4.6620 72.1170 ;
        RECT 4.5280 71.0235 4.5540 72.1170 ;
        RECT 4.4200 71.0235 4.4460 72.1170 ;
        RECT 4.3120 71.0235 4.3380 72.1170 ;
        RECT 4.2040 71.0235 4.2300 72.1170 ;
        RECT 4.0960 71.0235 4.1220 72.1170 ;
        RECT 3.9880 71.0235 4.0140 72.1170 ;
        RECT 3.8800 71.0235 3.9060 72.1170 ;
        RECT 3.7720 71.0235 3.7980 72.1170 ;
        RECT 3.6640 71.0235 3.6900 72.1170 ;
        RECT 3.5560 71.0235 3.5820 72.1170 ;
        RECT 3.4480 71.0235 3.4740 72.1170 ;
        RECT 3.3400 71.0235 3.3660 72.1170 ;
        RECT 3.2320 71.0235 3.2580 72.1170 ;
        RECT 3.1240 71.0235 3.1500 72.1170 ;
        RECT 3.0160 71.0235 3.0420 72.1170 ;
        RECT 2.9080 71.0235 2.9340 72.1170 ;
        RECT 2.8000 71.0235 2.8260 72.1170 ;
        RECT 2.6920 71.0235 2.7180 72.1170 ;
        RECT 2.5840 71.0235 2.6100 72.1170 ;
        RECT 2.4760 71.0235 2.5020 72.1170 ;
        RECT 2.3680 71.0235 2.3940 72.1170 ;
        RECT 2.2600 71.0235 2.2860 72.1170 ;
        RECT 2.1520 71.0235 2.1780 72.1170 ;
        RECT 2.0440 71.0235 2.0700 72.1170 ;
        RECT 1.9360 71.0235 1.9620 72.1170 ;
        RECT 1.8280 71.0235 1.8540 72.1170 ;
        RECT 1.7200 71.0235 1.7460 72.1170 ;
        RECT 1.6120 71.0235 1.6380 72.1170 ;
        RECT 1.5040 71.0235 1.5300 72.1170 ;
        RECT 1.3960 71.0235 1.4220 72.1170 ;
        RECT 1.2880 71.0235 1.3140 72.1170 ;
        RECT 1.1800 71.0235 1.2060 72.1170 ;
        RECT 1.0720 71.0235 1.0980 72.1170 ;
        RECT 0.9640 71.0235 0.9900 72.1170 ;
        RECT 0.8560 71.0235 0.8820 72.1170 ;
        RECT 0.7480 71.0235 0.7740 72.1170 ;
        RECT 0.6400 71.0235 0.6660 72.1170 ;
        RECT 0.5320 71.0235 0.5580 72.1170 ;
        RECT 0.4240 71.0235 0.4500 72.1170 ;
        RECT 0.3160 71.0235 0.3420 72.1170 ;
        RECT 0.2080 71.0235 0.2340 72.1170 ;
        RECT 0.0050 71.0235 0.0900 72.1170 ;
        RECT 8.6410 72.1035 8.7690 73.1970 ;
        RECT 8.6270 72.7690 8.7690 73.0915 ;
        RECT 8.4790 72.4960 8.5410 73.1970 ;
        RECT 8.4650 72.8055 8.5410 72.9590 ;
        RECT 8.4790 72.1035 8.5050 73.1970 ;
        RECT 8.4790 72.2245 8.5190 72.4640 ;
        RECT 8.4790 72.1035 8.5410 72.1925 ;
        RECT 8.1820 72.5540 8.3880 73.1970 ;
        RECT 8.3620 72.1035 8.3880 73.1970 ;
        RECT 8.1820 72.8310 8.4020 73.0890 ;
        RECT 8.1820 72.1035 8.2800 73.1970 ;
        RECT 7.7650 72.1035 7.8480 73.1970 ;
        RECT 7.7650 72.1920 7.8620 73.1275 ;
        RECT 16.4440 72.1035 16.5290 73.1970 ;
        RECT 16.3000 72.1035 16.3260 73.1970 ;
        RECT 16.1920 72.1035 16.2180 73.1970 ;
        RECT 16.0840 72.1035 16.1100 73.1970 ;
        RECT 15.9760 72.1035 16.0020 73.1970 ;
        RECT 15.8680 72.1035 15.8940 73.1970 ;
        RECT 15.7600 72.1035 15.7860 73.1970 ;
        RECT 15.6520 72.1035 15.6780 73.1970 ;
        RECT 15.5440 72.1035 15.5700 73.1970 ;
        RECT 15.4360 72.1035 15.4620 73.1970 ;
        RECT 15.3280 72.1035 15.3540 73.1970 ;
        RECT 15.2200 72.1035 15.2460 73.1970 ;
        RECT 15.1120 72.1035 15.1380 73.1970 ;
        RECT 15.0040 72.1035 15.0300 73.1970 ;
        RECT 14.8960 72.1035 14.9220 73.1970 ;
        RECT 14.7880 72.1035 14.8140 73.1970 ;
        RECT 14.6800 72.1035 14.7060 73.1970 ;
        RECT 14.5720 72.1035 14.5980 73.1970 ;
        RECT 14.4640 72.1035 14.4900 73.1970 ;
        RECT 14.3560 72.1035 14.3820 73.1970 ;
        RECT 14.2480 72.1035 14.2740 73.1970 ;
        RECT 14.1400 72.1035 14.1660 73.1970 ;
        RECT 14.0320 72.1035 14.0580 73.1970 ;
        RECT 13.9240 72.1035 13.9500 73.1970 ;
        RECT 13.8160 72.1035 13.8420 73.1970 ;
        RECT 13.7080 72.1035 13.7340 73.1970 ;
        RECT 13.6000 72.1035 13.6260 73.1970 ;
        RECT 13.4920 72.1035 13.5180 73.1970 ;
        RECT 13.3840 72.1035 13.4100 73.1970 ;
        RECT 13.2760 72.1035 13.3020 73.1970 ;
        RECT 13.1680 72.1035 13.1940 73.1970 ;
        RECT 13.0600 72.1035 13.0860 73.1970 ;
        RECT 12.9520 72.1035 12.9780 73.1970 ;
        RECT 12.8440 72.1035 12.8700 73.1970 ;
        RECT 12.7360 72.1035 12.7620 73.1970 ;
        RECT 12.6280 72.1035 12.6540 73.1970 ;
        RECT 12.5200 72.1035 12.5460 73.1970 ;
        RECT 12.4120 72.1035 12.4380 73.1970 ;
        RECT 12.3040 72.1035 12.3300 73.1970 ;
        RECT 12.1960 72.1035 12.2220 73.1970 ;
        RECT 12.0880 72.1035 12.1140 73.1970 ;
        RECT 11.9800 72.1035 12.0060 73.1970 ;
        RECT 11.8720 72.1035 11.8980 73.1970 ;
        RECT 11.7640 72.1035 11.7900 73.1970 ;
        RECT 11.6560 72.1035 11.6820 73.1970 ;
        RECT 11.5480 72.1035 11.5740 73.1970 ;
        RECT 11.4400 72.1035 11.4660 73.1970 ;
        RECT 11.3320 72.1035 11.3580 73.1970 ;
        RECT 11.2240 72.1035 11.2500 73.1970 ;
        RECT 11.1160 72.1035 11.1420 73.1970 ;
        RECT 11.0080 72.1035 11.0340 73.1970 ;
        RECT 10.9000 72.1035 10.9260 73.1970 ;
        RECT 10.7920 72.1035 10.8180 73.1970 ;
        RECT 10.6840 72.1035 10.7100 73.1970 ;
        RECT 10.5760 72.1035 10.6020 73.1970 ;
        RECT 10.4680 72.1035 10.4940 73.1970 ;
        RECT 10.3600 72.1035 10.3860 73.1970 ;
        RECT 10.2520 72.1035 10.2780 73.1970 ;
        RECT 10.1440 72.1035 10.1700 73.1970 ;
        RECT 10.0360 72.1035 10.0620 73.1970 ;
        RECT 9.9280 72.1035 9.9540 73.1970 ;
        RECT 9.8200 72.1035 9.8460 73.1970 ;
        RECT 9.7120 72.1035 9.7380 73.1970 ;
        RECT 9.6040 72.1035 9.6300 73.1970 ;
        RECT 9.4960 72.1035 9.5220 73.1970 ;
        RECT 9.3880 72.1035 9.4140 73.1970 ;
        RECT 9.1750 72.1035 9.2520 73.1970 ;
        RECT 7.2820 72.1035 7.3590 73.1970 ;
        RECT 7.1200 72.1035 7.1460 73.1970 ;
        RECT 7.0120 72.1035 7.0380 73.1970 ;
        RECT 6.9040 72.1035 6.9300 73.1970 ;
        RECT 6.7960 72.1035 6.8220 73.1970 ;
        RECT 6.6880 72.1035 6.7140 73.1970 ;
        RECT 6.5800 72.1035 6.6060 73.1970 ;
        RECT 6.4720 72.1035 6.4980 73.1970 ;
        RECT 6.3640 72.1035 6.3900 73.1970 ;
        RECT 6.2560 72.1035 6.2820 73.1970 ;
        RECT 6.1480 72.1035 6.1740 73.1970 ;
        RECT 6.0400 72.1035 6.0660 73.1970 ;
        RECT 5.9320 72.1035 5.9580 73.1970 ;
        RECT 5.8240 72.1035 5.8500 73.1970 ;
        RECT 5.7160 72.1035 5.7420 73.1970 ;
        RECT 5.6080 72.1035 5.6340 73.1970 ;
        RECT 5.5000 72.1035 5.5260 73.1970 ;
        RECT 5.3920 72.1035 5.4180 73.1970 ;
        RECT 5.2840 72.1035 5.3100 73.1970 ;
        RECT 5.1760 72.1035 5.2020 73.1970 ;
        RECT 5.0680 72.1035 5.0940 73.1970 ;
        RECT 4.9600 72.1035 4.9860 73.1970 ;
        RECT 4.8520 72.1035 4.8780 73.1970 ;
        RECT 4.7440 72.1035 4.7700 73.1970 ;
        RECT 4.6360 72.1035 4.6620 73.1970 ;
        RECT 4.5280 72.1035 4.5540 73.1970 ;
        RECT 4.4200 72.1035 4.4460 73.1970 ;
        RECT 4.3120 72.1035 4.3380 73.1970 ;
        RECT 4.2040 72.1035 4.2300 73.1970 ;
        RECT 4.0960 72.1035 4.1220 73.1970 ;
        RECT 3.9880 72.1035 4.0140 73.1970 ;
        RECT 3.8800 72.1035 3.9060 73.1970 ;
        RECT 3.7720 72.1035 3.7980 73.1970 ;
        RECT 3.6640 72.1035 3.6900 73.1970 ;
        RECT 3.5560 72.1035 3.5820 73.1970 ;
        RECT 3.4480 72.1035 3.4740 73.1970 ;
        RECT 3.3400 72.1035 3.3660 73.1970 ;
        RECT 3.2320 72.1035 3.2580 73.1970 ;
        RECT 3.1240 72.1035 3.1500 73.1970 ;
        RECT 3.0160 72.1035 3.0420 73.1970 ;
        RECT 2.9080 72.1035 2.9340 73.1970 ;
        RECT 2.8000 72.1035 2.8260 73.1970 ;
        RECT 2.6920 72.1035 2.7180 73.1970 ;
        RECT 2.5840 72.1035 2.6100 73.1970 ;
        RECT 2.4760 72.1035 2.5020 73.1970 ;
        RECT 2.3680 72.1035 2.3940 73.1970 ;
        RECT 2.2600 72.1035 2.2860 73.1970 ;
        RECT 2.1520 72.1035 2.1780 73.1970 ;
        RECT 2.0440 72.1035 2.0700 73.1970 ;
        RECT 1.9360 72.1035 1.9620 73.1970 ;
        RECT 1.8280 72.1035 1.8540 73.1970 ;
        RECT 1.7200 72.1035 1.7460 73.1970 ;
        RECT 1.6120 72.1035 1.6380 73.1970 ;
        RECT 1.5040 72.1035 1.5300 73.1970 ;
        RECT 1.3960 72.1035 1.4220 73.1970 ;
        RECT 1.2880 72.1035 1.3140 73.1970 ;
        RECT 1.1800 72.1035 1.2060 73.1970 ;
        RECT 1.0720 72.1035 1.0980 73.1970 ;
        RECT 0.9640 72.1035 0.9900 73.1970 ;
        RECT 0.8560 72.1035 0.8820 73.1970 ;
        RECT 0.7480 72.1035 0.7740 73.1970 ;
        RECT 0.6400 72.1035 0.6660 73.1970 ;
        RECT 0.5320 72.1035 0.5580 73.1970 ;
        RECT 0.4240 72.1035 0.4500 73.1970 ;
        RECT 0.3160 72.1035 0.3420 73.1970 ;
        RECT 0.2080 72.1035 0.2340 73.1970 ;
        RECT 0.0050 72.1035 0.0900 73.1970 ;
        RECT 8.6410 73.1835 8.7690 74.2770 ;
        RECT 8.6270 73.8490 8.7690 74.1715 ;
        RECT 8.4790 73.5760 8.5410 74.2770 ;
        RECT 8.4650 73.8855 8.5410 74.0390 ;
        RECT 8.4790 73.1835 8.5050 74.2770 ;
        RECT 8.4790 73.3045 8.5190 73.5440 ;
        RECT 8.4790 73.1835 8.5410 73.2725 ;
        RECT 8.1820 73.6340 8.3880 74.2770 ;
        RECT 8.3620 73.1835 8.3880 74.2770 ;
        RECT 8.1820 73.9110 8.4020 74.1690 ;
        RECT 8.1820 73.1835 8.2800 74.2770 ;
        RECT 7.7650 73.1835 7.8480 74.2770 ;
        RECT 7.7650 73.2720 7.8620 74.2075 ;
        RECT 16.4440 73.1835 16.5290 74.2770 ;
        RECT 16.3000 73.1835 16.3260 74.2770 ;
        RECT 16.1920 73.1835 16.2180 74.2770 ;
        RECT 16.0840 73.1835 16.1100 74.2770 ;
        RECT 15.9760 73.1835 16.0020 74.2770 ;
        RECT 15.8680 73.1835 15.8940 74.2770 ;
        RECT 15.7600 73.1835 15.7860 74.2770 ;
        RECT 15.6520 73.1835 15.6780 74.2770 ;
        RECT 15.5440 73.1835 15.5700 74.2770 ;
        RECT 15.4360 73.1835 15.4620 74.2770 ;
        RECT 15.3280 73.1835 15.3540 74.2770 ;
        RECT 15.2200 73.1835 15.2460 74.2770 ;
        RECT 15.1120 73.1835 15.1380 74.2770 ;
        RECT 15.0040 73.1835 15.0300 74.2770 ;
        RECT 14.8960 73.1835 14.9220 74.2770 ;
        RECT 14.7880 73.1835 14.8140 74.2770 ;
        RECT 14.6800 73.1835 14.7060 74.2770 ;
        RECT 14.5720 73.1835 14.5980 74.2770 ;
        RECT 14.4640 73.1835 14.4900 74.2770 ;
        RECT 14.3560 73.1835 14.3820 74.2770 ;
        RECT 14.2480 73.1835 14.2740 74.2770 ;
        RECT 14.1400 73.1835 14.1660 74.2770 ;
        RECT 14.0320 73.1835 14.0580 74.2770 ;
        RECT 13.9240 73.1835 13.9500 74.2770 ;
        RECT 13.8160 73.1835 13.8420 74.2770 ;
        RECT 13.7080 73.1835 13.7340 74.2770 ;
        RECT 13.6000 73.1835 13.6260 74.2770 ;
        RECT 13.4920 73.1835 13.5180 74.2770 ;
        RECT 13.3840 73.1835 13.4100 74.2770 ;
        RECT 13.2760 73.1835 13.3020 74.2770 ;
        RECT 13.1680 73.1835 13.1940 74.2770 ;
        RECT 13.0600 73.1835 13.0860 74.2770 ;
        RECT 12.9520 73.1835 12.9780 74.2770 ;
        RECT 12.8440 73.1835 12.8700 74.2770 ;
        RECT 12.7360 73.1835 12.7620 74.2770 ;
        RECT 12.6280 73.1835 12.6540 74.2770 ;
        RECT 12.5200 73.1835 12.5460 74.2770 ;
        RECT 12.4120 73.1835 12.4380 74.2770 ;
        RECT 12.3040 73.1835 12.3300 74.2770 ;
        RECT 12.1960 73.1835 12.2220 74.2770 ;
        RECT 12.0880 73.1835 12.1140 74.2770 ;
        RECT 11.9800 73.1835 12.0060 74.2770 ;
        RECT 11.8720 73.1835 11.8980 74.2770 ;
        RECT 11.7640 73.1835 11.7900 74.2770 ;
        RECT 11.6560 73.1835 11.6820 74.2770 ;
        RECT 11.5480 73.1835 11.5740 74.2770 ;
        RECT 11.4400 73.1835 11.4660 74.2770 ;
        RECT 11.3320 73.1835 11.3580 74.2770 ;
        RECT 11.2240 73.1835 11.2500 74.2770 ;
        RECT 11.1160 73.1835 11.1420 74.2770 ;
        RECT 11.0080 73.1835 11.0340 74.2770 ;
        RECT 10.9000 73.1835 10.9260 74.2770 ;
        RECT 10.7920 73.1835 10.8180 74.2770 ;
        RECT 10.6840 73.1835 10.7100 74.2770 ;
        RECT 10.5760 73.1835 10.6020 74.2770 ;
        RECT 10.4680 73.1835 10.4940 74.2770 ;
        RECT 10.3600 73.1835 10.3860 74.2770 ;
        RECT 10.2520 73.1835 10.2780 74.2770 ;
        RECT 10.1440 73.1835 10.1700 74.2770 ;
        RECT 10.0360 73.1835 10.0620 74.2770 ;
        RECT 9.9280 73.1835 9.9540 74.2770 ;
        RECT 9.8200 73.1835 9.8460 74.2770 ;
        RECT 9.7120 73.1835 9.7380 74.2770 ;
        RECT 9.6040 73.1835 9.6300 74.2770 ;
        RECT 9.4960 73.1835 9.5220 74.2770 ;
        RECT 9.3880 73.1835 9.4140 74.2770 ;
        RECT 9.1750 73.1835 9.2520 74.2770 ;
        RECT 7.2820 73.1835 7.3590 74.2770 ;
        RECT 7.1200 73.1835 7.1460 74.2770 ;
        RECT 7.0120 73.1835 7.0380 74.2770 ;
        RECT 6.9040 73.1835 6.9300 74.2770 ;
        RECT 6.7960 73.1835 6.8220 74.2770 ;
        RECT 6.6880 73.1835 6.7140 74.2770 ;
        RECT 6.5800 73.1835 6.6060 74.2770 ;
        RECT 6.4720 73.1835 6.4980 74.2770 ;
        RECT 6.3640 73.1835 6.3900 74.2770 ;
        RECT 6.2560 73.1835 6.2820 74.2770 ;
        RECT 6.1480 73.1835 6.1740 74.2770 ;
        RECT 6.0400 73.1835 6.0660 74.2770 ;
        RECT 5.9320 73.1835 5.9580 74.2770 ;
        RECT 5.8240 73.1835 5.8500 74.2770 ;
        RECT 5.7160 73.1835 5.7420 74.2770 ;
        RECT 5.6080 73.1835 5.6340 74.2770 ;
        RECT 5.5000 73.1835 5.5260 74.2770 ;
        RECT 5.3920 73.1835 5.4180 74.2770 ;
        RECT 5.2840 73.1835 5.3100 74.2770 ;
        RECT 5.1760 73.1835 5.2020 74.2770 ;
        RECT 5.0680 73.1835 5.0940 74.2770 ;
        RECT 4.9600 73.1835 4.9860 74.2770 ;
        RECT 4.8520 73.1835 4.8780 74.2770 ;
        RECT 4.7440 73.1835 4.7700 74.2770 ;
        RECT 4.6360 73.1835 4.6620 74.2770 ;
        RECT 4.5280 73.1835 4.5540 74.2770 ;
        RECT 4.4200 73.1835 4.4460 74.2770 ;
        RECT 4.3120 73.1835 4.3380 74.2770 ;
        RECT 4.2040 73.1835 4.2300 74.2770 ;
        RECT 4.0960 73.1835 4.1220 74.2770 ;
        RECT 3.9880 73.1835 4.0140 74.2770 ;
        RECT 3.8800 73.1835 3.9060 74.2770 ;
        RECT 3.7720 73.1835 3.7980 74.2770 ;
        RECT 3.6640 73.1835 3.6900 74.2770 ;
        RECT 3.5560 73.1835 3.5820 74.2770 ;
        RECT 3.4480 73.1835 3.4740 74.2770 ;
        RECT 3.3400 73.1835 3.3660 74.2770 ;
        RECT 3.2320 73.1835 3.2580 74.2770 ;
        RECT 3.1240 73.1835 3.1500 74.2770 ;
        RECT 3.0160 73.1835 3.0420 74.2770 ;
        RECT 2.9080 73.1835 2.9340 74.2770 ;
        RECT 2.8000 73.1835 2.8260 74.2770 ;
        RECT 2.6920 73.1835 2.7180 74.2770 ;
        RECT 2.5840 73.1835 2.6100 74.2770 ;
        RECT 2.4760 73.1835 2.5020 74.2770 ;
        RECT 2.3680 73.1835 2.3940 74.2770 ;
        RECT 2.2600 73.1835 2.2860 74.2770 ;
        RECT 2.1520 73.1835 2.1780 74.2770 ;
        RECT 2.0440 73.1835 2.0700 74.2770 ;
        RECT 1.9360 73.1835 1.9620 74.2770 ;
        RECT 1.8280 73.1835 1.8540 74.2770 ;
        RECT 1.7200 73.1835 1.7460 74.2770 ;
        RECT 1.6120 73.1835 1.6380 74.2770 ;
        RECT 1.5040 73.1835 1.5300 74.2770 ;
        RECT 1.3960 73.1835 1.4220 74.2770 ;
        RECT 1.2880 73.1835 1.3140 74.2770 ;
        RECT 1.1800 73.1835 1.2060 74.2770 ;
        RECT 1.0720 73.1835 1.0980 74.2770 ;
        RECT 0.9640 73.1835 0.9900 74.2770 ;
        RECT 0.8560 73.1835 0.8820 74.2770 ;
        RECT 0.7480 73.1835 0.7740 74.2770 ;
        RECT 0.6400 73.1835 0.6660 74.2770 ;
        RECT 0.5320 73.1835 0.5580 74.2770 ;
        RECT 0.4240 73.1835 0.4500 74.2770 ;
        RECT 0.3160 73.1835 0.3420 74.2770 ;
        RECT 0.2080 73.1835 0.2340 74.2770 ;
        RECT 0.0050 73.1835 0.0900 74.2770 ;
        RECT 8.6410 74.2635 8.7690 75.3570 ;
        RECT 8.6270 74.9290 8.7690 75.2515 ;
        RECT 8.4790 74.6560 8.5410 75.3570 ;
        RECT 8.4650 74.9655 8.5410 75.1190 ;
        RECT 8.4790 74.2635 8.5050 75.3570 ;
        RECT 8.4790 74.3845 8.5190 74.6240 ;
        RECT 8.4790 74.2635 8.5410 74.3525 ;
        RECT 8.1820 74.7140 8.3880 75.3570 ;
        RECT 8.3620 74.2635 8.3880 75.3570 ;
        RECT 8.1820 74.9910 8.4020 75.2490 ;
        RECT 8.1820 74.2635 8.2800 75.3570 ;
        RECT 7.7650 74.2635 7.8480 75.3570 ;
        RECT 7.7650 74.3520 7.8620 75.2875 ;
        RECT 16.4440 74.2635 16.5290 75.3570 ;
        RECT 16.3000 74.2635 16.3260 75.3570 ;
        RECT 16.1920 74.2635 16.2180 75.3570 ;
        RECT 16.0840 74.2635 16.1100 75.3570 ;
        RECT 15.9760 74.2635 16.0020 75.3570 ;
        RECT 15.8680 74.2635 15.8940 75.3570 ;
        RECT 15.7600 74.2635 15.7860 75.3570 ;
        RECT 15.6520 74.2635 15.6780 75.3570 ;
        RECT 15.5440 74.2635 15.5700 75.3570 ;
        RECT 15.4360 74.2635 15.4620 75.3570 ;
        RECT 15.3280 74.2635 15.3540 75.3570 ;
        RECT 15.2200 74.2635 15.2460 75.3570 ;
        RECT 15.1120 74.2635 15.1380 75.3570 ;
        RECT 15.0040 74.2635 15.0300 75.3570 ;
        RECT 14.8960 74.2635 14.9220 75.3570 ;
        RECT 14.7880 74.2635 14.8140 75.3570 ;
        RECT 14.6800 74.2635 14.7060 75.3570 ;
        RECT 14.5720 74.2635 14.5980 75.3570 ;
        RECT 14.4640 74.2635 14.4900 75.3570 ;
        RECT 14.3560 74.2635 14.3820 75.3570 ;
        RECT 14.2480 74.2635 14.2740 75.3570 ;
        RECT 14.1400 74.2635 14.1660 75.3570 ;
        RECT 14.0320 74.2635 14.0580 75.3570 ;
        RECT 13.9240 74.2635 13.9500 75.3570 ;
        RECT 13.8160 74.2635 13.8420 75.3570 ;
        RECT 13.7080 74.2635 13.7340 75.3570 ;
        RECT 13.6000 74.2635 13.6260 75.3570 ;
        RECT 13.4920 74.2635 13.5180 75.3570 ;
        RECT 13.3840 74.2635 13.4100 75.3570 ;
        RECT 13.2760 74.2635 13.3020 75.3570 ;
        RECT 13.1680 74.2635 13.1940 75.3570 ;
        RECT 13.0600 74.2635 13.0860 75.3570 ;
        RECT 12.9520 74.2635 12.9780 75.3570 ;
        RECT 12.8440 74.2635 12.8700 75.3570 ;
        RECT 12.7360 74.2635 12.7620 75.3570 ;
        RECT 12.6280 74.2635 12.6540 75.3570 ;
        RECT 12.5200 74.2635 12.5460 75.3570 ;
        RECT 12.4120 74.2635 12.4380 75.3570 ;
        RECT 12.3040 74.2635 12.3300 75.3570 ;
        RECT 12.1960 74.2635 12.2220 75.3570 ;
        RECT 12.0880 74.2635 12.1140 75.3570 ;
        RECT 11.9800 74.2635 12.0060 75.3570 ;
        RECT 11.8720 74.2635 11.8980 75.3570 ;
        RECT 11.7640 74.2635 11.7900 75.3570 ;
        RECT 11.6560 74.2635 11.6820 75.3570 ;
        RECT 11.5480 74.2635 11.5740 75.3570 ;
        RECT 11.4400 74.2635 11.4660 75.3570 ;
        RECT 11.3320 74.2635 11.3580 75.3570 ;
        RECT 11.2240 74.2635 11.2500 75.3570 ;
        RECT 11.1160 74.2635 11.1420 75.3570 ;
        RECT 11.0080 74.2635 11.0340 75.3570 ;
        RECT 10.9000 74.2635 10.9260 75.3570 ;
        RECT 10.7920 74.2635 10.8180 75.3570 ;
        RECT 10.6840 74.2635 10.7100 75.3570 ;
        RECT 10.5760 74.2635 10.6020 75.3570 ;
        RECT 10.4680 74.2635 10.4940 75.3570 ;
        RECT 10.3600 74.2635 10.3860 75.3570 ;
        RECT 10.2520 74.2635 10.2780 75.3570 ;
        RECT 10.1440 74.2635 10.1700 75.3570 ;
        RECT 10.0360 74.2635 10.0620 75.3570 ;
        RECT 9.9280 74.2635 9.9540 75.3570 ;
        RECT 9.8200 74.2635 9.8460 75.3570 ;
        RECT 9.7120 74.2635 9.7380 75.3570 ;
        RECT 9.6040 74.2635 9.6300 75.3570 ;
        RECT 9.4960 74.2635 9.5220 75.3570 ;
        RECT 9.3880 74.2635 9.4140 75.3570 ;
        RECT 9.1750 74.2635 9.2520 75.3570 ;
        RECT 7.2820 74.2635 7.3590 75.3570 ;
        RECT 7.1200 74.2635 7.1460 75.3570 ;
        RECT 7.0120 74.2635 7.0380 75.3570 ;
        RECT 6.9040 74.2635 6.9300 75.3570 ;
        RECT 6.7960 74.2635 6.8220 75.3570 ;
        RECT 6.6880 74.2635 6.7140 75.3570 ;
        RECT 6.5800 74.2635 6.6060 75.3570 ;
        RECT 6.4720 74.2635 6.4980 75.3570 ;
        RECT 6.3640 74.2635 6.3900 75.3570 ;
        RECT 6.2560 74.2635 6.2820 75.3570 ;
        RECT 6.1480 74.2635 6.1740 75.3570 ;
        RECT 6.0400 74.2635 6.0660 75.3570 ;
        RECT 5.9320 74.2635 5.9580 75.3570 ;
        RECT 5.8240 74.2635 5.8500 75.3570 ;
        RECT 5.7160 74.2635 5.7420 75.3570 ;
        RECT 5.6080 74.2635 5.6340 75.3570 ;
        RECT 5.5000 74.2635 5.5260 75.3570 ;
        RECT 5.3920 74.2635 5.4180 75.3570 ;
        RECT 5.2840 74.2635 5.3100 75.3570 ;
        RECT 5.1760 74.2635 5.2020 75.3570 ;
        RECT 5.0680 74.2635 5.0940 75.3570 ;
        RECT 4.9600 74.2635 4.9860 75.3570 ;
        RECT 4.8520 74.2635 4.8780 75.3570 ;
        RECT 4.7440 74.2635 4.7700 75.3570 ;
        RECT 4.6360 74.2635 4.6620 75.3570 ;
        RECT 4.5280 74.2635 4.5540 75.3570 ;
        RECT 4.4200 74.2635 4.4460 75.3570 ;
        RECT 4.3120 74.2635 4.3380 75.3570 ;
        RECT 4.2040 74.2635 4.2300 75.3570 ;
        RECT 4.0960 74.2635 4.1220 75.3570 ;
        RECT 3.9880 74.2635 4.0140 75.3570 ;
        RECT 3.8800 74.2635 3.9060 75.3570 ;
        RECT 3.7720 74.2635 3.7980 75.3570 ;
        RECT 3.6640 74.2635 3.6900 75.3570 ;
        RECT 3.5560 74.2635 3.5820 75.3570 ;
        RECT 3.4480 74.2635 3.4740 75.3570 ;
        RECT 3.3400 74.2635 3.3660 75.3570 ;
        RECT 3.2320 74.2635 3.2580 75.3570 ;
        RECT 3.1240 74.2635 3.1500 75.3570 ;
        RECT 3.0160 74.2635 3.0420 75.3570 ;
        RECT 2.9080 74.2635 2.9340 75.3570 ;
        RECT 2.8000 74.2635 2.8260 75.3570 ;
        RECT 2.6920 74.2635 2.7180 75.3570 ;
        RECT 2.5840 74.2635 2.6100 75.3570 ;
        RECT 2.4760 74.2635 2.5020 75.3570 ;
        RECT 2.3680 74.2635 2.3940 75.3570 ;
        RECT 2.2600 74.2635 2.2860 75.3570 ;
        RECT 2.1520 74.2635 2.1780 75.3570 ;
        RECT 2.0440 74.2635 2.0700 75.3570 ;
        RECT 1.9360 74.2635 1.9620 75.3570 ;
        RECT 1.8280 74.2635 1.8540 75.3570 ;
        RECT 1.7200 74.2635 1.7460 75.3570 ;
        RECT 1.6120 74.2635 1.6380 75.3570 ;
        RECT 1.5040 74.2635 1.5300 75.3570 ;
        RECT 1.3960 74.2635 1.4220 75.3570 ;
        RECT 1.2880 74.2635 1.3140 75.3570 ;
        RECT 1.1800 74.2635 1.2060 75.3570 ;
        RECT 1.0720 74.2635 1.0980 75.3570 ;
        RECT 0.9640 74.2635 0.9900 75.3570 ;
        RECT 0.8560 74.2635 0.8820 75.3570 ;
        RECT 0.7480 74.2635 0.7740 75.3570 ;
        RECT 0.6400 74.2635 0.6660 75.3570 ;
        RECT 0.5320 74.2635 0.5580 75.3570 ;
        RECT 0.4240 74.2635 0.4500 75.3570 ;
        RECT 0.3160 74.2635 0.3420 75.3570 ;
        RECT 0.2080 74.2635 0.2340 75.3570 ;
        RECT 0.0050 74.2635 0.0900 75.3570 ;
        RECT 8.6410 75.3435 8.7690 76.4370 ;
        RECT 8.6270 76.0090 8.7690 76.3315 ;
        RECT 8.4790 75.7360 8.5410 76.4370 ;
        RECT 8.4650 76.0455 8.5410 76.1990 ;
        RECT 8.4790 75.3435 8.5050 76.4370 ;
        RECT 8.4790 75.4645 8.5190 75.7040 ;
        RECT 8.4790 75.3435 8.5410 75.4325 ;
        RECT 8.1820 75.7940 8.3880 76.4370 ;
        RECT 8.3620 75.3435 8.3880 76.4370 ;
        RECT 8.1820 76.0710 8.4020 76.3290 ;
        RECT 8.1820 75.3435 8.2800 76.4370 ;
        RECT 7.7650 75.3435 7.8480 76.4370 ;
        RECT 7.7650 75.4320 7.8620 76.3675 ;
        RECT 16.4440 75.3435 16.5290 76.4370 ;
        RECT 16.3000 75.3435 16.3260 76.4370 ;
        RECT 16.1920 75.3435 16.2180 76.4370 ;
        RECT 16.0840 75.3435 16.1100 76.4370 ;
        RECT 15.9760 75.3435 16.0020 76.4370 ;
        RECT 15.8680 75.3435 15.8940 76.4370 ;
        RECT 15.7600 75.3435 15.7860 76.4370 ;
        RECT 15.6520 75.3435 15.6780 76.4370 ;
        RECT 15.5440 75.3435 15.5700 76.4370 ;
        RECT 15.4360 75.3435 15.4620 76.4370 ;
        RECT 15.3280 75.3435 15.3540 76.4370 ;
        RECT 15.2200 75.3435 15.2460 76.4370 ;
        RECT 15.1120 75.3435 15.1380 76.4370 ;
        RECT 15.0040 75.3435 15.0300 76.4370 ;
        RECT 14.8960 75.3435 14.9220 76.4370 ;
        RECT 14.7880 75.3435 14.8140 76.4370 ;
        RECT 14.6800 75.3435 14.7060 76.4370 ;
        RECT 14.5720 75.3435 14.5980 76.4370 ;
        RECT 14.4640 75.3435 14.4900 76.4370 ;
        RECT 14.3560 75.3435 14.3820 76.4370 ;
        RECT 14.2480 75.3435 14.2740 76.4370 ;
        RECT 14.1400 75.3435 14.1660 76.4370 ;
        RECT 14.0320 75.3435 14.0580 76.4370 ;
        RECT 13.9240 75.3435 13.9500 76.4370 ;
        RECT 13.8160 75.3435 13.8420 76.4370 ;
        RECT 13.7080 75.3435 13.7340 76.4370 ;
        RECT 13.6000 75.3435 13.6260 76.4370 ;
        RECT 13.4920 75.3435 13.5180 76.4370 ;
        RECT 13.3840 75.3435 13.4100 76.4370 ;
        RECT 13.2760 75.3435 13.3020 76.4370 ;
        RECT 13.1680 75.3435 13.1940 76.4370 ;
        RECT 13.0600 75.3435 13.0860 76.4370 ;
        RECT 12.9520 75.3435 12.9780 76.4370 ;
        RECT 12.8440 75.3435 12.8700 76.4370 ;
        RECT 12.7360 75.3435 12.7620 76.4370 ;
        RECT 12.6280 75.3435 12.6540 76.4370 ;
        RECT 12.5200 75.3435 12.5460 76.4370 ;
        RECT 12.4120 75.3435 12.4380 76.4370 ;
        RECT 12.3040 75.3435 12.3300 76.4370 ;
        RECT 12.1960 75.3435 12.2220 76.4370 ;
        RECT 12.0880 75.3435 12.1140 76.4370 ;
        RECT 11.9800 75.3435 12.0060 76.4370 ;
        RECT 11.8720 75.3435 11.8980 76.4370 ;
        RECT 11.7640 75.3435 11.7900 76.4370 ;
        RECT 11.6560 75.3435 11.6820 76.4370 ;
        RECT 11.5480 75.3435 11.5740 76.4370 ;
        RECT 11.4400 75.3435 11.4660 76.4370 ;
        RECT 11.3320 75.3435 11.3580 76.4370 ;
        RECT 11.2240 75.3435 11.2500 76.4370 ;
        RECT 11.1160 75.3435 11.1420 76.4370 ;
        RECT 11.0080 75.3435 11.0340 76.4370 ;
        RECT 10.9000 75.3435 10.9260 76.4370 ;
        RECT 10.7920 75.3435 10.8180 76.4370 ;
        RECT 10.6840 75.3435 10.7100 76.4370 ;
        RECT 10.5760 75.3435 10.6020 76.4370 ;
        RECT 10.4680 75.3435 10.4940 76.4370 ;
        RECT 10.3600 75.3435 10.3860 76.4370 ;
        RECT 10.2520 75.3435 10.2780 76.4370 ;
        RECT 10.1440 75.3435 10.1700 76.4370 ;
        RECT 10.0360 75.3435 10.0620 76.4370 ;
        RECT 9.9280 75.3435 9.9540 76.4370 ;
        RECT 9.8200 75.3435 9.8460 76.4370 ;
        RECT 9.7120 75.3435 9.7380 76.4370 ;
        RECT 9.6040 75.3435 9.6300 76.4370 ;
        RECT 9.4960 75.3435 9.5220 76.4370 ;
        RECT 9.3880 75.3435 9.4140 76.4370 ;
        RECT 9.1750 75.3435 9.2520 76.4370 ;
        RECT 7.2820 75.3435 7.3590 76.4370 ;
        RECT 7.1200 75.3435 7.1460 76.4370 ;
        RECT 7.0120 75.3435 7.0380 76.4370 ;
        RECT 6.9040 75.3435 6.9300 76.4370 ;
        RECT 6.7960 75.3435 6.8220 76.4370 ;
        RECT 6.6880 75.3435 6.7140 76.4370 ;
        RECT 6.5800 75.3435 6.6060 76.4370 ;
        RECT 6.4720 75.3435 6.4980 76.4370 ;
        RECT 6.3640 75.3435 6.3900 76.4370 ;
        RECT 6.2560 75.3435 6.2820 76.4370 ;
        RECT 6.1480 75.3435 6.1740 76.4370 ;
        RECT 6.0400 75.3435 6.0660 76.4370 ;
        RECT 5.9320 75.3435 5.9580 76.4370 ;
        RECT 5.8240 75.3435 5.8500 76.4370 ;
        RECT 5.7160 75.3435 5.7420 76.4370 ;
        RECT 5.6080 75.3435 5.6340 76.4370 ;
        RECT 5.5000 75.3435 5.5260 76.4370 ;
        RECT 5.3920 75.3435 5.4180 76.4370 ;
        RECT 5.2840 75.3435 5.3100 76.4370 ;
        RECT 5.1760 75.3435 5.2020 76.4370 ;
        RECT 5.0680 75.3435 5.0940 76.4370 ;
        RECT 4.9600 75.3435 4.9860 76.4370 ;
        RECT 4.8520 75.3435 4.8780 76.4370 ;
        RECT 4.7440 75.3435 4.7700 76.4370 ;
        RECT 4.6360 75.3435 4.6620 76.4370 ;
        RECT 4.5280 75.3435 4.5540 76.4370 ;
        RECT 4.4200 75.3435 4.4460 76.4370 ;
        RECT 4.3120 75.3435 4.3380 76.4370 ;
        RECT 4.2040 75.3435 4.2300 76.4370 ;
        RECT 4.0960 75.3435 4.1220 76.4370 ;
        RECT 3.9880 75.3435 4.0140 76.4370 ;
        RECT 3.8800 75.3435 3.9060 76.4370 ;
        RECT 3.7720 75.3435 3.7980 76.4370 ;
        RECT 3.6640 75.3435 3.6900 76.4370 ;
        RECT 3.5560 75.3435 3.5820 76.4370 ;
        RECT 3.4480 75.3435 3.4740 76.4370 ;
        RECT 3.3400 75.3435 3.3660 76.4370 ;
        RECT 3.2320 75.3435 3.2580 76.4370 ;
        RECT 3.1240 75.3435 3.1500 76.4370 ;
        RECT 3.0160 75.3435 3.0420 76.4370 ;
        RECT 2.9080 75.3435 2.9340 76.4370 ;
        RECT 2.8000 75.3435 2.8260 76.4370 ;
        RECT 2.6920 75.3435 2.7180 76.4370 ;
        RECT 2.5840 75.3435 2.6100 76.4370 ;
        RECT 2.4760 75.3435 2.5020 76.4370 ;
        RECT 2.3680 75.3435 2.3940 76.4370 ;
        RECT 2.2600 75.3435 2.2860 76.4370 ;
        RECT 2.1520 75.3435 2.1780 76.4370 ;
        RECT 2.0440 75.3435 2.0700 76.4370 ;
        RECT 1.9360 75.3435 1.9620 76.4370 ;
        RECT 1.8280 75.3435 1.8540 76.4370 ;
        RECT 1.7200 75.3435 1.7460 76.4370 ;
        RECT 1.6120 75.3435 1.6380 76.4370 ;
        RECT 1.5040 75.3435 1.5300 76.4370 ;
        RECT 1.3960 75.3435 1.4220 76.4370 ;
        RECT 1.2880 75.3435 1.3140 76.4370 ;
        RECT 1.1800 75.3435 1.2060 76.4370 ;
        RECT 1.0720 75.3435 1.0980 76.4370 ;
        RECT 0.9640 75.3435 0.9900 76.4370 ;
        RECT 0.8560 75.3435 0.8820 76.4370 ;
        RECT 0.7480 75.3435 0.7740 76.4370 ;
        RECT 0.6400 75.3435 0.6660 76.4370 ;
        RECT 0.5320 75.3435 0.5580 76.4370 ;
        RECT 0.4240 75.3435 0.4500 76.4370 ;
        RECT 0.3160 75.3435 0.3420 76.4370 ;
        RECT 0.2080 75.3435 0.2340 76.4370 ;
        RECT 0.0050 75.3435 0.0900 76.4370 ;
        RECT 8.6410 76.4235 8.7690 77.5170 ;
        RECT 8.6270 77.0890 8.7690 77.4115 ;
        RECT 8.4790 76.8160 8.5410 77.5170 ;
        RECT 8.4650 77.1255 8.5410 77.2790 ;
        RECT 8.4790 76.4235 8.5050 77.5170 ;
        RECT 8.4790 76.5445 8.5190 76.7840 ;
        RECT 8.4790 76.4235 8.5410 76.5125 ;
        RECT 8.1820 76.8740 8.3880 77.5170 ;
        RECT 8.3620 76.4235 8.3880 77.5170 ;
        RECT 8.1820 77.1510 8.4020 77.4090 ;
        RECT 8.1820 76.4235 8.2800 77.5170 ;
        RECT 7.7650 76.4235 7.8480 77.5170 ;
        RECT 7.7650 76.5120 7.8620 77.4475 ;
        RECT 16.4440 76.4235 16.5290 77.5170 ;
        RECT 16.3000 76.4235 16.3260 77.5170 ;
        RECT 16.1920 76.4235 16.2180 77.5170 ;
        RECT 16.0840 76.4235 16.1100 77.5170 ;
        RECT 15.9760 76.4235 16.0020 77.5170 ;
        RECT 15.8680 76.4235 15.8940 77.5170 ;
        RECT 15.7600 76.4235 15.7860 77.5170 ;
        RECT 15.6520 76.4235 15.6780 77.5170 ;
        RECT 15.5440 76.4235 15.5700 77.5170 ;
        RECT 15.4360 76.4235 15.4620 77.5170 ;
        RECT 15.3280 76.4235 15.3540 77.5170 ;
        RECT 15.2200 76.4235 15.2460 77.5170 ;
        RECT 15.1120 76.4235 15.1380 77.5170 ;
        RECT 15.0040 76.4235 15.0300 77.5170 ;
        RECT 14.8960 76.4235 14.9220 77.5170 ;
        RECT 14.7880 76.4235 14.8140 77.5170 ;
        RECT 14.6800 76.4235 14.7060 77.5170 ;
        RECT 14.5720 76.4235 14.5980 77.5170 ;
        RECT 14.4640 76.4235 14.4900 77.5170 ;
        RECT 14.3560 76.4235 14.3820 77.5170 ;
        RECT 14.2480 76.4235 14.2740 77.5170 ;
        RECT 14.1400 76.4235 14.1660 77.5170 ;
        RECT 14.0320 76.4235 14.0580 77.5170 ;
        RECT 13.9240 76.4235 13.9500 77.5170 ;
        RECT 13.8160 76.4235 13.8420 77.5170 ;
        RECT 13.7080 76.4235 13.7340 77.5170 ;
        RECT 13.6000 76.4235 13.6260 77.5170 ;
        RECT 13.4920 76.4235 13.5180 77.5170 ;
        RECT 13.3840 76.4235 13.4100 77.5170 ;
        RECT 13.2760 76.4235 13.3020 77.5170 ;
        RECT 13.1680 76.4235 13.1940 77.5170 ;
        RECT 13.0600 76.4235 13.0860 77.5170 ;
        RECT 12.9520 76.4235 12.9780 77.5170 ;
        RECT 12.8440 76.4235 12.8700 77.5170 ;
        RECT 12.7360 76.4235 12.7620 77.5170 ;
        RECT 12.6280 76.4235 12.6540 77.5170 ;
        RECT 12.5200 76.4235 12.5460 77.5170 ;
        RECT 12.4120 76.4235 12.4380 77.5170 ;
        RECT 12.3040 76.4235 12.3300 77.5170 ;
        RECT 12.1960 76.4235 12.2220 77.5170 ;
        RECT 12.0880 76.4235 12.1140 77.5170 ;
        RECT 11.9800 76.4235 12.0060 77.5170 ;
        RECT 11.8720 76.4235 11.8980 77.5170 ;
        RECT 11.7640 76.4235 11.7900 77.5170 ;
        RECT 11.6560 76.4235 11.6820 77.5170 ;
        RECT 11.5480 76.4235 11.5740 77.5170 ;
        RECT 11.4400 76.4235 11.4660 77.5170 ;
        RECT 11.3320 76.4235 11.3580 77.5170 ;
        RECT 11.2240 76.4235 11.2500 77.5170 ;
        RECT 11.1160 76.4235 11.1420 77.5170 ;
        RECT 11.0080 76.4235 11.0340 77.5170 ;
        RECT 10.9000 76.4235 10.9260 77.5170 ;
        RECT 10.7920 76.4235 10.8180 77.5170 ;
        RECT 10.6840 76.4235 10.7100 77.5170 ;
        RECT 10.5760 76.4235 10.6020 77.5170 ;
        RECT 10.4680 76.4235 10.4940 77.5170 ;
        RECT 10.3600 76.4235 10.3860 77.5170 ;
        RECT 10.2520 76.4235 10.2780 77.5170 ;
        RECT 10.1440 76.4235 10.1700 77.5170 ;
        RECT 10.0360 76.4235 10.0620 77.5170 ;
        RECT 9.9280 76.4235 9.9540 77.5170 ;
        RECT 9.8200 76.4235 9.8460 77.5170 ;
        RECT 9.7120 76.4235 9.7380 77.5170 ;
        RECT 9.6040 76.4235 9.6300 77.5170 ;
        RECT 9.4960 76.4235 9.5220 77.5170 ;
        RECT 9.3880 76.4235 9.4140 77.5170 ;
        RECT 9.1750 76.4235 9.2520 77.5170 ;
        RECT 7.2820 76.4235 7.3590 77.5170 ;
        RECT 7.1200 76.4235 7.1460 77.5170 ;
        RECT 7.0120 76.4235 7.0380 77.5170 ;
        RECT 6.9040 76.4235 6.9300 77.5170 ;
        RECT 6.7960 76.4235 6.8220 77.5170 ;
        RECT 6.6880 76.4235 6.7140 77.5170 ;
        RECT 6.5800 76.4235 6.6060 77.5170 ;
        RECT 6.4720 76.4235 6.4980 77.5170 ;
        RECT 6.3640 76.4235 6.3900 77.5170 ;
        RECT 6.2560 76.4235 6.2820 77.5170 ;
        RECT 6.1480 76.4235 6.1740 77.5170 ;
        RECT 6.0400 76.4235 6.0660 77.5170 ;
        RECT 5.9320 76.4235 5.9580 77.5170 ;
        RECT 5.8240 76.4235 5.8500 77.5170 ;
        RECT 5.7160 76.4235 5.7420 77.5170 ;
        RECT 5.6080 76.4235 5.6340 77.5170 ;
        RECT 5.5000 76.4235 5.5260 77.5170 ;
        RECT 5.3920 76.4235 5.4180 77.5170 ;
        RECT 5.2840 76.4235 5.3100 77.5170 ;
        RECT 5.1760 76.4235 5.2020 77.5170 ;
        RECT 5.0680 76.4235 5.0940 77.5170 ;
        RECT 4.9600 76.4235 4.9860 77.5170 ;
        RECT 4.8520 76.4235 4.8780 77.5170 ;
        RECT 4.7440 76.4235 4.7700 77.5170 ;
        RECT 4.6360 76.4235 4.6620 77.5170 ;
        RECT 4.5280 76.4235 4.5540 77.5170 ;
        RECT 4.4200 76.4235 4.4460 77.5170 ;
        RECT 4.3120 76.4235 4.3380 77.5170 ;
        RECT 4.2040 76.4235 4.2300 77.5170 ;
        RECT 4.0960 76.4235 4.1220 77.5170 ;
        RECT 3.9880 76.4235 4.0140 77.5170 ;
        RECT 3.8800 76.4235 3.9060 77.5170 ;
        RECT 3.7720 76.4235 3.7980 77.5170 ;
        RECT 3.6640 76.4235 3.6900 77.5170 ;
        RECT 3.5560 76.4235 3.5820 77.5170 ;
        RECT 3.4480 76.4235 3.4740 77.5170 ;
        RECT 3.3400 76.4235 3.3660 77.5170 ;
        RECT 3.2320 76.4235 3.2580 77.5170 ;
        RECT 3.1240 76.4235 3.1500 77.5170 ;
        RECT 3.0160 76.4235 3.0420 77.5170 ;
        RECT 2.9080 76.4235 2.9340 77.5170 ;
        RECT 2.8000 76.4235 2.8260 77.5170 ;
        RECT 2.6920 76.4235 2.7180 77.5170 ;
        RECT 2.5840 76.4235 2.6100 77.5170 ;
        RECT 2.4760 76.4235 2.5020 77.5170 ;
        RECT 2.3680 76.4235 2.3940 77.5170 ;
        RECT 2.2600 76.4235 2.2860 77.5170 ;
        RECT 2.1520 76.4235 2.1780 77.5170 ;
        RECT 2.0440 76.4235 2.0700 77.5170 ;
        RECT 1.9360 76.4235 1.9620 77.5170 ;
        RECT 1.8280 76.4235 1.8540 77.5170 ;
        RECT 1.7200 76.4235 1.7460 77.5170 ;
        RECT 1.6120 76.4235 1.6380 77.5170 ;
        RECT 1.5040 76.4235 1.5300 77.5170 ;
        RECT 1.3960 76.4235 1.4220 77.5170 ;
        RECT 1.2880 76.4235 1.3140 77.5170 ;
        RECT 1.1800 76.4235 1.2060 77.5170 ;
        RECT 1.0720 76.4235 1.0980 77.5170 ;
        RECT 0.9640 76.4235 0.9900 77.5170 ;
        RECT 0.8560 76.4235 0.8820 77.5170 ;
        RECT 0.7480 76.4235 0.7740 77.5170 ;
        RECT 0.6400 76.4235 0.6660 77.5170 ;
        RECT 0.5320 76.4235 0.5580 77.5170 ;
        RECT 0.4240 76.4235 0.4500 77.5170 ;
        RECT 0.3160 76.4235 0.3420 77.5170 ;
        RECT 0.2080 76.4235 0.2340 77.5170 ;
        RECT 0.0050 76.4235 0.0900 77.5170 ;
        RECT 8.6410 77.5035 8.7690 78.5970 ;
        RECT 8.6270 78.1690 8.7690 78.4915 ;
        RECT 8.4790 77.8960 8.5410 78.5970 ;
        RECT 8.4650 78.2055 8.5410 78.3590 ;
        RECT 8.4790 77.5035 8.5050 78.5970 ;
        RECT 8.4790 77.6245 8.5190 77.8640 ;
        RECT 8.4790 77.5035 8.5410 77.5925 ;
        RECT 8.1820 77.9540 8.3880 78.5970 ;
        RECT 8.3620 77.5035 8.3880 78.5970 ;
        RECT 8.1820 78.2310 8.4020 78.4890 ;
        RECT 8.1820 77.5035 8.2800 78.5970 ;
        RECT 7.7650 77.5035 7.8480 78.5970 ;
        RECT 7.7650 77.5920 7.8620 78.5275 ;
        RECT 16.4440 77.5035 16.5290 78.5970 ;
        RECT 16.3000 77.5035 16.3260 78.5970 ;
        RECT 16.1920 77.5035 16.2180 78.5970 ;
        RECT 16.0840 77.5035 16.1100 78.5970 ;
        RECT 15.9760 77.5035 16.0020 78.5970 ;
        RECT 15.8680 77.5035 15.8940 78.5970 ;
        RECT 15.7600 77.5035 15.7860 78.5970 ;
        RECT 15.6520 77.5035 15.6780 78.5970 ;
        RECT 15.5440 77.5035 15.5700 78.5970 ;
        RECT 15.4360 77.5035 15.4620 78.5970 ;
        RECT 15.3280 77.5035 15.3540 78.5970 ;
        RECT 15.2200 77.5035 15.2460 78.5970 ;
        RECT 15.1120 77.5035 15.1380 78.5970 ;
        RECT 15.0040 77.5035 15.0300 78.5970 ;
        RECT 14.8960 77.5035 14.9220 78.5970 ;
        RECT 14.7880 77.5035 14.8140 78.5970 ;
        RECT 14.6800 77.5035 14.7060 78.5970 ;
        RECT 14.5720 77.5035 14.5980 78.5970 ;
        RECT 14.4640 77.5035 14.4900 78.5970 ;
        RECT 14.3560 77.5035 14.3820 78.5970 ;
        RECT 14.2480 77.5035 14.2740 78.5970 ;
        RECT 14.1400 77.5035 14.1660 78.5970 ;
        RECT 14.0320 77.5035 14.0580 78.5970 ;
        RECT 13.9240 77.5035 13.9500 78.5970 ;
        RECT 13.8160 77.5035 13.8420 78.5970 ;
        RECT 13.7080 77.5035 13.7340 78.5970 ;
        RECT 13.6000 77.5035 13.6260 78.5970 ;
        RECT 13.4920 77.5035 13.5180 78.5970 ;
        RECT 13.3840 77.5035 13.4100 78.5970 ;
        RECT 13.2760 77.5035 13.3020 78.5970 ;
        RECT 13.1680 77.5035 13.1940 78.5970 ;
        RECT 13.0600 77.5035 13.0860 78.5970 ;
        RECT 12.9520 77.5035 12.9780 78.5970 ;
        RECT 12.8440 77.5035 12.8700 78.5970 ;
        RECT 12.7360 77.5035 12.7620 78.5970 ;
        RECT 12.6280 77.5035 12.6540 78.5970 ;
        RECT 12.5200 77.5035 12.5460 78.5970 ;
        RECT 12.4120 77.5035 12.4380 78.5970 ;
        RECT 12.3040 77.5035 12.3300 78.5970 ;
        RECT 12.1960 77.5035 12.2220 78.5970 ;
        RECT 12.0880 77.5035 12.1140 78.5970 ;
        RECT 11.9800 77.5035 12.0060 78.5970 ;
        RECT 11.8720 77.5035 11.8980 78.5970 ;
        RECT 11.7640 77.5035 11.7900 78.5970 ;
        RECT 11.6560 77.5035 11.6820 78.5970 ;
        RECT 11.5480 77.5035 11.5740 78.5970 ;
        RECT 11.4400 77.5035 11.4660 78.5970 ;
        RECT 11.3320 77.5035 11.3580 78.5970 ;
        RECT 11.2240 77.5035 11.2500 78.5970 ;
        RECT 11.1160 77.5035 11.1420 78.5970 ;
        RECT 11.0080 77.5035 11.0340 78.5970 ;
        RECT 10.9000 77.5035 10.9260 78.5970 ;
        RECT 10.7920 77.5035 10.8180 78.5970 ;
        RECT 10.6840 77.5035 10.7100 78.5970 ;
        RECT 10.5760 77.5035 10.6020 78.5970 ;
        RECT 10.4680 77.5035 10.4940 78.5970 ;
        RECT 10.3600 77.5035 10.3860 78.5970 ;
        RECT 10.2520 77.5035 10.2780 78.5970 ;
        RECT 10.1440 77.5035 10.1700 78.5970 ;
        RECT 10.0360 77.5035 10.0620 78.5970 ;
        RECT 9.9280 77.5035 9.9540 78.5970 ;
        RECT 9.8200 77.5035 9.8460 78.5970 ;
        RECT 9.7120 77.5035 9.7380 78.5970 ;
        RECT 9.6040 77.5035 9.6300 78.5970 ;
        RECT 9.4960 77.5035 9.5220 78.5970 ;
        RECT 9.3880 77.5035 9.4140 78.5970 ;
        RECT 9.1750 77.5035 9.2520 78.5970 ;
        RECT 7.2820 77.5035 7.3590 78.5970 ;
        RECT 7.1200 77.5035 7.1460 78.5970 ;
        RECT 7.0120 77.5035 7.0380 78.5970 ;
        RECT 6.9040 77.5035 6.9300 78.5970 ;
        RECT 6.7960 77.5035 6.8220 78.5970 ;
        RECT 6.6880 77.5035 6.7140 78.5970 ;
        RECT 6.5800 77.5035 6.6060 78.5970 ;
        RECT 6.4720 77.5035 6.4980 78.5970 ;
        RECT 6.3640 77.5035 6.3900 78.5970 ;
        RECT 6.2560 77.5035 6.2820 78.5970 ;
        RECT 6.1480 77.5035 6.1740 78.5970 ;
        RECT 6.0400 77.5035 6.0660 78.5970 ;
        RECT 5.9320 77.5035 5.9580 78.5970 ;
        RECT 5.8240 77.5035 5.8500 78.5970 ;
        RECT 5.7160 77.5035 5.7420 78.5970 ;
        RECT 5.6080 77.5035 5.6340 78.5970 ;
        RECT 5.5000 77.5035 5.5260 78.5970 ;
        RECT 5.3920 77.5035 5.4180 78.5970 ;
        RECT 5.2840 77.5035 5.3100 78.5970 ;
        RECT 5.1760 77.5035 5.2020 78.5970 ;
        RECT 5.0680 77.5035 5.0940 78.5970 ;
        RECT 4.9600 77.5035 4.9860 78.5970 ;
        RECT 4.8520 77.5035 4.8780 78.5970 ;
        RECT 4.7440 77.5035 4.7700 78.5970 ;
        RECT 4.6360 77.5035 4.6620 78.5970 ;
        RECT 4.5280 77.5035 4.5540 78.5970 ;
        RECT 4.4200 77.5035 4.4460 78.5970 ;
        RECT 4.3120 77.5035 4.3380 78.5970 ;
        RECT 4.2040 77.5035 4.2300 78.5970 ;
        RECT 4.0960 77.5035 4.1220 78.5970 ;
        RECT 3.9880 77.5035 4.0140 78.5970 ;
        RECT 3.8800 77.5035 3.9060 78.5970 ;
        RECT 3.7720 77.5035 3.7980 78.5970 ;
        RECT 3.6640 77.5035 3.6900 78.5970 ;
        RECT 3.5560 77.5035 3.5820 78.5970 ;
        RECT 3.4480 77.5035 3.4740 78.5970 ;
        RECT 3.3400 77.5035 3.3660 78.5970 ;
        RECT 3.2320 77.5035 3.2580 78.5970 ;
        RECT 3.1240 77.5035 3.1500 78.5970 ;
        RECT 3.0160 77.5035 3.0420 78.5970 ;
        RECT 2.9080 77.5035 2.9340 78.5970 ;
        RECT 2.8000 77.5035 2.8260 78.5970 ;
        RECT 2.6920 77.5035 2.7180 78.5970 ;
        RECT 2.5840 77.5035 2.6100 78.5970 ;
        RECT 2.4760 77.5035 2.5020 78.5970 ;
        RECT 2.3680 77.5035 2.3940 78.5970 ;
        RECT 2.2600 77.5035 2.2860 78.5970 ;
        RECT 2.1520 77.5035 2.1780 78.5970 ;
        RECT 2.0440 77.5035 2.0700 78.5970 ;
        RECT 1.9360 77.5035 1.9620 78.5970 ;
        RECT 1.8280 77.5035 1.8540 78.5970 ;
        RECT 1.7200 77.5035 1.7460 78.5970 ;
        RECT 1.6120 77.5035 1.6380 78.5970 ;
        RECT 1.5040 77.5035 1.5300 78.5970 ;
        RECT 1.3960 77.5035 1.4220 78.5970 ;
        RECT 1.2880 77.5035 1.3140 78.5970 ;
        RECT 1.1800 77.5035 1.2060 78.5970 ;
        RECT 1.0720 77.5035 1.0980 78.5970 ;
        RECT 0.9640 77.5035 0.9900 78.5970 ;
        RECT 0.8560 77.5035 0.8820 78.5970 ;
        RECT 0.7480 77.5035 0.7740 78.5970 ;
        RECT 0.6400 77.5035 0.6660 78.5970 ;
        RECT 0.5320 77.5035 0.5580 78.5970 ;
        RECT 0.4240 77.5035 0.4500 78.5970 ;
        RECT 0.3160 77.5035 0.3420 78.5970 ;
        RECT 0.2080 77.5035 0.2340 78.5970 ;
        RECT 0.0050 77.5035 0.0900 78.5970 ;
        RECT 8.6410 78.5835 8.7690 79.6770 ;
        RECT 8.6270 79.2490 8.7690 79.5715 ;
        RECT 8.4790 78.9760 8.5410 79.6770 ;
        RECT 8.4650 79.2855 8.5410 79.4390 ;
        RECT 8.4790 78.5835 8.5050 79.6770 ;
        RECT 8.4790 78.7045 8.5190 78.9440 ;
        RECT 8.4790 78.5835 8.5410 78.6725 ;
        RECT 8.1820 79.0340 8.3880 79.6770 ;
        RECT 8.3620 78.5835 8.3880 79.6770 ;
        RECT 8.1820 79.3110 8.4020 79.5690 ;
        RECT 8.1820 78.5835 8.2800 79.6770 ;
        RECT 7.7650 78.5835 7.8480 79.6770 ;
        RECT 7.7650 78.6720 7.8620 79.6075 ;
        RECT 16.4440 78.5835 16.5290 79.6770 ;
        RECT 16.3000 78.5835 16.3260 79.6770 ;
        RECT 16.1920 78.5835 16.2180 79.6770 ;
        RECT 16.0840 78.5835 16.1100 79.6770 ;
        RECT 15.9760 78.5835 16.0020 79.6770 ;
        RECT 15.8680 78.5835 15.8940 79.6770 ;
        RECT 15.7600 78.5835 15.7860 79.6770 ;
        RECT 15.6520 78.5835 15.6780 79.6770 ;
        RECT 15.5440 78.5835 15.5700 79.6770 ;
        RECT 15.4360 78.5835 15.4620 79.6770 ;
        RECT 15.3280 78.5835 15.3540 79.6770 ;
        RECT 15.2200 78.5835 15.2460 79.6770 ;
        RECT 15.1120 78.5835 15.1380 79.6770 ;
        RECT 15.0040 78.5835 15.0300 79.6770 ;
        RECT 14.8960 78.5835 14.9220 79.6770 ;
        RECT 14.7880 78.5835 14.8140 79.6770 ;
        RECT 14.6800 78.5835 14.7060 79.6770 ;
        RECT 14.5720 78.5835 14.5980 79.6770 ;
        RECT 14.4640 78.5835 14.4900 79.6770 ;
        RECT 14.3560 78.5835 14.3820 79.6770 ;
        RECT 14.2480 78.5835 14.2740 79.6770 ;
        RECT 14.1400 78.5835 14.1660 79.6770 ;
        RECT 14.0320 78.5835 14.0580 79.6770 ;
        RECT 13.9240 78.5835 13.9500 79.6770 ;
        RECT 13.8160 78.5835 13.8420 79.6770 ;
        RECT 13.7080 78.5835 13.7340 79.6770 ;
        RECT 13.6000 78.5835 13.6260 79.6770 ;
        RECT 13.4920 78.5835 13.5180 79.6770 ;
        RECT 13.3840 78.5835 13.4100 79.6770 ;
        RECT 13.2760 78.5835 13.3020 79.6770 ;
        RECT 13.1680 78.5835 13.1940 79.6770 ;
        RECT 13.0600 78.5835 13.0860 79.6770 ;
        RECT 12.9520 78.5835 12.9780 79.6770 ;
        RECT 12.8440 78.5835 12.8700 79.6770 ;
        RECT 12.7360 78.5835 12.7620 79.6770 ;
        RECT 12.6280 78.5835 12.6540 79.6770 ;
        RECT 12.5200 78.5835 12.5460 79.6770 ;
        RECT 12.4120 78.5835 12.4380 79.6770 ;
        RECT 12.3040 78.5835 12.3300 79.6770 ;
        RECT 12.1960 78.5835 12.2220 79.6770 ;
        RECT 12.0880 78.5835 12.1140 79.6770 ;
        RECT 11.9800 78.5835 12.0060 79.6770 ;
        RECT 11.8720 78.5835 11.8980 79.6770 ;
        RECT 11.7640 78.5835 11.7900 79.6770 ;
        RECT 11.6560 78.5835 11.6820 79.6770 ;
        RECT 11.5480 78.5835 11.5740 79.6770 ;
        RECT 11.4400 78.5835 11.4660 79.6770 ;
        RECT 11.3320 78.5835 11.3580 79.6770 ;
        RECT 11.2240 78.5835 11.2500 79.6770 ;
        RECT 11.1160 78.5835 11.1420 79.6770 ;
        RECT 11.0080 78.5835 11.0340 79.6770 ;
        RECT 10.9000 78.5835 10.9260 79.6770 ;
        RECT 10.7920 78.5835 10.8180 79.6770 ;
        RECT 10.6840 78.5835 10.7100 79.6770 ;
        RECT 10.5760 78.5835 10.6020 79.6770 ;
        RECT 10.4680 78.5835 10.4940 79.6770 ;
        RECT 10.3600 78.5835 10.3860 79.6770 ;
        RECT 10.2520 78.5835 10.2780 79.6770 ;
        RECT 10.1440 78.5835 10.1700 79.6770 ;
        RECT 10.0360 78.5835 10.0620 79.6770 ;
        RECT 9.9280 78.5835 9.9540 79.6770 ;
        RECT 9.8200 78.5835 9.8460 79.6770 ;
        RECT 9.7120 78.5835 9.7380 79.6770 ;
        RECT 9.6040 78.5835 9.6300 79.6770 ;
        RECT 9.4960 78.5835 9.5220 79.6770 ;
        RECT 9.3880 78.5835 9.4140 79.6770 ;
        RECT 9.1750 78.5835 9.2520 79.6770 ;
        RECT 7.2820 78.5835 7.3590 79.6770 ;
        RECT 7.1200 78.5835 7.1460 79.6770 ;
        RECT 7.0120 78.5835 7.0380 79.6770 ;
        RECT 6.9040 78.5835 6.9300 79.6770 ;
        RECT 6.7960 78.5835 6.8220 79.6770 ;
        RECT 6.6880 78.5835 6.7140 79.6770 ;
        RECT 6.5800 78.5835 6.6060 79.6770 ;
        RECT 6.4720 78.5835 6.4980 79.6770 ;
        RECT 6.3640 78.5835 6.3900 79.6770 ;
        RECT 6.2560 78.5835 6.2820 79.6770 ;
        RECT 6.1480 78.5835 6.1740 79.6770 ;
        RECT 6.0400 78.5835 6.0660 79.6770 ;
        RECT 5.9320 78.5835 5.9580 79.6770 ;
        RECT 5.8240 78.5835 5.8500 79.6770 ;
        RECT 5.7160 78.5835 5.7420 79.6770 ;
        RECT 5.6080 78.5835 5.6340 79.6770 ;
        RECT 5.5000 78.5835 5.5260 79.6770 ;
        RECT 5.3920 78.5835 5.4180 79.6770 ;
        RECT 5.2840 78.5835 5.3100 79.6770 ;
        RECT 5.1760 78.5835 5.2020 79.6770 ;
        RECT 5.0680 78.5835 5.0940 79.6770 ;
        RECT 4.9600 78.5835 4.9860 79.6770 ;
        RECT 4.8520 78.5835 4.8780 79.6770 ;
        RECT 4.7440 78.5835 4.7700 79.6770 ;
        RECT 4.6360 78.5835 4.6620 79.6770 ;
        RECT 4.5280 78.5835 4.5540 79.6770 ;
        RECT 4.4200 78.5835 4.4460 79.6770 ;
        RECT 4.3120 78.5835 4.3380 79.6770 ;
        RECT 4.2040 78.5835 4.2300 79.6770 ;
        RECT 4.0960 78.5835 4.1220 79.6770 ;
        RECT 3.9880 78.5835 4.0140 79.6770 ;
        RECT 3.8800 78.5835 3.9060 79.6770 ;
        RECT 3.7720 78.5835 3.7980 79.6770 ;
        RECT 3.6640 78.5835 3.6900 79.6770 ;
        RECT 3.5560 78.5835 3.5820 79.6770 ;
        RECT 3.4480 78.5835 3.4740 79.6770 ;
        RECT 3.3400 78.5835 3.3660 79.6770 ;
        RECT 3.2320 78.5835 3.2580 79.6770 ;
        RECT 3.1240 78.5835 3.1500 79.6770 ;
        RECT 3.0160 78.5835 3.0420 79.6770 ;
        RECT 2.9080 78.5835 2.9340 79.6770 ;
        RECT 2.8000 78.5835 2.8260 79.6770 ;
        RECT 2.6920 78.5835 2.7180 79.6770 ;
        RECT 2.5840 78.5835 2.6100 79.6770 ;
        RECT 2.4760 78.5835 2.5020 79.6770 ;
        RECT 2.3680 78.5835 2.3940 79.6770 ;
        RECT 2.2600 78.5835 2.2860 79.6770 ;
        RECT 2.1520 78.5835 2.1780 79.6770 ;
        RECT 2.0440 78.5835 2.0700 79.6770 ;
        RECT 1.9360 78.5835 1.9620 79.6770 ;
        RECT 1.8280 78.5835 1.8540 79.6770 ;
        RECT 1.7200 78.5835 1.7460 79.6770 ;
        RECT 1.6120 78.5835 1.6380 79.6770 ;
        RECT 1.5040 78.5835 1.5300 79.6770 ;
        RECT 1.3960 78.5835 1.4220 79.6770 ;
        RECT 1.2880 78.5835 1.3140 79.6770 ;
        RECT 1.1800 78.5835 1.2060 79.6770 ;
        RECT 1.0720 78.5835 1.0980 79.6770 ;
        RECT 0.9640 78.5835 0.9900 79.6770 ;
        RECT 0.8560 78.5835 0.8820 79.6770 ;
        RECT 0.7480 78.5835 0.7740 79.6770 ;
        RECT 0.6400 78.5835 0.6660 79.6770 ;
        RECT 0.5320 78.5835 0.5580 79.6770 ;
        RECT 0.4240 78.5835 0.4500 79.6770 ;
        RECT 0.3160 78.5835 0.3420 79.6770 ;
        RECT 0.2080 78.5835 0.2340 79.6770 ;
        RECT 0.0050 78.5835 0.0900 79.6770 ;
        RECT 8.6410 79.6635 8.7690 80.7570 ;
        RECT 8.6270 80.3290 8.7690 80.6515 ;
        RECT 8.4790 80.0560 8.5410 80.7570 ;
        RECT 8.4650 80.3655 8.5410 80.5190 ;
        RECT 8.4790 79.6635 8.5050 80.7570 ;
        RECT 8.4790 79.7845 8.5190 80.0240 ;
        RECT 8.4790 79.6635 8.5410 79.7525 ;
        RECT 8.1820 80.1140 8.3880 80.7570 ;
        RECT 8.3620 79.6635 8.3880 80.7570 ;
        RECT 8.1820 80.3910 8.4020 80.6490 ;
        RECT 8.1820 79.6635 8.2800 80.7570 ;
        RECT 7.7650 79.6635 7.8480 80.7570 ;
        RECT 7.7650 79.7520 7.8620 80.6875 ;
        RECT 16.4440 79.6635 16.5290 80.7570 ;
        RECT 16.3000 79.6635 16.3260 80.7570 ;
        RECT 16.1920 79.6635 16.2180 80.7570 ;
        RECT 16.0840 79.6635 16.1100 80.7570 ;
        RECT 15.9760 79.6635 16.0020 80.7570 ;
        RECT 15.8680 79.6635 15.8940 80.7570 ;
        RECT 15.7600 79.6635 15.7860 80.7570 ;
        RECT 15.6520 79.6635 15.6780 80.7570 ;
        RECT 15.5440 79.6635 15.5700 80.7570 ;
        RECT 15.4360 79.6635 15.4620 80.7570 ;
        RECT 15.3280 79.6635 15.3540 80.7570 ;
        RECT 15.2200 79.6635 15.2460 80.7570 ;
        RECT 15.1120 79.6635 15.1380 80.7570 ;
        RECT 15.0040 79.6635 15.0300 80.7570 ;
        RECT 14.8960 79.6635 14.9220 80.7570 ;
        RECT 14.7880 79.6635 14.8140 80.7570 ;
        RECT 14.6800 79.6635 14.7060 80.7570 ;
        RECT 14.5720 79.6635 14.5980 80.7570 ;
        RECT 14.4640 79.6635 14.4900 80.7570 ;
        RECT 14.3560 79.6635 14.3820 80.7570 ;
        RECT 14.2480 79.6635 14.2740 80.7570 ;
        RECT 14.1400 79.6635 14.1660 80.7570 ;
        RECT 14.0320 79.6635 14.0580 80.7570 ;
        RECT 13.9240 79.6635 13.9500 80.7570 ;
        RECT 13.8160 79.6635 13.8420 80.7570 ;
        RECT 13.7080 79.6635 13.7340 80.7570 ;
        RECT 13.6000 79.6635 13.6260 80.7570 ;
        RECT 13.4920 79.6635 13.5180 80.7570 ;
        RECT 13.3840 79.6635 13.4100 80.7570 ;
        RECT 13.2760 79.6635 13.3020 80.7570 ;
        RECT 13.1680 79.6635 13.1940 80.7570 ;
        RECT 13.0600 79.6635 13.0860 80.7570 ;
        RECT 12.9520 79.6635 12.9780 80.7570 ;
        RECT 12.8440 79.6635 12.8700 80.7570 ;
        RECT 12.7360 79.6635 12.7620 80.7570 ;
        RECT 12.6280 79.6635 12.6540 80.7570 ;
        RECT 12.5200 79.6635 12.5460 80.7570 ;
        RECT 12.4120 79.6635 12.4380 80.7570 ;
        RECT 12.3040 79.6635 12.3300 80.7570 ;
        RECT 12.1960 79.6635 12.2220 80.7570 ;
        RECT 12.0880 79.6635 12.1140 80.7570 ;
        RECT 11.9800 79.6635 12.0060 80.7570 ;
        RECT 11.8720 79.6635 11.8980 80.7570 ;
        RECT 11.7640 79.6635 11.7900 80.7570 ;
        RECT 11.6560 79.6635 11.6820 80.7570 ;
        RECT 11.5480 79.6635 11.5740 80.7570 ;
        RECT 11.4400 79.6635 11.4660 80.7570 ;
        RECT 11.3320 79.6635 11.3580 80.7570 ;
        RECT 11.2240 79.6635 11.2500 80.7570 ;
        RECT 11.1160 79.6635 11.1420 80.7570 ;
        RECT 11.0080 79.6635 11.0340 80.7570 ;
        RECT 10.9000 79.6635 10.9260 80.7570 ;
        RECT 10.7920 79.6635 10.8180 80.7570 ;
        RECT 10.6840 79.6635 10.7100 80.7570 ;
        RECT 10.5760 79.6635 10.6020 80.7570 ;
        RECT 10.4680 79.6635 10.4940 80.7570 ;
        RECT 10.3600 79.6635 10.3860 80.7570 ;
        RECT 10.2520 79.6635 10.2780 80.7570 ;
        RECT 10.1440 79.6635 10.1700 80.7570 ;
        RECT 10.0360 79.6635 10.0620 80.7570 ;
        RECT 9.9280 79.6635 9.9540 80.7570 ;
        RECT 9.8200 79.6635 9.8460 80.7570 ;
        RECT 9.7120 79.6635 9.7380 80.7570 ;
        RECT 9.6040 79.6635 9.6300 80.7570 ;
        RECT 9.4960 79.6635 9.5220 80.7570 ;
        RECT 9.3880 79.6635 9.4140 80.7570 ;
        RECT 9.1750 79.6635 9.2520 80.7570 ;
        RECT 7.2820 79.6635 7.3590 80.7570 ;
        RECT 7.1200 79.6635 7.1460 80.7570 ;
        RECT 7.0120 79.6635 7.0380 80.7570 ;
        RECT 6.9040 79.6635 6.9300 80.7570 ;
        RECT 6.7960 79.6635 6.8220 80.7570 ;
        RECT 6.6880 79.6635 6.7140 80.7570 ;
        RECT 6.5800 79.6635 6.6060 80.7570 ;
        RECT 6.4720 79.6635 6.4980 80.7570 ;
        RECT 6.3640 79.6635 6.3900 80.7570 ;
        RECT 6.2560 79.6635 6.2820 80.7570 ;
        RECT 6.1480 79.6635 6.1740 80.7570 ;
        RECT 6.0400 79.6635 6.0660 80.7570 ;
        RECT 5.9320 79.6635 5.9580 80.7570 ;
        RECT 5.8240 79.6635 5.8500 80.7570 ;
        RECT 5.7160 79.6635 5.7420 80.7570 ;
        RECT 5.6080 79.6635 5.6340 80.7570 ;
        RECT 5.5000 79.6635 5.5260 80.7570 ;
        RECT 5.3920 79.6635 5.4180 80.7570 ;
        RECT 5.2840 79.6635 5.3100 80.7570 ;
        RECT 5.1760 79.6635 5.2020 80.7570 ;
        RECT 5.0680 79.6635 5.0940 80.7570 ;
        RECT 4.9600 79.6635 4.9860 80.7570 ;
        RECT 4.8520 79.6635 4.8780 80.7570 ;
        RECT 4.7440 79.6635 4.7700 80.7570 ;
        RECT 4.6360 79.6635 4.6620 80.7570 ;
        RECT 4.5280 79.6635 4.5540 80.7570 ;
        RECT 4.4200 79.6635 4.4460 80.7570 ;
        RECT 4.3120 79.6635 4.3380 80.7570 ;
        RECT 4.2040 79.6635 4.2300 80.7570 ;
        RECT 4.0960 79.6635 4.1220 80.7570 ;
        RECT 3.9880 79.6635 4.0140 80.7570 ;
        RECT 3.8800 79.6635 3.9060 80.7570 ;
        RECT 3.7720 79.6635 3.7980 80.7570 ;
        RECT 3.6640 79.6635 3.6900 80.7570 ;
        RECT 3.5560 79.6635 3.5820 80.7570 ;
        RECT 3.4480 79.6635 3.4740 80.7570 ;
        RECT 3.3400 79.6635 3.3660 80.7570 ;
        RECT 3.2320 79.6635 3.2580 80.7570 ;
        RECT 3.1240 79.6635 3.1500 80.7570 ;
        RECT 3.0160 79.6635 3.0420 80.7570 ;
        RECT 2.9080 79.6635 2.9340 80.7570 ;
        RECT 2.8000 79.6635 2.8260 80.7570 ;
        RECT 2.6920 79.6635 2.7180 80.7570 ;
        RECT 2.5840 79.6635 2.6100 80.7570 ;
        RECT 2.4760 79.6635 2.5020 80.7570 ;
        RECT 2.3680 79.6635 2.3940 80.7570 ;
        RECT 2.2600 79.6635 2.2860 80.7570 ;
        RECT 2.1520 79.6635 2.1780 80.7570 ;
        RECT 2.0440 79.6635 2.0700 80.7570 ;
        RECT 1.9360 79.6635 1.9620 80.7570 ;
        RECT 1.8280 79.6635 1.8540 80.7570 ;
        RECT 1.7200 79.6635 1.7460 80.7570 ;
        RECT 1.6120 79.6635 1.6380 80.7570 ;
        RECT 1.5040 79.6635 1.5300 80.7570 ;
        RECT 1.3960 79.6635 1.4220 80.7570 ;
        RECT 1.2880 79.6635 1.3140 80.7570 ;
        RECT 1.1800 79.6635 1.2060 80.7570 ;
        RECT 1.0720 79.6635 1.0980 80.7570 ;
        RECT 0.9640 79.6635 0.9900 80.7570 ;
        RECT 0.8560 79.6635 0.8820 80.7570 ;
        RECT 0.7480 79.6635 0.7740 80.7570 ;
        RECT 0.6400 79.6635 0.6660 80.7570 ;
        RECT 0.5320 79.6635 0.5580 80.7570 ;
        RECT 0.4240 79.6635 0.4500 80.7570 ;
        RECT 0.3160 79.6635 0.3420 80.7570 ;
        RECT 0.2080 79.6635 0.2340 80.7570 ;
        RECT 0.0050 79.6635 0.0900 80.7570 ;
        RECT 8.6410 80.7435 8.7690 81.8370 ;
        RECT 8.6270 81.4090 8.7690 81.7315 ;
        RECT 8.4790 81.1360 8.5410 81.8370 ;
        RECT 8.4650 81.4455 8.5410 81.5990 ;
        RECT 8.4790 80.7435 8.5050 81.8370 ;
        RECT 8.4790 80.8645 8.5190 81.1040 ;
        RECT 8.4790 80.7435 8.5410 80.8325 ;
        RECT 8.1820 81.1940 8.3880 81.8370 ;
        RECT 8.3620 80.7435 8.3880 81.8370 ;
        RECT 8.1820 81.4710 8.4020 81.7290 ;
        RECT 8.1820 80.7435 8.2800 81.8370 ;
        RECT 7.7650 80.7435 7.8480 81.8370 ;
        RECT 7.7650 80.8320 7.8620 81.7675 ;
        RECT 16.4440 80.7435 16.5290 81.8370 ;
        RECT 16.3000 80.7435 16.3260 81.8370 ;
        RECT 16.1920 80.7435 16.2180 81.8370 ;
        RECT 16.0840 80.7435 16.1100 81.8370 ;
        RECT 15.9760 80.7435 16.0020 81.8370 ;
        RECT 15.8680 80.7435 15.8940 81.8370 ;
        RECT 15.7600 80.7435 15.7860 81.8370 ;
        RECT 15.6520 80.7435 15.6780 81.8370 ;
        RECT 15.5440 80.7435 15.5700 81.8370 ;
        RECT 15.4360 80.7435 15.4620 81.8370 ;
        RECT 15.3280 80.7435 15.3540 81.8370 ;
        RECT 15.2200 80.7435 15.2460 81.8370 ;
        RECT 15.1120 80.7435 15.1380 81.8370 ;
        RECT 15.0040 80.7435 15.0300 81.8370 ;
        RECT 14.8960 80.7435 14.9220 81.8370 ;
        RECT 14.7880 80.7435 14.8140 81.8370 ;
        RECT 14.6800 80.7435 14.7060 81.8370 ;
        RECT 14.5720 80.7435 14.5980 81.8370 ;
        RECT 14.4640 80.7435 14.4900 81.8370 ;
        RECT 14.3560 80.7435 14.3820 81.8370 ;
        RECT 14.2480 80.7435 14.2740 81.8370 ;
        RECT 14.1400 80.7435 14.1660 81.8370 ;
        RECT 14.0320 80.7435 14.0580 81.8370 ;
        RECT 13.9240 80.7435 13.9500 81.8370 ;
        RECT 13.8160 80.7435 13.8420 81.8370 ;
        RECT 13.7080 80.7435 13.7340 81.8370 ;
        RECT 13.6000 80.7435 13.6260 81.8370 ;
        RECT 13.4920 80.7435 13.5180 81.8370 ;
        RECT 13.3840 80.7435 13.4100 81.8370 ;
        RECT 13.2760 80.7435 13.3020 81.8370 ;
        RECT 13.1680 80.7435 13.1940 81.8370 ;
        RECT 13.0600 80.7435 13.0860 81.8370 ;
        RECT 12.9520 80.7435 12.9780 81.8370 ;
        RECT 12.8440 80.7435 12.8700 81.8370 ;
        RECT 12.7360 80.7435 12.7620 81.8370 ;
        RECT 12.6280 80.7435 12.6540 81.8370 ;
        RECT 12.5200 80.7435 12.5460 81.8370 ;
        RECT 12.4120 80.7435 12.4380 81.8370 ;
        RECT 12.3040 80.7435 12.3300 81.8370 ;
        RECT 12.1960 80.7435 12.2220 81.8370 ;
        RECT 12.0880 80.7435 12.1140 81.8370 ;
        RECT 11.9800 80.7435 12.0060 81.8370 ;
        RECT 11.8720 80.7435 11.8980 81.8370 ;
        RECT 11.7640 80.7435 11.7900 81.8370 ;
        RECT 11.6560 80.7435 11.6820 81.8370 ;
        RECT 11.5480 80.7435 11.5740 81.8370 ;
        RECT 11.4400 80.7435 11.4660 81.8370 ;
        RECT 11.3320 80.7435 11.3580 81.8370 ;
        RECT 11.2240 80.7435 11.2500 81.8370 ;
        RECT 11.1160 80.7435 11.1420 81.8370 ;
        RECT 11.0080 80.7435 11.0340 81.8370 ;
        RECT 10.9000 80.7435 10.9260 81.8370 ;
        RECT 10.7920 80.7435 10.8180 81.8370 ;
        RECT 10.6840 80.7435 10.7100 81.8370 ;
        RECT 10.5760 80.7435 10.6020 81.8370 ;
        RECT 10.4680 80.7435 10.4940 81.8370 ;
        RECT 10.3600 80.7435 10.3860 81.8370 ;
        RECT 10.2520 80.7435 10.2780 81.8370 ;
        RECT 10.1440 80.7435 10.1700 81.8370 ;
        RECT 10.0360 80.7435 10.0620 81.8370 ;
        RECT 9.9280 80.7435 9.9540 81.8370 ;
        RECT 9.8200 80.7435 9.8460 81.8370 ;
        RECT 9.7120 80.7435 9.7380 81.8370 ;
        RECT 9.6040 80.7435 9.6300 81.8370 ;
        RECT 9.4960 80.7435 9.5220 81.8370 ;
        RECT 9.3880 80.7435 9.4140 81.8370 ;
        RECT 9.1750 80.7435 9.2520 81.8370 ;
        RECT 7.2820 80.7435 7.3590 81.8370 ;
        RECT 7.1200 80.7435 7.1460 81.8370 ;
        RECT 7.0120 80.7435 7.0380 81.8370 ;
        RECT 6.9040 80.7435 6.9300 81.8370 ;
        RECT 6.7960 80.7435 6.8220 81.8370 ;
        RECT 6.6880 80.7435 6.7140 81.8370 ;
        RECT 6.5800 80.7435 6.6060 81.8370 ;
        RECT 6.4720 80.7435 6.4980 81.8370 ;
        RECT 6.3640 80.7435 6.3900 81.8370 ;
        RECT 6.2560 80.7435 6.2820 81.8370 ;
        RECT 6.1480 80.7435 6.1740 81.8370 ;
        RECT 6.0400 80.7435 6.0660 81.8370 ;
        RECT 5.9320 80.7435 5.9580 81.8370 ;
        RECT 5.8240 80.7435 5.8500 81.8370 ;
        RECT 5.7160 80.7435 5.7420 81.8370 ;
        RECT 5.6080 80.7435 5.6340 81.8370 ;
        RECT 5.5000 80.7435 5.5260 81.8370 ;
        RECT 5.3920 80.7435 5.4180 81.8370 ;
        RECT 5.2840 80.7435 5.3100 81.8370 ;
        RECT 5.1760 80.7435 5.2020 81.8370 ;
        RECT 5.0680 80.7435 5.0940 81.8370 ;
        RECT 4.9600 80.7435 4.9860 81.8370 ;
        RECT 4.8520 80.7435 4.8780 81.8370 ;
        RECT 4.7440 80.7435 4.7700 81.8370 ;
        RECT 4.6360 80.7435 4.6620 81.8370 ;
        RECT 4.5280 80.7435 4.5540 81.8370 ;
        RECT 4.4200 80.7435 4.4460 81.8370 ;
        RECT 4.3120 80.7435 4.3380 81.8370 ;
        RECT 4.2040 80.7435 4.2300 81.8370 ;
        RECT 4.0960 80.7435 4.1220 81.8370 ;
        RECT 3.9880 80.7435 4.0140 81.8370 ;
        RECT 3.8800 80.7435 3.9060 81.8370 ;
        RECT 3.7720 80.7435 3.7980 81.8370 ;
        RECT 3.6640 80.7435 3.6900 81.8370 ;
        RECT 3.5560 80.7435 3.5820 81.8370 ;
        RECT 3.4480 80.7435 3.4740 81.8370 ;
        RECT 3.3400 80.7435 3.3660 81.8370 ;
        RECT 3.2320 80.7435 3.2580 81.8370 ;
        RECT 3.1240 80.7435 3.1500 81.8370 ;
        RECT 3.0160 80.7435 3.0420 81.8370 ;
        RECT 2.9080 80.7435 2.9340 81.8370 ;
        RECT 2.8000 80.7435 2.8260 81.8370 ;
        RECT 2.6920 80.7435 2.7180 81.8370 ;
        RECT 2.5840 80.7435 2.6100 81.8370 ;
        RECT 2.4760 80.7435 2.5020 81.8370 ;
        RECT 2.3680 80.7435 2.3940 81.8370 ;
        RECT 2.2600 80.7435 2.2860 81.8370 ;
        RECT 2.1520 80.7435 2.1780 81.8370 ;
        RECT 2.0440 80.7435 2.0700 81.8370 ;
        RECT 1.9360 80.7435 1.9620 81.8370 ;
        RECT 1.8280 80.7435 1.8540 81.8370 ;
        RECT 1.7200 80.7435 1.7460 81.8370 ;
        RECT 1.6120 80.7435 1.6380 81.8370 ;
        RECT 1.5040 80.7435 1.5300 81.8370 ;
        RECT 1.3960 80.7435 1.4220 81.8370 ;
        RECT 1.2880 80.7435 1.3140 81.8370 ;
        RECT 1.1800 80.7435 1.2060 81.8370 ;
        RECT 1.0720 80.7435 1.0980 81.8370 ;
        RECT 0.9640 80.7435 0.9900 81.8370 ;
        RECT 0.8560 80.7435 0.8820 81.8370 ;
        RECT 0.7480 80.7435 0.7740 81.8370 ;
        RECT 0.6400 80.7435 0.6660 81.8370 ;
        RECT 0.5320 80.7435 0.5580 81.8370 ;
        RECT 0.4240 80.7435 0.4500 81.8370 ;
        RECT 0.3160 80.7435 0.3420 81.8370 ;
        RECT 0.2080 80.7435 0.2340 81.8370 ;
        RECT 0.0050 80.7435 0.0900 81.8370 ;
        RECT 8.6410 81.8235 8.7690 82.9170 ;
        RECT 8.6270 82.4890 8.7690 82.8115 ;
        RECT 8.4790 82.2160 8.5410 82.9170 ;
        RECT 8.4650 82.5255 8.5410 82.6790 ;
        RECT 8.4790 81.8235 8.5050 82.9170 ;
        RECT 8.4790 81.9445 8.5190 82.1840 ;
        RECT 8.4790 81.8235 8.5410 81.9125 ;
        RECT 8.1820 82.2740 8.3880 82.9170 ;
        RECT 8.3620 81.8235 8.3880 82.9170 ;
        RECT 8.1820 82.5510 8.4020 82.8090 ;
        RECT 8.1820 81.8235 8.2800 82.9170 ;
        RECT 7.7650 81.8235 7.8480 82.9170 ;
        RECT 7.7650 81.9120 7.8620 82.8475 ;
        RECT 16.4440 81.8235 16.5290 82.9170 ;
        RECT 16.3000 81.8235 16.3260 82.9170 ;
        RECT 16.1920 81.8235 16.2180 82.9170 ;
        RECT 16.0840 81.8235 16.1100 82.9170 ;
        RECT 15.9760 81.8235 16.0020 82.9170 ;
        RECT 15.8680 81.8235 15.8940 82.9170 ;
        RECT 15.7600 81.8235 15.7860 82.9170 ;
        RECT 15.6520 81.8235 15.6780 82.9170 ;
        RECT 15.5440 81.8235 15.5700 82.9170 ;
        RECT 15.4360 81.8235 15.4620 82.9170 ;
        RECT 15.3280 81.8235 15.3540 82.9170 ;
        RECT 15.2200 81.8235 15.2460 82.9170 ;
        RECT 15.1120 81.8235 15.1380 82.9170 ;
        RECT 15.0040 81.8235 15.0300 82.9170 ;
        RECT 14.8960 81.8235 14.9220 82.9170 ;
        RECT 14.7880 81.8235 14.8140 82.9170 ;
        RECT 14.6800 81.8235 14.7060 82.9170 ;
        RECT 14.5720 81.8235 14.5980 82.9170 ;
        RECT 14.4640 81.8235 14.4900 82.9170 ;
        RECT 14.3560 81.8235 14.3820 82.9170 ;
        RECT 14.2480 81.8235 14.2740 82.9170 ;
        RECT 14.1400 81.8235 14.1660 82.9170 ;
        RECT 14.0320 81.8235 14.0580 82.9170 ;
        RECT 13.9240 81.8235 13.9500 82.9170 ;
        RECT 13.8160 81.8235 13.8420 82.9170 ;
        RECT 13.7080 81.8235 13.7340 82.9170 ;
        RECT 13.6000 81.8235 13.6260 82.9170 ;
        RECT 13.4920 81.8235 13.5180 82.9170 ;
        RECT 13.3840 81.8235 13.4100 82.9170 ;
        RECT 13.2760 81.8235 13.3020 82.9170 ;
        RECT 13.1680 81.8235 13.1940 82.9170 ;
        RECT 13.0600 81.8235 13.0860 82.9170 ;
        RECT 12.9520 81.8235 12.9780 82.9170 ;
        RECT 12.8440 81.8235 12.8700 82.9170 ;
        RECT 12.7360 81.8235 12.7620 82.9170 ;
        RECT 12.6280 81.8235 12.6540 82.9170 ;
        RECT 12.5200 81.8235 12.5460 82.9170 ;
        RECT 12.4120 81.8235 12.4380 82.9170 ;
        RECT 12.3040 81.8235 12.3300 82.9170 ;
        RECT 12.1960 81.8235 12.2220 82.9170 ;
        RECT 12.0880 81.8235 12.1140 82.9170 ;
        RECT 11.9800 81.8235 12.0060 82.9170 ;
        RECT 11.8720 81.8235 11.8980 82.9170 ;
        RECT 11.7640 81.8235 11.7900 82.9170 ;
        RECT 11.6560 81.8235 11.6820 82.9170 ;
        RECT 11.5480 81.8235 11.5740 82.9170 ;
        RECT 11.4400 81.8235 11.4660 82.9170 ;
        RECT 11.3320 81.8235 11.3580 82.9170 ;
        RECT 11.2240 81.8235 11.2500 82.9170 ;
        RECT 11.1160 81.8235 11.1420 82.9170 ;
        RECT 11.0080 81.8235 11.0340 82.9170 ;
        RECT 10.9000 81.8235 10.9260 82.9170 ;
        RECT 10.7920 81.8235 10.8180 82.9170 ;
        RECT 10.6840 81.8235 10.7100 82.9170 ;
        RECT 10.5760 81.8235 10.6020 82.9170 ;
        RECT 10.4680 81.8235 10.4940 82.9170 ;
        RECT 10.3600 81.8235 10.3860 82.9170 ;
        RECT 10.2520 81.8235 10.2780 82.9170 ;
        RECT 10.1440 81.8235 10.1700 82.9170 ;
        RECT 10.0360 81.8235 10.0620 82.9170 ;
        RECT 9.9280 81.8235 9.9540 82.9170 ;
        RECT 9.8200 81.8235 9.8460 82.9170 ;
        RECT 9.7120 81.8235 9.7380 82.9170 ;
        RECT 9.6040 81.8235 9.6300 82.9170 ;
        RECT 9.4960 81.8235 9.5220 82.9170 ;
        RECT 9.3880 81.8235 9.4140 82.9170 ;
        RECT 9.1750 81.8235 9.2520 82.9170 ;
        RECT 7.2820 81.8235 7.3590 82.9170 ;
        RECT 7.1200 81.8235 7.1460 82.9170 ;
        RECT 7.0120 81.8235 7.0380 82.9170 ;
        RECT 6.9040 81.8235 6.9300 82.9170 ;
        RECT 6.7960 81.8235 6.8220 82.9170 ;
        RECT 6.6880 81.8235 6.7140 82.9170 ;
        RECT 6.5800 81.8235 6.6060 82.9170 ;
        RECT 6.4720 81.8235 6.4980 82.9170 ;
        RECT 6.3640 81.8235 6.3900 82.9170 ;
        RECT 6.2560 81.8235 6.2820 82.9170 ;
        RECT 6.1480 81.8235 6.1740 82.9170 ;
        RECT 6.0400 81.8235 6.0660 82.9170 ;
        RECT 5.9320 81.8235 5.9580 82.9170 ;
        RECT 5.8240 81.8235 5.8500 82.9170 ;
        RECT 5.7160 81.8235 5.7420 82.9170 ;
        RECT 5.6080 81.8235 5.6340 82.9170 ;
        RECT 5.5000 81.8235 5.5260 82.9170 ;
        RECT 5.3920 81.8235 5.4180 82.9170 ;
        RECT 5.2840 81.8235 5.3100 82.9170 ;
        RECT 5.1760 81.8235 5.2020 82.9170 ;
        RECT 5.0680 81.8235 5.0940 82.9170 ;
        RECT 4.9600 81.8235 4.9860 82.9170 ;
        RECT 4.8520 81.8235 4.8780 82.9170 ;
        RECT 4.7440 81.8235 4.7700 82.9170 ;
        RECT 4.6360 81.8235 4.6620 82.9170 ;
        RECT 4.5280 81.8235 4.5540 82.9170 ;
        RECT 4.4200 81.8235 4.4460 82.9170 ;
        RECT 4.3120 81.8235 4.3380 82.9170 ;
        RECT 4.2040 81.8235 4.2300 82.9170 ;
        RECT 4.0960 81.8235 4.1220 82.9170 ;
        RECT 3.9880 81.8235 4.0140 82.9170 ;
        RECT 3.8800 81.8235 3.9060 82.9170 ;
        RECT 3.7720 81.8235 3.7980 82.9170 ;
        RECT 3.6640 81.8235 3.6900 82.9170 ;
        RECT 3.5560 81.8235 3.5820 82.9170 ;
        RECT 3.4480 81.8235 3.4740 82.9170 ;
        RECT 3.3400 81.8235 3.3660 82.9170 ;
        RECT 3.2320 81.8235 3.2580 82.9170 ;
        RECT 3.1240 81.8235 3.1500 82.9170 ;
        RECT 3.0160 81.8235 3.0420 82.9170 ;
        RECT 2.9080 81.8235 2.9340 82.9170 ;
        RECT 2.8000 81.8235 2.8260 82.9170 ;
        RECT 2.6920 81.8235 2.7180 82.9170 ;
        RECT 2.5840 81.8235 2.6100 82.9170 ;
        RECT 2.4760 81.8235 2.5020 82.9170 ;
        RECT 2.3680 81.8235 2.3940 82.9170 ;
        RECT 2.2600 81.8235 2.2860 82.9170 ;
        RECT 2.1520 81.8235 2.1780 82.9170 ;
        RECT 2.0440 81.8235 2.0700 82.9170 ;
        RECT 1.9360 81.8235 1.9620 82.9170 ;
        RECT 1.8280 81.8235 1.8540 82.9170 ;
        RECT 1.7200 81.8235 1.7460 82.9170 ;
        RECT 1.6120 81.8235 1.6380 82.9170 ;
        RECT 1.5040 81.8235 1.5300 82.9170 ;
        RECT 1.3960 81.8235 1.4220 82.9170 ;
        RECT 1.2880 81.8235 1.3140 82.9170 ;
        RECT 1.1800 81.8235 1.2060 82.9170 ;
        RECT 1.0720 81.8235 1.0980 82.9170 ;
        RECT 0.9640 81.8235 0.9900 82.9170 ;
        RECT 0.8560 81.8235 0.8820 82.9170 ;
        RECT 0.7480 81.8235 0.7740 82.9170 ;
        RECT 0.6400 81.8235 0.6660 82.9170 ;
        RECT 0.5320 81.8235 0.5580 82.9170 ;
        RECT 0.4240 81.8235 0.4500 82.9170 ;
        RECT 0.3160 81.8235 0.3420 82.9170 ;
        RECT 0.2080 81.8235 0.2340 82.9170 ;
        RECT 0.0050 81.8235 0.0900 82.9170 ;
        RECT 8.6410 82.9035 8.7690 83.9970 ;
        RECT 8.6270 83.5690 8.7690 83.8915 ;
        RECT 8.4790 83.2960 8.5410 83.9970 ;
        RECT 8.4650 83.6055 8.5410 83.7590 ;
        RECT 8.4790 82.9035 8.5050 83.9970 ;
        RECT 8.4790 83.0245 8.5190 83.2640 ;
        RECT 8.4790 82.9035 8.5410 82.9925 ;
        RECT 8.1820 83.3540 8.3880 83.9970 ;
        RECT 8.3620 82.9035 8.3880 83.9970 ;
        RECT 8.1820 83.6310 8.4020 83.8890 ;
        RECT 8.1820 82.9035 8.2800 83.9970 ;
        RECT 7.7650 82.9035 7.8480 83.9970 ;
        RECT 7.7650 82.9920 7.8620 83.9275 ;
        RECT 16.4440 82.9035 16.5290 83.9970 ;
        RECT 16.3000 82.9035 16.3260 83.9970 ;
        RECT 16.1920 82.9035 16.2180 83.9970 ;
        RECT 16.0840 82.9035 16.1100 83.9970 ;
        RECT 15.9760 82.9035 16.0020 83.9970 ;
        RECT 15.8680 82.9035 15.8940 83.9970 ;
        RECT 15.7600 82.9035 15.7860 83.9970 ;
        RECT 15.6520 82.9035 15.6780 83.9970 ;
        RECT 15.5440 82.9035 15.5700 83.9970 ;
        RECT 15.4360 82.9035 15.4620 83.9970 ;
        RECT 15.3280 82.9035 15.3540 83.9970 ;
        RECT 15.2200 82.9035 15.2460 83.9970 ;
        RECT 15.1120 82.9035 15.1380 83.9970 ;
        RECT 15.0040 82.9035 15.0300 83.9970 ;
        RECT 14.8960 82.9035 14.9220 83.9970 ;
        RECT 14.7880 82.9035 14.8140 83.9970 ;
        RECT 14.6800 82.9035 14.7060 83.9970 ;
        RECT 14.5720 82.9035 14.5980 83.9970 ;
        RECT 14.4640 82.9035 14.4900 83.9970 ;
        RECT 14.3560 82.9035 14.3820 83.9970 ;
        RECT 14.2480 82.9035 14.2740 83.9970 ;
        RECT 14.1400 82.9035 14.1660 83.9970 ;
        RECT 14.0320 82.9035 14.0580 83.9970 ;
        RECT 13.9240 82.9035 13.9500 83.9970 ;
        RECT 13.8160 82.9035 13.8420 83.9970 ;
        RECT 13.7080 82.9035 13.7340 83.9970 ;
        RECT 13.6000 82.9035 13.6260 83.9970 ;
        RECT 13.4920 82.9035 13.5180 83.9970 ;
        RECT 13.3840 82.9035 13.4100 83.9970 ;
        RECT 13.2760 82.9035 13.3020 83.9970 ;
        RECT 13.1680 82.9035 13.1940 83.9970 ;
        RECT 13.0600 82.9035 13.0860 83.9970 ;
        RECT 12.9520 82.9035 12.9780 83.9970 ;
        RECT 12.8440 82.9035 12.8700 83.9970 ;
        RECT 12.7360 82.9035 12.7620 83.9970 ;
        RECT 12.6280 82.9035 12.6540 83.9970 ;
        RECT 12.5200 82.9035 12.5460 83.9970 ;
        RECT 12.4120 82.9035 12.4380 83.9970 ;
        RECT 12.3040 82.9035 12.3300 83.9970 ;
        RECT 12.1960 82.9035 12.2220 83.9970 ;
        RECT 12.0880 82.9035 12.1140 83.9970 ;
        RECT 11.9800 82.9035 12.0060 83.9970 ;
        RECT 11.8720 82.9035 11.8980 83.9970 ;
        RECT 11.7640 82.9035 11.7900 83.9970 ;
        RECT 11.6560 82.9035 11.6820 83.9970 ;
        RECT 11.5480 82.9035 11.5740 83.9970 ;
        RECT 11.4400 82.9035 11.4660 83.9970 ;
        RECT 11.3320 82.9035 11.3580 83.9970 ;
        RECT 11.2240 82.9035 11.2500 83.9970 ;
        RECT 11.1160 82.9035 11.1420 83.9970 ;
        RECT 11.0080 82.9035 11.0340 83.9970 ;
        RECT 10.9000 82.9035 10.9260 83.9970 ;
        RECT 10.7920 82.9035 10.8180 83.9970 ;
        RECT 10.6840 82.9035 10.7100 83.9970 ;
        RECT 10.5760 82.9035 10.6020 83.9970 ;
        RECT 10.4680 82.9035 10.4940 83.9970 ;
        RECT 10.3600 82.9035 10.3860 83.9970 ;
        RECT 10.2520 82.9035 10.2780 83.9970 ;
        RECT 10.1440 82.9035 10.1700 83.9970 ;
        RECT 10.0360 82.9035 10.0620 83.9970 ;
        RECT 9.9280 82.9035 9.9540 83.9970 ;
        RECT 9.8200 82.9035 9.8460 83.9970 ;
        RECT 9.7120 82.9035 9.7380 83.9970 ;
        RECT 9.6040 82.9035 9.6300 83.9970 ;
        RECT 9.4960 82.9035 9.5220 83.9970 ;
        RECT 9.3880 82.9035 9.4140 83.9970 ;
        RECT 9.1750 82.9035 9.2520 83.9970 ;
        RECT 7.2820 82.9035 7.3590 83.9970 ;
        RECT 7.1200 82.9035 7.1460 83.9970 ;
        RECT 7.0120 82.9035 7.0380 83.9970 ;
        RECT 6.9040 82.9035 6.9300 83.9970 ;
        RECT 6.7960 82.9035 6.8220 83.9970 ;
        RECT 6.6880 82.9035 6.7140 83.9970 ;
        RECT 6.5800 82.9035 6.6060 83.9970 ;
        RECT 6.4720 82.9035 6.4980 83.9970 ;
        RECT 6.3640 82.9035 6.3900 83.9970 ;
        RECT 6.2560 82.9035 6.2820 83.9970 ;
        RECT 6.1480 82.9035 6.1740 83.9970 ;
        RECT 6.0400 82.9035 6.0660 83.9970 ;
        RECT 5.9320 82.9035 5.9580 83.9970 ;
        RECT 5.8240 82.9035 5.8500 83.9970 ;
        RECT 5.7160 82.9035 5.7420 83.9970 ;
        RECT 5.6080 82.9035 5.6340 83.9970 ;
        RECT 5.5000 82.9035 5.5260 83.9970 ;
        RECT 5.3920 82.9035 5.4180 83.9970 ;
        RECT 5.2840 82.9035 5.3100 83.9970 ;
        RECT 5.1760 82.9035 5.2020 83.9970 ;
        RECT 5.0680 82.9035 5.0940 83.9970 ;
        RECT 4.9600 82.9035 4.9860 83.9970 ;
        RECT 4.8520 82.9035 4.8780 83.9970 ;
        RECT 4.7440 82.9035 4.7700 83.9970 ;
        RECT 4.6360 82.9035 4.6620 83.9970 ;
        RECT 4.5280 82.9035 4.5540 83.9970 ;
        RECT 4.4200 82.9035 4.4460 83.9970 ;
        RECT 4.3120 82.9035 4.3380 83.9970 ;
        RECT 4.2040 82.9035 4.2300 83.9970 ;
        RECT 4.0960 82.9035 4.1220 83.9970 ;
        RECT 3.9880 82.9035 4.0140 83.9970 ;
        RECT 3.8800 82.9035 3.9060 83.9970 ;
        RECT 3.7720 82.9035 3.7980 83.9970 ;
        RECT 3.6640 82.9035 3.6900 83.9970 ;
        RECT 3.5560 82.9035 3.5820 83.9970 ;
        RECT 3.4480 82.9035 3.4740 83.9970 ;
        RECT 3.3400 82.9035 3.3660 83.9970 ;
        RECT 3.2320 82.9035 3.2580 83.9970 ;
        RECT 3.1240 82.9035 3.1500 83.9970 ;
        RECT 3.0160 82.9035 3.0420 83.9970 ;
        RECT 2.9080 82.9035 2.9340 83.9970 ;
        RECT 2.8000 82.9035 2.8260 83.9970 ;
        RECT 2.6920 82.9035 2.7180 83.9970 ;
        RECT 2.5840 82.9035 2.6100 83.9970 ;
        RECT 2.4760 82.9035 2.5020 83.9970 ;
        RECT 2.3680 82.9035 2.3940 83.9970 ;
        RECT 2.2600 82.9035 2.2860 83.9970 ;
        RECT 2.1520 82.9035 2.1780 83.9970 ;
        RECT 2.0440 82.9035 2.0700 83.9970 ;
        RECT 1.9360 82.9035 1.9620 83.9970 ;
        RECT 1.8280 82.9035 1.8540 83.9970 ;
        RECT 1.7200 82.9035 1.7460 83.9970 ;
        RECT 1.6120 82.9035 1.6380 83.9970 ;
        RECT 1.5040 82.9035 1.5300 83.9970 ;
        RECT 1.3960 82.9035 1.4220 83.9970 ;
        RECT 1.2880 82.9035 1.3140 83.9970 ;
        RECT 1.1800 82.9035 1.2060 83.9970 ;
        RECT 1.0720 82.9035 1.0980 83.9970 ;
        RECT 0.9640 82.9035 0.9900 83.9970 ;
        RECT 0.8560 82.9035 0.8820 83.9970 ;
        RECT 0.7480 82.9035 0.7740 83.9970 ;
        RECT 0.6400 82.9035 0.6660 83.9970 ;
        RECT 0.5320 82.9035 0.5580 83.9970 ;
        RECT 0.4240 82.9035 0.4500 83.9970 ;
        RECT 0.3160 82.9035 0.3420 83.9970 ;
        RECT 0.2080 82.9035 0.2340 83.9970 ;
        RECT 0.0050 82.9035 0.0900 83.9970 ;
        RECT 8.6410 83.9835 8.7690 85.0770 ;
        RECT 8.6270 84.6490 8.7690 84.9715 ;
        RECT 8.4790 84.3760 8.5410 85.0770 ;
        RECT 8.4650 84.6855 8.5410 84.8390 ;
        RECT 8.4790 83.9835 8.5050 85.0770 ;
        RECT 8.4790 84.1045 8.5190 84.3440 ;
        RECT 8.4790 83.9835 8.5410 84.0725 ;
        RECT 8.1820 84.4340 8.3880 85.0770 ;
        RECT 8.3620 83.9835 8.3880 85.0770 ;
        RECT 8.1820 84.7110 8.4020 84.9690 ;
        RECT 8.1820 83.9835 8.2800 85.0770 ;
        RECT 7.7650 83.9835 7.8480 85.0770 ;
        RECT 7.7650 84.0720 7.8620 85.0075 ;
        RECT 16.4440 83.9835 16.5290 85.0770 ;
        RECT 16.3000 83.9835 16.3260 85.0770 ;
        RECT 16.1920 83.9835 16.2180 85.0770 ;
        RECT 16.0840 83.9835 16.1100 85.0770 ;
        RECT 15.9760 83.9835 16.0020 85.0770 ;
        RECT 15.8680 83.9835 15.8940 85.0770 ;
        RECT 15.7600 83.9835 15.7860 85.0770 ;
        RECT 15.6520 83.9835 15.6780 85.0770 ;
        RECT 15.5440 83.9835 15.5700 85.0770 ;
        RECT 15.4360 83.9835 15.4620 85.0770 ;
        RECT 15.3280 83.9835 15.3540 85.0770 ;
        RECT 15.2200 83.9835 15.2460 85.0770 ;
        RECT 15.1120 83.9835 15.1380 85.0770 ;
        RECT 15.0040 83.9835 15.0300 85.0770 ;
        RECT 14.8960 83.9835 14.9220 85.0770 ;
        RECT 14.7880 83.9835 14.8140 85.0770 ;
        RECT 14.6800 83.9835 14.7060 85.0770 ;
        RECT 14.5720 83.9835 14.5980 85.0770 ;
        RECT 14.4640 83.9835 14.4900 85.0770 ;
        RECT 14.3560 83.9835 14.3820 85.0770 ;
        RECT 14.2480 83.9835 14.2740 85.0770 ;
        RECT 14.1400 83.9835 14.1660 85.0770 ;
        RECT 14.0320 83.9835 14.0580 85.0770 ;
        RECT 13.9240 83.9835 13.9500 85.0770 ;
        RECT 13.8160 83.9835 13.8420 85.0770 ;
        RECT 13.7080 83.9835 13.7340 85.0770 ;
        RECT 13.6000 83.9835 13.6260 85.0770 ;
        RECT 13.4920 83.9835 13.5180 85.0770 ;
        RECT 13.3840 83.9835 13.4100 85.0770 ;
        RECT 13.2760 83.9835 13.3020 85.0770 ;
        RECT 13.1680 83.9835 13.1940 85.0770 ;
        RECT 13.0600 83.9835 13.0860 85.0770 ;
        RECT 12.9520 83.9835 12.9780 85.0770 ;
        RECT 12.8440 83.9835 12.8700 85.0770 ;
        RECT 12.7360 83.9835 12.7620 85.0770 ;
        RECT 12.6280 83.9835 12.6540 85.0770 ;
        RECT 12.5200 83.9835 12.5460 85.0770 ;
        RECT 12.4120 83.9835 12.4380 85.0770 ;
        RECT 12.3040 83.9835 12.3300 85.0770 ;
        RECT 12.1960 83.9835 12.2220 85.0770 ;
        RECT 12.0880 83.9835 12.1140 85.0770 ;
        RECT 11.9800 83.9835 12.0060 85.0770 ;
        RECT 11.8720 83.9835 11.8980 85.0770 ;
        RECT 11.7640 83.9835 11.7900 85.0770 ;
        RECT 11.6560 83.9835 11.6820 85.0770 ;
        RECT 11.5480 83.9835 11.5740 85.0770 ;
        RECT 11.4400 83.9835 11.4660 85.0770 ;
        RECT 11.3320 83.9835 11.3580 85.0770 ;
        RECT 11.2240 83.9835 11.2500 85.0770 ;
        RECT 11.1160 83.9835 11.1420 85.0770 ;
        RECT 11.0080 83.9835 11.0340 85.0770 ;
        RECT 10.9000 83.9835 10.9260 85.0770 ;
        RECT 10.7920 83.9835 10.8180 85.0770 ;
        RECT 10.6840 83.9835 10.7100 85.0770 ;
        RECT 10.5760 83.9835 10.6020 85.0770 ;
        RECT 10.4680 83.9835 10.4940 85.0770 ;
        RECT 10.3600 83.9835 10.3860 85.0770 ;
        RECT 10.2520 83.9835 10.2780 85.0770 ;
        RECT 10.1440 83.9835 10.1700 85.0770 ;
        RECT 10.0360 83.9835 10.0620 85.0770 ;
        RECT 9.9280 83.9835 9.9540 85.0770 ;
        RECT 9.8200 83.9835 9.8460 85.0770 ;
        RECT 9.7120 83.9835 9.7380 85.0770 ;
        RECT 9.6040 83.9835 9.6300 85.0770 ;
        RECT 9.4960 83.9835 9.5220 85.0770 ;
        RECT 9.3880 83.9835 9.4140 85.0770 ;
        RECT 9.1750 83.9835 9.2520 85.0770 ;
        RECT 7.2820 83.9835 7.3590 85.0770 ;
        RECT 7.1200 83.9835 7.1460 85.0770 ;
        RECT 7.0120 83.9835 7.0380 85.0770 ;
        RECT 6.9040 83.9835 6.9300 85.0770 ;
        RECT 6.7960 83.9835 6.8220 85.0770 ;
        RECT 6.6880 83.9835 6.7140 85.0770 ;
        RECT 6.5800 83.9835 6.6060 85.0770 ;
        RECT 6.4720 83.9835 6.4980 85.0770 ;
        RECT 6.3640 83.9835 6.3900 85.0770 ;
        RECT 6.2560 83.9835 6.2820 85.0770 ;
        RECT 6.1480 83.9835 6.1740 85.0770 ;
        RECT 6.0400 83.9835 6.0660 85.0770 ;
        RECT 5.9320 83.9835 5.9580 85.0770 ;
        RECT 5.8240 83.9835 5.8500 85.0770 ;
        RECT 5.7160 83.9835 5.7420 85.0770 ;
        RECT 5.6080 83.9835 5.6340 85.0770 ;
        RECT 5.5000 83.9835 5.5260 85.0770 ;
        RECT 5.3920 83.9835 5.4180 85.0770 ;
        RECT 5.2840 83.9835 5.3100 85.0770 ;
        RECT 5.1760 83.9835 5.2020 85.0770 ;
        RECT 5.0680 83.9835 5.0940 85.0770 ;
        RECT 4.9600 83.9835 4.9860 85.0770 ;
        RECT 4.8520 83.9835 4.8780 85.0770 ;
        RECT 4.7440 83.9835 4.7700 85.0770 ;
        RECT 4.6360 83.9835 4.6620 85.0770 ;
        RECT 4.5280 83.9835 4.5540 85.0770 ;
        RECT 4.4200 83.9835 4.4460 85.0770 ;
        RECT 4.3120 83.9835 4.3380 85.0770 ;
        RECT 4.2040 83.9835 4.2300 85.0770 ;
        RECT 4.0960 83.9835 4.1220 85.0770 ;
        RECT 3.9880 83.9835 4.0140 85.0770 ;
        RECT 3.8800 83.9835 3.9060 85.0770 ;
        RECT 3.7720 83.9835 3.7980 85.0770 ;
        RECT 3.6640 83.9835 3.6900 85.0770 ;
        RECT 3.5560 83.9835 3.5820 85.0770 ;
        RECT 3.4480 83.9835 3.4740 85.0770 ;
        RECT 3.3400 83.9835 3.3660 85.0770 ;
        RECT 3.2320 83.9835 3.2580 85.0770 ;
        RECT 3.1240 83.9835 3.1500 85.0770 ;
        RECT 3.0160 83.9835 3.0420 85.0770 ;
        RECT 2.9080 83.9835 2.9340 85.0770 ;
        RECT 2.8000 83.9835 2.8260 85.0770 ;
        RECT 2.6920 83.9835 2.7180 85.0770 ;
        RECT 2.5840 83.9835 2.6100 85.0770 ;
        RECT 2.4760 83.9835 2.5020 85.0770 ;
        RECT 2.3680 83.9835 2.3940 85.0770 ;
        RECT 2.2600 83.9835 2.2860 85.0770 ;
        RECT 2.1520 83.9835 2.1780 85.0770 ;
        RECT 2.0440 83.9835 2.0700 85.0770 ;
        RECT 1.9360 83.9835 1.9620 85.0770 ;
        RECT 1.8280 83.9835 1.8540 85.0770 ;
        RECT 1.7200 83.9835 1.7460 85.0770 ;
        RECT 1.6120 83.9835 1.6380 85.0770 ;
        RECT 1.5040 83.9835 1.5300 85.0770 ;
        RECT 1.3960 83.9835 1.4220 85.0770 ;
        RECT 1.2880 83.9835 1.3140 85.0770 ;
        RECT 1.1800 83.9835 1.2060 85.0770 ;
        RECT 1.0720 83.9835 1.0980 85.0770 ;
        RECT 0.9640 83.9835 0.9900 85.0770 ;
        RECT 0.8560 83.9835 0.8820 85.0770 ;
        RECT 0.7480 83.9835 0.7740 85.0770 ;
        RECT 0.6400 83.9835 0.6660 85.0770 ;
        RECT 0.5320 83.9835 0.5580 85.0770 ;
        RECT 0.4240 83.9835 0.4500 85.0770 ;
        RECT 0.3160 83.9835 0.3420 85.0770 ;
        RECT 0.2080 83.9835 0.2340 85.0770 ;
        RECT 0.0050 83.9835 0.0900 85.0770 ;
        RECT 8.6410 85.0635 8.7690 86.1570 ;
        RECT 8.6270 85.7290 8.7690 86.0515 ;
        RECT 8.4790 85.4560 8.5410 86.1570 ;
        RECT 8.4650 85.7655 8.5410 85.9190 ;
        RECT 8.4790 85.0635 8.5050 86.1570 ;
        RECT 8.4790 85.1845 8.5190 85.4240 ;
        RECT 8.4790 85.0635 8.5410 85.1525 ;
        RECT 8.1820 85.5140 8.3880 86.1570 ;
        RECT 8.3620 85.0635 8.3880 86.1570 ;
        RECT 8.1820 85.7910 8.4020 86.0490 ;
        RECT 8.1820 85.0635 8.2800 86.1570 ;
        RECT 7.7650 85.0635 7.8480 86.1570 ;
        RECT 7.7650 85.1520 7.8620 86.0875 ;
        RECT 16.4440 85.0635 16.5290 86.1570 ;
        RECT 16.3000 85.0635 16.3260 86.1570 ;
        RECT 16.1920 85.0635 16.2180 86.1570 ;
        RECT 16.0840 85.0635 16.1100 86.1570 ;
        RECT 15.9760 85.0635 16.0020 86.1570 ;
        RECT 15.8680 85.0635 15.8940 86.1570 ;
        RECT 15.7600 85.0635 15.7860 86.1570 ;
        RECT 15.6520 85.0635 15.6780 86.1570 ;
        RECT 15.5440 85.0635 15.5700 86.1570 ;
        RECT 15.4360 85.0635 15.4620 86.1570 ;
        RECT 15.3280 85.0635 15.3540 86.1570 ;
        RECT 15.2200 85.0635 15.2460 86.1570 ;
        RECT 15.1120 85.0635 15.1380 86.1570 ;
        RECT 15.0040 85.0635 15.0300 86.1570 ;
        RECT 14.8960 85.0635 14.9220 86.1570 ;
        RECT 14.7880 85.0635 14.8140 86.1570 ;
        RECT 14.6800 85.0635 14.7060 86.1570 ;
        RECT 14.5720 85.0635 14.5980 86.1570 ;
        RECT 14.4640 85.0635 14.4900 86.1570 ;
        RECT 14.3560 85.0635 14.3820 86.1570 ;
        RECT 14.2480 85.0635 14.2740 86.1570 ;
        RECT 14.1400 85.0635 14.1660 86.1570 ;
        RECT 14.0320 85.0635 14.0580 86.1570 ;
        RECT 13.9240 85.0635 13.9500 86.1570 ;
        RECT 13.8160 85.0635 13.8420 86.1570 ;
        RECT 13.7080 85.0635 13.7340 86.1570 ;
        RECT 13.6000 85.0635 13.6260 86.1570 ;
        RECT 13.4920 85.0635 13.5180 86.1570 ;
        RECT 13.3840 85.0635 13.4100 86.1570 ;
        RECT 13.2760 85.0635 13.3020 86.1570 ;
        RECT 13.1680 85.0635 13.1940 86.1570 ;
        RECT 13.0600 85.0635 13.0860 86.1570 ;
        RECT 12.9520 85.0635 12.9780 86.1570 ;
        RECT 12.8440 85.0635 12.8700 86.1570 ;
        RECT 12.7360 85.0635 12.7620 86.1570 ;
        RECT 12.6280 85.0635 12.6540 86.1570 ;
        RECT 12.5200 85.0635 12.5460 86.1570 ;
        RECT 12.4120 85.0635 12.4380 86.1570 ;
        RECT 12.3040 85.0635 12.3300 86.1570 ;
        RECT 12.1960 85.0635 12.2220 86.1570 ;
        RECT 12.0880 85.0635 12.1140 86.1570 ;
        RECT 11.9800 85.0635 12.0060 86.1570 ;
        RECT 11.8720 85.0635 11.8980 86.1570 ;
        RECT 11.7640 85.0635 11.7900 86.1570 ;
        RECT 11.6560 85.0635 11.6820 86.1570 ;
        RECT 11.5480 85.0635 11.5740 86.1570 ;
        RECT 11.4400 85.0635 11.4660 86.1570 ;
        RECT 11.3320 85.0635 11.3580 86.1570 ;
        RECT 11.2240 85.0635 11.2500 86.1570 ;
        RECT 11.1160 85.0635 11.1420 86.1570 ;
        RECT 11.0080 85.0635 11.0340 86.1570 ;
        RECT 10.9000 85.0635 10.9260 86.1570 ;
        RECT 10.7920 85.0635 10.8180 86.1570 ;
        RECT 10.6840 85.0635 10.7100 86.1570 ;
        RECT 10.5760 85.0635 10.6020 86.1570 ;
        RECT 10.4680 85.0635 10.4940 86.1570 ;
        RECT 10.3600 85.0635 10.3860 86.1570 ;
        RECT 10.2520 85.0635 10.2780 86.1570 ;
        RECT 10.1440 85.0635 10.1700 86.1570 ;
        RECT 10.0360 85.0635 10.0620 86.1570 ;
        RECT 9.9280 85.0635 9.9540 86.1570 ;
        RECT 9.8200 85.0635 9.8460 86.1570 ;
        RECT 9.7120 85.0635 9.7380 86.1570 ;
        RECT 9.6040 85.0635 9.6300 86.1570 ;
        RECT 9.4960 85.0635 9.5220 86.1570 ;
        RECT 9.3880 85.0635 9.4140 86.1570 ;
        RECT 9.1750 85.0635 9.2520 86.1570 ;
        RECT 7.2820 85.0635 7.3590 86.1570 ;
        RECT 7.1200 85.0635 7.1460 86.1570 ;
        RECT 7.0120 85.0635 7.0380 86.1570 ;
        RECT 6.9040 85.0635 6.9300 86.1570 ;
        RECT 6.7960 85.0635 6.8220 86.1570 ;
        RECT 6.6880 85.0635 6.7140 86.1570 ;
        RECT 6.5800 85.0635 6.6060 86.1570 ;
        RECT 6.4720 85.0635 6.4980 86.1570 ;
        RECT 6.3640 85.0635 6.3900 86.1570 ;
        RECT 6.2560 85.0635 6.2820 86.1570 ;
        RECT 6.1480 85.0635 6.1740 86.1570 ;
        RECT 6.0400 85.0635 6.0660 86.1570 ;
        RECT 5.9320 85.0635 5.9580 86.1570 ;
        RECT 5.8240 85.0635 5.8500 86.1570 ;
        RECT 5.7160 85.0635 5.7420 86.1570 ;
        RECT 5.6080 85.0635 5.6340 86.1570 ;
        RECT 5.5000 85.0635 5.5260 86.1570 ;
        RECT 5.3920 85.0635 5.4180 86.1570 ;
        RECT 5.2840 85.0635 5.3100 86.1570 ;
        RECT 5.1760 85.0635 5.2020 86.1570 ;
        RECT 5.0680 85.0635 5.0940 86.1570 ;
        RECT 4.9600 85.0635 4.9860 86.1570 ;
        RECT 4.8520 85.0635 4.8780 86.1570 ;
        RECT 4.7440 85.0635 4.7700 86.1570 ;
        RECT 4.6360 85.0635 4.6620 86.1570 ;
        RECT 4.5280 85.0635 4.5540 86.1570 ;
        RECT 4.4200 85.0635 4.4460 86.1570 ;
        RECT 4.3120 85.0635 4.3380 86.1570 ;
        RECT 4.2040 85.0635 4.2300 86.1570 ;
        RECT 4.0960 85.0635 4.1220 86.1570 ;
        RECT 3.9880 85.0635 4.0140 86.1570 ;
        RECT 3.8800 85.0635 3.9060 86.1570 ;
        RECT 3.7720 85.0635 3.7980 86.1570 ;
        RECT 3.6640 85.0635 3.6900 86.1570 ;
        RECT 3.5560 85.0635 3.5820 86.1570 ;
        RECT 3.4480 85.0635 3.4740 86.1570 ;
        RECT 3.3400 85.0635 3.3660 86.1570 ;
        RECT 3.2320 85.0635 3.2580 86.1570 ;
        RECT 3.1240 85.0635 3.1500 86.1570 ;
        RECT 3.0160 85.0635 3.0420 86.1570 ;
        RECT 2.9080 85.0635 2.9340 86.1570 ;
        RECT 2.8000 85.0635 2.8260 86.1570 ;
        RECT 2.6920 85.0635 2.7180 86.1570 ;
        RECT 2.5840 85.0635 2.6100 86.1570 ;
        RECT 2.4760 85.0635 2.5020 86.1570 ;
        RECT 2.3680 85.0635 2.3940 86.1570 ;
        RECT 2.2600 85.0635 2.2860 86.1570 ;
        RECT 2.1520 85.0635 2.1780 86.1570 ;
        RECT 2.0440 85.0635 2.0700 86.1570 ;
        RECT 1.9360 85.0635 1.9620 86.1570 ;
        RECT 1.8280 85.0635 1.8540 86.1570 ;
        RECT 1.7200 85.0635 1.7460 86.1570 ;
        RECT 1.6120 85.0635 1.6380 86.1570 ;
        RECT 1.5040 85.0635 1.5300 86.1570 ;
        RECT 1.3960 85.0635 1.4220 86.1570 ;
        RECT 1.2880 85.0635 1.3140 86.1570 ;
        RECT 1.1800 85.0635 1.2060 86.1570 ;
        RECT 1.0720 85.0635 1.0980 86.1570 ;
        RECT 0.9640 85.0635 0.9900 86.1570 ;
        RECT 0.8560 85.0635 0.8820 86.1570 ;
        RECT 0.7480 85.0635 0.7740 86.1570 ;
        RECT 0.6400 85.0635 0.6660 86.1570 ;
        RECT 0.5320 85.0635 0.5580 86.1570 ;
        RECT 0.4240 85.0635 0.4500 86.1570 ;
        RECT 0.3160 85.0635 0.3420 86.1570 ;
        RECT 0.2080 85.0635 0.2340 86.1570 ;
        RECT 0.0050 85.0635 0.0900 86.1570 ;
        RECT 8.6410 86.1435 8.7690 87.2370 ;
        RECT 8.6270 86.8090 8.7690 87.1315 ;
        RECT 8.4790 86.5360 8.5410 87.2370 ;
        RECT 8.4650 86.8455 8.5410 86.9990 ;
        RECT 8.4790 86.1435 8.5050 87.2370 ;
        RECT 8.4790 86.2645 8.5190 86.5040 ;
        RECT 8.4790 86.1435 8.5410 86.2325 ;
        RECT 8.1820 86.5940 8.3880 87.2370 ;
        RECT 8.3620 86.1435 8.3880 87.2370 ;
        RECT 8.1820 86.8710 8.4020 87.1290 ;
        RECT 8.1820 86.1435 8.2800 87.2370 ;
        RECT 7.7650 86.1435 7.8480 87.2370 ;
        RECT 7.7650 86.2320 7.8620 87.1675 ;
        RECT 16.4440 86.1435 16.5290 87.2370 ;
        RECT 16.3000 86.1435 16.3260 87.2370 ;
        RECT 16.1920 86.1435 16.2180 87.2370 ;
        RECT 16.0840 86.1435 16.1100 87.2370 ;
        RECT 15.9760 86.1435 16.0020 87.2370 ;
        RECT 15.8680 86.1435 15.8940 87.2370 ;
        RECT 15.7600 86.1435 15.7860 87.2370 ;
        RECT 15.6520 86.1435 15.6780 87.2370 ;
        RECT 15.5440 86.1435 15.5700 87.2370 ;
        RECT 15.4360 86.1435 15.4620 87.2370 ;
        RECT 15.3280 86.1435 15.3540 87.2370 ;
        RECT 15.2200 86.1435 15.2460 87.2370 ;
        RECT 15.1120 86.1435 15.1380 87.2370 ;
        RECT 15.0040 86.1435 15.0300 87.2370 ;
        RECT 14.8960 86.1435 14.9220 87.2370 ;
        RECT 14.7880 86.1435 14.8140 87.2370 ;
        RECT 14.6800 86.1435 14.7060 87.2370 ;
        RECT 14.5720 86.1435 14.5980 87.2370 ;
        RECT 14.4640 86.1435 14.4900 87.2370 ;
        RECT 14.3560 86.1435 14.3820 87.2370 ;
        RECT 14.2480 86.1435 14.2740 87.2370 ;
        RECT 14.1400 86.1435 14.1660 87.2370 ;
        RECT 14.0320 86.1435 14.0580 87.2370 ;
        RECT 13.9240 86.1435 13.9500 87.2370 ;
        RECT 13.8160 86.1435 13.8420 87.2370 ;
        RECT 13.7080 86.1435 13.7340 87.2370 ;
        RECT 13.6000 86.1435 13.6260 87.2370 ;
        RECT 13.4920 86.1435 13.5180 87.2370 ;
        RECT 13.3840 86.1435 13.4100 87.2370 ;
        RECT 13.2760 86.1435 13.3020 87.2370 ;
        RECT 13.1680 86.1435 13.1940 87.2370 ;
        RECT 13.0600 86.1435 13.0860 87.2370 ;
        RECT 12.9520 86.1435 12.9780 87.2370 ;
        RECT 12.8440 86.1435 12.8700 87.2370 ;
        RECT 12.7360 86.1435 12.7620 87.2370 ;
        RECT 12.6280 86.1435 12.6540 87.2370 ;
        RECT 12.5200 86.1435 12.5460 87.2370 ;
        RECT 12.4120 86.1435 12.4380 87.2370 ;
        RECT 12.3040 86.1435 12.3300 87.2370 ;
        RECT 12.1960 86.1435 12.2220 87.2370 ;
        RECT 12.0880 86.1435 12.1140 87.2370 ;
        RECT 11.9800 86.1435 12.0060 87.2370 ;
        RECT 11.8720 86.1435 11.8980 87.2370 ;
        RECT 11.7640 86.1435 11.7900 87.2370 ;
        RECT 11.6560 86.1435 11.6820 87.2370 ;
        RECT 11.5480 86.1435 11.5740 87.2370 ;
        RECT 11.4400 86.1435 11.4660 87.2370 ;
        RECT 11.3320 86.1435 11.3580 87.2370 ;
        RECT 11.2240 86.1435 11.2500 87.2370 ;
        RECT 11.1160 86.1435 11.1420 87.2370 ;
        RECT 11.0080 86.1435 11.0340 87.2370 ;
        RECT 10.9000 86.1435 10.9260 87.2370 ;
        RECT 10.7920 86.1435 10.8180 87.2370 ;
        RECT 10.6840 86.1435 10.7100 87.2370 ;
        RECT 10.5760 86.1435 10.6020 87.2370 ;
        RECT 10.4680 86.1435 10.4940 87.2370 ;
        RECT 10.3600 86.1435 10.3860 87.2370 ;
        RECT 10.2520 86.1435 10.2780 87.2370 ;
        RECT 10.1440 86.1435 10.1700 87.2370 ;
        RECT 10.0360 86.1435 10.0620 87.2370 ;
        RECT 9.9280 86.1435 9.9540 87.2370 ;
        RECT 9.8200 86.1435 9.8460 87.2370 ;
        RECT 9.7120 86.1435 9.7380 87.2370 ;
        RECT 9.6040 86.1435 9.6300 87.2370 ;
        RECT 9.4960 86.1435 9.5220 87.2370 ;
        RECT 9.3880 86.1435 9.4140 87.2370 ;
        RECT 9.1750 86.1435 9.2520 87.2370 ;
        RECT 7.2820 86.1435 7.3590 87.2370 ;
        RECT 7.1200 86.1435 7.1460 87.2370 ;
        RECT 7.0120 86.1435 7.0380 87.2370 ;
        RECT 6.9040 86.1435 6.9300 87.2370 ;
        RECT 6.7960 86.1435 6.8220 87.2370 ;
        RECT 6.6880 86.1435 6.7140 87.2370 ;
        RECT 6.5800 86.1435 6.6060 87.2370 ;
        RECT 6.4720 86.1435 6.4980 87.2370 ;
        RECT 6.3640 86.1435 6.3900 87.2370 ;
        RECT 6.2560 86.1435 6.2820 87.2370 ;
        RECT 6.1480 86.1435 6.1740 87.2370 ;
        RECT 6.0400 86.1435 6.0660 87.2370 ;
        RECT 5.9320 86.1435 5.9580 87.2370 ;
        RECT 5.8240 86.1435 5.8500 87.2370 ;
        RECT 5.7160 86.1435 5.7420 87.2370 ;
        RECT 5.6080 86.1435 5.6340 87.2370 ;
        RECT 5.5000 86.1435 5.5260 87.2370 ;
        RECT 5.3920 86.1435 5.4180 87.2370 ;
        RECT 5.2840 86.1435 5.3100 87.2370 ;
        RECT 5.1760 86.1435 5.2020 87.2370 ;
        RECT 5.0680 86.1435 5.0940 87.2370 ;
        RECT 4.9600 86.1435 4.9860 87.2370 ;
        RECT 4.8520 86.1435 4.8780 87.2370 ;
        RECT 4.7440 86.1435 4.7700 87.2370 ;
        RECT 4.6360 86.1435 4.6620 87.2370 ;
        RECT 4.5280 86.1435 4.5540 87.2370 ;
        RECT 4.4200 86.1435 4.4460 87.2370 ;
        RECT 4.3120 86.1435 4.3380 87.2370 ;
        RECT 4.2040 86.1435 4.2300 87.2370 ;
        RECT 4.0960 86.1435 4.1220 87.2370 ;
        RECT 3.9880 86.1435 4.0140 87.2370 ;
        RECT 3.8800 86.1435 3.9060 87.2370 ;
        RECT 3.7720 86.1435 3.7980 87.2370 ;
        RECT 3.6640 86.1435 3.6900 87.2370 ;
        RECT 3.5560 86.1435 3.5820 87.2370 ;
        RECT 3.4480 86.1435 3.4740 87.2370 ;
        RECT 3.3400 86.1435 3.3660 87.2370 ;
        RECT 3.2320 86.1435 3.2580 87.2370 ;
        RECT 3.1240 86.1435 3.1500 87.2370 ;
        RECT 3.0160 86.1435 3.0420 87.2370 ;
        RECT 2.9080 86.1435 2.9340 87.2370 ;
        RECT 2.8000 86.1435 2.8260 87.2370 ;
        RECT 2.6920 86.1435 2.7180 87.2370 ;
        RECT 2.5840 86.1435 2.6100 87.2370 ;
        RECT 2.4760 86.1435 2.5020 87.2370 ;
        RECT 2.3680 86.1435 2.3940 87.2370 ;
        RECT 2.2600 86.1435 2.2860 87.2370 ;
        RECT 2.1520 86.1435 2.1780 87.2370 ;
        RECT 2.0440 86.1435 2.0700 87.2370 ;
        RECT 1.9360 86.1435 1.9620 87.2370 ;
        RECT 1.8280 86.1435 1.8540 87.2370 ;
        RECT 1.7200 86.1435 1.7460 87.2370 ;
        RECT 1.6120 86.1435 1.6380 87.2370 ;
        RECT 1.5040 86.1435 1.5300 87.2370 ;
        RECT 1.3960 86.1435 1.4220 87.2370 ;
        RECT 1.2880 86.1435 1.3140 87.2370 ;
        RECT 1.1800 86.1435 1.2060 87.2370 ;
        RECT 1.0720 86.1435 1.0980 87.2370 ;
        RECT 0.9640 86.1435 0.9900 87.2370 ;
        RECT 0.8560 86.1435 0.8820 87.2370 ;
        RECT 0.7480 86.1435 0.7740 87.2370 ;
        RECT 0.6400 86.1435 0.6660 87.2370 ;
        RECT 0.5320 86.1435 0.5580 87.2370 ;
        RECT 0.4240 86.1435 0.4500 87.2370 ;
        RECT 0.3160 86.1435 0.3420 87.2370 ;
        RECT 0.2080 86.1435 0.2340 87.2370 ;
        RECT 0.0050 86.1435 0.0900 87.2370 ;
        RECT 8.6410 87.2235 8.7690 88.3170 ;
        RECT 8.6270 87.8890 8.7690 88.2115 ;
        RECT 8.4790 87.6160 8.5410 88.3170 ;
        RECT 8.4650 87.9255 8.5410 88.0790 ;
        RECT 8.4790 87.2235 8.5050 88.3170 ;
        RECT 8.4790 87.3445 8.5190 87.5840 ;
        RECT 8.4790 87.2235 8.5410 87.3125 ;
        RECT 8.1820 87.6740 8.3880 88.3170 ;
        RECT 8.3620 87.2235 8.3880 88.3170 ;
        RECT 8.1820 87.9510 8.4020 88.2090 ;
        RECT 8.1820 87.2235 8.2800 88.3170 ;
        RECT 7.7650 87.2235 7.8480 88.3170 ;
        RECT 7.7650 87.3120 7.8620 88.2475 ;
        RECT 16.4440 87.2235 16.5290 88.3170 ;
        RECT 16.3000 87.2235 16.3260 88.3170 ;
        RECT 16.1920 87.2235 16.2180 88.3170 ;
        RECT 16.0840 87.2235 16.1100 88.3170 ;
        RECT 15.9760 87.2235 16.0020 88.3170 ;
        RECT 15.8680 87.2235 15.8940 88.3170 ;
        RECT 15.7600 87.2235 15.7860 88.3170 ;
        RECT 15.6520 87.2235 15.6780 88.3170 ;
        RECT 15.5440 87.2235 15.5700 88.3170 ;
        RECT 15.4360 87.2235 15.4620 88.3170 ;
        RECT 15.3280 87.2235 15.3540 88.3170 ;
        RECT 15.2200 87.2235 15.2460 88.3170 ;
        RECT 15.1120 87.2235 15.1380 88.3170 ;
        RECT 15.0040 87.2235 15.0300 88.3170 ;
        RECT 14.8960 87.2235 14.9220 88.3170 ;
        RECT 14.7880 87.2235 14.8140 88.3170 ;
        RECT 14.6800 87.2235 14.7060 88.3170 ;
        RECT 14.5720 87.2235 14.5980 88.3170 ;
        RECT 14.4640 87.2235 14.4900 88.3170 ;
        RECT 14.3560 87.2235 14.3820 88.3170 ;
        RECT 14.2480 87.2235 14.2740 88.3170 ;
        RECT 14.1400 87.2235 14.1660 88.3170 ;
        RECT 14.0320 87.2235 14.0580 88.3170 ;
        RECT 13.9240 87.2235 13.9500 88.3170 ;
        RECT 13.8160 87.2235 13.8420 88.3170 ;
        RECT 13.7080 87.2235 13.7340 88.3170 ;
        RECT 13.6000 87.2235 13.6260 88.3170 ;
        RECT 13.4920 87.2235 13.5180 88.3170 ;
        RECT 13.3840 87.2235 13.4100 88.3170 ;
        RECT 13.2760 87.2235 13.3020 88.3170 ;
        RECT 13.1680 87.2235 13.1940 88.3170 ;
        RECT 13.0600 87.2235 13.0860 88.3170 ;
        RECT 12.9520 87.2235 12.9780 88.3170 ;
        RECT 12.8440 87.2235 12.8700 88.3170 ;
        RECT 12.7360 87.2235 12.7620 88.3170 ;
        RECT 12.6280 87.2235 12.6540 88.3170 ;
        RECT 12.5200 87.2235 12.5460 88.3170 ;
        RECT 12.4120 87.2235 12.4380 88.3170 ;
        RECT 12.3040 87.2235 12.3300 88.3170 ;
        RECT 12.1960 87.2235 12.2220 88.3170 ;
        RECT 12.0880 87.2235 12.1140 88.3170 ;
        RECT 11.9800 87.2235 12.0060 88.3170 ;
        RECT 11.8720 87.2235 11.8980 88.3170 ;
        RECT 11.7640 87.2235 11.7900 88.3170 ;
        RECT 11.6560 87.2235 11.6820 88.3170 ;
        RECT 11.5480 87.2235 11.5740 88.3170 ;
        RECT 11.4400 87.2235 11.4660 88.3170 ;
        RECT 11.3320 87.2235 11.3580 88.3170 ;
        RECT 11.2240 87.2235 11.2500 88.3170 ;
        RECT 11.1160 87.2235 11.1420 88.3170 ;
        RECT 11.0080 87.2235 11.0340 88.3170 ;
        RECT 10.9000 87.2235 10.9260 88.3170 ;
        RECT 10.7920 87.2235 10.8180 88.3170 ;
        RECT 10.6840 87.2235 10.7100 88.3170 ;
        RECT 10.5760 87.2235 10.6020 88.3170 ;
        RECT 10.4680 87.2235 10.4940 88.3170 ;
        RECT 10.3600 87.2235 10.3860 88.3170 ;
        RECT 10.2520 87.2235 10.2780 88.3170 ;
        RECT 10.1440 87.2235 10.1700 88.3170 ;
        RECT 10.0360 87.2235 10.0620 88.3170 ;
        RECT 9.9280 87.2235 9.9540 88.3170 ;
        RECT 9.8200 87.2235 9.8460 88.3170 ;
        RECT 9.7120 87.2235 9.7380 88.3170 ;
        RECT 9.6040 87.2235 9.6300 88.3170 ;
        RECT 9.4960 87.2235 9.5220 88.3170 ;
        RECT 9.3880 87.2235 9.4140 88.3170 ;
        RECT 9.1750 87.2235 9.2520 88.3170 ;
        RECT 7.2820 87.2235 7.3590 88.3170 ;
        RECT 7.1200 87.2235 7.1460 88.3170 ;
        RECT 7.0120 87.2235 7.0380 88.3170 ;
        RECT 6.9040 87.2235 6.9300 88.3170 ;
        RECT 6.7960 87.2235 6.8220 88.3170 ;
        RECT 6.6880 87.2235 6.7140 88.3170 ;
        RECT 6.5800 87.2235 6.6060 88.3170 ;
        RECT 6.4720 87.2235 6.4980 88.3170 ;
        RECT 6.3640 87.2235 6.3900 88.3170 ;
        RECT 6.2560 87.2235 6.2820 88.3170 ;
        RECT 6.1480 87.2235 6.1740 88.3170 ;
        RECT 6.0400 87.2235 6.0660 88.3170 ;
        RECT 5.9320 87.2235 5.9580 88.3170 ;
        RECT 5.8240 87.2235 5.8500 88.3170 ;
        RECT 5.7160 87.2235 5.7420 88.3170 ;
        RECT 5.6080 87.2235 5.6340 88.3170 ;
        RECT 5.5000 87.2235 5.5260 88.3170 ;
        RECT 5.3920 87.2235 5.4180 88.3170 ;
        RECT 5.2840 87.2235 5.3100 88.3170 ;
        RECT 5.1760 87.2235 5.2020 88.3170 ;
        RECT 5.0680 87.2235 5.0940 88.3170 ;
        RECT 4.9600 87.2235 4.9860 88.3170 ;
        RECT 4.8520 87.2235 4.8780 88.3170 ;
        RECT 4.7440 87.2235 4.7700 88.3170 ;
        RECT 4.6360 87.2235 4.6620 88.3170 ;
        RECT 4.5280 87.2235 4.5540 88.3170 ;
        RECT 4.4200 87.2235 4.4460 88.3170 ;
        RECT 4.3120 87.2235 4.3380 88.3170 ;
        RECT 4.2040 87.2235 4.2300 88.3170 ;
        RECT 4.0960 87.2235 4.1220 88.3170 ;
        RECT 3.9880 87.2235 4.0140 88.3170 ;
        RECT 3.8800 87.2235 3.9060 88.3170 ;
        RECT 3.7720 87.2235 3.7980 88.3170 ;
        RECT 3.6640 87.2235 3.6900 88.3170 ;
        RECT 3.5560 87.2235 3.5820 88.3170 ;
        RECT 3.4480 87.2235 3.4740 88.3170 ;
        RECT 3.3400 87.2235 3.3660 88.3170 ;
        RECT 3.2320 87.2235 3.2580 88.3170 ;
        RECT 3.1240 87.2235 3.1500 88.3170 ;
        RECT 3.0160 87.2235 3.0420 88.3170 ;
        RECT 2.9080 87.2235 2.9340 88.3170 ;
        RECT 2.8000 87.2235 2.8260 88.3170 ;
        RECT 2.6920 87.2235 2.7180 88.3170 ;
        RECT 2.5840 87.2235 2.6100 88.3170 ;
        RECT 2.4760 87.2235 2.5020 88.3170 ;
        RECT 2.3680 87.2235 2.3940 88.3170 ;
        RECT 2.2600 87.2235 2.2860 88.3170 ;
        RECT 2.1520 87.2235 2.1780 88.3170 ;
        RECT 2.0440 87.2235 2.0700 88.3170 ;
        RECT 1.9360 87.2235 1.9620 88.3170 ;
        RECT 1.8280 87.2235 1.8540 88.3170 ;
        RECT 1.7200 87.2235 1.7460 88.3170 ;
        RECT 1.6120 87.2235 1.6380 88.3170 ;
        RECT 1.5040 87.2235 1.5300 88.3170 ;
        RECT 1.3960 87.2235 1.4220 88.3170 ;
        RECT 1.2880 87.2235 1.3140 88.3170 ;
        RECT 1.1800 87.2235 1.2060 88.3170 ;
        RECT 1.0720 87.2235 1.0980 88.3170 ;
        RECT 0.9640 87.2235 0.9900 88.3170 ;
        RECT 0.8560 87.2235 0.8820 88.3170 ;
        RECT 0.7480 87.2235 0.7740 88.3170 ;
        RECT 0.6400 87.2235 0.6660 88.3170 ;
        RECT 0.5320 87.2235 0.5580 88.3170 ;
        RECT 0.4240 87.2235 0.4500 88.3170 ;
        RECT 0.3160 87.2235 0.3420 88.3170 ;
        RECT 0.2080 87.2235 0.2340 88.3170 ;
        RECT 0.0050 87.2235 0.0900 88.3170 ;
  LAYER V3 SPACING 0.018  ;
      RECT 0.0050 1.2200 16.5290 1.3500 ;
      RECT 16.4120 0.2565 16.5290 1.3500 ;
      RECT 9.3020 1.1240 16.3940 1.3500 ;
      RECT 7.9700 1.1240 9.2840 1.3500 ;
      RECT 7.2500 0.2565 7.8800 1.3500 ;
      RECT 0.1400 1.1240 7.2320 1.3500 ;
      RECT 0.0050 0.2565 0.1220 1.3500 ;
      RECT 16.3760 0.2565 16.5290 1.1720 ;
      RECT 9.3560 0.2565 16.3580 1.3500 ;
      RECT 8.6090 0.2565 9.3380 1.1720 ;
      RECT 8.4470 0.4520 8.5730 1.3500 ;
      RECT 7.1960 0.3560 8.4200 1.1720 ;
      RECT 0.1760 0.2565 7.1780 1.3500 ;
      RECT 0.0050 0.2565 0.1580 1.1720 ;
      RECT 8.5550 0.2565 16.5290 1.0760 ;
      RECT 0.0050 0.3560 8.5370 1.0760 ;
      RECT 8.3300 0.2565 16.5290 0.4280 ;
      RECT 0.0050 0.2565 8.3120 1.0760 ;
      RECT 0.0050 0.2565 16.5290 0.3320 ;
      RECT 0.0050 2.3000 16.5290 2.4300 ;
      RECT 16.4120 1.3365 16.5290 2.4300 ;
      RECT 9.3020 2.2040 16.3940 2.4300 ;
      RECT 7.9700 2.2040 9.2840 2.4300 ;
      RECT 7.2500 1.3365 7.8800 2.4300 ;
      RECT 0.1400 2.2040 7.2320 2.4300 ;
      RECT 0.0050 1.3365 0.1220 2.4300 ;
      RECT 16.3760 1.3365 16.5290 2.2520 ;
      RECT 9.3560 1.3365 16.3580 2.4300 ;
      RECT 8.6090 1.3365 9.3380 2.2520 ;
      RECT 8.4470 1.5320 8.5730 2.4300 ;
      RECT 7.1960 1.4360 8.4200 2.2520 ;
      RECT 0.1760 1.3365 7.1780 2.4300 ;
      RECT 0.0050 1.3365 0.1580 2.2520 ;
      RECT 8.5550 1.3365 16.5290 2.1560 ;
      RECT 0.0050 1.4360 8.5370 2.1560 ;
      RECT 8.3300 1.3365 16.5290 1.5080 ;
      RECT 0.0050 1.3365 8.3120 2.1560 ;
      RECT 0.0050 1.3365 16.5290 1.4120 ;
      RECT 0.0050 3.3800 16.5290 3.5100 ;
      RECT 16.4120 2.4165 16.5290 3.5100 ;
      RECT 9.3020 3.2840 16.3940 3.5100 ;
      RECT 7.9700 3.2840 9.2840 3.5100 ;
      RECT 7.2500 2.4165 7.8800 3.5100 ;
      RECT 0.1400 3.2840 7.2320 3.5100 ;
      RECT 0.0050 2.4165 0.1220 3.5100 ;
      RECT 16.3760 2.4165 16.5290 3.3320 ;
      RECT 9.3560 2.4165 16.3580 3.5100 ;
      RECT 8.6090 2.4165 9.3380 3.3320 ;
      RECT 8.4470 2.6120 8.5730 3.5100 ;
      RECT 7.1960 2.5160 8.4200 3.3320 ;
      RECT 0.1760 2.4165 7.1780 3.5100 ;
      RECT 0.0050 2.4165 0.1580 3.3320 ;
      RECT 8.5550 2.4165 16.5290 3.2360 ;
      RECT 0.0050 2.5160 8.5370 3.2360 ;
      RECT 8.3300 2.4165 16.5290 2.5880 ;
      RECT 0.0050 2.4165 8.3120 3.2360 ;
      RECT 0.0050 2.4165 16.5290 2.4920 ;
      RECT 0.0050 4.4600 16.5290 4.5900 ;
      RECT 16.4120 3.4965 16.5290 4.5900 ;
      RECT 9.3020 4.3640 16.3940 4.5900 ;
      RECT 7.9700 4.3640 9.2840 4.5900 ;
      RECT 7.2500 3.4965 7.8800 4.5900 ;
      RECT 0.1400 4.3640 7.2320 4.5900 ;
      RECT 0.0050 3.4965 0.1220 4.5900 ;
      RECT 16.3760 3.4965 16.5290 4.4120 ;
      RECT 9.3560 3.4965 16.3580 4.5900 ;
      RECT 8.6090 3.4965 9.3380 4.4120 ;
      RECT 8.4470 3.6920 8.5730 4.5900 ;
      RECT 7.1960 3.5960 8.4200 4.4120 ;
      RECT 0.1760 3.4965 7.1780 4.5900 ;
      RECT 0.0050 3.4965 0.1580 4.4120 ;
      RECT 8.5550 3.4965 16.5290 4.3160 ;
      RECT 0.0050 3.5960 8.5370 4.3160 ;
      RECT 8.3300 3.4965 16.5290 3.6680 ;
      RECT 0.0050 3.4965 8.3120 4.3160 ;
      RECT 0.0050 3.4965 16.5290 3.5720 ;
      RECT 0.0050 5.5400 16.5290 5.6700 ;
      RECT 16.4120 4.5765 16.5290 5.6700 ;
      RECT 9.3020 5.4440 16.3940 5.6700 ;
      RECT 7.9700 5.4440 9.2840 5.6700 ;
      RECT 7.2500 4.5765 7.8800 5.6700 ;
      RECT 0.1400 5.4440 7.2320 5.6700 ;
      RECT 0.0050 4.5765 0.1220 5.6700 ;
      RECT 16.3760 4.5765 16.5290 5.4920 ;
      RECT 9.3560 4.5765 16.3580 5.6700 ;
      RECT 8.6090 4.5765 9.3380 5.4920 ;
      RECT 8.4470 4.7720 8.5730 5.6700 ;
      RECT 7.1960 4.6760 8.4200 5.4920 ;
      RECT 0.1760 4.5765 7.1780 5.6700 ;
      RECT 0.0050 4.5765 0.1580 5.4920 ;
      RECT 8.5550 4.5765 16.5290 5.3960 ;
      RECT 0.0050 4.6760 8.5370 5.3960 ;
      RECT 8.3300 4.5765 16.5290 4.7480 ;
      RECT 0.0050 4.5765 8.3120 5.3960 ;
      RECT 0.0050 4.5765 16.5290 4.6520 ;
      RECT 0.0050 6.6200 16.5290 6.7500 ;
      RECT 16.4120 5.6565 16.5290 6.7500 ;
      RECT 9.3020 6.5240 16.3940 6.7500 ;
      RECT 7.9700 6.5240 9.2840 6.7500 ;
      RECT 7.2500 5.6565 7.8800 6.7500 ;
      RECT 0.1400 6.5240 7.2320 6.7500 ;
      RECT 0.0050 5.6565 0.1220 6.7500 ;
      RECT 16.3760 5.6565 16.5290 6.5720 ;
      RECT 9.3560 5.6565 16.3580 6.7500 ;
      RECT 8.6090 5.6565 9.3380 6.5720 ;
      RECT 8.4470 5.8520 8.5730 6.7500 ;
      RECT 7.1960 5.7560 8.4200 6.5720 ;
      RECT 0.1760 5.6565 7.1780 6.7500 ;
      RECT 0.0050 5.6565 0.1580 6.5720 ;
      RECT 8.5550 5.6565 16.5290 6.4760 ;
      RECT 0.0050 5.7560 8.5370 6.4760 ;
      RECT 8.3300 5.6565 16.5290 5.8280 ;
      RECT 0.0050 5.6565 8.3120 6.4760 ;
      RECT 0.0050 5.6565 16.5290 5.7320 ;
      RECT 0.0050 7.7000 16.5290 7.8300 ;
      RECT 16.4120 6.7365 16.5290 7.8300 ;
      RECT 9.3020 7.6040 16.3940 7.8300 ;
      RECT 7.9700 7.6040 9.2840 7.8300 ;
      RECT 7.2500 6.7365 7.8800 7.8300 ;
      RECT 0.1400 7.6040 7.2320 7.8300 ;
      RECT 0.0050 6.7365 0.1220 7.8300 ;
      RECT 16.3760 6.7365 16.5290 7.6520 ;
      RECT 9.3560 6.7365 16.3580 7.8300 ;
      RECT 8.6090 6.7365 9.3380 7.6520 ;
      RECT 8.4470 6.9320 8.5730 7.8300 ;
      RECT 7.1960 6.8360 8.4200 7.6520 ;
      RECT 0.1760 6.7365 7.1780 7.8300 ;
      RECT 0.0050 6.7365 0.1580 7.6520 ;
      RECT 8.5550 6.7365 16.5290 7.5560 ;
      RECT 0.0050 6.8360 8.5370 7.5560 ;
      RECT 8.3300 6.7365 16.5290 6.9080 ;
      RECT 0.0050 6.7365 8.3120 7.5560 ;
      RECT 0.0050 6.7365 16.5290 6.8120 ;
      RECT 0.0050 8.7800 16.5290 8.9100 ;
      RECT 16.4120 7.8165 16.5290 8.9100 ;
      RECT 9.3020 8.6840 16.3940 8.9100 ;
      RECT 7.9700 8.6840 9.2840 8.9100 ;
      RECT 7.2500 7.8165 7.8800 8.9100 ;
      RECT 0.1400 8.6840 7.2320 8.9100 ;
      RECT 0.0050 7.8165 0.1220 8.9100 ;
      RECT 16.3760 7.8165 16.5290 8.7320 ;
      RECT 9.3560 7.8165 16.3580 8.9100 ;
      RECT 8.6090 7.8165 9.3380 8.7320 ;
      RECT 8.4470 8.0120 8.5730 8.9100 ;
      RECT 7.1960 7.9160 8.4200 8.7320 ;
      RECT 0.1760 7.8165 7.1780 8.9100 ;
      RECT 0.0050 7.8165 0.1580 8.7320 ;
      RECT 8.5550 7.8165 16.5290 8.6360 ;
      RECT 0.0050 7.9160 8.5370 8.6360 ;
      RECT 8.3300 7.8165 16.5290 7.9880 ;
      RECT 0.0050 7.8165 8.3120 8.6360 ;
      RECT 0.0050 7.8165 16.5290 7.8920 ;
      RECT 0.0050 9.8600 16.5290 9.9900 ;
      RECT 16.4120 8.8965 16.5290 9.9900 ;
      RECT 9.3020 9.7640 16.3940 9.9900 ;
      RECT 7.9700 9.7640 9.2840 9.9900 ;
      RECT 7.2500 8.8965 7.8800 9.9900 ;
      RECT 0.1400 9.7640 7.2320 9.9900 ;
      RECT 0.0050 8.8965 0.1220 9.9900 ;
      RECT 16.3760 8.8965 16.5290 9.8120 ;
      RECT 9.3560 8.8965 16.3580 9.9900 ;
      RECT 8.6090 8.8965 9.3380 9.8120 ;
      RECT 8.4470 9.0920 8.5730 9.9900 ;
      RECT 7.1960 8.9960 8.4200 9.8120 ;
      RECT 0.1760 8.8965 7.1780 9.9900 ;
      RECT 0.0050 8.8965 0.1580 9.8120 ;
      RECT 8.5550 8.8965 16.5290 9.7160 ;
      RECT 0.0050 8.9960 8.5370 9.7160 ;
      RECT 8.3300 8.8965 16.5290 9.0680 ;
      RECT 0.0050 8.8965 8.3120 9.7160 ;
      RECT 0.0050 8.8965 16.5290 8.9720 ;
      RECT 0.0050 10.9400 16.5290 11.0700 ;
      RECT 16.4120 9.9765 16.5290 11.0700 ;
      RECT 9.3020 10.8440 16.3940 11.0700 ;
      RECT 7.9700 10.8440 9.2840 11.0700 ;
      RECT 7.2500 9.9765 7.8800 11.0700 ;
      RECT 0.1400 10.8440 7.2320 11.0700 ;
      RECT 0.0050 9.9765 0.1220 11.0700 ;
      RECT 16.3760 9.9765 16.5290 10.8920 ;
      RECT 9.3560 9.9765 16.3580 11.0700 ;
      RECT 8.6090 9.9765 9.3380 10.8920 ;
      RECT 8.4470 10.1720 8.5730 11.0700 ;
      RECT 7.1960 10.0760 8.4200 10.8920 ;
      RECT 0.1760 9.9765 7.1780 11.0700 ;
      RECT 0.0050 9.9765 0.1580 10.8920 ;
      RECT 8.5550 9.9765 16.5290 10.7960 ;
      RECT 0.0050 10.0760 8.5370 10.7960 ;
      RECT 8.3300 9.9765 16.5290 10.1480 ;
      RECT 0.0050 9.9765 8.3120 10.7960 ;
      RECT 0.0050 9.9765 16.5290 10.0520 ;
      RECT 0.0050 12.0200 16.5290 12.1500 ;
      RECT 16.4120 11.0565 16.5290 12.1500 ;
      RECT 9.3020 11.9240 16.3940 12.1500 ;
      RECT 7.9700 11.9240 9.2840 12.1500 ;
      RECT 7.2500 11.0565 7.8800 12.1500 ;
      RECT 0.1400 11.9240 7.2320 12.1500 ;
      RECT 0.0050 11.0565 0.1220 12.1500 ;
      RECT 16.3760 11.0565 16.5290 11.9720 ;
      RECT 9.3560 11.0565 16.3580 12.1500 ;
      RECT 8.6090 11.0565 9.3380 11.9720 ;
      RECT 8.4470 11.2520 8.5730 12.1500 ;
      RECT 7.1960 11.1560 8.4200 11.9720 ;
      RECT 0.1760 11.0565 7.1780 12.1500 ;
      RECT 0.0050 11.0565 0.1580 11.9720 ;
      RECT 8.5550 11.0565 16.5290 11.8760 ;
      RECT 0.0050 11.1560 8.5370 11.8760 ;
      RECT 8.3300 11.0565 16.5290 11.2280 ;
      RECT 0.0050 11.0565 8.3120 11.8760 ;
      RECT 0.0050 11.0565 16.5290 11.1320 ;
      RECT 0.0050 13.1000 16.5290 13.2300 ;
      RECT 16.4120 12.1365 16.5290 13.2300 ;
      RECT 9.3020 13.0040 16.3940 13.2300 ;
      RECT 7.9700 13.0040 9.2840 13.2300 ;
      RECT 7.2500 12.1365 7.8800 13.2300 ;
      RECT 0.1400 13.0040 7.2320 13.2300 ;
      RECT 0.0050 12.1365 0.1220 13.2300 ;
      RECT 16.3760 12.1365 16.5290 13.0520 ;
      RECT 9.3560 12.1365 16.3580 13.2300 ;
      RECT 8.6090 12.1365 9.3380 13.0520 ;
      RECT 8.4470 12.3320 8.5730 13.2300 ;
      RECT 7.1960 12.2360 8.4200 13.0520 ;
      RECT 0.1760 12.1365 7.1780 13.2300 ;
      RECT 0.0050 12.1365 0.1580 13.0520 ;
      RECT 8.5550 12.1365 16.5290 12.9560 ;
      RECT 0.0050 12.2360 8.5370 12.9560 ;
      RECT 8.3300 12.1365 16.5290 12.3080 ;
      RECT 0.0050 12.1365 8.3120 12.9560 ;
      RECT 0.0050 12.1365 16.5290 12.2120 ;
      RECT 0.0050 14.1800 16.5290 14.3100 ;
      RECT 16.4120 13.2165 16.5290 14.3100 ;
      RECT 9.3020 14.0840 16.3940 14.3100 ;
      RECT 7.9700 14.0840 9.2840 14.3100 ;
      RECT 7.2500 13.2165 7.8800 14.3100 ;
      RECT 0.1400 14.0840 7.2320 14.3100 ;
      RECT 0.0050 13.2165 0.1220 14.3100 ;
      RECT 16.3760 13.2165 16.5290 14.1320 ;
      RECT 9.3560 13.2165 16.3580 14.3100 ;
      RECT 8.6090 13.2165 9.3380 14.1320 ;
      RECT 8.4470 13.4120 8.5730 14.3100 ;
      RECT 7.1960 13.3160 8.4200 14.1320 ;
      RECT 0.1760 13.2165 7.1780 14.3100 ;
      RECT 0.0050 13.2165 0.1580 14.1320 ;
      RECT 8.5550 13.2165 16.5290 14.0360 ;
      RECT 0.0050 13.3160 8.5370 14.0360 ;
      RECT 8.3300 13.2165 16.5290 13.3880 ;
      RECT 0.0050 13.2165 8.3120 14.0360 ;
      RECT 0.0050 13.2165 16.5290 13.2920 ;
      RECT 0.0050 15.2600 16.5290 15.3900 ;
      RECT 16.4120 14.2965 16.5290 15.3900 ;
      RECT 9.3020 15.1640 16.3940 15.3900 ;
      RECT 7.9700 15.1640 9.2840 15.3900 ;
      RECT 7.2500 14.2965 7.8800 15.3900 ;
      RECT 0.1400 15.1640 7.2320 15.3900 ;
      RECT 0.0050 14.2965 0.1220 15.3900 ;
      RECT 16.3760 14.2965 16.5290 15.2120 ;
      RECT 9.3560 14.2965 16.3580 15.3900 ;
      RECT 8.6090 14.2965 9.3380 15.2120 ;
      RECT 8.4470 14.4920 8.5730 15.3900 ;
      RECT 7.1960 14.3960 8.4200 15.2120 ;
      RECT 0.1760 14.2965 7.1780 15.3900 ;
      RECT 0.0050 14.2965 0.1580 15.2120 ;
      RECT 8.5550 14.2965 16.5290 15.1160 ;
      RECT 0.0050 14.3960 8.5370 15.1160 ;
      RECT 8.3300 14.2965 16.5290 14.4680 ;
      RECT 0.0050 14.2965 8.3120 15.1160 ;
      RECT 0.0050 14.2965 16.5290 14.3720 ;
      RECT 0.0050 16.3400 16.5290 16.4700 ;
      RECT 16.4120 15.3765 16.5290 16.4700 ;
      RECT 9.3020 16.2440 16.3940 16.4700 ;
      RECT 7.9700 16.2440 9.2840 16.4700 ;
      RECT 7.2500 15.3765 7.8800 16.4700 ;
      RECT 0.1400 16.2440 7.2320 16.4700 ;
      RECT 0.0050 15.3765 0.1220 16.4700 ;
      RECT 16.3760 15.3765 16.5290 16.2920 ;
      RECT 9.3560 15.3765 16.3580 16.4700 ;
      RECT 8.6090 15.3765 9.3380 16.2920 ;
      RECT 8.4470 15.5720 8.5730 16.4700 ;
      RECT 7.1960 15.4760 8.4200 16.2920 ;
      RECT 0.1760 15.3765 7.1780 16.4700 ;
      RECT 0.0050 15.3765 0.1580 16.2920 ;
      RECT 8.5550 15.3765 16.5290 16.1960 ;
      RECT 0.0050 15.4760 8.5370 16.1960 ;
      RECT 8.3300 15.3765 16.5290 15.5480 ;
      RECT 0.0050 15.3765 8.3120 16.1960 ;
      RECT 0.0050 15.3765 16.5290 15.4520 ;
      RECT 0.0050 17.4200 16.5290 17.5500 ;
      RECT 16.4120 16.4565 16.5290 17.5500 ;
      RECT 9.3020 17.3240 16.3940 17.5500 ;
      RECT 7.9700 17.3240 9.2840 17.5500 ;
      RECT 7.2500 16.4565 7.8800 17.5500 ;
      RECT 0.1400 17.3240 7.2320 17.5500 ;
      RECT 0.0050 16.4565 0.1220 17.5500 ;
      RECT 16.3760 16.4565 16.5290 17.3720 ;
      RECT 9.3560 16.4565 16.3580 17.5500 ;
      RECT 8.6090 16.4565 9.3380 17.3720 ;
      RECT 8.4470 16.6520 8.5730 17.5500 ;
      RECT 7.1960 16.5560 8.4200 17.3720 ;
      RECT 0.1760 16.4565 7.1780 17.5500 ;
      RECT 0.0050 16.4565 0.1580 17.3720 ;
      RECT 8.5550 16.4565 16.5290 17.2760 ;
      RECT 0.0050 16.5560 8.5370 17.2760 ;
      RECT 8.3300 16.4565 16.5290 16.6280 ;
      RECT 0.0050 16.4565 8.3120 17.2760 ;
      RECT 0.0050 16.4565 16.5290 16.5320 ;
      RECT 0.0050 18.5000 16.5290 18.6300 ;
      RECT 16.4120 17.5365 16.5290 18.6300 ;
      RECT 9.3020 18.4040 16.3940 18.6300 ;
      RECT 7.9700 18.4040 9.2840 18.6300 ;
      RECT 7.2500 17.5365 7.8800 18.6300 ;
      RECT 0.1400 18.4040 7.2320 18.6300 ;
      RECT 0.0050 17.5365 0.1220 18.6300 ;
      RECT 16.3760 17.5365 16.5290 18.4520 ;
      RECT 9.3560 17.5365 16.3580 18.6300 ;
      RECT 8.6090 17.5365 9.3380 18.4520 ;
      RECT 8.4470 17.7320 8.5730 18.6300 ;
      RECT 7.1960 17.6360 8.4200 18.4520 ;
      RECT 0.1760 17.5365 7.1780 18.6300 ;
      RECT 0.0050 17.5365 0.1580 18.4520 ;
      RECT 8.5550 17.5365 16.5290 18.3560 ;
      RECT 0.0050 17.6360 8.5370 18.3560 ;
      RECT 8.3300 17.5365 16.5290 17.7080 ;
      RECT 0.0050 17.5365 8.3120 18.3560 ;
      RECT 0.0050 17.5365 16.5290 17.6120 ;
      RECT 0.0050 19.5800 16.5290 19.7100 ;
      RECT 16.4120 18.6165 16.5290 19.7100 ;
      RECT 9.3020 19.4840 16.3940 19.7100 ;
      RECT 7.9700 19.4840 9.2840 19.7100 ;
      RECT 7.2500 18.6165 7.8800 19.7100 ;
      RECT 0.1400 19.4840 7.2320 19.7100 ;
      RECT 0.0050 18.6165 0.1220 19.7100 ;
      RECT 16.3760 18.6165 16.5290 19.5320 ;
      RECT 9.3560 18.6165 16.3580 19.7100 ;
      RECT 8.6090 18.6165 9.3380 19.5320 ;
      RECT 8.4470 18.8120 8.5730 19.7100 ;
      RECT 7.1960 18.7160 8.4200 19.5320 ;
      RECT 0.1760 18.6165 7.1780 19.7100 ;
      RECT 0.0050 18.6165 0.1580 19.5320 ;
      RECT 8.5550 18.6165 16.5290 19.4360 ;
      RECT 0.0050 18.7160 8.5370 19.4360 ;
      RECT 8.3300 18.6165 16.5290 18.7880 ;
      RECT 0.0050 18.6165 8.3120 19.4360 ;
      RECT 0.0050 18.6165 16.5290 18.6920 ;
      RECT 0.0050 20.6600 16.5290 20.7900 ;
      RECT 16.4120 19.6965 16.5290 20.7900 ;
      RECT 9.3020 20.5640 16.3940 20.7900 ;
      RECT 7.9700 20.5640 9.2840 20.7900 ;
      RECT 7.2500 19.6965 7.8800 20.7900 ;
      RECT 0.1400 20.5640 7.2320 20.7900 ;
      RECT 0.0050 19.6965 0.1220 20.7900 ;
      RECT 16.3760 19.6965 16.5290 20.6120 ;
      RECT 9.3560 19.6965 16.3580 20.7900 ;
      RECT 8.6090 19.6965 9.3380 20.6120 ;
      RECT 8.4470 19.8920 8.5730 20.7900 ;
      RECT 7.1960 19.7960 8.4200 20.6120 ;
      RECT 0.1760 19.6965 7.1780 20.7900 ;
      RECT 0.0050 19.6965 0.1580 20.6120 ;
      RECT 8.5550 19.6965 16.5290 20.5160 ;
      RECT 0.0050 19.7960 8.5370 20.5160 ;
      RECT 8.3300 19.6965 16.5290 19.8680 ;
      RECT 0.0050 19.6965 8.3120 20.5160 ;
      RECT 0.0050 19.6965 16.5290 19.7720 ;
      RECT 0.0050 21.7400 16.5290 21.8700 ;
      RECT 16.4120 20.7765 16.5290 21.8700 ;
      RECT 9.3020 21.6440 16.3940 21.8700 ;
      RECT 7.9700 21.6440 9.2840 21.8700 ;
      RECT 7.2500 20.7765 7.8800 21.8700 ;
      RECT 0.1400 21.6440 7.2320 21.8700 ;
      RECT 0.0050 20.7765 0.1220 21.8700 ;
      RECT 16.3760 20.7765 16.5290 21.6920 ;
      RECT 9.3560 20.7765 16.3580 21.8700 ;
      RECT 8.6090 20.7765 9.3380 21.6920 ;
      RECT 8.4470 20.9720 8.5730 21.8700 ;
      RECT 7.1960 20.8760 8.4200 21.6920 ;
      RECT 0.1760 20.7765 7.1780 21.8700 ;
      RECT 0.0050 20.7765 0.1580 21.6920 ;
      RECT 8.5550 20.7765 16.5290 21.5960 ;
      RECT 0.0050 20.8760 8.5370 21.5960 ;
      RECT 8.3300 20.7765 16.5290 20.9480 ;
      RECT 0.0050 20.7765 8.3120 21.5960 ;
      RECT 0.0050 20.7765 16.5290 20.8520 ;
      RECT 0.0050 22.8200 16.5290 22.9500 ;
      RECT 16.4120 21.8565 16.5290 22.9500 ;
      RECT 9.3020 22.7240 16.3940 22.9500 ;
      RECT 7.9700 22.7240 9.2840 22.9500 ;
      RECT 7.2500 21.8565 7.8800 22.9500 ;
      RECT 0.1400 22.7240 7.2320 22.9500 ;
      RECT 0.0050 21.8565 0.1220 22.9500 ;
      RECT 16.3760 21.8565 16.5290 22.7720 ;
      RECT 9.3560 21.8565 16.3580 22.9500 ;
      RECT 8.6090 21.8565 9.3380 22.7720 ;
      RECT 8.4470 22.0520 8.5730 22.9500 ;
      RECT 7.1960 21.9560 8.4200 22.7720 ;
      RECT 0.1760 21.8565 7.1780 22.9500 ;
      RECT 0.0050 21.8565 0.1580 22.7720 ;
      RECT 8.5550 21.8565 16.5290 22.6760 ;
      RECT 0.0050 21.9560 8.5370 22.6760 ;
      RECT 8.3300 21.8565 16.5290 22.0280 ;
      RECT 0.0050 21.8565 8.3120 22.6760 ;
      RECT 0.0050 21.8565 16.5290 21.9320 ;
      RECT 0.0050 23.9000 16.5290 24.0300 ;
      RECT 16.4120 22.9365 16.5290 24.0300 ;
      RECT 9.3020 23.8040 16.3940 24.0300 ;
      RECT 7.9700 23.8040 9.2840 24.0300 ;
      RECT 7.2500 22.9365 7.8800 24.0300 ;
      RECT 0.1400 23.8040 7.2320 24.0300 ;
      RECT 0.0050 22.9365 0.1220 24.0300 ;
      RECT 16.3760 22.9365 16.5290 23.8520 ;
      RECT 9.3560 22.9365 16.3580 24.0300 ;
      RECT 8.6090 22.9365 9.3380 23.8520 ;
      RECT 8.4470 23.1320 8.5730 24.0300 ;
      RECT 7.1960 23.0360 8.4200 23.8520 ;
      RECT 0.1760 22.9365 7.1780 24.0300 ;
      RECT 0.0050 22.9365 0.1580 23.8520 ;
      RECT 8.5550 22.9365 16.5290 23.7560 ;
      RECT 0.0050 23.0360 8.5370 23.7560 ;
      RECT 8.3300 22.9365 16.5290 23.1080 ;
      RECT 0.0050 22.9365 8.3120 23.7560 ;
      RECT 0.0050 22.9365 16.5290 23.0120 ;
      RECT 0.0050 24.9800 16.5290 25.1100 ;
      RECT 16.4120 24.0165 16.5290 25.1100 ;
      RECT 9.3020 24.8840 16.3940 25.1100 ;
      RECT 7.9700 24.8840 9.2840 25.1100 ;
      RECT 7.2500 24.0165 7.8800 25.1100 ;
      RECT 0.1400 24.8840 7.2320 25.1100 ;
      RECT 0.0050 24.0165 0.1220 25.1100 ;
      RECT 16.3760 24.0165 16.5290 24.9320 ;
      RECT 9.3560 24.0165 16.3580 25.1100 ;
      RECT 8.6090 24.0165 9.3380 24.9320 ;
      RECT 8.4470 24.2120 8.5730 25.1100 ;
      RECT 7.1960 24.1160 8.4200 24.9320 ;
      RECT 0.1760 24.0165 7.1780 25.1100 ;
      RECT 0.0050 24.0165 0.1580 24.9320 ;
      RECT 8.5550 24.0165 16.5290 24.8360 ;
      RECT 0.0050 24.1160 8.5370 24.8360 ;
      RECT 8.3300 24.0165 16.5290 24.1880 ;
      RECT 0.0050 24.0165 8.3120 24.8360 ;
      RECT 0.0050 24.0165 16.5290 24.0920 ;
      RECT 0.0050 26.0600 16.5290 26.1900 ;
      RECT 16.4120 25.0965 16.5290 26.1900 ;
      RECT 9.3020 25.9640 16.3940 26.1900 ;
      RECT 7.9700 25.9640 9.2840 26.1900 ;
      RECT 7.2500 25.0965 7.8800 26.1900 ;
      RECT 0.1400 25.9640 7.2320 26.1900 ;
      RECT 0.0050 25.0965 0.1220 26.1900 ;
      RECT 16.3760 25.0965 16.5290 26.0120 ;
      RECT 9.3560 25.0965 16.3580 26.1900 ;
      RECT 8.6090 25.0965 9.3380 26.0120 ;
      RECT 8.4470 25.2920 8.5730 26.1900 ;
      RECT 7.1960 25.1960 8.4200 26.0120 ;
      RECT 0.1760 25.0965 7.1780 26.1900 ;
      RECT 0.0050 25.0965 0.1580 26.0120 ;
      RECT 8.5550 25.0965 16.5290 25.9160 ;
      RECT 0.0050 25.1960 8.5370 25.9160 ;
      RECT 8.3300 25.0965 16.5290 25.2680 ;
      RECT 0.0050 25.0965 8.3120 25.9160 ;
      RECT 0.0050 25.0965 16.5290 25.1720 ;
      RECT 0.0050 27.1400 16.5290 27.2700 ;
      RECT 16.4120 26.1765 16.5290 27.2700 ;
      RECT 9.3020 27.0440 16.3940 27.2700 ;
      RECT 7.9700 27.0440 9.2840 27.2700 ;
      RECT 7.2500 26.1765 7.8800 27.2700 ;
      RECT 0.1400 27.0440 7.2320 27.2700 ;
      RECT 0.0050 26.1765 0.1220 27.2700 ;
      RECT 16.3760 26.1765 16.5290 27.0920 ;
      RECT 9.3560 26.1765 16.3580 27.2700 ;
      RECT 8.6090 26.1765 9.3380 27.0920 ;
      RECT 8.4470 26.3720 8.5730 27.2700 ;
      RECT 7.1960 26.2760 8.4200 27.0920 ;
      RECT 0.1760 26.1765 7.1780 27.2700 ;
      RECT 0.0050 26.1765 0.1580 27.0920 ;
      RECT 8.5550 26.1765 16.5290 26.9960 ;
      RECT 0.0050 26.2760 8.5370 26.9960 ;
      RECT 8.3300 26.1765 16.5290 26.3480 ;
      RECT 0.0050 26.1765 8.3120 26.9960 ;
      RECT 0.0050 26.1765 16.5290 26.2520 ;
      RECT 0.0050 28.2200 16.5290 28.3500 ;
      RECT 16.4120 27.2565 16.5290 28.3500 ;
      RECT 9.3020 28.1240 16.3940 28.3500 ;
      RECT 7.9700 28.1240 9.2840 28.3500 ;
      RECT 7.2500 27.2565 7.8800 28.3500 ;
      RECT 0.1400 28.1240 7.2320 28.3500 ;
      RECT 0.0050 27.2565 0.1220 28.3500 ;
      RECT 16.3760 27.2565 16.5290 28.1720 ;
      RECT 9.3560 27.2565 16.3580 28.3500 ;
      RECT 8.6090 27.2565 9.3380 28.1720 ;
      RECT 8.4470 27.4520 8.5730 28.3500 ;
      RECT 7.1960 27.3560 8.4200 28.1720 ;
      RECT 0.1760 27.2565 7.1780 28.3500 ;
      RECT 0.0050 27.2565 0.1580 28.1720 ;
      RECT 8.5550 27.2565 16.5290 28.0760 ;
      RECT 0.0050 27.3560 8.5370 28.0760 ;
      RECT 8.3300 27.2565 16.5290 27.4280 ;
      RECT 0.0050 27.2565 8.3120 28.0760 ;
      RECT 0.0050 27.2565 16.5290 27.3320 ;
      RECT 0.0050 29.3000 16.5290 29.4300 ;
      RECT 16.4120 28.3365 16.5290 29.4300 ;
      RECT 9.3020 29.2040 16.3940 29.4300 ;
      RECT 7.9700 29.2040 9.2840 29.4300 ;
      RECT 7.2500 28.3365 7.8800 29.4300 ;
      RECT 0.1400 29.2040 7.2320 29.4300 ;
      RECT 0.0050 28.3365 0.1220 29.4300 ;
      RECT 16.3760 28.3365 16.5290 29.2520 ;
      RECT 9.3560 28.3365 16.3580 29.4300 ;
      RECT 8.6090 28.3365 9.3380 29.2520 ;
      RECT 8.4470 28.5320 8.5730 29.4300 ;
      RECT 7.1960 28.4360 8.4200 29.2520 ;
      RECT 0.1760 28.3365 7.1780 29.4300 ;
      RECT 0.0050 28.3365 0.1580 29.2520 ;
      RECT 8.5550 28.3365 16.5290 29.1560 ;
      RECT 0.0050 28.4360 8.5370 29.1560 ;
      RECT 8.3300 28.3365 16.5290 28.5080 ;
      RECT 0.0050 28.3365 8.3120 29.1560 ;
      RECT 0.0050 28.3365 16.5290 28.4120 ;
      RECT 0.0050 30.3800 16.5290 30.5100 ;
      RECT 16.4120 29.4165 16.5290 30.5100 ;
      RECT 9.3020 30.2840 16.3940 30.5100 ;
      RECT 7.9700 30.2840 9.2840 30.5100 ;
      RECT 7.2500 29.4165 7.8800 30.5100 ;
      RECT 0.1400 30.2840 7.2320 30.5100 ;
      RECT 0.0050 29.4165 0.1220 30.5100 ;
      RECT 16.3760 29.4165 16.5290 30.3320 ;
      RECT 9.3560 29.4165 16.3580 30.5100 ;
      RECT 8.6090 29.4165 9.3380 30.3320 ;
      RECT 8.4470 29.6120 8.5730 30.5100 ;
      RECT 7.1960 29.5160 8.4200 30.3320 ;
      RECT 0.1760 29.4165 7.1780 30.5100 ;
      RECT 0.0050 29.4165 0.1580 30.3320 ;
      RECT 8.5550 29.4165 16.5290 30.2360 ;
      RECT 0.0050 29.5160 8.5370 30.2360 ;
      RECT 8.3300 29.4165 16.5290 29.5880 ;
      RECT 0.0050 29.4165 8.3120 30.2360 ;
      RECT 0.0050 29.4165 16.5290 29.4920 ;
      RECT 0.0050 31.4600 16.5290 31.5900 ;
      RECT 16.4120 30.4965 16.5290 31.5900 ;
      RECT 9.3020 31.3640 16.3940 31.5900 ;
      RECT 7.9700 31.3640 9.2840 31.5900 ;
      RECT 7.2500 30.4965 7.8800 31.5900 ;
      RECT 0.1400 31.3640 7.2320 31.5900 ;
      RECT 0.0050 30.4965 0.1220 31.5900 ;
      RECT 16.3760 30.4965 16.5290 31.4120 ;
      RECT 9.3560 30.4965 16.3580 31.5900 ;
      RECT 8.6090 30.4965 9.3380 31.4120 ;
      RECT 8.4470 30.6920 8.5730 31.5900 ;
      RECT 7.1960 30.5960 8.4200 31.4120 ;
      RECT 0.1760 30.4965 7.1780 31.5900 ;
      RECT 0.0050 30.4965 0.1580 31.4120 ;
      RECT 8.5550 30.4965 16.5290 31.3160 ;
      RECT 0.0050 30.5960 8.5370 31.3160 ;
      RECT 8.3300 30.4965 16.5290 30.6680 ;
      RECT 0.0050 30.4965 8.3120 31.3160 ;
      RECT 0.0050 30.4965 16.5290 30.5720 ;
      RECT 0.0050 32.5400 16.5290 32.6700 ;
      RECT 16.4120 31.5765 16.5290 32.6700 ;
      RECT 9.3020 32.4440 16.3940 32.6700 ;
      RECT 7.9700 32.4440 9.2840 32.6700 ;
      RECT 7.2500 31.5765 7.8800 32.6700 ;
      RECT 0.1400 32.4440 7.2320 32.6700 ;
      RECT 0.0050 31.5765 0.1220 32.6700 ;
      RECT 16.3760 31.5765 16.5290 32.4920 ;
      RECT 9.3560 31.5765 16.3580 32.6700 ;
      RECT 8.6090 31.5765 9.3380 32.4920 ;
      RECT 8.4470 31.7720 8.5730 32.6700 ;
      RECT 7.1960 31.6760 8.4200 32.4920 ;
      RECT 0.1760 31.5765 7.1780 32.6700 ;
      RECT 0.0050 31.5765 0.1580 32.4920 ;
      RECT 8.5550 31.5765 16.5290 32.3960 ;
      RECT 0.0050 31.6760 8.5370 32.3960 ;
      RECT 8.3300 31.5765 16.5290 31.7480 ;
      RECT 0.0050 31.5765 8.3120 32.3960 ;
      RECT 0.0050 31.5765 16.5290 31.6520 ;
      RECT 0.0050 33.6200 16.5290 33.7500 ;
      RECT 16.4120 32.6565 16.5290 33.7500 ;
      RECT 9.3020 33.5240 16.3940 33.7500 ;
      RECT 7.9700 33.5240 9.2840 33.7500 ;
      RECT 7.2500 32.6565 7.8800 33.7500 ;
      RECT 0.1400 33.5240 7.2320 33.7500 ;
      RECT 0.0050 32.6565 0.1220 33.7500 ;
      RECT 16.3760 32.6565 16.5290 33.5720 ;
      RECT 9.3560 32.6565 16.3580 33.7500 ;
      RECT 8.6090 32.6565 9.3380 33.5720 ;
      RECT 8.4470 32.8520 8.5730 33.7500 ;
      RECT 7.1960 32.7560 8.4200 33.5720 ;
      RECT 0.1760 32.6565 7.1780 33.7500 ;
      RECT 0.0050 32.6565 0.1580 33.5720 ;
      RECT 8.5550 32.6565 16.5290 33.4760 ;
      RECT 0.0050 32.7560 8.5370 33.4760 ;
      RECT 8.3300 32.6565 16.5290 32.8280 ;
      RECT 0.0050 32.6565 8.3120 33.4760 ;
      RECT 0.0050 32.6565 16.5290 32.7320 ;
      RECT 0.0050 34.7000 16.5290 34.8300 ;
      RECT 16.4120 33.7365 16.5290 34.8300 ;
      RECT 9.3020 34.6040 16.3940 34.8300 ;
      RECT 7.9700 34.6040 9.2840 34.8300 ;
      RECT 7.2500 33.7365 7.8800 34.8300 ;
      RECT 0.1400 34.6040 7.2320 34.8300 ;
      RECT 0.0050 33.7365 0.1220 34.8300 ;
      RECT 16.3760 33.7365 16.5290 34.6520 ;
      RECT 9.3560 33.7365 16.3580 34.8300 ;
      RECT 8.6090 33.7365 9.3380 34.6520 ;
      RECT 8.4470 33.9320 8.5730 34.8300 ;
      RECT 7.1960 33.8360 8.4200 34.6520 ;
      RECT 0.1760 33.7365 7.1780 34.8300 ;
      RECT 0.0050 33.7365 0.1580 34.6520 ;
      RECT 8.5550 33.7365 16.5290 34.5560 ;
      RECT 0.0050 33.8360 8.5370 34.5560 ;
      RECT 8.3300 33.7365 16.5290 33.9080 ;
      RECT 0.0050 33.7365 8.3120 34.5560 ;
      RECT 0.0050 33.7365 16.5290 33.8120 ;
      RECT 0.0050 35.7800 16.5290 35.9100 ;
      RECT 16.4120 34.8165 16.5290 35.9100 ;
      RECT 9.3020 35.6840 16.3940 35.9100 ;
      RECT 7.9700 35.6840 9.2840 35.9100 ;
      RECT 7.2500 34.8165 7.8800 35.9100 ;
      RECT 0.1400 35.6840 7.2320 35.9100 ;
      RECT 0.0050 34.8165 0.1220 35.9100 ;
      RECT 16.3760 34.8165 16.5290 35.7320 ;
      RECT 9.3560 34.8165 16.3580 35.9100 ;
      RECT 8.6090 34.8165 9.3380 35.7320 ;
      RECT 8.4470 35.0120 8.5730 35.9100 ;
      RECT 7.1960 34.9160 8.4200 35.7320 ;
      RECT 0.1760 34.8165 7.1780 35.9100 ;
      RECT 0.0050 34.8165 0.1580 35.7320 ;
      RECT 8.5550 34.8165 16.5290 35.6360 ;
      RECT 0.0050 34.9160 8.5370 35.6360 ;
      RECT 8.3300 34.8165 16.5290 34.9880 ;
      RECT 0.0050 34.8165 8.3120 35.6360 ;
      RECT 0.0050 34.8165 16.5290 34.8920 ;
      RECT 0.0050 36.8600 16.5290 36.9900 ;
      RECT 16.4120 35.8965 16.5290 36.9900 ;
      RECT 9.3020 36.7640 16.3940 36.9900 ;
      RECT 7.9700 36.7640 9.2840 36.9900 ;
      RECT 7.2500 35.8965 7.8800 36.9900 ;
      RECT 0.1400 36.7640 7.2320 36.9900 ;
      RECT 0.0050 35.8965 0.1220 36.9900 ;
      RECT 16.3760 35.8965 16.5290 36.8120 ;
      RECT 9.3560 35.8965 16.3580 36.9900 ;
      RECT 8.6090 35.8965 9.3380 36.8120 ;
      RECT 8.4470 36.0920 8.5730 36.9900 ;
      RECT 7.1960 35.9960 8.4200 36.8120 ;
      RECT 0.1760 35.8965 7.1780 36.9900 ;
      RECT 0.0050 35.8965 0.1580 36.8120 ;
      RECT 8.5550 35.8965 16.5290 36.7160 ;
      RECT 0.0050 35.9960 8.5370 36.7160 ;
      RECT 8.3300 35.8965 16.5290 36.0680 ;
      RECT 0.0050 35.8965 8.3120 36.7160 ;
      RECT 0.0050 35.8965 16.5290 35.9720 ;
      RECT 0.0050 37.9400 16.5290 38.0700 ;
      RECT 16.4120 36.9765 16.5290 38.0700 ;
      RECT 9.3020 37.8440 16.3940 38.0700 ;
      RECT 7.9700 37.8440 9.2840 38.0700 ;
      RECT 7.2500 36.9765 7.8800 38.0700 ;
      RECT 0.1400 37.8440 7.2320 38.0700 ;
      RECT 0.0050 36.9765 0.1220 38.0700 ;
      RECT 16.3760 36.9765 16.5290 37.8920 ;
      RECT 9.3560 36.9765 16.3580 38.0700 ;
      RECT 8.6090 36.9765 9.3380 37.8920 ;
      RECT 8.4470 37.1720 8.5730 38.0700 ;
      RECT 7.1960 37.0760 8.4200 37.8920 ;
      RECT 0.1760 36.9765 7.1780 38.0700 ;
      RECT 0.0050 36.9765 0.1580 37.8920 ;
      RECT 8.5550 36.9765 16.5290 37.7960 ;
      RECT 0.0050 37.0760 8.5370 37.7960 ;
      RECT 8.3300 36.9765 16.5290 37.1480 ;
      RECT 0.0050 36.9765 8.3120 37.7960 ;
      RECT 0.0050 36.9765 16.5290 37.0520 ;
      RECT 0.0050 39.0200 16.5290 39.1500 ;
      RECT 16.4120 38.0565 16.5290 39.1500 ;
      RECT 9.3020 38.9240 16.3940 39.1500 ;
      RECT 7.9700 38.9240 9.2840 39.1500 ;
      RECT 7.2500 38.0565 7.8800 39.1500 ;
      RECT 0.1400 38.9240 7.2320 39.1500 ;
      RECT 0.0050 38.0565 0.1220 39.1500 ;
      RECT 16.3760 38.0565 16.5290 38.9720 ;
      RECT 9.3560 38.0565 16.3580 39.1500 ;
      RECT 8.6090 38.0565 9.3380 38.9720 ;
      RECT 8.4470 38.2520 8.5730 39.1500 ;
      RECT 7.1960 38.1560 8.4200 38.9720 ;
      RECT 0.1760 38.0565 7.1780 39.1500 ;
      RECT 0.0050 38.0565 0.1580 38.9720 ;
      RECT 8.5550 38.0565 16.5290 38.8760 ;
      RECT 0.0050 38.1560 8.5370 38.8760 ;
      RECT 8.3300 38.0565 16.5290 38.2280 ;
      RECT 0.0050 38.0565 8.3120 38.8760 ;
      RECT 0.0050 38.0565 16.5290 38.1320 ;
      RECT 0.0050 40.1000 16.5290 40.2300 ;
      RECT 16.4120 39.1365 16.5290 40.2300 ;
      RECT 9.3020 40.0040 16.3940 40.2300 ;
      RECT 7.9700 40.0040 9.2840 40.2300 ;
      RECT 7.2500 39.1365 7.8800 40.2300 ;
      RECT 0.1400 40.0040 7.2320 40.2300 ;
      RECT 0.0050 39.1365 0.1220 40.2300 ;
      RECT 16.3760 39.1365 16.5290 40.0520 ;
      RECT 9.3560 39.1365 16.3580 40.2300 ;
      RECT 8.6090 39.1365 9.3380 40.0520 ;
      RECT 8.4470 39.3320 8.5730 40.2300 ;
      RECT 7.1960 39.2360 8.4200 40.0520 ;
      RECT 0.1760 39.1365 7.1780 40.2300 ;
      RECT 0.0050 39.1365 0.1580 40.0520 ;
      RECT 8.5550 39.1365 16.5290 39.9560 ;
      RECT 0.0050 39.2360 8.5370 39.9560 ;
      RECT 8.3300 39.1365 16.5290 39.3080 ;
      RECT 0.0050 39.1365 8.3120 39.9560 ;
      RECT 0.0050 39.1365 16.5290 39.2120 ;
      RECT 0.0000 47.5170 16.5240 48.8505 ;
      RECT 10.8090 40.1970 16.5240 48.8505 ;
      RECT 8.6090 44.0610 16.5240 48.8505 ;
      RECT 9.5130 41.4690 16.5240 48.8505 ;
      RECT 8.5570 40.1970 8.5910 48.8505 ;
      RECT 8.5050 40.1970 8.5390 48.8505 ;
      RECT 8.4530 40.1970 8.4870 48.8505 ;
      RECT 8.4010 40.1970 8.4350 48.8505 ;
      RECT 0.0000 47.0850 8.3830 48.8505 ;
      RECT 8.1410 44.3490 16.5240 47.3010 ;
      RECT 8.0890 40.1970 8.1230 48.8505 ;
      RECT 8.0370 40.1970 8.0710 48.8505 ;
      RECT 7.9850 40.1970 8.0190 48.8505 ;
      RECT 7.9330 40.1970 7.9670 48.8505 ;
      RECT 0.0000 41.7570 7.9150 48.8505 ;
      RECT 0.0000 43.9170 8.3830 46.8690 ;
      RECT 8.1410 41.1810 9.2790 44.1330 ;
      RECT 9.3150 41.6610 16.5240 48.8505 ;
      RECT 0.0000 43.9170 9.2970 44.1330 ;
      RECT 8.1410 41.6610 16.5240 44.0370 ;
      RECT 7.4610 40.7490 8.2350 43.7010 ;
      RECT 7.2450 40.8930 7.9150 48.8505 ;
      RECT 0.0000 41.4690 7.2270 48.8505 ;
      RECT 6.8130 40.1970 7.2630 41.7330 ;
      RECT 0.0000 41.5650 9.4950 41.7330 ;
      RECT 9.2970 41.4690 16.5240 41.6370 ;
      RECT 10.5930 40.1970 10.7910 48.8505 ;
      RECT 6.8130 41.2770 10.5750 41.5410 ;
      RECT 5.9490 40.8930 6.7950 48.8505 ;
      RECT 0.0000 40.1970 5.9310 48.8505 ;
      RECT 10.3770 40.1970 16.5240 41.4450 ;
      RECT 10.1610 40.8930 16.5240 41.4450 ;
      RECT 0.0000 41.1815 10.1430 41.4450 ;
      RECT 9.9450 40.1970 10.3590 41.2530 ;
      RECT 9.3510 40.8930 16.5240 41.2530 ;
      RECT 8.6090 40.8930 9.3330 41.5410 ;
      RECT 8.1410 40.8450 8.3830 48.8505 ;
      RECT 8.2530 40.1970 8.6310 40.9650 ;
      RECT 8.6490 40.8450 9.9270 40.9655 ;
      RECT 6.5970 40.8450 7.4430 41.4450 ;
      RECT 6.1650 40.8450 6.5790 48.8505 ;
      RECT 0.0000 40.1970 6.1470 41.4450 ;
      RECT 9.7290 40.1970 16.5240 40.8690 ;
      RECT 8.2530 40.2770 9.7110 40.8690 ;
      RECT 7.2810 40.7490 8.2350 40.8690 ;
      RECT 6.3810 40.1970 7.2630 40.8690 ;
      RECT 0.0000 40.1970 6.3630 40.8690 ;
      RECT 9.2970 40.1970 16.5240 40.8210 ;
      RECT 8.1410 40.2770 16.5240 40.8210 ;
      RECT 0.0000 40.1970 7.9150 40.8210 ;
      RECT 0.0000 40.1970 9.2790 40.5330 ;
      RECT 0.0000 40.1970 16.5240 40.2530 ;
        RECT 0.0050 49.3070 16.5290 49.4370 ;
        RECT 16.4120 48.3435 16.5290 49.4370 ;
        RECT 9.3020 49.2110 16.3940 49.4370 ;
        RECT 7.9700 49.2110 9.2840 49.4370 ;
        RECT 7.2500 48.3435 7.8800 49.4370 ;
        RECT 0.1400 49.2110 7.2320 49.4370 ;
        RECT 0.0050 48.3435 0.1220 49.4370 ;
        RECT 16.3760 48.3435 16.5290 49.2590 ;
        RECT 9.3560 48.3435 16.3580 49.4370 ;
        RECT 8.6090 48.3435 9.3380 49.2590 ;
        RECT 8.4470 48.5390 8.5730 49.4370 ;
        RECT 7.1960 48.4430 8.4200 49.2590 ;
        RECT 0.1760 48.3435 7.1780 49.4370 ;
        RECT 0.0050 48.3435 0.1580 49.2590 ;
        RECT 8.5550 48.3435 16.5290 49.1630 ;
        RECT 0.0050 48.4430 8.5370 49.1630 ;
        RECT 8.3300 48.3435 16.5290 48.5150 ;
        RECT 0.0050 48.3435 8.3120 49.1630 ;
        RECT 0.0050 48.3435 16.5290 48.4190 ;
        RECT 0.0050 50.3870 16.5290 50.5170 ;
        RECT 16.4120 49.4235 16.5290 50.5170 ;
        RECT 9.3020 50.2910 16.3940 50.5170 ;
        RECT 7.9700 50.2910 9.2840 50.5170 ;
        RECT 7.2500 49.4235 7.8800 50.5170 ;
        RECT 0.1400 50.2910 7.2320 50.5170 ;
        RECT 0.0050 49.4235 0.1220 50.5170 ;
        RECT 16.3760 49.4235 16.5290 50.3390 ;
        RECT 9.3560 49.4235 16.3580 50.5170 ;
        RECT 8.6090 49.4235 9.3380 50.3390 ;
        RECT 8.4470 49.6190 8.5730 50.5170 ;
        RECT 7.1960 49.5230 8.4200 50.3390 ;
        RECT 0.1760 49.4235 7.1780 50.5170 ;
        RECT 0.0050 49.4235 0.1580 50.3390 ;
        RECT 8.5550 49.4235 16.5290 50.2430 ;
        RECT 0.0050 49.5230 8.5370 50.2430 ;
        RECT 8.3300 49.4235 16.5290 49.5950 ;
        RECT 0.0050 49.4235 8.3120 50.2430 ;
        RECT 0.0050 49.4235 16.5290 49.4990 ;
        RECT 0.0050 51.4670 16.5290 51.5970 ;
        RECT 16.4120 50.5035 16.5290 51.5970 ;
        RECT 9.3020 51.3710 16.3940 51.5970 ;
        RECT 7.9700 51.3710 9.2840 51.5970 ;
        RECT 7.2500 50.5035 7.8800 51.5970 ;
        RECT 0.1400 51.3710 7.2320 51.5970 ;
        RECT 0.0050 50.5035 0.1220 51.5970 ;
        RECT 16.3760 50.5035 16.5290 51.4190 ;
        RECT 9.3560 50.5035 16.3580 51.5970 ;
        RECT 8.6090 50.5035 9.3380 51.4190 ;
        RECT 8.4470 50.6990 8.5730 51.5970 ;
        RECT 7.1960 50.6030 8.4200 51.4190 ;
        RECT 0.1760 50.5035 7.1780 51.5970 ;
        RECT 0.0050 50.5035 0.1580 51.4190 ;
        RECT 8.5550 50.5035 16.5290 51.3230 ;
        RECT 0.0050 50.6030 8.5370 51.3230 ;
        RECT 8.3300 50.5035 16.5290 50.6750 ;
        RECT 0.0050 50.5035 8.3120 51.3230 ;
        RECT 0.0050 50.5035 16.5290 50.5790 ;
        RECT 0.0050 52.5470 16.5290 52.6770 ;
        RECT 16.4120 51.5835 16.5290 52.6770 ;
        RECT 9.3020 52.4510 16.3940 52.6770 ;
        RECT 7.9700 52.4510 9.2840 52.6770 ;
        RECT 7.2500 51.5835 7.8800 52.6770 ;
        RECT 0.1400 52.4510 7.2320 52.6770 ;
        RECT 0.0050 51.5835 0.1220 52.6770 ;
        RECT 16.3760 51.5835 16.5290 52.4990 ;
        RECT 9.3560 51.5835 16.3580 52.6770 ;
        RECT 8.6090 51.5835 9.3380 52.4990 ;
        RECT 8.4470 51.7790 8.5730 52.6770 ;
        RECT 7.1960 51.6830 8.4200 52.4990 ;
        RECT 0.1760 51.5835 7.1780 52.6770 ;
        RECT 0.0050 51.5835 0.1580 52.4990 ;
        RECT 8.5550 51.5835 16.5290 52.4030 ;
        RECT 0.0050 51.6830 8.5370 52.4030 ;
        RECT 8.3300 51.5835 16.5290 51.7550 ;
        RECT 0.0050 51.5835 8.3120 52.4030 ;
        RECT 0.0050 51.5835 16.5290 51.6590 ;
        RECT 0.0050 53.6270 16.5290 53.7570 ;
        RECT 16.4120 52.6635 16.5290 53.7570 ;
        RECT 9.3020 53.5310 16.3940 53.7570 ;
        RECT 7.9700 53.5310 9.2840 53.7570 ;
        RECT 7.2500 52.6635 7.8800 53.7570 ;
        RECT 0.1400 53.5310 7.2320 53.7570 ;
        RECT 0.0050 52.6635 0.1220 53.7570 ;
        RECT 16.3760 52.6635 16.5290 53.5790 ;
        RECT 9.3560 52.6635 16.3580 53.7570 ;
        RECT 8.6090 52.6635 9.3380 53.5790 ;
        RECT 8.4470 52.8590 8.5730 53.7570 ;
        RECT 7.1960 52.7630 8.4200 53.5790 ;
        RECT 0.1760 52.6635 7.1780 53.7570 ;
        RECT 0.0050 52.6635 0.1580 53.5790 ;
        RECT 8.5550 52.6635 16.5290 53.4830 ;
        RECT 0.0050 52.7630 8.5370 53.4830 ;
        RECT 8.3300 52.6635 16.5290 52.8350 ;
        RECT 0.0050 52.6635 8.3120 53.4830 ;
        RECT 0.0050 52.6635 16.5290 52.7390 ;
        RECT 0.0050 54.7070 16.5290 54.8370 ;
        RECT 16.4120 53.7435 16.5290 54.8370 ;
        RECT 9.3020 54.6110 16.3940 54.8370 ;
        RECT 7.9700 54.6110 9.2840 54.8370 ;
        RECT 7.2500 53.7435 7.8800 54.8370 ;
        RECT 0.1400 54.6110 7.2320 54.8370 ;
        RECT 0.0050 53.7435 0.1220 54.8370 ;
        RECT 16.3760 53.7435 16.5290 54.6590 ;
        RECT 9.3560 53.7435 16.3580 54.8370 ;
        RECT 8.6090 53.7435 9.3380 54.6590 ;
        RECT 8.4470 53.9390 8.5730 54.8370 ;
        RECT 7.1960 53.8430 8.4200 54.6590 ;
        RECT 0.1760 53.7435 7.1780 54.8370 ;
        RECT 0.0050 53.7435 0.1580 54.6590 ;
        RECT 8.5550 53.7435 16.5290 54.5630 ;
        RECT 0.0050 53.8430 8.5370 54.5630 ;
        RECT 8.3300 53.7435 16.5290 53.9150 ;
        RECT 0.0050 53.7435 8.3120 54.5630 ;
        RECT 0.0050 53.7435 16.5290 53.8190 ;
        RECT 0.0050 55.7870 16.5290 55.9170 ;
        RECT 16.4120 54.8235 16.5290 55.9170 ;
        RECT 9.3020 55.6910 16.3940 55.9170 ;
        RECT 7.9700 55.6910 9.2840 55.9170 ;
        RECT 7.2500 54.8235 7.8800 55.9170 ;
        RECT 0.1400 55.6910 7.2320 55.9170 ;
        RECT 0.0050 54.8235 0.1220 55.9170 ;
        RECT 16.3760 54.8235 16.5290 55.7390 ;
        RECT 9.3560 54.8235 16.3580 55.9170 ;
        RECT 8.6090 54.8235 9.3380 55.7390 ;
        RECT 8.4470 55.0190 8.5730 55.9170 ;
        RECT 7.1960 54.9230 8.4200 55.7390 ;
        RECT 0.1760 54.8235 7.1780 55.9170 ;
        RECT 0.0050 54.8235 0.1580 55.7390 ;
        RECT 8.5550 54.8235 16.5290 55.6430 ;
        RECT 0.0050 54.9230 8.5370 55.6430 ;
        RECT 8.3300 54.8235 16.5290 54.9950 ;
        RECT 0.0050 54.8235 8.3120 55.6430 ;
        RECT 0.0050 54.8235 16.5290 54.8990 ;
        RECT 0.0050 56.8670 16.5290 56.9970 ;
        RECT 16.4120 55.9035 16.5290 56.9970 ;
        RECT 9.3020 56.7710 16.3940 56.9970 ;
        RECT 7.9700 56.7710 9.2840 56.9970 ;
        RECT 7.2500 55.9035 7.8800 56.9970 ;
        RECT 0.1400 56.7710 7.2320 56.9970 ;
        RECT 0.0050 55.9035 0.1220 56.9970 ;
        RECT 16.3760 55.9035 16.5290 56.8190 ;
        RECT 9.3560 55.9035 16.3580 56.9970 ;
        RECT 8.6090 55.9035 9.3380 56.8190 ;
        RECT 8.4470 56.0990 8.5730 56.9970 ;
        RECT 7.1960 56.0030 8.4200 56.8190 ;
        RECT 0.1760 55.9035 7.1780 56.9970 ;
        RECT 0.0050 55.9035 0.1580 56.8190 ;
        RECT 8.5550 55.9035 16.5290 56.7230 ;
        RECT 0.0050 56.0030 8.5370 56.7230 ;
        RECT 8.3300 55.9035 16.5290 56.0750 ;
        RECT 0.0050 55.9035 8.3120 56.7230 ;
        RECT 0.0050 55.9035 16.5290 55.9790 ;
        RECT 0.0050 57.9470 16.5290 58.0770 ;
        RECT 16.4120 56.9835 16.5290 58.0770 ;
        RECT 9.3020 57.8510 16.3940 58.0770 ;
        RECT 7.9700 57.8510 9.2840 58.0770 ;
        RECT 7.2500 56.9835 7.8800 58.0770 ;
        RECT 0.1400 57.8510 7.2320 58.0770 ;
        RECT 0.0050 56.9835 0.1220 58.0770 ;
        RECT 16.3760 56.9835 16.5290 57.8990 ;
        RECT 9.3560 56.9835 16.3580 58.0770 ;
        RECT 8.6090 56.9835 9.3380 57.8990 ;
        RECT 8.4470 57.1790 8.5730 58.0770 ;
        RECT 7.1960 57.0830 8.4200 57.8990 ;
        RECT 0.1760 56.9835 7.1780 58.0770 ;
        RECT 0.0050 56.9835 0.1580 57.8990 ;
        RECT 8.5550 56.9835 16.5290 57.8030 ;
        RECT 0.0050 57.0830 8.5370 57.8030 ;
        RECT 8.3300 56.9835 16.5290 57.1550 ;
        RECT 0.0050 56.9835 8.3120 57.8030 ;
        RECT 0.0050 56.9835 16.5290 57.0590 ;
        RECT 0.0050 59.0270 16.5290 59.1570 ;
        RECT 16.4120 58.0635 16.5290 59.1570 ;
        RECT 9.3020 58.9310 16.3940 59.1570 ;
        RECT 7.9700 58.9310 9.2840 59.1570 ;
        RECT 7.2500 58.0635 7.8800 59.1570 ;
        RECT 0.1400 58.9310 7.2320 59.1570 ;
        RECT 0.0050 58.0635 0.1220 59.1570 ;
        RECT 16.3760 58.0635 16.5290 58.9790 ;
        RECT 9.3560 58.0635 16.3580 59.1570 ;
        RECT 8.6090 58.0635 9.3380 58.9790 ;
        RECT 8.4470 58.2590 8.5730 59.1570 ;
        RECT 7.1960 58.1630 8.4200 58.9790 ;
        RECT 0.1760 58.0635 7.1780 59.1570 ;
        RECT 0.0050 58.0635 0.1580 58.9790 ;
        RECT 8.5550 58.0635 16.5290 58.8830 ;
        RECT 0.0050 58.1630 8.5370 58.8830 ;
        RECT 8.3300 58.0635 16.5290 58.2350 ;
        RECT 0.0050 58.0635 8.3120 58.8830 ;
        RECT 0.0050 58.0635 16.5290 58.1390 ;
        RECT 0.0050 60.1070 16.5290 60.2370 ;
        RECT 16.4120 59.1435 16.5290 60.2370 ;
        RECT 9.3020 60.0110 16.3940 60.2370 ;
        RECT 7.9700 60.0110 9.2840 60.2370 ;
        RECT 7.2500 59.1435 7.8800 60.2370 ;
        RECT 0.1400 60.0110 7.2320 60.2370 ;
        RECT 0.0050 59.1435 0.1220 60.2370 ;
        RECT 16.3760 59.1435 16.5290 60.0590 ;
        RECT 9.3560 59.1435 16.3580 60.2370 ;
        RECT 8.6090 59.1435 9.3380 60.0590 ;
        RECT 8.4470 59.3390 8.5730 60.2370 ;
        RECT 7.1960 59.2430 8.4200 60.0590 ;
        RECT 0.1760 59.1435 7.1780 60.2370 ;
        RECT 0.0050 59.1435 0.1580 60.0590 ;
        RECT 8.5550 59.1435 16.5290 59.9630 ;
        RECT 0.0050 59.2430 8.5370 59.9630 ;
        RECT 8.3300 59.1435 16.5290 59.3150 ;
        RECT 0.0050 59.1435 8.3120 59.9630 ;
        RECT 0.0050 59.1435 16.5290 59.2190 ;
        RECT 0.0050 61.1870 16.5290 61.3170 ;
        RECT 16.4120 60.2235 16.5290 61.3170 ;
        RECT 9.3020 61.0910 16.3940 61.3170 ;
        RECT 7.9700 61.0910 9.2840 61.3170 ;
        RECT 7.2500 60.2235 7.8800 61.3170 ;
        RECT 0.1400 61.0910 7.2320 61.3170 ;
        RECT 0.0050 60.2235 0.1220 61.3170 ;
        RECT 16.3760 60.2235 16.5290 61.1390 ;
        RECT 9.3560 60.2235 16.3580 61.3170 ;
        RECT 8.6090 60.2235 9.3380 61.1390 ;
        RECT 8.4470 60.4190 8.5730 61.3170 ;
        RECT 7.1960 60.3230 8.4200 61.1390 ;
        RECT 0.1760 60.2235 7.1780 61.3170 ;
        RECT 0.0050 60.2235 0.1580 61.1390 ;
        RECT 8.5550 60.2235 16.5290 61.0430 ;
        RECT 0.0050 60.3230 8.5370 61.0430 ;
        RECT 8.3300 60.2235 16.5290 60.3950 ;
        RECT 0.0050 60.2235 8.3120 61.0430 ;
        RECT 0.0050 60.2235 16.5290 60.2990 ;
        RECT 0.0050 62.2670 16.5290 62.3970 ;
        RECT 16.4120 61.3035 16.5290 62.3970 ;
        RECT 9.3020 62.1710 16.3940 62.3970 ;
        RECT 7.9700 62.1710 9.2840 62.3970 ;
        RECT 7.2500 61.3035 7.8800 62.3970 ;
        RECT 0.1400 62.1710 7.2320 62.3970 ;
        RECT 0.0050 61.3035 0.1220 62.3970 ;
        RECT 16.3760 61.3035 16.5290 62.2190 ;
        RECT 9.3560 61.3035 16.3580 62.3970 ;
        RECT 8.6090 61.3035 9.3380 62.2190 ;
        RECT 8.4470 61.4990 8.5730 62.3970 ;
        RECT 7.1960 61.4030 8.4200 62.2190 ;
        RECT 0.1760 61.3035 7.1780 62.3970 ;
        RECT 0.0050 61.3035 0.1580 62.2190 ;
        RECT 8.5550 61.3035 16.5290 62.1230 ;
        RECT 0.0050 61.4030 8.5370 62.1230 ;
        RECT 8.3300 61.3035 16.5290 61.4750 ;
        RECT 0.0050 61.3035 8.3120 62.1230 ;
        RECT 0.0050 61.3035 16.5290 61.3790 ;
        RECT 0.0050 63.3470 16.5290 63.4770 ;
        RECT 16.4120 62.3835 16.5290 63.4770 ;
        RECT 9.3020 63.2510 16.3940 63.4770 ;
        RECT 7.9700 63.2510 9.2840 63.4770 ;
        RECT 7.2500 62.3835 7.8800 63.4770 ;
        RECT 0.1400 63.2510 7.2320 63.4770 ;
        RECT 0.0050 62.3835 0.1220 63.4770 ;
        RECT 16.3760 62.3835 16.5290 63.2990 ;
        RECT 9.3560 62.3835 16.3580 63.4770 ;
        RECT 8.6090 62.3835 9.3380 63.2990 ;
        RECT 8.4470 62.5790 8.5730 63.4770 ;
        RECT 7.1960 62.4830 8.4200 63.2990 ;
        RECT 0.1760 62.3835 7.1780 63.4770 ;
        RECT 0.0050 62.3835 0.1580 63.2990 ;
        RECT 8.5550 62.3835 16.5290 63.2030 ;
        RECT 0.0050 62.4830 8.5370 63.2030 ;
        RECT 8.3300 62.3835 16.5290 62.5550 ;
        RECT 0.0050 62.3835 8.3120 63.2030 ;
        RECT 0.0050 62.3835 16.5290 62.4590 ;
        RECT 0.0050 64.4270 16.5290 64.5570 ;
        RECT 16.4120 63.4635 16.5290 64.5570 ;
        RECT 9.3020 64.3310 16.3940 64.5570 ;
        RECT 7.9700 64.3310 9.2840 64.5570 ;
        RECT 7.2500 63.4635 7.8800 64.5570 ;
        RECT 0.1400 64.3310 7.2320 64.5570 ;
        RECT 0.0050 63.4635 0.1220 64.5570 ;
        RECT 16.3760 63.4635 16.5290 64.3790 ;
        RECT 9.3560 63.4635 16.3580 64.5570 ;
        RECT 8.6090 63.4635 9.3380 64.3790 ;
        RECT 8.4470 63.6590 8.5730 64.5570 ;
        RECT 7.1960 63.5630 8.4200 64.3790 ;
        RECT 0.1760 63.4635 7.1780 64.5570 ;
        RECT 0.0050 63.4635 0.1580 64.3790 ;
        RECT 8.5550 63.4635 16.5290 64.2830 ;
        RECT 0.0050 63.5630 8.5370 64.2830 ;
        RECT 8.3300 63.4635 16.5290 63.6350 ;
        RECT 0.0050 63.4635 8.3120 64.2830 ;
        RECT 0.0050 63.4635 16.5290 63.5390 ;
        RECT 0.0050 65.5070 16.5290 65.6370 ;
        RECT 16.4120 64.5435 16.5290 65.6370 ;
        RECT 9.3020 65.4110 16.3940 65.6370 ;
        RECT 7.9700 65.4110 9.2840 65.6370 ;
        RECT 7.2500 64.5435 7.8800 65.6370 ;
        RECT 0.1400 65.4110 7.2320 65.6370 ;
        RECT 0.0050 64.5435 0.1220 65.6370 ;
        RECT 16.3760 64.5435 16.5290 65.4590 ;
        RECT 9.3560 64.5435 16.3580 65.6370 ;
        RECT 8.6090 64.5435 9.3380 65.4590 ;
        RECT 8.4470 64.7390 8.5730 65.6370 ;
        RECT 7.1960 64.6430 8.4200 65.4590 ;
        RECT 0.1760 64.5435 7.1780 65.6370 ;
        RECT 0.0050 64.5435 0.1580 65.4590 ;
        RECT 8.5550 64.5435 16.5290 65.3630 ;
        RECT 0.0050 64.6430 8.5370 65.3630 ;
        RECT 8.3300 64.5435 16.5290 64.7150 ;
        RECT 0.0050 64.5435 8.3120 65.3630 ;
        RECT 0.0050 64.5435 16.5290 64.6190 ;
        RECT 0.0050 66.5870 16.5290 66.7170 ;
        RECT 16.4120 65.6235 16.5290 66.7170 ;
        RECT 9.3020 66.4910 16.3940 66.7170 ;
        RECT 7.9700 66.4910 9.2840 66.7170 ;
        RECT 7.2500 65.6235 7.8800 66.7170 ;
        RECT 0.1400 66.4910 7.2320 66.7170 ;
        RECT 0.0050 65.6235 0.1220 66.7170 ;
        RECT 16.3760 65.6235 16.5290 66.5390 ;
        RECT 9.3560 65.6235 16.3580 66.7170 ;
        RECT 8.6090 65.6235 9.3380 66.5390 ;
        RECT 8.4470 65.8190 8.5730 66.7170 ;
        RECT 7.1960 65.7230 8.4200 66.5390 ;
        RECT 0.1760 65.6235 7.1780 66.7170 ;
        RECT 0.0050 65.6235 0.1580 66.5390 ;
        RECT 8.5550 65.6235 16.5290 66.4430 ;
        RECT 0.0050 65.7230 8.5370 66.4430 ;
        RECT 8.3300 65.6235 16.5290 65.7950 ;
        RECT 0.0050 65.6235 8.3120 66.4430 ;
        RECT 0.0050 65.6235 16.5290 65.6990 ;
        RECT 0.0050 67.6670 16.5290 67.7970 ;
        RECT 16.4120 66.7035 16.5290 67.7970 ;
        RECT 9.3020 67.5710 16.3940 67.7970 ;
        RECT 7.9700 67.5710 9.2840 67.7970 ;
        RECT 7.2500 66.7035 7.8800 67.7970 ;
        RECT 0.1400 67.5710 7.2320 67.7970 ;
        RECT 0.0050 66.7035 0.1220 67.7970 ;
        RECT 16.3760 66.7035 16.5290 67.6190 ;
        RECT 9.3560 66.7035 16.3580 67.7970 ;
        RECT 8.6090 66.7035 9.3380 67.6190 ;
        RECT 8.4470 66.8990 8.5730 67.7970 ;
        RECT 7.1960 66.8030 8.4200 67.6190 ;
        RECT 0.1760 66.7035 7.1780 67.7970 ;
        RECT 0.0050 66.7035 0.1580 67.6190 ;
        RECT 8.5550 66.7035 16.5290 67.5230 ;
        RECT 0.0050 66.8030 8.5370 67.5230 ;
        RECT 8.3300 66.7035 16.5290 66.8750 ;
        RECT 0.0050 66.7035 8.3120 67.5230 ;
        RECT 0.0050 66.7035 16.5290 66.7790 ;
        RECT 0.0050 68.7470 16.5290 68.8770 ;
        RECT 16.4120 67.7835 16.5290 68.8770 ;
        RECT 9.3020 68.6510 16.3940 68.8770 ;
        RECT 7.9700 68.6510 9.2840 68.8770 ;
        RECT 7.2500 67.7835 7.8800 68.8770 ;
        RECT 0.1400 68.6510 7.2320 68.8770 ;
        RECT 0.0050 67.7835 0.1220 68.8770 ;
        RECT 16.3760 67.7835 16.5290 68.6990 ;
        RECT 9.3560 67.7835 16.3580 68.8770 ;
        RECT 8.6090 67.7835 9.3380 68.6990 ;
        RECT 8.4470 67.9790 8.5730 68.8770 ;
        RECT 7.1960 67.8830 8.4200 68.6990 ;
        RECT 0.1760 67.7835 7.1780 68.8770 ;
        RECT 0.0050 67.7835 0.1580 68.6990 ;
        RECT 8.5550 67.7835 16.5290 68.6030 ;
        RECT 0.0050 67.8830 8.5370 68.6030 ;
        RECT 8.3300 67.7835 16.5290 67.9550 ;
        RECT 0.0050 67.7835 8.3120 68.6030 ;
        RECT 0.0050 67.7835 16.5290 67.8590 ;
        RECT 0.0050 69.8270 16.5290 69.9570 ;
        RECT 16.4120 68.8635 16.5290 69.9570 ;
        RECT 9.3020 69.7310 16.3940 69.9570 ;
        RECT 7.9700 69.7310 9.2840 69.9570 ;
        RECT 7.2500 68.8635 7.8800 69.9570 ;
        RECT 0.1400 69.7310 7.2320 69.9570 ;
        RECT 0.0050 68.8635 0.1220 69.9570 ;
        RECT 16.3760 68.8635 16.5290 69.7790 ;
        RECT 9.3560 68.8635 16.3580 69.9570 ;
        RECT 8.6090 68.8635 9.3380 69.7790 ;
        RECT 8.4470 69.0590 8.5730 69.9570 ;
        RECT 7.1960 68.9630 8.4200 69.7790 ;
        RECT 0.1760 68.8635 7.1780 69.9570 ;
        RECT 0.0050 68.8635 0.1580 69.7790 ;
        RECT 8.5550 68.8635 16.5290 69.6830 ;
        RECT 0.0050 68.9630 8.5370 69.6830 ;
        RECT 8.3300 68.8635 16.5290 69.0350 ;
        RECT 0.0050 68.8635 8.3120 69.6830 ;
        RECT 0.0050 68.8635 16.5290 68.9390 ;
        RECT 0.0050 70.9070 16.5290 71.0370 ;
        RECT 16.4120 69.9435 16.5290 71.0370 ;
        RECT 9.3020 70.8110 16.3940 71.0370 ;
        RECT 7.9700 70.8110 9.2840 71.0370 ;
        RECT 7.2500 69.9435 7.8800 71.0370 ;
        RECT 0.1400 70.8110 7.2320 71.0370 ;
        RECT 0.0050 69.9435 0.1220 71.0370 ;
        RECT 16.3760 69.9435 16.5290 70.8590 ;
        RECT 9.3560 69.9435 16.3580 71.0370 ;
        RECT 8.6090 69.9435 9.3380 70.8590 ;
        RECT 8.4470 70.1390 8.5730 71.0370 ;
        RECT 7.1960 70.0430 8.4200 70.8590 ;
        RECT 0.1760 69.9435 7.1780 71.0370 ;
        RECT 0.0050 69.9435 0.1580 70.8590 ;
        RECT 8.5550 69.9435 16.5290 70.7630 ;
        RECT 0.0050 70.0430 8.5370 70.7630 ;
        RECT 8.3300 69.9435 16.5290 70.1150 ;
        RECT 0.0050 69.9435 8.3120 70.7630 ;
        RECT 0.0050 69.9435 16.5290 70.0190 ;
        RECT 0.0050 71.9870 16.5290 72.1170 ;
        RECT 16.4120 71.0235 16.5290 72.1170 ;
        RECT 9.3020 71.8910 16.3940 72.1170 ;
        RECT 7.9700 71.8910 9.2840 72.1170 ;
        RECT 7.2500 71.0235 7.8800 72.1170 ;
        RECT 0.1400 71.8910 7.2320 72.1170 ;
        RECT 0.0050 71.0235 0.1220 72.1170 ;
        RECT 16.3760 71.0235 16.5290 71.9390 ;
        RECT 9.3560 71.0235 16.3580 72.1170 ;
        RECT 8.6090 71.0235 9.3380 71.9390 ;
        RECT 8.4470 71.2190 8.5730 72.1170 ;
        RECT 7.1960 71.1230 8.4200 71.9390 ;
        RECT 0.1760 71.0235 7.1780 72.1170 ;
        RECT 0.0050 71.0235 0.1580 71.9390 ;
        RECT 8.5550 71.0235 16.5290 71.8430 ;
        RECT 0.0050 71.1230 8.5370 71.8430 ;
        RECT 8.3300 71.0235 16.5290 71.1950 ;
        RECT 0.0050 71.0235 8.3120 71.8430 ;
        RECT 0.0050 71.0235 16.5290 71.0990 ;
        RECT 0.0050 73.0670 16.5290 73.1970 ;
        RECT 16.4120 72.1035 16.5290 73.1970 ;
        RECT 9.3020 72.9710 16.3940 73.1970 ;
        RECT 7.9700 72.9710 9.2840 73.1970 ;
        RECT 7.2500 72.1035 7.8800 73.1970 ;
        RECT 0.1400 72.9710 7.2320 73.1970 ;
        RECT 0.0050 72.1035 0.1220 73.1970 ;
        RECT 16.3760 72.1035 16.5290 73.0190 ;
        RECT 9.3560 72.1035 16.3580 73.1970 ;
        RECT 8.6090 72.1035 9.3380 73.0190 ;
        RECT 8.4470 72.2990 8.5730 73.1970 ;
        RECT 7.1960 72.2030 8.4200 73.0190 ;
        RECT 0.1760 72.1035 7.1780 73.1970 ;
        RECT 0.0050 72.1035 0.1580 73.0190 ;
        RECT 8.5550 72.1035 16.5290 72.9230 ;
        RECT 0.0050 72.2030 8.5370 72.9230 ;
        RECT 8.3300 72.1035 16.5290 72.2750 ;
        RECT 0.0050 72.1035 8.3120 72.9230 ;
        RECT 0.0050 72.1035 16.5290 72.1790 ;
        RECT 0.0050 74.1470 16.5290 74.2770 ;
        RECT 16.4120 73.1835 16.5290 74.2770 ;
        RECT 9.3020 74.0510 16.3940 74.2770 ;
        RECT 7.9700 74.0510 9.2840 74.2770 ;
        RECT 7.2500 73.1835 7.8800 74.2770 ;
        RECT 0.1400 74.0510 7.2320 74.2770 ;
        RECT 0.0050 73.1835 0.1220 74.2770 ;
        RECT 16.3760 73.1835 16.5290 74.0990 ;
        RECT 9.3560 73.1835 16.3580 74.2770 ;
        RECT 8.6090 73.1835 9.3380 74.0990 ;
        RECT 8.4470 73.3790 8.5730 74.2770 ;
        RECT 7.1960 73.2830 8.4200 74.0990 ;
        RECT 0.1760 73.1835 7.1780 74.2770 ;
        RECT 0.0050 73.1835 0.1580 74.0990 ;
        RECT 8.5550 73.1835 16.5290 74.0030 ;
        RECT 0.0050 73.2830 8.5370 74.0030 ;
        RECT 8.3300 73.1835 16.5290 73.3550 ;
        RECT 0.0050 73.1835 8.3120 74.0030 ;
        RECT 0.0050 73.1835 16.5290 73.2590 ;
        RECT 0.0050 75.2270 16.5290 75.3570 ;
        RECT 16.4120 74.2635 16.5290 75.3570 ;
        RECT 9.3020 75.1310 16.3940 75.3570 ;
        RECT 7.9700 75.1310 9.2840 75.3570 ;
        RECT 7.2500 74.2635 7.8800 75.3570 ;
        RECT 0.1400 75.1310 7.2320 75.3570 ;
        RECT 0.0050 74.2635 0.1220 75.3570 ;
        RECT 16.3760 74.2635 16.5290 75.1790 ;
        RECT 9.3560 74.2635 16.3580 75.3570 ;
        RECT 8.6090 74.2635 9.3380 75.1790 ;
        RECT 8.4470 74.4590 8.5730 75.3570 ;
        RECT 7.1960 74.3630 8.4200 75.1790 ;
        RECT 0.1760 74.2635 7.1780 75.3570 ;
        RECT 0.0050 74.2635 0.1580 75.1790 ;
        RECT 8.5550 74.2635 16.5290 75.0830 ;
        RECT 0.0050 74.3630 8.5370 75.0830 ;
        RECT 8.3300 74.2635 16.5290 74.4350 ;
        RECT 0.0050 74.2635 8.3120 75.0830 ;
        RECT 0.0050 74.2635 16.5290 74.3390 ;
        RECT 0.0050 76.3070 16.5290 76.4370 ;
        RECT 16.4120 75.3435 16.5290 76.4370 ;
        RECT 9.3020 76.2110 16.3940 76.4370 ;
        RECT 7.9700 76.2110 9.2840 76.4370 ;
        RECT 7.2500 75.3435 7.8800 76.4370 ;
        RECT 0.1400 76.2110 7.2320 76.4370 ;
        RECT 0.0050 75.3435 0.1220 76.4370 ;
        RECT 16.3760 75.3435 16.5290 76.2590 ;
        RECT 9.3560 75.3435 16.3580 76.4370 ;
        RECT 8.6090 75.3435 9.3380 76.2590 ;
        RECT 8.4470 75.5390 8.5730 76.4370 ;
        RECT 7.1960 75.4430 8.4200 76.2590 ;
        RECT 0.1760 75.3435 7.1780 76.4370 ;
        RECT 0.0050 75.3435 0.1580 76.2590 ;
        RECT 8.5550 75.3435 16.5290 76.1630 ;
        RECT 0.0050 75.4430 8.5370 76.1630 ;
        RECT 8.3300 75.3435 16.5290 75.5150 ;
        RECT 0.0050 75.3435 8.3120 76.1630 ;
        RECT 0.0050 75.3435 16.5290 75.4190 ;
        RECT 0.0050 77.3870 16.5290 77.5170 ;
        RECT 16.4120 76.4235 16.5290 77.5170 ;
        RECT 9.3020 77.2910 16.3940 77.5170 ;
        RECT 7.9700 77.2910 9.2840 77.5170 ;
        RECT 7.2500 76.4235 7.8800 77.5170 ;
        RECT 0.1400 77.2910 7.2320 77.5170 ;
        RECT 0.0050 76.4235 0.1220 77.5170 ;
        RECT 16.3760 76.4235 16.5290 77.3390 ;
        RECT 9.3560 76.4235 16.3580 77.5170 ;
        RECT 8.6090 76.4235 9.3380 77.3390 ;
        RECT 8.4470 76.6190 8.5730 77.5170 ;
        RECT 7.1960 76.5230 8.4200 77.3390 ;
        RECT 0.1760 76.4235 7.1780 77.5170 ;
        RECT 0.0050 76.4235 0.1580 77.3390 ;
        RECT 8.5550 76.4235 16.5290 77.2430 ;
        RECT 0.0050 76.5230 8.5370 77.2430 ;
        RECT 8.3300 76.4235 16.5290 76.5950 ;
        RECT 0.0050 76.4235 8.3120 77.2430 ;
        RECT 0.0050 76.4235 16.5290 76.4990 ;
        RECT 0.0050 78.4670 16.5290 78.5970 ;
        RECT 16.4120 77.5035 16.5290 78.5970 ;
        RECT 9.3020 78.3710 16.3940 78.5970 ;
        RECT 7.9700 78.3710 9.2840 78.5970 ;
        RECT 7.2500 77.5035 7.8800 78.5970 ;
        RECT 0.1400 78.3710 7.2320 78.5970 ;
        RECT 0.0050 77.5035 0.1220 78.5970 ;
        RECT 16.3760 77.5035 16.5290 78.4190 ;
        RECT 9.3560 77.5035 16.3580 78.5970 ;
        RECT 8.6090 77.5035 9.3380 78.4190 ;
        RECT 8.4470 77.6990 8.5730 78.5970 ;
        RECT 7.1960 77.6030 8.4200 78.4190 ;
        RECT 0.1760 77.5035 7.1780 78.5970 ;
        RECT 0.0050 77.5035 0.1580 78.4190 ;
        RECT 8.5550 77.5035 16.5290 78.3230 ;
        RECT 0.0050 77.6030 8.5370 78.3230 ;
        RECT 8.3300 77.5035 16.5290 77.6750 ;
        RECT 0.0050 77.5035 8.3120 78.3230 ;
        RECT 0.0050 77.5035 16.5290 77.5790 ;
        RECT 0.0050 79.5470 16.5290 79.6770 ;
        RECT 16.4120 78.5835 16.5290 79.6770 ;
        RECT 9.3020 79.4510 16.3940 79.6770 ;
        RECT 7.9700 79.4510 9.2840 79.6770 ;
        RECT 7.2500 78.5835 7.8800 79.6770 ;
        RECT 0.1400 79.4510 7.2320 79.6770 ;
        RECT 0.0050 78.5835 0.1220 79.6770 ;
        RECT 16.3760 78.5835 16.5290 79.4990 ;
        RECT 9.3560 78.5835 16.3580 79.6770 ;
        RECT 8.6090 78.5835 9.3380 79.4990 ;
        RECT 8.4470 78.7790 8.5730 79.6770 ;
        RECT 7.1960 78.6830 8.4200 79.4990 ;
        RECT 0.1760 78.5835 7.1780 79.6770 ;
        RECT 0.0050 78.5835 0.1580 79.4990 ;
        RECT 8.5550 78.5835 16.5290 79.4030 ;
        RECT 0.0050 78.6830 8.5370 79.4030 ;
        RECT 8.3300 78.5835 16.5290 78.7550 ;
        RECT 0.0050 78.5835 8.3120 79.4030 ;
        RECT 0.0050 78.5835 16.5290 78.6590 ;
        RECT 0.0050 80.6270 16.5290 80.7570 ;
        RECT 16.4120 79.6635 16.5290 80.7570 ;
        RECT 9.3020 80.5310 16.3940 80.7570 ;
        RECT 7.9700 80.5310 9.2840 80.7570 ;
        RECT 7.2500 79.6635 7.8800 80.7570 ;
        RECT 0.1400 80.5310 7.2320 80.7570 ;
        RECT 0.0050 79.6635 0.1220 80.7570 ;
        RECT 16.3760 79.6635 16.5290 80.5790 ;
        RECT 9.3560 79.6635 16.3580 80.7570 ;
        RECT 8.6090 79.6635 9.3380 80.5790 ;
        RECT 8.4470 79.8590 8.5730 80.7570 ;
        RECT 7.1960 79.7630 8.4200 80.5790 ;
        RECT 0.1760 79.6635 7.1780 80.7570 ;
        RECT 0.0050 79.6635 0.1580 80.5790 ;
        RECT 8.5550 79.6635 16.5290 80.4830 ;
        RECT 0.0050 79.7630 8.5370 80.4830 ;
        RECT 8.3300 79.6635 16.5290 79.8350 ;
        RECT 0.0050 79.6635 8.3120 80.4830 ;
        RECT 0.0050 79.6635 16.5290 79.7390 ;
        RECT 0.0050 81.7070 16.5290 81.8370 ;
        RECT 16.4120 80.7435 16.5290 81.8370 ;
        RECT 9.3020 81.6110 16.3940 81.8370 ;
        RECT 7.9700 81.6110 9.2840 81.8370 ;
        RECT 7.2500 80.7435 7.8800 81.8370 ;
        RECT 0.1400 81.6110 7.2320 81.8370 ;
        RECT 0.0050 80.7435 0.1220 81.8370 ;
        RECT 16.3760 80.7435 16.5290 81.6590 ;
        RECT 9.3560 80.7435 16.3580 81.8370 ;
        RECT 8.6090 80.7435 9.3380 81.6590 ;
        RECT 8.4470 80.9390 8.5730 81.8370 ;
        RECT 7.1960 80.8430 8.4200 81.6590 ;
        RECT 0.1760 80.7435 7.1780 81.8370 ;
        RECT 0.0050 80.7435 0.1580 81.6590 ;
        RECT 8.5550 80.7435 16.5290 81.5630 ;
        RECT 0.0050 80.8430 8.5370 81.5630 ;
        RECT 8.3300 80.7435 16.5290 80.9150 ;
        RECT 0.0050 80.7435 8.3120 81.5630 ;
        RECT 0.0050 80.7435 16.5290 80.8190 ;
        RECT 0.0050 82.7870 16.5290 82.9170 ;
        RECT 16.4120 81.8235 16.5290 82.9170 ;
        RECT 9.3020 82.6910 16.3940 82.9170 ;
        RECT 7.9700 82.6910 9.2840 82.9170 ;
        RECT 7.2500 81.8235 7.8800 82.9170 ;
        RECT 0.1400 82.6910 7.2320 82.9170 ;
        RECT 0.0050 81.8235 0.1220 82.9170 ;
        RECT 16.3760 81.8235 16.5290 82.7390 ;
        RECT 9.3560 81.8235 16.3580 82.9170 ;
        RECT 8.6090 81.8235 9.3380 82.7390 ;
        RECT 8.4470 82.0190 8.5730 82.9170 ;
        RECT 7.1960 81.9230 8.4200 82.7390 ;
        RECT 0.1760 81.8235 7.1780 82.9170 ;
        RECT 0.0050 81.8235 0.1580 82.7390 ;
        RECT 8.5550 81.8235 16.5290 82.6430 ;
        RECT 0.0050 81.9230 8.5370 82.6430 ;
        RECT 8.3300 81.8235 16.5290 81.9950 ;
        RECT 0.0050 81.8235 8.3120 82.6430 ;
        RECT 0.0050 81.8235 16.5290 81.8990 ;
        RECT 0.0050 83.8670 16.5290 83.9970 ;
        RECT 16.4120 82.9035 16.5290 83.9970 ;
        RECT 9.3020 83.7710 16.3940 83.9970 ;
        RECT 7.9700 83.7710 9.2840 83.9970 ;
        RECT 7.2500 82.9035 7.8800 83.9970 ;
        RECT 0.1400 83.7710 7.2320 83.9970 ;
        RECT 0.0050 82.9035 0.1220 83.9970 ;
        RECT 16.3760 82.9035 16.5290 83.8190 ;
        RECT 9.3560 82.9035 16.3580 83.9970 ;
        RECT 8.6090 82.9035 9.3380 83.8190 ;
        RECT 8.4470 83.0990 8.5730 83.9970 ;
        RECT 7.1960 83.0030 8.4200 83.8190 ;
        RECT 0.1760 82.9035 7.1780 83.9970 ;
        RECT 0.0050 82.9035 0.1580 83.8190 ;
        RECT 8.5550 82.9035 16.5290 83.7230 ;
        RECT 0.0050 83.0030 8.5370 83.7230 ;
        RECT 8.3300 82.9035 16.5290 83.0750 ;
        RECT 0.0050 82.9035 8.3120 83.7230 ;
        RECT 0.0050 82.9035 16.5290 82.9790 ;
        RECT 0.0050 84.9470 16.5290 85.0770 ;
        RECT 16.4120 83.9835 16.5290 85.0770 ;
        RECT 9.3020 84.8510 16.3940 85.0770 ;
        RECT 7.9700 84.8510 9.2840 85.0770 ;
        RECT 7.2500 83.9835 7.8800 85.0770 ;
        RECT 0.1400 84.8510 7.2320 85.0770 ;
        RECT 0.0050 83.9835 0.1220 85.0770 ;
        RECT 16.3760 83.9835 16.5290 84.8990 ;
        RECT 9.3560 83.9835 16.3580 85.0770 ;
        RECT 8.6090 83.9835 9.3380 84.8990 ;
        RECT 8.4470 84.1790 8.5730 85.0770 ;
        RECT 7.1960 84.0830 8.4200 84.8990 ;
        RECT 0.1760 83.9835 7.1780 85.0770 ;
        RECT 0.0050 83.9835 0.1580 84.8990 ;
        RECT 8.5550 83.9835 16.5290 84.8030 ;
        RECT 0.0050 84.0830 8.5370 84.8030 ;
        RECT 8.3300 83.9835 16.5290 84.1550 ;
        RECT 0.0050 83.9835 8.3120 84.8030 ;
        RECT 0.0050 83.9835 16.5290 84.0590 ;
        RECT 0.0050 86.0270 16.5290 86.1570 ;
        RECT 16.4120 85.0635 16.5290 86.1570 ;
        RECT 9.3020 85.9310 16.3940 86.1570 ;
        RECT 7.9700 85.9310 9.2840 86.1570 ;
        RECT 7.2500 85.0635 7.8800 86.1570 ;
        RECT 0.1400 85.9310 7.2320 86.1570 ;
        RECT 0.0050 85.0635 0.1220 86.1570 ;
        RECT 16.3760 85.0635 16.5290 85.9790 ;
        RECT 9.3560 85.0635 16.3580 86.1570 ;
        RECT 8.6090 85.0635 9.3380 85.9790 ;
        RECT 8.4470 85.2590 8.5730 86.1570 ;
        RECT 7.1960 85.1630 8.4200 85.9790 ;
        RECT 0.1760 85.0635 7.1780 86.1570 ;
        RECT 0.0050 85.0635 0.1580 85.9790 ;
        RECT 8.5550 85.0635 16.5290 85.8830 ;
        RECT 0.0050 85.1630 8.5370 85.8830 ;
        RECT 8.3300 85.0635 16.5290 85.2350 ;
        RECT 0.0050 85.0635 8.3120 85.8830 ;
        RECT 0.0050 85.0635 16.5290 85.1390 ;
        RECT 0.0050 87.1070 16.5290 87.2370 ;
        RECT 16.4120 86.1435 16.5290 87.2370 ;
        RECT 9.3020 87.0110 16.3940 87.2370 ;
        RECT 7.9700 87.0110 9.2840 87.2370 ;
        RECT 7.2500 86.1435 7.8800 87.2370 ;
        RECT 0.1400 87.0110 7.2320 87.2370 ;
        RECT 0.0050 86.1435 0.1220 87.2370 ;
        RECT 16.3760 86.1435 16.5290 87.0590 ;
        RECT 9.3560 86.1435 16.3580 87.2370 ;
        RECT 8.6090 86.1435 9.3380 87.0590 ;
        RECT 8.4470 86.3390 8.5730 87.2370 ;
        RECT 7.1960 86.2430 8.4200 87.0590 ;
        RECT 0.1760 86.1435 7.1780 87.2370 ;
        RECT 0.0050 86.1435 0.1580 87.0590 ;
        RECT 8.5550 86.1435 16.5290 86.9630 ;
        RECT 0.0050 86.2430 8.5370 86.9630 ;
        RECT 8.3300 86.1435 16.5290 86.3150 ;
        RECT 0.0050 86.1435 8.3120 86.9630 ;
        RECT 0.0050 86.1435 16.5290 86.2190 ;
        RECT 0.0050 88.1870 16.5290 88.3170 ;
        RECT 16.4120 87.2235 16.5290 88.3170 ;
        RECT 9.3020 88.0910 16.3940 88.3170 ;
        RECT 7.9700 88.0910 9.2840 88.3170 ;
        RECT 7.2500 87.2235 7.8800 88.3170 ;
        RECT 0.1400 88.0910 7.2320 88.3170 ;
        RECT 0.0050 87.2235 0.1220 88.3170 ;
        RECT 16.3760 87.2235 16.5290 88.1390 ;
        RECT 9.3560 87.2235 16.3580 88.3170 ;
        RECT 8.6090 87.2235 9.3380 88.1390 ;
        RECT 8.4470 87.4190 8.5730 88.3170 ;
        RECT 7.1960 87.3230 8.4200 88.1390 ;
        RECT 0.1760 87.2235 7.1780 88.3170 ;
        RECT 0.0050 87.2235 0.1580 88.1390 ;
        RECT 8.5550 87.2235 16.5290 88.0430 ;
        RECT 0.0050 87.3230 8.5370 88.0430 ;
        RECT 8.3300 87.2235 16.5290 87.3950 ;
        RECT 0.0050 87.2235 8.3120 88.0430 ;
        RECT 0.0050 87.2235 16.5290 87.2990 ;
  LAYER M4  ;
      RECT 1.5690 41.9100 15.0095 41.9340 ;
      RECT 1.5690 42.1980 15.0095 42.2220 ;
      RECT 1.5690 42.5820 15.0095 42.6060 ;
      RECT 1.5690 42.6780 15.0095 42.7020 ;
      RECT 1.5690 43.0140 15.0095 43.0380 ;
      RECT 1.5690 43.3980 15.0095 43.4220 ;
      RECT 10.9550 40.8690 11.0390 40.8930 ;
      RECT 10.7670 41.3010 10.8970 41.3250 ;
      RECT 10.7750 41.9585 10.8920 41.9825 ;
      RECT 10.7750 42.2460 10.8920 42.2700 ;
      RECT 10.1360 41.3010 10.7070 41.3250 ;
      RECT 10.1960 42.0780 10.3040 42.1020 ;
      RECT 8.8630 42.4530 9.9560 42.4770 ;
      RECT 9.5510 42.0210 9.6350 42.0450 ;
      RECT 8.7670 43.2210 9.6350 43.2450 ;
      RECT 9.5510 43.3170 9.6350 43.3410 ;
      RECT 9.3730 41.5410 9.4570 41.5650 ;
      RECT 9.3350 42.8850 9.4190 42.9090 ;
      RECT 9.3350 43.6050 9.4190 43.6290 ;
      RECT 9.1570 41.4450 9.2410 41.4690 ;
      RECT 8.9430 40.1570 9.2060 40.1810 ;
      RECT 8.9430 48.7810 9.2060 48.8050 ;
      RECT 8.9590 42.9330 9.2030 42.9570 ;
      RECT 9.1190 43.0770 9.2030 43.1010 ;
      RECT 7.6630 43.3170 9.2030 43.3410 ;
      RECT 9.1190 43.6050 9.2030 43.6290 ;
      RECT 8.8850 48.6850 9.1480 48.7090 ;
      RECT 8.8840 40.0610 9.1470 40.0850 ;
      RECT 8.8460 39.9650 9.1090 39.9890 ;
      RECT 8.8460 48.4930 9.1090 48.5170 ;
      RECT 9.0110 44.0370 9.0950 44.0610 ;
      RECT 8.2390 44.4210 9.0950 44.4450 ;
      RECT 8.6230 46.6770 9.0950 46.7010 ;
      RECT 9.0110 46.7730 9.0950 46.7970 ;
      RECT 8.7980 39.8690 9.0610 39.8930 ;
      RECT 8.7980 48.3970 9.0610 48.4210 ;
      RECT 8.5750 45.7650 9.0200 45.7890 ;
      RECT 8.7540 39.7730 9.0170 39.7970 ;
      RECT 8.7540 48.7330 9.0170 48.7570 ;
      RECT 8.7050 40.1090 8.9680 40.1330 ;
      RECT 8.7050 48.6370 8.9680 48.6610 ;
      RECT 8.8360 43.0770 8.9570 43.1010 ;
      RECT 8.8150 45.1890 8.9480 45.2130 ;
      RECT 8.6580 40.0130 8.9210 40.0370 ;
      RECT 8.6580 48.5410 8.9210 48.5650 ;
      RECT 8.6230 39.7250 8.8860 39.7490 ;
      RECT 8.6230 48.4450 8.8860 48.4690 ;
      RECT 7.8070 46.7730 8.8760 46.7970 ;
      RECT 8.7920 47.9250 8.8760 47.9490 ;
      RECT 8.5670 39.5810 8.8300 39.6050 ;
      RECT 8.5670 48.3490 8.8300 48.3730 ;
      RECT 8.7190 44.0370 8.8040 44.0610 ;
      RECT 7.6150 44.6130 8.7320 44.6370 ;
      RECT 8.2600 42.4530 8.7170 42.4770 ;
      RECT 8.0870 40.3010 8.3540 40.3250 ;
      RECT 8.0870 48.2050 8.3540 48.2290 ;
      RECT 8.2240 43.9890 8.3330 44.0130 ;
      RECT 8.0640 40.2050 8.3060 40.2290 ;
      RECT 8.0640 48.8290 8.3060 48.8530 ;
      RECT 8.0080 39.7250 8.2500 39.7490 ;
      RECT 8.0370 48.9250 8.2500 48.9490 ;
      RECT 8.1530 43.6050 8.2370 43.6290 ;
      RECT 7.9540 39.8210 8.2020 39.8450 ;
      RECT 7.9540 48.7810 8.2020 48.8050 ;
      RECT 7.7200 46.1970 8.1410 46.2210 ;
      RECT 7.6880 40.1570 7.9550 40.1810 ;
      RECT 7.6880 48.9250 7.9550 48.9490 ;
      RECT 7.8280 44.7570 7.9490 44.7810 ;
      RECT 7.8200 47.9250 7.9040 47.9490 ;
      RECT 7.6540 40.0610 7.9010 40.0850 ;
      RECT 7.5870 48.4930 7.9010 48.5170 ;
      RECT 7.6280 39.9650 7.8580 39.9890 ;
      RECT 7.6160 48.8290 7.8580 48.8530 ;
      RECT 7.5750 39.8690 7.8050 39.8930 ;
      RECT 7.7210 46.3410 7.8050 46.3650 ;
      RECT 7.5250 48.3970 7.8050 48.4210 ;
      RECT 7.5300 39.7730 7.7600 39.7970 ;
      RECT 7.5300 48.7330 7.7600 48.7570 ;
      RECT 6.5680 43.6050 7.7570 43.6290 ;
      RECT 7.4920 40.0130 7.7220 40.0370 ;
      RECT 7.4920 48.6370 7.7220 48.6610 ;
      RECT 7.4740 39.9170 7.6670 39.9410 ;
      RECT 7.4740 48.5410 7.6670 48.5650 ;
      RECT 7.4250 39.8210 7.6180 39.8450 ;
      RECT 7.4250 48.4450 7.6180 48.4690 ;
      RECT 7.4290 44.5170 7.6130 44.5410 ;
      RECT 7.3730 39.7250 7.5660 39.7490 ;
      RECT 7.3730 48.3490 7.5660 48.3730 ;
      RECT 6.8890 41.8290 7.5650 41.8530 ;
      RECT 7.4290 44.6130 7.5130 44.6370 ;
      RECT 7.1600 40.2530 7.4230 40.2770 ;
      RECT 7.1925 44.0370 7.3260 44.0610 ;
      RECT 6.8510 42.0210 6.9350 42.0450 ;
  LAYER V4  ;
      RECT 11.0040 40.8690 11.0280 40.8930 ;
      RECT 11.0040 41.9100 11.0280 41.9340 ;
      RECT 10.8360 41.3010 10.8600 41.3250 ;
      RECT 10.8360 41.9585 10.8600 41.9825 ;
      RECT 10.8360 42.2460 10.8600 42.2700 ;
      RECT 10.2120 41.3010 10.2360 41.3250 ;
      RECT 10.2120 42.0780 10.2360 42.1020 ;
      RECT 9.6000 42.0210 9.6240 42.0450 ;
      RECT 9.6000 42.1980 9.6240 42.2220 ;
      RECT 9.6000 43.2210 9.6240 43.2450 ;
      RECT 9.6000 43.3170 9.6240 43.3410 ;
      RECT 9.3840 41.5410 9.4080 41.5650 ;
      RECT 9.3840 42.5820 9.4080 42.6060 ;
      RECT 9.3840 42.8850 9.4080 42.9090 ;
      RECT 9.3840 43.0140 9.4080 43.0380 ;
      RECT 9.3840 43.3980 9.4080 43.4220 ;
      RECT 9.3840 43.6050 9.4080 43.6290 ;
      RECT 9.1680 41.4450 9.1920 41.4690 ;
      RECT 9.1680 42.6780 9.1920 42.7020 ;
      RECT 9.1680 42.9330 9.1920 42.9570 ;
      RECT 9.1680 43.0770 9.1920 43.1010 ;
      RECT 9.1680 43.3170 9.1920 43.3410 ;
      RECT 9.1680 43.6050 9.1920 43.6290 ;
      RECT 9.0600 44.0370 9.0840 44.0610 ;
      RECT 9.0600 44.4210 9.0840 44.4450 ;
      RECT 9.0600 46.6770 9.0840 46.7010 ;
      RECT 9.0600 46.7730 9.0840 46.7970 ;
      RECT 8.9700 40.1570 8.9940 40.1810 ;
      RECT 8.9700 42.9330 8.9940 42.9570 ;
      RECT 8.9700 48.7810 8.9940 48.8050 ;
      RECT 8.9220 40.0610 8.9460 40.0850 ;
      RECT 8.9220 43.0770 8.9460 43.1010 ;
      RECT 8.9220 48.6850 8.9460 48.7090 ;
      RECT 8.8740 39.9650 8.8980 39.9890 ;
      RECT 8.8740 42.4530 8.8980 42.4770 ;
      RECT 8.8740 48.4930 8.8980 48.5170 ;
      RECT 8.8260 39.8690 8.8500 39.8930 ;
      RECT 8.8260 45.1890 8.8500 45.2130 ;
      RECT 8.8260 47.9250 8.8500 47.9490 ;
      RECT 8.8260 48.3970 8.8500 48.4210 ;
      RECT 8.7780 39.7730 8.8020 39.7970 ;
      RECT 8.7780 43.2210 8.8020 43.2450 ;
      RECT 8.7780 48.7330 8.8020 48.7570 ;
      RECT 8.7300 40.1090 8.7540 40.1330 ;
      RECT 8.7300 44.0370 8.7540 44.0610 ;
      RECT 8.7300 48.6370 8.7540 48.6610 ;
      RECT 8.6820 40.0130 8.7060 40.0370 ;
      RECT 8.6820 42.4530 8.7060 42.4770 ;
      RECT 8.6820 48.5410 8.7060 48.5650 ;
      RECT 8.6340 39.7250 8.6580 39.7490 ;
      RECT 8.6340 46.6770 8.6580 46.7010 ;
      RECT 8.6340 48.4450 8.6580 48.4690 ;
      RECT 8.5860 39.5810 8.6100 39.6050 ;
      RECT 8.5860 45.7650 8.6100 45.7890 ;
      RECT 8.5860 48.3490 8.6100 48.3730 ;
      RECT 8.2980 40.3010 8.3220 40.3250 ;
      RECT 8.2980 43.9890 8.3220 44.0130 ;
      RECT 8.2980 48.2050 8.3220 48.2290 ;
      RECT 8.2500 40.2050 8.2740 40.2290 ;
      RECT 8.2500 44.4210 8.2740 44.4450 ;
      RECT 8.2500 48.8290 8.2740 48.8530 ;
      RECT 8.2020 39.7250 8.2260 39.7490 ;
      RECT 8.2020 43.6050 8.2260 43.6290 ;
      RECT 8.2020 48.9250 8.2260 48.9490 ;
      RECT 8.1060 39.8210 8.1300 39.8450 ;
      RECT 8.1060 46.1970 8.1300 46.2210 ;
      RECT 8.1060 48.7810 8.1300 48.8050 ;
      RECT 7.9140 40.1570 7.9380 40.1810 ;
      RECT 7.9140 44.7570 7.9380 44.7810 ;
      RECT 7.9140 48.9250 7.9380 48.9490 ;
      RECT 7.8660 40.0610 7.8900 40.0850 ;
      RECT 7.8660 47.9250 7.8900 47.9490 ;
      RECT 7.8660 48.4930 7.8900 48.5170 ;
      RECT 7.8180 39.9650 7.8420 39.9890 ;
      RECT 7.8180 46.7730 7.8420 46.7970 ;
      RECT 7.8180 48.8290 7.8420 48.8530 ;
      RECT 7.7700 39.8690 7.7940 39.8930 ;
      RECT 7.7700 46.3410 7.7940 46.3650 ;
      RECT 7.7700 48.3970 7.7940 48.4210 ;
      RECT 7.7220 39.7730 7.7460 39.7970 ;
      RECT 7.7220 43.6050 7.7460 43.6290 ;
      RECT 7.7220 48.7330 7.7460 48.7570 ;
      RECT 7.6740 40.0130 7.6980 40.0370 ;
      RECT 7.6740 43.3170 7.6980 43.3410 ;
      RECT 7.6740 48.6370 7.6980 48.6610 ;
      RECT 7.6260 39.9170 7.6500 39.9410 ;
      RECT 7.6260 44.6130 7.6500 44.6370 ;
      RECT 7.6260 48.5410 7.6500 48.5650 ;
      RECT 7.5780 39.8210 7.6020 39.8450 ;
      RECT 7.5780 44.5170 7.6020 44.5410 ;
      RECT 7.5780 48.4450 7.6020 48.4690 ;
      RECT 7.5300 39.7250 7.5540 39.7490 ;
      RECT 7.5300 41.8290 7.5540 41.8530 ;
      RECT 7.5300 48.3490 7.5540 48.3730 ;
      RECT 7.4400 44.5170 7.4640 44.5410 ;
      RECT 7.4400 44.6130 7.4640 44.6370 ;
      RECT 7.2720 40.2530 7.2960 40.2770 ;
      RECT 7.2720 44.0370 7.2960 44.0610 ;
      RECT 6.9000 41.8290 6.9240 41.8530 ;
      RECT 6.9000 42.0210 6.9240 42.0450 ;
  LAYER M5  ;
      RECT 11.0040 40.8580 11.0280 41.9450 ;
      RECT 10.8360 41.2730 10.8600 42.3335 ;
      RECT 10.2120 41.2815 10.2360 42.1140 ;
      RECT 9.6000 42.0100 9.6240 42.2330 ;
      RECT 9.6000 43.2100 9.6240 43.3520 ;
      RECT 9.3840 41.5300 9.4080 42.6170 ;
      RECT 9.3840 42.8740 9.4080 43.0490 ;
      RECT 9.3840 43.3870 9.4080 43.6400 ;
      RECT 9.1680 41.4340 9.1920 42.7130 ;
      RECT 9.1680 42.9220 9.1920 43.1120 ;
      RECT 9.1680 43.3060 9.1920 43.6400 ;
      RECT 9.0600 44.0260 9.0840 44.4560 ;
      RECT 9.0600 46.6660 9.0840 46.8080 ;
      RECT 8.9700 40.4940 8.9940 48.0770 ;
      RECT 8.9220 40.4940 8.9460 48.0770 ;
      RECT 8.8740 40.4940 8.8980 48.0770 ;
      RECT 8.8260 40.4940 8.8500 48.0770 ;
      RECT 8.7780 40.4940 8.8020 48.0770 ;
      RECT 8.7300 40.4940 8.7540 48.0770 ;
      RECT 8.6820 40.4940 8.7060 48.0770 ;
      RECT 8.6340 40.4940 8.6580 48.0770 ;
      RECT 8.5860 40.4940 8.6100 48.0770 ;
      RECT 8.2980 40.4940 8.3220 48.0770 ;
      RECT 8.2500 40.4940 8.2740 48.0770 ;
      RECT 8.2020 40.4940 8.2260 48.0770 ;
      RECT 8.1060 40.4940 8.1300 48.0770 ;
      RECT 7.9140 40.4940 7.9380 48.0770 ;
      RECT 7.8660 40.4940 7.8900 48.0770 ;
      RECT 7.8180 40.4940 7.8420 48.0770 ;
      RECT 7.7700 40.4940 7.7940 48.0770 ;
      RECT 7.7220 40.4940 7.7460 48.0770 ;
      RECT 7.6740 40.4940 7.6980 48.0770 ;
      RECT 7.6260 39.6520 7.6500 48.7070 ;
      RECT 7.5780 39.6150 7.6020 48.6610 ;
      RECT 7.5300 39.5610 7.5540 48.6070 ;
      RECT 7.4400 44.5060 7.4640 44.6480 ;
      RECT 7.2720 40.2350 7.2960 44.0790 ;
      RECT 6.9000 41.8180 6.9240 42.0560 ;
  LAYER M2  ;
    RECT 0.108 0.036 15.8920 88.5240 ;
  LAYER M1  ;
    RECT 0.108 0.036 15.8920 88.5240 ;
  END
END srambank_128x4x74_6t122 
