VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_64x4x16_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_64x4x16_6t122 0 0 ;
  SIZE 9.612 BY 25.92 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1010 1.1720 9.5090 1.2200 ;
        RECT 0.1010 2.2520 9.5090 2.3000 ;
        RECT 0.1010 3.3320 9.5090 3.3800 ;
        RECT 0.1010 4.4120 9.5090 4.4600 ;
        RECT 0.1010 5.4920 9.5090 5.5400 ;
        RECT 0.1010 6.5720 9.5090 6.6200 ;
        RECT 0.1010 7.6520 9.5090 7.7000 ;
        RECT 0.1010 8.7320 9.5090 8.7800 ;
        RECT 0.1080 9.2190 9.5040 9.4350 ;
        RECT 5.6100 8.9390 5.8730 8.9630 ;
        RECT 5.7410 12.7230 5.8530 12.7470 ;
        RECT 3.9420 12.3870 5.6700 12.6030 ;
        RECT 3.9420 15.5550 5.6700 15.7710 ;
        RECT 0.1010 17.9390 9.5090 17.9870 ;
        RECT 0.1010 19.0190 9.5090 19.0670 ;
        RECT 0.1010 20.0990 9.5090 20.1470 ;
        RECT 0.1010 21.1790 9.5090 21.2270 ;
        RECT 0.1010 22.2590 9.5090 22.3070 ;
        RECT 0.1010 23.3390 9.5090 23.3870 ;
        RECT 0.1010 24.4190 9.5090 24.4670 ;
        RECT 0.1010 25.4990 9.5090 25.5470 ;
      LAYER M3  ;
        RECT 9.4770 0.2165 9.4950 1.3765 ;
        RECT 5.8230 0.2170 5.8410 1.3760 ;
        RECT 4.4190 0.2530 4.5090 1.3670 ;
        RECT 3.7710 0.2170 3.7890 1.3760 ;
        RECT 0.1170 0.2165 0.1350 1.3765 ;
        RECT 9.4770 1.2965 9.4950 2.4565 ;
        RECT 5.8230 1.2970 5.8410 2.4560 ;
        RECT 4.4190 1.3330 4.5090 2.4470 ;
        RECT 3.7710 1.2970 3.7890 2.4560 ;
        RECT 0.1170 1.2965 0.1350 2.4565 ;
        RECT 9.4770 2.3765 9.4950 3.5365 ;
        RECT 5.8230 2.3770 5.8410 3.5360 ;
        RECT 4.4190 2.4130 4.5090 3.5270 ;
        RECT 3.7710 2.3770 3.7890 3.5360 ;
        RECT 0.1170 2.3765 0.1350 3.5365 ;
        RECT 9.4770 3.4565 9.4950 4.6165 ;
        RECT 5.8230 3.4570 5.8410 4.6160 ;
        RECT 4.4190 3.4930 4.5090 4.6070 ;
        RECT 3.7710 3.4570 3.7890 4.6160 ;
        RECT 0.1170 3.4565 0.1350 4.6165 ;
        RECT 9.4770 4.5365 9.4950 5.6965 ;
        RECT 5.8230 4.5370 5.8410 5.6960 ;
        RECT 4.4190 4.5730 4.5090 5.6870 ;
        RECT 3.7710 4.5370 3.7890 5.6960 ;
        RECT 0.1170 4.5365 0.1350 5.6965 ;
        RECT 9.4770 5.6165 9.4950 6.7765 ;
        RECT 5.8230 5.6170 5.8410 6.7760 ;
        RECT 4.4190 5.6530 4.5090 6.7670 ;
        RECT 3.7710 5.6170 3.7890 6.7760 ;
        RECT 0.1170 5.6165 0.1350 6.7765 ;
        RECT 9.4770 6.6965 9.4950 7.8565 ;
        RECT 5.8230 6.6970 5.8410 7.8560 ;
        RECT 4.4190 6.7330 4.5090 7.8470 ;
        RECT 3.7710 6.6970 3.7890 7.8560 ;
        RECT 0.1170 6.6965 0.1350 7.8565 ;
        RECT 9.4770 7.7765 9.4950 8.9365 ;
        RECT 5.8230 7.7770 5.8410 8.9360 ;
        RECT 4.4190 7.8130 4.5090 8.9270 ;
        RECT 3.7710 7.7770 3.7890 8.9360 ;
        RECT 0.1170 7.7765 0.1350 8.9365 ;
        RECT 9.4770 8.8565 9.4950 17.0635 ;
        RECT 5.8230 8.9360 5.8410 9.0275 ;
        RECT 5.8230 12.6760 5.8410 17.0360 ;
        RECT 4.4550 9.1800 4.6890 16.7630 ;
        RECT 4.4190 16.6770 4.5090 17.2120 ;
        RECT 4.4190 8.9000 4.5090 9.4350 ;
        RECT 0.1170 8.8565 0.1350 17.0635 ;
        RECT 9.4770 16.9835 9.4950 18.1435 ;
        RECT 5.8230 16.9840 5.8410 18.1430 ;
        RECT 4.4190 17.0200 4.5090 18.1340 ;
        RECT 3.7710 16.9840 3.7890 18.1430 ;
        RECT 0.1170 16.9835 0.1350 18.1435 ;
        RECT 9.4770 18.0635 9.4950 19.2235 ;
        RECT 5.8230 18.0640 5.8410 19.2230 ;
        RECT 4.4190 18.1000 4.5090 19.2140 ;
        RECT 3.7710 18.0640 3.7890 19.2230 ;
        RECT 0.1170 18.0635 0.1350 19.2235 ;
        RECT 9.4770 19.1435 9.4950 20.3035 ;
        RECT 5.8230 19.1440 5.8410 20.3030 ;
        RECT 4.4190 19.1800 4.5090 20.2940 ;
        RECT 3.7710 19.1440 3.7890 20.3030 ;
        RECT 0.1170 19.1435 0.1350 20.3035 ;
        RECT 9.4770 20.2235 9.4950 21.3835 ;
        RECT 5.8230 20.2240 5.8410 21.3830 ;
        RECT 4.4190 20.2600 4.5090 21.3740 ;
        RECT 3.7710 20.2240 3.7890 21.3830 ;
        RECT 0.1170 20.2235 0.1350 21.3835 ;
        RECT 9.4770 21.3035 9.4950 22.4635 ;
        RECT 5.8230 21.3040 5.8410 22.4630 ;
        RECT 4.4190 21.3400 4.5090 22.4540 ;
        RECT 3.7710 21.3040 3.7890 22.4630 ;
        RECT 0.1170 21.3035 0.1350 22.4635 ;
        RECT 9.4770 22.3835 9.4950 23.5435 ;
        RECT 5.8230 22.3840 5.8410 23.5430 ;
        RECT 4.4190 22.4200 4.5090 23.5340 ;
        RECT 3.7710 22.3840 3.7890 23.5430 ;
        RECT 0.1170 22.3835 0.1350 23.5435 ;
        RECT 9.4770 23.4635 9.4950 24.6235 ;
        RECT 5.8230 23.4640 5.8410 24.6230 ;
        RECT 4.4190 23.5000 4.5090 24.6140 ;
        RECT 3.7710 23.4640 3.7890 24.6230 ;
        RECT 0.1170 23.4635 0.1350 24.6235 ;
        RECT 9.4770 24.5435 9.4950 25.7035 ;
        RECT 5.8230 24.5440 5.8410 25.7030 ;
        RECT 4.4190 24.5800 4.5090 25.6940 ;
        RECT 3.7710 24.5440 3.7890 25.7030 ;
        RECT 0.1170 24.5435 0.1350 25.7035 ;
      LAYER V3  ;
        RECT 0.1170 1.1720 0.1350 1.2200 ;
        RECT 3.7710 1.1720 3.7890 1.2200 ;
        RECT 4.4190 1.1720 4.5090 1.2200 ;
        RECT 5.8230 1.1720 5.8410 1.2200 ;
        RECT 9.4770 1.1720 9.4950 1.2200 ;
        RECT 0.1170 2.2520 0.1350 2.3000 ;
        RECT 3.7710 2.2520 3.7890 2.3000 ;
        RECT 4.4190 2.2520 4.5090 2.3000 ;
        RECT 5.8230 2.2520 5.8410 2.3000 ;
        RECT 9.4770 2.2520 9.4950 2.3000 ;
        RECT 0.1170 3.3320 0.1350 3.3800 ;
        RECT 3.7710 3.3320 3.7890 3.3800 ;
        RECT 4.4190 3.3320 4.5090 3.3800 ;
        RECT 5.8230 3.3320 5.8410 3.3800 ;
        RECT 9.4770 3.3320 9.4950 3.3800 ;
        RECT 0.1170 4.4120 0.1350 4.4600 ;
        RECT 3.7710 4.4120 3.7890 4.4600 ;
        RECT 4.4190 4.4120 4.5090 4.4600 ;
        RECT 5.8230 4.4120 5.8410 4.4600 ;
        RECT 9.4770 4.4120 9.4950 4.4600 ;
        RECT 0.1170 5.4920 0.1350 5.5400 ;
        RECT 3.7710 5.4920 3.7890 5.5400 ;
        RECT 4.4190 5.4920 4.5090 5.5400 ;
        RECT 5.8230 5.4920 5.8410 5.5400 ;
        RECT 9.4770 5.4920 9.4950 5.5400 ;
        RECT 0.1170 6.5720 0.1350 6.6200 ;
        RECT 3.7710 6.5720 3.7890 6.6200 ;
        RECT 4.4190 6.5720 4.5090 6.6200 ;
        RECT 5.8230 6.5720 5.8410 6.6200 ;
        RECT 9.4770 6.5720 9.4950 6.6200 ;
        RECT 0.1170 7.6520 0.1350 7.7000 ;
        RECT 3.7710 7.6520 3.7890 7.7000 ;
        RECT 4.4190 7.6520 4.5090 7.7000 ;
        RECT 5.8230 7.6520 5.8410 7.7000 ;
        RECT 9.4770 7.6520 9.4950 7.7000 ;
        RECT 0.1170 8.7320 0.1350 8.7800 ;
        RECT 3.7710 8.7320 3.7890 8.7800 ;
        RECT 4.4190 8.7320 4.5090 8.7800 ;
        RECT 5.8230 8.7320 5.8410 8.7800 ;
        RECT 9.4770 8.7320 9.4950 8.7800 ;
        RECT 0.1170 9.2190 0.1350 9.4350 ;
        RECT 4.4590 15.5550 4.4770 15.7710 ;
        RECT 4.4590 12.3870 4.4770 12.6030 ;
        RECT 4.4590 9.2190 4.4770 9.4350 ;
        RECT 4.5110 15.5550 4.5290 15.7710 ;
        RECT 4.5110 12.3870 4.5290 12.6030 ;
        RECT 4.5110 9.2190 4.5290 9.4350 ;
        RECT 4.5630 15.5550 4.5810 15.7710 ;
        RECT 4.5630 12.3870 4.5810 12.6030 ;
        RECT 4.5630 9.2190 4.5810 9.4350 ;
        RECT 4.6150 15.5550 4.6330 15.7710 ;
        RECT 4.6150 12.3870 4.6330 12.6030 ;
        RECT 4.6150 9.2190 4.6330 9.4350 ;
        RECT 4.6670 15.5550 4.6850 15.7710 ;
        RECT 4.6670 12.3870 4.6850 12.6030 ;
        RECT 4.6670 9.2190 4.6850 9.4350 ;
        RECT 5.8230 12.7230 5.8410 12.7470 ;
        RECT 5.8230 8.9390 5.8410 8.9630 ;
        RECT 0.1170 17.9390 0.1350 17.9870 ;
        RECT 3.7710 17.9390 3.7890 17.9870 ;
        RECT 4.4190 17.9390 4.5090 17.9870 ;
        RECT 5.8230 17.9390 5.8410 17.9870 ;
        RECT 9.4770 17.9390 9.4950 17.9870 ;
        RECT 0.1170 19.0190 0.1350 19.0670 ;
        RECT 3.7710 19.0190 3.7890 19.0670 ;
        RECT 4.4190 19.0190 4.5090 19.0670 ;
        RECT 5.8230 19.0190 5.8410 19.0670 ;
        RECT 9.4770 19.0190 9.4950 19.0670 ;
        RECT 0.1170 20.0990 0.1350 20.1470 ;
        RECT 3.7710 20.0990 3.7890 20.1470 ;
        RECT 4.4190 20.0990 4.5090 20.1470 ;
        RECT 5.8230 20.0990 5.8410 20.1470 ;
        RECT 9.4770 20.0990 9.4950 20.1470 ;
        RECT 0.1170 21.1790 0.1350 21.2270 ;
        RECT 3.7710 21.1790 3.7890 21.2270 ;
        RECT 4.4190 21.1790 4.5090 21.2270 ;
        RECT 5.8230 21.1790 5.8410 21.2270 ;
        RECT 9.4770 21.1790 9.4950 21.2270 ;
        RECT 0.1170 22.2590 0.1350 22.3070 ;
        RECT 3.7710 22.2590 3.7890 22.3070 ;
        RECT 4.4190 22.2590 4.5090 22.3070 ;
        RECT 5.8230 22.2590 5.8410 22.3070 ;
        RECT 9.4770 22.2590 9.4950 22.3070 ;
        RECT 0.1170 23.3390 0.1350 23.3870 ;
        RECT 3.7710 23.3390 3.7890 23.3870 ;
        RECT 4.4190 23.3390 4.5090 23.3870 ;
        RECT 5.8230 23.3390 5.8410 23.3870 ;
        RECT 9.4770 23.3390 9.4950 23.3870 ;
        RECT 0.1170 24.4190 0.1350 24.4670 ;
        RECT 3.7710 24.4190 3.7890 24.4670 ;
        RECT 4.4190 24.4190 4.5090 24.4670 ;
        RECT 5.8230 24.4190 5.8410 24.4670 ;
        RECT 9.4770 24.4190 9.4950 24.4670 ;
        RECT 0.1170 25.4990 0.1350 25.5470 ;
        RECT 3.7710 25.4990 3.7890 25.5470 ;
        RECT 4.4190 25.4990 4.5090 25.5470 ;
        RECT 5.8230 25.4990 5.8410 25.5470 ;
        RECT 9.4770 25.4990 9.4950 25.5470 ;
      LAYER M5  ;
        RECT 5.7590 8.9210 5.7830 12.7650 ;
      LAYER V4  ;
        RECT 5.7590 12.7230 5.7830 12.7470 ;
        RECT 5.7590 8.9390 5.7830 8.9630 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1010 1.0760 9.5040 1.1240 ;
        RECT 0.1010 2.1560 9.5040 2.2040 ;
        RECT 0.1010 3.2360 9.5040 3.2840 ;
        RECT 0.1010 4.3160 9.5040 4.3640 ;
        RECT 0.1010 5.3960 9.5040 5.4440 ;
        RECT 0.1010 6.4760 9.5040 6.5240 ;
        RECT 0.1010 7.5560 9.5040 7.6040 ;
        RECT 0.1010 8.6360 9.5040 8.6840 ;
        RECT 0.1080 9.6510 9.5040 9.8670 ;
        RECT 3.9420 12.8190 5.6700 13.0350 ;
        RECT 3.9420 15.9870 5.6700 16.2030 ;
        RECT 0.1010 17.8430 9.5040 17.8910 ;
        RECT 0.1010 18.9230 9.5040 18.9710 ;
        RECT 0.1010 20.0030 9.5040 20.0510 ;
        RECT 0.1010 21.0830 9.5040 21.1310 ;
        RECT 0.1010 22.1630 9.5040 22.2110 ;
        RECT 0.1010 23.2430 9.5040 23.2910 ;
        RECT 0.1010 24.3230 9.5040 24.3710 ;
        RECT 0.1010 25.4030 9.5040 25.4510 ;
      LAYER M3  ;
        RECT 9.4410 0.2165 9.4590 1.3765 ;
        RECT 5.8770 0.2165 5.8950 1.3765 ;
        RECT 5.1120 0.2530 5.1480 1.3670 ;
        RECT 4.9590 0.2530 4.9860 1.3670 ;
        RECT 3.7170 0.2165 3.7350 1.3765 ;
        RECT 0.1530 0.2165 0.1710 1.3765 ;
        RECT 9.4410 1.2965 9.4590 2.4565 ;
        RECT 5.8770 1.2965 5.8950 2.4565 ;
        RECT 5.1120 1.3330 5.1480 2.4470 ;
        RECT 4.9590 1.3330 4.9860 2.4470 ;
        RECT 3.7170 1.2965 3.7350 2.4565 ;
        RECT 0.1530 1.2965 0.1710 2.4565 ;
        RECT 9.4410 2.3765 9.4590 3.5365 ;
        RECT 5.8770 2.3765 5.8950 3.5365 ;
        RECT 5.1120 2.4130 5.1480 3.5270 ;
        RECT 4.9590 2.4130 4.9860 3.5270 ;
        RECT 3.7170 2.3765 3.7350 3.5365 ;
        RECT 0.1530 2.3765 0.1710 3.5365 ;
        RECT 9.4410 3.4565 9.4590 4.6165 ;
        RECT 5.8770 3.4565 5.8950 4.6165 ;
        RECT 5.1120 3.4930 5.1480 4.6070 ;
        RECT 4.9590 3.4930 4.9860 4.6070 ;
        RECT 3.7170 3.4565 3.7350 4.6165 ;
        RECT 0.1530 3.4565 0.1710 4.6165 ;
        RECT 9.4410 4.5365 9.4590 5.6965 ;
        RECT 5.8770 4.5365 5.8950 5.6965 ;
        RECT 5.1120 4.5730 5.1480 5.6870 ;
        RECT 4.9590 4.5730 4.9860 5.6870 ;
        RECT 3.7170 4.5365 3.7350 5.6965 ;
        RECT 0.1530 4.5365 0.1710 5.6965 ;
        RECT 9.4410 5.6165 9.4590 6.7765 ;
        RECT 5.8770 5.6165 5.8950 6.7765 ;
        RECT 5.1120 5.6530 5.1480 6.7670 ;
        RECT 4.9590 5.6530 4.9860 6.7670 ;
        RECT 3.7170 5.6165 3.7350 6.7765 ;
        RECT 0.1530 5.6165 0.1710 6.7765 ;
        RECT 9.4410 6.6965 9.4590 7.8565 ;
        RECT 5.8770 6.6965 5.8950 7.8565 ;
        RECT 5.1120 6.7330 5.1480 7.8470 ;
        RECT 4.9590 6.7330 4.9860 7.8470 ;
        RECT 3.7170 6.6965 3.7350 7.8565 ;
        RECT 0.1530 6.6965 0.1710 7.8565 ;
        RECT 9.4410 7.7765 9.4590 8.9365 ;
        RECT 5.8770 7.7765 5.8950 8.9365 ;
        RECT 5.1120 7.8130 5.1480 8.9270 ;
        RECT 4.9590 7.8130 4.9860 8.9270 ;
        RECT 3.7170 7.7765 3.7350 8.9365 ;
        RECT 0.1530 7.7765 0.1710 8.9365 ;
        RECT 9.4410 8.8565 9.4590 17.0635 ;
        RECT 5.8770 8.8565 5.8950 17.0635 ;
        RECT 4.9230 9.0800 5.1570 16.7630 ;
        RECT 5.1120 8.9000 5.1480 17.0370 ;
        RECT 4.9590 8.9000 4.9860 17.0340 ;
        RECT 3.7170 8.8565 3.7350 17.0635 ;
        RECT 0.1530 8.8565 0.1710 17.0635 ;
        RECT 9.4410 16.9835 9.4590 18.1435 ;
        RECT 5.8770 16.9835 5.8950 18.1435 ;
        RECT 5.1120 17.0200 5.1480 18.1340 ;
        RECT 4.9590 17.0200 4.9860 18.1340 ;
        RECT 3.7170 16.9835 3.7350 18.1435 ;
        RECT 0.1530 16.9835 0.1710 18.1435 ;
        RECT 9.4410 18.0635 9.4590 19.2235 ;
        RECT 5.8770 18.0635 5.8950 19.2235 ;
        RECT 5.1120 18.1000 5.1480 19.2140 ;
        RECT 4.9590 18.1000 4.9860 19.2140 ;
        RECT 3.7170 18.0635 3.7350 19.2235 ;
        RECT 0.1530 18.0635 0.1710 19.2235 ;
        RECT 9.4410 19.1435 9.4590 20.3035 ;
        RECT 5.8770 19.1435 5.8950 20.3035 ;
        RECT 5.1120 19.1800 5.1480 20.2940 ;
        RECT 4.9590 19.1800 4.9860 20.2940 ;
        RECT 3.7170 19.1435 3.7350 20.3035 ;
        RECT 0.1530 19.1435 0.1710 20.3035 ;
        RECT 9.4410 20.2235 9.4590 21.3835 ;
        RECT 5.8770 20.2235 5.8950 21.3835 ;
        RECT 5.1120 20.2600 5.1480 21.3740 ;
        RECT 4.9590 20.2600 4.9860 21.3740 ;
        RECT 3.7170 20.2235 3.7350 21.3835 ;
        RECT 0.1530 20.2235 0.1710 21.3835 ;
        RECT 9.4410 21.3035 9.4590 22.4635 ;
        RECT 5.8770 21.3035 5.8950 22.4635 ;
        RECT 5.1120 21.3400 5.1480 22.4540 ;
        RECT 4.9590 21.3400 4.9860 22.4540 ;
        RECT 3.7170 21.3035 3.7350 22.4635 ;
        RECT 0.1530 21.3035 0.1710 22.4635 ;
        RECT 9.4410 22.3835 9.4590 23.5435 ;
        RECT 5.8770 22.3835 5.8950 23.5435 ;
        RECT 5.1120 22.4200 5.1480 23.5340 ;
        RECT 4.9590 22.4200 4.9860 23.5340 ;
        RECT 3.7170 22.3835 3.7350 23.5435 ;
        RECT 0.1530 22.3835 0.1710 23.5435 ;
        RECT 9.4410 23.4635 9.4590 24.6235 ;
        RECT 5.8770 23.4635 5.8950 24.6235 ;
        RECT 5.1120 23.5000 5.1480 24.6140 ;
        RECT 4.9590 23.5000 4.9860 24.6140 ;
        RECT 3.7170 23.4635 3.7350 24.6235 ;
        RECT 0.1530 23.4635 0.1710 24.6235 ;
        RECT 9.4410 24.5435 9.4590 25.7035 ;
        RECT 5.8770 24.5435 5.8950 25.7035 ;
        RECT 5.1120 24.5800 5.1480 25.6940 ;
        RECT 4.9590 24.5800 4.9860 25.6940 ;
        RECT 3.7170 24.5435 3.7350 25.7035 ;
        RECT 0.1530 24.5435 0.1710 25.7035 ;
      LAYER V3  ;
        RECT 0.1530 1.0760 0.1710 1.1240 ;
        RECT 3.7170 1.0760 3.7350 1.1240 ;
        RECT 4.9590 1.0760 4.9860 1.1240 ;
        RECT 5.1120 1.0760 5.1480 1.1240 ;
        RECT 5.8770 1.0760 5.8950 1.1240 ;
        RECT 9.4410 1.0760 9.4590 1.1240 ;
        RECT 0.1530 2.1560 0.1710 2.2040 ;
        RECT 3.7170 2.1560 3.7350 2.2040 ;
        RECT 4.9590 2.1560 4.9860 2.2040 ;
        RECT 5.1120 2.1560 5.1480 2.2040 ;
        RECT 5.8770 2.1560 5.8950 2.2040 ;
        RECT 9.4410 2.1560 9.4590 2.2040 ;
        RECT 0.1530 3.2360 0.1710 3.2840 ;
        RECT 3.7170 3.2360 3.7350 3.2840 ;
        RECT 4.9590 3.2360 4.9860 3.2840 ;
        RECT 5.1120 3.2360 5.1480 3.2840 ;
        RECT 5.8770 3.2360 5.8950 3.2840 ;
        RECT 9.4410 3.2360 9.4590 3.2840 ;
        RECT 0.1530 4.3160 0.1710 4.3640 ;
        RECT 3.7170 4.3160 3.7350 4.3640 ;
        RECT 4.9590 4.3160 4.9860 4.3640 ;
        RECT 5.1120 4.3160 5.1480 4.3640 ;
        RECT 5.8770 4.3160 5.8950 4.3640 ;
        RECT 9.4410 4.3160 9.4590 4.3640 ;
        RECT 0.1530 5.3960 0.1710 5.4440 ;
        RECT 3.7170 5.3960 3.7350 5.4440 ;
        RECT 4.9590 5.3960 4.9860 5.4440 ;
        RECT 5.1120 5.3960 5.1480 5.4440 ;
        RECT 5.8770 5.3960 5.8950 5.4440 ;
        RECT 9.4410 5.3960 9.4590 5.4440 ;
        RECT 0.1530 6.4760 0.1710 6.5240 ;
        RECT 3.7170 6.4760 3.7350 6.5240 ;
        RECT 4.9590 6.4760 4.9860 6.5240 ;
        RECT 5.1120 6.4760 5.1480 6.5240 ;
        RECT 5.8770 6.4760 5.8950 6.5240 ;
        RECT 9.4410 6.4760 9.4590 6.5240 ;
        RECT 0.1530 7.5560 0.1710 7.6040 ;
        RECT 3.7170 7.5560 3.7350 7.6040 ;
        RECT 4.9590 7.5560 4.9860 7.6040 ;
        RECT 5.1120 7.5560 5.1480 7.6040 ;
        RECT 5.8770 7.5560 5.8950 7.6040 ;
        RECT 9.4410 7.5560 9.4590 7.6040 ;
        RECT 0.1530 8.6360 0.1710 8.6840 ;
        RECT 3.7170 8.6360 3.7350 8.6840 ;
        RECT 4.9590 8.6360 4.9860 8.6840 ;
        RECT 5.1120 8.6360 5.1480 8.6840 ;
        RECT 5.8770 8.6360 5.8950 8.6840 ;
        RECT 9.4410 8.6360 9.4590 8.6840 ;
        RECT 0.1530 9.6510 0.1710 9.8670 ;
        RECT 4.9270 15.9870 4.9450 16.2030 ;
        RECT 4.9270 12.8190 4.9450 13.0350 ;
        RECT 4.9270 9.6510 4.9450 9.8670 ;
        RECT 4.9790 15.9870 4.9970 16.2030 ;
        RECT 4.9790 12.8190 4.9970 13.0350 ;
        RECT 4.9790 9.6510 4.9970 9.8670 ;
        RECT 5.0310 15.9870 5.0490 16.2030 ;
        RECT 5.0310 12.8190 5.0490 13.0350 ;
        RECT 5.0310 9.6510 5.0490 9.8670 ;
        RECT 5.0830 15.9870 5.1010 16.2030 ;
        RECT 5.0830 12.8190 5.1010 13.0350 ;
        RECT 5.0830 9.6510 5.1010 9.8670 ;
        RECT 5.1350 15.9870 5.1530 16.2030 ;
        RECT 5.1350 12.8190 5.1530 13.0350 ;
        RECT 5.1350 9.6510 5.1530 9.8670 ;
        RECT 0.1530 17.8430 0.1710 17.8910 ;
        RECT 3.7170 17.8430 3.7350 17.8910 ;
        RECT 4.9590 17.8430 4.9860 17.8910 ;
        RECT 5.1120 17.8430 5.1480 17.8910 ;
        RECT 5.8770 17.8430 5.8950 17.8910 ;
        RECT 9.4410 17.8430 9.4590 17.8910 ;
        RECT 0.1530 18.9230 0.1710 18.9710 ;
        RECT 3.7170 18.9230 3.7350 18.9710 ;
        RECT 4.9590 18.9230 4.9860 18.9710 ;
        RECT 5.1120 18.9230 5.1480 18.9710 ;
        RECT 5.8770 18.9230 5.8950 18.9710 ;
        RECT 9.4410 18.9230 9.4590 18.9710 ;
        RECT 0.1530 20.0030 0.1710 20.0510 ;
        RECT 3.7170 20.0030 3.7350 20.0510 ;
        RECT 4.9590 20.0030 4.9860 20.0510 ;
        RECT 5.1120 20.0030 5.1480 20.0510 ;
        RECT 5.8770 20.0030 5.8950 20.0510 ;
        RECT 9.4410 20.0030 9.4590 20.0510 ;
        RECT 0.1530 21.0830 0.1710 21.1310 ;
        RECT 3.7170 21.0830 3.7350 21.1310 ;
        RECT 4.9590 21.0830 4.9860 21.1310 ;
        RECT 5.1120 21.0830 5.1480 21.1310 ;
        RECT 5.8770 21.0830 5.8950 21.1310 ;
        RECT 9.4410 21.0830 9.4590 21.1310 ;
        RECT 0.1530 22.1630 0.1710 22.2110 ;
        RECT 3.7170 22.1630 3.7350 22.2110 ;
        RECT 4.9590 22.1630 4.9860 22.2110 ;
        RECT 5.1120 22.1630 5.1480 22.2110 ;
        RECT 5.8770 22.1630 5.8950 22.2110 ;
        RECT 9.4410 22.1630 9.4590 22.2110 ;
        RECT 0.1530 23.2430 0.1710 23.2910 ;
        RECT 3.7170 23.2430 3.7350 23.2910 ;
        RECT 4.9590 23.2430 4.9860 23.2910 ;
        RECT 5.1120 23.2430 5.1480 23.2910 ;
        RECT 5.8770 23.2430 5.8950 23.2910 ;
        RECT 9.4410 23.2430 9.4590 23.2910 ;
        RECT 0.1530 24.3230 0.1710 24.3710 ;
        RECT 3.7170 24.3230 3.7350 24.3710 ;
        RECT 4.9590 24.3230 4.9860 24.3710 ;
        RECT 5.1120 24.3230 5.1480 24.3710 ;
        RECT 5.8770 24.3230 5.8950 24.3710 ;
        RECT 9.4410 24.3230 9.4590 24.3710 ;
        RECT 0.1530 25.4030 0.1710 25.4510 ;
        RECT 3.7170 25.4030 3.7350 25.4510 ;
        RECT 4.9590 25.4030 4.9860 25.4510 ;
        RECT 5.1120 25.4030 5.1480 25.4510 ;
        RECT 5.8770 25.4030 5.8950 25.4510 ;
        RECT 9.4410 25.4030 9.4590 25.4510 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.3350 10.1230 7.3530 10.1600 ;
      LAYER M4  ;
        RECT 7.2830 10.1310 7.3670 10.1550 ;
      LAYER M5  ;
        RECT 7.3320 9.1800 7.3560 12.4200 ;
      LAYER V3  ;
        RECT 7.3350 10.1310 7.3530 10.1550 ;
      LAYER V4  ;
        RECT 7.3320 10.1310 7.3560 10.1550 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.1190 10.1260 7.1370 10.1630 ;
      LAYER M4  ;
        RECT 7.0670 10.1310 7.1510 10.1550 ;
      LAYER M5  ;
        RECT 7.1160 9.1800 7.1400 12.4200 ;
      LAYER V3  ;
        RECT 7.1190 10.1310 7.1370 10.1550 ;
      LAYER V4  ;
        RECT 7.1160 10.1310 7.1400 10.1550 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.9030 9.5470 6.9210 9.5840 ;
      LAYER M4  ;
        RECT 6.8510 9.5550 6.9350 9.5790 ;
      LAYER M5  ;
        RECT 6.9000 9.1800 6.9240 12.4200 ;
      LAYER V3  ;
        RECT 6.9030 9.5550 6.9210 9.5790 ;
      LAYER V4  ;
        RECT 6.9000 9.5550 6.9240 9.5790 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.6870 9.7870 6.7050 9.9680 ;
      LAYER M4  ;
        RECT 6.6350 9.9390 6.7190 9.9630 ;
      LAYER M5  ;
        RECT 6.6840 9.1800 6.7080 12.4200 ;
      LAYER V3  ;
        RECT 6.6870 9.9390 6.7050 9.9630 ;
      LAYER V4  ;
        RECT 6.6840 9.9390 6.7080 9.9630 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.4710 9.5500 6.4890 9.6170 ;
      LAYER M4  ;
        RECT 6.4190 9.5550 6.5030 9.5790 ;
      LAYER M5  ;
        RECT 6.4680 9.1800 6.4920 12.4200 ;
      LAYER V3  ;
        RECT 6.4710 9.5550 6.4890 9.5790 ;
      LAYER V4  ;
        RECT 6.4680 9.5550 6.4920 9.5790 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.2550 9.2830 6.2730 9.5360 ;
      LAYER M4  ;
        RECT 6.2030 9.5070 6.2870 9.5310 ;
      LAYER M5  ;
        RECT 6.2520 9.1800 6.2760 12.4200 ;
      LAYER V3  ;
        RECT 6.2550 9.5070 6.2730 9.5310 ;
      LAYER V4  ;
        RECT 6.2520 9.5070 6.2760 9.5310 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.0390 10.3180 6.0570 10.3550 ;
      LAYER M4  ;
        RECT 5.9870 10.3230 6.0710 10.3470 ;
      LAYER M5  ;
        RECT 6.0360 9.1800 6.0600 12.4200 ;
      LAYER V3  ;
        RECT 6.0390 10.3230 6.0570 10.3470 ;
      LAYER V4  ;
        RECT 6.0360 10.3230 6.0600 10.3470 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 5.1750 9.5500 5.1930 9.6170 ;
      LAYER M4  ;
        RECT 4.8910 9.5550 5.2040 9.5790 ;
      LAYER M5  ;
        RECT 4.9020 9.1800 4.9260 12.4200 ;
      LAYER V3  ;
        RECT 5.1750 9.5550 5.1930 9.5790 ;
      LAYER V4  ;
        RECT 4.9020 9.5550 4.9260 9.5790 ;
    END
  END ADDRESS[7]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 4.7790 9.2830 4.7970 9.5360 ;
      LAYER M4  ;
        RECT 4.5670 9.5070 4.8080 9.5310 ;
      LAYER M5  ;
        RECT 4.5780 9.1800 4.6020 12.4200 ;
      LAYER V3  ;
        RECT 4.7790 9.5070 4.7970 9.5310 ;
      LAYER V4  ;
        RECT 4.5780 9.5070 4.6020 9.5310 ;
    END
  END banksel
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.9870 9.5500 4.0050 9.6170 ;
      LAYER M4  ;
        RECT 3.9350 9.5550 4.0190 9.5790 ;
      LAYER M5  ;
        RECT 3.9840 9.1800 4.0080 12.4200 ;
      LAYER V3  ;
        RECT 3.9870 9.5550 4.0050 9.5790 ;
      LAYER V4  ;
        RECT 3.9840 9.5550 4.0080 9.5790 ;
    END
  END write
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.7710 10.4140 3.7890 10.4630 ;
      LAYER M4  ;
        RECT 3.7190 10.4190 3.8030 10.4430 ;
      LAYER M5  ;
        RECT 3.7680 9.1800 3.7920 12.4200 ;
      LAYER V3  ;
        RECT 3.7710 10.4190 3.7890 10.4430 ;
      LAYER V4  ;
        RECT 3.7680 10.4190 3.7920 10.4430 ;
    END
  END clk
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.8070 9.2830 3.8250 9.5360 ;
      LAYER M4  ;
        RECT 3.5410 9.5070 3.8360 9.5310 ;
      LAYER M5  ;
        RECT 3.5520 9.1800 3.5760 12.4200 ;
      LAYER V3  ;
        RECT 3.8070 9.5070 3.8250 9.5310 ;
      LAYER V4  ;
        RECT 3.5520 9.5070 3.5760 9.5310 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.3390 10.1230 3.3570 10.1600 ;
      LAYER M4  ;
        RECT 3.2870 10.1310 3.3710 10.1550 ;
      LAYER M5  ;
        RECT 3.3360 9.1800 3.3600 12.4200 ;
      LAYER V3  ;
        RECT 3.3390 10.1310 3.3570 10.1550 ;
      LAYER V4  ;
        RECT 3.3360 10.1310 3.3600 10.1550 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 3.1230 9.5500 3.1410 9.7790 ;
      LAYER M4  ;
        RECT 3.0710 9.5550 3.1550 9.5790 ;
      LAYER M5  ;
        RECT 3.1200 9.1800 3.1440 12.4200 ;
      LAYER V3  ;
        RECT 3.1230 9.5550 3.1410 9.5790 ;
      LAYER V4  ;
        RECT 3.1200 9.5550 3.1440 9.5790 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.9070 9.2830 2.9250 9.5360 ;
      LAYER M4  ;
        RECT 2.8550 9.5070 2.9390 9.5310 ;
      LAYER M5  ;
        RECT 2.9040 9.1800 2.9280 12.4200 ;
      LAYER V3  ;
        RECT 2.9070 9.5070 2.9250 9.5310 ;
      LAYER V4  ;
        RECT 2.9040 9.5070 2.9280 9.5310 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.6910 9.5470 2.7090 9.5840 ;
      LAYER M4  ;
        RECT 2.6390 9.5550 2.7230 9.5790 ;
      LAYER M5  ;
        RECT 2.6880 9.1800 2.7120 12.4200 ;
      LAYER V3  ;
        RECT 2.6910 9.5550 2.7090 9.5790 ;
      LAYER V4  ;
        RECT 2.6880 9.5550 2.7120 9.5790 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 2.4750 10.1230 2.4930 10.1600 ;
      LAYER M4  ;
        RECT 2.4230 10.1310 2.5070 10.1550 ;
      LAYER M5  ;
        RECT 2.4720 9.1800 2.4960 12.4200 ;
      LAYER V3  ;
        RECT 2.4750 10.1310 2.4930 10.1550 ;
      LAYER V4  ;
        RECT 2.4720 10.1310 2.4960 10.1550 ;
    END
  END sdel[4]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 0.4280 5.1360 0.4520 ;
      LAYER M3  ;
        RECT 5.0760 0.3775 5.0940 0.6170 ;
      LAYER V3  ;
        RECT 5.0760 0.4280 5.0940 0.4520 ;
    END
  END dataout[0]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 0.3320 5.2040 0.3560 ;
      LAYER M3  ;
        RECT 4.8510 0.2700 4.8690 0.6750 ;
      LAYER V3  ;
        RECT 4.8510 0.3320 4.8690 0.3560 ;
    END
  END wd[0]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 1.5080 5.1360 1.5320 ;
      LAYER M3  ;
        RECT 5.0760 1.4575 5.0940 1.6970 ;
      LAYER V3  ;
        RECT 5.0760 1.5080 5.0940 1.5320 ;
    END
  END dataout[1]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 1.4120 5.2040 1.4360 ;
      LAYER M3  ;
        RECT 4.8510 1.3500 4.8690 1.7550 ;
      LAYER V3  ;
        RECT 4.8510 1.4120 4.8690 1.4360 ;
    END
  END wd[1]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 2.5880 5.1360 2.6120 ;
      LAYER M3  ;
        RECT 5.0760 2.5375 5.0940 2.7770 ;
      LAYER V3  ;
        RECT 5.0760 2.5880 5.0940 2.6120 ;
    END
  END dataout[2]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 2.4920 5.2040 2.5160 ;
      LAYER M3  ;
        RECT 4.8510 2.4300 4.8690 2.8350 ;
      LAYER V3  ;
        RECT 4.8510 2.4920 4.8690 2.5160 ;
    END
  END wd[2]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 3.6680 5.1360 3.6920 ;
      LAYER M3  ;
        RECT 5.0760 3.6175 5.0940 3.8570 ;
      LAYER V3  ;
        RECT 5.0760 3.6680 5.0940 3.6920 ;
    END
  END dataout[3]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 3.5720 5.2040 3.5960 ;
      LAYER M3  ;
        RECT 4.8510 3.5100 4.8690 3.9150 ;
      LAYER V3  ;
        RECT 4.8510 3.5720 4.8690 3.5960 ;
    END
  END wd[3]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 4.7480 5.1360 4.7720 ;
      LAYER M3  ;
        RECT 5.0760 4.6975 5.0940 4.9370 ;
      LAYER V3  ;
        RECT 5.0760 4.7480 5.0940 4.7720 ;
    END
  END dataout[4]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 4.6520 5.2040 4.6760 ;
      LAYER M3  ;
        RECT 4.8510 4.5900 4.8690 4.9950 ;
      LAYER V3  ;
        RECT 4.8510 4.6520 4.8690 4.6760 ;
    END
  END wd[4]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 5.8280 5.1360 5.8520 ;
      LAYER M3  ;
        RECT 5.0760 5.7775 5.0940 6.0170 ;
      LAYER V3  ;
        RECT 5.0760 5.8280 5.0940 5.8520 ;
    END
  END dataout[5]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 5.7320 5.2040 5.7560 ;
      LAYER M3  ;
        RECT 4.8510 5.6700 4.8690 6.0750 ;
      LAYER V3  ;
        RECT 4.8510 5.7320 4.8690 5.7560 ;
    END
  END wd[5]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 6.9080 5.1360 6.9320 ;
      LAYER M3  ;
        RECT 5.0760 6.8575 5.0940 7.0970 ;
      LAYER V3  ;
        RECT 5.0760 6.9080 5.0940 6.9320 ;
    END
  END dataout[6]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 6.8120 5.2040 6.8360 ;
      LAYER M3  ;
        RECT 4.8510 6.7500 4.8690 7.1550 ;
      LAYER V3  ;
        RECT 4.8510 6.8120 4.8690 6.8360 ;
    END
  END wd[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 7.9880 5.1360 8.0120 ;
      LAYER M3  ;
        RECT 5.0760 7.9375 5.0940 8.1770 ;
      LAYER V3  ;
        RECT 5.0760 7.9880 5.0940 8.0120 ;
    END
  END dataout[7]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 7.8920 5.2040 7.9160 ;
      LAYER M3  ;
        RECT 4.8510 7.8300 4.8690 8.2350 ;
      LAYER V3  ;
        RECT 4.8510 7.8920 4.8690 7.9160 ;
    END
  END wd[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 17.1950 5.1360 17.2190 ;
      LAYER M3  ;
        RECT 5.0760 17.1445 5.0940 17.3840 ;
      LAYER V3  ;
        RECT 5.0760 17.1950 5.0940 17.2190 ;
    END
  END dataout[8]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 17.0990 5.2040 17.1230 ;
      LAYER M3  ;
        RECT 4.8510 17.0370 4.8690 17.4420 ;
      LAYER V3  ;
        RECT 4.8510 17.0990 4.8690 17.1230 ;
    END
  END wd[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 18.2750 5.1360 18.2990 ;
      LAYER M3  ;
        RECT 5.0760 18.2245 5.0940 18.4640 ;
      LAYER V3  ;
        RECT 5.0760 18.2750 5.0940 18.2990 ;
    END
  END dataout[9]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 18.1790 5.2040 18.2030 ;
      LAYER M3  ;
        RECT 4.8510 18.1170 4.8690 18.5220 ;
      LAYER V3  ;
        RECT 4.8510 18.1790 4.8690 18.2030 ;
    END
  END wd[9]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 19.3550 5.1360 19.3790 ;
      LAYER M3  ;
        RECT 5.0760 19.3045 5.0940 19.5440 ;
      LAYER V3  ;
        RECT 5.0760 19.3550 5.0940 19.3790 ;
    END
  END dataout[10]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 19.2590 5.2040 19.2830 ;
      LAYER M3  ;
        RECT 4.8510 19.1970 4.8690 19.6020 ;
      LAYER V3  ;
        RECT 4.8510 19.2590 4.8690 19.2830 ;
    END
  END wd[10]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 20.4350 5.1360 20.4590 ;
      LAYER M3  ;
        RECT 5.0760 20.3845 5.0940 20.6240 ;
      LAYER V3  ;
        RECT 5.0760 20.4350 5.0940 20.4590 ;
    END
  END dataout[11]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 20.3390 5.2040 20.3630 ;
      LAYER M3  ;
        RECT 4.8510 20.2770 4.8690 20.6820 ;
      LAYER V3  ;
        RECT 4.8510 20.3390 4.8690 20.3630 ;
    END
  END wd[11]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 21.5150 5.1360 21.5390 ;
      LAYER M3  ;
        RECT 5.0760 21.4645 5.0940 21.7040 ;
      LAYER V3  ;
        RECT 5.0760 21.5150 5.0940 21.5390 ;
    END
  END dataout[12]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 21.4190 5.2040 21.4430 ;
      LAYER M3  ;
        RECT 4.8510 21.3570 4.8690 21.7620 ;
      LAYER V3  ;
        RECT 4.8510 21.4190 4.8690 21.4430 ;
    END
  END wd[12]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 22.5950 5.1360 22.6190 ;
      LAYER M3  ;
        RECT 5.0760 22.5445 5.0940 22.7840 ;
      LAYER V3  ;
        RECT 5.0760 22.5950 5.0940 22.6190 ;
    END
  END dataout[13]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 22.4990 5.2040 22.5230 ;
      LAYER M3  ;
        RECT 4.8510 22.4370 4.8690 22.8420 ;
      LAYER V3  ;
        RECT 4.8510 22.4990 4.8690 22.5230 ;
    END
  END wd[13]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 23.6750 5.1360 23.6990 ;
      LAYER M3  ;
        RECT 5.0760 23.6245 5.0940 23.8640 ;
      LAYER V3  ;
        RECT 5.0760 23.6750 5.0940 23.6990 ;
    END
  END dataout[14]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 23.5790 5.2040 23.6030 ;
      LAYER M3  ;
        RECT 4.8510 23.5170 4.8690 23.9220 ;
      LAYER V3  ;
        RECT 4.8510 23.5790 4.8690 23.6030 ;
    END
  END wd[14]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 24.7550 5.1360 24.7790 ;
      LAYER M3  ;
        RECT 5.0760 24.7045 5.0940 24.9440 ;
      LAYER V3  ;
        RECT 5.0760 24.7550 5.0940 24.7790 ;
    END
  END dataout[15]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 4.4880 24.6590 5.2040 24.6830 ;
      LAYER M3  ;
        RECT 4.8510 24.5970 4.8690 25.0020 ;
      LAYER V3  ;
        RECT 4.8510 24.6590 4.8690 24.6830 ;
    END
  END wd[15]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8830 9.6120 17.5365 ;
        RECT 0.0000 17.0235 9.6120 18.1170 ;
        RECT 0.0000 18.1035 9.6120 19.1970 ;
        RECT 0.0000 19.1835 9.6120 20.2770 ;
        RECT 0.0000 20.2635 9.6120 21.3570 ;
        RECT 0.0000 21.3435 9.6120 22.4370 ;
        RECT 0.0000 22.4235 9.6120 23.5170 ;
        RECT 0.0000 23.5035 9.6120 24.5970 ;
        RECT 0.0000 24.5835 9.6120 25.6770 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8830 9.6120 17.5365 ;
        RECT 0.0000 17.0235 9.6120 18.1170 ;
        RECT 0.0000 18.1035 9.6120 19.1970 ;
        RECT 0.0000 19.1835 9.6120 20.2770 ;
        RECT 0.0000 20.2635 9.6120 21.3570 ;
        RECT 0.0000 21.3435 9.6120 22.4370 ;
        RECT 0.0000 22.4235 9.6120 23.5170 ;
        RECT 0.0000 23.5035 9.6120 24.5970 ;
        RECT 0.0000 24.5835 9.6120 25.6770 ;
  LAYER V1  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8830 9.6120 17.5365 ;
        RECT 0.0000 17.0235 9.6120 18.1170 ;
        RECT 0.0000 18.1035 9.6120 19.1970 ;
        RECT 0.0000 19.1835 9.6120 20.2770 ;
        RECT 0.0000 20.2635 9.6120 21.3570 ;
        RECT 0.0000 21.3435 9.6120 22.4370 ;
        RECT 0.0000 22.4235 9.6120 23.5170 ;
        RECT 0.0000 23.5035 9.6120 24.5970 ;
        RECT 0.0000 24.5835 9.6120 25.6770 ;
  LAYER V2  ;
      RECT 0.0000 0.2565 9.6120 1.3500 ;
      RECT 0.0000 1.3365 9.6120 2.4300 ;
      RECT 0.0000 2.4165 9.6120 3.5100 ;
      RECT 0.0000 3.4965 9.6120 4.5900 ;
      RECT 0.0000 4.5765 9.6120 5.6700 ;
      RECT 0.0000 5.6565 9.6120 6.7500 ;
      RECT 0.0000 6.7365 9.6120 7.8300 ;
      RECT 0.0000 7.8165 9.6120 8.9100 ;
      RECT 0.0000 8.8830 9.6120 17.5365 ;
        RECT 0.0000 17.0235 9.6120 18.1170 ;
        RECT 0.0000 18.1035 9.6120 19.1970 ;
        RECT 0.0000 19.1835 9.6120 20.2770 ;
        RECT 0.0000 20.2635 9.6120 21.3570 ;
        RECT 0.0000 21.3435 9.6120 22.4370 ;
        RECT 0.0000 22.4235 9.6120 23.5170 ;
        RECT 0.0000 23.5035 9.6120 24.5970 ;
        RECT 0.0000 24.5835 9.6120 25.6770 ;
  LAYER M3  ;
      RECT 5.2380 0.3450 5.2560 1.2805 ;
      RECT 5.2020 0.3450 5.2200 1.2805 ;
      RECT 5.1660 0.9220 5.1840 1.2445 ;
      RECT 5.0490 1.1190 5.0670 1.2285 ;
      RECT 5.0400 0.3775 5.0580 0.6170 ;
      RECT 5.0040 0.9585 5.0220 1.1120 ;
      RECT 4.9230 0.9840 4.9410 1.2420 ;
      RECT 4.3830 0.3450 4.4010 1.2805 ;
      RECT 4.3470 0.3450 4.3650 1.2805 ;
      RECT 4.3110 0.5260 4.3290 1.0940 ;
      RECT 5.2380 1.4250 5.2560 2.3605 ;
      RECT 5.2020 1.4250 5.2200 2.3605 ;
      RECT 5.1660 2.0020 5.1840 2.3245 ;
      RECT 5.0490 2.1990 5.0670 2.3085 ;
      RECT 5.0400 1.4575 5.0580 1.6970 ;
      RECT 5.0040 2.0385 5.0220 2.1920 ;
      RECT 4.9230 2.0640 4.9410 2.3220 ;
      RECT 4.3830 1.4250 4.4010 2.3605 ;
      RECT 4.3470 1.4250 4.3650 2.3605 ;
      RECT 4.3110 1.6060 4.3290 2.1740 ;
      RECT 5.2380 2.5050 5.2560 3.4405 ;
      RECT 5.2020 2.5050 5.2200 3.4405 ;
      RECT 5.1660 3.0820 5.1840 3.4045 ;
      RECT 5.0490 3.2790 5.0670 3.3885 ;
      RECT 5.0400 2.5375 5.0580 2.7770 ;
      RECT 5.0040 3.1185 5.0220 3.2720 ;
      RECT 4.9230 3.1440 4.9410 3.4020 ;
      RECT 4.3830 2.5050 4.4010 3.4405 ;
      RECT 4.3470 2.5050 4.3650 3.4405 ;
      RECT 4.3110 2.6860 4.3290 3.2540 ;
      RECT 5.2380 3.5850 5.2560 4.5205 ;
      RECT 5.2020 3.5850 5.2200 4.5205 ;
      RECT 5.1660 4.1620 5.1840 4.4845 ;
      RECT 5.0490 4.3590 5.0670 4.4685 ;
      RECT 5.0400 3.6175 5.0580 3.8570 ;
      RECT 5.0040 4.1985 5.0220 4.3520 ;
      RECT 4.9230 4.2240 4.9410 4.4820 ;
      RECT 4.3830 3.5850 4.4010 4.5205 ;
      RECT 4.3470 3.5850 4.3650 4.5205 ;
      RECT 4.3110 3.7660 4.3290 4.3340 ;
      RECT 5.2380 4.6650 5.2560 5.6005 ;
      RECT 5.2020 4.6650 5.2200 5.6005 ;
      RECT 5.1660 5.2420 5.1840 5.5645 ;
      RECT 5.0490 5.4390 5.0670 5.5485 ;
      RECT 5.0400 4.6975 5.0580 4.9370 ;
      RECT 5.0040 5.2785 5.0220 5.4320 ;
      RECT 4.9230 5.3040 4.9410 5.5620 ;
      RECT 4.3830 4.6650 4.4010 5.6005 ;
      RECT 4.3470 4.6650 4.3650 5.6005 ;
      RECT 4.3110 4.8460 4.3290 5.4140 ;
      RECT 5.2380 5.7450 5.2560 6.6805 ;
      RECT 5.2020 5.7450 5.2200 6.6805 ;
      RECT 5.1660 6.3220 5.1840 6.6445 ;
      RECT 5.0490 6.5190 5.0670 6.6285 ;
      RECT 5.0400 5.7775 5.0580 6.0170 ;
      RECT 5.0040 6.3585 5.0220 6.5120 ;
      RECT 4.9230 6.3840 4.9410 6.6420 ;
      RECT 4.3830 5.7450 4.4010 6.6805 ;
      RECT 4.3470 5.7450 4.3650 6.6805 ;
      RECT 4.3110 5.9260 4.3290 6.4940 ;
      RECT 5.2380 6.8250 5.2560 7.7605 ;
      RECT 5.2020 6.8250 5.2200 7.7605 ;
      RECT 5.1660 7.4020 5.1840 7.7245 ;
      RECT 5.0490 7.5990 5.0670 7.7085 ;
      RECT 5.0400 6.8575 5.0580 7.0970 ;
      RECT 5.0040 7.4385 5.0220 7.5920 ;
      RECT 4.9230 7.4640 4.9410 7.7220 ;
      RECT 4.3830 6.8250 4.4010 7.7605 ;
      RECT 4.3470 6.8250 4.3650 7.7605 ;
      RECT 4.3110 7.0060 4.3290 7.5740 ;
      RECT 5.2380 7.9050 5.2560 8.8405 ;
      RECT 5.2020 7.9050 5.2200 8.8405 ;
      RECT 5.1660 8.4820 5.1840 8.8045 ;
      RECT 5.0490 8.6790 5.0670 8.7885 ;
      RECT 5.0400 7.9375 5.0580 8.1770 ;
      RECT 5.0040 8.5185 5.0220 8.6720 ;
      RECT 4.9230 8.5440 4.9410 8.8020 ;
      RECT 4.3830 7.9050 4.4010 8.8405 ;
      RECT 4.3470 7.9050 4.3650 8.8405 ;
      RECT 4.3110 8.0860 4.3290 8.6540 ;
      RECT 9.4050 12.6760 9.4230 17.0315 ;
      RECT 9.3690 11.3610 9.3870 11.4300 ;
      RECT 9.3690 13.1690 9.3870 13.6335 ;
      RECT 9.3330 8.8565 9.3510 17.0635 ;
      RECT 9.2970 12.6260 9.3150 13.3985 ;
      RECT 9.2970 13.4497 9.3150 13.9410 ;
      RECT 9.2970 13.9910 9.3150 14.3625 ;
      RECT 9.2970 14.4255 9.3150 15.2370 ;
      RECT 9.2610 12.7115 9.2790 13.3535 ;
      RECT 9.2610 14.0310 9.2790 14.5630 ;
      RECT 9.2250 8.8565 9.2430 9.2065 ;
      RECT 9.1170 8.8565 9.1350 9.2065 ;
      RECT 9.0090 8.8565 9.0270 9.2065 ;
      RECT 8.9010 8.8565 8.9190 9.2065 ;
      RECT 8.7930 8.8565 8.8110 9.2065 ;
      RECT 8.6850 8.8565 8.7030 9.2065 ;
      RECT 8.5770 8.8565 8.5950 9.2065 ;
      RECT 8.4690 8.8565 8.4870 9.2065 ;
      RECT 8.3610 8.8565 8.3790 9.2065 ;
      RECT 8.2530 8.8565 8.2710 9.2065 ;
      RECT 8.1450 8.8565 8.1630 9.2065 ;
      RECT 8.0370 8.8565 8.0550 9.2065 ;
      RECT 7.9290 8.8565 7.9470 9.2065 ;
      RECT 7.8210 8.8565 7.8390 9.2065 ;
      RECT 7.7130 8.8565 7.7310 9.2065 ;
      RECT 7.6050 8.8565 7.6230 9.2065 ;
      RECT 7.4970 8.8565 7.5150 9.2065 ;
      RECT 7.3890 8.8565 7.4070 9.2065 ;
      RECT 7.2810 8.8565 7.2990 9.2065 ;
      RECT 7.1730 8.8565 7.1910 9.2065 ;
      RECT 7.0650 8.8565 7.0830 9.2065 ;
      RECT 6.9570 8.8565 6.9750 9.2065 ;
      RECT 6.8490 8.8565 6.8670 9.2065 ;
      RECT 6.7410 8.8565 6.7590 9.2065 ;
      RECT 6.6330 8.8565 6.6510 9.2065 ;
      RECT 6.5250 8.8565 6.5430 9.2065 ;
      RECT 6.4170 8.8565 6.4350 9.2065 ;
      RECT 6.3090 8.8565 6.3270 9.2065 ;
      RECT 6.2010 8.8565 6.2190 9.2065 ;
      RECT 6.0930 8.8565 6.1110 9.2065 ;
      RECT 6.0570 12.6450 6.0750 13.3498 ;
      RECT 6.0570 14.0920 6.0750 15.2730 ;
      RECT 6.0390 9.5170 6.0570 10.1930 ;
      RECT 6.0390 10.9390 6.0570 11.2370 ;
      RECT 6.0210 12.7085 6.0390 13.3985 ;
      RECT 6.0210 13.4495 6.0390 14.4410 ;
      RECT 6.0210 14.4710 6.0390 15.2550 ;
      RECT 5.9850 8.8565 6.0030 17.0635 ;
      RECT 5.9490 12.9810 5.9670 13.0640 ;
      RECT 5.9310 9.6250 5.9490 10.2560 ;
      RECT 5.9310 10.6690 5.9490 10.8590 ;
      RECT 5.9310 11.5510 5.9490 11.6000 ;
      RECT 5.9130 12.6760 5.9310 17.0360 ;
      RECT 5.8230 9.2470 5.8410 10.0490 ;
      RECT 5.8230 10.5970 5.8410 11.1650 ;
      RECT 5.7870 10.6690 5.8050 11.0390 ;
      RECT 5.7510 10.0210 5.7690 10.1570 ;
      RECT 5.7510 11.0110 5.7690 11.2370 ;
      RECT 5.7510 12.2530 5.7690 12.3170 ;
      RECT 5.7150 10.1230 5.7330 10.1600 ;
      RECT 5.7150 11.7490 5.7330 11.7920 ;
      RECT 5.7150 12.2830 5.7330 12.3200 ;
      RECT 5.6790 10.4350 5.6970 10.9310 ;
      RECT 5.6790 10.9750 5.6970 11.1650 ;
      RECT 5.6790 11.9350 5.6970 12.2450 ;
      RECT 5.6430 14.2150 5.6610 14.9450 ;
      RECT 5.6430 15.2950 5.6610 16.0250 ;
      RECT 5.3190 10.0570 5.3370 10.3550 ;
      RECT 5.3190 11.2450 5.3370 11.3090 ;
      RECT 5.3190 11.5150 5.3370 11.9750 ;
      RECT 5.3190 12.7150 5.3370 12.7520 ;
      RECT 5.3190 14.7550 5.3370 15.0530 ;
      RECT 5.2830 10.1290 5.3010 10.6340 ;
      RECT 5.2830 10.9030 5.3010 11.7050 ;
      RECT 5.2830 12.7480 5.3010 13.0190 ;
      RECT 5.2830 13.0990 5.3010 13.3250 ;
      RECT 5.2470 10.0570 5.2650 10.7330 ;
      RECT 5.2470 10.8310 5.2650 11.1650 ;
      RECT 5.2470 11.3710 5.2650 11.5070 ;
      RECT 5.2470 12.0550 5.2650 12.8570 ;
      RECT 5.2470 13.2910 5.2650 13.3280 ;
      RECT 5.2470 15.4570 5.2650 15.7910 ;
      RECT 5.2110 10.2910 5.2290 10.4270 ;
      RECT 5.2110 12.1810 5.2290 13.1630 ;
      RECT 5.2110 13.6030 5.2290 13.9010 ;
      RECT 5.2110 15.2950 5.2290 15.5570 ;
      RECT 5.1750 9.3550 5.1930 9.5090 ;
      RECT 5.1750 10.1650 5.1930 11.9510 ;
      RECT 5.1750 12.9910 5.1930 15.3230 ;
      RECT 5.1750 15.5290 5.1930 16.6370 ;
      RECT 4.8870 9.6250 4.9050 9.8870 ;
      RECT 4.8870 10.0210 4.9050 10.0850 ;
      RECT 4.8870 10.1650 4.9050 10.3910 ;
      RECT 4.8870 10.4350 4.9050 10.6250 ;
      RECT 4.8870 10.7050 4.9050 13.3250 ;
      RECT 4.8870 13.3690 4.9050 14.6750 ;
      RECT 4.8870 15.7630 4.9050 16.0250 ;
      RECT 4.8510 10.6240 4.8690 10.8950 ;
      RECT 4.8510 10.9750 4.8690 11.8130 ;
      RECT 4.8510 11.9830 4.8690 12.8210 ;
      RECT 4.8510 12.8650 4.8690 14.1350 ;
      RECT 4.8510 14.3410 4.8690 14.5130 ;
      RECT 4.8510 15.2230 4.8690 16.2950 ;
      RECT 4.8150 10.7050 4.8330 10.9760 ;
      RECT 4.8150 11.1310 4.8330 11.1680 ;
      RECT 4.8150 11.9110 4.8330 12.8930 ;
      RECT 4.8150 13.1350 4.8330 13.5950 ;
      RECT 4.8150 13.9450 4.8330 14.6840 ;
      RECT 4.7790 9.8230 4.7970 10.8950 ;
      RECT 4.7790 12.4870 4.7970 12.7040 ;
      RECT 4.7790 13.8730 4.7970 14.1710 ;
      RECT 4.7430 10.4710 4.7610 10.9310 ;
      RECT 4.7430 12.0550 4.7610 12.2450 ;
      RECT 4.7430 12.2860 4.7610 12.3230 ;
      RECT 4.7430 12.5590 4.7610 12.8930 ;
      RECT 4.7430 13.0270 4.7610 14.3690 ;
      RECT 4.7430 14.4760 4.7610 15.5930 ;
      RECT 4.7070 9.8950 4.7250 10.0850 ;
      RECT 4.7070 10.2910 4.7250 10.4270 ;
      RECT 4.7070 10.7050 4.7250 13.8650 ;
      RECT 4.7070 13.9450 4.7250 14.4050 ;
      RECT 4.7070 15.0250 4.7250 15.4850 ;
      RECT 4.7070 16.3390 4.7250 16.5650 ;
      RECT 4.6710 8.8830 4.6890 9.0370 ;
      RECT 4.6710 16.8940 4.6890 17.0480 ;
      RECT 4.6350 8.8830 4.6530 8.9330 ;
      RECT 4.5630 8.8830 4.5810 8.9545 ;
      RECT 4.5630 16.9635 4.5810 17.0635 ;
      RECT 4.4190 10.3990 4.4370 10.5890 ;
      RECT 4.4190 11.1370 4.4370 11.5070 ;
      RECT 4.4190 13.0990 4.4370 13.3250 ;
      RECT 4.4190 13.6390 4.4370 14.7830 ;
      RECT 4.4190 15.5650 4.4370 16.0250 ;
      RECT 4.4190 16.6030 4.4370 16.6400 ;
      RECT 4.3830 9.3550 4.4010 9.8510 ;
      RECT 4.3830 13.4350 4.4010 13.4720 ;
      RECT 4.3830 14.5120 4.4010 15.3230 ;
      RECT 4.3470 9.8230 4.3650 10.0850 ;
      RECT 4.3470 10.3630 4.3650 10.6970 ;
      RECT 4.3470 10.9030 4.3650 11.0030 ;
      RECT 4.3470 11.7850 4.3650 14.5490 ;
      RECT 4.3470 14.6830 4.3650 14.9090 ;
      RECT 4.3110 9.4810 4.3290 10.6250 ;
      RECT 4.3110 14.2150 4.3290 14.4050 ;
      RECT 4.3110 15.0190 4.3290 15.0560 ;
      RECT 4.3110 15.2950 4.3290 16.0970 ;
      RECT 4.2750 10.4350 4.2930 11.4350 ;
      RECT 4.2750 14.8750 4.2930 14.9120 ;
      RECT 4.2390 9.6250 4.2570 9.6530 ;
      RECT 3.9150 10.0210 3.9330 10.4270 ;
      RECT 3.8430 10.0570 3.8610 10.6610 ;
      RECT 3.8070 9.8950 3.8250 9.9590 ;
      RECT 3.7710 8.9360 3.7890 8.9870 ;
      RECT 3.7710 12.0550 3.7890 12.2450 ;
      RECT 3.7710 12.6760 3.7890 17.0360 ;
      RECT 3.6810 12.6760 3.6990 17.0360 ;
      RECT 3.6630 9.3550 3.6810 9.5450 ;
      RECT 3.6630 10.1290 3.6810 12.3890 ;
      RECT 3.6450 12.9810 3.6630 13.0640 ;
      RECT 3.6090 8.8565 3.6270 17.0635 ;
      RECT 3.5730 12.7085 3.5910 13.3985 ;
      RECT 3.5730 13.4495 3.5910 14.4410 ;
      RECT 3.5730 14.4710 3.5910 15.2550 ;
      RECT 3.5550 9.3550 3.5730 9.8510 ;
      RECT 3.5550 10.6330 3.5730 11.2010 ;
      RECT 3.5550 11.5150 3.5730 12.2450 ;
      RECT 3.5370 12.6450 3.5550 13.3498 ;
      RECT 3.5370 14.0920 3.5550 15.2730 ;
      RECT 3.5010 8.8565 3.5190 9.2065 ;
      RECT 3.3930 8.8565 3.4110 9.2065 ;
      RECT 3.2850 8.8565 3.3030 9.2065 ;
      RECT 3.1770 8.8565 3.1950 9.2065 ;
      RECT 3.0690 8.8565 3.0870 9.2065 ;
      RECT 2.9610 8.8565 2.9790 9.2065 ;
      RECT 2.8530 8.8565 2.8710 9.2065 ;
      RECT 2.7450 8.8565 2.7630 9.2065 ;
      RECT 2.6370 8.8565 2.6550 9.2065 ;
      RECT 2.5290 8.8565 2.5470 9.2065 ;
      RECT 2.4210 8.8565 2.4390 9.2065 ;
      RECT 2.3130 8.8565 2.3310 9.2065 ;
      RECT 2.2050 8.8565 2.2230 9.2065 ;
      RECT 2.0970 8.8565 2.1150 9.2065 ;
      RECT 1.9890 8.8565 2.0070 9.2065 ;
      RECT 1.8810 8.8565 1.8990 9.2065 ;
      RECT 1.7730 8.8565 1.7910 9.2065 ;
      RECT 1.6650 8.8565 1.6830 9.2065 ;
      RECT 1.5570 8.8565 1.5750 9.2065 ;
      RECT 1.4490 8.8565 1.4670 9.2065 ;
      RECT 1.3410 8.8565 1.3590 9.2065 ;
      RECT 1.2330 8.8565 1.2510 9.2065 ;
      RECT 1.1250 8.8565 1.1430 9.2065 ;
      RECT 1.0170 8.8565 1.0350 9.2065 ;
      RECT 0.9090 8.8565 0.9270 9.2065 ;
      RECT 0.8010 8.8565 0.8190 9.2065 ;
      RECT 0.6930 8.8565 0.7110 9.2065 ;
      RECT 0.5850 8.8565 0.6030 9.2065 ;
      RECT 0.4770 8.8565 0.4950 9.2065 ;
      RECT 0.3690 8.8565 0.3870 9.2065 ;
      RECT 0.3330 12.7115 0.3510 13.3535 ;
      RECT 0.3330 14.0310 0.3510 14.5630 ;
      RECT 0.3150 9.8950 0.3330 10.1210 ;
      RECT 0.2970 12.6260 0.3150 13.3985 ;
      RECT 0.2970 13.4497 0.3150 13.9410 ;
      RECT 0.2970 13.9910 0.3150 14.3625 ;
      RECT 0.2970 14.4255 0.3150 15.2370 ;
      RECT 0.2610 8.8565 0.2790 17.0635 ;
      RECT 0.2250 11.3610 0.2430 11.4300 ;
      RECT 0.2250 13.1690 0.2430 13.6335 ;
      RECT 0.1890 12.6760 0.2070 17.0315 ;
        RECT 5.2380 17.1120 5.2560 18.0475 ;
        RECT 5.2020 17.1120 5.2200 18.0475 ;
        RECT 5.1660 17.6890 5.1840 18.0115 ;
        RECT 5.0490 17.8860 5.0670 17.9955 ;
        RECT 5.0400 17.1445 5.0580 17.3840 ;
        RECT 5.0040 17.7255 5.0220 17.8790 ;
        RECT 4.9230 17.7510 4.9410 18.0090 ;
        RECT 4.3830 17.1120 4.4010 18.0475 ;
        RECT 4.3470 17.1120 4.3650 18.0475 ;
        RECT 4.3110 17.2930 4.3290 17.8610 ;
        RECT 5.2380 18.1920 5.2560 19.1275 ;
        RECT 5.2020 18.1920 5.2200 19.1275 ;
        RECT 5.1660 18.7690 5.1840 19.0915 ;
        RECT 5.0490 18.9660 5.0670 19.0755 ;
        RECT 5.0400 18.2245 5.0580 18.4640 ;
        RECT 5.0040 18.8055 5.0220 18.9590 ;
        RECT 4.9230 18.8310 4.9410 19.0890 ;
        RECT 4.3830 18.1920 4.4010 19.1275 ;
        RECT 4.3470 18.1920 4.3650 19.1275 ;
        RECT 4.3110 18.3730 4.3290 18.9410 ;
        RECT 5.2380 19.2720 5.2560 20.2075 ;
        RECT 5.2020 19.2720 5.2200 20.2075 ;
        RECT 5.1660 19.8490 5.1840 20.1715 ;
        RECT 5.0490 20.0460 5.0670 20.1555 ;
        RECT 5.0400 19.3045 5.0580 19.5440 ;
        RECT 5.0040 19.8855 5.0220 20.0390 ;
        RECT 4.9230 19.9110 4.9410 20.1690 ;
        RECT 4.3830 19.2720 4.4010 20.2075 ;
        RECT 4.3470 19.2720 4.3650 20.2075 ;
        RECT 4.3110 19.4530 4.3290 20.0210 ;
        RECT 5.2380 20.3520 5.2560 21.2875 ;
        RECT 5.2020 20.3520 5.2200 21.2875 ;
        RECT 5.1660 20.9290 5.1840 21.2515 ;
        RECT 5.0490 21.1260 5.0670 21.2355 ;
        RECT 5.0400 20.3845 5.0580 20.6240 ;
        RECT 5.0040 20.9655 5.0220 21.1190 ;
        RECT 4.9230 20.9910 4.9410 21.2490 ;
        RECT 4.3830 20.3520 4.4010 21.2875 ;
        RECT 4.3470 20.3520 4.3650 21.2875 ;
        RECT 4.3110 20.5330 4.3290 21.1010 ;
        RECT 5.2380 21.4320 5.2560 22.3675 ;
        RECT 5.2020 21.4320 5.2200 22.3675 ;
        RECT 5.1660 22.0090 5.1840 22.3315 ;
        RECT 5.0490 22.2060 5.0670 22.3155 ;
        RECT 5.0400 21.4645 5.0580 21.7040 ;
        RECT 5.0040 22.0455 5.0220 22.1990 ;
        RECT 4.9230 22.0710 4.9410 22.3290 ;
        RECT 4.3830 21.4320 4.4010 22.3675 ;
        RECT 4.3470 21.4320 4.3650 22.3675 ;
        RECT 4.3110 21.6130 4.3290 22.1810 ;
        RECT 5.2380 22.5120 5.2560 23.4475 ;
        RECT 5.2020 22.5120 5.2200 23.4475 ;
        RECT 5.1660 23.0890 5.1840 23.4115 ;
        RECT 5.0490 23.2860 5.0670 23.3955 ;
        RECT 5.0400 22.5445 5.0580 22.7840 ;
        RECT 5.0040 23.1255 5.0220 23.2790 ;
        RECT 4.9230 23.1510 4.9410 23.4090 ;
        RECT 4.3830 22.5120 4.4010 23.4475 ;
        RECT 4.3470 22.5120 4.3650 23.4475 ;
        RECT 4.3110 22.6930 4.3290 23.2610 ;
        RECT 5.2380 23.5920 5.2560 24.5275 ;
        RECT 5.2020 23.5920 5.2200 24.5275 ;
        RECT 5.1660 24.1690 5.1840 24.4915 ;
        RECT 5.0490 24.3660 5.0670 24.4755 ;
        RECT 5.0400 23.6245 5.0580 23.8640 ;
        RECT 5.0040 24.2055 5.0220 24.3590 ;
        RECT 4.9230 24.2310 4.9410 24.4890 ;
        RECT 4.3830 23.5920 4.4010 24.5275 ;
        RECT 4.3470 23.5920 4.3650 24.5275 ;
        RECT 4.3110 23.7730 4.3290 24.3410 ;
        RECT 5.2380 24.6720 5.2560 25.6075 ;
        RECT 5.2020 24.6720 5.2200 25.6075 ;
        RECT 5.1660 25.2490 5.1840 25.5715 ;
        RECT 5.0490 25.4460 5.0670 25.5555 ;
        RECT 5.0400 24.7045 5.0580 24.9440 ;
        RECT 5.0040 25.2855 5.0220 25.4390 ;
        RECT 4.9230 25.3110 4.9410 25.5690 ;
        RECT 4.3830 24.6720 4.4010 25.6075 ;
        RECT 4.3470 24.6720 4.3650 25.6075 ;
        RECT 4.3110 24.8530 4.3290 25.4210 ;
  LAYER M3 SPACING 0.018  ;
      RECT 5.1800 0.2565 5.3080 1.3500 ;
      RECT 5.1660 0.9220 5.3080 1.2445 ;
      RECT 5.0180 0.6490 5.0800 1.3500 ;
      RECT 5.0040 0.9585 5.0800 1.1120 ;
      RECT 5.0180 0.2565 5.0440 1.3500 ;
      RECT 5.0180 0.3775 5.0580 0.6170 ;
      RECT 5.0180 0.2565 5.0800 0.3455 ;
      RECT 4.7210 0.7070 4.9270 1.3500 ;
      RECT 4.9010 0.2565 4.9270 1.3500 ;
      RECT 4.7210 0.9840 4.9410 1.2420 ;
      RECT 4.7210 0.2565 4.8190 1.3500 ;
      RECT 4.3040 0.2565 4.3870 1.3500 ;
      RECT 4.3040 0.3450 4.4010 1.2805 ;
      RECT 9.5270 0.2565 9.6120 1.3500 ;
      RECT 9.3830 0.2565 9.4090 1.3500 ;
      RECT 9.2750 0.2565 9.3010 1.3500 ;
      RECT 9.1670 0.2565 9.1930 1.3500 ;
      RECT 9.0590 0.2565 9.0850 1.3500 ;
      RECT 8.9510 0.2565 8.9770 1.3500 ;
      RECT 8.8430 0.2565 8.8690 1.3500 ;
      RECT 8.7350 0.2565 8.7610 1.3500 ;
      RECT 8.6270 0.2565 8.6530 1.3500 ;
      RECT 8.5190 0.2565 8.5450 1.3500 ;
      RECT 8.4110 0.2565 8.4370 1.3500 ;
      RECT 8.3030 0.2565 8.3290 1.3500 ;
      RECT 8.1950 0.2565 8.2210 1.3500 ;
      RECT 8.0870 0.2565 8.1130 1.3500 ;
      RECT 7.9790 0.2565 8.0050 1.3500 ;
      RECT 7.8710 0.2565 7.8970 1.3500 ;
      RECT 7.7630 0.2565 7.7890 1.3500 ;
      RECT 7.6550 0.2565 7.6810 1.3500 ;
      RECT 7.5470 0.2565 7.5730 1.3500 ;
      RECT 7.4390 0.2565 7.4650 1.3500 ;
      RECT 7.3310 0.2565 7.3570 1.3500 ;
      RECT 7.2230 0.2565 7.2490 1.3500 ;
      RECT 7.1150 0.2565 7.1410 1.3500 ;
      RECT 7.0070 0.2565 7.0330 1.3500 ;
      RECT 6.8990 0.2565 6.9250 1.3500 ;
      RECT 6.7910 0.2565 6.8170 1.3500 ;
      RECT 6.6830 0.2565 6.7090 1.3500 ;
      RECT 6.5750 0.2565 6.6010 1.3500 ;
      RECT 6.4670 0.2565 6.4930 1.3500 ;
      RECT 6.3590 0.2565 6.3850 1.3500 ;
      RECT 6.2510 0.2565 6.2770 1.3500 ;
      RECT 6.1430 0.2565 6.1690 1.3500 ;
      RECT 6.0350 0.2565 6.0610 1.3500 ;
      RECT 5.9270 0.2565 5.9530 1.3500 ;
      RECT 5.7140 0.2565 5.7910 1.3500 ;
      RECT 3.8210 0.2565 3.8980 1.3500 ;
      RECT 3.6590 0.2565 3.6850 1.3500 ;
      RECT 3.5510 0.2565 3.5770 1.3500 ;
      RECT 3.4430 0.2565 3.4690 1.3500 ;
      RECT 3.3350 0.2565 3.3610 1.3500 ;
      RECT 3.2270 0.2565 3.2530 1.3500 ;
      RECT 3.1190 0.2565 3.1450 1.3500 ;
      RECT 3.0110 0.2565 3.0370 1.3500 ;
      RECT 2.9030 0.2565 2.9290 1.3500 ;
      RECT 2.7950 0.2565 2.8210 1.3500 ;
      RECT 2.6870 0.2565 2.7130 1.3500 ;
      RECT 2.5790 0.2565 2.6050 1.3500 ;
      RECT 2.4710 0.2565 2.4970 1.3500 ;
      RECT 2.3630 0.2565 2.3890 1.3500 ;
      RECT 2.2550 0.2565 2.2810 1.3500 ;
      RECT 2.1470 0.2565 2.1730 1.3500 ;
      RECT 2.0390 0.2565 2.0650 1.3500 ;
      RECT 1.9310 0.2565 1.9570 1.3500 ;
      RECT 1.8230 0.2565 1.8490 1.3500 ;
      RECT 1.7150 0.2565 1.7410 1.3500 ;
      RECT 1.6070 0.2565 1.6330 1.3500 ;
      RECT 1.4990 0.2565 1.5250 1.3500 ;
      RECT 1.3910 0.2565 1.4170 1.3500 ;
      RECT 1.2830 0.2565 1.3090 1.3500 ;
      RECT 1.1750 0.2565 1.2010 1.3500 ;
      RECT 1.0670 0.2565 1.0930 1.3500 ;
      RECT 0.9590 0.2565 0.9850 1.3500 ;
      RECT 0.8510 0.2565 0.8770 1.3500 ;
      RECT 0.7430 0.2565 0.7690 1.3500 ;
      RECT 0.6350 0.2565 0.6610 1.3500 ;
      RECT 0.5270 0.2565 0.5530 1.3500 ;
      RECT 0.4190 0.2565 0.4450 1.3500 ;
      RECT 0.3110 0.2565 0.3370 1.3500 ;
      RECT 0.2030 0.2565 0.2290 1.3500 ;
      RECT 0.0000 0.2565 0.0850 1.3500 ;
      RECT 5.1800 1.3365 5.3080 2.4300 ;
      RECT 5.1660 2.0020 5.3080 2.3245 ;
      RECT 5.0180 1.7290 5.0800 2.4300 ;
      RECT 5.0040 2.0385 5.0800 2.1920 ;
      RECT 5.0180 1.3365 5.0440 2.4300 ;
      RECT 5.0180 1.4575 5.0580 1.6970 ;
      RECT 5.0180 1.3365 5.0800 1.4255 ;
      RECT 4.7210 1.7870 4.9270 2.4300 ;
      RECT 4.9010 1.3365 4.9270 2.4300 ;
      RECT 4.7210 2.0640 4.9410 2.3220 ;
      RECT 4.7210 1.3365 4.8190 2.4300 ;
      RECT 4.3040 1.3365 4.3870 2.4300 ;
      RECT 4.3040 1.4250 4.4010 2.3605 ;
      RECT 9.5270 1.3365 9.6120 2.4300 ;
      RECT 9.3830 1.3365 9.4090 2.4300 ;
      RECT 9.2750 1.3365 9.3010 2.4300 ;
      RECT 9.1670 1.3365 9.1930 2.4300 ;
      RECT 9.0590 1.3365 9.0850 2.4300 ;
      RECT 8.9510 1.3365 8.9770 2.4300 ;
      RECT 8.8430 1.3365 8.8690 2.4300 ;
      RECT 8.7350 1.3365 8.7610 2.4300 ;
      RECT 8.6270 1.3365 8.6530 2.4300 ;
      RECT 8.5190 1.3365 8.5450 2.4300 ;
      RECT 8.4110 1.3365 8.4370 2.4300 ;
      RECT 8.3030 1.3365 8.3290 2.4300 ;
      RECT 8.1950 1.3365 8.2210 2.4300 ;
      RECT 8.0870 1.3365 8.1130 2.4300 ;
      RECT 7.9790 1.3365 8.0050 2.4300 ;
      RECT 7.8710 1.3365 7.8970 2.4300 ;
      RECT 7.7630 1.3365 7.7890 2.4300 ;
      RECT 7.6550 1.3365 7.6810 2.4300 ;
      RECT 7.5470 1.3365 7.5730 2.4300 ;
      RECT 7.4390 1.3365 7.4650 2.4300 ;
      RECT 7.3310 1.3365 7.3570 2.4300 ;
      RECT 7.2230 1.3365 7.2490 2.4300 ;
      RECT 7.1150 1.3365 7.1410 2.4300 ;
      RECT 7.0070 1.3365 7.0330 2.4300 ;
      RECT 6.8990 1.3365 6.9250 2.4300 ;
      RECT 6.7910 1.3365 6.8170 2.4300 ;
      RECT 6.6830 1.3365 6.7090 2.4300 ;
      RECT 6.5750 1.3365 6.6010 2.4300 ;
      RECT 6.4670 1.3365 6.4930 2.4300 ;
      RECT 6.3590 1.3365 6.3850 2.4300 ;
      RECT 6.2510 1.3365 6.2770 2.4300 ;
      RECT 6.1430 1.3365 6.1690 2.4300 ;
      RECT 6.0350 1.3365 6.0610 2.4300 ;
      RECT 5.9270 1.3365 5.9530 2.4300 ;
      RECT 5.7140 1.3365 5.7910 2.4300 ;
      RECT 3.8210 1.3365 3.8980 2.4300 ;
      RECT 3.6590 1.3365 3.6850 2.4300 ;
      RECT 3.5510 1.3365 3.5770 2.4300 ;
      RECT 3.4430 1.3365 3.4690 2.4300 ;
      RECT 3.3350 1.3365 3.3610 2.4300 ;
      RECT 3.2270 1.3365 3.2530 2.4300 ;
      RECT 3.1190 1.3365 3.1450 2.4300 ;
      RECT 3.0110 1.3365 3.0370 2.4300 ;
      RECT 2.9030 1.3365 2.9290 2.4300 ;
      RECT 2.7950 1.3365 2.8210 2.4300 ;
      RECT 2.6870 1.3365 2.7130 2.4300 ;
      RECT 2.5790 1.3365 2.6050 2.4300 ;
      RECT 2.4710 1.3365 2.4970 2.4300 ;
      RECT 2.3630 1.3365 2.3890 2.4300 ;
      RECT 2.2550 1.3365 2.2810 2.4300 ;
      RECT 2.1470 1.3365 2.1730 2.4300 ;
      RECT 2.0390 1.3365 2.0650 2.4300 ;
      RECT 1.9310 1.3365 1.9570 2.4300 ;
      RECT 1.8230 1.3365 1.8490 2.4300 ;
      RECT 1.7150 1.3365 1.7410 2.4300 ;
      RECT 1.6070 1.3365 1.6330 2.4300 ;
      RECT 1.4990 1.3365 1.5250 2.4300 ;
      RECT 1.3910 1.3365 1.4170 2.4300 ;
      RECT 1.2830 1.3365 1.3090 2.4300 ;
      RECT 1.1750 1.3365 1.2010 2.4300 ;
      RECT 1.0670 1.3365 1.0930 2.4300 ;
      RECT 0.9590 1.3365 0.9850 2.4300 ;
      RECT 0.8510 1.3365 0.8770 2.4300 ;
      RECT 0.7430 1.3365 0.7690 2.4300 ;
      RECT 0.6350 1.3365 0.6610 2.4300 ;
      RECT 0.5270 1.3365 0.5530 2.4300 ;
      RECT 0.4190 1.3365 0.4450 2.4300 ;
      RECT 0.3110 1.3365 0.3370 2.4300 ;
      RECT 0.2030 1.3365 0.2290 2.4300 ;
      RECT 0.0000 1.3365 0.0850 2.4300 ;
      RECT 5.1800 2.4165 5.3080 3.5100 ;
      RECT 5.1660 3.0820 5.3080 3.4045 ;
      RECT 5.0180 2.8090 5.0800 3.5100 ;
      RECT 5.0040 3.1185 5.0800 3.2720 ;
      RECT 5.0180 2.4165 5.0440 3.5100 ;
      RECT 5.0180 2.5375 5.0580 2.7770 ;
      RECT 5.0180 2.4165 5.0800 2.5055 ;
      RECT 4.7210 2.8670 4.9270 3.5100 ;
      RECT 4.9010 2.4165 4.9270 3.5100 ;
      RECT 4.7210 3.1440 4.9410 3.4020 ;
      RECT 4.7210 2.4165 4.8190 3.5100 ;
      RECT 4.3040 2.4165 4.3870 3.5100 ;
      RECT 4.3040 2.5050 4.4010 3.4405 ;
      RECT 9.5270 2.4165 9.6120 3.5100 ;
      RECT 9.3830 2.4165 9.4090 3.5100 ;
      RECT 9.2750 2.4165 9.3010 3.5100 ;
      RECT 9.1670 2.4165 9.1930 3.5100 ;
      RECT 9.0590 2.4165 9.0850 3.5100 ;
      RECT 8.9510 2.4165 8.9770 3.5100 ;
      RECT 8.8430 2.4165 8.8690 3.5100 ;
      RECT 8.7350 2.4165 8.7610 3.5100 ;
      RECT 8.6270 2.4165 8.6530 3.5100 ;
      RECT 8.5190 2.4165 8.5450 3.5100 ;
      RECT 8.4110 2.4165 8.4370 3.5100 ;
      RECT 8.3030 2.4165 8.3290 3.5100 ;
      RECT 8.1950 2.4165 8.2210 3.5100 ;
      RECT 8.0870 2.4165 8.1130 3.5100 ;
      RECT 7.9790 2.4165 8.0050 3.5100 ;
      RECT 7.8710 2.4165 7.8970 3.5100 ;
      RECT 7.7630 2.4165 7.7890 3.5100 ;
      RECT 7.6550 2.4165 7.6810 3.5100 ;
      RECT 7.5470 2.4165 7.5730 3.5100 ;
      RECT 7.4390 2.4165 7.4650 3.5100 ;
      RECT 7.3310 2.4165 7.3570 3.5100 ;
      RECT 7.2230 2.4165 7.2490 3.5100 ;
      RECT 7.1150 2.4165 7.1410 3.5100 ;
      RECT 7.0070 2.4165 7.0330 3.5100 ;
      RECT 6.8990 2.4165 6.9250 3.5100 ;
      RECT 6.7910 2.4165 6.8170 3.5100 ;
      RECT 6.6830 2.4165 6.7090 3.5100 ;
      RECT 6.5750 2.4165 6.6010 3.5100 ;
      RECT 6.4670 2.4165 6.4930 3.5100 ;
      RECT 6.3590 2.4165 6.3850 3.5100 ;
      RECT 6.2510 2.4165 6.2770 3.5100 ;
      RECT 6.1430 2.4165 6.1690 3.5100 ;
      RECT 6.0350 2.4165 6.0610 3.5100 ;
      RECT 5.9270 2.4165 5.9530 3.5100 ;
      RECT 5.7140 2.4165 5.7910 3.5100 ;
      RECT 3.8210 2.4165 3.8980 3.5100 ;
      RECT 3.6590 2.4165 3.6850 3.5100 ;
      RECT 3.5510 2.4165 3.5770 3.5100 ;
      RECT 3.4430 2.4165 3.4690 3.5100 ;
      RECT 3.3350 2.4165 3.3610 3.5100 ;
      RECT 3.2270 2.4165 3.2530 3.5100 ;
      RECT 3.1190 2.4165 3.1450 3.5100 ;
      RECT 3.0110 2.4165 3.0370 3.5100 ;
      RECT 2.9030 2.4165 2.9290 3.5100 ;
      RECT 2.7950 2.4165 2.8210 3.5100 ;
      RECT 2.6870 2.4165 2.7130 3.5100 ;
      RECT 2.5790 2.4165 2.6050 3.5100 ;
      RECT 2.4710 2.4165 2.4970 3.5100 ;
      RECT 2.3630 2.4165 2.3890 3.5100 ;
      RECT 2.2550 2.4165 2.2810 3.5100 ;
      RECT 2.1470 2.4165 2.1730 3.5100 ;
      RECT 2.0390 2.4165 2.0650 3.5100 ;
      RECT 1.9310 2.4165 1.9570 3.5100 ;
      RECT 1.8230 2.4165 1.8490 3.5100 ;
      RECT 1.7150 2.4165 1.7410 3.5100 ;
      RECT 1.6070 2.4165 1.6330 3.5100 ;
      RECT 1.4990 2.4165 1.5250 3.5100 ;
      RECT 1.3910 2.4165 1.4170 3.5100 ;
      RECT 1.2830 2.4165 1.3090 3.5100 ;
      RECT 1.1750 2.4165 1.2010 3.5100 ;
      RECT 1.0670 2.4165 1.0930 3.5100 ;
      RECT 0.9590 2.4165 0.9850 3.5100 ;
      RECT 0.8510 2.4165 0.8770 3.5100 ;
      RECT 0.7430 2.4165 0.7690 3.5100 ;
      RECT 0.6350 2.4165 0.6610 3.5100 ;
      RECT 0.5270 2.4165 0.5530 3.5100 ;
      RECT 0.4190 2.4165 0.4450 3.5100 ;
      RECT 0.3110 2.4165 0.3370 3.5100 ;
      RECT 0.2030 2.4165 0.2290 3.5100 ;
      RECT 0.0000 2.4165 0.0850 3.5100 ;
      RECT 5.1800 3.4965 5.3080 4.5900 ;
      RECT 5.1660 4.1620 5.3080 4.4845 ;
      RECT 5.0180 3.8890 5.0800 4.5900 ;
      RECT 5.0040 4.1985 5.0800 4.3520 ;
      RECT 5.0180 3.4965 5.0440 4.5900 ;
      RECT 5.0180 3.6175 5.0580 3.8570 ;
      RECT 5.0180 3.4965 5.0800 3.5855 ;
      RECT 4.7210 3.9470 4.9270 4.5900 ;
      RECT 4.9010 3.4965 4.9270 4.5900 ;
      RECT 4.7210 4.2240 4.9410 4.4820 ;
      RECT 4.7210 3.4965 4.8190 4.5900 ;
      RECT 4.3040 3.4965 4.3870 4.5900 ;
      RECT 4.3040 3.5850 4.4010 4.5205 ;
      RECT 9.5270 3.4965 9.6120 4.5900 ;
      RECT 9.3830 3.4965 9.4090 4.5900 ;
      RECT 9.2750 3.4965 9.3010 4.5900 ;
      RECT 9.1670 3.4965 9.1930 4.5900 ;
      RECT 9.0590 3.4965 9.0850 4.5900 ;
      RECT 8.9510 3.4965 8.9770 4.5900 ;
      RECT 8.8430 3.4965 8.8690 4.5900 ;
      RECT 8.7350 3.4965 8.7610 4.5900 ;
      RECT 8.6270 3.4965 8.6530 4.5900 ;
      RECT 8.5190 3.4965 8.5450 4.5900 ;
      RECT 8.4110 3.4965 8.4370 4.5900 ;
      RECT 8.3030 3.4965 8.3290 4.5900 ;
      RECT 8.1950 3.4965 8.2210 4.5900 ;
      RECT 8.0870 3.4965 8.1130 4.5900 ;
      RECT 7.9790 3.4965 8.0050 4.5900 ;
      RECT 7.8710 3.4965 7.8970 4.5900 ;
      RECT 7.7630 3.4965 7.7890 4.5900 ;
      RECT 7.6550 3.4965 7.6810 4.5900 ;
      RECT 7.5470 3.4965 7.5730 4.5900 ;
      RECT 7.4390 3.4965 7.4650 4.5900 ;
      RECT 7.3310 3.4965 7.3570 4.5900 ;
      RECT 7.2230 3.4965 7.2490 4.5900 ;
      RECT 7.1150 3.4965 7.1410 4.5900 ;
      RECT 7.0070 3.4965 7.0330 4.5900 ;
      RECT 6.8990 3.4965 6.9250 4.5900 ;
      RECT 6.7910 3.4965 6.8170 4.5900 ;
      RECT 6.6830 3.4965 6.7090 4.5900 ;
      RECT 6.5750 3.4965 6.6010 4.5900 ;
      RECT 6.4670 3.4965 6.4930 4.5900 ;
      RECT 6.3590 3.4965 6.3850 4.5900 ;
      RECT 6.2510 3.4965 6.2770 4.5900 ;
      RECT 6.1430 3.4965 6.1690 4.5900 ;
      RECT 6.0350 3.4965 6.0610 4.5900 ;
      RECT 5.9270 3.4965 5.9530 4.5900 ;
      RECT 5.7140 3.4965 5.7910 4.5900 ;
      RECT 3.8210 3.4965 3.8980 4.5900 ;
      RECT 3.6590 3.4965 3.6850 4.5900 ;
      RECT 3.5510 3.4965 3.5770 4.5900 ;
      RECT 3.4430 3.4965 3.4690 4.5900 ;
      RECT 3.3350 3.4965 3.3610 4.5900 ;
      RECT 3.2270 3.4965 3.2530 4.5900 ;
      RECT 3.1190 3.4965 3.1450 4.5900 ;
      RECT 3.0110 3.4965 3.0370 4.5900 ;
      RECT 2.9030 3.4965 2.9290 4.5900 ;
      RECT 2.7950 3.4965 2.8210 4.5900 ;
      RECT 2.6870 3.4965 2.7130 4.5900 ;
      RECT 2.5790 3.4965 2.6050 4.5900 ;
      RECT 2.4710 3.4965 2.4970 4.5900 ;
      RECT 2.3630 3.4965 2.3890 4.5900 ;
      RECT 2.2550 3.4965 2.2810 4.5900 ;
      RECT 2.1470 3.4965 2.1730 4.5900 ;
      RECT 2.0390 3.4965 2.0650 4.5900 ;
      RECT 1.9310 3.4965 1.9570 4.5900 ;
      RECT 1.8230 3.4965 1.8490 4.5900 ;
      RECT 1.7150 3.4965 1.7410 4.5900 ;
      RECT 1.6070 3.4965 1.6330 4.5900 ;
      RECT 1.4990 3.4965 1.5250 4.5900 ;
      RECT 1.3910 3.4965 1.4170 4.5900 ;
      RECT 1.2830 3.4965 1.3090 4.5900 ;
      RECT 1.1750 3.4965 1.2010 4.5900 ;
      RECT 1.0670 3.4965 1.0930 4.5900 ;
      RECT 0.9590 3.4965 0.9850 4.5900 ;
      RECT 0.8510 3.4965 0.8770 4.5900 ;
      RECT 0.7430 3.4965 0.7690 4.5900 ;
      RECT 0.6350 3.4965 0.6610 4.5900 ;
      RECT 0.5270 3.4965 0.5530 4.5900 ;
      RECT 0.4190 3.4965 0.4450 4.5900 ;
      RECT 0.3110 3.4965 0.3370 4.5900 ;
      RECT 0.2030 3.4965 0.2290 4.5900 ;
      RECT 0.0000 3.4965 0.0850 4.5900 ;
      RECT 5.1800 4.5765 5.3080 5.6700 ;
      RECT 5.1660 5.2420 5.3080 5.5645 ;
      RECT 5.0180 4.9690 5.0800 5.6700 ;
      RECT 5.0040 5.2785 5.0800 5.4320 ;
      RECT 5.0180 4.5765 5.0440 5.6700 ;
      RECT 5.0180 4.6975 5.0580 4.9370 ;
      RECT 5.0180 4.5765 5.0800 4.6655 ;
      RECT 4.7210 5.0270 4.9270 5.6700 ;
      RECT 4.9010 4.5765 4.9270 5.6700 ;
      RECT 4.7210 5.3040 4.9410 5.5620 ;
      RECT 4.7210 4.5765 4.8190 5.6700 ;
      RECT 4.3040 4.5765 4.3870 5.6700 ;
      RECT 4.3040 4.6650 4.4010 5.6005 ;
      RECT 9.5270 4.5765 9.6120 5.6700 ;
      RECT 9.3830 4.5765 9.4090 5.6700 ;
      RECT 9.2750 4.5765 9.3010 5.6700 ;
      RECT 9.1670 4.5765 9.1930 5.6700 ;
      RECT 9.0590 4.5765 9.0850 5.6700 ;
      RECT 8.9510 4.5765 8.9770 5.6700 ;
      RECT 8.8430 4.5765 8.8690 5.6700 ;
      RECT 8.7350 4.5765 8.7610 5.6700 ;
      RECT 8.6270 4.5765 8.6530 5.6700 ;
      RECT 8.5190 4.5765 8.5450 5.6700 ;
      RECT 8.4110 4.5765 8.4370 5.6700 ;
      RECT 8.3030 4.5765 8.3290 5.6700 ;
      RECT 8.1950 4.5765 8.2210 5.6700 ;
      RECT 8.0870 4.5765 8.1130 5.6700 ;
      RECT 7.9790 4.5765 8.0050 5.6700 ;
      RECT 7.8710 4.5765 7.8970 5.6700 ;
      RECT 7.7630 4.5765 7.7890 5.6700 ;
      RECT 7.6550 4.5765 7.6810 5.6700 ;
      RECT 7.5470 4.5765 7.5730 5.6700 ;
      RECT 7.4390 4.5765 7.4650 5.6700 ;
      RECT 7.3310 4.5765 7.3570 5.6700 ;
      RECT 7.2230 4.5765 7.2490 5.6700 ;
      RECT 7.1150 4.5765 7.1410 5.6700 ;
      RECT 7.0070 4.5765 7.0330 5.6700 ;
      RECT 6.8990 4.5765 6.9250 5.6700 ;
      RECT 6.7910 4.5765 6.8170 5.6700 ;
      RECT 6.6830 4.5765 6.7090 5.6700 ;
      RECT 6.5750 4.5765 6.6010 5.6700 ;
      RECT 6.4670 4.5765 6.4930 5.6700 ;
      RECT 6.3590 4.5765 6.3850 5.6700 ;
      RECT 6.2510 4.5765 6.2770 5.6700 ;
      RECT 6.1430 4.5765 6.1690 5.6700 ;
      RECT 6.0350 4.5765 6.0610 5.6700 ;
      RECT 5.9270 4.5765 5.9530 5.6700 ;
      RECT 5.7140 4.5765 5.7910 5.6700 ;
      RECT 3.8210 4.5765 3.8980 5.6700 ;
      RECT 3.6590 4.5765 3.6850 5.6700 ;
      RECT 3.5510 4.5765 3.5770 5.6700 ;
      RECT 3.4430 4.5765 3.4690 5.6700 ;
      RECT 3.3350 4.5765 3.3610 5.6700 ;
      RECT 3.2270 4.5765 3.2530 5.6700 ;
      RECT 3.1190 4.5765 3.1450 5.6700 ;
      RECT 3.0110 4.5765 3.0370 5.6700 ;
      RECT 2.9030 4.5765 2.9290 5.6700 ;
      RECT 2.7950 4.5765 2.8210 5.6700 ;
      RECT 2.6870 4.5765 2.7130 5.6700 ;
      RECT 2.5790 4.5765 2.6050 5.6700 ;
      RECT 2.4710 4.5765 2.4970 5.6700 ;
      RECT 2.3630 4.5765 2.3890 5.6700 ;
      RECT 2.2550 4.5765 2.2810 5.6700 ;
      RECT 2.1470 4.5765 2.1730 5.6700 ;
      RECT 2.0390 4.5765 2.0650 5.6700 ;
      RECT 1.9310 4.5765 1.9570 5.6700 ;
      RECT 1.8230 4.5765 1.8490 5.6700 ;
      RECT 1.7150 4.5765 1.7410 5.6700 ;
      RECT 1.6070 4.5765 1.6330 5.6700 ;
      RECT 1.4990 4.5765 1.5250 5.6700 ;
      RECT 1.3910 4.5765 1.4170 5.6700 ;
      RECT 1.2830 4.5765 1.3090 5.6700 ;
      RECT 1.1750 4.5765 1.2010 5.6700 ;
      RECT 1.0670 4.5765 1.0930 5.6700 ;
      RECT 0.9590 4.5765 0.9850 5.6700 ;
      RECT 0.8510 4.5765 0.8770 5.6700 ;
      RECT 0.7430 4.5765 0.7690 5.6700 ;
      RECT 0.6350 4.5765 0.6610 5.6700 ;
      RECT 0.5270 4.5765 0.5530 5.6700 ;
      RECT 0.4190 4.5765 0.4450 5.6700 ;
      RECT 0.3110 4.5765 0.3370 5.6700 ;
      RECT 0.2030 4.5765 0.2290 5.6700 ;
      RECT 0.0000 4.5765 0.0850 5.6700 ;
      RECT 5.1800 5.6565 5.3080 6.7500 ;
      RECT 5.1660 6.3220 5.3080 6.6445 ;
      RECT 5.0180 6.0490 5.0800 6.7500 ;
      RECT 5.0040 6.3585 5.0800 6.5120 ;
      RECT 5.0180 5.6565 5.0440 6.7500 ;
      RECT 5.0180 5.7775 5.0580 6.0170 ;
      RECT 5.0180 5.6565 5.0800 5.7455 ;
      RECT 4.7210 6.1070 4.9270 6.7500 ;
      RECT 4.9010 5.6565 4.9270 6.7500 ;
      RECT 4.7210 6.3840 4.9410 6.6420 ;
      RECT 4.7210 5.6565 4.8190 6.7500 ;
      RECT 4.3040 5.6565 4.3870 6.7500 ;
      RECT 4.3040 5.7450 4.4010 6.6805 ;
      RECT 9.5270 5.6565 9.6120 6.7500 ;
      RECT 9.3830 5.6565 9.4090 6.7500 ;
      RECT 9.2750 5.6565 9.3010 6.7500 ;
      RECT 9.1670 5.6565 9.1930 6.7500 ;
      RECT 9.0590 5.6565 9.0850 6.7500 ;
      RECT 8.9510 5.6565 8.9770 6.7500 ;
      RECT 8.8430 5.6565 8.8690 6.7500 ;
      RECT 8.7350 5.6565 8.7610 6.7500 ;
      RECT 8.6270 5.6565 8.6530 6.7500 ;
      RECT 8.5190 5.6565 8.5450 6.7500 ;
      RECT 8.4110 5.6565 8.4370 6.7500 ;
      RECT 8.3030 5.6565 8.3290 6.7500 ;
      RECT 8.1950 5.6565 8.2210 6.7500 ;
      RECT 8.0870 5.6565 8.1130 6.7500 ;
      RECT 7.9790 5.6565 8.0050 6.7500 ;
      RECT 7.8710 5.6565 7.8970 6.7500 ;
      RECT 7.7630 5.6565 7.7890 6.7500 ;
      RECT 7.6550 5.6565 7.6810 6.7500 ;
      RECT 7.5470 5.6565 7.5730 6.7500 ;
      RECT 7.4390 5.6565 7.4650 6.7500 ;
      RECT 7.3310 5.6565 7.3570 6.7500 ;
      RECT 7.2230 5.6565 7.2490 6.7500 ;
      RECT 7.1150 5.6565 7.1410 6.7500 ;
      RECT 7.0070 5.6565 7.0330 6.7500 ;
      RECT 6.8990 5.6565 6.9250 6.7500 ;
      RECT 6.7910 5.6565 6.8170 6.7500 ;
      RECT 6.6830 5.6565 6.7090 6.7500 ;
      RECT 6.5750 5.6565 6.6010 6.7500 ;
      RECT 6.4670 5.6565 6.4930 6.7500 ;
      RECT 6.3590 5.6565 6.3850 6.7500 ;
      RECT 6.2510 5.6565 6.2770 6.7500 ;
      RECT 6.1430 5.6565 6.1690 6.7500 ;
      RECT 6.0350 5.6565 6.0610 6.7500 ;
      RECT 5.9270 5.6565 5.9530 6.7500 ;
      RECT 5.7140 5.6565 5.7910 6.7500 ;
      RECT 3.8210 5.6565 3.8980 6.7500 ;
      RECT 3.6590 5.6565 3.6850 6.7500 ;
      RECT 3.5510 5.6565 3.5770 6.7500 ;
      RECT 3.4430 5.6565 3.4690 6.7500 ;
      RECT 3.3350 5.6565 3.3610 6.7500 ;
      RECT 3.2270 5.6565 3.2530 6.7500 ;
      RECT 3.1190 5.6565 3.1450 6.7500 ;
      RECT 3.0110 5.6565 3.0370 6.7500 ;
      RECT 2.9030 5.6565 2.9290 6.7500 ;
      RECT 2.7950 5.6565 2.8210 6.7500 ;
      RECT 2.6870 5.6565 2.7130 6.7500 ;
      RECT 2.5790 5.6565 2.6050 6.7500 ;
      RECT 2.4710 5.6565 2.4970 6.7500 ;
      RECT 2.3630 5.6565 2.3890 6.7500 ;
      RECT 2.2550 5.6565 2.2810 6.7500 ;
      RECT 2.1470 5.6565 2.1730 6.7500 ;
      RECT 2.0390 5.6565 2.0650 6.7500 ;
      RECT 1.9310 5.6565 1.9570 6.7500 ;
      RECT 1.8230 5.6565 1.8490 6.7500 ;
      RECT 1.7150 5.6565 1.7410 6.7500 ;
      RECT 1.6070 5.6565 1.6330 6.7500 ;
      RECT 1.4990 5.6565 1.5250 6.7500 ;
      RECT 1.3910 5.6565 1.4170 6.7500 ;
      RECT 1.2830 5.6565 1.3090 6.7500 ;
      RECT 1.1750 5.6565 1.2010 6.7500 ;
      RECT 1.0670 5.6565 1.0930 6.7500 ;
      RECT 0.9590 5.6565 0.9850 6.7500 ;
      RECT 0.8510 5.6565 0.8770 6.7500 ;
      RECT 0.7430 5.6565 0.7690 6.7500 ;
      RECT 0.6350 5.6565 0.6610 6.7500 ;
      RECT 0.5270 5.6565 0.5530 6.7500 ;
      RECT 0.4190 5.6565 0.4450 6.7500 ;
      RECT 0.3110 5.6565 0.3370 6.7500 ;
      RECT 0.2030 5.6565 0.2290 6.7500 ;
      RECT 0.0000 5.6565 0.0850 6.7500 ;
      RECT 5.1800 6.7365 5.3080 7.8300 ;
      RECT 5.1660 7.4020 5.3080 7.7245 ;
      RECT 5.0180 7.1290 5.0800 7.8300 ;
      RECT 5.0040 7.4385 5.0800 7.5920 ;
      RECT 5.0180 6.7365 5.0440 7.8300 ;
      RECT 5.0180 6.8575 5.0580 7.0970 ;
      RECT 5.0180 6.7365 5.0800 6.8255 ;
      RECT 4.7210 7.1870 4.9270 7.8300 ;
      RECT 4.9010 6.7365 4.9270 7.8300 ;
      RECT 4.7210 7.4640 4.9410 7.7220 ;
      RECT 4.7210 6.7365 4.8190 7.8300 ;
      RECT 4.3040 6.7365 4.3870 7.8300 ;
      RECT 4.3040 6.8250 4.4010 7.7605 ;
      RECT 9.5270 6.7365 9.6120 7.8300 ;
      RECT 9.3830 6.7365 9.4090 7.8300 ;
      RECT 9.2750 6.7365 9.3010 7.8300 ;
      RECT 9.1670 6.7365 9.1930 7.8300 ;
      RECT 9.0590 6.7365 9.0850 7.8300 ;
      RECT 8.9510 6.7365 8.9770 7.8300 ;
      RECT 8.8430 6.7365 8.8690 7.8300 ;
      RECT 8.7350 6.7365 8.7610 7.8300 ;
      RECT 8.6270 6.7365 8.6530 7.8300 ;
      RECT 8.5190 6.7365 8.5450 7.8300 ;
      RECT 8.4110 6.7365 8.4370 7.8300 ;
      RECT 8.3030 6.7365 8.3290 7.8300 ;
      RECT 8.1950 6.7365 8.2210 7.8300 ;
      RECT 8.0870 6.7365 8.1130 7.8300 ;
      RECT 7.9790 6.7365 8.0050 7.8300 ;
      RECT 7.8710 6.7365 7.8970 7.8300 ;
      RECT 7.7630 6.7365 7.7890 7.8300 ;
      RECT 7.6550 6.7365 7.6810 7.8300 ;
      RECT 7.5470 6.7365 7.5730 7.8300 ;
      RECT 7.4390 6.7365 7.4650 7.8300 ;
      RECT 7.3310 6.7365 7.3570 7.8300 ;
      RECT 7.2230 6.7365 7.2490 7.8300 ;
      RECT 7.1150 6.7365 7.1410 7.8300 ;
      RECT 7.0070 6.7365 7.0330 7.8300 ;
      RECT 6.8990 6.7365 6.9250 7.8300 ;
      RECT 6.7910 6.7365 6.8170 7.8300 ;
      RECT 6.6830 6.7365 6.7090 7.8300 ;
      RECT 6.5750 6.7365 6.6010 7.8300 ;
      RECT 6.4670 6.7365 6.4930 7.8300 ;
      RECT 6.3590 6.7365 6.3850 7.8300 ;
      RECT 6.2510 6.7365 6.2770 7.8300 ;
      RECT 6.1430 6.7365 6.1690 7.8300 ;
      RECT 6.0350 6.7365 6.0610 7.8300 ;
      RECT 5.9270 6.7365 5.9530 7.8300 ;
      RECT 5.7140 6.7365 5.7910 7.8300 ;
      RECT 3.8210 6.7365 3.8980 7.8300 ;
      RECT 3.6590 6.7365 3.6850 7.8300 ;
      RECT 3.5510 6.7365 3.5770 7.8300 ;
      RECT 3.4430 6.7365 3.4690 7.8300 ;
      RECT 3.3350 6.7365 3.3610 7.8300 ;
      RECT 3.2270 6.7365 3.2530 7.8300 ;
      RECT 3.1190 6.7365 3.1450 7.8300 ;
      RECT 3.0110 6.7365 3.0370 7.8300 ;
      RECT 2.9030 6.7365 2.9290 7.8300 ;
      RECT 2.7950 6.7365 2.8210 7.8300 ;
      RECT 2.6870 6.7365 2.7130 7.8300 ;
      RECT 2.5790 6.7365 2.6050 7.8300 ;
      RECT 2.4710 6.7365 2.4970 7.8300 ;
      RECT 2.3630 6.7365 2.3890 7.8300 ;
      RECT 2.2550 6.7365 2.2810 7.8300 ;
      RECT 2.1470 6.7365 2.1730 7.8300 ;
      RECT 2.0390 6.7365 2.0650 7.8300 ;
      RECT 1.9310 6.7365 1.9570 7.8300 ;
      RECT 1.8230 6.7365 1.8490 7.8300 ;
      RECT 1.7150 6.7365 1.7410 7.8300 ;
      RECT 1.6070 6.7365 1.6330 7.8300 ;
      RECT 1.4990 6.7365 1.5250 7.8300 ;
      RECT 1.3910 6.7365 1.4170 7.8300 ;
      RECT 1.2830 6.7365 1.3090 7.8300 ;
      RECT 1.1750 6.7365 1.2010 7.8300 ;
      RECT 1.0670 6.7365 1.0930 7.8300 ;
      RECT 0.9590 6.7365 0.9850 7.8300 ;
      RECT 0.8510 6.7365 0.8770 7.8300 ;
      RECT 0.7430 6.7365 0.7690 7.8300 ;
      RECT 0.6350 6.7365 0.6610 7.8300 ;
      RECT 0.5270 6.7365 0.5530 7.8300 ;
      RECT 0.4190 6.7365 0.4450 7.8300 ;
      RECT 0.3110 6.7365 0.3370 7.8300 ;
      RECT 0.2030 6.7365 0.2290 7.8300 ;
      RECT 0.0000 6.7365 0.0850 7.8300 ;
      RECT 5.1800 7.8165 5.3080 8.9100 ;
      RECT 5.1660 8.4820 5.3080 8.8045 ;
      RECT 5.0180 8.2090 5.0800 8.9100 ;
      RECT 5.0040 8.5185 5.0800 8.6720 ;
      RECT 5.0180 7.8165 5.0440 8.9100 ;
      RECT 5.0180 7.9375 5.0580 8.1770 ;
      RECT 5.0180 7.8165 5.0800 7.9055 ;
      RECT 4.7210 8.2670 4.9270 8.9100 ;
      RECT 4.9010 7.8165 4.9270 8.9100 ;
      RECT 4.7210 8.5440 4.9410 8.8020 ;
      RECT 4.7210 7.8165 4.8190 8.9100 ;
      RECT 4.3040 7.8165 4.3870 8.9100 ;
      RECT 4.3040 7.9050 4.4010 8.8405 ;
      RECT 9.5270 7.8165 9.6120 8.9100 ;
      RECT 9.3830 7.8165 9.4090 8.9100 ;
      RECT 9.2750 7.8165 9.3010 8.9100 ;
      RECT 9.1670 7.8165 9.1930 8.9100 ;
      RECT 9.0590 7.8165 9.0850 8.9100 ;
      RECT 8.9510 7.8165 8.9770 8.9100 ;
      RECT 8.8430 7.8165 8.8690 8.9100 ;
      RECT 8.7350 7.8165 8.7610 8.9100 ;
      RECT 8.6270 7.8165 8.6530 8.9100 ;
      RECT 8.5190 7.8165 8.5450 8.9100 ;
      RECT 8.4110 7.8165 8.4370 8.9100 ;
      RECT 8.3030 7.8165 8.3290 8.9100 ;
      RECT 8.1950 7.8165 8.2210 8.9100 ;
      RECT 8.0870 7.8165 8.1130 8.9100 ;
      RECT 7.9790 7.8165 8.0050 8.9100 ;
      RECT 7.8710 7.8165 7.8970 8.9100 ;
      RECT 7.7630 7.8165 7.7890 8.9100 ;
      RECT 7.6550 7.8165 7.6810 8.9100 ;
      RECT 7.5470 7.8165 7.5730 8.9100 ;
      RECT 7.4390 7.8165 7.4650 8.9100 ;
      RECT 7.3310 7.8165 7.3570 8.9100 ;
      RECT 7.2230 7.8165 7.2490 8.9100 ;
      RECT 7.1150 7.8165 7.1410 8.9100 ;
      RECT 7.0070 7.8165 7.0330 8.9100 ;
      RECT 6.8990 7.8165 6.9250 8.9100 ;
      RECT 6.7910 7.8165 6.8170 8.9100 ;
      RECT 6.6830 7.8165 6.7090 8.9100 ;
      RECT 6.5750 7.8165 6.6010 8.9100 ;
      RECT 6.4670 7.8165 6.4930 8.9100 ;
      RECT 6.3590 7.8165 6.3850 8.9100 ;
      RECT 6.2510 7.8165 6.2770 8.9100 ;
      RECT 6.1430 7.8165 6.1690 8.9100 ;
      RECT 6.0350 7.8165 6.0610 8.9100 ;
      RECT 5.9270 7.8165 5.9530 8.9100 ;
      RECT 5.7140 7.8165 5.7910 8.9100 ;
      RECT 3.8210 7.8165 3.8980 8.9100 ;
      RECT 3.6590 7.8165 3.6850 8.9100 ;
      RECT 3.5510 7.8165 3.5770 8.9100 ;
      RECT 3.4430 7.8165 3.4690 8.9100 ;
      RECT 3.3350 7.8165 3.3610 8.9100 ;
      RECT 3.2270 7.8165 3.2530 8.9100 ;
      RECT 3.1190 7.8165 3.1450 8.9100 ;
      RECT 3.0110 7.8165 3.0370 8.9100 ;
      RECT 2.9030 7.8165 2.9290 8.9100 ;
      RECT 2.7950 7.8165 2.8210 8.9100 ;
      RECT 2.6870 7.8165 2.7130 8.9100 ;
      RECT 2.5790 7.8165 2.6050 8.9100 ;
      RECT 2.4710 7.8165 2.4970 8.9100 ;
      RECT 2.3630 7.8165 2.3890 8.9100 ;
      RECT 2.2550 7.8165 2.2810 8.9100 ;
      RECT 2.1470 7.8165 2.1730 8.9100 ;
      RECT 2.0390 7.8165 2.0650 8.9100 ;
      RECT 1.9310 7.8165 1.9570 8.9100 ;
      RECT 1.8230 7.8165 1.8490 8.9100 ;
      RECT 1.7150 7.8165 1.7410 8.9100 ;
      RECT 1.6070 7.8165 1.6330 8.9100 ;
      RECT 1.4990 7.8165 1.5250 8.9100 ;
      RECT 1.3910 7.8165 1.4170 8.9100 ;
      RECT 1.2830 7.8165 1.3090 8.9100 ;
      RECT 1.1750 7.8165 1.2010 8.9100 ;
      RECT 1.0670 7.8165 1.0930 8.9100 ;
      RECT 0.9590 7.8165 0.9850 8.9100 ;
      RECT 0.8510 7.8165 0.8770 8.9100 ;
      RECT 0.7430 7.8165 0.7690 8.9100 ;
      RECT 0.6350 7.8165 0.6610 8.9100 ;
      RECT 0.5270 7.8165 0.5530 8.9100 ;
      RECT 0.4190 7.8165 0.4450 8.9100 ;
      RECT 0.3110 7.8165 0.3370 8.9100 ;
      RECT 0.2030 7.8165 0.2290 8.9100 ;
      RECT 0.0000 7.8165 0.0850 8.9100 ;
      RECT 0.0000 17.2440 9.6120 17.5365 ;
      RECT 9.5270 8.8830 9.6120 17.5365 ;
      RECT 4.5410 17.0955 9.6120 17.5365 ;
      RECT 0.0000 17.0955 4.3870 17.5365 ;
      RECT 5.9270 10.3870 9.4090 17.5365 ;
      RECT 7.3850 8.8830 9.4090 17.5365 ;
      RECT 4.5410 17.0690 5.8450 17.5365 ;
      RECT 5.1800 17.0680 5.8450 17.5365 ;
      RECT 3.7670 10.4950 4.3870 17.5365 ;
      RECT 3.8210 9.6490 4.3870 17.5365 ;
      RECT 0.2030 10.1920 3.6850 17.5365 ;
      RECT 3.3890 8.8830 3.6850 17.5365 ;
      RECT 0.0000 8.8830 0.0850 17.5365 ;
      RECT 4.5410 17.0660 5.0800 17.5365 ;
      RECT 5.0180 16.7950 5.0800 17.5365 ;
      RECT 5.1800 16.7950 5.7910 17.5365 ;
      RECT 4.5410 16.7950 4.9270 17.5365 ;
      RECT 5.9130 12.6760 9.4090 17.0360 ;
      RECT 0.2030 12.6760 3.6990 17.0360 ;
      RECT 5.9130 12.6760 9.4230 17.0315 ;
      RECT 0.1890 12.6760 3.6990 17.0315 ;
      RECT 5.1890 9.6490 5.7910 17.5365 ;
      RECT 4.7210 9.5680 4.8910 17.5365 ;
      RECT 4.8290 8.8830 4.8910 17.5365 ;
      RECT 4.0370 9.4670 4.4230 16.6450 ;
      RECT 3.7670 16.6030 4.4370 16.6400 ;
      RECT 5.1750 15.5290 5.7910 16.6370 ;
      RECT 4.7070 16.3390 4.8910 16.5650 ;
      RECT 4.7210 15.7630 4.9050 16.0250 ;
      RECT 3.7670 15.5650 4.4370 16.0250 ;
      RECT 4.7070 15.0250 4.8910 15.4850 ;
      RECT 5.1750 12.9910 5.7910 15.3230 ;
      RECT 3.7670 13.6390 4.4370 14.7830 ;
      RECT 4.7210 13.3690 4.9050 14.6750 ;
      RECT 4.7070 13.9450 4.9050 14.4050 ;
      RECT 4.7070 10.7050 4.8910 13.8650 ;
      RECT 4.7070 10.7050 4.9050 13.3250 ;
      RECT 3.7670 13.0990 4.4370 13.3250 ;
      RECT 5.2250 9.0595 5.8450 12.6440 ;
      RECT 5.1750 10.1650 5.8450 11.9510 ;
      RECT 3.7670 11.1370 4.4370 11.5070 ;
      RECT 4.7210 10.4350 4.9050 10.6250 ;
      RECT 3.8210 10.3990 4.4370 10.5890 ;
      RECT 4.7070 10.2910 4.8910 10.4270 ;
      RECT 4.7210 10.1650 4.9050 10.3910 ;
      RECT 6.0890 10.1950 9.4090 17.5365 ;
      RECT 7.1690 10.1920 9.4090 17.5365 ;
      RECT 5.9270 8.8830 6.0070 17.5365 ;
      RECT 3.7670 9.5680 3.9550 10.3820 ;
      RECT 5.9270 8.8830 6.2230 10.2860 ;
      RECT 5.9270 10.0000 7.0870 10.2860 ;
      RECT 7.1690 8.8830 7.3030 17.5365 ;
      RECT 2.5250 9.8110 3.3070 17.5365 ;
      RECT 0.2030 8.8830 2.4430 17.5365 ;
      RECT 5.9270 10.0000 7.3030 10.0940 ;
      RECT 6.9530 8.8830 9.4090 10.0910 ;
      RECT 3.1730 8.8830 3.6850 10.0910 ;
      RECT 4.7070 10.0210 4.9050 10.0850 ;
      RECT 4.7070 9.8950 4.8910 10.0850 ;
      RECT 6.7370 9.6160 9.4090 10.0910 ;
      RECT 5.9270 9.6490 6.6550 10.2860 ;
      RECT 4.7210 9.6250 4.9050 9.8870 ;
      RECT 0.2030 9.6160 3.0910 10.0910 ;
      RECT 2.9570 8.8830 3.0910 17.5365 ;
      RECT 6.5210 8.8830 6.8710 9.7550 ;
      RECT 5.9270 9.5680 6.4390 10.2860 ;
      RECT 6.3050 8.8830 6.4390 17.5365 ;
      RECT 2.7410 9.5680 3.0910 17.5365 ;
      RECT 0.2030 8.8830 2.6590 10.0910 ;
      RECT 4.7210 8.8830 4.7470 17.5365 ;
      RECT 3.8570 8.8830 3.9550 17.5365 ;
      RECT 2.7410 8.8830 2.8750 17.5365 ;
      RECT 6.3050 8.8830 6.8710 9.5180 ;
      RECT 5.1890 8.8830 5.7910 9.5180 ;
      RECT 3.8570 8.8830 4.3870 9.5180 ;
      RECT 2.9570 8.8830 3.6850 9.5180 ;
      RECT 6.3050 8.8830 9.4090 9.5150 ;
      RECT 0.2030 8.8830 2.8750 9.5150 ;
      RECT 5.1750 9.3550 5.8450 9.5090 ;
      RECT 3.8570 9.3550 4.4010 9.5180 ;
      RECT 5.9270 8.8830 9.4090 9.2510 ;
      RECT 4.7210 8.8830 4.8910 9.2510 ;
      RECT 3.7670 8.8830 4.3870 9.2510 ;
      RECT 0.2030 8.8830 3.6850 9.2510 ;
      RECT 4.5410 8.8830 4.8910 9.1480 ;
      RECT 5.1800 8.8830 5.7910 9.0480 ;
      RECT 4.5410 8.8830 4.9270 9.0480 ;
      RECT 5.1800 8.8830 5.8450 8.9040 ;
      RECT 6.3090 8.8565 6.3270 17.5365 ;
      RECT 6.2010 8.8565 6.2190 17.5365 ;
      RECT 2.9610 8.8565 2.9790 17.5365 ;
      RECT 2.8530 8.8565 2.8710 17.5365 ;
      RECT 5.0180 8.8830 5.0800 9.0480 ;
        RECT 5.1800 17.0235 5.3080 18.1170 ;
        RECT 5.1660 17.6890 5.3080 18.0115 ;
        RECT 5.0180 17.4160 5.0800 18.1170 ;
        RECT 5.0040 17.7255 5.0800 17.8790 ;
        RECT 5.0180 17.0235 5.0440 18.1170 ;
        RECT 5.0180 17.1445 5.0580 17.3840 ;
        RECT 5.0180 17.0235 5.0800 17.1125 ;
        RECT 4.7210 17.4740 4.9270 18.1170 ;
        RECT 4.9010 17.0235 4.9270 18.1170 ;
        RECT 4.7210 17.7510 4.9410 18.0090 ;
        RECT 4.7210 17.0235 4.8190 18.1170 ;
        RECT 4.3040 17.0235 4.3870 18.1170 ;
        RECT 4.3040 17.1120 4.4010 18.0475 ;
        RECT 9.5270 17.0235 9.6120 18.1170 ;
        RECT 9.3830 17.0235 9.4090 18.1170 ;
        RECT 9.2750 17.0235 9.3010 18.1170 ;
        RECT 9.1670 17.0235 9.1930 18.1170 ;
        RECT 9.0590 17.0235 9.0850 18.1170 ;
        RECT 8.9510 17.0235 8.9770 18.1170 ;
        RECT 8.8430 17.0235 8.8690 18.1170 ;
        RECT 8.7350 17.0235 8.7610 18.1170 ;
        RECT 8.6270 17.0235 8.6530 18.1170 ;
        RECT 8.5190 17.0235 8.5450 18.1170 ;
        RECT 8.4110 17.0235 8.4370 18.1170 ;
        RECT 8.3030 17.0235 8.3290 18.1170 ;
        RECT 8.1950 17.0235 8.2210 18.1170 ;
        RECT 8.0870 17.0235 8.1130 18.1170 ;
        RECT 7.9790 17.0235 8.0050 18.1170 ;
        RECT 7.8710 17.0235 7.8970 18.1170 ;
        RECT 7.7630 17.0235 7.7890 18.1170 ;
        RECT 7.6550 17.0235 7.6810 18.1170 ;
        RECT 7.5470 17.0235 7.5730 18.1170 ;
        RECT 7.4390 17.0235 7.4650 18.1170 ;
        RECT 7.3310 17.0235 7.3570 18.1170 ;
        RECT 7.2230 17.0235 7.2490 18.1170 ;
        RECT 7.1150 17.0235 7.1410 18.1170 ;
        RECT 7.0070 17.0235 7.0330 18.1170 ;
        RECT 6.8990 17.0235 6.9250 18.1170 ;
        RECT 6.7910 17.0235 6.8170 18.1170 ;
        RECT 6.6830 17.0235 6.7090 18.1170 ;
        RECT 6.5750 17.0235 6.6010 18.1170 ;
        RECT 6.4670 17.0235 6.4930 18.1170 ;
        RECT 6.3590 17.0235 6.3850 18.1170 ;
        RECT 6.2510 17.0235 6.2770 18.1170 ;
        RECT 6.1430 17.0235 6.1690 18.1170 ;
        RECT 6.0350 17.0235 6.0610 18.1170 ;
        RECT 5.9270 17.0235 5.9530 18.1170 ;
        RECT 5.7140 17.0235 5.7910 18.1170 ;
        RECT 3.8210 17.0235 3.8980 18.1170 ;
        RECT 3.6590 17.0235 3.6850 18.1170 ;
        RECT 3.5510 17.0235 3.5770 18.1170 ;
        RECT 3.4430 17.0235 3.4690 18.1170 ;
        RECT 3.3350 17.0235 3.3610 18.1170 ;
        RECT 3.2270 17.0235 3.2530 18.1170 ;
        RECT 3.1190 17.0235 3.1450 18.1170 ;
        RECT 3.0110 17.0235 3.0370 18.1170 ;
        RECT 2.9030 17.0235 2.9290 18.1170 ;
        RECT 2.7950 17.0235 2.8210 18.1170 ;
        RECT 2.6870 17.0235 2.7130 18.1170 ;
        RECT 2.5790 17.0235 2.6050 18.1170 ;
        RECT 2.4710 17.0235 2.4970 18.1170 ;
        RECT 2.3630 17.0235 2.3890 18.1170 ;
        RECT 2.2550 17.0235 2.2810 18.1170 ;
        RECT 2.1470 17.0235 2.1730 18.1170 ;
        RECT 2.0390 17.0235 2.0650 18.1170 ;
        RECT 1.9310 17.0235 1.9570 18.1170 ;
        RECT 1.8230 17.0235 1.8490 18.1170 ;
        RECT 1.7150 17.0235 1.7410 18.1170 ;
        RECT 1.6070 17.0235 1.6330 18.1170 ;
        RECT 1.4990 17.0235 1.5250 18.1170 ;
        RECT 1.3910 17.0235 1.4170 18.1170 ;
        RECT 1.2830 17.0235 1.3090 18.1170 ;
        RECT 1.1750 17.0235 1.2010 18.1170 ;
        RECT 1.0670 17.0235 1.0930 18.1170 ;
        RECT 0.9590 17.0235 0.9850 18.1170 ;
        RECT 0.8510 17.0235 0.8770 18.1170 ;
        RECT 0.7430 17.0235 0.7690 18.1170 ;
        RECT 0.6350 17.0235 0.6610 18.1170 ;
        RECT 0.5270 17.0235 0.5530 18.1170 ;
        RECT 0.4190 17.0235 0.4450 18.1170 ;
        RECT 0.3110 17.0235 0.3370 18.1170 ;
        RECT 0.2030 17.0235 0.2290 18.1170 ;
        RECT 0.0000 17.0235 0.0850 18.1170 ;
        RECT 5.1800 18.1035 5.3080 19.1970 ;
        RECT 5.1660 18.7690 5.3080 19.0915 ;
        RECT 5.0180 18.4960 5.0800 19.1970 ;
        RECT 5.0040 18.8055 5.0800 18.9590 ;
        RECT 5.0180 18.1035 5.0440 19.1970 ;
        RECT 5.0180 18.2245 5.0580 18.4640 ;
        RECT 5.0180 18.1035 5.0800 18.1925 ;
        RECT 4.7210 18.5540 4.9270 19.1970 ;
        RECT 4.9010 18.1035 4.9270 19.1970 ;
        RECT 4.7210 18.8310 4.9410 19.0890 ;
        RECT 4.7210 18.1035 4.8190 19.1970 ;
        RECT 4.3040 18.1035 4.3870 19.1970 ;
        RECT 4.3040 18.1920 4.4010 19.1275 ;
        RECT 9.5270 18.1035 9.6120 19.1970 ;
        RECT 9.3830 18.1035 9.4090 19.1970 ;
        RECT 9.2750 18.1035 9.3010 19.1970 ;
        RECT 9.1670 18.1035 9.1930 19.1970 ;
        RECT 9.0590 18.1035 9.0850 19.1970 ;
        RECT 8.9510 18.1035 8.9770 19.1970 ;
        RECT 8.8430 18.1035 8.8690 19.1970 ;
        RECT 8.7350 18.1035 8.7610 19.1970 ;
        RECT 8.6270 18.1035 8.6530 19.1970 ;
        RECT 8.5190 18.1035 8.5450 19.1970 ;
        RECT 8.4110 18.1035 8.4370 19.1970 ;
        RECT 8.3030 18.1035 8.3290 19.1970 ;
        RECT 8.1950 18.1035 8.2210 19.1970 ;
        RECT 8.0870 18.1035 8.1130 19.1970 ;
        RECT 7.9790 18.1035 8.0050 19.1970 ;
        RECT 7.8710 18.1035 7.8970 19.1970 ;
        RECT 7.7630 18.1035 7.7890 19.1970 ;
        RECT 7.6550 18.1035 7.6810 19.1970 ;
        RECT 7.5470 18.1035 7.5730 19.1970 ;
        RECT 7.4390 18.1035 7.4650 19.1970 ;
        RECT 7.3310 18.1035 7.3570 19.1970 ;
        RECT 7.2230 18.1035 7.2490 19.1970 ;
        RECT 7.1150 18.1035 7.1410 19.1970 ;
        RECT 7.0070 18.1035 7.0330 19.1970 ;
        RECT 6.8990 18.1035 6.9250 19.1970 ;
        RECT 6.7910 18.1035 6.8170 19.1970 ;
        RECT 6.6830 18.1035 6.7090 19.1970 ;
        RECT 6.5750 18.1035 6.6010 19.1970 ;
        RECT 6.4670 18.1035 6.4930 19.1970 ;
        RECT 6.3590 18.1035 6.3850 19.1970 ;
        RECT 6.2510 18.1035 6.2770 19.1970 ;
        RECT 6.1430 18.1035 6.1690 19.1970 ;
        RECT 6.0350 18.1035 6.0610 19.1970 ;
        RECT 5.9270 18.1035 5.9530 19.1970 ;
        RECT 5.7140 18.1035 5.7910 19.1970 ;
        RECT 3.8210 18.1035 3.8980 19.1970 ;
        RECT 3.6590 18.1035 3.6850 19.1970 ;
        RECT 3.5510 18.1035 3.5770 19.1970 ;
        RECT 3.4430 18.1035 3.4690 19.1970 ;
        RECT 3.3350 18.1035 3.3610 19.1970 ;
        RECT 3.2270 18.1035 3.2530 19.1970 ;
        RECT 3.1190 18.1035 3.1450 19.1970 ;
        RECT 3.0110 18.1035 3.0370 19.1970 ;
        RECT 2.9030 18.1035 2.9290 19.1970 ;
        RECT 2.7950 18.1035 2.8210 19.1970 ;
        RECT 2.6870 18.1035 2.7130 19.1970 ;
        RECT 2.5790 18.1035 2.6050 19.1970 ;
        RECT 2.4710 18.1035 2.4970 19.1970 ;
        RECT 2.3630 18.1035 2.3890 19.1970 ;
        RECT 2.2550 18.1035 2.2810 19.1970 ;
        RECT 2.1470 18.1035 2.1730 19.1970 ;
        RECT 2.0390 18.1035 2.0650 19.1970 ;
        RECT 1.9310 18.1035 1.9570 19.1970 ;
        RECT 1.8230 18.1035 1.8490 19.1970 ;
        RECT 1.7150 18.1035 1.7410 19.1970 ;
        RECT 1.6070 18.1035 1.6330 19.1970 ;
        RECT 1.4990 18.1035 1.5250 19.1970 ;
        RECT 1.3910 18.1035 1.4170 19.1970 ;
        RECT 1.2830 18.1035 1.3090 19.1970 ;
        RECT 1.1750 18.1035 1.2010 19.1970 ;
        RECT 1.0670 18.1035 1.0930 19.1970 ;
        RECT 0.9590 18.1035 0.9850 19.1970 ;
        RECT 0.8510 18.1035 0.8770 19.1970 ;
        RECT 0.7430 18.1035 0.7690 19.1970 ;
        RECT 0.6350 18.1035 0.6610 19.1970 ;
        RECT 0.5270 18.1035 0.5530 19.1970 ;
        RECT 0.4190 18.1035 0.4450 19.1970 ;
        RECT 0.3110 18.1035 0.3370 19.1970 ;
        RECT 0.2030 18.1035 0.2290 19.1970 ;
        RECT 0.0000 18.1035 0.0850 19.1970 ;
        RECT 5.1800 19.1835 5.3080 20.2770 ;
        RECT 5.1660 19.8490 5.3080 20.1715 ;
        RECT 5.0180 19.5760 5.0800 20.2770 ;
        RECT 5.0040 19.8855 5.0800 20.0390 ;
        RECT 5.0180 19.1835 5.0440 20.2770 ;
        RECT 5.0180 19.3045 5.0580 19.5440 ;
        RECT 5.0180 19.1835 5.0800 19.2725 ;
        RECT 4.7210 19.6340 4.9270 20.2770 ;
        RECT 4.9010 19.1835 4.9270 20.2770 ;
        RECT 4.7210 19.9110 4.9410 20.1690 ;
        RECT 4.7210 19.1835 4.8190 20.2770 ;
        RECT 4.3040 19.1835 4.3870 20.2770 ;
        RECT 4.3040 19.2720 4.4010 20.2075 ;
        RECT 9.5270 19.1835 9.6120 20.2770 ;
        RECT 9.3830 19.1835 9.4090 20.2770 ;
        RECT 9.2750 19.1835 9.3010 20.2770 ;
        RECT 9.1670 19.1835 9.1930 20.2770 ;
        RECT 9.0590 19.1835 9.0850 20.2770 ;
        RECT 8.9510 19.1835 8.9770 20.2770 ;
        RECT 8.8430 19.1835 8.8690 20.2770 ;
        RECT 8.7350 19.1835 8.7610 20.2770 ;
        RECT 8.6270 19.1835 8.6530 20.2770 ;
        RECT 8.5190 19.1835 8.5450 20.2770 ;
        RECT 8.4110 19.1835 8.4370 20.2770 ;
        RECT 8.3030 19.1835 8.3290 20.2770 ;
        RECT 8.1950 19.1835 8.2210 20.2770 ;
        RECT 8.0870 19.1835 8.1130 20.2770 ;
        RECT 7.9790 19.1835 8.0050 20.2770 ;
        RECT 7.8710 19.1835 7.8970 20.2770 ;
        RECT 7.7630 19.1835 7.7890 20.2770 ;
        RECT 7.6550 19.1835 7.6810 20.2770 ;
        RECT 7.5470 19.1835 7.5730 20.2770 ;
        RECT 7.4390 19.1835 7.4650 20.2770 ;
        RECT 7.3310 19.1835 7.3570 20.2770 ;
        RECT 7.2230 19.1835 7.2490 20.2770 ;
        RECT 7.1150 19.1835 7.1410 20.2770 ;
        RECT 7.0070 19.1835 7.0330 20.2770 ;
        RECT 6.8990 19.1835 6.9250 20.2770 ;
        RECT 6.7910 19.1835 6.8170 20.2770 ;
        RECT 6.6830 19.1835 6.7090 20.2770 ;
        RECT 6.5750 19.1835 6.6010 20.2770 ;
        RECT 6.4670 19.1835 6.4930 20.2770 ;
        RECT 6.3590 19.1835 6.3850 20.2770 ;
        RECT 6.2510 19.1835 6.2770 20.2770 ;
        RECT 6.1430 19.1835 6.1690 20.2770 ;
        RECT 6.0350 19.1835 6.0610 20.2770 ;
        RECT 5.9270 19.1835 5.9530 20.2770 ;
        RECT 5.7140 19.1835 5.7910 20.2770 ;
        RECT 3.8210 19.1835 3.8980 20.2770 ;
        RECT 3.6590 19.1835 3.6850 20.2770 ;
        RECT 3.5510 19.1835 3.5770 20.2770 ;
        RECT 3.4430 19.1835 3.4690 20.2770 ;
        RECT 3.3350 19.1835 3.3610 20.2770 ;
        RECT 3.2270 19.1835 3.2530 20.2770 ;
        RECT 3.1190 19.1835 3.1450 20.2770 ;
        RECT 3.0110 19.1835 3.0370 20.2770 ;
        RECT 2.9030 19.1835 2.9290 20.2770 ;
        RECT 2.7950 19.1835 2.8210 20.2770 ;
        RECT 2.6870 19.1835 2.7130 20.2770 ;
        RECT 2.5790 19.1835 2.6050 20.2770 ;
        RECT 2.4710 19.1835 2.4970 20.2770 ;
        RECT 2.3630 19.1835 2.3890 20.2770 ;
        RECT 2.2550 19.1835 2.2810 20.2770 ;
        RECT 2.1470 19.1835 2.1730 20.2770 ;
        RECT 2.0390 19.1835 2.0650 20.2770 ;
        RECT 1.9310 19.1835 1.9570 20.2770 ;
        RECT 1.8230 19.1835 1.8490 20.2770 ;
        RECT 1.7150 19.1835 1.7410 20.2770 ;
        RECT 1.6070 19.1835 1.6330 20.2770 ;
        RECT 1.4990 19.1835 1.5250 20.2770 ;
        RECT 1.3910 19.1835 1.4170 20.2770 ;
        RECT 1.2830 19.1835 1.3090 20.2770 ;
        RECT 1.1750 19.1835 1.2010 20.2770 ;
        RECT 1.0670 19.1835 1.0930 20.2770 ;
        RECT 0.9590 19.1835 0.9850 20.2770 ;
        RECT 0.8510 19.1835 0.8770 20.2770 ;
        RECT 0.7430 19.1835 0.7690 20.2770 ;
        RECT 0.6350 19.1835 0.6610 20.2770 ;
        RECT 0.5270 19.1835 0.5530 20.2770 ;
        RECT 0.4190 19.1835 0.4450 20.2770 ;
        RECT 0.3110 19.1835 0.3370 20.2770 ;
        RECT 0.2030 19.1835 0.2290 20.2770 ;
        RECT 0.0000 19.1835 0.0850 20.2770 ;
        RECT 5.1800 20.2635 5.3080 21.3570 ;
        RECT 5.1660 20.9290 5.3080 21.2515 ;
        RECT 5.0180 20.6560 5.0800 21.3570 ;
        RECT 5.0040 20.9655 5.0800 21.1190 ;
        RECT 5.0180 20.2635 5.0440 21.3570 ;
        RECT 5.0180 20.3845 5.0580 20.6240 ;
        RECT 5.0180 20.2635 5.0800 20.3525 ;
        RECT 4.7210 20.7140 4.9270 21.3570 ;
        RECT 4.9010 20.2635 4.9270 21.3570 ;
        RECT 4.7210 20.9910 4.9410 21.2490 ;
        RECT 4.7210 20.2635 4.8190 21.3570 ;
        RECT 4.3040 20.2635 4.3870 21.3570 ;
        RECT 4.3040 20.3520 4.4010 21.2875 ;
        RECT 9.5270 20.2635 9.6120 21.3570 ;
        RECT 9.3830 20.2635 9.4090 21.3570 ;
        RECT 9.2750 20.2635 9.3010 21.3570 ;
        RECT 9.1670 20.2635 9.1930 21.3570 ;
        RECT 9.0590 20.2635 9.0850 21.3570 ;
        RECT 8.9510 20.2635 8.9770 21.3570 ;
        RECT 8.8430 20.2635 8.8690 21.3570 ;
        RECT 8.7350 20.2635 8.7610 21.3570 ;
        RECT 8.6270 20.2635 8.6530 21.3570 ;
        RECT 8.5190 20.2635 8.5450 21.3570 ;
        RECT 8.4110 20.2635 8.4370 21.3570 ;
        RECT 8.3030 20.2635 8.3290 21.3570 ;
        RECT 8.1950 20.2635 8.2210 21.3570 ;
        RECT 8.0870 20.2635 8.1130 21.3570 ;
        RECT 7.9790 20.2635 8.0050 21.3570 ;
        RECT 7.8710 20.2635 7.8970 21.3570 ;
        RECT 7.7630 20.2635 7.7890 21.3570 ;
        RECT 7.6550 20.2635 7.6810 21.3570 ;
        RECT 7.5470 20.2635 7.5730 21.3570 ;
        RECT 7.4390 20.2635 7.4650 21.3570 ;
        RECT 7.3310 20.2635 7.3570 21.3570 ;
        RECT 7.2230 20.2635 7.2490 21.3570 ;
        RECT 7.1150 20.2635 7.1410 21.3570 ;
        RECT 7.0070 20.2635 7.0330 21.3570 ;
        RECT 6.8990 20.2635 6.9250 21.3570 ;
        RECT 6.7910 20.2635 6.8170 21.3570 ;
        RECT 6.6830 20.2635 6.7090 21.3570 ;
        RECT 6.5750 20.2635 6.6010 21.3570 ;
        RECT 6.4670 20.2635 6.4930 21.3570 ;
        RECT 6.3590 20.2635 6.3850 21.3570 ;
        RECT 6.2510 20.2635 6.2770 21.3570 ;
        RECT 6.1430 20.2635 6.1690 21.3570 ;
        RECT 6.0350 20.2635 6.0610 21.3570 ;
        RECT 5.9270 20.2635 5.9530 21.3570 ;
        RECT 5.7140 20.2635 5.7910 21.3570 ;
        RECT 3.8210 20.2635 3.8980 21.3570 ;
        RECT 3.6590 20.2635 3.6850 21.3570 ;
        RECT 3.5510 20.2635 3.5770 21.3570 ;
        RECT 3.4430 20.2635 3.4690 21.3570 ;
        RECT 3.3350 20.2635 3.3610 21.3570 ;
        RECT 3.2270 20.2635 3.2530 21.3570 ;
        RECT 3.1190 20.2635 3.1450 21.3570 ;
        RECT 3.0110 20.2635 3.0370 21.3570 ;
        RECT 2.9030 20.2635 2.9290 21.3570 ;
        RECT 2.7950 20.2635 2.8210 21.3570 ;
        RECT 2.6870 20.2635 2.7130 21.3570 ;
        RECT 2.5790 20.2635 2.6050 21.3570 ;
        RECT 2.4710 20.2635 2.4970 21.3570 ;
        RECT 2.3630 20.2635 2.3890 21.3570 ;
        RECT 2.2550 20.2635 2.2810 21.3570 ;
        RECT 2.1470 20.2635 2.1730 21.3570 ;
        RECT 2.0390 20.2635 2.0650 21.3570 ;
        RECT 1.9310 20.2635 1.9570 21.3570 ;
        RECT 1.8230 20.2635 1.8490 21.3570 ;
        RECT 1.7150 20.2635 1.7410 21.3570 ;
        RECT 1.6070 20.2635 1.6330 21.3570 ;
        RECT 1.4990 20.2635 1.5250 21.3570 ;
        RECT 1.3910 20.2635 1.4170 21.3570 ;
        RECT 1.2830 20.2635 1.3090 21.3570 ;
        RECT 1.1750 20.2635 1.2010 21.3570 ;
        RECT 1.0670 20.2635 1.0930 21.3570 ;
        RECT 0.9590 20.2635 0.9850 21.3570 ;
        RECT 0.8510 20.2635 0.8770 21.3570 ;
        RECT 0.7430 20.2635 0.7690 21.3570 ;
        RECT 0.6350 20.2635 0.6610 21.3570 ;
        RECT 0.5270 20.2635 0.5530 21.3570 ;
        RECT 0.4190 20.2635 0.4450 21.3570 ;
        RECT 0.3110 20.2635 0.3370 21.3570 ;
        RECT 0.2030 20.2635 0.2290 21.3570 ;
        RECT 0.0000 20.2635 0.0850 21.3570 ;
        RECT 5.1800 21.3435 5.3080 22.4370 ;
        RECT 5.1660 22.0090 5.3080 22.3315 ;
        RECT 5.0180 21.7360 5.0800 22.4370 ;
        RECT 5.0040 22.0455 5.0800 22.1990 ;
        RECT 5.0180 21.3435 5.0440 22.4370 ;
        RECT 5.0180 21.4645 5.0580 21.7040 ;
        RECT 5.0180 21.3435 5.0800 21.4325 ;
        RECT 4.7210 21.7940 4.9270 22.4370 ;
        RECT 4.9010 21.3435 4.9270 22.4370 ;
        RECT 4.7210 22.0710 4.9410 22.3290 ;
        RECT 4.7210 21.3435 4.8190 22.4370 ;
        RECT 4.3040 21.3435 4.3870 22.4370 ;
        RECT 4.3040 21.4320 4.4010 22.3675 ;
        RECT 9.5270 21.3435 9.6120 22.4370 ;
        RECT 9.3830 21.3435 9.4090 22.4370 ;
        RECT 9.2750 21.3435 9.3010 22.4370 ;
        RECT 9.1670 21.3435 9.1930 22.4370 ;
        RECT 9.0590 21.3435 9.0850 22.4370 ;
        RECT 8.9510 21.3435 8.9770 22.4370 ;
        RECT 8.8430 21.3435 8.8690 22.4370 ;
        RECT 8.7350 21.3435 8.7610 22.4370 ;
        RECT 8.6270 21.3435 8.6530 22.4370 ;
        RECT 8.5190 21.3435 8.5450 22.4370 ;
        RECT 8.4110 21.3435 8.4370 22.4370 ;
        RECT 8.3030 21.3435 8.3290 22.4370 ;
        RECT 8.1950 21.3435 8.2210 22.4370 ;
        RECT 8.0870 21.3435 8.1130 22.4370 ;
        RECT 7.9790 21.3435 8.0050 22.4370 ;
        RECT 7.8710 21.3435 7.8970 22.4370 ;
        RECT 7.7630 21.3435 7.7890 22.4370 ;
        RECT 7.6550 21.3435 7.6810 22.4370 ;
        RECT 7.5470 21.3435 7.5730 22.4370 ;
        RECT 7.4390 21.3435 7.4650 22.4370 ;
        RECT 7.3310 21.3435 7.3570 22.4370 ;
        RECT 7.2230 21.3435 7.2490 22.4370 ;
        RECT 7.1150 21.3435 7.1410 22.4370 ;
        RECT 7.0070 21.3435 7.0330 22.4370 ;
        RECT 6.8990 21.3435 6.9250 22.4370 ;
        RECT 6.7910 21.3435 6.8170 22.4370 ;
        RECT 6.6830 21.3435 6.7090 22.4370 ;
        RECT 6.5750 21.3435 6.6010 22.4370 ;
        RECT 6.4670 21.3435 6.4930 22.4370 ;
        RECT 6.3590 21.3435 6.3850 22.4370 ;
        RECT 6.2510 21.3435 6.2770 22.4370 ;
        RECT 6.1430 21.3435 6.1690 22.4370 ;
        RECT 6.0350 21.3435 6.0610 22.4370 ;
        RECT 5.9270 21.3435 5.9530 22.4370 ;
        RECT 5.7140 21.3435 5.7910 22.4370 ;
        RECT 3.8210 21.3435 3.8980 22.4370 ;
        RECT 3.6590 21.3435 3.6850 22.4370 ;
        RECT 3.5510 21.3435 3.5770 22.4370 ;
        RECT 3.4430 21.3435 3.4690 22.4370 ;
        RECT 3.3350 21.3435 3.3610 22.4370 ;
        RECT 3.2270 21.3435 3.2530 22.4370 ;
        RECT 3.1190 21.3435 3.1450 22.4370 ;
        RECT 3.0110 21.3435 3.0370 22.4370 ;
        RECT 2.9030 21.3435 2.9290 22.4370 ;
        RECT 2.7950 21.3435 2.8210 22.4370 ;
        RECT 2.6870 21.3435 2.7130 22.4370 ;
        RECT 2.5790 21.3435 2.6050 22.4370 ;
        RECT 2.4710 21.3435 2.4970 22.4370 ;
        RECT 2.3630 21.3435 2.3890 22.4370 ;
        RECT 2.2550 21.3435 2.2810 22.4370 ;
        RECT 2.1470 21.3435 2.1730 22.4370 ;
        RECT 2.0390 21.3435 2.0650 22.4370 ;
        RECT 1.9310 21.3435 1.9570 22.4370 ;
        RECT 1.8230 21.3435 1.8490 22.4370 ;
        RECT 1.7150 21.3435 1.7410 22.4370 ;
        RECT 1.6070 21.3435 1.6330 22.4370 ;
        RECT 1.4990 21.3435 1.5250 22.4370 ;
        RECT 1.3910 21.3435 1.4170 22.4370 ;
        RECT 1.2830 21.3435 1.3090 22.4370 ;
        RECT 1.1750 21.3435 1.2010 22.4370 ;
        RECT 1.0670 21.3435 1.0930 22.4370 ;
        RECT 0.9590 21.3435 0.9850 22.4370 ;
        RECT 0.8510 21.3435 0.8770 22.4370 ;
        RECT 0.7430 21.3435 0.7690 22.4370 ;
        RECT 0.6350 21.3435 0.6610 22.4370 ;
        RECT 0.5270 21.3435 0.5530 22.4370 ;
        RECT 0.4190 21.3435 0.4450 22.4370 ;
        RECT 0.3110 21.3435 0.3370 22.4370 ;
        RECT 0.2030 21.3435 0.2290 22.4370 ;
        RECT 0.0000 21.3435 0.0850 22.4370 ;
        RECT 5.1800 22.4235 5.3080 23.5170 ;
        RECT 5.1660 23.0890 5.3080 23.4115 ;
        RECT 5.0180 22.8160 5.0800 23.5170 ;
        RECT 5.0040 23.1255 5.0800 23.2790 ;
        RECT 5.0180 22.4235 5.0440 23.5170 ;
        RECT 5.0180 22.5445 5.0580 22.7840 ;
        RECT 5.0180 22.4235 5.0800 22.5125 ;
        RECT 4.7210 22.8740 4.9270 23.5170 ;
        RECT 4.9010 22.4235 4.9270 23.5170 ;
        RECT 4.7210 23.1510 4.9410 23.4090 ;
        RECT 4.7210 22.4235 4.8190 23.5170 ;
        RECT 4.3040 22.4235 4.3870 23.5170 ;
        RECT 4.3040 22.5120 4.4010 23.4475 ;
        RECT 9.5270 22.4235 9.6120 23.5170 ;
        RECT 9.3830 22.4235 9.4090 23.5170 ;
        RECT 9.2750 22.4235 9.3010 23.5170 ;
        RECT 9.1670 22.4235 9.1930 23.5170 ;
        RECT 9.0590 22.4235 9.0850 23.5170 ;
        RECT 8.9510 22.4235 8.9770 23.5170 ;
        RECT 8.8430 22.4235 8.8690 23.5170 ;
        RECT 8.7350 22.4235 8.7610 23.5170 ;
        RECT 8.6270 22.4235 8.6530 23.5170 ;
        RECT 8.5190 22.4235 8.5450 23.5170 ;
        RECT 8.4110 22.4235 8.4370 23.5170 ;
        RECT 8.3030 22.4235 8.3290 23.5170 ;
        RECT 8.1950 22.4235 8.2210 23.5170 ;
        RECT 8.0870 22.4235 8.1130 23.5170 ;
        RECT 7.9790 22.4235 8.0050 23.5170 ;
        RECT 7.8710 22.4235 7.8970 23.5170 ;
        RECT 7.7630 22.4235 7.7890 23.5170 ;
        RECT 7.6550 22.4235 7.6810 23.5170 ;
        RECT 7.5470 22.4235 7.5730 23.5170 ;
        RECT 7.4390 22.4235 7.4650 23.5170 ;
        RECT 7.3310 22.4235 7.3570 23.5170 ;
        RECT 7.2230 22.4235 7.2490 23.5170 ;
        RECT 7.1150 22.4235 7.1410 23.5170 ;
        RECT 7.0070 22.4235 7.0330 23.5170 ;
        RECT 6.8990 22.4235 6.9250 23.5170 ;
        RECT 6.7910 22.4235 6.8170 23.5170 ;
        RECT 6.6830 22.4235 6.7090 23.5170 ;
        RECT 6.5750 22.4235 6.6010 23.5170 ;
        RECT 6.4670 22.4235 6.4930 23.5170 ;
        RECT 6.3590 22.4235 6.3850 23.5170 ;
        RECT 6.2510 22.4235 6.2770 23.5170 ;
        RECT 6.1430 22.4235 6.1690 23.5170 ;
        RECT 6.0350 22.4235 6.0610 23.5170 ;
        RECT 5.9270 22.4235 5.9530 23.5170 ;
        RECT 5.7140 22.4235 5.7910 23.5170 ;
        RECT 3.8210 22.4235 3.8980 23.5170 ;
        RECT 3.6590 22.4235 3.6850 23.5170 ;
        RECT 3.5510 22.4235 3.5770 23.5170 ;
        RECT 3.4430 22.4235 3.4690 23.5170 ;
        RECT 3.3350 22.4235 3.3610 23.5170 ;
        RECT 3.2270 22.4235 3.2530 23.5170 ;
        RECT 3.1190 22.4235 3.1450 23.5170 ;
        RECT 3.0110 22.4235 3.0370 23.5170 ;
        RECT 2.9030 22.4235 2.9290 23.5170 ;
        RECT 2.7950 22.4235 2.8210 23.5170 ;
        RECT 2.6870 22.4235 2.7130 23.5170 ;
        RECT 2.5790 22.4235 2.6050 23.5170 ;
        RECT 2.4710 22.4235 2.4970 23.5170 ;
        RECT 2.3630 22.4235 2.3890 23.5170 ;
        RECT 2.2550 22.4235 2.2810 23.5170 ;
        RECT 2.1470 22.4235 2.1730 23.5170 ;
        RECT 2.0390 22.4235 2.0650 23.5170 ;
        RECT 1.9310 22.4235 1.9570 23.5170 ;
        RECT 1.8230 22.4235 1.8490 23.5170 ;
        RECT 1.7150 22.4235 1.7410 23.5170 ;
        RECT 1.6070 22.4235 1.6330 23.5170 ;
        RECT 1.4990 22.4235 1.5250 23.5170 ;
        RECT 1.3910 22.4235 1.4170 23.5170 ;
        RECT 1.2830 22.4235 1.3090 23.5170 ;
        RECT 1.1750 22.4235 1.2010 23.5170 ;
        RECT 1.0670 22.4235 1.0930 23.5170 ;
        RECT 0.9590 22.4235 0.9850 23.5170 ;
        RECT 0.8510 22.4235 0.8770 23.5170 ;
        RECT 0.7430 22.4235 0.7690 23.5170 ;
        RECT 0.6350 22.4235 0.6610 23.5170 ;
        RECT 0.5270 22.4235 0.5530 23.5170 ;
        RECT 0.4190 22.4235 0.4450 23.5170 ;
        RECT 0.3110 22.4235 0.3370 23.5170 ;
        RECT 0.2030 22.4235 0.2290 23.5170 ;
        RECT 0.0000 22.4235 0.0850 23.5170 ;
        RECT 5.1800 23.5035 5.3080 24.5970 ;
        RECT 5.1660 24.1690 5.3080 24.4915 ;
        RECT 5.0180 23.8960 5.0800 24.5970 ;
        RECT 5.0040 24.2055 5.0800 24.3590 ;
        RECT 5.0180 23.5035 5.0440 24.5970 ;
        RECT 5.0180 23.6245 5.0580 23.8640 ;
        RECT 5.0180 23.5035 5.0800 23.5925 ;
        RECT 4.7210 23.9540 4.9270 24.5970 ;
        RECT 4.9010 23.5035 4.9270 24.5970 ;
        RECT 4.7210 24.2310 4.9410 24.4890 ;
        RECT 4.7210 23.5035 4.8190 24.5970 ;
        RECT 4.3040 23.5035 4.3870 24.5970 ;
        RECT 4.3040 23.5920 4.4010 24.5275 ;
        RECT 9.5270 23.5035 9.6120 24.5970 ;
        RECT 9.3830 23.5035 9.4090 24.5970 ;
        RECT 9.2750 23.5035 9.3010 24.5970 ;
        RECT 9.1670 23.5035 9.1930 24.5970 ;
        RECT 9.0590 23.5035 9.0850 24.5970 ;
        RECT 8.9510 23.5035 8.9770 24.5970 ;
        RECT 8.8430 23.5035 8.8690 24.5970 ;
        RECT 8.7350 23.5035 8.7610 24.5970 ;
        RECT 8.6270 23.5035 8.6530 24.5970 ;
        RECT 8.5190 23.5035 8.5450 24.5970 ;
        RECT 8.4110 23.5035 8.4370 24.5970 ;
        RECT 8.3030 23.5035 8.3290 24.5970 ;
        RECT 8.1950 23.5035 8.2210 24.5970 ;
        RECT 8.0870 23.5035 8.1130 24.5970 ;
        RECT 7.9790 23.5035 8.0050 24.5970 ;
        RECT 7.8710 23.5035 7.8970 24.5970 ;
        RECT 7.7630 23.5035 7.7890 24.5970 ;
        RECT 7.6550 23.5035 7.6810 24.5970 ;
        RECT 7.5470 23.5035 7.5730 24.5970 ;
        RECT 7.4390 23.5035 7.4650 24.5970 ;
        RECT 7.3310 23.5035 7.3570 24.5970 ;
        RECT 7.2230 23.5035 7.2490 24.5970 ;
        RECT 7.1150 23.5035 7.1410 24.5970 ;
        RECT 7.0070 23.5035 7.0330 24.5970 ;
        RECT 6.8990 23.5035 6.9250 24.5970 ;
        RECT 6.7910 23.5035 6.8170 24.5970 ;
        RECT 6.6830 23.5035 6.7090 24.5970 ;
        RECT 6.5750 23.5035 6.6010 24.5970 ;
        RECT 6.4670 23.5035 6.4930 24.5970 ;
        RECT 6.3590 23.5035 6.3850 24.5970 ;
        RECT 6.2510 23.5035 6.2770 24.5970 ;
        RECT 6.1430 23.5035 6.1690 24.5970 ;
        RECT 6.0350 23.5035 6.0610 24.5970 ;
        RECT 5.9270 23.5035 5.9530 24.5970 ;
        RECT 5.7140 23.5035 5.7910 24.5970 ;
        RECT 3.8210 23.5035 3.8980 24.5970 ;
        RECT 3.6590 23.5035 3.6850 24.5970 ;
        RECT 3.5510 23.5035 3.5770 24.5970 ;
        RECT 3.4430 23.5035 3.4690 24.5970 ;
        RECT 3.3350 23.5035 3.3610 24.5970 ;
        RECT 3.2270 23.5035 3.2530 24.5970 ;
        RECT 3.1190 23.5035 3.1450 24.5970 ;
        RECT 3.0110 23.5035 3.0370 24.5970 ;
        RECT 2.9030 23.5035 2.9290 24.5970 ;
        RECT 2.7950 23.5035 2.8210 24.5970 ;
        RECT 2.6870 23.5035 2.7130 24.5970 ;
        RECT 2.5790 23.5035 2.6050 24.5970 ;
        RECT 2.4710 23.5035 2.4970 24.5970 ;
        RECT 2.3630 23.5035 2.3890 24.5970 ;
        RECT 2.2550 23.5035 2.2810 24.5970 ;
        RECT 2.1470 23.5035 2.1730 24.5970 ;
        RECT 2.0390 23.5035 2.0650 24.5970 ;
        RECT 1.9310 23.5035 1.9570 24.5970 ;
        RECT 1.8230 23.5035 1.8490 24.5970 ;
        RECT 1.7150 23.5035 1.7410 24.5970 ;
        RECT 1.6070 23.5035 1.6330 24.5970 ;
        RECT 1.4990 23.5035 1.5250 24.5970 ;
        RECT 1.3910 23.5035 1.4170 24.5970 ;
        RECT 1.2830 23.5035 1.3090 24.5970 ;
        RECT 1.1750 23.5035 1.2010 24.5970 ;
        RECT 1.0670 23.5035 1.0930 24.5970 ;
        RECT 0.9590 23.5035 0.9850 24.5970 ;
        RECT 0.8510 23.5035 0.8770 24.5970 ;
        RECT 0.7430 23.5035 0.7690 24.5970 ;
        RECT 0.6350 23.5035 0.6610 24.5970 ;
        RECT 0.5270 23.5035 0.5530 24.5970 ;
        RECT 0.4190 23.5035 0.4450 24.5970 ;
        RECT 0.3110 23.5035 0.3370 24.5970 ;
        RECT 0.2030 23.5035 0.2290 24.5970 ;
        RECT 0.0000 23.5035 0.0850 24.5970 ;
        RECT 5.1800 24.5835 5.3080 25.6770 ;
        RECT 5.1660 25.2490 5.3080 25.5715 ;
        RECT 5.0180 24.9760 5.0800 25.6770 ;
        RECT 5.0040 25.2855 5.0800 25.4390 ;
        RECT 5.0180 24.5835 5.0440 25.6770 ;
        RECT 5.0180 24.7045 5.0580 24.9440 ;
        RECT 5.0180 24.5835 5.0800 24.6725 ;
        RECT 4.7210 25.0340 4.9270 25.6770 ;
        RECT 4.9010 24.5835 4.9270 25.6770 ;
        RECT 4.7210 25.3110 4.9410 25.5690 ;
        RECT 4.7210 24.5835 4.8190 25.6770 ;
        RECT 4.3040 24.5835 4.3870 25.6770 ;
        RECT 4.3040 24.6720 4.4010 25.6075 ;
        RECT 9.5270 24.5835 9.6120 25.6770 ;
        RECT 9.3830 24.5835 9.4090 25.6770 ;
        RECT 9.2750 24.5835 9.3010 25.6770 ;
        RECT 9.1670 24.5835 9.1930 25.6770 ;
        RECT 9.0590 24.5835 9.0850 25.6770 ;
        RECT 8.9510 24.5835 8.9770 25.6770 ;
        RECT 8.8430 24.5835 8.8690 25.6770 ;
        RECT 8.7350 24.5835 8.7610 25.6770 ;
        RECT 8.6270 24.5835 8.6530 25.6770 ;
        RECT 8.5190 24.5835 8.5450 25.6770 ;
        RECT 8.4110 24.5835 8.4370 25.6770 ;
        RECT 8.3030 24.5835 8.3290 25.6770 ;
        RECT 8.1950 24.5835 8.2210 25.6770 ;
        RECT 8.0870 24.5835 8.1130 25.6770 ;
        RECT 7.9790 24.5835 8.0050 25.6770 ;
        RECT 7.8710 24.5835 7.8970 25.6770 ;
        RECT 7.7630 24.5835 7.7890 25.6770 ;
        RECT 7.6550 24.5835 7.6810 25.6770 ;
        RECT 7.5470 24.5835 7.5730 25.6770 ;
        RECT 7.4390 24.5835 7.4650 25.6770 ;
        RECT 7.3310 24.5835 7.3570 25.6770 ;
        RECT 7.2230 24.5835 7.2490 25.6770 ;
        RECT 7.1150 24.5835 7.1410 25.6770 ;
        RECT 7.0070 24.5835 7.0330 25.6770 ;
        RECT 6.8990 24.5835 6.9250 25.6770 ;
        RECT 6.7910 24.5835 6.8170 25.6770 ;
        RECT 6.6830 24.5835 6.7090 25.6770 ;
        RECT 6.5750 24.5835 6.6010 25.6770 ;
        RECT 6.4670 24.5835 6.4930 25.6770 ;
        RECT 6.3590 24.5835 6.3850 25.6770 ;
        RECT 6.2510 24.5835 6.2770 25.6770 ;
        RECT 6.1430 24.5835 6.1690 25.6770 ;
        RECT 6.0350 24.5835 6.0610 25.6770 ;
        RECT 5.9270 24.5835 5.9530 25.6770 ;
        RECT 5.7140 24.5835 5.7910 25.6770 ;
        RECT 3.8210 24.5835 3.8980 25.6770 ;
        RECT 3.6590 24.5835 3.6850 25.6770 ;
        RECT 3.5510 24.5835 3.5770 25.6770 ;
        RECT 3.4430 24.5835 3.4690 25.6770 ;
        RECT 3.3350 24.5835 3.3610 25.6770 ;
        RECT 3.2270 24.5835 3.2530 25.6770 ;
        RECT 3.1190 24.5835 3.1450 25.6770 ;
        RECT 3.0110 24.5835 3.0370 25.6770 ;
        RECT 2.9030 24.5835 2.9290 25.6770 ;
        RECT 2.7950 24.5835 2.8210 25.6770 ;
        RECT 2.6870 24.5835 2.7130 25.6770 ;
        RECT 2.5790 24.5835 2.6050 25.6770 ;
        RECT 2.4710 24.5835 2.4970 25.6770 ;
        RECT 2.3630 24.5835 2.3890 25.6770 ;
        RECT 2.2550 24.5835 2.2810 25.6770 ;
        RECT 2.1470 24.5835 2.1730 25.6770 ;
        RECT 2.0390 24.5835 2.0650 25.6770 ;
        RECT 1.9310 24.5835 1.9570 25.6770 ;
        RECT 1.8230 24.5835 1.8490 25.6770 ;
        RECT 1.7150 24.5835 1.7410 25.6770 ;
        RECT 1.6070 24.5835 1.6330 25.6770 ;
        RECT 1.4990 24.5835 1.5250 25.6770 ;
        RECT 1.3910 24.5835 1.4170 25.6770 ;
        RECT 1.2830 24.5835 1.3090 25.6770 ;
        RECT 1.1750 24.5835 1.2010 25.6770 ;
        RECT 1.0670 24.5835 1.0930 25.6770 ;
        RECT 0.9590 24.5835 0.9850 25.6770 ;
        RECT 0.8510 24.5835 0.8770 25.6770 ;
        RECT 0.7430 24.5835 0.7690 25.6770 ;
        RECT 0.6350 24.5835 0.6610 25.6770 ;
        RECT 0.5270 24.5835 0.5530 25.6770 ;
        RECT 0.4190 24.5835 0.4450 25.6770 ;
        RECT 0.3110 24.5835 0.3370 25.6770 ;
        RECT 0.2030 24.5835 0.2290 25.6770 ;
        RECT 0.0000 24.5835 0.0850 25.6770 ;
  LAYER V3  ;
      RECT 0.0000 1.2200 9.6120 1.3500 ;
      RECT 9.4950 0.2565 9.6120 1.3500 ;
      RECT 5.8410 1.1240 9.4770 1.3500 ;
      RECT 4.5090 1.1240 5.8230 1.3500 ;
      RECT 3.7890 0.2565 4.4190 1.3500 ;
      RECT 0.1350 1.1240 3.7710 1.3500 ;
      RECT 0.0000 0.2565 0.1170 1.3500 ;
      RECT 9.4590 0.2565 9.6120 1.1720 ;
      RECT 5.8950 0.2565 9.4410 1.3500 ;
      RECT 5.1480 0.2565 5.8770 1.1720 ;
      RECT 4.9860 0.4520 5.1120 1.3500 ;
      RECT 3.7350 0.3560 4.9590 1.1720 ;
      RECT 0.1710 0.2565 3.7170 1.3500 ;
      RECT 0.0000 0.2565 0.1530 1.1720 ;
      RECT 5.0940 0.2565 9.6120 1.0760 ;
      RECT 0.0000 0.3560 5.0760 1.0760 ;
      RECT 4.8690 0.2565 9.6120 0.4280 ;
      RECT 0.0000 0.2565 4.8510 1.0760 ;
      RECT 0.0000 0.2565 9.6120 0.3320 ;
      RECT 0.0000 2.3000 9.6120 2.4300 ;
      RECT 9.4950 1.3365 9.6120 2.4300 ;
      RECT 5.8410 2.2040 9.4770 2.4300 ;
      RECT 4.5090 2.2040 5.8230 2.4300 ;
      RECT 3.7890 1.3365 4.4190 2.4300 ;
      RECT 0.1350 2.2040 3.7710 2.4300 ;
      RECT 0.0000 1.3365 0.1170 2.4300 ;
      RECT 9.4590 1.3365 9.6120 2.2520 ;
      RECT 5.8950 1.3365 9.4410 2.4300 ;
      RECT 5.1480 1.3365 5.8770 2.2520 ;
      RECT 4.9860 1.5320 5.1120 2.4300 ;
      RECT 3.7350 1.4360 4.9590 2.2520 ;
      RECT 0.1710 1.3365 3.7170 2.4300 ;
      RECT 0.0000 1.3365 0.1530 2.2520 ;
      RECT 5.0940 1.3365 9.6120 2.1560 ;
      RECT 0.0000 1.4360 5.0760 2.1560 ;
      RECT 4.8690 1.3365 9.6120 1.5080 ;
      RECT 0.0000 1.3365 4.8510 2.1560 ;
      RECT 0.0000 1.3365 9.6120 1.4120 ;
      RECT 0.0000 3.3800 9.6120 3.5100 ;
      RECT 9.4950 2.4165 9.6120 3.5100 ;
      RECT 5.8410 3.2840 9.4770 3.5100 ;
      RECT 4.5090 3.2840 5.8230 3.5100 ;
      RECT 3.7890 2.4165 4.4190 3.5100 ;
      RECT 0.1350 3.2840 3.7710 3.5100 ;
      RECT 0.0000 2.4165 0.1170 3.5100 ;
      RECT 9.4590 2.4165 9.6120 3.3320 ;
      RECT 5.8950 2.4165 9.4410 3.5100 ;
      RECT 5.1480 2.4165 5.8770 3.3320 ;
      RECT 4.9860 2.6120 5.1120 3.5100 ;
      RECT 3.7350 2.5160 4.9590 3.3320 ;
      RECT 0.1710 2.4165 3.7170 3.5100 ;
      RECT 0.0000 2.4165 0.1530 3.3320 ;
      RECT 5.0940 2.4165 9.6120 3.2360 ;
      RECT 0.0000 2.5160 5.0760 3.2360 ;
      RECT 4.8690 2.4165 9.6120 2.5880 ;
      RECT 0.0000 2.4165 4.8510 3.2360 ;
      RECT 0.0000 2.4165 9.6120 2.4920 ;
      RECT 0.0000 4.4600 9.6120 4.5900 ;
      RECT 9.4950 3.4965 9.6120 4.5900 ;
      RECT 5.8410 4.3640 9.4770 4.5900 ;
      RECT 4.5090 4.3640 5.8230 4.5900 ;
      RECT 3.7890 3.4965 4.4190 4.5900 ;
      RECT 0.1350 4.3640 3.7710 4.5900 ;
      RECT 0.0000 3.4965 0.1170 4.5900 ;
      RECT 9.4590 3.4965 9.6120 4.4120 ;
      RECT 5.8950 3.4965 9.4410 4.5900 ;
      RECT 5.1480 3.4965 5.8770 4.4120 ;
      RECT 4.9860 3.6920 5.1120 4.5900 ;
      RECT 3.7350 3.5960 4.9590 4.4120 ;
      RECT 0.1710 3.4965 3.7170 4.5900 ;
      RECT 0.0000 3.4965 0.1530 4.4120 ;
      RECT 5.0940 3.4965 9.6120 4.3160 ;
      RECT 0.0000 3.5960 5.0760 4.3160 ;
      RECT 4.8690 3.4965 9.6120 3.6680 ;
      RECT 0.0000 3.4965 4.8510 4.3160 ;
      RECT 0.0000 3.4965 9.6120 3.5720 ;
      RECT 0.0000 5.5400 9.6120 5.6700 ;
      RECT 9.4950 4.5765 9.6120 5.6700 ;
      RECT 5.8410 5.4440 9.4770 5.6700 ;
      RECT 4.5090 5.4440 5.8230 5.6700 ;
      RECT 3.7890 4.5765 4.4190 5.6700 ;
      RECT 0.1350 5.4440 3.7710 5.6700 ;
      RECT 0.0000 4.5765 0.1170 5.6700 ;
      RECT 9.4590 4.5765 9.6120 5.4920 ;
      RECT 5.8950 4.5765 9.4410 5.6700 ;
      RECT 5.1480 4.5765 5.8770 5.4920 ;
      RECT 4.9860 4.7720 5.1120 5.6700 ;
      RECT 3.7350 4.6760 4.9590 5.4920 ;
      RECT 0.1710 4.5765 3.7170 5.6700 ;
      RECT 0.0000 4.5765 0.1530 5.4920 ;
      RECT 5.0940 4.5765 9.6120 5.3960 ;
      RECT 0.0000 4.6760 5.0760 5.3960 ;
      RECT 4.8690 4.5765 9.6120 4.7480 ;
      RECT 0.0000 4.5765 4.8510 5.3960 ;
      RECT 0.0000 4.5765 9.6120 4.6520 ;
      RECT 0.0000 6.6200 9.6120 6.7500 ;
      RECT 9.4950 5.6565 9.6120 6.7500 ;
      RECT 5.8410 6.5240 9.4770 6.7500 ;
      RECT 4.5090 6.5240 5.8230 6.7500 ;
      RECT 3.7890 5.6565 4.4190 6.7500 ;
      RECT 0.1350 6.5240 3.7710 6.7500 ;
      RECT 0.0000 5.6565 0.1170 6.7500 ;
      RECT 9.4590 5.6565 9.6120 6.5720 ;
      RECT 5.8950 5.6565 9.4410 6.7500 ;
      RECT 5.1480 5.6565 5.8770 6.5720 ;
      RECT 4.9860 5.8520 5.1120 6.7500 ;
      RECT 3.7350 5.7560 4.9590 6.5720 ;
      RECT 0.1710 5.6565 3.7170 6.7500 ;
      RECT 0.0000 5.6565 0.1530 6.5720 ;
      RECT 5.0940 5.6565 9.6120 6.4760 ;
      RECT 0.0000 5.7560 5.0760 6.4760 ;
      RECT 4.8690 5.6565 9.6120 5.8280 ;
      RECT 0.0000 5.6565 4.8510 6.4760 ;
      RECT 0.0000 5.6565 9.6120 5.7320 ;
      RECT 0.0000 7.7000 9.6120 7.8300 ;
      RECT 9.4950 6.7365 9.6120 7.8300 ;
      RECT 5.8410 7.6040 9.4770 7.8300 ;
      RECT 4.5090 7.6040 5.8230 7.8300 ;
      RECT 3.7890 6.7365 4.4190 7.8300 ;
      RECT 0.1350 7.6040 3.7710 7.8300 ;
      RECT 0.0000 6.7365 0.1170 7.8300 ;
      RECT 9.4590 6.7365 9.6120 7.6520 ;
      RECT 5.8950 6.7365 9.4410 7.8300 ;
      RECT 5.1480 6.7365 5.8770 7.6520 ;
      RECT 4.9860 6.9320 5.1120 7.8300 ;
      RECT 3.7350 6.8360 4.9590 7.6520 ;
      RECT 0.1710 6.7365 3.7170 7.8300 ;
      RECT 0.0000 6.7365 0.1530 7.6520 ;
      RECT 5.0940 6.7365 9.6120 7.5560 ;
      RECT 0.0000 6.8360 5.0760 7.5560 ;
      RECT 4.8690 6.7365 9.6120 6.9080 ;
      RECT 0.0000 6.7365 4.8510 7.5560 ;
      RECT 0.0000 6.7365 9.6120 6.8120 ;
      RECT 0.0000 8.7800 9.6120 8.9100 ;
      RECT 9.4950 7.8165 9.6120 8.9100 ;
      RECT 5.8410 8.6840 9.4770 8.9100 ;
      RECT 4.5090 8.6840 5.8230 8.9100 ;
      RECT 3.7890 7.8165 4.4190 8.9100 ;
      RECT 0.1350 8.6840 3.7710 8.9100 ;
      RECT 0.0000 7.8165 0.1170 8.9100 ;
      RECT 9.4590 7.8165 9.6120 8.7320 ;
      RECT 5.8950 7.8165 9.4410 8.9100 ;
      RECT 5.1480 7.8165 5.8770 8.7320 ;
      RECT 4.9860 8.0120 5.1120 8.9100 ;
      RECT 3.7350 7.9160 4.9590 8.7320 ;
      RECT 0.1710 7.8165 3.7170 8.9100 ;
      RECT 0.0000 7.8165 0.1530 8.7320 ;
      RECT 5.0940 7.8165 9.6120 8.6360 ;
      RECT 0.0000 7.9160 5.0760 8.6360 ;
      RECT 4.8690 7.8165 9.6120 7.9880 ;
      RECT 0.0000 7.8165 4.8510 8.6360 ;
      RECT 0.0000 7.8165 9.6120 7.8920 ;
      RECT 0.0000 16.2030 9.6120 17.5365 ;
      RECT 7.3530 8.8830 9.6120 17.5365 ;
      RECT 5.1530 12.7470 9.6120 17.5365 ;
      RECT 6.0570 10.1550 9.6120 17.5365 ;
      RECT 5.1010 8.8830 5.1350 17.5365 ;
      RECT 5.0490 8.8830 5.0830 17.5365 ;
      RECT 4.9970 8.8830 5.0310 17.5365 ;
      RECT 4.9450 8.8830 4.9790 17.5365 ;
      RECT 0.0000 15.7710 4.9270 17.5365 ;
      RECT 4.6850 13.0350 9.6120 15.9870 ;
      RECT 4.6330 8.8830 4.6670 17.5365 ;
      RECT 4.5810 8.8830 4.6150 17.5365 ;
      RECT 4.5290 8.8830 4.5630 17.5365 ;
      RECT 4.4770 8.8830 4.5110 17.5365 ;
      RECT 0.0000 10.4430 4.4590 17.5365 ;
      RECT 0.0000 12.6030 4.9270 15.5550 ;
      RECT 4.6850 9.8670 5.8230 12.8190 ;
      RECT 5.8410 10.3470 9.6120 17.5365 ;
      RECT 5.1930 8.9630 6.0390 12.7230 ;
      RECT 4.0050 9.4350 4.7790 12.3870 ;
      RECT 3.7890 9.5790 4.4590 17.5365 ;
      RECT 0.0000 10.1550 3.7710 17.5365 ;
      RECT 3.3570 8.8830 3.8070 10.4190 ;
      RECT 7.1370 8.8830 7.3350 17.5365 ;
      RECT 3.3570 9.9630 7.1190 10.3230 ;
      RECT 2.4930 9.5790 3.3390 17.5365 ;
      RECT 0.0000 9.8670 2.4750 17.5365 ;
      RECT 6.9210 8.8830 9.6120 10.1310 ;
      RECT 6.7050 9.5790 9.6120 10.1310 ;
      RECT 0.0000 9.8670 6.6870 10.1310 ;
      RECT 6.4890 8.8830 6.9030 9.9390 ;
      RECT 5.1530 9.5790 9.6120 9.9390 ;
      RECT 0.1710 9.5790 4.9270 10.1310 ;
      RECT 4.6850 9.5310 4.9270 17.5365 ;
      RECT 0.0000 9.4350 0.1530 17.5365 ;
      RECT 4.7970 8.8830 5.1750 9.6510 ;
      RECT 5.1930 9.5310 6.4710 10.3230 ;
      RECT 3.1410 9.5310 3.9870 10.1310 ;
      RECT 2.7090 9.5310 3.1230 17.5365 ;
      RECT 0.0000 9.4350 2.6910 9.6510 ;
      RECT 6.2730 8.8830 9.6120 9.5550 ;
      RECT 4.7970 8.9630 6.2550 9.5550 ;
      RECT 3.8250 9.4350 4.7790 9.5550 ;
      RECT 2.9250 8.8830 3.8070 9.5550 ;
      RECT 0.0000 9.4350 2.9070 9.5550 ;
      RECT 5.8410 8.8830 9.6120 9.5070 ;
      RECT 4.6850 8.9630 9.6120 9.5070 ;
      RECT 0.1350 8.8830 4.4590 9.5070 ;
      RECT 0.0000 8.8830 0.1170 17.5365 ;
      RECT 0.0000 8.8830 5.8230 9.2190 ;
      RECT 0.0000 8.8830 9.6120 8.9390 ;
        RECT 0.0000 17.9870 9.6120 18.1170 ;
        RECT 9.4950 17.0235 9.6120 18.1170 ;
        RECT 5.8410 17.8910 9.4770 18.1170 ;
        RECT 4.5090 17.8910 5.8230 18.1170 ;
        RECT 3.7890 17.0235 4.4190 18.1170 ;
        RECT 0.1350 17.8910 3.7710 18.1170 ;
        RECT 0.0000 17.0235 0.1170 18.1170 ;
        RECT 9.4590 17.0235 9.6120 17.9390 ;
        RECT 5.8950 17.0235 9.4410 18.1170 ;
        RECT 5.1480 17.0235 5.8770 17.9390 ;
        RECT 4.9860 17.2190 5.1120 18.1170 ;
        RECT 3.7350 17.1230 4.9590 17.9390 ;
        RECT 0.1710 17.0235 3.7170 18.1170 ;
        RECT 0.0000 17.0235 0.1530 17.9390 ;
        RECT 5.0940 17.0235 9.6120 17.8430 ;
        RECT 0.0000 17.1230 5.0760 17.8430 ;
        RECT 4.8690 17.0235 9.6120 17.1950 ;
        RECT 0.0000 17.0235 4.8510 17.8430 ;
        RECT 0.0000 17.0235 9.6120 17.0990 ;
        RECT 0.0000 19.0670 9.6120 19.1970 ;
        RECT 9.4950 18.1035 9.6120 19.1970 ;
        RECT 5.8410 18.9710 9.4770 19.1970 ;
        RECT 4.5090 18.9710 5.8230 19.1970 ;
        RECT 3.7890 18.1035 4.4190 19.1970 ;
        RECT 0.1350 18.9710 3.7710 19.1970 ;
        RECT 0.0000 18.1035 0.1170 19.1970 ;
        RECT 9.4590 18.1035 9.6120 19.0190 ;
        RECT 5.8950 18.1035 9.4410 19.1970 ;
        RECT 5.1480 18.1035 5.8770 19.0190 ;
        RECT 4.9860 18.2990 5.1120 19.1970 ;
        RECT 3.7350 18.2030 4.9590 19.0190 ;
        RECT 0.1710 18.1035 3.7170 19.1970 ;
        RECT 0.0000 18.1035 0.1530 19.0190 ;
        RECT 5.0940 18.1035 9.6120 18.9230 ;
        RECT 0.0000 18.2030 5.0760 18.9230 ;
        RECT 4.8690 18.1035 9.6120 18.2750 ;
        RECT 0.0000 18.1035 4.8510 18.9230 ;
        RECT 0.0000 18.1035 9.6120 18.1790 ;
        RECT 0.0000 20.1470 9.6120 20.2770 ;
        RECT 9.4950 19.1835 9.6120 20.2770 ;
        RECT 5.8410 20.0510 9.4770 20.2770 ;
        RECT 4.5090 20.0510 5.8230 20.2770 ;
        RECT 3.7890 19.1835 4.4190 20.2770 ;
        RECT 0.1350 20.0510 3.7710 20.2770 ;
        RECT 0.0000 19.1835 0.1170 20.2770 ;
        RECT 9.4590 19.1835 9.6120 20.0990 ;
        RECT 5.8950 19.1835 9.4410 20.2770 ;
        RECT 5.1480 19.1835 5.8770 20.0990 ;
        RECT 4.9860 19.3790 5.1120 20.2770 ;
        RECT 3.7350 19.2830 4.9590 20.0990 ;
        RECT 0.1710 19.1835 3.7170 20.2770 ;
        RECT 0.0000 19.1835 0.1530 20.0990 ;
        RECT 5.0940 19.1835 9.6120 20.0030 ;
        RECT 0.0000 19.2830 5.0760 20.0030 ;
        RECT 4.8690 19.1835 9.6120 19.3550 ;
        RECT 0.0000 19.1835 4.8510 20.0030 ;
        RECT 0.0000 19.1835 9.6120 19.2590 ;
        RECT 0.0000 21.2270 9.6120 21.3570 ;
        RECT 9.4950 20.2635 9.6120 21.3570 ;
        RECT 5.8410 21.1310 9.4770 21.3570 ;
        RECT 4.5090 21.1310 5.8230 21.3570 ;
        RECT 3.7890 20.2635 4.4190 21.3570 ;
        RECT 0.1350 21.1310 3.7710 21.3570 ;
        RECT 0.0000 20.2635 0.1170 21.3570 ;
        RECT 9.4590 20.2635 9.6120 21.1790 ;
        RECT 5.8950 20.2635 9.4410 21.3570 ;
        RECT 5.1480 20.2635 5.8770 21.1790 ;
        RECT 4.9860 20.4590 5.1120 21.3570 ;
        RECT 3.7350 20.3630 4.9590 21.1790 ;
        RECT 0.1710 20.2635 3.7170 21.3570 ;
        RECT 0.0000 20.2635 0.1530 21.1790 ;
        RECT 5.0940 20.2635 9.6120 21.0830 ;
        RECT 0.0000 20.3630 5.0760 21.0830 ;
        RECT 4.8690 20.2635 9.6120 20.4350 ;
        RECT 0.0000 20.2635 4.8510 21.0830 ;
        RECT 0.0000 20.2635 9.6120 20.3390 ;
        RECT 0.0000 22.3070 9.6120 22.4370 ;
        RECT 9.4950 21.3435 9.6120 22.4370 ;
        RECT 5.8410 22.2110 9.4770 22.4370 ;
        RECT 4.5090 22.2110 5.8230 22.4370 ;
        RECT 3.7890 21.3435 4.4190 22.4370 ;
        RECT 0.1350 22.2110 3.7710 22.4370 ;
        RECT 0.0000 21.3435 0.1170 22.4370 ;
        RECT 9.4590 21.3435 9.6120 22.2590 ;
        RECT 5.8950 21.3435 9.4410 22.4370 ;
        RECT 5.1480 21.3435 5.8770 22.2590 ;
        RECT 4.9860 21.5390 5.1120 22.4370 ;
        RECT 3.7350 21.4430 4.9590 22.2590 ;
        RECT 0.1710 21.3435 3.7170 22.4370 ;
        RECT 0.0000 21.3435 0.1530 22.2590 ;
        RECT 5.0940 21.3435 9.6120 22.1630 ;
        RECT 0.0000 21.4430 5.0760 22.1630 ;
        RECT 4.8690 21.3435 9.6120 21.5150 ;
        RECT 0.0000 21.3435 4.8510 22.1630 ;
        RECT 0.0000 21.3435 9.6120 21.4190 ;
        RECT 0.0000 23.3870 9.6120 23.5170 ;
        RECT 9.4950 22.4235 9.6120 23.5170 ;
        RECT 5.8410 23.2910 9.4770 23.5170 ;
        RECT 4.5090 23.2910 5.8230 23.5170 ;
        RECT 3.7890 22.4235 4.4190 23.5170 ;
        RECT 0.1350 23.2910 3.7710 23.5170 ;
        RECT 0.0000 22.4235 0.1170 23.5170 ;
        RECT 9.4590 22.4235 9.6120 23.3390 ;
        RECT 5.8950 22.4235 9.4410 23.5170 ;
        RECT 5.1480 22.4235 5.8770 23.3390 ;
        RECT 4.9860 22.6190 5.1120 23.5170 ;
        RECT 3.7350 22.5230 4.9590 23.3390 ;
        RECT 0.1710 22.4235 3.7170 23.5170 ;
        RECT 0.0000 22.4235 0.1530 23.3390 ;
        RECT 5.0940 22.4235 9.6120 23.2430 ;
        RECT 0.0000 22.5230 5.0760 23.2430 ;
        RECT 4.8690 22.4235 9.6120 22.5950 ;
        RECT 0.0000 22.4235 4.8510 23.2430 ;
        RECT 0.0000 22.4235 9.6120 22.4990 ;
        RECT 0.0000 24.4670 9.6120 24.5970 ;
        RECT 9.4950 23.5035 9.6120 24.5970 ;
        RECT 5.8410 24.3710 9.4770 24.5970 ;
        RECT 4.5090 24.3710 5.8230 24.5970 ;
        RECT 3.7890 23.5035 4.4190 24.5970 ;
        RECT 0.1350 24.3710 3.7710 24.5970 ;
        RECT 0.0000 23.5035 0.1170 24.5970 ;
        RECT 9.4590 23.5035 9.6120 24.4190 ;
        RECT 5.8950 23.5035 9.4410 24.5970 ;
        RECT 5.1480 23.5035 5.8770 24.4190 ;
        RECT 4.9860 23.6990 5.1120 24.5970 ;
        RECT 3.7350 23.6030 4.9590 24.4190 ;
        RECT 0.1710 23.5035 3.7170 24.5970 ;
        RECT 0.0000 23.5035 0.1530 24.4190 ;
        RECT 5.0940 23.5035 9.6120 24.3230 ;
        RECT 0.0000 23.6030 5.0760 24.3230 ;
        RECT 4.8690 23.5035 9.6120 23.6750 ;
        RECT 0.0000 23.5035 4.8510 24.3230 ;
        RECT 0.0000 23.5035 9.6120 23.5790 ;
        RECT 0.0000 25.5470 9.6120 25.6770 ;
        RECT 9.4950 24.5835 9.6120 25.6770 ;
        RECT 5.8410 25.4510 9.4770 25.6770 ;
        RECT 4.5090 25.4510 5.8230 25.6770 ;
        RECT 3.7890 24.5835 4.4190 25.6770 ;
        RECT 0.1350 25.4510 3.7710 25.6770 ;
        RECT 0.0000 24.5835 0.1170 25.6770 ;
        RECT 9.4590 24.5835 9.6120 25.4990 ;
        RECT 5.8950 24.5835 9.4410 25.6770 ;
        RECT 5.1480 24.5835 5.8770 25.4990 ;
        RECT 4.9860 24.7790 5.1120 25.6770 ;
        RECT 3.7350 24.6830 4.9590 25.4990 ;
        RECT 0.1710 24.5835 3.7170 25.6770 ;
        RECT 0.0000 24.5835 0.1530 25.4990 ;
        RECT 5.0940 24.5835 9.6120 25.4030 ;
        RECT 0.0000 24.6830 5.0760 25.4030 ;
        RECT 4.8690 24.5835 9.6120 24.7550 ;
        RECT 0.0000 24.5835 4.8510 25.4030 ;
        RECT 0.0000 24.5835 9.6120 24.6590 ;
  LAYER M4  ;
      RECT 1.6070 10.5960 8.0025 10.6200 ;
      RECT 1.6070 10.8840 8.0025 10.9080 ;
      RECT 1.6070 11.2680 8.0025 11.2920 ;
      RECT 1.6070 11.3640 8.0025 11.3880 ;
      RECT 1.6070 11.7000 8.0025 11.7240 ;
      RECT 7.4990 9.5550 7.5830 9.5790 ;
      RECT 7.3190 9.9870 7.4360 10.0110 ;
      RECT 7.3190 10.6440 7.4360 10.6680 ;
      RECT 7.3190 10.9320 7.4360 10.9560 ;
      RECT 6.6785 9.9870 7.2480 10.0110 ;
      RECT 6.7430 10.7640 6.8510 10.7880 ;
      RECT 5.4070 11.1390 6.5000 11.1630 ;
      RECT 6.0950 10.7070 6.1790 10.7310 ;
      RECT 5.3110 11.9070 6.1790 11.9310 ;
      RECT 6.0950 12.0030 6.1790 12.0270 ;
      RECT 5.9170 10.2270 6.0010 10.2510 ;
      RECT 5.8790 11.5710 5.9630 11.5950 ;
      RECT 5.7010 10.1310 5.7850 10.1550 ;
      RECT 5.4870 8.8430 5.7500 8.8670 ;
      RECT 5.4870 17.4830 5.7500 17.5070 ;
      RECT 5.5030 11.6190 5.7470 11.6430 ;
      RECT 5.6630 11.7630 5.7470 11.7870 ;
      RECT 4.2070 12.0030 5.7470 12.0270 ;
      RECT 5.6630 12.2910 5.7470 12.3150 ;
      RECT 5.4290 17.3870 5.6920 17.4110 ;
      RECT 5.4280 8.7470 5.6910 8.7710 ;
      RECT 5.3900 8.6510 5.6530 8.6750 ;
      RECT 5.3900 17.1950 5.6530 17.2190 ;
      RECT 5.5550 12.7230 5.6390 12.7470 ;
      RECT 4.7830 13.1070 5.6390 13.1310 ;
      RECT 5.1670 15.3630 5.6390 15.3870 ;
      RECT 5.5550 15.4590 5.6390 15.4830 ;
      RECT 5.3420 8.5550 5.6050 8.5790 ;
      RECT 5.3420 17.0990 5.6050 17.1230 ;
      RECT 5.1190 14.4510 5.5640 14.4750 ;
      RECT 5.2980 8.4590 5.5610 8.4830 ;
      RECT 5.2980 17.4350 5.5610 17.4590 ;
      RECT 5.2490 8.7950 5.5120 8.8190 ;
      RECT 5.2490 17.3390 5.5120 17.3630 ;
      RECT 5.3800 11.7630 5.5010 11.7870 ;
      RECT 5.3590 13.8750 5.4920 13.8990 ;
      RECT 5.2020 8.6990 5.4650 8.7230 ;
      RECT 5.2020 17.2430 5.4650 17.2670 ;
      RECT 5.1670 8.4110 5.4300 8.4350 ;
      RECT 5.1670 17.1470 5.4300 17.1710 ;
      RECT 4.3510 15.4590 5.4200 15.4830 ;
      RECT 5.3360 16.6110 5.4200 16.6350 ;
      RECT 5.1110 8.2670 5.3740 8.2910 ;
      RECT 5.1110 17.0510 5.3740 17.0750 ;
      RECT 5.2630 12.7230 5.3480 12.7470 ;
      RECT 4.1590 13.2990 5.2760 13.3230 ;
      RECT 4.8040 11.1390 5.2610 11.1630 ;
      RECT 4.6310 8.9870 4.8980 9.0110 ;
      RECT 4.6310 16.9070 4.8980 16.9310 ;
      RECT 4.7680 12.6750 4.8770 12.6990 ;
      RECT 4.6080 8.8910 4.8500 8.9150 ;
      RECT 4.6080 17.5310 4.8500 17.5550 ;
      RECT 4.5520 8.4110 4.7940 8.4350 ;
      RECT 4.5810 17.6270 4.7940 17.6510 ;
      RECT 4.6970 12.2910 4.7810 12.3150 ;
      RECT 4.4980 8.5070 4.7460 8.5310 ;
      RECT 4.4980 17.4830 4.7460 17.5070 ;
      RECT 4.2640 14.8830 4.6850 14.9070 ;
      RECT 4.2320 8.8430 4.4990 8.8670 ;
      RECT 4.2320 17.6270 4.4990 17.6510 ;
      RECT 4.3720 13.4430 4.4930 13.4670 ;
      RECT 4.3640 16.6110 4.4480 16.6350 ;
      RECT 4.1980 8.7470 4.4450 8.7710 ;
      RECT 4.1310 17.1950 4.4450 17.2190 ;
      RECT 4.1720 8.6510 4.4020 8.6750 ;
      RECT 4.1600 17.5310 4.4020 17.5550 ;
      RECT 4.1190 8.5550 4.3490 8.5790 ;
      RECT 4.2650 15.0270 4.3490 15.0510 ;
      RECT 4.0690 17.0990 4.3490 17.1230 ;
      RECT 4.0740 8.4590 4.3040 8.4830 ;
      RECT 4.0740 17.4350 4.3040 17.4590 ;
      RECT 3.1120 12.2910 4.3010 12.3150 ;
      RECT 4.0360 8.6990 4.2660 8.7230 ;
      RECT 4.0360 17.3390 4.2660 17.3630 ;
      RECT 4.0180 8.6030 4.2110 8.6270 ;
      RECT 4.0180 17.2430 4.2110 17.2670 ;
      RECT 3.9690 8.5070 4.1620 8.5310 ;
      RECT 3.9690 17.1470 4.1620 17.1710 ;
      RECT 3.9730 13.2030 4.1570 13.2270 ;
      RECT 3.9170 8.4110 4.1100 8.4350 ;
      RECT 3.9170 17.0510 4.1100 17.0750 ;
      RECT 3.4330 10.5150 4.1090 10.5390 ;
      RECT 3.9730 13.2990 4.0570 13.3230 ;
      RECT 3.7040 8.9390 3.9670 8.9630 ;
      RECT 3.7580 12.7230 3.8700 12.7470 ;
      RECT 3.3950 10.7070 3.4790 10.7310 ;
  LAYER V4  ;
      RECT 7.5480 9.5550 7.5720 9.5790 ;
      RECT 7.5480 10.5960 7.5720 10.6200 ;
      RECT 7.3800 9.9870 7.4040 10.0110 ;
      RECT 7.3800 10.6440 7.4040 10.6680 ;
      RECT 7.3800 10.9320 7.4040 10.9560 ;
      RECT 6.7560 9.9870 6.7800 10.0110 ;
      RECT 6.7560 10.7640 6.7800 10.7880 ;
      RECT 6.1440 10.7070 6.1680 10.7310 ;
      RECT 6.1440 10.8840 6.1680 10.9080 ;
      RECT 6.1440 11.9070 6.1680 11.9310 ;
      RECT 6.1440 12.0030 6.1680 12.0270 ;
      RECT 5.9280 10.2270 5.9520 10.2510 ;
      RECT 5.9280 11.2680 5.9520 11.2920 ;
      RECT 5.9280 11.5710 5.9520 11.5950 ;
      RECT 5.9280 11.7000 5.9520 11.7240 ;
      RECT 5.7120 10.1310 5.7360 10.1550 ;
      RECT 5.7120 11.3640 5.7360 11.3880 ;
      RECT 5.7120 11.6190 5.7360 11.6430 ;
      RECT 5.7120 11.7630 5.7360 11.7870 ;
      RECT 5.7120 12.0030 5.7360 12.0270 ;
      RECT 5.7120 12.2910 5.7360 12.3150 ;
      RECT 5.6040 12.7230 5.6280 12.7470 ;
      RECT 5.6040 13.1070 5.6280 13.1310 ;
      RECT 5.6040 15.3630 5.6280 15.3870 ;
      RECT 5.6040 15.4590 5.6280 15.4830 ;
      RECT 5.5140 8.8430 5.5380 8.8670 ;
      RECT 5.5140 11.6190 5.5380 11.6430 ;
      RECT 5.5140 17.4830 5.5380 17.5070 ;
      RECT 5.4660 8.7470 5.4900 8.7710 ;
      RECT 5.4660 11.7630 5.4900 11.7870 ;
      RECT 5.4660 17.3870 5.4900 17.4110 ;
      RECT 5.4180 8.6510 5.4420 8.6750 ;
      RECT 5.4180 11.1390 5.4420 11.1630 ;
      RECT 5.4180 17.1950 5.4420 17.2190 ;
      RECT 5.3700 8.5550 5.3940 8.5790 ;
      RECT 5.3700 13.8750 5.3940 13.8990 ;
      RECT 5.3700 16.6110 5.3940 16.6350 ;
      RECT 5.3700 17.0990 5.3940 17.1230 ;
      RECT 5.3220 8.4590 5.3460 8.4830 ;
      RECT 5.3220 11.9070 5.3460 11.9310 ;
      RECT 5.3220 17.4350 5.3460 17.4590 ;
      RECT 5.2740 8.7950 5.2980 8.8190 ;
      RECT 5.2740 12.7230 5.2980 12.7470 ;
      RECT 5.2740 17.3390 5.2980 17.3630 ;
      RECT 5.2260 8.6990 5.2500 8.7230 ;
      RECT 5.2260 11.1390 5.2500 11.1630 ;
      RECT 5.2260 17.2430 5.2500 17.2670 ;
      RECT 5.1780 8.4110 5.2020 8.4350 ;
      RECT 5.1780 15.3630 5.2020 15.3870 ;
      RECT 5.1780 17.1470 5.2020 17.1710 ;
      RECT 5.1300 8.2670 5.1540 8.2910 ;
      RECT 5.1300 14.4510 5.1540 14.4750 ;
      RECT 5.1300 17.0510 5.1540 17.0750 ;
      RECT 4.8420 8.9870 4.8660 9.0110 ;
      RECT 4.8420 12.6750 4.8660 12.6990 ;
      RECT 4.8420 16.9070 4.8660 16.9310 ;
      RECT 4.7940 8.8910 4.8180 8.9150 ;
      RECT 4.7940 13.1070 4.8180 13.1310 ;
      RECT 4.7940 17.5310 4.8180 17.5550 ;
      RECT 4.7460 8.4110 4.7700 8.4350 ;
      RECT 4.7460 12.2910 4.7700 12.3150 ;
      RECT 4.7460 17.6270 4.7700 17.6510 ;
      RECT 4.6500 8.5070 4.6740 8.5310 ;
      RECT 4.6500 14.8830 4.6740 14.9070 ;
      RECT 4.6500 17.4830 4.6740 17.5070 ;
      RECT 4.4580 8.8430 4.4820 8.8670 ;
      RECT 4.4580 13.4430 4.4820 13.4670 ;
      RECT 4.4580 17.6270 4.4820 17.6510 ;
      RECT 4.4100 8.7470 4.4340 8.7710 ;
      RECT 4.4100 16.6110 4.4340 16.6350 ;
      RECT 4.4100 17.1950 4.4340 17.2190 ;
      RECT 4.3620 8.6510 4.3860 8.6750 ;
      RECT 4.3620 15.4590 4.3860 15.4830 ;
      RECT 4.3620 17.5310 4.3860 17.5550 ;
      RECT 4.3140 8.5550 4.3380 8.5790 ;
      RECT 4.3140 15.0270 4.3380 15.0510 ;
      RECT 4.3140 17.0990 4.3380 17.1230 ;
      RECT 4.2660 8.4590 4.2900 8.4830 ;
      RECT 4.2660 12.2910 4.2900 12.3150 ;
      RECT 4.2660 17.4350 4.2900 17.4590 ;
      RECT 4.2180 8.6990 4.2420 8.7230 ;
      RECT 4.2180 12.0030 4.2420 12.0270 ;
      RECT 4.2180 17.3390 4.2420 17.3630 ;
      RECT 4.1700 8.6030 4.1940 8.6270 ;
      RECT 4.1700 13.2990 4.1940 13.3230 ;
      RECT 4.1700 17.2430 4.1940 17.2670 ;
      RECT 4.1220 8.5070 4.1460 8.5310 ;
      RECT 4.1220 13.2030 4.1460 13.2270 ;
      RECT 4.1220 17.1470 4.1460 17.1710 ;
      RECT 4.0740 8.4110 4.0980 8.4350 ;
      RECT 4.0740 10.5150 4.0980 10.5390 ;
      RECT 4.0740 17.0510 4.0980 17.0750 ;
      RECT 3.9840 13.2030 4.0080 13.2270 ;
      RECT 3.9840 13.2990 4.0080 13.3230 ;
      RECT 3.8170 8.9390 3.8410 8.9630 ;
      RECT 3.8170 12.7230 3.8410 12.7470 ;
      RECT 3.4440 10.5150 3.4680 10.5390 ;
      RECT 3.4440 10.7070 3.4680 10.7310 ;
  LAYER M5  ;
      RECT 7.5480 9.5440 7.5720 10.6310 ;
      RECT 7.3800 9.9735 7.4040 11.0060 ;
      RECT 6.7560 9.9675 6.7800 10.8000 ;
      RECT 6.1440 10.6960 6.1680 10.9190 ;
      RECT 6.1440 11.8960 6.1680 12.0380 ;
      RECT 5.9280 10.2160 5.9520 11.3030 ;
      RECT 5.9280 11.5600 5.9520 11.7350 ;
      RECT 5.7120 10.1200 5.7360 11.3990 ;
      RECT 5.7120 11.6080 5.7360 11.7980 ;
      RECT 5.7120 11.9920 5.7360 12.3260 ;
      RECT 5.6040 12.7120 5.6280 13.1420 ;
      RECT 5.6040 15.3520 5.6280 15.4940 ;
      RECT 5.5140 9.1800 5.5380 16.7630 ;
      RECT 5.4660 9.1800 5.4900 16.7630 ;
      RECT 5.4180 9.1800 5.4420 16.7630 ;
      RECT 5.3700 9.1800 5.3940 16.7630 ;
      RECT 5.3220 9.1800 5.3460 16.7630 ;
      RECT 5.2740 9.1800 5.2980 16.7630 ;
      RECT 5.2260 9.1800 5.2500 16.7630 ;
      RECT 5.1780 9.1800 5.2020 16.7630 ;
      RECT 5.1300 9.1800 5.1540 16.7630 ;
      RECT 4.8420 8.9180 4.8660 16.9510 ;
      RECT 4.7940 8.3970 4.8180 17.7260 ;
      RECT 4.7460 8.3660 4.7700 17.7250 ;
      RECT 4.6500 8.4120 4.6740 17.7260 ;
      RECT 4.4580 8.4110 4.4820 17.6790 ;
      RECT 4.4100 8.4110 4.4340 17.6790 ;
      RECT 4.3620 8.4110 4.3860 17.6790 ;
      RECT 4.3140 8.4110 4.3380 17.6790 ;
      RECT 4.2660 8.4110 4.2900 17.6790 ;
      RECT 4.2180 8.3820 4.2420 17.6790 ;
      RECT 4.1700 8.3380 4.1940 17.6800 ;
      RECT 4.1220 8.3010 4.1460 17.6810 ;
      RECT 4.0740 8.2410 4.0980 17.6810 ;
      RECT 3.9840 13.1920 4.0080 13.3340 ;
      RECT 3.8170 8.9210 3.8410 12.7650 ;
      RECT 3.4440 10.5040 3.4680 10.7420 ;
  LAYER M2  ;
    RECT 0.108 0.036 9.5040 25.8840 ;
  LAYER M1  ;
    RECT 0.108 0.036 9.5040 25.8840 ;
  END
END srambank_64x4x16_6t122 
