VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_128x4x18_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_128x4x18_6t122 0 0 ;
  SIZE 16.0 BY 28.080000000000002 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.1720 16.4420 1.2200 ;
        RECT 0.0940 2.2520 16.4420 2.3000 ;
        RECT 0.0940 3.3320 16.4420 3.3800 ;
        RECT 0.0940 4.4120 16.4420 4.4600 ;
        RECT 0.0940 5.4920 16.4420 5.5400 ;
        RECT 0.0940 6.5720 16.4420 6.6200 ;
        RECT 0.0940 7.6520 16.4420 7.7000 ;
        RECT 0.0940 8.7320 16.4420 8.7800 ;
        RECT 0.0940 9.8120 16.4420 9.8600 ;
        RECT 3.5640 10.2930 12.9600 10.5090 ;
        RECT 9.1970 13.7970 9.3380 13.8210 ;
        RECT 9.0660 10.0130 9.3290 10.0370 ;
        RECT 7.3980 13.4610 9.1260 13.6770 ;
        RECT 7.3980 16.6290 9.1260 16.8450 ;
        RECT 0.0940 19.0190 16.4420 19.0670 ;
        RECT 0.0940 20.0990 16.4420 20.1470 ;
        RECT 0.0940 21.1790 16.4420 21.2270 ;
        RECT 0.0940 22.2590 16.4420 22.3070 ;
        RECT 0.0940 23.3390 16.4420 23.3870 ;
        RECT 0.0940 24.4190 16.4420 24.4670 ;
        RECT 0.0940 25.4990 16.4420 25.5470 ;
        RECT 0.0940 26.5790 16.4420 26.6270 ;
        RECT 0.0940 27.6590 16.4420 27.7070 ;
      LAYER M3  ;
        RECT 16.3940 0.2165 16.4120 1.3765 ;
        RECT 9.2840 0.2170 9.3020 1.3760 ;
        RECT 7.8800 0.2570 7.9700 1.3710 ;
        RECT 7.2320 0.2170 7.2500 1.3760 ;
        RECT 0.1220 0.2165 0.1400 1.3765 ;
        RECT 16.3940 1.2965 16.4120 2.4565 ;
        RECT 9.2840 1.2970 9.3020 2.4560 ;
        RECT 7.8800 1.3370 7.9700 2.4510 ;
        RECT 7.2320 1.2970 7.2500 2.4560 ;
        RECT 0.1220 1.2965 0.1400 2.4565 ;
        RECT 16.3940 2.3765 16.4120 3.5365 ;
        RECT 9.2840 2.3770 9.3020 3.5360 ;
        RECT 7.8800 2.4170 7.9700 3.5310 ;
        RECT 7.2320 2.3770 7.2500 3.5360 ;
        RECT 0.1220 2.3765 0.1400 3.5365 ;
        RECT 16.3940 3.4565 16.4120 4.6165 ;
        RECT 9.2840 3.4570 9.3020 4.6160 ;
        RECT 7.8800 3.4970 7.9700 4.6110 ;
        RECT 7.2320 3.4570 7.2500 4.6160 ;
        RECT 0.1220 3.4565 0.1400 4.6165 ;
        RECT 16.3940 4.5365 16.4120 5.6965 ;
        RECT 9.2840 4.5370 9.3020 5.6960 ;
        RECT 7.8800 4.5770 7.9700 5.6910 ;
        RECT 7.2320 4.5370 7.2500 5.6960 ;
        RECT 0.1220 4.5365 0.1400 5.6965 ;
        RECT 16.3940 5.6165 16.4120 6.7765 ;
        RECT 9.2840 5.6170 9.3020 6.7760 ;
        RECT 7.8800 5.6570 7.9700 6.7710 ;
        RECT 7.2320 5.6170 7.2500 6.7760 ;
        RECT 0.1220 5.6165 0.1400 6.7765 ;
        RECT 16.3940 6.6965 16.4120 7.8565 ;
        RECT 9.2840 6.6970 9.3020 7.8560 ;
        RECT 7.8800 6.7370 7.9700 7.8510 ;
        RECT 7.2320 6.6970 7.2500 7.8560 ;
        RECT 0.1220 6.6965 0.1400 7.8565 ;
        RECT 16.3940 7.7765 16.4120 8.9365 ;
        RECT 9.2840 7.7770 9.3020 8.9360 ;
        RECT 7.8800 7.8170 7.9700 8.9310 ;
        RECT 7.2320 7.7770 7.2500 8.9360 ;
        RECT 0.1220 7.7765 0.1400 8.9365 ;
        RECT 16.3940 8.8565 16.4120 10.0165 ;
        RECT 9.2840 8.8570 9.3020 10.0160 ;
        RECT 7.8800 8.8970 7.9700 10.0110 ;
        RECT 7.2320 8.8570 7.2500 10.0160 ;
        RECT 0.1220 8.8565 0.1400 10.0165 ;
        RECT 16.3890 9.9305 16.4070 18.1375 ;
        RECT 9.2970 13.7500 9.3150 18.0985 ;
        RECT 9.2790 9.9635 9.2970 10.1015 ;
        RECT 7.9110 10.2540 8.1450 17.8370 ;
        RECT 7.8750 17.7540 7.9650 18.1300 ;
        RECT 7.8750 9.9700 7.9650 10.3460 ;
        RECT 0.1170 9.9305 0.1350 18.1375 ;
        RECT 16.3940 18.0635 16.4120 19.2235 ;
        RECT 9.2840 18.0640 9.3020 19.2230 ;
        RECT 7.8800 18.1040 7.9700 19.2180 ;
        RECT 7.2320 18.0640 7.2500 19.2230 ;
        RECT 0.1220 18.0635 0.1400 19.2235 ;
        RECT 16.3940 19.1435 16.4120 20.3035 ;
        RECT 9.2840 19.1440 9.3020 20.3030 ;
        RECT 7.8800 19.1840 7.9700 20.2980 ;
        RECT 7.2320 19.1440 7.2500 20.3030 ;
        RECT 0.1220 19.1435 0.1400 20.3035 ;
        RECT 16.3940 20.2235 16.4120 21.3835 ;
        RECT 9.2840 20.2240 9.3020 21.3830 ;
        RECT 7.8800 20.2640 7.9700 21.3780 ;
        RECT 7.2320 20.2240 7.2500 21.3830 ;
        RECT 0.1220 20.2235 0.1400 21.3835 ;
        RECT 16.3940 21.3035 16.4120 22.4635 ;
        RECT 9.2840 21.3040 9.3020 22.4630 ;
        RECT 7.8800 21.3440 7.9700 22.4580 ;
        RECT 7.2320 21.3040 7.2500 22.4630 ;
        RECT 0.1220 21.3035 0.1400 22.4635 ;
        RECT 16.3940 22.3835 16.4120 23.5435 ;
        RECT 9.2840 22.3840 9.3020 23.5430 ;
        RECT 7.8800 22.4240 7.9700 23.5380 ;
        RECT 7.2320 22.3840 7.2500 23.5430 ;
        RECT 0.1220 22.3835 0.1400 23.5435 ;
        RECT 16.3940 23.4635 16.4120 24.6235 ;
        RECT 9.2840 23.4640 9.3020 24.6230 ;
        RECT 7.8800 23.5040 7.9700 24.6180 ;
        RECT 7.2320 23.4640 7.2500 24.6230 ;
        RECT 0.1220 23.4635 0.1400 24.6235 ;
        RECT 16.3940 24.5435 16.4120 25.7035 ;
        RECT 9.2840 24.5440 9.3020 25.7030 ;
        RECT 7.8800 24.5840 7.9700 25.6980 ;
        RECT 7.2320 24.5440 7.2500 25.7030 ;
        RECT 0.1220 24.5435 0.1400 25.7035 ;
        RECT 16.3940 25.6235 16.4120 26.7835 ;
        RECT 9.2840 25.6240 9.3020 26.7830 ;
        RECT 7.8800 25.6640 7.9700 26.7780 ;
        RECT 7.2320 25.6240 7.2500 26.7830 ;
        RECT 0.1220 25.6235 0.1400 26.7835 ;
        RECT 16.3940 26.7035 16.4120 27.8635 ;
        RECT 9.2840 26.7040 9.3020 27.8630 ;
        RECT 7.8800 26.7440 7.9700 27.8580 ;
        RECT 7.2320 26.7040 7.2500 27.8630 ;
        RECT 0.1220 26.7035 0.1400 27.8635 ;
      LAYER V3  ;
        RECT 0.1220 1.1720 0.1400 1.2200 ;
        RECT 7.2320 1.1720 7.2500 1.2200 ;
        RECT 7.8800 1.1720 7.9700 1.2200 ;
        RECT 9.2840 1.1720 9.3020 1.2200 ;
        RECT 16.3940 1.1720 16.4120 1.2200 ;
        RECT 0.1220 2.2520 0.1400 2.3000 ;
        RECT 7.2320 2.2520 7.2500 2.3000 ;
        RECT 7.8800 2.2520 7.9700 2.3000 ;
        RECT 9.2840 2.2520 9.3020 2.3000 ;
        RECT 16.3940 2.2520 16.4120 2.3000 ;
        RECT 0.1220 3.3320 0.1400 3.3800 ;
        RECT 7.2320 3.3320 7.2500 3.3800 ;
        RECT 7.8800 3.3320 7.9700 3.3800 ;
        RECT 9.2840 3.3320 9.3020 3.3800 ;
        RECT 16.3940 3.3320 16.4120 3.3800 ;
        RECT 0.1220 4.4120 0.1400 4.4600 ;
        RECT 7.2320 4.4120 7.2500 4.4600 ;
        RECT 7.8800 4.4120 7.9700 4.4600 ;
        RECT 9.2840 4.4120 9.3020 4.4600 ;
        RECT 16.3940 4.4120 16.4120 4.4600 ;
        RECT 0.1220 5.4920 0.1400 5.5400 ;
        RECT 7.2320 5.4920 7.2500 5.5400 ;
        RECT 7.8800 5.4920 7.9700 5.5400 ;
        RECT 9.2840 5.4920 9.3020 5.5400 ;
        RECT 16.3940 5.4920 16.4120 5.5400 ;
        RECT 0.1220 6.5720 0.1400 6.6200 ;
        RECT 7.2320 6.5720 7.2500 6.6200 ;
        RECT 7.8800 6.5720 7.9700 6.6200 ;
        RECT 9.2840 6.5720 9.3020 6.6200 ;
        RECT 16.3940 6.5720 16.4120 6.6200 ;
        RECT 0.1220 7.6520 0.1400 7.7000 ;
        RECT 7.2320 7.6520 7.2500 7.7000 ;
        RECT 7.8800 7.6520 7.9700 7.7000 ;
        RECT 9.2840 7.6520 9.3020 7.7000 ;
        RECT 16.3940 7.6520 16.4120 7.7000 ;
        RECT 0.1220 8.7320 0.1400 8.7800 ;
        RECT 7.2320 8.7320 7.2500 8.7800 ;
        RECT 7.8800 8.7320 7.9700 8.7800 ;
        RECT 9.2840 8.7320 9.3020 8.7800 ;
        RECT 16.3940 8.7320 16.4120 8.7800 ;
        RECT 0.1220 9.8120 0.1400 9.8600 ;
        RECT 7.2320 9.8120 7.2500 9.8600 ;
        RECT 7.8800 9.8120 7.9700 9.8600 ;
        RECT 9.2840 9.8120 9.3020 9.8600 ;
        RECT 16.3940 9.8120 16.4120 9.8600 ;
        RECT 7.9150 16.6290 7.9330 16.8450 ;
        RECT 7.9150 13.4610 7.9330 13.6770 ;
        RECT 7.9150 10.2930 7.9330 10.5090 ;
        RECT 7.9670 16.6290 7.9850 16.8450 ;
        RECT 7.9670 13.4610 7.9850 13.6770 ;
        RECT 7.9670 10.2930 7.9850 10.5090 ;
        RECT 8.0190 16.6290 8.0370 16.8450 ;
        RECT 8.0190 13.4610 8.0370 13.6770 ;
        RECT 8.0190 10.2930 8.0370 10.5090 ;
        RECT 8.0710 16.6290 8.0890 16.8450 ;
        RECT 8.0710 13.4610 8.0890 13.6770 ;
        RECT 8.0710 10.2930 8.0890 10.5090 ;
        RECT 8.1230 16.6290 8.1410 16.8450 ;
        RECT 8.1230 13.4610 8.1410 13.6770 ;
        RECT 8.1230 10.2930 8.1410 10.5090 ;
        RECT 9.2790 10.0130 9.2970 10.0370 ;
        RECT 9.2970 13.7970 9.3150 13.8210 ;
        RECT 0.1220 19.0190 0.1400 19.0670 ;
        RECT 7.2320 19.0190 7.2500 19.0670 ;
        RECT 7.8800 19.0190 7.9700 19.0670 ;
        RECT 9.2840 19.0190 9.3020 19.0670 ;
        RECT 16.3940 19.0190 16.4120 19.0670 ;
        RECT 0.1220 20.0990 0.1400 20.1470 ;
        RECT 7.2320 20.0990 7.2500 20.1470 ;
        RECT 7.8800 20.0990 7.9700 20.1470 ;
        RECT 9.2840 20.0990 9.3020 20.1470 ;
        RECT 16.3940 20.0990 16.4120 20.1470 ;
        RECT 0.1220 21.1790 0.1400 21.2270 ;
        RECT 7.2320 21.1790 7.2500 21.2270 ;
        RECT 7.8800 21.1790 7.9700 21.2270 ;
        RECT 9.2840 21.1790 9.3020 21.2270 ;
        RECT 16.3940 21.1790 16.4120 21.2270 ;
        RECT 0.1220 22.2590 0.1400 22.3070 ;
        RECT 7.2320 22.2590 7.2500 22.3070 ;
        RECT 7.8800 22.2590 7.9700 22.3070 ;
        RECT 9.2840 22.2590 9.3020 22.3070 ;
        RECT 16.3940 22.2590 16.4120 22.3070 ;
        RECT 0.1220 23.3390 0.1400 23.3870 ;
        RECT 7.2320 23.3390 7.2500 23.3870 ;
        RECT 7.8800 23.3390 7.9700 23.3870 ;
        RECT 9.2840 23.3390 9.3020 23.3870 ;
        RECT 16.3940 23.3390 16.4120 23.3870 ;
        RECT 0.1220 24.4190 0.1400 24.4670 ;
        RECT 7.2320 24.4190 7.2500 24.4670 ;
        RECT 7.8800 24.4190 7.9700 24.4670 ;
        RECT 9.2840 24.4190 9.3020 24.4670 ;
        RECT 16.3940 24.4190 16.4120 24.4670 ;
        RECT 0.1220 25.4990 0.1400 25.5470 ;
        RECT 7.2320 25.4990 7.2500 25.5470 ;
        RECT 7.8800 25.4990 7.9700 25.5470 ;
        RECT 9.2840 25.4990 9.3020 25.5470 ;
        RECT 16.3940 25.4990 16.4120 25.5470 ;
        RECT 0.1220 26.5790 0.1400 26.6270 ;
        RECT 7.2320 26.5790 7.2500 26.6270 ;
        RECT 7.8800 26.5790 7.9700 26.6270 ;
        RECT 9.2840 26.5790 9.3020 26.6270 ;
        RECT 16.3940 26.5790 16.4120 26.6270 ;
        RECT 0.1220 27.6590 0.1400 27.7070 ;
        RECT 7.2320 27.6590 7.2500 27.7070 ;
        RECT 7.8800 27.6590 7.9700 27.7070 ;
        RECT 9.2840 27.6590 9.3020 27.7070 ;
        RECT 16.3940 27.6590 16.4120 27.7070 ;
      LAYER M5  ;
        RECT 9.2160 9.9950 9.2400 13.8390 ;
      LAYER V4  ;
        RECT 9.2160 13.7970 9.2400 13.8210 ;
        RECT 9.2160 10.2930 9.2400 10.5090 ;
        RECT 9.2160 10.0130 9.2400 10.0370 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.0760 16.4370 1.1240 ;
        RECT 0.0940 2.1560 16.4370 2.2040 ;
        RECT 0.0940 3.2360 16.4370 3.2840 ;
        RECT 0.0940 4.3160 16.4370 4.3640 ;
        RECT 0.0940 5.3960 16.4370 5.4440 ;
        RECT 0.0940 6.4760 16.4370 6.5240 ;
        RECT 0.0940 7.5560 16.4370 7.6040 ;
        RECT 0.0940 8.6360 16.4370 8.6840 ;
        RECT 0.0940 9.7160 16.4370 9.7640 ;
        RECT 3.5640 10.7250 12.9600 10.9410 ;
        RECT 7.3980 13.8930 9.1260 14.1090 ;
        RECT 7.3980 17.0610 9.1260 17.2770 ;
        RECT 0.0940 18.9230 16.4370 18.9710 ;
        RECT 0.0940 20.0030 16.4370 20.0510 ;
        RECT 0.0940 21.0830 16.4370 21.1310 ;
        RECT 0.0940 22.1630 16.4370 22.2110 ;
        RECT 0.0940 23.2430 16.4370 23.2910 ;
        RECT 0.0940 24.3230 16.4370 24.3710 ;
        RECT 0.0940 25.4030 16.4370 25.4510 ;
        RECT 0.0940 26.4830 16.4370 26.5310 ;
        RECT 0.0940 27.5630 16.4370 27.6110 ;
      LAYER M3  ;
        RECT 16.3580 0.2165 16.3760 1.3765 ;
        RECT 9.3380 0.2165 9.3560 1.3765 ;
        RECT 8.5730 0.2530 8.6090 1.3670 ;
        RECT 8.4200 0.2530 8.4470 1.3670 ;
        RECT 7.1780 0.2165 7.1960 1.3765 ;
        RECT 0.1580 0.2165 0.1760 1.3765 ;
        RECT 16.3580 1.2965 16.3760 2.4565 ;
        RECT 9.3380 1.2965 9.3560 2.4565 ;
        RECT 8.5730 1.3330 8.6090 2.4470 ;
        RECT 8.4200 1.3330 8.4470 2.4470 ;
        RECT 7.1780 1.2965 7.1960 2.4565 ;
        RECT 0.1580 1.2965 0.1760 2.4565 ;
        RECT 16.3580 2.3765 16.3760 3.5365 ;
        RECT 9.3380 2.3765 9.3560 3.5365 ;
        RECT 8.5730 2.4130 8.6090 3.5270 ;
        RECT 8.4200 2.4130 8.4470 3.5270 ;
        RECT 7.1780 2.3765 7.1960 3.5365 ;
        RECT 0.1580 2.3765 0.1760 3.5365 ;
        RECT 16.3580 3.4565 16.3760 4.6165 ;
        RECT 9.3380 3.4565 9.3560 4.6165 ;
        RECT 8.5730 3.4930 8.6090 4.6070 ;
        RECT 8.4200 3.4930 8.4470 4.6070 ;
        RECT 7.1780 3.4565 7.1960 4.6165 ;
        RECT 0.1580 3.4565 0.1760 4.6165 ;
        RECT 16.3580 4.5365 16.3760 5.6965 ;
        RECT 9.3380 4.5365 9.3560 5.6965 ;
        RECT 8.5730 4.5730 8.6090 5.6870 ;
        RECT 8.4200 4.5730 8.4470 5.6870 ;
        RECT 7.1780 4.5365 7.1960 5.6965 ;
        RECT 0.1580 4.5365 0.1760 5.6965 ;
        RECT 16.3580 5.6165 16.3760 6.7765 ;
        RECT 9.3380 5.6165 9.3560 6.7765 ;
        RECT 8.5730 5.6530 8.6090 6.7670 ;
        RECT 8.4200 5.6530 8.4470 6.7670 ;
        RECT 7.1780 5.6165 7.1960 6.7765 ;
        RECT 0.1580 5.6165 0.1760 6.7765 ;
        RECT 16.3580 6.6965 16.3760 7.8565 ;
        RECT 9.3380 6.6965 9.3560 7.8565 ;
        RECT 8.5730 6.7330 8.6090 7.8470 ;
        RECT 8.4200 6.7330 8.4470 7.8470 ;
        RECT 7.1780 6.6965 7.1960 7.8565 ;
        RECT 0.1580 6.6965 0.1760 7.8565 ;
        RECT 16.3580 7.7765 16.3760 8.9365 ;
        RECT 9.3380 7.7765 9.3560 8.9365 ;
        RECT 8.5730 7.8130 8.6090 8.9270 ;
        RECT 8.4200 7.8130 8.4470 8.9270 ;
        RECT 7.1780 7.7765 7.1960 8.9365 ;
        RECT 0.1580 7.7765 0.1760 8.9365 ;
        RECT 16.3580 8.8565 16.3760 10.0165 ;
        RECT 9.3380 8.8565 9.3560 10.0165 ;
        RECT 8.5730 8.8930 8.6090 10.0070 ;
        RECT 8.4200 8.8930 8.4470 10.0070 ;
        RECT 7.1780 8.8565 7.1960 10.0165 ;
        RECT 0.1580 8.8565 0.1760 10.0165 ;
        RECT 16.3530 9.9305 16.3710 18.1375 ;
        RECT 9.3330 9.9305 9.3510 18.1375 ;
        RECT 8.3790 10.1540 8.6130 17.8370 ;
        RECT 8.5680 9.9745 8.6040 18.0940 ;
        RECT 8.4150 9.9740 8.4420 18.0940 ;
        RECT 7.1730 9.9305 7.1910 18.1375 ;
        RECT 0.1530 9.9305 0.1710 18.1375 ;
        RECT 16.3580 18.0635 16.3760 19.2235 ;
        RECT 9.3380 18.0635 9.3560 19.2235 ;
        RECT 8.5730 18.1000 8.6090 19.2140 ;
        RECT 8.4200 18.1000 8.4470 19.2140 ;
        RECT 7.1780 18.0635 7.1960 19.2235 ;
        RECT 0.1580 18.0635 0.1760 19.2235 ;
        RECT 16.3580 19.1435 16.3760 20.3035 ;
        RECT 9.3380 19.1435 9.3560 20.3035 ;
        RECT 8.5730 19.1800 8.6090 20.2940 ;
        RECT 8.4200 19.1800 8.4470 20.2940 ;
        RECT 7.1780 19.1435 7.1960 20.3035 ;
        RECT 0.1580 19.1435 0.1760 20.3035 ;
        RECT 16.3580 20.2235 16.3760 21.3835 ;
        RECT 9.3380 20.2235 9.3560 21.3835 ;
        RECT 8.5730 20.2600 8.6090 21.3740 ;
        RECT 8.4200 20.2600 8.4470 21.3740 ;
        RECT 7.1780 20.2235 7.1960 21.3835 ;
        RECT 0.1580 20.2235 0.1760 21.3835 ;
        RECT 16.3580 21.3035 16.3760 22.4635 ;
        RECT 9.3380 21.3035 9.3560 22.4635 ;
        RECT 8.5730 21.3400 8.6090 22.4540 ;
        RECT 8.4200 21.3400 8.4470 22.4540 ;
        RECT 7.1780 21.3035 7.1960 22.4635 ;
        RECT 0.1580 21.3035 0.1760 22.4635 ;
        RECT 16.3580 22.3835 16.3760 23.5435 ;
        RECT 9.3380 22.3835 9.3560 23.5435 ;
        RECT 8.5730 22.4200 8.6090 23.5340 ;
        RECT 8.4200 22.4200 8.4470 23.5340 ;
        RECT 7.1780 22.3835 7.1960 23.5435 ;
        RECT 0.1580 22.3835 0.1760 23.5435 ;
        RECT 16.3580 23.4635 16.3760 24.6235 ;
        RECT 9.3380 23.4635 9.3560 24.6235 ;
        RECT 8.5730 23.5000 8.6090 24.6140 ;
        RECT 8.4200 23.5000 8.4470 24.6140 ;
        RECT 7.1780 23.4635 7.1960 24.6235 ;
        RECT 0.1580 23.4635 0.1760 24.6235 ;
        RECT 16.3580 24.5435 16.3760 25.7035 ;
        RECT 9.3380 24.5435 9.3560 25.7035 ;
        RECT 8.5730 24.5800 8.6090 25.6940 ;
        RECT 8.4200 24.5800 8.4470 25.6940 ;
        RECT 7.1780 24.5435 7.1960 25.7035 ;
        RECT 0.1580 24.5435 0.1760 25.7035 ;
        RECT 16.3580 25.6235 16.3760 26.7835 ;
        RECT 9.3380 25.6235 9.3560 26.7835 ;
        RECT 8.5730 25.6600 8.6090 26.7740 ;
        RECT 8.4200 25.6600 8.4470 26.7740 ;
        RECT 7.1780 25.6235 7.1960 26.7835 ;
        RECT 0.1580 25.6235 0.1760 26.7835 ;
        RECT 16.3580 26.7035 16.3760 27.8635 ;
        RECT 9.3380 26.7035 9.3560 27.8635 ;
        RECT 8.5730 26.7400 8.6090 27.8540 ;
        RECT 8.4200 26.7400 8.4470 27.8540 ;
        RECT 7.1780 26.7035 7.1960 27.8635 ;
        RECT 0.1580 26.7035 0.1760 27.8635 ;
      LAYER V3  ;
        RECT 0.1580 1.0760 0.1760 1.1240 ;
        RECT 7.1780 1.0760 7.1960 1.1240 ;
        RECT 8.4200 1.0760 8.4470 1.1240 ;
        RECT 8.5730 1.0760 8.6090 1.1240 ;
        RECT 9.3380 1.0760 9.3560 1.1240 ;
        RECT 16.3580 1.0760 16.3760 1.1240 ;
        RECT 0.1580 2.1560 0.1760 2.2040 ;
        RECT 7.1780 2.1560 7.1960 2.2040 ;
        RECT 8.4200 2.1560 8.4470 2.2040 ;
        RECT 8.5730 2.1560 8.6090 2.2040 ;
        RECT 9.3380 2.1560 9.3560 2.2040 ;
        RECT 16.3580 2.1560 16.3760 2.2040 ;
        RECT 0.1580 3.2360 0.1760 3.2840 ;
        RECT 7.1780 3.2360 7.1960 3.2840 ;
        RECT 8.4200 3.2360 8.4470 3.2840 ;
        RECT 8.5730 3.2360 8.6090 3.2840 ;
        RECT 9.3380 3.2360 9.3560 3.2840 ;
        RECT 16.3580 3.2360 16.3760 3.2840 ;
        RECT 0.1580 4.3160 0.1760 4.3640 ;
        RECT 7.1780 4.3160 7.1960 4.3640 ;
        RECT 8.4200 4.3160 8.4470 4.3640 ;
        RECT 8.5730 4.3160 8.6090 4.3640 ;
        RECT 9.3380 4.3160 9.3560 4.3640 ;
        RECT 16.3580 4.3160 16.3760 4.3640 ;
        RECT 0.1580 5.3960 0.1760 5.4440 ;
        RECT 7.1780 5.3960 7.1960 5.4440 ;
        RECT 8.4200 5.3960 8.4470 5.4440 ;
        RECT 8.5730 5.3960 8.6090 5.4440 ;
        RECT 9.3380 5.3960 9.3560 5.4440 ;
        RECT 16.3580 5.3960 16.3760 5.4440 ;
        RECT 0.1580 6.4760 0.1760 6.5240 ;
        RECT 7.1780 6.4760 7.1960 6.5240 ;
        RECT 8.4200 6.4760 8.4470 6.5240 ;
        RECT 8.5730 6.4760 8.6090 6.5240 ;
        RECT 9.3380 6.4760 9.3560 6.5240 ;
        RECT 16.3580 6.4760 16.3760 6.5240 ;
        RECT 0.1580 7.5560 0.1760 7.6040 ;
        RECT 7.1780 7.5560 7.1960 7.6040 ;
        RECT 8.4200 7.5560 8.4470 7.6040 ;
        RECT 8.5730 7.5560 8.6090 7.6040 ;
        RECT 9.3380 7.5560 9.3560 7.6040 ;
        RECT 16.3580 7.5560 16.3760 7.6040 ;
        RECT 0.1580 8.6360 0.1760 8.6840 ;
        RECT 7.1780 8.6360 7.1960 8.6840 ;
        RECT 8.4200 8.6360 8.4470 8.6840 ;
        RECT 8.5730 8.6360 8.6090 8.6840 ;
        RECT 9.3380 8.6360 9.3560 8.6840 ;
        RECT 16.3580 8.6360 16.3760 8.6840 ;
        RECT 0.1580 9.7160 0.1760 9.7640 ;
        RECT 7.1780 9.7160 7.1960 9.7640 ;
        RECT 8.4200 9.7160 8.4470 9.7640 ;
        RECT 8.5730 9.7160 8.6090 9.7640 ;
        RECT 9.3380 9.7160 9.3560 9.7640 ;
        RECT 16.3580 9.7160 16.3760 9.7640 ;
        RECT 8.3830 17.0610 8.4010 17.2770 ;
        RECT 8.3830 13.8930 8.4010 14.1090 ;
        RECT 8.3830 10.7250 8.4010 10.9410 ;
        RECT 8.4350 17.0610 8.4530 17.2770 ;
        RECT 8.4350 13.8930 8.4530 14.1090 ;
        RECT 8.4350 10.7250 8.4530 10.9410 ;
        RECT 8.4870 17.0610 8.5050 17.2770 ;
        RECT 8.4870 13.8930 8.5050 14.1090 ;
        RECT 8.4870 10.7250 8.5050 10.9410 ;
        RECT 8.5390 17.0610 8.5570 17.2770 ;
        RECT 8.5390 13.8930 8.5570 14.1090 ;
        RECT 8.5390 10.7250 8.5570 10.9410 ;
        RECT 8.5910 17.0610 8.6090 17.2770 ;
        RECT 8.5910 13.8930 8.6090 14.1090 ;
        RECT 8.5910 10.7250 8.6090 10.9410 ;
        RECT 9.3330 10.7255 9.3510 10.9415 ;
        RECT 0.1580 18.9230 0.1760 18.9710 ;
        RECT 7.1780 18.9230 7.1960 18.9710 ;
        RECT 8.4200 18.9230 8.4470 18.9710 ;
        RECT 8.5730 18.9230 8.6090 18.9710 ;
        RECT 9.3380 18.9230 9.3560 18.9710 ;
        RECT 16.3580 18.9230 16.3760 18.9710 ;
        RECT 0.1580 20.0030 0.1760 20.0510 ;
        RECT 7.1780 20.0030 7.1960 20.0510 ;
        RECT 8.4200 20.0030 8.4470 20.0510 ;
        RECT 8.5730 20.0030 8.6090 20.0510 ;
        RECT 9.3380 20.0030 9.3560 20.0510 ;
        RECT 16.3580 20.0030 16.3760 20.0510 ;
        RECT 0.1580 21.0830 0.1760 21.1310 ;
        RECT 7.1780 21.0830 7.1960 21.1310 ;
        RECT 8.4200 21.0830 8.4470 21.1310 ;
        RECT 8.5730 21.0830 8.6090 21.1310 ;
        RECT 9.3380 21.0830 9.3560 21.1310 ;
        RECT 16.3580 21.0830 16.3760 21.1310 ;
        RECT 0.1580 22.1630 0.1760 22.2110 ;
        RECT 7.1780 22.1630 7.1960 22.2110 ;
        RECT 8.4200 22.1630 8.4470 22.2110 ;
        RECT 8.5730 22.1630 8.6090 22.2110 ;
        RECT 9.3380 22.1630 9.3560 22.2110 ;
        RECT 16.3580 22.1630 16.3760 22.2110 ;
        RECT 0.1580 23.2430 0.1760 23.2910 ;
        RECT 7.1780 23.2430 7.1960 23.2910 ;
        RECT 8.4200 23.2430 8.4470 23.2910 ;
        RECT 8.5730 23.2430 8.6090 23.2910 ;
        RECT 9.3380 23.2430 9.3560 23.2910 ;
        RECT 16.3580 23.2430 16.3760 23.2910 ;
        RECT 0.1580 24.3230 0.1760 24.3710 ;
        RECT 7.1780 24.3230 7.1960 24.3710 ;
        RECT 8.4200 24.3230 8.4470 24.3710 ;
        RECT 8.5730 24.3230 8.6090 24.3710 ;
        RECT 9.3380 24.3230 9.3560 24.3710 ;
        RECT 16.3580 24.3230 16.3760 24.3710 ;
        RECT 0.1580 25.4030 0.1760 25.4510 ;
        RECT 7.1780 25.4030 7.1960 25.4510 ;
        RECT 8.4200 25.4030 8.4470 25.4510 ;
        RECT 8.5730 25.4030 8.6090 25.4510 ;
        RECT 9.3380 25.4030 9.3560 25.4510 ;
        RECT 16.3580 25.4030 16.3760 25.4510 ;
        RECT 0.1580 26.4830 0.1760 26.5310 ;
        RECT 7.1780 26.4830 7.1960 26.5310 ;
        RECT 8.4200 26.4830 8.4470 26.5310 ;
        RECT 8.5730 26.4830 8.6090 26.5310 ;
        RECT 9.3380 26.4830 9.3560 26.5310 ;
        RECT 16.3580 26.4830 16.3760 26.5310 ;
        RECT 0.1580 27.5630 0.1760 27.6110 ;
        RECT 7.1780 27.5630 7.1960 27.6110 ;
        RECT 8.4200 27.5630 8.4470 27.6110 ;
        RECT 8.5730 27.5630 8.6090 27.6110 ;
        RECT 9.3380 27.5630 9.3560 27.6110 ;
        RECT 16.3580 27.5630 16.3760 27.6110 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.7910 11.1970 10.8090 11.2340 ;
      LAYER M4  ;
        RECT 10.7390 11.2050 10.8230 11.2290 ;
      LAYER M5  ;
        RECT 10.7880 10.2540 10.8120 13.4940 ;
      LAYER V3  ;
        RECT 10.7910 11.2050 10.8090 11.2290 ;
      LAYER V4  ;
        RECT 10.7880 11.2050 10.8120 11.2290 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.5750 11.2000 10.5930 11.2370 ;
      LAYER M4  ;
        RECT 10.5230 11.2050 10.6070 11.2290 ;
      LAYER M5  ;
        RECT 10.5720 10.2540 10.5960 13.4940 ;
      LAYER V3  ;
        RECT 10.5750 11.2050 10.5930 11.2290 ;
      LAYER V4  ;
        RECT 10.5720 11.2050 10.5960 11.2290 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.3590 10.6210 10.3770 10.6580 ;
      LAYER M4  ;
        RECT 10.3070 10.6290 10.3910 10.6530 ;
      LAYER M5  ;
        RECT 10.3560 10.2540 10.3800 13.4940 ;
      LAYER V3  ;
        RECT 10.3590 10.6290 10.3770 10.6530 ;
      LAYER V4  ;
        RECT 10.3560 10.6290 10.3800 10.6530 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.1430 10.8610 10.1610 11.0420 ;
      LAYER M4  ;
        RECT 10.0910 11.0130 10.1750 11.0370 ;
      LAYER M5  ;
        RECT 10.1400 10.2540 10.1640 13.4940 ;
      LAYER V3  ;
        RECT 10.1430 11.0130 10.1610 11.0370 ;
      LAYER V4  ;
        RECT 10.1400 11.0130 10.1640 11.0370 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.9270 10.6240 9.9450 10.6910 ;
      LAYER M4  ;
        RECT 9.8750 10.6290 9.9590 10.6530 ;
      LAYER M5  ;
        RECT 9.9240 10.2540 9.9480 13.4940 ;
      LAYER V3  ;
        RECT 9.9270 10.6290 9.9450 10.6530 ;
      LAYER V4  ;
        RECT 9.9240 10.6290 9.9480 10.6530 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.7110 10.3570 9.7290 10.6100 ;
      LAYER M4  ;
        RECT 9.6590 10.5810 9.7430 10.6050 ;
      LAYER M5  ;
        RECT 9.7080 10.2540 9.7320 13.4940 ;
      LAYER V3  ;
        RECT 9.7110 10.5810 9.7290 10.6050 ;
      LAYER V4  ;
        RECT 9.7080 10.5810 9.7320 10.6050 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.4950 11.3920 9.5130 11.4290 ;
      LAYER M4  ;
        RECT 9.4430 11.3970 9.5270 11.4210 ;
      LAYER M5  ;
        RECT 9.4920 10.2540 9.5160 13.4940 ;
      LAYER V3  ;
        RECT 9.4950 11.3970 9.5130 11.4210 ;
      LAYER V4  ;
        RECT 9.4920 11.3970 9.5160 11.4210 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.2790 11.2390 9.2970 11.3300 ;
      LAYER M4  ;
        RECT 9.2270 11.3010 9.3110 11.3250 ;
      LAYER M5  ;
        RECT 9.2760 10.2540 9.3000 13.4940 ;
      LAYER V3  ;
        RECT 9.2790 11.3010 9.2970 11.3250 ;
      LAYER V4  ;
        RECT 9.2760 11.3010 9.3000 11.3250 ;
    END
  END ADDRESS[7]
  PIN ADDRESS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.6310 10.6240 8.6490 10.6910 ;
      LAYER M4  ;
        RECT 8.3470 10.6290 8.6600 10.6530 ;
      LAYER M5  ;
        RECT 8.3580 10.2540 8.3820 13.4940 ;
      LAYER V3  ;
        RECT 8.6310 10.6290 8.6490 10.6530 ;
      LAYER V4  ;
        RECT 8.3580 10.6290 8.3820 10.6530 ;
    END
  END ADDRESS[8]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.2350 10.3570 8.2530 10.6100 ;
      LAYER M4  ;
        RECT 8.0230 10.5810 8.2640 10.6050 ;
      LAYER M5  ;
        RECT 8.0340 10.2540 8.0580 13.4940 ;
      LAYER V3  ;
        RECT 8.2350 10.5810 8.2530 10.6050 ;
      LAYER V4  ;
        RECT 8.0340 10.5810 8.0580 10.6050 ;
    END
  END banksel
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.4430 10.6240 7.4610 10.6910 ;
      LAYER M4  ;
        RECT 7.3910 10.6290 7.4750 10.6530 ;
      LAYER M5  ;
        RECT 7.4400 10.2540 7.4640 13.4940 ;
      LAYER V3  ;
        RECT 7.4430 10.6290 7.4610 10.6530 ;
      LAYER V4  ;
        RECT 7.4400 10.6290 7.4640 10.6530 ;
    END
  END write
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2270 11.4880 7.2450 11.5370 ;
      LAYER M4  ;
        RECT 7.1750 11.4930 7.2590 11.5170 ;
      LAYER M5  ;
        RECT 7.2240 10.2540 7.2480 13.4940 ;
      LAYER V3  ;
        RECT 7.2270 11.4930 7.2450 11.5170 ;
      LAYER V4  ;
        RECT 7.2240 11.4930 7.2480 11.5170 ;
    END
  END clk
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2630 10.3570 7.2810 10.6100 ;
      LAYER M4  ;
        RECT 6.9970 10.5810 7.2920 10.6050 ;
      LAYER M5  ;
        RECT 7.0080 10.2540 7.0320 13.4940 ;
      LAYER V3  ;
        RECT 7.2630 10.5810 7.2810 10.6050 ;
      LAYER V4  ;
        RECT 7.0080 10.5810 7.0320 10.6050 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.7950 11.1970 6.8130 11.2340 ;
      LAYER M4  ;
        RECT 6.7430 11.2050 6.8270 11.2290 ;
      LAYER M5  ;
        RECT 6.7920 10.2540 6.8160 13.4940 ;
      LAYER V3  ;
        RECT 6.7950 11.2050 6.8130 11.2290 ;
      LAYER V4  ;
        RECT 6.7920 11.2050 6.8160 11.2290 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.5790 10.6240 6.5970 10.8530 ;
      LAYER M4  ;
        RECT 6.5270 10.6290 6.6110 10.6530 ;
      LAYER M5  ;
        RECT 6.5760 10.2540 6.6000 13.4940 ;
      LAYER V3  ;
        RECT 6.5790 10.6290 6.5970 10.6530 ;
      LAYER V4  ;
        RECT 6.5760 10.6290 6.6000 10.6530 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.3630 10.3570 6.3810 10.6100 ;
      LAYER M4  ;
        RECT 6.3110 10.5810 6.3950 10.6050 ;
      LAYER M5  ;
        RECT 6.3600 10.2540 6.3840 13.4940 ;
      LAYER V3  ;
        RECT 6.3630 10.5810 6.3810 10.6050 ;
      LAYER V4  ;
        RECT 6.3600 10.5810 6.3840 10.6050 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.1470 10.6210 6.1650 10.6580 ;
      LAYER M4  ;
        RECT 6.0950 10.6290 6.1790 10.6530 ;
      LAYER M5  ;
        RECT 6.1440 10.2540 6.1680 13.4940 ;
      LAYER V3  ;
        RECT 6.1470 10.6290 6.1650 10.6530 ;
      LAYER V4  ;
        RECT 6.1440 10.6290 6.1680 10.6530 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 5.9310 11.1970 5.9490 11.2340 ;
      LAYER M4  ;
        RECT 5.8790 11.2050 5.9630 11.2290 ;
      LAYER M5  ;
        RECT 5.9280 10.2540 5.9520 13.4940 ;
      LAYER V3  ;
        RECT 5.9310 11.2050 5.9490 11.2290 ;
      LAYER V4  ;
        RECT 5.9280 11.2050 5.9520 11.2290 ;
    END
  END sdel[4]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.4280 8.5970 0.4520 ;
      LAYER M3  ;
        RECT 8.5370 0.3775 8.5550 0.6170 ;
      LAYER V3  ;
        RECT 8.5370 0.4280 8.5550 0.4520 ;
    END
  END dataout[0]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.3320 8.6650 0.3560 ;
      LAYER M3  ;
        RECT 8.3120 0.2700 8.3300 0.6750 ;
      LAYER V3  ;
        RECT 8.3120 0.3320 8.3300 0.3560 ;
    END
  END wd[0]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.5080 8.5970 1.5320 ;
      LAYER M3  ;
        RECT 8.5370 1.4575 8.5550 1.6970 ;
      LAYER V3  ;
        RECT 8.5370 1.5080 8.5550 1.5320 ;
    END
  END dataout[1]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.4120 8.6650 1.4360 ;
      LAYER M3  ;
        RECT 8.3120 1.3500 8.3300 1.7550 ;
      LAYER V3  ;
        RECT 8.3120 1.4120 8.3300 1.4360 ;
    END
  END wd[1]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.5880 8.5970 2.6120 ;
      LAYER M3  ;
        RECT 8.5370 2.5375 8.5550 2.7770 ;
      LAYER V3  ;
        RECT 8.5370 2.5880 8.5550 2.6120 ;
    END
  END dataout[2]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.4920 8.6650 2.5160 ;
      LAYER M3  ;
        RECT 8.3120 2.4300 8.3300 2.8350 ;
      LAYER V3  ;
        RECT 8.3120 2.4920 8.3300 2.5160 ;
    END
  END wd[2]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.6680 8.5970 3.6920 ;
      LAYER M3  ;
        RECT 8.5370 3.6175 8.5550 3.8570 ;
      LAYER V3  ;
        RECT 8.5370 3.6680 8.5550 3.6920 ;
    END
  END dataout[3]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.5720 8.6650 3.5960 ;
      LAYER M3  ;
        RECT 8.3120 3.5100 8.3300 3.9150 ;
      LAYER V3  ;
        RECT 8.3120 3.5720 8.3300 3.5960 ;
    END
  END wd[3]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.7480 8.5970 4.7720 ;
      LAYER M3  ;
        RECT 8.5370 4.6975 8.5550 4.9370 ;
      LAYER V3  ;
        RECT 8.5370 4.7480 8.5550 4.7720 ;
    END
  END dataout[4]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.6520 8.6650 4.6760 ;
      LAYER M3  ;
        RECT 8.3120 4.5900 8.3300 4.9950 ;
      LAYER V3  ;
        RECT 8.3120 4.6520 8.3300 4.6760 ;
    END
  END wd[4]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.8280 8.5970 5.8520 ;
      LAYER M3  ;
        RECT 8.5370 5.7775 8.5550 6.0170 ;
      LAYER V3  ;
        RECT 8.5370 5.8280 8.5550 5.8520 ;
    END
  END dataout[5]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.7320 8.6650 5.7560 ;
      LAYER M3  ;
        RECT 8.3120 5.6700 8.3300 6.0750 ;
      LAYER V3  ;
        RECT 8.3120 5.7320 8.3300 5.7560 ;
    END
  END wd[5]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.9080 8.5970 6.9320 ;
      LAYER M3  ;
        RECT 8.5370 6.8575 8.5550 7.0970 ;
      LAYER V3  ;
        RECT 8.5370 6.9080 8.5550 6.9320 ;
    END
  END dataout[6]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.8120 8.6650 6.8360 ;
      LAYER M3  ;
        RECT 8.3120 6.7500 8.3300 7.1550 ;
      LAYER V3  ;
        RECT 8.3120 6.8120 8.3300 6.8360 ;
    END
  END wd[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.9880 8.5970 8.0120 ;
      LAYER M3  ;
        RECT 8.5370 7.9375 8.5550 8.1770 ;
      LAYER V3  ;
        RECT 8.5370 7.9880 8.5550 8.0120 ;
    END
  END dataout[7]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.8920 8.6650 7.9160 ;
      LAYER M3  ;
        RECT 8.3120 7.8300 8.3300 8.2350 ;
      LAYER V3  ;
        RECT 8.3120 7.8920 8.3300 7.9160 ;
    END
  END wd[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 9.0680 8.5970 9.0920 ;
      LAYER M3  ;
        RECT 8.5370 9.0175 8.5550 9.2570 ;
      LAYER V3  ;
        RECT 8.5370 9.0680 8.5550 9.0920 ;
    END
  END dataout[8]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 8.9720 8.6650 8.9960 ;
      LAYER M3  ;
        RECT 8.3120 8.9100 8.3300 9.3150 ;
      LAYER V3  ;
        RECT 8.3120 8.9720 8.3300 8.9960 ;
    END
  END wd[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 18.2750 8.5970 18.2990 ;
      LAYER M3  ;
        RECT 8.5370 18.2245 8.5550 18.4640 ;
      LAYER V3  ;
        RECT 8.5370 18.2750 8.5550 18.2990 ;
    END
  END dataout[9]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 18.1790 8.6650 18.2030 ;
      LAYER M3  ;
        RECT 8.3120 18.1170 8.3300 18.5220 ;
      LAYER V3  ;
        RECT 8.3120 18.1790 8.3300 18.2030 ;
    END
  END wd[9]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.3550 8.5970 19.3790 ;
      LAYER M3  ;
        RECT 8.5370 19.3045 8.5550 19.5440 ;
      LAYER V3  ;
        RECT 8.5370 19.3550 8.5550 19.3790 ;
    END
  END dataout[10]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.2590 8.6650 19.2830 ;
      LAYER M3  ;
        RECT 8.3120 19.1970 8.3300 19.6020 ;
      LAYER V3  ;
        RECT 8.3120 19.2590 8.3300 19.2830 ;
    END
  END wd[10]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.4350 8.5970 20.4590 ;
      LAYER M3  ;
        RECT 8.5370 20.3845 8.5550 20.6240 ;
      LAYER V3  ;
        RECT 8.5370 20.4350 8.5550 20.4590 ;
    END
  END dataout[11]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.3390 8.6650 20.3630 ;
      LAYER M3  ;
        RECT 8.3120 20.2770 8.3300 20.6820 ;
      LAYER V3  ;
        RECT 8.3120 20.3390 8.3300 20.3630 ;
    END
  END wd[11]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 21.5150 8.5970 21.5390 ;
      LAYER M3  ;
        RECT 8.5370 21.4645 8.5550 21.7040 ;
      LAYER V3  ;
        RECT 8.5370 21.5150 8.5550 21.5390 ;
    END
  END dataout[12]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 21.4190 8.6650 21.4430 ;
      LAYER M3  ;
        RECT 8.3120 21.3570 8.3300 21.7620 ;
      LAYER V3  ;
        RECT 8.3120 21.4190 8.3300 21.4430 ;
    END
  END wd[12]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 22.5950 8.5970 22.6190 ;
      LAYER M3  ;
        RECT 8.5370 22.5445 8.5550 22.7840 ;
      LAYER V3  ;
        RECT 8.5370 22.5950 8.5550 22.6190 ;
    END
  END dataout[13]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 22.4990 8.6650 22.5230 ;
      LAYER M3  ;
        RECT 8.3120 22.4370 8.3300 22.8420 ;
      LAYER V3  ;
        RECT 8.3120 22.4990 8.3300 22.5230 ;
    END
  END wd[13]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.6750 8.5970 23.6990 ;
      LAYER M3  ;
        RECT 8.5370 23.6245 8.5550 23.8640 ;
      LAYER V3  ;
        RECT 8.5370 23.6750 8.5550 23.6990 ;
    END
  END dataout[14]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.5790 8.6650 23.6030 ;
      LAYER M3  ;
        RECT 8.3120 23.5170 8.3300 23.9220 ;
      LAYER V3  ;
        RECT 8.3120 23.5790 8.3300 23.6030 ;
    END
  END wd[14]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.7550 8.5970 24.7790 ;
      LAYER M3  ;
        RECT 8.5370 24.7045 8.5550 24.9440 ;
      LAYER V3  ;
        RECT 8.5370 24.7550 8.5550 24.7790 ;
    END
  END dataout[15]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.6590 8.6650 24.6830 ;
      LAYER M3  ;
        RECT 8.3120 24.5970 8.3300 25.0020 ;
      LAYER V3  ;
        RECT 8.3120 24.6590 8.3300 24.6830 ;
    END
  END wd[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.8350 8.5970 25.8590 ;
      LAYER M3  ;
        RECT 8.5370 25.7845 8.5550 26.0240 ;
      LAYER V3  ;
        RECT 8.5370 25.8350 8.5550 25.8590 ;
    END
  END dataout[16]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.7390 8.6650 25.7630 ;
      LAYER M3  ;
        RECT 8.3120 25.6770 8.3300 26.0820 ;
      LAYER V3  ;
        RECT 8.3120 25.7390 8.3300 25.7630 ;
    END
  END wd[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 26.9150 8.5970 26.9390 ;
      LAYER M3  ;
        RECT 8.5370 26.8645 8.5550 27.1040 ;
      LAYER V3  ;
        RECT 8.5370 26.9150 8.5550 26.9390 ;
    END
  END dataout[17]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 26.8190 8.6650 26.8430 ;
      LAYER M3  ;
        RECT 8.3120 26.7570 8.3300 27.1620 ;
      LAYER V3  ;
        RECT 8.3120 26.8190 8.3300 26.8430 ;
    END
  END wd[17]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0000 9.9570 16.5240 18.6105 ;
        RECT 0.0050 18.1035 16.5290 19.1970 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0000 9.9570 16.5240 18.6105 ;
        RECT 0.0050 18.1035 16.5290 19.1970 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
  LAYER V1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0000 9.9570 16.5240 18.6105 ;
        RECT 0.0050 18.1035 16.5290 19.1970 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
  LAYER V2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0000 9.9570 16.5240 18.6105 ;
        RECT 0.0050 18.1035 16.5290 19.1970 ;
        RECT 0.0050 19.1835 16.5290 20.2770 ;
        RECT 0.0050 20.2635 16.5290 21.3570 ;
        RECT 0.0050 21.3435 16.5290 22.4370 ;
        RECT 0.0050 22.4235 16.5290 23.5170 ;
        RECT 0.0050 23.5035 16.5290 24.5970 ;
        RECT 0.0050 24.5835 16.5290 25.6770 ;
        RECT 0.0050 25.6635 16.5290 26.7570 ;
        RECT 0.0050 26.7435 16.5290 27.8370 ;
  LAYER M3  ;
      RECT 8.6990 0.3450 8.7170 1.2805 ;
      RECT 8.6630 0.3450 8.6810 1.2805 ;
      RECT 8.6270 0.9220 8.6450 1.2445 ;
      RECT 8.5100 1.1190 8.5280 1.2285 ;
      RECT 8.5010 0.3775 8.5190 0.6170 ;
      RECT 8.4650 0.9585 8.4830 1.1120 ;
      RECT 8.3840 0.9840 8.4020 1.2420 ;
      RECT 7.8440 0.3450 7.8620 1.2805 ;
      RECT 7.8080 0.3450 7.8260 1.2805 ;
      RECT 7.7720 0.5260 7.7900 1.0940 ;
      RECT 8.6990 1.4250 8.7170 2.3605 ;
      RECT 8.6630 1.4250 8.6810 2.3605 ;
      RECT 8.6270 2.0020 8.6450 2.3245 ;
      RECT 8.5100 2.1990 8.5280 2.3085 ;
      RECT 8.5010 1.4575 8.5190 1.6970 ;
      RECT 8.4650 2.0385 8.4830 2.1920 ;
      RECT 8.3840 2.0640 8.4020 2.3220 ;
      RECT 7.8440 1.4250 7.8620 2.3605 ;
      RECT 7.8080 1.4250 7.8260 2.3605 ;
      RECT 7.7720 1.6060 7.7900 2.1740 ;
      RECT 8.6990 2.5050 8.7170 3.4405 ;
      RECT 8.6630 2.5050 8.6810 3.4405 ;
      RECT 8.6270 3.0820 8.6450 3.4045 ;
      RECT 8.5100 3.2790 8.5280 3.3885 ;
      RECT 8.5010 2.5375 8.5190 2.7770 ;
      RECT 8.4650 3.1185 8.4830 3.2720 ;
      RECT 8.3840 3.1440 8.4020 3.4020 ;
      RECT 7.8440 2.5050 7.8620 3.4405 ;
      RECT 7.8080 2.5050 7.8260 3.4405 ;
      RECT 7.7720 2.6860 7.7900 3.2540 ;
      RECT 8.6990 3.5850 8.7170 4.5205 ;
      RECT 8.6630 3.5850 8.6810 4.5205 ;
      RECT 8.6270 4.1620 8.6450 4.4845 ;
      RECT 8.5100 4.3590 8.5280 4.4685 ;
      RECT 8.5010 3.6175 8.5190 3.8570 ;
      RECT 8.4650 4.1985 8.4830 4.3520 ;
      RECT 8.3840 4.2240 8.4020 4.4820 ;
      RECT 7.8440 3.5850 7.8620 4.5205 ;
      RECT 7.8080 3.5850 7.8260 4.5205 ;
      RECT 7.7720 3.7660 7.7900 4.3340 ;
      RECT 8.6990 4.6650 8.7170 5.6005 ;
      RECT 8.6630 4.6650 8.6810 5.6005 ;
      RECT 8.6270 5.2420 8.6450 5.5645 ;
      RECT 8.5100 5.4390 8.5280 5.5485 ;
      RECT 8.5010 4.6975 8.5190 4.9370 ;
      RECT 8.4650 5.2785 8.4830 5.4320 ;
      RECT 8.3840 5.3040 8.4020 5.5620 ;
      RECT 7.8440 4.6650 7.8620 5.6005 ;
      RECT 7.8080 4.6650 7.8260 5.6005 ;
      RECT 7.7720 4.8460 7.7900 5.4140 ;
      RECT 8.6990 5.7450 8.7170 6.6805 ;
      RECT 8.6630 5.7450 8.6810 6.6805 ;
      RECT 8.6270 6.3220 8.6450 6.6445 ;
      RECT 8.5100 6.5190 8.5280 6.6285 ;
      RECT 8.5010 5.7775 8.5190 6.0170 ;
      RECT 8.4650 6.3585 8.4830 6.5120 ;
      RECT 8.3840 6.3840 8.4020 6.6420 ;
      RECT 7.8440 5.7450 7.8620 6.6805 ;
      RECT 7.8080 5.7450 7.8260 6.6805 ;
      RECT 7.7720 5.9260 7.7900 6.4940 ;
      RECT 8.6990 6.8250 8.7170 7.7605 ;
      RECT 8.6630 6.8250 8.6810 7.7605 ;
      RECT 8.6270 7.4020 8.6450 7.7245 ;
      RECT 8.5100 7.5990 8.5280 7.7085 ;
      RECT 8.5010 6.8575 8.5190 7.0970 ;
      RECT 8.4650 7.4385 8.4830 7.5920 ;
      RECT 8.3840 7.4640 8.4020 7.7220 ;
      RECT 7.8440 6.8250 7.8620 7.7605 ;
      RECT 7.8080 6.8250 7.8260 7.7605 ;
      RECT 7.7720 7.0060 7.7900 7.5740 ;
      RECT 8.6990 7.9050 8.7170 8.8405 ;
      RECT 8.6630 7.9050 8.6810 8.8405 ;
      RECT 8.6270 8.4820 8.6450 8.8045 ;
      RECT 8.5100 8.6790 8.5280 8.7885 ;
      RECT 8.5010 7.9375 8.5190 8.1770 ;
      RECT 8.4650 8.5185 8.4830 8.6720 ;
      RECT 8.3840 8.5440 8.4020 8.8020 ;
      RECT 7.8440 7.9050 7.8620 8.8405 ;
      RECT 7.8080 7.9050 7.8260 8.8405 ;
      RECT 7.7720 8.0860 7.7900 8.6540 ;
      RECT 8.6990 8.9850 8.7170 9.9205 ;
      RECT 8.6630 8.9850 8.6810 9.9205 ;
      RECT 8.6270 9.5620 8.6450 9.8845 ;
      RECT 8.5100 9.7590 8.5280 9.8685 ;
      RECT 8.5010 9.0175 8.5190 9.2570 ;
      RECT 8.4650 9.5985 8.4830 9.7520 ;
      RECT 8.3840 9.6240 8.4020 9.8820 ;
      RECT 7.8440 8.9850 7.8620 9.9205 ;
      RECT 7.8080 8.9850 7.8260 9.9205 ;
      RECT 7.7720 9.1660 7.7900 9.7340 ;
      RECT 16.3170 13.7500 16.3350 18.1040 ;
      RECT 16.2810 12.4350 16.2990 12.5040 ;
      RECT 16.2810 14.0550 16.2990 14.1380 ;
      RECT 16.2450 9.9305 16.2630 18.1375 ;
      RECT 16.2090 13.7825 16.2270 14.4725 ;
      RECT 16.2090 14.5235 16.2270 15.5100 ;
      RECT 16.2090 15.5500 16.2270 16.1670 ;
      RECT 16.1730 13.7190 16.1910 14.4238 ;
      RECT 16.1730 15.1770 16.1910 16.3470 ;
      RECT 16.1370 9.9305 16.1550 13.5270 ;
      RECT 16.0290 9.9305 16.0470 13.5270 ;
      RECT 15.9210 9.9305 15.9390 13.5270 ;
      RECT 15.8130 9.9305 15.8310 13.5270 ;
      RECT 15.7050 9.9305 15.7230 13.5270 ;
      RECT 15.5970 9.9305 15.6150 13.5270 ;
      RECT 15.4890 9.9305 15.5070 13.5270 ;
      RECT 15.3810 9.9305 15.3990 13.5270 ;
      RECT 15.2730 9.9305 15.2910 13.5270 ;
      RECT 15.1650 9.9305 15.1830 13.5270 ;
      RECT 15.0570 9.9305 15.0750 13.5270 ;
      RECT 14.9490 9.9305 14.9670 13.5270 ;
      RECT 14.8410 9.9305 14.8590 13.5270 ;
      RECT 14.7330 9.9305 14.7510 13.5270 ;
      RECT 14.6250 9.9305 14.6430 13.5270 ;
      RECT 14.5170 9.9305 14.5350 13.5270 ;
      RECT 14.4090 9.9305 14.4270 13.5270 ;
      RECT 14.3010 9.9305 14.3190 13.5270 ;
      RECT 14.1930 9.9305 14.2110 13.5270 ;
      RECT 14.0850 9.9305 14.1030 13.5270 ;
      RECT 13.9770 9.9305 13.9950 13.5270 ;
      RECT 13.8690 9.9305 13.8870 13.5270 ;
      RECT 13.7610 9.9305 13.7790 13.5270 ;
      RECT 13.6530 9.9305 13.6710 13.5270 ;
      RECT 13.5450 9.9305 13.5630 13.5270 ;
      RECT 13.4370 9.9305 13.4550 13.5270 ;
      RECT 13.3290 9.9305 13.3470 13.5270 ;
      RECT 13.2210 9.9305 13.2390 13.5270 ;
      RECT 13.1130 9.9305 13.1310 13.5270 ;
      RECT 13.0050 9.9305 13.0230 13.5270 ;
      RECT 12.8970 9.9305 12.9150 13.5270 ;
      RECT 12.7890 9.9305 12.8070 13.5270 ;
      RECT 12.6810 9.9305 12.6990 13.5270 ;
      RECT 12.5730 9.9305 12.5910 13.5270 ;
      RECT 12.4650 9.9305 12.4830 13.5270 ;
      RECT 12.3570 9.9305 12.3750 13.5270 ;
      RECT 12.2490 9.9305 12.2670 13.5270 ;
      RECT 12.1410 9.9305 12.1590 13.5270 ;
      RECT 12.0330 9.9305 12.0510 13.5270 ;
      RECT 11.9250 9.9305 11.9430 13.5270 ;
      RECT 11.8170 9.9305 11.8350 13.5270 ;
      RECT 11.7090 9.9305 11.7270 13.5270 ;
      RECT 11.6010 9.9305 11.6190 13.5270 ;
      RECT 11.4930 9.9305 11.5110 13.5270 ;
      RECT 11.3850 9.9305 11.4030 13.5270 ;
      RECT 11.2770 9.9305 11.2950 13.5270 ;
      RECT 11.1690 9.9305 11.1870 13.5270 ;
      RECT 11.0610 9.9305 11.0790 13.5270 ;
      RECT 10.9530 9.9305 10.9710 13.5270 ;
      RECT 10.8450 9.9305 10.8630 13.5270 ;
      RECT 10.7370 9.9305 10.7550 13.5270 ;
      RECT 10.6290 9.9305 10.6470 13.5270 ;
      RECT 10.5210 9.9305 10.5390 13.5270 ;
      RECT 10.4130 9.9305 10.4310 13.5270 ;
      RECT 10.3050 9.9305 10.3230 13.5270 ;
      RECT 10.1970 9.9305 10.2150 13.5270 ;
      RECT 10.0890 9.9305 10.1070 13.5270 ;
      RECT 9.9810 9.9305 9.9990 13.5270 ;
      RECT 9.8730 9.9305 9.8910 13.5270 ;
      RECT 9.7650 9.9305 9.7830 13.5270 ;
      RECT 9.6570 9.9305 9.6750 13.5270 ;
      RECT 9.5490 9.9305 9.5670 13.5270 ;
      RECT 9.5130 13.7855 9.5310 14.4275 ;
      RECT 9.5130 15.1050 9.5310 15.6370 ;
      RECT 9.4950 10.5910 9.5130 11.2670 ;
      RECT 9.4950 12.0130 9.5130 12.3110 ;
      RECT 9.4950 13.1290 9.5130 13.3910 ;
      RECT 9.4770 13.7000 9.4950 14.4725 ;
      RECT 9.4770 14.5237 9.4950 15.0150 ;
      RECT 9.4770 15.0600 9.4950 15.4310 ;
      RECT 9.4770 15.5070 9.4950 16.1670 ;
      RECT 9.4410 9.9305 9.4590 18.1375 ;
      RECT 9.4050 14.2430 9.4230 14.7075 ;
      RECT 9.3870 10.6990 9.4050 11.3300 ;
      RECT 9.3870 11.7430 9.4050 11.9330 ;
      RECT 9.3870 12.6250 9.4050 12.6740 ;
      RECT 9.3870 13.3570 9.4050 13.3940 ;
      RECT 9.3690 13.7500 9.3870 18.0995 ;
      RECT 9.2790 10.3210 9.2970 11.1230 ;
      RECT 9.2790 11.6710 9.2970 12.2390 ;
      RECT 9.2430 11.7430 9.2610 12.1130 ;
      RECT 9.2070 11.0950 9.2250 11.2310 ;
      RECT 9.2070 12.0850 9.2250 12.3110 ;
      RECT 9.2070 13.3270 9.2250 13.3910 ;
      RECT 9.1710 11.1970 9.1890 11.2340 ;
      RECT 9.1710 12.8230 9.1890 12.8660 ;
      RECT 9.1710 13.3570 9.1890 13.3940 ;
      RECT 9.1350 11.5090 9.1530 12.0050 ;
      RECT 9.1350 12.0490 9.1530 12.2390 ;
      RECT 9.1350 13.0090 9.1530 13.3190 ;
      RECT 9.0990 11.4010 9.1170 12.6480 ;
      RECT 9.0990 15.2890 9.1170 16.0190 ;
      RECT 9.0990 16.3690 9.1170 17.0990 ;
      RECT 8.7750 11.1310 8.7930 11.4290 ;
      RECT 8.7750 12.3190 8.7930 12.3830 ;
      RECT 8.7750 12.5890 8.7930 13.0490 ;
      RECT 8.7750 13.7890 8.7930 13.8260 ;
      RECT 8.7750 15.8290 8.7930 16.1270 ;
      RECT 8.7390 11.2030 8.7570 11.7080 ;
      RECT 8.7390 11.9770 8.7570 12.7790 ;
      RECT 8.7390 13.8220 8.7570 14.0930 ;
      RECT 8.7390 14.1730 8.7570 14.3990 ;
      RECT 8.7030 11.1310 8.7210 11.8070 ;
      RECT 8.7030 11.9050 8.7210 12.2390 ;
      RECT 8.7030 12.4450 8.7210 12.5810 ;
      RECT 8.7030 13.1290 8.7210 13.9310 ;
      RECT 8.7030 14.3650 8.7210 14.4020 ;
      RECT 8.7030 16.5310 8.7210 16.8650 ;
      RECT 8.6670 11.3650 8.6850 11.5010 ;
      RECT 8.6670 13.2550 8.6850 14.2370 ;
      RECT 8.6670 14.6770 8.6850 14.9750 ;
      RECT 8.6670 16.3690 8.6850 16.6310 ;
      RECT 8.6310 10.4290 8.6490 10.5830 ;
      RECT 8.6310 11.2390 8.6490 13.0250 ;
      RECT 8.6310 14.0650 8.6490 16.3970 ;
      RECT 8.6310 16.6030 8.6490 17.7110 ;
      RECT 8.3430 10.6990 8.3610 10.9610 ;
      RECT 8.3430 11.0950 8.3610 11.1590 ;
      RECT 8.3430 11.2390 8.3610 11.4650 ;
      RECT 8.3430 11.5090 8.3610 11.6990 ;
      RECT 8.3430 11.7790 8.3610 14.3990 ;
      RECT 8.3430 14.4430 8.3610 15.7490 ;
      RECT 8.3430 16.8370 8.3610 17.0990 ;
      RECT 8.3070 11.6980 8.3250 11.9690 ;
      RECT 8.3070 12.0490 8.3250 12.8870 ;
      RECT 8.3070 13.0570 8.3250 13.8950 ;
      RECT 8.3070 13.9390 8.3250 15.2090 ;
      RECT 8.3070 15.4150 8.3250 15.5870 ;
      RECT 8.3070 16.2970 8.3250 17.3690 ;
      RECT 8.2710 11.7790 8.2890 12.0500 ;
      RECT 8.2710 12.2050 8.2890 12.2420 ;
      RECT 8.2710 12.9850 8.2890 13.9670 ;
      RECT 8.2710 14.2090 8.2890 14.6690 ;
      RECT 8.2710 15.0190 8.2890 15.7580 ;
      RECT 8.2350 10.8970 8.2530 11.9690 ;
      RECT 8.2350 13.5610 8.2530 13.7780 ;
      RECT 8.2350 14.9470 8.2530 15.2450 ;
      RECT 8.1990 11.5450 8.2170 12.0050 ;
      RECT 8.1990 13.1290 8.2170 13.3190 ;
      RECT 8.1990 13.3600 8.2170 13.3970 ;
      RECT 8.1990 13.6330 8.2170 13.9670 ;
      RECT 8.1990 14.1010 8.2170 15.4430 ;
      RECT 8.1990 15.5500 8.2170 16.6670 ;
      RECT 8.1630 10.9690 8.1810 11.1590 ;
      RECT 8.1630 11.3650 8.1810 11.5010 ;
      RECT 8.1630 11.7790 8.1810 14.9390 ;
      RECT 8.1630 15.0190 8.1810 15.4790 ;
      RECT 8.1630 16.0990 8.1810 16.5590 ;
      RECT 8.1630 17.4130 8.1810 17.6390 ;
      RECT 8.1270 9.9570 8.1450 10.1110 ;
      RECT 8.1270 17.9520 8.1450 18.1180 ;
      RECT 8.0910 9.9570 8.1090 10.0070 ;
      RECT 8.0190 9.9570 8.0370 10.0285 ;
      RECT 8.0190 18.0215 8.0370 18.1375 ;
      RECT 7.8750 11.4730 7.8930 11.6630 ;
      RECT 7.8750 12.2110 7.8930 12.5810 ;
      RECT 7.8750 14.1730 7.8930 14.3990 ;
      RECT 7.8750 14.7130 7.8930 15.8570 ;
      RECT 7.8750 16.6390 7.8930 17.0990 ;
      RECT 7.8750 17.6770 7.8930 17.7140 ;
      RECT 7.8390 10.4290 7.8570 10.9250 ;
      RECT 7.8390 14.5090 7.8570 14.5460 ;
      RECT 7.8390 15.5860 7.8570 16.3970 ;
      RECT 7.8030 10.8970 7.8210 11.1590 ;
      RECT 7.8030 11.4370 7.8210 11.7710 ;
      RECT 7.8030 11.9770 7.8210 12.0770 ;
      RECT 7.8030 12.8590 7.8210 15.6230 ;
      RECT 7.8030 15.7570 7.8210 15.9830 ;
      RECT 7.7670 10.5550 7.7850 11.6990 ;
      RECT 7.7670 15.2890 7.7850 15.4790 ;
      RECT 7.7670 16.0930 7.7850 16.1300 ;
      RECT 7.7670 16.3690 7.7850 17.1710 ;
      RECT 7.7310 11.5090 7.7490 12.5090 ;
      RECT 7.7310 15.9490 7.7490 15.9860 ;
      RECT 7.3710 11.0950 7.3890 11.5010 ;
      RECT 7.2990 11.1310 7.3170 11.7350 ;
      RECT 7.2630 10.9690 7.2810 11.0330 ;
      RECT 7.2270 10.0100 7.2450 10.0610 ;
      RECT 7.2270 13.1290 7.2450 13.3190 ;
      RECT 7.2090 13.7500 7.2270 18.0985 ;
      RECT 7.1370 13.7500 7.1550 18.0995 ;
      RECT 7.1190 10.4290 7.1370 10.6190 ;
      RECT 7.1190 11.2030 7.1370 13.4630 ;
      RECT 7.1010 14.2430 7.1190 14.7075 ;
      RECT 7.0650 9.9305 7.0830 18.1375 ;
      RECT 7.0290 13.7000 7.0470 14.4725 ;
      RECT 7.0290 14.5237 7.0470 15.0150 ;
      RECT 7.0290 15.0600 7.0470 15.4310 ;
      RECT 7.0290 15.5070 7.0470 16.1670 ;
      RECT 7.0110 10.4290 7.0290 10.9250 ;
      RECT 7.0110 11.7070 7.0290 12.2750 ;
      RECT 7.0110 12.5890 7.0290 13.3190 ;
      RECT 6.9930 13.7855 7.0110 14.4275 ;
      RECT 6.9930 15.1050 7.0110 15.6370 ;
      RECT 6.9570 9.9305 6.9750 13.5270 ;
      RECT 6.8490 9.9305 6.8670 13.5270 ;
      RECT 6.7410 9.9305 6.7590 13.5270 ;
      RECT 6.6330 9.9305 6.6510 13.5270 ;
      RECT 6.5250 9.9305 6.5430 13.5270 ;
      RECT 6.4170 9.9305 6.4350 13.5270 ;
      RECT 6.3090 9.9305 6.3270 13.5270 ;
      RECT 6.2010 9.9305 6.2190 13.5270 ;
      RECT 6.0930 9.9305 6.1110 13.5270 ;
      RECT 5.9850 9.9305 6.0030 13.5270 ;
      RECT 5.8770 9.9305 5.8950 13.5270 ;
      RECT 5.7690 9.9305 5.7870 13.5270 ;
      RECT 5.6610 9.9305 5.6790 13.5270 ;
      RECT 5.5530 9.9305 5.5710 13.5270 ;
      RECT 5.4450 9.9305 5.4630 13.5270 ;
      RECT 5.3370 9.9305 5.3550 13.5270 ;
      RECT 5.2290 9.9305 5.2470 13.5270 ;
      RECT 5.1210 9.9305 5.1390 13.5270 ;
      RECT 5.0130 9.9305 5.0310 13.5270 ;
      RECT 4.9050 9.9305 4.9230 13.5270 ;
      RECT 4.7970 9.9305 4.8150 13.5270 ;
      RECT 4.6890 9.9305 4.7070 13.5270 ;
      RECT 4.5810 9.9305 4.5990 13.5270 ;
      RECT 4.4730 9.9305 4.4910 13.5270 ;
      RECT 4.3650 9.9305 4.3830 13.5270 ;
      RECT 4.2570 9.9305 4.2750 13.5270 ;
      RECT 4.1490 9.9305 4.1670 13.5270 ;
      RECT 4.0410 9.9305 4.0590 13.5270 ;
      RECT 3.9330 9.9305 3.9510 13.5270 ;
      RECT 3.8250 9.9305 3.8430 13.5270 ;
      RECT 3.7170 9.9305 3.7350 13.5270 ;
      RECT 3.6090 9.9305 3.6270 13.5270 ;
      RECT 3.5010 9.9305 3.5190 13.5270 ;
      RECT 3.3930 9.9305 3.4110 13.5270 ;
      RECT 3.2850 9.9305 3.3030 13.5270 ;
      RECT 3.1770 9.9305 3.1950 13.5270 ;
      RECT 3.0690 9.9305 3.0870 13.5270 ;
      RECT 2.9610 9.9305 2.9790 13.5270 ;
      RECT 2.8530 9.9305 2.8710 13.5270 ;
      RECT 2.7450 9.9305 2.7630 13.5270 ;
      RECT 2.6370 9.9305 2.6550 13.5270 ;
      RECT 2.5290 9.9305 2.5470 13.5270 ;
      RECT 2.4210 9.9305 2.4390 13.5270 ;
      RECT 2.3130 9.9305 2.3310 13.5270 ;
      RECT 2.2050 9.9305 2.2230 13.5270 ;
      RECT 2.0970 9.9305 2.1150 13.5270 ;
      RECT 1.9890 9.9305 2.0070 13.5270 ;
      RECT 1.8810 9.9305 1.8990 13.5270 ;
      RECT 1.7730 9.9305 1.7910 13.5270 ;
      RECT 1.6650 9.9305 1.6830 13.5270 ;
      RECT 1.5570 9.9305 1.5750 13.5270 ;
      RECT 1.4490 9.9305 1.4670 13.5270 ;
      RECT 1.3410 9.9305 1.3590 13.5270 ;
      RECT 1.2330 9.9305 1.2510 13.5270 ;
      RECT 1.1250 9.9305 1.1430 13.5270 ;
      RECT 1.0170 9.9305 1.0350 13.5270 ;
      RECT 0.9090 9.9305 0.9270 13.5270 ;
      RECT 0.8010 9.9305 0.8190 13.5270 ;
      RECT 0.6930 9.9305 0.7110 13.5270 ;
      RECT 0.5850 9.9305 0.6030 13.5270 ;
      RECT 0.4770 9.9305 0.4950 13.5270 ;
      RECT 0.3690 9.9305 0.3870 13.5270 ;
      RECT 0.3330 13.7190 0.3510 14.4238 ;
      RECT 0.3330 15.1770 0.3510 16.3470 ;
      RECT 0.2970 13.7825 0.3150 14.4725 ;
      RECT 0.2970 14.5235 0.3150 15.5100 ;
      RECT 0.2970 15.5500 0.3150 16.1670 ;
      RECT 0.2610 9.9305 0.2790 18.1375 ;
      RECT 0.2250 12.4350 0.2430 12.5040 ;
      RECT 0.2250 14.0550 0.2430 14.1380 ;
      RECT 0.1890 13.7500 0.2070 18.1040 ;
        RECT 8.6990 18.1920 8.7170 19.1275 ;
        RECT 8.6630 18.1920 8.6810 19.1275 ;
        RECT 8.6270 18.7690 8.6450 19.0915 ;
        RECT 8.5100 18.9660 8.5280 19.0755 ;
        RECT 8.5010 18.2245 8.5190 18.4640 ;
        RECT 8.4650 18.8055 8.4830 18.9590 ;
        RECT 8.3840 18.8310 8.4020 19.0890 ;
        RECT 7.8440 18.1920 7.8620 19.1275 ;
        RECT 7.8080 18.1920 7.8260 19.1275 ;
        RECT 7.7720 18.3730 7.7900 18.9410 ;
        RECT 8.6990 19.2720 8.7170 20.2075 ;
        RECT 8.6630 19.2720 8.6810 20.2075 ;
        RECT 8.6270 19.8490 8.6450 20.1715 ;
        RECT 8.5100 20.0460 8.5280 20.1555 ;
        RECT 8.5010 19.3045 8.5190 19.5440 ;
        RECT 8.4650 19.8855 8.4830 20.0390 ;
        RECT 8.3840 19.9110 8.4020 20.1690 ;
        RECT 7.8440 19.2720 7.8620 20.2075 ;
        RECT 7.8080 19.2720 7.8260 20.2075 ;
        RECT 7.7720 19.4530 7.7900 20.0210 ;
        RECT 8.6990 20.3520 8.7170 21.2875 ;
        RECT 8.6630 20.3520 8.6810 21.2875 ;
        RECT 8.6270 20.9290 8.6450 21.2515 ;
        RECT 8.5100 21.1260 8.5280 21.2355 ;
        RECT 8.5010 20.3845 8.5190 20.6240 ;
        RECT 8.4650 20.9655 8.4830 21.1190 ;
        RECT 8.3840 20.9910 8.4020 21.2490 ;
        RECT 7.8440 20.3520 7.8620 21.2875 ;
        RECT 7.8080 20.3520 7.8260 21.2875 ;
        RECT 7.7720 20.5330 7.7900 21.1010 ;
        RECT 8.6990 21.4320 8.7170 22.3675 ;
        RECT 8.6630 21.4320 8.6810 22.3675 ;
        RECT 8.6270 22.0090 8.6450 22.3315 ;
        RECT 8.5100 22.2060 8.5280 22.3155 ;
        RECT 8.5010 21.4645 8.5190 21.7040 ;
        RECT 8.4650 22.0455 8.4830 22.1990 ;
        RECT 8.3840 22.0710 8.4020 22.3290 ;
        RECT 7.8440 21.4320 7.8620 22.3675 ;
        RECT 7.8080 21.4320 7.8260 22.3675 ;
        RECT 7.7720 21.6130 7.7900 22.1810 ;
        RECT 8.6990 22.5120 8.7170 23.4475 ;
        RECT 8.6630 22.5120 8.6810 23.4475 ;
        RECT 8.6270 23.0890 8.6450 23.4115 ;
        RECT 8.5100 23.2860 8.5280 23.3955 ;
        RECT 8.5010 22.5445 8.5190 22.7840 ;
        RECT 8.4650 23.1255 8.4830 23.2790 ;
        RECT 8.3840 23.1510 8.4020 23.4090 ;
        RECT 7.8440 22.5120 7.8620 23.4475 ;
        RECT 7.8080 22.5120 7.8260 23.4475 ;
        RECT 7.7720 22.6930 7.7900 23.2610 ;
        RECT 8.6990 23.5920 8.7170 24.5275 ;
        RECT 8.6630 23.5920 8.6810 24.5275 ;
        RECT 8.6270 24.1690 8.6450 24.4915 ;
        RECT 8.5100 24.3660 8.5280 24.4755 ;
        RECT 8.5010 23.6245 8.5190 23.8640 ;
        RECT 8.4650 24.2055 8.4830 24.3590 ;
        RECT 8.3840 24.2310 8.4020 24.4890 ;
        RECT 7.8440 23.5920 7.8620 24.5275 ;
        RECT 7.8080 23.5920 7.8260 24.5275 ;
        RECT 7.7720 23.7730 7.7900 24.3410 ;
        RECT 8.6990 24.6720 8.7170 25.6075 ;
        RECT 8.6630 24.6720 8.6810 25.6075 ;
        RECT 8.6270 25.2490 8.6450 25.5715 ;
        RECT 8.5100 25.4460 8.5280 25.5555 ;
        RECT 8.5010 24.7045 8.5190 24.9440 ;
        RECT 8.4650 25.2855 8.4830 25.4390 ;
        RECT 8.3840 25.3110 8.4020 25.5690 ;
        RECT 7.8440 24.6720 7.8620 25.6075 ;
        RECT 7.8080 24.6720 7.8260 25.6075 ;
        RECT 7.7720 24.8530 7.7900 25.4210 ;
        RECT 8.6990 25.7520 8.7170 26.6875 ;
        RECT 8.6630 25.7520 8.6810 26.6875 ;
        RECT 8.6270 26.3290 8.6450 26.6515 ;
        RECT 8.5100 26.5260 8.5280 26.6355 ;
        RECT 8.5010 25.7845 8.5190 26.0240 ;
        RECT 8.4650 26.3655 8.4830 26.5190 ;
        RECT 8.3840 26.3910 8.4020 26.6490 ;
        RECT 7.8440 25.7520 7.8620 26.6875 ;
        RECT 7.8080 25.7520 7.8260 26.6875 ;
        RECT 7.7720 25.9330 7.7900 26.5010 ;
        RECT 8.6990 26.8320 8.7170 27.7675 ;
        RECT 8.6630 26.8320 8.6810 27.7675 ;
        RECT 8.6270 27.4090 8.6450 27.7315 ;
        RECT 8.5100 27.6060 8.5280 27.7155 ;
        RECT 8.5010 26.8645 8.5190 27.1040 ;
        RECT 8.4650 27.4455 8.4830 27.5990 ;
        RECT 8.3840 27.4710 8.4020 27.7290 ;
        RECT 7.8440 26.8320 7.8620 27.7675 ;
        RECT 7.8080 26.8320 7.8260 27.7675 ;
        RECT 7.7720 27.0130 7.7900 27.5810 ;
  LAYER M3 SPACING 0.018  ;
      RECT 8.6410 0.2565 8.7690 1.3500 ;
      RECT 8.6270 0.9220 8.7690 1.2445 ;
      RECT 8.4790 0.6490 8.5410 1.3500 ;
      RECT 8.4650 0.9585 8.5410 1.1120 ;
      RECT 8.4790 0.2565 8.5050 1.3500 ;
      RECT 8.4790 0.3775 8.5190 0.6170 ;
      RECT 8.4790 0.2565 8.5410 0.3455 ;
      RECT 8.1820 0.7070 8.3880 1.3500 ;
      RECT 8.3620 0.2565 8.3880 1.3500 ;
      RECT 8.1820 0.9840 8.4020 1.2420 ;
      RECT 8.1820 0.2565 8.2800 1.3500 ;
      RECT 7.7650 0.2565 7.8480 1.3500 ;
      RECT 7.7650 0.3450 7.8620 1.2805 ;
      RECT 16.4440 0.2565 16.5290 1.3500 ;
      RECT 16.3000 0.2565 16.3260 1.3500 ;
      RECT 16.1920 0.2565 16.2180 1.3500 ;
      RECT 16.0840 0.2565 16.1100 1.3500 ;
      RECT 15.9760 0.2565 16.0020 1.3500 ;
      RECT 15.8680 0.2565 15.8940 1.3500 ;
      RECT 15.7600 0.2565 15.7860 1.3500 ;
      RECT 15.6520 0.2565 15.6780 1.3500 ;
      RECT 15.5440 0.2565 15.5700 1.3500 ;
      RECT 15.4360 0.2565 15.4620 1.3500 ;
      RECT 15.3280 0.2565 15.3540 1.3500 ;
      RECT 15.2200 0.2565 15.2460 1.3500 ;
      RECT 15.1120 0.2565 15.1380 1.3500 ;
      RECT 15.0040 0.2565 15.0300 1.3500 ;
      RECT 14.8960 0.2565 14.9220 1.3500 ;
      RECT 14.7880 0.2565 14.8140 1.3500 ;
      RECT 14.6800 0.2565 14.7060 1.3500 ;
      RECT 14.5720 0.2565 14.5980 1.3500 ;
      RECT 14.4640 0.2565 14.4900 1.3500 ;
      RECT 14.3560 0.2565 14.3820 1.3500 ;
      RECT 14.2480 0.2565 14.2740 1.3500 ;
      RECT 14.1400 0.2565 14.1660 1.3500 ;
      RECT 14.0320 0.2565 14.0580 1.3500 ;
      RECT 13.9240 0.2565 13.9500 1.3500 ;
      RECT 13.8160 0.2565 13.8420 1.3500 ;
      RECT 13.7080 0.2565 13.7340 1.3500 ;
      RECT 13.6000 0.2565 13.6260 1.3500 ;
      RECT 13.4920 0.2565 13.5180 1.3500 ;
      RECT 13.3840 0.2565 13.4100 1.3500 ;
      RECT 13.2760 0.2565 13.3020 1.3500 ;
      RECT 13.1680 0.2565 13.1940 1.3500 ;
      RECT 13.0600 0.2565 13.0860 1.3500 ;
      RECT 12.9520 0.2565 12.9780 1.3500 ;
      RECT 12.8440 0.2565 12.8700 1.3500 ;
      RECT 12.7360 0.2565 12.7620 1.3500 ;
      RECT 12.6280 0.2565 12.6540 1.3500 ;
      RECT 12.5200 0.2565 12.5460 1.3500 ;
      RECT 12.4120 0.2565 12.4380 1.3500 ;
      RECT 12.3040 0.2565 12.3300 1.3500 ;
      RECT 12.1960 0.2565 12.2220 1.3500 ;
      RECT 12.0880 0.2565 12.1140 1.3500 ;
      RECT 11.9800 0.2565 12.0060 1.3500 ;
      RECT 11.8720 0.2565 11.8980 1.3500 ;
      RECT 11.7640 0.2565 11.7900 1.3500 ;
      RECT 11.6560 0.2565 11.6820 1.3500 ;
      RECT 11.5480 0.2565 11.5740 1.3500 ;
      RECT 11.4400 0.2565 11.4660 1.3500 ;
      RECT 11.3320 0.2565 11.3580 1.3500 ;
      RECT 11.2240 0.2565 11.2500 1.3500 ;
      RECT 11.1160 0.2565 11.1420 1.3500 ;
      RECT 11.0080 0.2565 11.0340 1.3500 ;
      RECT 10.9000 0.2565 10.9260 1.3500 ;
      RECT 10.7920 0.2565 10.8180 1.3500 ;
      RECT 10.6840 0.2565 10.7100 1.3500 ;
      RECT 10.5760 0.2565 10.6020 1.3500 ;
      RECT 10.4680 0.2565 10.4940 1.3500 ;
      RECT 10.3600 0.2565 10.3860 1.3500 ;
      RECT 10.2520 0.2565 10.2780 1.3500 ;
      RECT 10.1440 0.2565 10.1700 1.3500 ;
      RECT 10.0360 0.2565 10.0620 1.3500 ;
      RECT 9.9280 0.2565 9.9540 1.3500 ;
      RECT 9.8200 0.2565 9.8460 1.3500 ;
      RECT 9.7120 0.2565 9.7380 1.3500 ;
      RECT 9.6040 0.2565 9.6300 1.3500 ;
      RECT 9.4960 0.2565 9.5220 1.3500 ;
      RECT 9.3880 0.2565 9.4140 1.3500 ;
      RECT 9.1750 0.2565 9.2520 1.3500 ;
      RECT 7.2820 0.2565 7.3590 1.3500 ;
      RECT 7.1200 0.2565 7.1460 1.3500 ;
      RECT 7.0120 0.2565 7.0380 1.3500 ;
      RECT 6.9040 0.2565 6.9300 1.3500 ;
      RECT 6.7960 0.2565 6.8220 1.3500 ;
      RECT 6.6880 0.2565 6.7140 1.3500 ;
      RECT 6.5800 0.2565 6.6060 1.3500 ;
      RECT 6.4720 0.2565 6.4980 1.3500 ;
      RECT 6.3640 0.2565 6.3900 1.3500 ;
      RECT 6.2560 0.2565 6.2820 1.3500 ;
      RECT 6.1480 0.2565 6.1740 1.3500 ;
      RECT 6.0400 0.2565 6.0660 1.3500 ;
      RECT 5.9320 0.2565 5.9580 1.3500 ;
      RECT 5.8240 0.2565 5.8500 1.3500 ;
      RECT 5.7160 0.2565 5.7420 1.3500 ;
      RECT 5.6080 0.2565 5.6340 1.3500 ;
      RECT 5.5000 0.2565 5.5260 1.3500 ;
      RECT 5.3920 0.2565 5.4180 1.3500 ;
      RECT 5.2840 0.2565 5.3100 1.3500 ;
      RECT 5.1760 0.2565 5.2020 1.3500 ;
      RECT 5.0680 0.2565 5.0940 1.3500 ;
      RECT 4.9600 0.2565 4.9860 1.3500 ;
      RECT 4.8520 0.2565 4.8780 1.3500 ;
      RECT 4.7440 0.2565 4.7700 1.3500 ;
      RECT 4.6360 0.2565 4.6620 1.3500 ;
      RECT 4.5280 0.2565 4.5540 1.3500 ;
      RECT 4.4200 0.2565 4.4460 1.3500 ;
      RECT 4.3120 0.2565 4.3380 1.3500 ;
      RECT 4.2040 0.2565 4.2300 1.3500 ;
      RECT 4.0960 0.2565 4.1220 1.3500 ;
      RECT 3.9880 0.2565 4.0140 1.3500 ;
      RECT 3.8800 0.2565 3.9060 1.3500 ;
      RECT 3.7720 0.2565 3.7980 1.3500 ;
      RECT 3.6640 0.2565 3.6900 1.3500 ;
      RECT 3.5560 0.2565 3.5820 1.3500 ;
      RECT 3.4480 0.2565 3.4740 1.3500 ;
      RECT 3.3400 0.2565 3.3660 1.3500 ;
      RECT 3.2320 0.2565 3.2580 1.3500 ;
      RECT 3.1240 0.2565 3.1500 1.3500 ;
      RECT 3.0160 0.2565 3.0420 1.3500 ;
      RECT 2.9080 0.2565 2.9340 1.3500 ;
      RECT 2.8000 0.2565 2.8260 1.3500 ;
      RECT 2.6920 0.2565 2.7180 1.3500 ;
      RECT 2.5840 0.2565 2.6100 1.3500 ;
      RECT 2.4760 0.2565 2.5020 1.3500 ;
      RECT 2.3680 0.2565 2.3940 1.3500 ;
      RECT 2.2600 0.2565 2.2860 1.3500 ;
      RECT 2.1520 0.2565 2.1780 1.3500 ;
      RECT 2.0440 0.2565 2.0700 1.3500 ;
      RECT 1.9360 0.2565 1.9620 1.3500 ;
      RECT 1.8280 0.2565 1.8540 1.3500 ;
      RECT 1.7200 0.2565 1.7460 1.3500 ;
      RECT 1.6120 0.2565 1.6380 1.3500 ;
      RECT 1.5040 0.2565 1.5300 1.3500 ;
      RECT 1.3960 0.2565 1.4220 1.3500 ;
      RECT 1.2880 0.2565 1.3140 1.3500 ;
      RECT 1.1800 0.2565 1.2060 1.3500 ;
      RECT 1.0720 0.2565 1.0980 1.3500 ;
      RECT 0.9640 0.2565 0.9900 1.3500 ;
      RECT 0.8560 0.2565 0.8820 1.3500 ;
      RECT 0.7480 0.2565 0.7740 1.3500 ;
      RECT 0.6400 0.2565 0.6660 1.3500 ;
      RECT 0.5320 0.2565 0.5580 1.3500 ;
      RECT 0.4240 0.2565 0.4500 1.3500 ;
      RECT 0.3160 0.2565 0.3420 1.3500 ;
      RECT 0.2080 0.2565 0.2340 1.3500 ;
      RECT 0.0050 0.2565 0.0900 1.3500 ;
      RECT 8.6410 1.3365 8.7690 2.4300 ;
      RECT 8.6270 2.0020 8.7690 2.3245 ;
      RECT 8.4790 1.7290 8.5410 2.4300 ;
      RECT 8.4650 2.0385 8.5410 2.1920 ;
      RECT 8.4790 1.3365 8.5050 2.4300 ;
      RECT 8.4790 1.4575 8.5190 1.6970 ;
      RECT 8.4790 1.3365 8.5410 1.4255 ;
      RECT 8.1820 1.7870 8.3880 2.4300 ;
      RECT 8.3620 1.3365 8.3880 2.4300 ;
      RECT 8.1820 2.0640 8.4020 2.3220 ;
      RECT 8.1820 1.3365 8.2800 2.4300 ;
      RECT 7.7650 1.3365 7.8480 2.4300 ;
      RECT 7.7650 1.4250 7.8620 2.3605 ;
      RECT 16.4440 1.3365 16.5290 2.4300 ;
      RECT 16.3000 1.3365 16.3260 2.4300 ;
      RECT 16.1920 1.3365 16.2180 2.4300 ;
      RECT 16.0840 1.3365 16.1100 2.4300 ;
      RECT 15.9760 1.3365 16.0020 2.4300 ;
      RECT 15.8680 1.3365 15.8940 2.4300 ;
      RECT 15.7600 1.3365 15.7860 2.4300 ;
      RECT 15.6520 1.3365 15.6780 2.4300 ;
      RECT 15.5440 1.3365 15.5700 2.4300 ;
      RECT 15.4360 1.3365 15.4620 2.4300 ;
      RECT 15.3280 1.3365 15.3540 2.4300 ;
      RECT 15.2200 1.3365 15.2460 2.4300 ;
      RECT 15.1120 1.3365 15.1380 2.4300 ;
      RECT 15.0040 1.3365 15.0300 2.4300 ;
      RECT 14.8960 1.3365 14.9220 2.4300 ;
      RECT 14.7880 1.3365 14.8140 2.4300 ;
      RECT 14.6800 1.3365 14.7060 2.4300 ;
      RECT 14.5720 1.3365 14.5980 2.4300 ;
      RECT 14.4640 1.3365 14.4900 2.4300 ;
      RECT 14.3560 1.3365 14.3820 2.4300 ;
      RECT 14.2480 1.3365 14.2740 2.4300 ;
      RECT 14.1400 1.3365 14.1660 2.4300 ;
      RECT 14.0320 1.3365 14.0580 2.4300 ;
      RECT 13.9240 1.3365 13.9500 2.4300 ;
      RECT 13.8160 1.3365 13.8420 2.4300 ;
      RECT 13.7080 1.3365 13.7340 2.4300 ;
      RECT 13.6000 1.3365 13.6260 2.4300 ;
      RECT 13.4920 1.3365 13.5180 2.4300 ;
      RECT 13.3840 1.3365 13.4100 2.4300 ;
      RECT 13.2760 1.3365 13.3020 2.4300 ;
      RECT 13.1680 1.3365 13.1940 2.4300 ;
      RECT 13.0600 1.3365 13.0860 2.4300 ;
      RECT 12.9520 1.3365 12.9780 2.4300 ;
      RECT 12.8440 1.3365 12.8700 2.4300 ;
      RECT 12.7360 1.3365 12.7620 2.4300 ;
      RECT 12.6280 1.3365 12.6540 2.4300 ;
      RECT 12.5200 1.3365 12.5460 2.4300 ;
      RECT 12.4120 1.3365 12.4380 2.4300 ;
      RECT 12.3040 1.3365 12.3300 2.4300 ;
      RECT 12.1960 1.3365 12.2220 2.4300 ;
      RECT 12.0880 1.3365 12.1140 2.4300 ;
      RECT 11.9800 1.3365 12.0060 2.4300 ;
      RECT 11.8720 1.3365 11.8980 2.4300 ;
      RECT 11.7640 1.3365 11.7900 2.4300 ;
      RECT 11.6560 1.3365 11.6820 2.4300 ;
      RECT 11.5480 1.3365 11.5740 2.4300 ;
      RECT 11.4400 1.3365 11.4660 2.4300 ;
      RECT 11.3320 1.3365 11.3580 2.4300 ;
      RECT 11.2240 1.3365 11.2500 2.4300 ;
      RECT 11.1160 1.3365 11.1420 2.4300 ;
      RECT 11.0080 1.3365 11.0340 2.4300 ;
      RECT 10.9000 1.3365 10.9260 2.4300 ;
      RECT 10.7920 1.3365 10.8180 2.4300 ;
      RECT 10.6840 1.3365 10.7100 2.4300 ;
      RECT 10.5760 1.3365 10.6020 2.4300 ;
      RECT 10.4680 1.3365 10.4940 2.4300 ;
      RECT 10.3600 1.3365 10.3860 2.4300 ;
      RECT 10.2520 1.3365 10.2780 2.4300 ;
      RECT 10.1440 1.3365 10.1700 2.4300 ;
      RECT 10.0360 1.3365 10.0620 2.4300 ;
      RECT 9.9280 1.3365 9.9540 2.4300 ;
      RECT 9.8200 1.3365 9.8460 2.4300 ;
      RECT 9.7120 1.3365 9.7380 2.4300 ;
      RECT 9.6040 1.3365 9.6300 2.4300 ;
      RECT 9.4960 1.3365 9.5220 2.4300 ;
      RECT 9.3880 1.3365 9.4140 2.4300 ;
      RECT 9.1750 1.3365 9.2520 2.4300 ;
      RECT 7.2820 1.3365 7.3590 2.4300 ;
      RECT 7.1200 1.3365 7.1460 2.4300 ;
      RECT 7.0120 1.3365 7.0380 2.4300 ;
      RECT 6.9040 1.3365 6.9300 2.4300 ;
      RECT 6.7960 1.3365 6.8220 2.4300 ;
      RECT 6.6880 1.3365 6.7140 2.4300 ;
      RECT 6.5800 1.3365 6.6060 2.4300 ;
      RECT 6.4720 1.3365 6.4980 2.4300 ;
      RECT 6.3640 1.3365 6.3900 2.4300 ;
      RECT 6.2560 1.3365 6.2820 2.4300 ;
      RECT 6.1480 1.3365 6.1740 2.4300 ;
      RECT 6.0400 1.3365 6.0660 2.4300 ;
      RECT 5.9320 1.3365 5.9580 2.4300 ;
      RECT 5.8240 1.3365 5.8500 2.4300 ;
      RECT 5.7160 1.3365 5.7420 2.4300 ;
      RECT 5.6080 1.3365 5.6340 2.4300 ;
      RECT 5.5000 1.3365 5.5260 2.4300 ;
      RECT 5.3920 1.3365 5.4180 2.4300 ;
      RECT 5.2840 1.3365 5.3100 2.4300 ;
      RECT 5.1760 1.3365 5.2020 2.4300 ;
      RECT 5.0680 1.3365 5.0940 2.4300 ;
      RECT 4.9600 1.3365 4.9860 2.4300 ;
      RECT 4.8520 1.3365 4.8780 2.4300 ;
      RECT 4.7440 1.3365 4.7700 2.4300 ;
      RECT 4.6360 1.3365 4.6620 2.4300 ;
      RECT 4.5280 1.3365 4.5540 2.4300 ;
      RECT 4.4200 1.3365 4.4460 2.4300 ;
      RECT 4.3120 1.3365 4.3380 2.4300 ;
      RECT 4.2040 1.3365 4.2300 2.4300 ;
      RECT 4.0960 1.3365 4.1220 2.4300 ;
      RECT 3.9880 1.3365 4.0140 2.4300 ;
      RECT 3.8800 1.3365 3.9060 2.4300 ;
      RECT 3.7720 1.3365 3.7980 2.4300 ;
      RECT 3.6640 1.3365 3.6900 2.4300 ;
      RECT 3.5560 1.3365 3.5820 2.4300 ;
      RECT 3.4480 1.3365 3.4740 2.4300 ;
      RECT 3.3400 1.3365 3.3660 2.4300 ;
      RECT 3.2320 1.3365 3.2580 2.4300 ;
      RECT 3.1240 1.3365 3.1500 2.4300 ;
      RECT 3.0160 1.3365 3.0420 2.4300 ;
      RECT 2.9080 1.3365 2.9340 2.4300 ;
      RECT 2.8000 1.3365 2.8260 2.4300 ;
      RECT 2.6920 1.3365 2.7180 2.4300 ;
      RECT 2.5840 1.3365 2.6100 2.4300 ;
      RECT 2.4760 1.3365 2.5020 2.4300 ;
      RECT 2.3680 1.3365 2.3940 2.4300 ;
      RECT 2.2600 1.3365 2.2860 2.4300 ;
      RECT 2.1520 1.3365 2.1780 2.4300 ;
      RECT 2.0440 1.3365 2.0700 2.4300 ;
      RECT 1.9360 1.3365 1.9620 2.4300 ;
      RECT 1.8280 1.3365 1.8540 2.4300 ;
      RECT 1.7200 1.3365 1.7460 2.4300 ;
      RECT 1.6120 1.3365 1.6380 2.4300 ;
      RECT 1.5040 1.3365 1.5300 2.4300 ;
      RECT 1.3960 1.3365 1.4220 2.4300 ;
      RECT 1.2880 1.3365 1.3140 2.4300 ;
      RECT 1.1800 1.3365 1.2060 2.4300 ;
      RECT 1.0720 1.3365 1.0980 2.4300 ;
      RECT 0.9640 1.3365 0.9900 2.4300 ;
      RECT 0.8560 1.3365 0.8820 2.4300 ;
      RECT 0.7480 1.3365 0.7740 2.4300 ;
      RECT 0.6400 1.3365 0.6660 2.4300 ;
      RECT 0.5320 1.3365 0.5580 2.4300 ;
      RECT 0.4240 1.3365 0.4500 2.4300 ;
      RECT 0.3160 1.3365 0.3420 2.4300 ;
      RECT 0.2080 1.3365 0.2340 2.4300 ;
      RECT 0.0050 1.3365 0.0900 2.4300 ;
      RECT 8.6410 2.4165 8.7690 3.5100 ;
      RECT 8.6270 3.0820 8.7690 3.4045 ;
      RECT 8.4790 2.8090 8.5410 3.5100 ;
      RECT 8.4650 3.1185 8.5410 3.2720 ;
      RECT 8.4790 2.4165 8.5050 3.5100 ;
      RECT 8.4790 2.5375 8.5190 2.7770 ;
      RECT 8.4790 2.4165 8.5410 2.5055 ;
      RECT 8.1820 2.8670 8.3880 3.5100 ;
      RECT 8.3620 2.4165 8.3880 3.5100 ;
      RECT 8.1820 3.1440 8.4020 3.4020 ;
      RECT 8.1820 2.4165 8.2800 3.5100 ;
      RECT 7.7650 2.4165 7.8480 3.5100 ;
      RECT 7.7650 2.5050 7.8620 3.4405 ;
      RECT 16.4440 2.4165 16.5290 3.5100 ;
      RECT 16.3000 2.4165 16.3260 3.5100 ;
      RECT 16.1920 2.4165 16.2180 3.5100 ;
      RECT 16.0840 2.4165 16.1100 3.5100 ;
      RECT 15.9760 2.4165 16.0020 3.5100 ;
      RECT 15.8680 2.4165 15.8940 3.5100 ;
      RECT 15.7600 2.4165 15.7860 3.5100 ;
      RECT 15.6520 2.4165 15.6780 3.5100 ;
      RECT 15.5440 2.4165 15.5700 3.5100 ;
      RECT 15.4360 2.4165 15.4620 3.5100 ;
      RECT 15.3280 2.4165 15.3540 3.5100 ;
      RECT 15.2200 2.4165 15.2460 3.5100 ;
      RECT 15.1120 2.4165 15.1380 3.5100 ;
      RECT 15.0040 2.4165 15.0300 3.5100 ;
      RECT 14.8960 2.4165 14.9220 3.5100 ;
      RECT 14.7880 2.4165 14.8140 3.5100 ;
      RECT 14.6800 2.4165 14.7060 3.5100 ;
      RECT 14.5720 2.4165 14.5980 3.5100 ;
      RECT 14.4640 2.4165 14.4900 3.5100 ;
      RECT 14.3560 2.4165 14.3820 3.5100 ;
      RECT 14.2480 2.4165 14.2740 3.5100 ;
      RECT 14.1400 2.4165 14.1660 3.5100 ;
      RECT 14.0320 2.4165 14.0580 3.5100 ;
      RECT 13.9240 2.4165 13.9500 3.5100 ;
      RECT 13.8160 2.4165 13.8420 3.5100 ;
      RECT 13.7080 2.4165 13.7340 3.5100 ;
      RECT 13.6000 2.4165 13.6260 3.5100 ;
      RECT 13.4920 2.4165 13.5180 3.5100 ;
      RECT 13.3840 2.4165 13.4100 3.5100 ;
      RECT 13.2760 2.4165 13.3020 3.5100 ;
      RECT 13.1680 2.4165 13.1940 3.5100 ;
      RECT 13.0600 2.4165 13.0860 3.5100 ;
      RECT 12.9520 2.4165 12.9780 3.5100 ;
      RECT 12.8440 2.4165 12.8700 3.5100 ;
      RECT 12.7360 2.4165 12.7620 3.5100 ;
      RECT 12.6280 2.4165 12.6540 3.5100 ;
      RECT 12.5200 2.4165 12.5460 3.5100 ;
      RECT 12.4120 2.4165 12.4380 3.5100 ;
      RECT 12.3040 2.4165 12.3300 3.5100 ;
      RECT 12.1960 2.4165 12.2220 3.5100 ;
      RECT 12.0880 2.4165 12.1140 3.5100 ;
      RECT 11.9800 2.4165 12.0060 3.5100 ;
      RECT 11.8720 2.4165 11.8980 3.5100 ;
      RECT 11.7640 2.4165 11.7900 3.5100 ;
      RECT 11.6560 2.4165 11.6820 3.5100 ;
      RECT 11.5480 2.4165 11.5740 3.5100 ;
      RECT 11.4400 2.4165 11.4660 3.5100 ;
      RECT 11.3320 2.4165 11.3580 3.5100 ;
      RECT 11.2240 2.4165 11.2500 3.5100 ;
      RECT 11.1160 2.4165 11.1420 3.5100 ;
      RECT 11.0080 2.4165 11.0340 3.5100 ;
      RECT 10.9000 2.4165 10.9260 3.5100 ;
      RECT 10.7920 2.4165 10.8180 3.5100 ;
      RECT 10.6840 2.4165 10.7100 3.5100 ;
      RECT 10.5760 2.4165 10.6020 3.5100 ;
      RECT 10.4680 2.4165 10.4940 3.5100 ;
      RECT 10.3600 2.4165 10.3860 3.5100 ;
      RECT 10.2520 2.4165 10.2780 3.5100 ;
      RECT 10.1440 2.4165 10.1700 3.5100 ;
      RECT 10.0360 2.4165 10.0620 3.5100 ;
      RECT 9.9280 2.4165 9.9540 3.5100 ;
      RECT 9.8200 2.4165 9.8460 3.5100 ;
      RECT 9.7120 2.4165 9.7380 3.5100 ;
      RECT 9.6040 2.4165 9.6300 3.5100 ;
      RECT 9.4960 2.4165 9.5220 3.5100 ;
      RECT 9.3880 2.4165 9.4140 3.5100 ;
      RECT 9.1750 2.4165 9.2520 3.5100 ;
      RECT 7.2820 2.4165 7.3590 3.5100 ;
      RECT 7.1200 2.4165 7.1460 3.5100 ;
      RECT 7.0120 2.4165 7.0380 3.5100 ;
      RECT 6.9040 2.4165 6.9300 3.5100 ;
      RECT 6.7960 2.4165 6.8220 3.5100 ;
      RECT 6.6880 2.4165 6.7140 3.5100 ;
      RECT 6.5800 2.4165 6.6060 3.5100 ;
      RECT 6.4720 2.4165 6.4980 3.5100 ;
      RECT 6.3640 2.4165 6.3900 3.5100 ;
      RECT 6.2560 2.4165 6.2820 3.5100 ;
      RECT 6.1480 2.4165 6.1740 3.5100 ;
      RECT 6.0400 2.4165 6.0660 3.5100 ;
      RECT 5.9320 2.4165 5.9580 3.5100 ;
      RECT 5.8240 2.4165 5.8500 3.5100 ;
      RECT 5.7160 2.4165 5.7420 3.5100 ;
      RECT 5.6080 2.4165 5.6340 3.5100 ;
      RECT 5.5000 2.4165 5.5260 3.5100 ;
      RECT 5.3920 2.4165 5.4180 3.5100 ;
      RECT 5.2840 2.4165 5.3100 3.5100 ;
      RECT 5.1760 2.4165 5.2020 3.5100 ;
      RECT 5.0680 2.4165 5.0940 3.5100 ;
      RECT 4.9600 2.4165 4.9860 3.5100 ;
      RECT 4.8520 2.4165 4.8780 3.5100 ;
      RECT 4.7440 2.4165 4.7700 3.5100 ;
      RECT 4.6360 2.4165 4.6620 3.5100 ;
      RECT 4.5280 2.4165 4.5540 3.5100 ;
      RECT 4.4200 2.4165 4.4460 3.5100 ;
      RECT 4.3120 2.4165 4.3380 3.5100 ;
      RECT 4.2040 2.4165 4.2300 3.5100 ;
      RECT 4.0960 2.4165 4.1220 3.5100 ;
      RECT 3.9880 2.4165 4.0140 3.5100 ;
      RECT 3.8800 2.4165 3.9060 3.5100 ;
      RECT 3.7720 2.4165 3.7980 3.5100 ;
      RECT 3.6640 2.4165 3.6900 3.5100 ;
      RECT 3.5560 2.4165 3.5820 3.5100 ;
      RECT 3.4480 2.4165 3.4740 3.5100 ;
      RECT 3.3400 2.4165 3.3660 3.5100 ;
      RECT 3.2320 2.4165 3.2580 3.5100 ;
      RECT 3.1240 2.4165 3.1500 3.5100 ;
      RECT 3.0160 2.4165 3.0420 3.5100 ;
      RECT 2.9080 2.4165 2.9340 3.5100 ;
      RECT 2.8000 2.4165 2.8260 3.5100 ;
      RECT 2.6920 2.4165 2.7180 3.5100 ;
      RECT 2.5840 2.4165 2.6100 3.5100 ;
      RECT 2.4760 2.4165 2.5020 3.5100 ;
      RECT 2.3680 2.4165 2.3940 3.5100 ;
      RECT 2.2600 2.4165 2.2860 3.5100 ;
      RECT 2.1520 2.4165 2.1780 3.5100 ;
      RECT 2.0440 2.4165 2.0700 3.5100 ;
      RECT 1.9360 2.4165 1.9620 3.5100 ;
      RECT 1.8280 2.4165 1.8540 3.5100 ;
      RECT 1.7200 2.4165 1.7460 3.5100 ;
      RECT 1.6120 2.4165 1.6380 3.5100 ;
      RECT 1.5040 2.4165 1.5300 3.5100 ;
      RECT 1.3960 2.4165 1.4220 3.5100 ;
      RECT 1.2880 2.4165 1.3140 3.5100 ;
      RECT 1.1800 2.4165 1.2060 3.5100 ;
      RECT 1.0720 2.4165 1.0980 3.5100 ;
      RECT 0.9640 2.4165 0.9900 3.5100 ;
      RECT 0.8560 2.4165 0.8820 3.5100 ;
      RECT 0.7480 2.4165 0.7740 3.5100 ;
      RECT 0.6400 2.4165 0.6660 3.5100 ;
      RECT 0.5320 2.4165 0.5580 3.5100 ;
      RECT 0.4240 2.4165 0.4500 3.5100 ;
      RECT 0.3160 2.4165 0.3420 3.5100 ;
      RECT 0.2080 2.4165 0.2340 3.5100 ;
      RECT 0.0050 2.4165 0.0900 3.5100 ;
      RECT 8.6410 3.4965 8.7690 4.5900 ;
      RECT 8.6270 4.1620 8.7690 4.4845 ;
      RECT 8.4790 3.8890 8.5410 4.5900 ;
      RECT 8.4650 4.1985 8.5410 4.3520 ;
      RECT 8.4790 3.4965 8.5050 4.5900 ;
      RECT 8.4790 3.6175 8.5190 3.8570 ;
      RECT 8.4790 3.4965 8.5410 3.5855 ;
      RECT 8.1820 3.9470 8.3880 4.5900 ;
      RECT 8.3620 3.4965 8.3880 4.5900 ;
      RECT 8.1820 4.2240 8.4020 4.4820 ;
      RECT 8.1820 3.4965 8.2800 4.5900 ;
      RECT 7.7650 3.4965 7.8480 4.5900 ;
      RECT 7.7650 3.5850 7.8620 4.5205 ;
      RECT 16.4440 3.4965 16.5290 4.5900 ;
      RECT 16.3000 3.4965 16.3260 4.5900 ;
      RECT 16.1920 3.4965 16.2180 4.5900 ;
      RECT 16.0840 3.4965 16.1100 4.5900 ;
      RECT 15.9760 3.4965 16.0020 4.5900 ;
      RECT 15.8680 3.4965 15.8940 4.5900 ;
      RECT 15.7600 3.4965 15.7860 4.5900 ;
      RECT 15.6520 3.4965 15.6780 4.5900 ;
      RECT 15.5440 3.4965 15.5700 4.5900 ;
      RECT 15.4360 3.4965 15.4620 4.5900 ;
      RECT 15.3280 3.4965 15.3540 4.5900 ;
      RECT 15.2200 3.4965 15.2460 4.5900 ;
      RECT 15.1120 3.4965 15.1380 4.5900 ;
      RECT 15.0040 3.4965 15.0300 4.5900 ;
      RECT 14.8960 3.4965 14.9220 4.5900 ;
      RECT 14.7880 3.4965 14.8140 4.5900 ;
      RECT 14.6800 3.4965 14.7060 4.5900 ;
      RECT 14.5720 3.4965 14.5980 4.5900 ;
      RECT 14.4640 3.4965 14.4900 4.5900 ;
      RECT 14.3560 3.4965 14.3820 4.5900 ;
      RECT 14.2480 3.4965 14.2740 4.5900 ;
      RECT 14.1400 3.4965 14.1660 4.5900 ;
      RECT 14.0320 3.4965 14.0580 4.5900 ;
      RECT 13.9240 3.4965 13.9500 4.5900 ;
      RECT 13.8160 3.4965 13.8420 4.5900 ;
      RECT 13.7080 3.4965 13.7340 4.5900 ;
      RECT 13.6000 3.4965 13.6260 4.5900 ;
      RECT 13.4920 3.4965 13.5180 4.5900 ;
      RECT 13.3840 3.4965 13.4100 4.5900 ;
      RECT 13.2760 3.4965 13.3020 4.5900 ;
      RECT 13.1680 3.4965 13.1940 4.5900 ;
      RECT 13.0600 3.4965 13.0860 4.5900 ;
      RECT 12.9520 3.4965 12.9780 4.5900 ;
      RECT 12.8440 3.4965 12.8700 4.5900 ;
      RECT 12.7360 3.4965 12.7620 4.5900 ;
      RECT 12.6280 3.4965 12.6540 4.5900 ;
      RECT 12.5200 3.4965 12.5460 4.5900 ;
      RECT 12.4120 3.4965 12.4380 4.5900 ;
      RECT 12.3040 3.4965 12.3300 4.5900 ;
      RECT 12.1960 3.4965 12.2220 4.5900 ;
      RECT 12.0880 3.4965 12.1140 4.5900 ;
      RECT 11.9800 3.4965 12.0060 4.5900 ;
      RECT 11.8720 3.4965 11.8980 4.5900 ;
      RECT 11.7640 3.4965 11.7900 4.5900 ;
      RECT 11.6560 3.4965 11.6820 4.5900 ;
      RECT 11.5480 3.4965 11.5740 4.5900 ;
      RECT 11.4400 3.4965 11.4660 4.5900 ;
      RECT 11.3320 3.4965 11.3580 4.5900 ;
      RECT 11.2240 3.4965 11.2500 4.5900 ;
      RECT 11.1160 3.4965 11.1420 4.5900 ;
      RECT 11.0080 3.4965 11.0340 4.5900 ;
      RECT 10.9000 3.4965 10.9260 4.5900 ;
      RECT 10.7920 3.4965 10.8180 4.5900 ;
      RECT 10.6840 3.4965 10.7100 4.5900 ;
      RECT 10.5760 3.4965 10.6020 4.5900 ;
      RECT 10.4680 3.4965 10.4940 4.5900 ;
      RECT 10.3600 3.4965 10.3860 4.5900 ;
      RECT 10.2520 3.4965 10.2780 4.5900 ;
      RECT 10.1440 3.4965 10.1700 4.5900 ;
      RECT 10.0360 3.4965 10.0620 4.5900 ;
      RECT 9.9280 3.4965 9.9540 4.5900 ;
      RECT 9.8200 3.4965 9.8460 4.5900 ;
      RECT 9.7120 3.4965 9.7380 4.5900 ;
      RECT 9.6040 3.4965 9.6300 4.5900 ;
      RECT 9.4960 3.4965 9.5220 4.5900 ;
      RECT 9.3880 3.4965 9.4140 4.5900 ;
      RECT 9.1750 3.4965 9.2520 4.5900 ;
      RECT 7.2820 3.4965 7.3590 4.5900 ;
      RECT 7.1200 3.4965 7.1460 4.5900 ;
      RECT 7.0120 3.4965 7.0380 4.5900 ;
      RECT 6.9040 3.4965 6.9300 4.5900 ;
      RECT 6.7960 3.4965 6.8220 4.5900 ;
      RECT 6.6880 3.4965 6.7140 4.5900 ;
      RECT 6.5800 3.4965 6.6060 4.5900 ;
      RECT 6.4720 3.4965 6.4980 4.5900 ;
      RECT 6.3640 3.4965 6.3900 4.5900 ;
      RECT 6.2560 3.4965 6.2820 4.5900 ;
      RECT 6.1480 3.4965 6.1740 4.5900 ;
      RECT 6.0400 3.4965 6.0660 4.5900 ;
      RECT 5.9320 3.4965 5.9580 4.5900 ;
      RECT 5.8240 3.4965 5.8500 4.5900 ;
      RECT 5.7160 3.4965 5.7420 4.5900 ;
      RECT 5.6080 3.4965 5.6340 4.5900 ;
      RECT 5.5000 3.4965 5.5260 4.5900 ;
      RECT 5.3920 3.4965 5.4180 4.5900 ;
      RECT 5.2840 3.4965 5.3100 4.5900 ;
      RECT 5.1760 3.4965 5.2020 4.5900 ;
      RECT 5.0680 3.4965 5.0940 4.5900 ;
      RECT 4.9600 3.4965 4.9860 4.5900 ;
      RECT 4.8520 3.4965 4.8780 4.5900 ;
      RECT 4.7440 3.4965 4.7700 4.5900 ;
      RECT 4.6360 3.4965 4.6620 4.5900 ;
      RECT 4.5280 3.4965 4.5540 4.5900 ;
      RECT 4.4200 3.4965 4.4460 4.5900 ;
      RECT 4.3120 3.4965 4.3380 4.5900 ;
      RECT 4.2040 3.4965 4.2300 4.5900 ;
      RECT 4.0960 3.4965 4.1220 4.5900 ;
      RECT 3.9880 3.4965 4.0140 4.5900 ;
      RECT 3.8800 3.4965 3.9060 4.5900 ;
      RECT 3.7720 3.4965 3.7980 4.5900 ;
      RECT 3.6640 3.4965 3.6900 4.5900 ;
      RECT 3.5560 3.4965 3.5820 4.5900 ;
      RECT 3.4480 3.4965 3.4740 4.5900 ;
      RECT 3.3400 3.4965 3.3660 4.5900 ;
      RECT 3.2320 3.4965 3.2580 4.5900 ;
      RECT 3.1240 3.4965 3.1500 4.5900 ;
      RECT 3.0160 3.4965 3.0420 4.5900 ;
      RECT 2.9080 3.4965 2.9340 4.5900 ;
      RECT 2.8000 3.4965 2.8260 4.5900 ;
      RECT 2.6920 3.4965 2.7180 4.5900 ;
      RECT 2.5840 3.4965 2.6100 4.5900 ;
      RECT 2.4760 3.4965 2.5020 4.5900 ;
      RECT 2.3680 3.4965 2.3940 4.5900 ;
      RECT 2.2600 3.4965 2.2860 4.5900 ;
      RECT 2.1520 3.4965 2.1780 4.5900 ;
      RECT 2.0440 3.4965 2.0700 4.5900 ;
      RECT 1.9360 3.4965 1.9620 4.5900 ;
      RECT 1.8280 3.4965 1.8540 4.5900 ;
      RECT 1.7200 3.4965 1.7460 4.5900 ;
      RECT 1.6120 3.4965 1.6380 4.5900 ;
      RECT 1.5040 3.4965 1.5300 4.5900 ;
      RECT 1.3960 3.4965 1.4220 4.5900 ;
      RECT 1.2880 3.4965 1.3140 4.5900 ;
      RECT 1.1800 3.4965 1.2060 4.5900 ;
      RECT 1.0720 3.4965 1.0980 4.5900 ;
      RECT 0.9640 3.4965 0.9900 4.5900 ;
      RECT 0.8560 3.4965 0.8820 4.5900 ;
      RECT 0.7480 3.4965 0.7740 4.5900 ;
      RECT 0.6400 3.4965 0.6660 4.5900 ;
      RECT 0.5320 3.4965 0.5580 4.5900 ;
      RECT 0.4240 3.4965 0.4500 4.5900 ;
      RECT 0.3160 3.4965 0.3420 4.5900 ;
      RECT 0.2080 3.4965 0.2340 4.5900 ;
      RECT 0.0050 3.4965 0.0900 4.5900 ;
      RECT 8.6410 4.5765 8.7690 5.6700 ;
      RECT 8.6270 5.2420 8.7690 5.5645 ;
      RECT 8.4790 4.9690 8.5410 5.6700 ;
      RECT 8.4650 5.2785 8.5410 5.4320 ;
      RECT 8.4790 4.5765 8.5050 5.6700 ;
      RECT 8.4790 4.6975 8.5190 4.9370 ;
      RECT 8.4790 4.5765 8.5410 4.6655 ;
      RECT 8.1820 5.0270 8.3880 5.6700 ;
      RECT 8.3620 4.5765 8.3880 5.6700 ;
      RECT 8.1820 5.3040 8.4020 5.5620 ;
      RECT 8.1820 4.5765 8.2800 5.6700 ;
      RECT 7.7650 4.5765 7.8480 5.6700 ;
      RECT 7.7650 4.6650 7.8620 5.6005 ;
      RECT 16.4440 4.5765 16.5290 5.6700 ;
      RECT 16.3000 4.5765 16.3260 5.6700 ;
      RECT 16.1920 4.5765 16.2180 5.6700 ;
      RECT 16.0840 4.5765 16.1100 5.6700 ;
      RECT 15.9760 4.5765 16.0020 5.6700 ;
      RECT 15.8680 4.5765 15.8940 5.6700 ;
      RECT 15.7600 4.5765 15.7860 5.6700 ;
      RECT 15.6520 4.5765 15.6780 5.6700 ;
      RECT 15.5440 4.5765 15.5700 5.6700 ;
      RECT 15.4360 4.5765 15.4620 5.6700 ;
      RECT 15.3280 4.5765 15.3540 5.6700 ;
      RECT 15.2200 4.5765 15.2460 5.6700 ;
      RECT 15.1120 4.5765 15.1380 5.6700 ;
      RECT 15.0040 4.5765 15.0300 5.6700 ;
      RECT 14.8960 4.5765 14.9220 5.6700 ;
      RECT 14.7880 4.5765 14.8140 5.6700 ;
      RECT 14.6800 4.5765 14.7060 5.6700 ;
      RECT 14.5720 4.5765 14.5980 5.6700 ;
      RECT 14.4640 4.5765 14.4900 5.6700 ;
      RECT 14.3560 4.5765 14.3820 5.6700 ;
      RECT 14.2480 4.5765 14.2740 5.6700 ;
      RECT 14.1400 4.5765 14.1660 5.6700 ;
      RECT 14.0320 4.5765 14.0580 5.6700 ;
      RECT 13.9240 4.5765 13.9500 5.6700 ;
      RECT 13.8160 4.5765 13.8420 5.6700 ;
      RECT 13.7080 4.5765 13.7340 5.6700 ;
      RECT 13.6000 4.5765 13.6260 5.6700 ;
      RECT 13.4920 4.5765 13.5180 5.6700 ;
      RECT 13.3840 4.5765 13.4100 5.6700 ;
      RECT 13.2760 4.5765 13.3020 5.6700 ;
      RECT 13.1680 4.5765 13.1940 5.6700 ;
      RECT 13.0600 4.5765 13.0860 5.6700 ;
      RECT 12.9520 4.5765 12.9780 5.6700 ;
      RECT 12.8440 4.5765 12.8700 5.6700 ;
      RECT 12.7360 4.5765 12.7620 5.6700 ;
      RECT 12.6280 4.5765 12.6540 5.6700 ;
      RECT 12.5200 4.5765 12.5460 5.6700 ;
      RECT 12.4120 4.5765 12.4380 5.6700 ;
      RECT 12.3040 4.5765 12.3300 5.6700 ;
      RECT 12.1960 4.5765 12.2220 5.6700 ;
      RECT 12.0880 4.5765 12.1140 5.6700 ;
      RECT 11.9800 4.5765 12.0060 5.6700 ;
      RECT 11.8720 4.5765 11.8980 5.6700 ;
      RECT 11.7640 4.5765 11.7900 5.6700 ;
      RECT 11.6560 4.5765 11.6820 5.6700 ;
      RECT 11.5480 4.5765 11.5740 5.6700 ;
      RECT 11.4400 4.5765 11.4660 5.6700 ;
      RECT 11.3320 4.5765 11.3580 5.6700 ;
      RECT 11.2240 4.5765 11.2500 5.6700 ;
      RECT 11.1160 4.5765 11.1420 5.6700 ;
      RECT 11.0080 4.5765 11.0340 5.6700 ;
      RECT 10.9000 4.5765 10.9260 5.6700 ;
      RECT 10.7920 4.5765 10.8180 5.6700 ;
      RECT 10.6840 4.5765 10.7100 5.6700 ;
      RECT 10.5760 4.5765 10.6020 5.6700 ;
      RECT 10.4680 4.5765 10.4940 5.6700 ;
      RECT 10.3600 4.5765 10.3860 5.6700 ;
      RECT 10.2520 4.5765 10.2780 5.6700 ;
      RECT 10.1440 4.5765 10.1700 5.6700 ;
      RECT 10.0360 4.5765 10.0620 5.6700 ;
      RECT 9.9280 4.5765 9.9540 5.6700 ;
      RECT 9.8200 4.5765 9.8460 5.6700 ;
      RECT 9.7120 4.5765 9.7380 5.6700 ;
      RECT 9.6040 4.5765 9.6300 5.6700 ;
      RECT 9.4960 4.5765 9.5220 5.6700 ;
      RECT 9.3880 4.5765 9.4140 5.6700 ;
      RECT 9.1750 4.5765 9.2520 5.6700 ;
      RECT 7.2820 4.5765 7.3590 5.6700 ;
      RECT 7.1200 4.5765 7.1460 5.6700 ;
      RECT 7.0120 4.5765 7.0380 5.6700 ;
      RECT 6.9040 4.5765 6.9300 5.6700 ;
      RECT 6.7960 4.5765 6.8220 5.6700 ;
      RECT 6.6880 4.5765 6.7140 5.6700 ;
      RECT 6.5800 4.5765 6.6060 5.6700 ;
      RECT 6.4720 4.5765 6.4980 5.6700 ;
      RECT 6.3640 4.5765 6.3900 5.6700 ;
      RECT 6.2560 4.5765 6.2820 5.6700 ;
      RECT 6.1480 4.5765 6.1740 5.6700 ;
      RECT 6.0400 4.5765 6.0660 5.6700 ;
      RECT 5.9320 4.5765 5.9580 5.6700 ;
      RECT 5.8240 4.5765 5.8500 5.6700 ;
      RECT 5.7160 4.5765 5.7420 5.6700 ;
      RECT 5.6080 4.5765 5.6340 5.6700 ;
      RECT 5.5000 4.5765 5.5260 5.6700 ;
      RECT 5.3920 4.5765 5.4180 5.6700 ;
      RECT 5.2840 4.5765 5.3100 5.6700 ;
      RECT 5.1760 4.5765 5.2020 5.6700 ;
      RECT 5.0680 4.5765 5.0940 5.6700 ;
      RECT 4.9600 4.5765 4.9860 5.6700 ;
      RECT 4.8520 4.5765 4.8780 5.6700 ;
      RECT 4.7440 4.5765 4.7700 5.6700 ;
      RECT 4.6360 4.5765 4.6620 5.6700 ;
      RECT 4.5280 4.5765 4.5540 5.6700 ;
      RECT 4.4200 4.5765 4.4460 5.6700 ;
      RECT 4.3120 4.5765 4.3380 5.6700 ;
      RECT 4.2040 4.5765 4.2300 5.6700 ;
      RECT 4.0960 4.5765 4.1220 5.6700 ;
      RECT 3.9880 4.5765 4.0140 5.6700 ;
      RECT 3.8800 4.5765 3.9060 5.6700 ;
      RECT 3.7720 4.5765 3.7980 5.6700 ;
      RECT 3.6640 4.5765 3.6900 5.6700 ;
      RECT 3.5560 4.5765 3.5820 5.6700 ;
      RECT 3.4480 4.5765 3.4740 5.6700 ;
      RECT 3.3400 4.5765 3.3660 5.6700 ;
      RECT 3.2320 4.5765 3.2580 5.6700 ;
      RECT 3.1240 4.5765 3.1500 5.6700 ;
      RECT 3.0160 4.5765 3.0420 5.6700 ;
      RECT 2.9080 4.5765 2.9340 5.6700 ;
      RECT 2.8000 4.5765 2.8260 5.6700 ;
      RECT 2.6920 4.5765 2.7180 5.6700 ;
      RECT 2.5840 4.5765 2.6100 5.6700 ;
      RECT 2.4760 4.5765 2.5020 5.6700 ;
      RECT 2.3680 4.5765 2.3940 5.6700 ;
      RECT 2.2600 4.5765 2.2860 5.6700 ;
      RECT 2.1520 4.5765 2.1780 5.6700 ;
      RECT 2.0440 4.5765 2.0700 5.6700 ;
      RECT 1.9360 4.5765 1.9620 5.6700 ;
      RECT 1.8280 4.5765 1.8540 5.6700 ;
      RECT 1.7200 4.5765 1.7460 5.6700 ;
      RECT 1.6120 4.5765 1.6380 5.6700 ;
      RECT 1.5040 4.5765 1.5300 5.6700 ;
      RECT 1.3960 4.5765 1.4220 5.6700 ;
      RECT 1.2880 4.5765 1.3140 5.6700 ;
      RECT 1.1800 4.5765 1.2060 5.6700 ;
      RECT 1.0720 4.5765 1.0980 5.6700 ;
      RECT 0.9640 4.5765 0.9900 5.6700 ;
      RECT 0.8560 4.5765 0.8820 5.6700 ;
      RECT 0.7480 4.5765 0.7740 5.6700 ;
      RECT 0.6400 4.5765 0.6660 5.6700 ;
      RECT 0.5320 4.5765 0.5580 5.6700 ;
      RECT 0.4240 4.5765 0.4500 5.6700 ;
      RECT 0.3160 4.5765 0.3420 5.6700 ;
      RECT 0.2080 4.5765 0.2340 5.6700 ;
      RECT 0.0050 4.5765 0.0900 5.6700 ;
      RECT 8.6410 5.6565 8.7690 6.7500 ;
      RECT 8.6270 6.3220 8.7690 6.6445 ;
      RECT 8.4790 6.0490 8.5410 6.7500 ;
      RECT 8.4650 6.3585 8.5410 6.5120 ;
      RECT 8.4790 5.6565 8.5050 6.7500 ;
      RECT 8.4790 5.7775 8.5190 6.0170 ;
      RECT 8.4790 5.6565 8.5410 5.7455 ;
      RECT 8.1820 6.1070 8.3880 6.7500 ;
      RECT 8.3620 5.6565 8.3880 6.7500 ;
      RECT 8.1820 6.3840 8.4020 6.6420 ;
      RECT 8.1820 5.6565 8.2800 6.7500 ;
      RECT 7.7650 5.6565 7.8480 6.7500 ;
      RECT 7.7650 5.7450 7.8620 6.6805 ;
      RECT 16.4440 5.6565 16.5290 6.7500 ;
      RECT 16.3000 5.6565 16.3260 6.7500 ;
      RECT 16.1920 5.6565 16.2180 6.7500 ;
      RECT 16.0840 5.6565 16.1100 6.7500 ;
      RECT 15.9760 5.6565 16.0020 6.7500 ;
      RECT 15.8680 5.6565 15.8940 6.7500 ;
      RECT 15.7600 5.6565 15.7860 6.7500 ;
      RECT 15.6520 5.6565 15.6780 6.7500 ;
      RECT 15.5440 5.6565 15.5700 6.7500 ;
      RECT 15.4360 5.6565 15.4620 6.7500 ;
      RECT 15.3280 5.6565 15.3540 6.7500 ;
      RECT 15.2200 5.6565 15.2460 6.7500 ;
      RECT 15.1120 5.6565 15.1380 6.7500 ;
      RECT 15.0040 5.6565 15.0300 6.7500 ;
      RECT 14.8960 5.6565 14.9220 6.7500 ;
      RECT 14.7880 5.6565 14.8140 6.7500 ;
      RECT 14.6800 5.6565 14.7060 6.7500 ;
      RECT 14.5720 5.6565 14.5980 6.7500 ;
      RECT 14.4640 5.6565 14.4900 6.7500 ;
      RECT 14.3560 5.6565 14.3820 6.7500 ;
      RECT 14.2480 5.6565 14.2740 6.7500 ;
      RECT 14.1400 5.6565 14.1660 6.7500 ;
      RECT 14.0320 5.6565 14.0580 6.7500 ;
      RECT 13.9240 5.6565 13.9500 6.7500 ;
      RECT 13.8160 5.6565 13.8420 6.7500 ;
      RECT 13.7080 5.6565 13.7340 6.7500 ;
      RECT 13.6000 5.6565 13.6260 6.7500 ;
      RECT 13.4920 5.6565 13.5180 6.7500 ;
      RECT 13.3840 5.6565 13.4100 6.7500 ;
      RECT 13.2760 5.6565 13.3020 6.7500 ;
      RECT 13.1680 5.6565 13.1940 6.7500 ;
      RECT 13.0600 5.6565 13.0860 6.7500 ;
      RECT 12.9520 5.6565 12.9780 6.7500 ;
      RECT 12.8440 5.6565 12.8700 6.7500 ;
      RECT 12.7360 5.6565 12.7620 6.7500 ;
      RECT 12.6280 5.6565 12.6540 6.7500 ;
      RECT 12.5200 5.6565 12.5460 6.7500 ;
      RECT 12.4120 5.6565 12.4380 6.7500 ;
      RECT 12.3040 5.6565 12.3300 6.7500 ;
      RECT 12.1960 5.6565 12.2220 6.7500 ;
      RECT 12.0880 5.6565 12.1140 6.7500 ;
      RECT 11.9800 5.6565 12.0060 6.7500 ;
      RECT 11.8720 5.6565 11.8980 6.7500 ;
      RECT 11.7640 5.6565 11.7900 6.7500 ;
      RECT 11.6560 5.6565 11.6820 6.7500 ;
      RECT 11.5480 5.6565 11.5740 6.7500 ;
      RECT 11.4400 5.6565 11.4660 6.7500 ;
      RECT 11.3320 5.6565 11.3580 6.7500 ;
      RECT 11.2240 5.6565 11.2500 6.7500 ;
      RECT 11.1160 5.6565 11.1420 6.7500 ;
      RECT 11.0080 5.6565 11.0340 6.7500 ;
      RECT 10.9000 5.6565 10.9260 6.7500 ;
      RECT 10.7920 5.6565 10.8180 6.7500 ;
      RECT 10.6840 5.6565 10.7100 6.7500 ;
      RECT 10.5760 5.6565 10.6020 6.7500 ;
      RECT 10.4680 5.6565 10.4940 6.7500 ;
      RECT 10.3600 5.6565 10.3860 6.7500 ;
      RECT 10.2520 5.6565 10.2780 6.7500 ;
      RECT 10.1440 5.6565 10.1700 6.7500 ;
      RECT 10.0360 5.6565 10.0620 6.7500 ;
      RECT 9.9280 5.6565 9.9540 6.7500 ;
      RECT 9.8200 5.6565 9.8460 6.7500 ;
      RECT 9.7120 5.6565 9.7380 6.7500 ;
      RECT 9.6040 5.6565 9.6300 6.7500 ;
      RECT 9.4960 5.6565 9.5220 6.7500 ;
      RECT 9.3880 5.6565 9.4140 6.7500 ;
      RECT 9.1750 5.6565 9.2520 6.7500 ;
      RECT 7.2820 5.6565 7.3590 6.7500 ;
      RECT 7.1200 5.6565 7.1460 6.7500 ;
      RECT 7.0120 5.6565 7.0380 6.7500 ;
      RECT 6.9040 5.6565 6.9300 6.7500 ;
      RECT 6.7960 5.6565 6.8220 6.7500 ;
      RECT 6.6880 5.6565 6.7140 6.7500 ;
      RECT 6.5800 5.6565 6.6060 6.7500 ;
      RECT 6.4720 5.6565 6.4980 6.7500 ;
      RECT 6.3640 5.6565 6.3900 6.7500 ;
      RECT 6.2560 5.6565 6.2820 6.7500 ;
      RECT 6.1480 5.6565 6.1740 6.7500 ;
      RECT 6.0400 5.6565 6.0660 6.7500 ;
      RECT 5.9320 5.6565 5.9580 6.7500 ;
      RECT 5.8240 5.6565 5.8500 6.7500 ;
      RECT 5.7160 5.6565 5.7420 6.7500 ;
      RECT 5.6080 5.6565 5.6340 6.7500 ;
      RECT 5.5000 5.6565 5.5260 6.7500 ;
      RECT 5.3920 5.6565 5.4180 6.7500 ;
      RECT 5.2840 5.6565 5.3100 6.7500 ;
      RECT 5.1760 5.6565 5.2020 6.7500 ;
      RECT 5.0680 5.6565 5.0940 6.7500 ;
      RECT 4.9600 5.6565 4.9860 6.7500 ;
      RECT 4.8520 5.6565 4.8780 6.7500 ;
      RECT 4.7440 5.6565 4.7700 6.7500 ;
      RECT 4.6360 5.6565 4.6620 6.7500 ;
      RECT 4.5280 5.6565 4.5540 6.7500 ;
      RECT 4.4200 5.6565 4.4460 6.7500 ;
      RECT 4.3120 5.6565 4.3380 6.7500 ;
      RECT 4.2040 5.6565 4.2300 6.7500 ;
      RECT 4.0960 5.6565 4.1220 6.7500 ;
      RECT 3.9880 5.6565 4.0140 6.7500 ;
      RECT 3.8800 5.6565 3.9060 6.7500 ;
      RECT 3.7720 5.6565 3.7980 6.7500 ;
      RECT 3.6640 5.6565 3.6900 6.7500 ;
      RECT 3.5560 5.6565 3.5820 6.7500 ;
      RECT 3.4480 5.6565 3.4740 6.7500 ;
      RECT 3.3400 5.6565 3.3660 6.7500 ;
      RECT 3.2320 5.6565 3.2580 6.7500 ;
      RECT 3.1240 5.6565 3.1500 6.7500 ;
      RECT 3.0160 5.6565 3.0420 6.7500 ;
      RECT 2.9080 5.6565 2.9340 6.7500 ;
      RECT 2.8000 5.6565 2.8260 6.7500 ;
      RECT 2.6920 5.6565 2.7180 6.7500 ;
      RECT 2.5840 5.6565 2.6100 6.7500 ;
      RECT 2.4760 5.6565 2.5020 6.7500 ;
      RECT 2.3680 5.6565 2.3940 6.7500 ;
      RECT 2.2600 5.6565 2.2860 6.7500 ;
      RECT 2.1520 5.6565 2.1780 6.7500 ;
      RECT 2.0440 5.6565 2.0700 6.7500 ;
      RECT 1.9360 5.6565 1.9620 6.7500 ;
      RECT 1.8280 5.6565 1.8540 6.7500 ;
      RECT 1.7200 5.6565 1.7460 6.7500 ;
      RECT 1.6120 5.6565 1.6380 6.7500 ;
      RECT 1.5040 5.6565 1.5300 6.7500 ;
      RECT 1.3960 5.6565 1.4220 6.7500 ;
      RECT 1.2880 5.6565 1.3140 6.7500 ;
      RECT 1.1800 5.6565 1.2060 6.7500 ;
      RECT 1.0720 5.6565 1.0980 6.7500 ;
      RECT 0.9640 5.6565 0.9900 6.7500 ;
      RECT 0.8560 5.6565 0.8820 6.7500 ;
      RECT 0.7480 5.6565 0.7740 6.7500 ;
      RECT 0.6400 5.6565 0.6660 6.7500 ;
      RECT 0.5320 5.6565 0.5580 6.7500 ;
      RECT 0.4240 5.6565 0.4500 6.7500 ;
      RECT 0.3160 5.6565 0.3420 6.7500 ;
      RECT 0.2080 5.6565 0.2340 6.7500 ;
      RECT 0.0050 5.6565 0.0900 6.7500 ;
      RECT 8.6410 6.7365 8.7690 7.8300 ;
      RECT 8.6270 7.4020 8.7690 7.7245 ;
      RECT 8.4790 7.1290 8.5410 7.8300 ;
      RECT 8.4650 7.4385 8.5410 7.5920 ;
      RECT 8.4790 6.7365 8.5050 7.8300 ;
      RECT 8.4790 6.8575 8.5190 7.0970 ;
      RECT 8.4790 6.7365 8.5410 6.8255 ;
      RECT 8.1820 7.1870 8.3880 7.8300 ;
      RECT 8.3620 6.7365 8.3880 7.8300 ;
      RECT 8.1820 7.4640 8.4020 7.7220 ;
      RECT 8.1820 6.7365 8.2800 7.8300 ;
      RECT 7.7650 6.7365 7.8480 7.8300 ;
      RECT 7.7650 6.8250 7.8620 7.7605 ;
      RECT 16.4440 6.7365 16.5290 7.8300 ;
      RECT 16.3000 6.7365 16.3260 7.8300 ;
      RECT 16.1920 6.7365 16.2180 7.8300 ;
      RECT 16.0840 6.7365 16.1100 7.8300 ;
      RECT 15.9760 6.7365 16.0020 7.8300 ;
      RECT 15.8680 6.7365 15.8940 7.8300 ;
      RECT 15.7600 6.7365 15.7860 7.8300 ;
      RECT 15.6520 6.7365 15.6780 7.8300 ;
      RECT 15.5440 6.7365 15.5700 7.8300 ;
      RECT 15.4360 6.7365 15.4620 7.8300 ;
      RECT 15.3280 6.7365 15.3540 7.8300 ;
      RECT 15.2200 6.7365 15.2460 7.8300 ;
      RECT 15.1120 6.7365 15.1380 7.8300 ;
      RECT 15.0040 6.7365 15.0300 7.8300 ;
      RECT 14.8960 6.7365 14.9220 7.8300 ;
      RECT 14.7880 6.7365 14.8140 7.8300 ;
      RECT 14.6800 6.7365 14.7060 7.8300 ;
      RECT 14.5720 6.7365 14.5980 7.8300 ;
      RECT 14.4640 6.7365 14.4900 7.8300 ;
      RECT 14.3560 6.7365 14.3820 7.8300 ;
      RECT 14.2480 6.7365 14.2740 7.8300 ;
      RECT 14.1400 6.7365 14.1660 7.8300 ;
      RECT 14.0320 6.7365 14.0580 7.8300 ;
      RECT 13.9240 6.7365 13.9500 7.8300 ;
      RECT 13.8160 6.7365 13.8420 7.8300 ;
      RECT 13.7080 6.7365 13.7340 7.8300 ;
      RECT 13.6000 6.7365 13.6260 7.8300 ;
      RECT 13.4920 6.7365 13.5180 7.8300 ;
      RECT 13.3840 6.7365 13.4100 7.8300 ;
      RECT 13.2760 6.7365 13.3020 7.8300 ;
      RECT 13.1680 6.7365 13.1940 7.8300 ;
      RECT 13.0600 6.7365 13.0860 7.8300 ;
      RECT 12.9520 6.7365 12.9780 7.8300 ;
      RECT 12.8440 6.7365 12.8700 7.8300 ;
      RECT 12.7360 6.7365 12.7620 7.8300 ;
      RECT 12.6280 6.7365 12.6540 7.8300 ;
      RECT 12.5200 6.7365 12.5460 7.8300 ;
      RECT 12.4120 6.7365 12.4380 7.8300 ;
      RECT 12.3040 6.7365 12.3300 7.8300 ;
      RECT 12.1960 6.7365 12.2220 7.8300 ;
      RECT 12.0880 6.7365 12.1140 7.8300 ;
      RECT 11.9800 6.7365 12.0060 7.8300 ;
      RECT 11.8720 6.7365 11.8980 7.8300 ;
      RECT 11.7640 6.7365 11.7900 7.8300 ;
      RECT 11.6560 6.7365 11.6820 7.8300 ;
      RECT 11.5480 6.7365 11.5740 7.8300 ;
      RECT 11.4400 6.7365 11.4660 7.8300 ;
      RECT 11.3320 6.7365 11.3580 7.8300 ;
      RECT 11.2240 6.7365 11.2500 7.8300 ;
      RECT 11.1160 6.7365 11.1420 7.8300 ;
      RECT 11.0080 6.7365 11.0340 7.8300 ;
      RECT 10.9000 6.7365 10.9260 7.8300 ;
      RECT 10.7920 6.7365 10.8180 7.8300 ;
      RECT 10.6840 6.7365 10.7100 7.8300 ;
      RECT 10.5760 6.7365 10.6020 7.8300 ;
      RECT 10.4680 6.7365 10.4940 7.8300 ;
      RECT 10.3600 6.7365 10.3860 7.8300 ;
      RECT 10.2520 6.7365 10.2780 7.8300 ;
      RECT 10.1440 6.7365 10.1700 7.8300 ;
      RECT 10.0360 6.7365 10.0620 7.8300 ;
      RECT 9.9280 6.7365 9.9540 7.8300 ;
      RECT 9.8200 6.7365 9.8460 7.8300 ;
      RECT 9.7120 6.7365 9.7380 7.8300 ;
      RECT 9.6040 6.7365 9.6300 7.8300 ;
      RECT 9.4960 6.7365 9.5220 7.8300 ;
      RECT 9.3880 6.7365 9.4140 7.8300 ;
      RECT 9.1750 6.7365 9.2520 7.8300 ;
      RECT 7.2820 6.7365 7.3590 7.8300 ;
      RECT 7.1200 6.7365 7.1460 7.8300 ;
      RECT 7.0120 6.7365 7.0380 7.8300 ;
      RECT 6.9040 6.7365 6.9300 7.8300 ;
      RECT 6.7960 6.7365 6.8220 7.8300 ;
      RECT 6.6880 6.7365 6.7140 7.8300 ;
      RECT 6.5800 6.7365 6.6060 7.8300 ;
      RECT 6.4720 6.7365 6.4980 7.8300 ;
      RECT 6.3640 6.7365 6.3900 7.8300 ;
      RECT 6.2560 6.7365 6.2820 7.8300 ;
      RECT 6.1480 6.7365 6.1740 7.8300 ;
      RECT 6.0400 6.7365 6.0660 7.8300 ;
      RECT 5.9320 6.7365 5.9580 7.8300 ;
      RECT 5.8240 6.7365 5.8500 7.8300 ;
      RECT 5.7160 6.7365 5.7420 7.8300 ;
      RECT 5.6080 6.7365 5.6340 7.8300 ;
      RECT 5.5000 6.7365 5.5260 7.8300 ;
      RECT 5.3920 6.7365 5.4180 7.8300 ;
      RECT 5.2840 6.7365 5.3100 7.8300 ;
      RECT 5.1760 6.7365 5.2020 7.8300 ;
      RECT 5.0680 6.7365 5.0940 7.8300 ;
      RECT 4.9600 6.7365 4.9860 7.8300 ;
      RECT 4.8520 6.7365 4.8780 7.8300 ;
      RECT 4.7440 6.7365 4.7700 7.8300 ;
      RECT 4.6360 6.7365 4.6620 7.8300 ;
      RECT 4.5280 6.7365 4.5540 7.8300 ;
      RECT 4.4200 6.7365 4.4460 7.8300 ;
      RECT 4.3120 6.7365 4.3380 7.8300 ;
      RECT 4.2040 6.7365 4.2300 7.8300 ;
      RECT 4.0960 6.7365 4.1220 7.8300 ;
      RECT 3.9880 6.7365 4.0140 7.8300 ;
      RECT 3.8800 6.7365 3.9060 7.8300 ;
      RECT 3.7720 6.7365 3.7980 7.8300 ;
      RECT 3.6640 6.7365 3.6900 7.8300 ;
      RECT 3.5560 6.7365 3.5820 7.8300 ;
      RECT 3.4480 6.7365 3.4740 7.8300 ;
      RECT 3.3400 6.7365 3.3660 7.8300 ;
      RECT 3.2320 6.7365 3.2580 7.8300 ;
      RECT 3.1240 6.7365 3.1500 7.8300 ;
      RECT 3.0160 6.7365 3.0420 7.8300 ;
      RECT 2.9080 6.7365 2.9340 7.8300 ;
      RECT 2.8000 6.7365 2.8260 7.8300 ;
      RECT 2.6920 6.7365 2.7180 7.8300 ;
      RECT 2.5840 6.7365 2.6100 7.8300 ;
      RECT 2.4760 6.7365 2.5020 7.8300 ;
      RECT 2.3680 6.7365 2.3940 7.8300 ;
      RECT 2.2600 6.7365 2.2860 7.8300 ;
      RECT 2.1520 6.7365 2.1780 7.8300 ;
      RECT 2.0440 6.7365 2.0700 7.8300 ;
      RECT 1.9360 6.7365 1.9620 7.8300 ;
      RECT 1.8280 6.7365 1.8540 7.8300 ;
      RECT 1.7200 6.7365 1.7460 7.8300 ;
      RECT 1.6120 6.7365 1.6380 7.8300 ;
      RECT 1.5040 6.7365 1.5300 7.8300 ;
      RECT 1.3960 6.7365 1.4220 7.8300 ;
      RECT 1.2880 6.7365 1.3140 7.8300 ;
      RECT 1.1800 6.7365 1.2060 7.8300 ;
      RECT 1.0720 6.7365 1.0980 7.8300 ;
      RECT 0.9640 6.7365 0.9900 7.8300 ;
      RECT 0.8560 6.7365 0.8820 7.8300 ;
      RECT 0.7480 6.7365 0.7740 7.8300 ;
      RECT 0.6400 6.7365 0.6660 7.8300 ;
      RECT 0.5320 6.7365 0.5580 7.8300 ;
      RECT 0.4240 6.7365 0.4500 7.8300 ;
      RECT 0.3160 6.7365 0.3420 7.8300 ;
      RECT 0.2080 6.7365 0.2340 7.8300 ;
      RECT 0.0050 6.7365 0.0900 7.8300 ;
      RECT 8.6410 7.8165 8.7690 8.9100 ;
      RECT 8.6270 8.4820 8.7690 8.8045 ;
      RECT 8.4790 8.2090 8.5410 8.9100 ;
      RECT 8.4650 8.5185 8.5410 8.6720 ;
      RECT 8.4790 7.8165 8.5050 8.9100 ;
      RECT 8.4790 7.9375 8.5190 8.1770 ;
      RECT 8.4790 7.8165 8.5410 7.9055 ;
      RECT 8.1820 8.2670 8.3880 8.9100 ;
      RECT 8.3620 7.8165 8.3880 8.9100 ;
      RECT 8.1820 8.5440 8.4020 8.8020 ;
      RECT 8.1820 7.8165 8.2800 8.9100 ;
      RECT 7.7650 7.8165 7.8480 8.9100 ;
      RECT 7.7650 7.9050 7.8620 8.8405 ;
      RECT 16.4440 7.8165 16.5290 8.9100 ;
      RECT 16.3000 7.8165 16.3260 8.9100 ;
      RECT 16.1920 7.8165 16.2180 8.9100 ;
      RECT 16.0840 7.8165 16.1100 8.9100 ;
      RECT 15.9760 7.8165 16.0020 8.9100 ;
      RECT 15.8680 7.8165 15.8940 8.9100 ;
      RECT 15.7600 7.8165 15.7860 8.9100 ;
      RECT 15.6520 7.8165 15.6780 8.9100 ;
      RECT 15.5440 7.8165 15.5700 8.9100 ;
      RECT 15.4360 7.8165 15.4620 8.9100 ;
      RECT 15.3280 7.8165 15.3540 8.9100 ;
      RECT 15.2200 7.8165 15.2460 8.9100 ;
      RECT 15.1120 7.8165 15.1380 8.9100 ;
      RECT 15.0040 7.8165 15.0300 8.9100 ;
      RECT 14.8960 7.8165 14.9220 8.9100 ;
      RECT 14.7880 7.8165 14.8140 8.9100 ;
      RECT 14.6800 7.8165 14.7060 8.9100 ;
      RECT 14.5720 7.8165 14.5980 8.9100 ;
      RECT 14.4640 7.8165 14.4900 8.9100 ;
      RECT 14.3560 7.8165 14.3820 8.9100 ;
      RECT 14.2480 7.8165 14.2740 8.9100 ;
      RECT 14.1400 7.8165 14.1660 8.9100 ;
      RECT 14.0320 7.8165 14.0580 8.9100 ;
      RECT 13.9240 7.8165 13.9500 8.9100 ;
      RECT 13.8160 7.8165 13.8420 8.9100 ;
      RECT 13.7080 7.8165 13.7340 8.9100 ;
      RECT 13.6000 7.8165 13.6260 8.9100 ;
      RECT 13.4920 7.8165 13.5180 8.9100 ;
      RECT 13.3840 7.8165 13.4100 8.9100 ;
      RECT 13.2760 7.8165 13.3020 8.9100 ;
      RECT 13.1680 7.8165 13.1940 8.9100 ;
      RECT 13.0600 7.8165 13.0860 8.9100 ;
      RECT 12.9520 7.8165 12.9780 8.9100 ;
      RECT 12.8440 7.8165 12.8700 8.9100 ;
      RECT 12.7360 7.8165 12.7620 8.9100 ;
      RECT 12.6280 7.8165 12.6540 8.9100 ;
      RECT 12.5200 7.8165 12.5460 8.9100 ;
      RECT 12.4120 7.8165 12.4380 8.9100 ;
      RECT 12.3040 7.8165 12.3300 8.9100 ;
      RECT 12.1960 7.8165 12.2220 8.9100 ;
      RECT 12.0880 7.8165 12.1140 8.9100 ;
      RECT 11.9800 7.8165 12.0060 8.9100 ;
      RECT 11.8720 7.8165 11.8980 8.9100 ;
      RECT 11.7640 7.8165 11.7900 8.9100 ;
      RECT 11.6560 7.8165 11.6820 8.9100 ;
      RECT 11.5480 7.8165 11.5740 8.9100 ;
      RECT 11.4400 7.8165 11.4660 8.9100 ;
      RECT 11.3320 7.8165 11.3580 8.9100 ;
      RECT 11.2240 7.8165 11.2500 8.9100 ;
      RECT 11.1160 7.8165 11.1420 8.9100 ;
      RECT 11.0080 7.8165 11.0340 8.9100 ;
      RECT 10.9000 7.8165 10.9260 8.9100 ;
      RECT 10.7920 7.8165 10.8180 8.9100 ;
      RECT 10.6840 7.8165 10.7100 8.9100 ;
      RECT 10.5760 7.8165 10.6020 8.9100 ;
      RECT 10.4680 7.8165 10.4940 8.9100 ;
      RECT 10.3600 7.8165 10.3860 8.9100 ;
      RECT 10.2520 7.8165 10.2780 8.9100 ;
      RECT 10.1440 7.8165 10.1700 8.9100 ;
      RECT 10.0360 7.8165 10.0620 8.9100 ;
      RECT 9.9280 7.8165 9.9540 8.9100 ;
      RECT 9.8200 7.8165 9.8460 8.9100 ;
      RECT 9.7120 7.8165 9.7380 8.9100 ;
      RECT 9.6040 7.8165 9.6300 8.9100 ;
      RECT 9.4960 7.8165 9.5220 8.9100 ;
      RECT 9.3880 7.8165 9.4140 8.9100 ;
      RECT 9.1750 7.8165 9.2520 8.9100 ;
      RECT 7.2820 7.8165 7.3590 8.9100 ;
      RECT 7.1200 7.8165 7.1460 8.9100 ;
      RECT 7.0120 7.8165 7.0380 8.9100 ;
      RECT 6.9040 7.8165 6.9300 8.9100 ;
      RECT 6.7960 7.8165 6.8220 8.9100 ;
      RECT 6.6880 7.8165 6.7140 8.9100 ;
      RECT 6.5800 7.8165 6.6060 8.9100 ;
      RECT 6.4720 7.8165 6.4980 8.9100 ;
      RECT 6.3640 7.8165 6.3900 8.9100 ;
      RECT 6.2560 7.8165 6.2820 8.9100 ;
      RECT 6.1480 7.8165 6.1740 8.9100 ;
      RECT 6.0400 7.8165 6.0660 8.9100 ;
      RECT 5.9320 7.8165 5.9580 8.9100 ;
      RECT 5.8240 7.8165 5.8500 8.9100 ;
      RECT 5.7160 7.8165 5.7420 8.9100 ;
      RECT 5.6080 7.8165 5.6340 8.9100 ;
      RECT 5.5000 7.8165 5.5260 8.9100 ;
      RECT 5.3920 7.8165 5.4180 8.9100 ;
      RECT 5.2840 7.8165 5.3100 8.9100 ;
      RECT 5.1760 7.8165 5.2020 8.9100 ;
      RECT 5.0680 7.8165 5.0940 8.9100 ;
      RECT 4.9600 7.8165 4.9860 8.9100 ;
      RECT 4.8520 7.8165 4.8780 8.9100 ;
      RECT 4.7440 7.8165 4.7700 8.9100 ;
      RECT 4.6360 7.8165 4.6620 8.9100 ;
      RECT 4.5280 7.8165 4.5540 8.9100 ;
      RECT 4.4200 7.8165 4.4460 8.9100 ;
      RECT 4.3120 7.8165 4.3380 8.9100 ;
      RECT 4.2040 7.8165 4.2300 8.9100 ;
      RECT 4.0960 7.8165 4.1220 8.9100 ;
      RECT 3.9880 7.8165 4.0140 8.9100 ;
      RECT 3.8800 7.8165 3.9060 8.9100 ;
      RECT 3.7720 7.8165 3.7980 8.9100 ;
      RECT 3.6640 7.8165 3.6900 8.9100 ;
      RECT 3.5560 7.8165 3.5820 8.9100 ;
      RECT 3.4480 7.8165 3.4740 8.9100 ;
      RECT 3.3400 7.8165 3.3660 8.9100 ;
      RECT 3.2320 7.8165 3.2580 8.9100 ;
      RECT 3.1240 7.8165 3.1500 8.9100 ;
      RECT 3.0160 7.8165 3.0420 8.9100 ;
      RECT 2.9080 7.8165 2.9340 8.9100 ;
      RECT 2.8000 7.8165 2.8260 8.9100 ;
      RECT 2.6920 7.8165 2.7180 8.9100 ;
      RECT 2.5840 7.8165 2.6100 8.9100 ;
      RECT 2.4760 7.8165 2.5020 8.9100 ;
      RECT 2.3680 7.8165 2.3940 8.9100 ;
      RECT 2.2600 7.8165 2.2860 8.9100 ;
      RECT 2.1520 7.8165 2.1780 8.9100 ;
      RECT 2.0440 7.8165 2.0700 8.9100 ;
      RECT 1.9360 7.8165 1.9620 8.9100 ;
      RECT 1.8280 7.8165 1.8540 8.9100 ;
      RECT 1.7200 7.8165 1.7460 8.9100 ;
      RECT 1.6120 7.8165 1.6380 8.9100 ;
      RECT 1.5040 7.8165 1.5300 8.9100 ;
      RECT 1.3960 7.8165 1.4220 8.9100 ;
      RECT 1.2880 7.8165 1.3140 8.9100 ;
      RECT 1.1800 7.8165 1.2060 8.9100 ;
      RECT 1.0720 7.8165 1.0980 8.9100 ;
      RECT 0.9640 7.8165 0.9900 8.9100 ;
      RECT 0.8560 7.8165 0.8820 8.9100 ;
      RECT 0.7480 7.8165 0.7740 8.9100 ;
      RECT 0.6400 7.8165 0.6660 8.9100 ;
      RECT 0.5320 7.8165 0.5580 8.9100 ;
      RECT 0.4240 7.8165 0.4500 8.9100 ;
      RECT 0.3160 7.8165 0.3420 8.9100 ;
      RECT 0.2080 7.8165 0.2340 8.9100 ;
      RECT 0.0050 7.8165 0.0900 8.9100 ;
      RECT 8.6410 8.8965 8.7690 9.9900 ;
      RECT 8.6270 9.5620 8.7690 9.8845 ;
      RECT 8.4790 9.2890 8.5410 9.9900 ;
      RECT 8.4650 9.5985 8.5410 9.7520 ;
      RECT 8.4790 8.8965 8.5050 9.9900 ;
      RECT 8.4790 9.0175 8.5190 9.2570 ;
      RECT 8.4790 8.8965 8.5410 8.9855 ;
      RECT 8.1820 9.3470 8.3880 9.9900 ;
      RECT 8.3620 8.8965 8.3880 9.9900 ;
      RECT 8.1820 9.6240 8.4020 9.8820 ;
      RECT 8.1820 8.8965 8.2800 9.9900 ;
      RECT 7.7650 8.8965 7.8480 9.9900 ;
      RECT 7.7650 8.9850 7.8620 9.9205 ;
      RECT 16.4440 8.8965 16.5290 9.9900 ;
      RECT 16.3000 8.8965 16.3260 9.9900 ;
      RECT 16.1920 8.8965 16.2180 9.9900 ;
      RECT 16.0840 8.8965 16.1100 9.9900 ;
      RECT 15.9760 8.8965 16.0020 9.9900 ;
      RECT 15.8680 8.8965 15.8940 9.9900 ;
      RECT 15.7600 8.8965 15.7860 9.9900 ;
      RECT 15.6520 8.8965 15.6780 9.9900 ;
      RECT 15.5440 8.8965 15.5700 9.9900 ;
      RECT 15.4360 8.8965 15.4620 9.9900 ;
      RECT 15.3280 8.8965 15.3540 9.9900 ;
      RECT 15.2200 8.8965 15.2460 9.9900 ;
      RECT 15.1120 8.8965 15.1380 9.9900 ;
      RECT 15.0040 8.8965 15.0300 9.9900 ;
      RECT 14.8960 8.8965 14.9220 9.9900 ;
      RECT 14.7880 8.8965 14.8140 9.9900 ;
      RECT 14.6800 8.8965 14.7060 9.9900 ;
      RECT 14.5720 8.8965 14.5980 9.9900 ;
      RECT 14.4640 8.8965 14.4900 9.9900 ;
      RECT 14.3560 8.8965 14.3820 9.9900 ;
      RECT 14.2480 8.8965 14.2740 9.9900 ;
      RECT 14.1400 8.8965 14.1660 9.9900 ;
      RECT 14.0320 8.8965 14.0580 9.9900 ;
      RECT 13.9240 8.8965 13.9500 9.9900 ;
      RECT 13.8160 8.8965 13.8420 9.9900 ;
      RECT 13.7080 8.8965 13.7340 9.9900 ;
      RECT 13.6000 8.8965 13.6260 9.9900 ;
      RECT 13.4920 8.8965 13.5180 9.9900 ;
      RECT 13.3840 8.8965 13.4100 9.9900 ;
      RECT 13.2760 8.8965 13.3020 9.9900 ;
      RECT 13.1680 8.8965 13.1940 9.9900 ;
      RECT 13.0600 8.8965 13.0860 9.9900 ;
      RECT 12.9520 8.8965 12.9780 9.9900 ;
      RECT 12.8440 8.8965 12.8700 9.9900 ;
      RECT 12.7360 8.8965 12.7620 9.9900 ;
      RECT 12.6280 8.8965 12.6540 9.9900 ;
      RECT 12.5200 8.8965 12.5460 9.9900 ;
      RECT 12.4120 8.8965 12.4380 9.9900 ;
      RECT 12.3040 8.8965 12.3300 9.9900 ;
      RECT 12.1960 8.8965 12.2220 9.9900 ;
      RECT 12.0880 8.8965 12.1140 9.9900 ;
      RECT 11.9800 8.8965 12.0060 9.9900 ;
      RECT 11.8720 8.8965 11.8980 9.9900 ;
      RECT 11.7640 8.8965 11.7900 9.9900 ;
      RECT 11.6560 8.8965 11.6820 9.9900 ;
      RECT 11.5480 8.8965 11.5740 9.9900 ;
      RECT 11.4400 8.8965 11.4660 9.9900 ;
      RECT 11.3320 8.8965 11.3580 9.9900 ;
      RECT 11.2240 8.8965 11.2500 9.9900 ;
      RECT 11.1160 8.8965 11.1420 9.9900 ;
      RECT 11.0080 8.8965 11.0340 9.9900 ;
      RECT 10.9000 8.8965 10.9260 9.9900 ;
      RECT 10.7920 8.8965 10.8180 9.9900 ;
      RECT 10.6840 8.8965 10.7100 9.9900 ;
      RECT 10.5760 8.8965 10.6020 9.9900 ;
      RECT 10.4680 8.8965 10.4940 9.9900 ;
      RECT 10.3600 8.8965 10.3860 9.9900 ;
      RECT 10.2520 8.8965 10.2780 9.9900 ;
      RECT 10.1440 8.8965 10.1700 9.9900 ;
      RECT 10.0360 8.8965 10.0620 9.9900 ;
      RECT 9.9280 8.8965 9.9540 9.9900 ;
      RECT 9.8200 8.8965 9.8460 9.9900 ;
      RECT 9.7120 8.8965 9.7380 9.9900 ;
      RECT 9.6040 8.8965 9.6300 9.9900 ;
      RECT 9.4960 8.8965 9.5220 9.9900 ;
      RECT 9.3880 8.8965 9.4140 9.9900 ;
      RECT 9.1750 8.8965 9.2520 9.9900 ;
      RECT 7.2820 8.8965 7.3590 9.9900 ;
      RECT 7.1200 8.8965 7.1460 9.9900 ;
      RECT 7.0120 8.8965 7.0380 9.9900 ;
      RECT 6.9040 8.8965 6.9300 9.9900 ;
      RECT 6.7960 8.8965 6.8220 9.9900 ;
      RECT 6.6880 8.8965 6.7140 9.9900 ;
      RECT 6.5800 8.8965 6.6060 9.9900 ;
      RECT 6.4720 8.8965 6.4980 9.9900 ;
      RECT 6.3640 8.8965 6.3900 9.9900 ;
      RECT 6.2560 8.8965 6.2820 9.9900 ;
      RECT 6.1480 8.8965 6.1740 9.9900 ;
      RECT 6.0400 8.8965 6.0660 9.9900 ;
      RECT 5.9320 8.8965 5.9580 9.9900 ;
      RECT 5.8240 8.8965 5.8500 9.9900 ;
      RECT 5.7160 8.8965 5.7420 9.9900 ;
      RECT 5.6080 8.8965 5.6340 9.9900 ;
      RECT 5.5000 8.8965 5.5260 9.9900 ;
      RECT 5.3920 8.8965 5.4180 9.9900 ;
      RECT 5.2840 8.8965 5.3100 9.9900 ;
      RECT 5.1760 8.8965 5.2020 9.9900 ;
      RECT 5.0680 8.8965 5.0940 9.9900 ;
      RECT 4.9600 8.8965 4.9860 9.9900 ;
      RECT 4.8520 8.8965 4.8780 9.9900 ;
      RECT 4.7440 8.8965 4.7700 9.9900 ;
      RECT 4.6360 8.8965 4.6620 9.9900 ;
      RECT 4.5280 8.8965 4.5540 9.9900 ;
      RECT 4.4200 8.8965 4.4460 9.9900 ;
      RECT 4.3120 8.8965 4.3380 9.9900 ;
      RECT 4.2040 8.8965 4.2300 9.9900 ;
      RECT 4.0960 8.8965 4.1220 9.9900 ;
      RECT 3.9880 8.8965 4.0140 9.9900 ;
      RECT 3.8800 8.8965 3.9060 9.9900 ;
      RECT 3.7720 8.8965 3.7980 9.9900 ;
      RECT 3.6640 8.8965 3.6900 9.9900 ;
      RECT 3.5560 8.8965 3.5820 9.9900 ;
      RECT 3.4480 8.8965 3.4740 9.9900 ;
      RECT 3.3400 8.8965 3.3660 9.9900 ;
      RECT 3.2320 8.8965 3.2580 9.9900 ;
      RECT 3.1240 8.8965 3.1500 9.9900 ;
      RECT 3.0160 8.8965 3.0420 9.9900 ;
      RECT 2.9080 8.8965 2.9340 9.9900 ;
      RECT 2.8000 8.8965 2.8260 9.9900 ;
      RECT 2.6920 8.8965 2.7180 9.9900 ;
      RECT 2.5840 8.8965 2.6100 9.9900 ;
      RECT 2.4760 8.8965 2.5020 9.9900 ;
      RECT 2.3680 8.8965 2.3940 9.9900 ;
      RECT 2.2600 8.8965 2.2860 9.9900 ;
      RECT 2.1520 8.8965 2.1780 9.9900 ;
      RECT 2.0440 8.8965 2.0700 9.9900 ;
      RECT 1.9360 8.8965 1.9620 9.9900 ;
      RECT 1.8280 8.8965 1.8540 9.9900 ;
      RECT 1.7200 8.8965 1.7460 9.9900 ;
      RECT 1.6120 8.8965 1.6380 9.9900 ;
      RECT 1.5040 8.8965 1.5300 9.9900 ;
      RECT 1.3960 8.8965 1.4220 9.9900 ;
      RECT 1.2880 8.8965 1.3140 9.9900 ;
      RECT 1.1800 8.8965 1.2060 9.9900 ;
      RECT 1.0720 8.8965 1.0980 9.9900 ;
      RECT 0.9640 8.8965 0.9900 9.9900 ;
      RECT 0.8560 8.8965 0.8820 9.9900 ;
      RECT 0.7480 8.8965 0.7740 9.9900 ;
      RECT 0.6400 8.8965 0.6660 9.9900 ;
      RECT 0.5320 8.8965 0.5580 9.9900 ;
      RECT 0.4240 8.8965 0.4500 9.9900 ;
      RECT 0.3160 8.8965 0.3420 9.9900 ;
      RECT 0.2080 8.8965 0.2340 9.9900 ;
      RECT 0.0050 8.8965 0.0900 9.9900 ;
      RECT 0.0000 18.1695 16.5240 18.6105 ;
      RECT 16.4390 9.9570 16.5240 18.6105 ;
      RECT 9.3830 11.4610 16.3210 18.6105 ;
      RECT 10.8410 9.9570 16.3210 18.6105 ;
      RECT 7.2230 18.1620 9.3010 18.6105 ;
      RECT 7.9970 18.1305 9.3010 18.6105 ;
      RECT 0.2030 11.2660 7.1410 18.6105 ;
      RECT 6.8450 9.9570 7.1410 18.6105 ;
      RECT 0.0000 9.9570 0.0850 18.6105 ;
      RECT 7.2230 11.5690 7.8430 18.6105 ;
      RECT 7.9970 18.1260 9.2650 18.6105 ;
      RECT 8.6450 11.3620 9.2650 18.6105 ;
      RECT 8.6360 17.8690 9.2650 18.6105 ;
      RECT 8.4740 17.8690 8.5360 18.6105 ;
      RECT 7.9970 17.8690 8.3830 18.6105 ;
      RECT 9.3830 13.7500 16.3350 18.1040 ;
      RECT 0.1890 13.7500 7.1410 18.1040 ;
      RECT 9.3690 13.7500 16.3350 18.0995 ;
      RECT 0.1890 13.7500 7.1550 18.0995 ;
      RECT 7.2090 13.7500 7.8430 18.0985 ;
      RECT 8.1770 10.6420 8.3470 18.6105 ;
      RECT 8.2850 9.9570 8.3470 18.6105 ;
      RECT 7.4930 10.3780 7.8790 17.7220 ;
      RECT 7.2090 17.6770 7.8930 17.7140 ;
      RECT 8.6310 16.6030 9.2650 17.7110 ;
      RECT 8.1630 17.4130 8.3470 17.6390 ;
      RECT 8.1770 16.8370 8.3610 17.0990 ;
      RECT 7.2090 16.6390 7.8930 17.0990 ;
      RECT 8.1630 16.0990 8.3470 16.5590 ;
      RECT 8.6310 14.0650 9.2650 16.3970 ;
      RECT 7.2090 14.7130 7.8930 15.8570 ;
      RECT 8.1770 14.4430 8.3610 15.7490 ;
      RECT 8.1630 15.0190 8.3610 15.4790 ;
      RECT 8.1630 11.7790 8.3470 14.9390 ;
      RECT 8.1630 11.7790 8.3610 14.3990 ;
      RECT 7.2090 14.1730 7.8930 14.3990 ;
      RECT 8.6450 11.3620 9.3010 13.7180 ;
      RECT 8.6310 11.2390 9.2470 13.0250 ;
      RECT 7.2230 12.2110 7.8930 12.5810 ;
      RECT 8.1770 11.5090 8.3610 11.6990 ;
      RECT 7.2770 11.4730 7.8930 11.6630 ;
      RECT 8.1630 11.3650 8.3470 11.5010 ;
      RECT 7.2770 10.7230 7.8790 17.7220 ;
      RECT 8.1770 11.2390 8.3610 11.4650 ;
      RECT 9.5450 11.2690 16.3210 18.6105 ;
      RECT 10.6250 11.2660 16.3210 18.6105 ;
      RECT 9.3830 9.9570 9.4630 18.6105 ;
      RECT 7.2230 10.6420 7.4110 11.4560 ;
      RECT 9.3830 9.9570 9.6790 11.3600 ;
      RECT 9.3830 11.0740 10.5430 11.3600 ;
      RECT 10.6250 9.9570 10.7590 18.6105 ;
      RECT 5.9810 10.8850 6.7630 18.6105 ;
      RECT 0.2030 9.9570 5.8990 18.6105 ;
      RECT 8.6450 10.7230 9.2470 18.6105 ;
      RECT 8.6810 10.1335 9.3010 11.2070 ;
      RECT 9.3830 11.0740 10.7590 11.1680 ;
      RECT 10.4090 9.9570 16.3210 11.1650 ;
      RECT 6.6290 9.9570 7.1410 11.1650 ;
      RECT 8.1630 11.0950 8.3610 11.1590 ;
      RECT 8.1630 10.9690 8.3470 11.1590 ;
      RECT 10.1930 10.6900 16.3210 11.1650 ;
      RECT 9.3830 10.7230 10.1110 11.3600 ;
      RECT 8.1770 10.6990 8.3610 10.9610 ;
      RECT 0.2030 10.6900 6.5470 11.1650 ;
      RECT 6.4130 9.9570 6.5470 18.6105 ;
      RECT 9.9770 9.9570 10.3270 10.8290 ;
      RECT 9.3830 10.6420 9.8950 11.3600 ;
      RECT 9.7610 9.9570 9.8950 18.6105 ;
      RECT 6.1970 10.6420 6.5470 18.6105 ;
      RECT 0.2030 9.9570 6.1150 11.1650 ;
      RECT 8.1770 9.9570 8.2030 18.6105 ;
      RECT 7.3130 9.9570 7.4110 18.6105 ;
      RECT 6.1970 9.9570 6.3310 18.6105 ;
      RECT 9.7610 9.9570 10.3270 10.5920 ;
      RECT 8.6450 9.9570 9.2470 10.5920 ;
      RECT 7.3130 9.9570 7.8430 10.5920 ;
      RECT 6.4130 9.9570 7.1410 10.5920 ;
      RECT 9.7610 9.9570 16.3210 10.5890 ;
      RECT 0.2030 9.9570 6.3310 10.5890 ;
      RECT 8.6310 10.4290 9.3010 10.5830 ;
      RECT 9.3830 9.9570 16.3210 10.3250 ;
      RECT 8.1770 9.9570 8.3470 10.3250 ;
      RECT 7.2230 9.9570 7.8430 10.3250 ;
      RECT 0.2030 9.9570 7.1410 10.3250 ;
      RECT 7.9970 9.9570 8.3470 10.2220 ;
      RECT 8.6360 9.9570 9.2470 10.1220 ;
      RECT 7.9970 9.9570 8.3830 10.1220 ;
      RECT 9.7650 9.9305 9.7830 18.6105 ;
      RECT 9.6570 9.9305 9.6750 18.6105 ;
      RECT 6.8490 9.9430 6.8670 18.6105 ;
      RECT 6.7410 9.9430 6.7590 18.6105 ;
      RECT 6.6330 9.9430 6.6510 18.6105 ;
      RECT 6.5250 9.9430 6.5430 18.6105 ;
      RECT 6.4170 9.9305 6.4350 18.6105 ;
      RECT 6.3090 9.9305 6.3270 18.6105 ;
      RECT 6.2010 9.9430 6.2190 18.6105 ;
      RECT 6.0930 9.9430 6.1110 18.6105 ;
      RECT 5.9850 9.9430 6.0030 18.6105 ;
      RECT 5.8770 9.9430 5.8950 18.6105 ;
      RECT 8.4740 9.9570 8.5360 10.1220 ;
        RECT 8.6410 18.1035 8.7690 19.1970 ;
        RECT 8.6270 18.7690 8.7690 19.0915 ;
        RECT 8.4790 18.4960 8.5410 19.1970 ;
        RECT 8.4650 18.8055 8.5410 18.9590 ;
        RECT 8.4790 18.1035 8.5050 19.1970 ;
        RECT 8.4790 18.2245 8.5190 18.4640 ;
        RECT 8.4790 18.1035 8.5410 18.1925 ;
        RECT 8.1820 18.5540 8.3880 19.1970 ;
        RECT 8.3620 18.1035 8.3880 19.1970 ;
        RECT 8.1820 18.8310 8.4020 19.0890 ;
        RECT 8.1820 18.1035 8.2800 19.1970 ;
        RECT 7.7650 18.1035 7.8480 19.1970 ;
        RECT 7.7650 18.1920 7.8620 19.1275 ;
        RECT 16.4440 18.1035 16.5290 19.1970 ;
        RECT 16.3000 18.1035 16.3260 19.1970 ;
        RECT 16.1920 18.1035 16.2180 19.1970 ;
        RECT 16.0840 18.1035 16.1100 19.1970 ;
        RECT 15.9760 18.1035 16.0020 19.1970 ;
        RECT 15.8680 18.1035 15.8940 19.1970 ;
        RECT 15.7600 18.1035 15.7860 19.1970 ;
        RECT 15.6520 18.1035 15.6780 19.1970 ;
        RECT 15.5440 18.1035 15.5700 19.1970 ;
        RECT 15.4360 18.1035 15.4620 19.1970 ;
        RECT 15.3280 18.1035 15.3540 19.1970 ;
        RECT 15.2200 18.1035 15.2460 19.1970 ;
        RECT 15.1120 18.1035 15.1380 19.1970 ;
        RECT 15.0040 18.1035 15.0300 19.1970 ;
        RECT 14.8960 18.1035 14.9220 19.1970 ;
        RECT 14.7880 18.1035 14.8140 19.1970 ;
        RECT 14.6800 18.1035 14.7060 19.1970 ;
        RECT 14.5720 18.1035 14.5980 19.1970 ;
        RECT 14.4640 18.1035 14.4900 19.1970 ;
        RECT 14.3560 18.1035 14.3820 19.1970 ;
        RECT 14.2480 18.1035 14.2740 19.1970 ;
        RECT 14.1400 18.1035 14.1660 19.1970 ;
        RECT 14.0320 18.1035 14.0580 19.1970 ;
        RECT 13.9240 18.1035 13.9500 19.1970 ;
        RECT 13.8160 18.1035 13.8420 19.1970 ;
        RECT 13.7080 18.1035 13.7340 19.1970 ;
        RECT 13.6000 18.1035 13.6260 19.1970 ;
        RECT 13.4920 18.1035 13.5180 19.1970 ;
        RECT 13.3840 18.1035 13.4100 19.1970 ;
        RECT 13.2760 18.1035 13.3020 19.1970 ;
        RECT 13.1680 18.1035 13.1940 19.1970 ;
        RECT 13.0600 18.1035 13.0860 19.1970 ;
        RECT 12.9520 18.1035 12.9780 19.1970 ;
        RECT 12.8440 18.1035 12.8700 19.1970 ;
        RECT 12.7360 18.1035 12.7620 19.1970 ;
        RECT 12.6280 18.1035 12.6540 19.1970 ;
        RECT 12.5200 18.1035 12.5460 19.1970 ;
        RECT 12.4120 18.1035 12.4380 19.1970 ;
        RECT 12.3040 18.1035 12.3300 19.1970 ;
        RECT 12.1960 18.1035 12.2220 19.1970 ;
        RECT 12.0880 18.1035 12.1140 19.1970 ;
        RECT 11.9800 18.1035 12.0060 19.1970 ;
        RECT 11.8720 18.1035 11.8980 19.1970 ;
        RECT 11.7640 18.1035 11.7900 19.1970 ;
        RECT 11.6560 18.1035 11.6820 19.1970 ;
        RECT 11.5480 18.1035 11.5740 19.1970 ;
        RECT 11.4400 18.1035 11.4660 19.1970 ;
        RECT 11.3320 18.1035 11.3580 19.1970 ;
        RECT 11.2240 18.1035 11.2500 19.1970 ;
        RECT 11.1160 18.1035 11.1420 19.1970 ;
        RECT 11.0080 18.1035 11.0340 19.1970 ;
        RECT 10.9000 18.1035 10.9260 19.1970 ;
        RECT 10.7920 18.1035 10.8180 19.1970 ;
        RECT 10.6840 18.1035 10.7100 19.1970 ;
        RECT 10.5760 18.1035 10.6020 19.1970 ;
        RECT 10.4680 18.1035 10.4940 19.1970 ;
        RECT 10.3600 18.1035 10.3860 19.1970 ;
        RECT 10.2520 18.1035 10.2780 19.1970 ;
        RECT 10.1440 18.1035 10.1700 19.1970 ;
        RECT 10.0360 18.1035 10.0620 19.1970 ;
        RECT 9.9280 18.1035 9.9540 19.1970 ;
        RECT 9.8200 18.1035 9.8460 19.1970 ;
        RECT 9.7120 18.1035 9.7380 19.1970 ;
        RECT 9.6040 18.1035 9.6300 19.1970 ;
        RECT 9.4960 18.1035 9.5220 19.1970 ;
        RECT 9.3880 18.1035 9.4140 19.1970 ;
        RECT 9.1750 18.1035 9.2520 19.1970 ;
        RECT 7.2820 18.1035 7.3590 19.1970 ;
        RECT 7.1200 18.1035 7.1460 19.1970 ;
        RECT 7.0120 18.1035 7.0380 19.1970 ;
        RECT 6.9040 18.1035 6.9300 19.1970 ;
        RECT 6.7960 18.1035 6.8220 19.1970 ;
        RECT 6.6880 18.1035 6.7140 19.1970 ;
        RECT 6.5800 18.1035 6.6060 19.1970 ;
        RECT 6.4720 18.1035 6.4980 19.1970 ;
        RECT 6.3640 18.1035 6.3900 19.1970 ;
        RECT 6.2560 18.1035 6.2820 19.1970 ;
        RECT 6.1480 18.1035 6.1740 19.1970 ;
        RECT 6.0400 18.1035 6.0660 19.1970 ;
        RECT 5.9320 18.1035 5.9580 19.1970 ;
        RECT 5.8240 18.1035 5.8500 19.1970 ;
        RECT 5.7160 18.1035 5.7420 19.1970 ;
        RECT 5.6080 18.1035 5.6340 19.1970 ;
        RECT 5.5000 18.1035 5.5260 19.1970 ;
        RECT 5.3920 18.1035 5.4180 19.1970 ;
        RECT 5.2840 18.1035 5.3100 19.1970 ;
        RECT 5.1760 18.1035 5.2020 19.1970 ;
        RECT 5.0680 18.1035 5.0940 19.1970 ;
        RECT 4.9600 18.1035 4.9860 19.1970 ;
        RECT 4.8520 18.1035 4.8780 19.1970 ;
        RECT 4.7440 18.1035 4.7700 19.1970 ;
        RECT 4.6360 18.1035 4.6620 19.1970 ;
        RECT 4.5280 18.1035 4.5540 19.1970 ;
        RECT 4.4200 18.1035 4.4460 19.1970 ;
        RECT 4.3120 18.1035 4.3380 19.1970 ;
        RECT 4.2040 18.1035 4.2300 19.1970 ;
        RECT 4.0960 18.1035 4.1220 19.1970 ;
        RECT 3.9880 18.1035 4.0140 19.1970 ;
        RECT 3.8800 18.1035 3.9060 19.1970 ;
        RECT 3.7720 18.1035 3.7980 19.1970 ;
        RECT 3.6640 18.1035 3.6900 19.1970 ;
        RECT 3.5560 18.1035 3.5820 19.1970 ;
        RECT 3.4480 18.1035 3.4740 19.1970 ;
        RECT 3.3400 18.1035 3.3660 19.1970 ;
        RECT 3.2320 18.1035 3.2580 19.1970 ;
        RECT 3.1240 18.1035 3.1500 19.1970 ;
        RECT 3.0160 18.1035 3.0420 19.1970 ;
        RECT 2.9080 18.1035 2.9340 19.1970 ;
        RECT 2.8000 18.1035 2.8260 19.1970 ;
        RECT 2.6920 18.1035 2.7180 19.1970 ;
        RECT 2.5840 18.1035 2.6100 19.1970 ;
        RECT 2.4760 18.1035 2.5020 19.1970 ;
        RECT 2.3680 18.1035 2.3940 19.1970 ;
        RECT 2.2600 18.1035 2.2860 19.1970 ;
        RECT 2.1520 18.1035 2.1780 19.1970 ;
        RECT 2.0440 18.1035 2.0700 19.1970 ;
        RECT 1.9360 18.1035 1.9620 19.1970 ;
        RECT 1.8280 18.1035 1.8540 19.1970 ;
        RECT 1.7200 18.1035 1.7460 19.1970 ;
        RECT 1.6120 18.1035 1.6380 19.1970 ;
        RECT 1.5040 18.1035 1.5300 19.1970 ;
        RECT 1.3960 18.1035 1.4220 19.1970 ;
        RECT 1.2880 18.1035 1.3140 19.1970 ;
        RECT 1.1800 18.1035 1.2060 19.1970 ;
        RECT 1.0720 18.1035 1.0980 19.1970 ;
        RECT 0.9640 18.1035 0.9900 19.1970 ;
        RECT 0.8560 18.1035 0.8820 19.1970 ;
        RECT 0.7480 18.1035 0.7740 19.1970 ;
        RECT 0.6400 18.1035 0.6660 19.1970 ;
        RECT 0.5320 18.1035 0.5580 19.1970 ;
        RECT 0.4240 18.1035 0.4500 19.1970 ;
        RECT 0.3160 18.1035 0.3420 19.1970 ;
        RECT 0.2080 18.1035 0.2340 19.1970 ;
        RECT 0.0050 18.1035 0.0900 19.1970 ;
        RECT 8.6410 19.1835 8.7690 20.2770 ;
        RECT 8.6270 19.8490 8.7690 20.1715 ;
        RECT 8.4790 19.5760 8.5410 20.2770 ;
        RECT 8.4650 19.8855 8.5410 20.0390 ;
        RECT 8.4790 19.1835 8.5050 20.2770 ;
        RECT 8.4790 19.3045 8.5190 19.5440 ;
        RECT 8.4790 19.1835 8.5410 19.2725 ;
        RECT 8.1820 19.6340 8.3880 20.2770 ;
        RECT 8.3620 19.1835 8.3880 20.2770 ;
        RECT 8.1820 19.9110 8.4020 20.1690 ;
        RECT 8.1820 19.1835 8.2800 20.2770 ;
        RECT 7.7650 19.1835 7.8480 20.2770 ;
        RECT 7.7650 19.2720 7.8620 20.2075 ;
        RECT 16.4440 19.1835 16.5290 20.2770 ;
        RECT 16.3000 19.1835 16.3260 20.2770 ;
        RECT 16.1920 19.1835 16.2180 20.2770 ;
        RECT 16.0840 19.1835 16.1100 20.2770 ;
        RECT 15.9760 19.1835 16.0020 20.2770 ;
        RECT 15.8680 19.1835 15.8940 20.2770 ;
        RECT 15.7600 19.1835 15.7860 20.2770 ;
        RECT 15.6520 19.1835 15.6780 20.2770 ;
        RECT 15.5440 19.1835 15.5700 20.2770 ;
        RECT 15.4360 19.1835 15.4620 20.2770 ;
        RECT 15.3280 19.1835 15.3540 20.2770 ;
        RECT 15.2200 19.1835 15.2460 20.2770 ;
        RECT 15.1120 19.1835 15.1380 20.2770 ;
        RECT 15.0040 19.1835 15.0300 20.2770 ;
        RECT 14.8960 19.1835 14.9220 20.2770 ;
        RECT 14.7880 19.1835 14.8140 20.2770 ;
        RECT 14.6800 19.1835 14.7060 20.2770 ;
        RECT 14.5720 19.1835 14.5980 20.2770 ;
        RECT 14.4640 19.1835 14.4900 20.2770 ;
        RECT 14.3560 19.1835 14.3820 20.2770 ;
        RECT 14.2480 19.1835 14.2740 20.2770 ;
        RECT 14.1400 19.1835 14.1660 20.2770 ;
        RECT 14.0320 19.1835 14.0580 20.2770 ;
        RECT 13.9240 19.1835 13.9500 20.2770 ;
        RECT 13.8160 19.1835 13.8420 20.2770 ;
        RECT 13.7080 19.1835 13.7340 20.2770 ;
        RECT 13.6000 19.1835 13.6260 20.2770 ;
        RECT 13.4920 19.1835 13.5180 20.2770 ;
        RECT 13.3840 19.1835 13.4100 20.2770 ;
        RECT 13.2760 19.1835 13.3020 20.2770 ;
        RECT 13.1680 19.1835 13.1940 20.2770 ;
        RECT 13.0600 19.1835 13.0860 20.2770 ;
        RECT 12.9520 19.1835 12.9780 20.2770 ;
        RECT 12.8440 19.1835 12.8700 20.2770 ;
        RECT 12.7360 19.1835 12.7620 20.2770 ;
        RECT 12.6280 19.1835 12.6540 20.2770 ;
        RECT 12.5200 19.1835 12.5460 20.2770 ;
        RECT 12.4120 19.1835 12.4380 20.2770 ;
        RECT 12.3040 19.1835 12.3300 20.2770 ;
        RECT 12.1960 19.1835 12.2220 20.2770 ;
        RECT 12.0880 19.1835 12.1140 20.2770 ;
        RECT 11.9800 19.1835 12.0060 20.2770 ;
        RECT 11.8720 19.1835 11.8980 20.2770 ;
        RECT 11.7640 19.1835 11.7900 20.2770 ;
        RECT 11.6560 19.1835 11.6820 20.2770 ;
        RECT 11.5480 19.1835 11.5740 20.2770 ;
        RECT 11.4400 19.1835 11.4660 20.2770 ;
        RECT 11.3320 19.1835 11.3580 20.2770 ;
        RECT 11.2240 19.1835 11.2500 20.2770 ;
        RECT 11.1160 19.1835 11.1420 20.2770 ;
        RECT 11.0080 19.1835 11.0340 20.2770 ;
        RECT 10.9000 19.1835 10.9260 20.2770 ;
        RECT 10.7920 19.1835 10.8180 20.2770 ;
        RECT 10.6840 19.1835 10.7100 20.2770 ;
        RECT 10.5760 19.1835 10.6020 20.2770 ;
        RECT 10.4680 19.1835 10.4940 20.2770 ;
        RECT 10.3600 19.1835 10.3860 20.2770 ;
        RECT 10.2520 19.1835 10.2780 20.2770 ;
        RECT 10.1440 19.1835 10.1700 20.2770 ;
        RECT 10.0360 19.1835 10.0620 20.2770 ;
        RECT 9.9280 19.1835 9.9540 20.2770 ;
        RECT 9.8200 19.1835 9.8460 20.2770 ;
        RECT 9.7120 19.1835 9.7380 20.2770 ;
        RECT 9.6040 19.1835 9.6300 20.2770 ;
        RECT 9.4960 19.1835 9.5220 20.2770 ;
        RECT 9.3880 19.1835 9.4140 20.2770 ;
        RECT 9.1750 19.1835 9.2520 20.2770 ;
        RECT 7.2820 19.1835 7.3590 20.2770 ;
        RECT 7.1200 19.1835 7.1460 20.2770 ;
        RECT 7.0120 19.1835 7.0380 20.2770 ;
        RECT 6.9040 19.1835 6.9300 20.2770 ;
        RECT 6.7960 19.1835 6.8220 20.2770 ;
        RECT 6.6880 19.1835 6.7140 20.2770 ;
        RECT 6.5800 19.1835 6.6060 20.2770 ;
        RECT 6.4720 19.1835 6.4980 20.2770 ;
        RECT 6.3640 19.1835 6.3900 20.2770 ;
        RECT 6.2560 19.1835 6.2820 20.2770 ;
        RECT 6.1480 19.1835 6.1740 20.2770 ;
        RECT 6.0400 19.1835 6.0660 20.2770 ;
        RECT 5.9320 19.1835 5.9580 20.2770 ;
        RECT 5.8240 19.1835 5.8500 20.2770 ;
        RECT 5.7160 19.1835 5.7420 20.2770 ;
        RECT 5.6080 19.1835 5.6340 20.2770 ;
        RECT 5.5000 19.1835 5.5260 20.2770 ;
        RECT 5.3920 19.1835 5.4180 20.2770 ;
        RECT 5.2840 19.1835 5.3100 20.2770 ;
        RECT 5.1760 19.1835 5.2020 20.2770 ;
        RECT 5.0680 19.1835 5.0940 20.2770 ;
        RECT 4.9600 19.1835 4.9860 20.2770 ;
        RECT 4.8520 19.1835 4.8780 20.2770 ;
        RECT 4.7440 19.1835 4.7700 20.2770 ;
        RECT 4.6360 19.1835 4.6620 20.2770 ;
        RECT 4.5280 19.1835 4.5540 20.2770 ;
        RECT 4.4200 19.1835 4.4460 20.2770 ;
        RECT 4.3120 19.1835 4.3380 20.2770 ;
        RECT 4.2040 19.1835 4.2300 20.2770 ;
        RECT 4.0960 19.1835 4.1220 20.2770 ;
        RECT 3.9880 19.1835 4.0140 20.2770 ;
        RECT 3.8800 19.1835 3.9060 20.2770 ;
        RECT 3.7720 19.1835 3.7980 20.2770 ;
        RECT 3.6640 19.1835 3.6900 20.2770 ;
        RECT 3.5560 19.1835 3.5820 20.2770 ;
        RECT 3.4480 19.1835 3.4740 20.2770 ;
        RECT 3.3400 19.1835 3.3660 20.2770 ;
        RECT 3.2320 19.1835 3.2580 20.2770 ;
        RECT 3.1240 19.1835 3.1500 20.2770 ;
        RECT 3.0160 19.1835 3.0420 20.2770 ;
        RECT 2.9080 19.1835 2.9340 20.2770 ;
        RECT 2.8000 19.1835 2.8260 20.2770 ;
        RECT 2.6920 19.1835 2.7180 20.2770 ;
        RECT 2.5840 19.1835 2.6100 20.2770 ;
        RECT 2.4760 19.1835 2.5020 20.2770 ;
        RECT 2.3680 19.1835 2.3940 20.2770 ;
        RECT 2.2600 19.1835 2.2860 20.2770 ;
        RECT 2.1520 19.1835 2.1780 20.2770 ;
        RECT 2.0440 19.1835 2.0700 20.2770 ;
        RECT 1.9360 19.1835 1.9620 20.2770 ;
        RECT 1.8280 19.1835 1.8540 20.2770 ;
        RECT 1.7200 19.1835 1.7460 20.2770 ;
        RECT 1.6120 19.1835 1.6380 20.2770 ;
        RECT 1.5040 19.1835 1.5300 20.2770 ;
        RECT 1.3960 19.1835 1.4220 20.2770 ;
        RECT 1.2880 19.1835 1.3140 20.2770 ;
        RECT 1.1800 19.1835 1.2060 20.2770 ;
        RECT 1.0720 19.1835 1.0980 20.2770 ;
        RECT 0.9640 19.1835 0.9900 20.2770 ;
        RECT 0.8560 19.1835 0.8820 20.2770 ;
        RECT 0.7480 19.1835 0.7740 20.2770 ;
        RECT 0.6400 19.1835 0.6660 20.2770 ;
        RECT 0.5320 19.1835 0.5580 20.2770 ;
        RECT 0.4240 19.1835 0.4500 20.2770 ;
        RECT 0.3160 19.1835 0.3420 20.2770 ;
        RECT 0.2080 19.1835 0.2340 20.2770 ;
        RECT 0.0050 19.1835 0.0900 20.2770 ;
        RECT 8.6410 20.2635 8.7690 21.3570 ;
        RECT 8.6270 20.9290 8.7690 21.2515 ;
        RECT 8.4790 20.6560 8.5410 21.3570 ;
        RECT 8.4650 20.9655 8.5410 21.1190 ;
        RECT 8.4790 20.2635 8.5050 21.3570 ;
        RECT 8.4790 20.3845 8.5190 20.6240 ;
        RECT 8.4790 20.2635 8.5410 20.3525 ;
        RECT 8.1820 20.7140 8.3880 21.3570 ;
        RECT 8.3620 20.2635 8.3880 21.3570 ;
        RECT 8.1820 20.9910 8.4020 21.2490 ;
        RECT 8.1820 20.2635 8.2800 21.3570 ;
        RECT 7.7650 20.2635 7.8480 21.3570 ;
        RECT 7.7650 20.3520 7.8620 21.2875 ;
        RECT 16.4440 20.2635 16.5290 21.3570 ;
        RECT 16.3000 20.2635 16.3260 21.3570 ;
        RECT 16.1920 20.2635 16.2180 21.3570 ;
        RECT 16.0840 20.2635 16.1100 21.3570 ;
        RECT 15.9760 20.2635 16.0020 21.3570 ;
        RECT 15.8680 20.2635 15.8940 21.3570 ;
        RECT 15.7600 20.2635 15.7860 21.3570 ;
        RECT 15.6520 20.2635 15.6780 21.3570 ;
        RECT 15.5440 20.2635 15.5700 21.3570 ;
        RECT 15.4360 20.2635 15.4620 21.3570 ;
        RECT 15.3280 20.2635 15.3540 21.3570 ;
        RECT 15.2200 20.2635 15.2460 21.3570 ;
        RECT 15.1120 20.2635 15.1380 21.3570 ;
        RECT 15.0040 20.2635 15.0300 21.3570 ;
        RECT 14.8960 20.2635 14.9220 21.3570 ;
        RECT 14.7880 20.2635 14.8140 21.3570 ;
        RECT 14.6800 20.2635 14.7060 21.3570 ;
        RECT 14.5720 20.2635 14.5980 21.3570 ;
        RECT 14.4640 20.2635 14.4900 21.3570 ;
        RECT 14.3560 20.2635 14.3820 21.3570 ;
        RECT 14.2480 20.2635 14.2740 21.3570 ;
        RECT 14.1400 20.2635 14.1660 21.3570 ;
        RECT 14.0320 20.2635 14.0580 21.3570 ;
        RECT 13.9240 20.2635 13.9500 21.3570 ;
        RECT 13.8160 20.2635 13.8420 21.3570 ;
        RECT 13.7080 20.2635 13.7340 21.3570 ;
        RECT 13.6000 20.2635 13.6260 21.3570 ;
        RECT 13.4920 20.2635 13.5180 21.3570 ;
        RECT 13.3840 20.2635 13.4100 21.3570 ;
        RECT 13.2760 20.2635 13.3020 21.3570 ;
        RECT 13.1680 20.2635 13.1940 21.3570 ;
        RECT 13.0600 20.2635 13.0860 21.3570 ;
        RECT 12.9520 20.2635 12.9780 21.3570 ;
        RECT 12.8440 20.2635 12.8700 21.3570 ;
        RECT 12.7360 20.2635 12.7620 21.3570 ;
        RECT 12.6280 20.2635 12.6540 21.3570 ;
        RECT 12.5200 20.2635 12.5460 21.3570 ;
        RECT 12.4120 20.2635 12.4380 21.3570 ;
        RECT 12.3040 20.2635 12.3300 21.3570 ;
        RECT 12.1960 20.2635 12.2220 21.3570 ;
        RECT 12.0880 20.2635 12.1140 21.3570 ;
        RECT 11.9800 20.2635 12.0060 21.3570 ;
        RECT 11.8720 20.2635 11.8980 21.3570 ;
        RECT 11.7640 20.2635 11.7900 21.3570 ;
        RECT 11.6560 20.2635 11.6820 21.3570 ;
        RECT 11.5480 20.2635 11.5740 21.3570 ;
        RECT 11.4400 20.2635 11.4660 21.3570 ;
        RECT 11.3320 20.2635 11.3580 21.3570 ;
        RECT 11.2240 20.2635 11.2500 21.3570 ;
        RECT 11.1160 20.2635 11.1420 21.3570 ;
        RECT 11.0080 20.2635 11.0340 21.3570 ;
        RECT 10.9000 20.2635 10.9260 21.3570 ;
        RECT 10.7920 20.2635 10.8180 21.3570 ;
        RECT 10.6840 20.2635 10.7100 21.3570 ;
        RECT 10.5760 20.2635 10.6020 21.3570 ;
        RECT 10.4680 20.2635 10.4940 21.3570 ;
        RECT 10.3600 20.2635 10.3860 21.3570 ;
        RECT 10.2520 20.2635 10.2780 21.3570 ;
        RECT 10.1440 20.2635 10.1700 21.3570 ;
        RECT 10.0360 20.2635 10.0620 21.3570 ;
        RECT 9.9280 20.2635 9.9540 21.3570 ;
        RECT 9.8200 20.2635 9.8460 21.3570 ;
        RECT 9.7120 20.2635 9.7380 21.3570 ;
        RECT 9.6040 20.2635 9.6300 21.3570 ;
        RECT 9.4960 20.2635 9.5220 21.3570 ;
        RECT 9.3880 20.2635 9.4140 21.3570 ;
        RECT 9.1750 20.2635 9.2520 21.3570 ;
        RECT 7.2820 20.2635 7.3590 21.3570 ;
        RECT 7.1200 20.2635 7.1460 21.3570 ;
        RECT 7.0120 20.2635 7.0380 21.3570 ;
        RECT 6.9040 20.2635 6.9300 21.3570 ;
        RECT 6.7960 20.2635 6.8220 21.3570 ;
        RECT 6.6880 20.2635 6.7140 21.3570 ;
        RECT 6.5800 20.2635 6.6060 21.3570 ;
        RECT 6.4720 20.2635 6.4980 21.3570 ;
        RECT 6.3640 20.2635 6.3900 21.3570 ;
        RECT 6.2560 20.2635 6.2820 21.3570 ;
        RECT 6.1480 20.2635 6.1740 21.3570 ;
        RECT 6.0400 20.2635 6.0660 21.3570 ;
        RECT 5.9320 20.2635 5.9580 21.3570 ;
        RECT 5.8240 20.2635 5.8500 21.3570 ;
        RECT 5.7160 20.2635 5.7420 21.3570 ;
        RECT 5.6080 20.2635 5.6340 21.3570 ;
        RECT 5.5000 20.2635 5.5260 21.3570 ;
        RECT 5.3920 20.2635 5.4180 21.3570 ;
        RECT 5.2840 20.2635 5.3100 21.3570 ;
        RECT 5.1760 20.2635 5.2020 21.3570 ;
        RECT 5.0680 20.2635 5.0940 21.3570 ;
        RECT 4.9600 20.2635 4.9860 21.3570 ;
        RECT 4.8520 20.2635 4.8780 21.3570 ;
        RECT 4.7440 20.2635 4.7700 21.3570 ;
        RECT 4.6360 20.2635 4.6620 21.3570 ;
        RECT 4.5280 20.2635 4.5540 21.3570 ;
        RECT 4.4200 20.2635 4.4460 21.3570 ;
        RECT 4.3120 20.2635 4.3380 21.3570 ;
        RECT 4.2040 20.2635 4.2300 21.3570 ;
        RECT 4.0960 20.2635 4.1220 21.3570 ;
        RECT 3.9880 20.2635 4.0140 21.3570 ;
        RECT 3.8800 20.2635 3.9060 21.3570 ;
        RECT 3.7720 20.2635 3.7980 21.3570 ;
        RECT 3.6640 20.2635 3.6900 21.3570 ;
        RECT 3.5560 20.2635 3.5820 21.3570 ;
        RECT 3.4480 20.2635 3.4740 21.3570 ;
        RECT 3.3400 20.2635 3.3660 21.3570 ;
        RECT 3.2320 20.2635 3.2580 21.3570 ;
        RECT 3.1240 20.2635 3.1500 21.3570 ;
        RECT 3.0160 20.2635 3.0420 21.3570 ;
        RECT 2.9080 20.2635 2.9340 21.3570 ;
        RECT 2.8000 20.2635 2.8260 21.3570 ;
        RECT 2.6920 20.2635 2.7180 21.3570 ;
        RECT 2.5840 20.2635 2.6100 21.3570 ;
        RECT 2.4760 20.2635 2.5020 21.3570 ;
        RECT 2.3680 20.2635 2.3940 21.3570 ;
        RECT 2.2600 20.2635 2.2860 21.3570 ;
        RECT 2.1520 20.2635 2.1780 21.3570 ;
        RECT 2.0440 20.2635 2.0700 21.3570 ;
        RECT 1.9360 20.2635 1.9620 21.3570 ;
        RECT 1.8280 20.2635 1.8540 21.3570 ;
        RECT 1.7200 20.2635 1.7460 21.3570 ;
        RECT 1.6120 20.2635 1.6380 21.3570 ;
        RECT 1.5040 20.2635 1.5300 21.3570 ;
        RECT 1.3960 20.2635 1.4220 21.3570 ;
        RECT 1.2880 20.2635 1.3140 21.3570 ;
        RECT 1.1800 20.2635 1.2060 21.3570 ;
        RECT 1.0720 20.2635 1.0980 21.3570 ;
        RECT 0.9640 20.2635 0.9900 21.3570 ;
        RECT 0.8560 20.2635 0.8820 21.3570 ;
        RECT 0.7480 20.2635 0.7740 21.3570 ;
        RECT 0.6400 20.2635 0.6660 21.3570 ;
        RECT 0.5320 20.2635 0.5580 21.3570 ;
        RECT 0.4240 20.2635 0.4500 21.3570 ;
        RECT 0.3160 20.2635 0.3420 21.3570 ;
        RECT 0.2080 20.2635 0.2340 21.3570 ;
        RECT 0.0050 20.2635 0.0900 21.3570 ;
        RECT 8.6410 21.3435 8.7690 22.4370 ;
        RECT 8.6270 22.0090 8.7690 22.3315 ;
        RECT 8.4790 21.7360 8.5410 22.4370 ;
        RECT 8.4650 22.0455 8.5410 22.1990 ;
        RECT 8.4790 21.3435 8.5050 22.4370 ;
        RECT 8.4790 21.4645 8.5190 21.7040 ;
        RECT 8.4790 21.3435 8.5410 21.4325 ;
        RECT 8.1820 21.7940 8.3880 22.4370 ;
        RECT 8.3620 21.3435 8.3880 22.4370 ;
        RECT 8.1820 22.0710 8.4020 22.3290 ;
        RECT 8.1820 21.3435 8.2800 22.4370 ;
        RECT 7.7650 21.3435 7.8480 22.4370 ;
        RECT 7.7650 21.4320 7.8620 22.3675 ;
        RECT 16.4440 21.3435 16.5290 22.4370 ;
        RECT 16.3000 21.3435 16.3260 22.4370 ;
        RECT 16.1920 21.3435 16.2180 22.4370 ;
        RECT 16.0840 21.3435 16.1100 22.4370 ;
        RECT 15.9760 21.3435 16.0020 22.4370 ;
        RECT 15.8680 21.3435 15.8940 22.4370 ;
        RECT 15.7600 21.3435 15.7860 22.4370 ;
        RECT 15.6520 21.3435 15.6780 22.4370 ;
        RECT 15.5440 21.3435 15.5700 22.4370 ;
        RECT 15.4360 21.3435 15.4620 22.4370 ;
        RECT 15.3280 21.3435 15.3540 22.4370 ;
        RECT 15.2200 21.3435 15.2460 22.4370 ;
        RECT 15.1120 21.3435 15.1380 22.4370 ;
        RECT 15.0040 21.3435 15.0300 22.4370 ;
        RECT 14.8960 21.3435 14.9220 22.4370 ;
        RECT 14.7880 21.3435 14.8140 22.4370 ;
        RECT 14.6800 21.3435 14.7060 22.4370 ;
        RECT 14.5720 21.3435 14.5980 22.4370 ;
        RECT 14.4640 21.3435 14.4900 22.4370 ;
        RECT 14.3560 21.3435 14.3820 22.4370 ;
        RECT 14.2480 21.3435 14.2740 22.4370 ;
        RECT 14.1400 21.3435 14.1660 22.4370 ;
        RECT 14.0320 21.3435 14.0580 22.4370 ;
        RECT 13.9240 21.3435 13.9500 22.4370 ;
        RECT 13.8160 21.3435 13.8420 22.4370 ;
        RECT 13.7080 21.3435 13.7340 22.4370 ;
        RECT 13.6000 21.3435 13.6260 22.4370 ;
        RECT 13.4920 21.3435 13.5180 22.4370 ;
        RECT 13.3840 21.3435 13.4100 22.4370 ;
        RECT 13.2760 21.3435 13.3020 22.4370 ;
        RECT 13.1680 21.3435 13.1940 22.4370 ;
        RECT 13.0600 21.3435 13.0860 22.4370 ;
        RECT 12.9520 21.3435 12.9780 22.4370 ;
        RECT 12.8440 21.3435 12.8700 22.4370 ;
        RECT 12.7360 21.3435 12.7620 22.4370 ;
        RECT 12.6280 21.3435 12.6540 22.4370 ;
        RECT 12.5200 21.3435 12.5460 22.4370 ;
        RECT 12.4120 21.3435 12.4380 22.4370 ;
        RECT 12.3040 21.3435 12.3300 22.4370 ;
        RECT 12.1960 21.3435 12.2220 22.4370 ;
        RECT 12.0880 21.3435 12.1140 22.4370 ;
        RECT 11.9800 21.3435 12.0060 22.4370 ;
        RECT 11.8720 21.3435 11.8980 22.4370 ;
        RECT 11.7640 21.3435 11.7900 22.4370 ;
        RECT 11.6560 21.3435 11.6820 22.4370 ;
        RECT 11.5480 21.3435 11.5740 22.4370 ;
        RECT 11.4400 21.3435 11.4660 22.4370 ;
        RECT 11.3320 21.3435 11.3580 22.4370 ;
        RECT 11.2240 21.3435 11.2500 22.4370 ;
        RECT 11.1160 21.3435 11.1420 22.4370 ;
        RECT 11.0080 21.3435 11.0340 22.4370 ;
        RECT 10.9000 21.3435 10.9260 22.4370 ;
        RECT 10.7920 21.3435 10.8180 22.4370 ;
        RECT 10.6840 21.3435 10.7100 22.4370 ;
        RECT 10.5760 21.3435 10.6020 22.4370 ;
        RECT 10.4680 21.3435 10.4940 22.4370 ;
        RECT 10.3600 21.3435 10.3860 22.4370 ;
        RECT 10.2520 21.3435 10.2780 22.4370 ;
        RECT 10.1440 21.3435 10.1700 22.4370 ;
        RECT 10.0360 21.3435 10.0620 22.4370 ;
        RECT 9.9280 21.3435 9.9540 22.4370 ;
        RECT 9.8200 21.3435 9.8460 22.4370 ;
        RECT 9.7120 21.3435 9.7380 22.4370 ;
        RECT 9.6040 21.3435 9.6300 22.4370 ;
        RECT 9.4960 21.3435 9.5220 22.4370 ;
        RECT 9.3880 21.3435 9.4140 22.4370 ;
        RECT 9.1750 21.3435 9.2520 22.4370 ;
        RECT 7.2820 21.3435 7.3590 22.4370 ;
        RECT 7.1200 21.3435 7.1460 22.4370 ;
        RECT 7.0120 21.3435 7.0380 22.4370 ;
        RECT 6.9040 21.3435 6.9300 22.4370 ;
        RECT 6.7960 21.3435 6.8220 22.4370 ;
        RECT 6.6880 21.3435 6.7140 22.4370 ;
        RECT 6.5800 21.3435 6.6060 22.4370 ;
        RECT 6.4720 21.3435 6.4980 22.4370 ;
        RECT 6.3640 21.3435 6.3900 22.4370 ;
        RECT 6.2560 21.3435 6.2820 22.4370 ;
        RECT 6.1480 21.3435 6.1740 22.4370 ;
        RECT 6.0400 21.3435 6.0660 22.4370 ;
        RECT 5.9320 21.3435 5.9580 22.4370 ;
        RECT 5.8240 21.3435 5.8500 22.4370 ;
        RECT 5.7160 21.3435 5.7420 22.4370 ;
        RECT 5.6080 21.3435 5.6340 22.4370 ;
        RECT 5.5000 21.3435 5.5260 22.4370 ;
        RECT 5.3920 21.3435 5.4180 22.4370 ;
        RECT 5.2840 21.3435 5.3100 22.4370 ;
        RECT 5.1760 21.3435 5.2020 22.4370 ;
        RECT 5.0680 21.3435 5.0940 22.4370 ;
        RECT 4.9600 21.3435 4.9860 22.4370 ;
        RECT 4.8520 21.3435 4.8780 22.4370 ;
        RECT 4.7440 21.3435 4.7700 22.4370 ;
        RECT 4.6360 21.3435 4.6620 22.4370 ;
        RECT 4.5280 21.3435 4.5540 22.4370 ;
        RECT 4.4200 21.3435 4.4460 22.4370 ;
        RECT 4.3120 21.3435 4.3380 22.4370 ;
        RECT 4.2040 21.3435 4.2300 22.4370 ;
        RECT 4.0960 21.3435 4.1220 22.4370 ;
        RECT 3.9880 21.3435 4.0140 22.4370 ;
        RECT 3.8800 21.3435 3.9060 22.4370 ;
        RECT 3.7720 21.3435 3.7980 22.4370 ;
        RECT 3.6640 21.3435 3.6900 22.4370 ;
        RECT 3.5560 21.3435 3.5820 22.4370 ;
        RECT 3.4480 21.3435 3.4740 22.4370 ;
        RECT 3.3400 21.3435 3.3660 22.4370 ;
        RECT 3.2320 21.3435 3.2580 22.4370 ;
        RECT 3.1240 21.3435 3.1500 22.4370 ;
        RECT 3.0160 21.3435 3.0420 22.4370 ;
        RECT 2.9080 21.3435 2.9340 22.4370 ;
        RECT 2.8000 21.3435 2.8260 22.4370 ;
        RECT 2.6920 21.3435 2.7180 22.4370 ;
        RECT 2.5840 21.3435 2.6100 22.4370 ;
        RECT 2.4760 21.3435 2.5020 22.4370 ;
        RECT 2.3680 21.3435 2.3940 22.4370 ;
        RECT 2.2600 21.3435 2.2860 22.4370 ;
        RECT 2.1520 21.3435 2.1780 22.4370 ;
        RECT 2.0440 21.3435 2.0700 22.4370 ;
        RECT 1.9360 21.3435 1.9620 22.4370 ;
        RECT 1.8280 21.3435 1.8540 22.4370 ;
        RECT 1.7200 21.3435 1.7460 22.4370 ;
        RECT 1.6120 21.3435 1.6380 22.4370 ;
        RECT 1.5040 21.3435 1.5300 22.4370 ;
        RECT 1.3960 21.3435 1.4220 22.4370 ;
        RECT 1.2880 21.3435 1.3140 22.4370 ;
        RECT 1.1800 21.3435 1.2060 22.4370 ;
        RECT 1.0720 21.3435 1.0980 22.4370 ;
        RECT 0.9640 21.3435 0.9900 22.4370 ;
        RECT 0.8560 21.3435 0.8820 22.4370 ;
        RECT 0.7480 21.3435 0.7740 22.4370 ;
        RECT 0.6400 21.3435 0.6660 22.4370 ;
        RECT 0.5320 21.3435 0.5580 22.4370 ;
        RECT 0.4240 21.3435 0.4500 22.4370 ;
        RECT 0.3160 21.3435 0.3420 22.4370 ;
        RECT 0.2080 21.3435 0.2340 22.4370 ;
        RECT 0.0050 21.3435 0.0900 22.4370 ;
        RECT 8.6410 22.4235 8.7690 23.5170 ;
        RECT 8.6270 23.0890 8.7690 23.4115 ;
        RECT 8.4790 22.8160 8.5410 23.5170 ;
        RECT 8.4650 23.1255 8.5410 23.2790 ;
        RECT 8.4790 22.4235 8.5050 23.5170 ;
        RECT 8.4790 22.5445 8.5190 22.7840 ;
        RECT 8.4790 22.4235 8.5410 22.5125 ;
        RECT 8.1820 22.8740 8.3880 23.5170 ;
        RECT 8.3620 22.4235 8.3880 23.5170 ;
        RECT 8.1820 23.1510 8.4020 23.4090 ;
        RECT 8.1820 22.4235 8.2800 23.5170 ;
        RECT 7.7650 22.4235 7.8480 23.5170 ;
        RECT 7.7650 22.5120 7.8620 23.4475 ;
        RECT 16.4440 22.4235 16.5290 23.5170 ;
        RECT 16.3000 22.4235 16.3260 23.5170 ;
        RECT 16.1920 22.4235 16.2180 23.5170 ;
        RECT 16.0840 22.4235 16.1100 23.5170 ;
        RECT 15.9760 22.4235 16.0020 23.5170 ;
        RECT 15.8680 22.4235 15.8940 23.5170 ;
        RECT 15.7600 22.4235 15.7860 23.5170 ;
        RECT 15.6520 22.4235 15.6780 23.5170 ;
        RECT 15.5440 22.4235 15.5700 23.5170 ;
        RECT 15.4360 22.4235 15.4620 23.5170 ;
        RECT 15.3280 22.4235 15.3540 23.5170 ;
        RECT 15.2200 22.4235 15.2460 23.5170 ;
        RECT 15.1120 22.4235 15.1380 23.5170 ;
        RECT 15.0040 22.4235 15.0300 23.5170 ;
        RECT 14.8960 22.4235 14.9220 23.5170 ;
        RECT 14.7880 22.4235 14.8140 23.5170 ;
        RECT 14.6800 22.4235 14.7060 23.5170 ;
        RECT 14.5720 22.4235 14.5980 23.5170 ;
        RECT 14.4640 22.4235 14.4900 23.5170 ;
        RECT 14.3560 22.4235 14.3820 23.5170 ;
        RECT 14.2480 22.4235 14.2740 23.5170 ;
        RECT 14.1400 22.4235 14.1660 23.5170 ;
        RECT 14.0320 22.4235 14.0580 23.5170 ;
        RECT 13.9240 22.4235 13.9500 23.5170 ;
        RECT 13.8160 22.4235 13.8420 23.5170 ;
        RECT 13.7080 22.4235 13.7340 23.5170 ;
        RECT 13.6000 22.4235 13.6260 23.5170 ;
        RECT 13.4920 22.4235 13.5180 23.5170 ;
        RECT 13.3840 22.4235 13.4100 23.5170 ;
        RECT 13.2760 22.4235 13.3020 23.5170 ;
        RECT 13.1680 22.4235 13.1940 23.5170 ;
        RECT 13.0600 22.4235 13.0860 23.5170 ;
        RECT 12.9520 22.4235 12.9780 23.5170 ;
        RECT 12.8440 22.4235 12.8700 23.5170 ;
        RECT 12.7360 22.4235 12.7620 23.5170 ;
        RECT 12.6280 22.4235 12.6540 23.5170 ;
        RECT 12.5200 22.4235 12.5460 23.5170 ;
        RECT 12.4120 22.4235 12.4380 23.5170 ;
        RECT 12.3040 22.4235 12.3300 23.5170 ;
        RECT 12.1960 22.4235 12.2220 23.5170 ;
        RECT 12.0880 22.4235 12.1140 23.5170 ;
        RECT 11.9800 22.4235 12.0060 23.5170 ;
        RECT 11.8720 22.4235 11.8980 23.5170 ;
        RECT 11.7640 22.4235 11.7900 23.5170 ;
        RECT 11.6560 22.4235 11.6820 23.5170 ;
        RECT 11.5480 22.4235 11.5740 23.5170 ;
        RECT 11.4400 22.4235 11.4660 23.5170 ;
        RECT 11.3320 22.4235 11.3580 23.5170 ;
        RECT 11.2240 22.4235 11.2500 23.5170 ;
        RECT 11.1160 22.4235 11.1420 23.5170 ;
        RECT 11.0080 22.4235 11.0340 23.5170 ;
        RECT 10.9000 22.4235 10.9260 23.5170 ;
        RECT 10.7920 22.4235 10.8180 23.5170 ;
        RECT 10.6840 22.4235 10.7100 23.5170 ;
        RECT 10.5760 22.4235 10.6020 23.5170 ;
        RECT 10.4680 22.4235 10.4940 23.5170 ;
        RECT 10.3600 22.4235 10.3860 23.5170 ;
        RECT 10.2520 22.4235 10.2780 23.5170 ;
        RECT 10.1440 22.4235 10.1700 23.5170 ;
        RECT 10.0360 22.4235 10.0620 23.5170 ;
        RECT 9.9280 22.4235 9.9540 23.5170 ;
        RECT 9.8200 22.4235 9.8460 23.5170 ;
        RECT 9.7120 22.4235 9.7380 23.5170 ;
        RECT 9.6040 22.4235 9.6300 23.5170 ;
        RECT 9.4960 22.4235 9.5220 23.5170 ;
        RECT 9.3880 22.4235 9.4140 23.5170 ;
        RECT 9.1750 22.4235 9.2520 23.5170 ;
        RECT 7.2820 22.4235 7.3590 23.5170 ;
        RECT 7.1200 22.4235 7.1460 23.5170 ;
        RECT 7.0120 22.4235 7.0380 23.5170 ;
        RECT 6.9040 22.4235 6.9300 23.5170 ;
        RECT 6.7960 22.4235 6.8220 23.5170 ;
        RECT 6.6880 22.4235 6.7140 23.5170 ;
        RECT 6.5800 22.4235 6.6060 23.5170 ;
        RECT 6.4720 22.4235 6.4980 23.5170 ;
        RECT 6.3640 22.4235 6.3900 23.5170 ;
        RECT 6.2560 22.4235 6.2820 23.5170 ;
        RECT 6.1480 22.4235 6.1740 23.5170 ;
        RECT 6.0400 22.4235 6.0660 23.5170 ;
        RECT 5.9320 22.4235 5.9580 23.5170 ;
        RECT 5.8240 22.4235 5.8500 23.5170 ;
        RECT 5.7160 22.4235 5.7420 23.5170 ;
        RECT 5.6080 22.4235 5.6340 23.5170 ;
        RECT 5.5000 22.4235 5.5260 23.5170 ;
        RECT 5.3920 22.4235 5.4180 23.5170 ;
        RECT 5.2840 22.4235 5.3100 23.5170 ;
        RECT 5.1760 22.4235 5.2020 23.5170 ;
        RECT 5.0680 22.4235 5.0940 23.5170 ;
        RECT 4.9600 22.4235 4.9860 23.5170 ;
        RECT 4.8520 22.4235 4.8780 23.5170 ;
        RECT 4.7440 22.4235 4.7700 23.5170 ;
        RECT 4.6360 22.4235 4.6620 23.5170 ;
        RECT 4.5280 22.4235 4.5540 23.5170 ;
        RECT 4.4200 22.4235 4.4460 23.5170 ;
        RECT 4.3120 22.4235 4.3380 23.5170 ;
        RECT 4.2040 22.4235 4.2300 23.5170 ;
        RECT 4.0960 22.4235 4.1220 23.5170 ;
        RECT 3.9880 22.4235 4.0140 23.5170 ;
        RECT 3.8800 22.4235 3.9060 23.5170 ;
        RECT 3.7720 22.4235 3.7980 23.5170 ;
        RECT 3.6640 22.4235 3.6900 23.5170 ;
        RECT 3.5560 22.4235 3.5820 23.5170 ;
        RECT 3.4480 22.4235 3.4740 23.5170 ;
        RECT 3.3400 22.4235 3.3660 23.5170 ;
        RECT 3.2320 22.4235 3.2580 23.5170 ;
        RECT 3.1240 22.4235 3.1500 23.5170 ;
        RECT 3.0160 22.4235 3.0420 23.5170 ;
        RECT 2.9080 22.4235 2.9340 23.5170 ;
        RECT 2.8000 22.4235 2.8260 23.5170 ;
        RECT 2.6920 22.4235 2.7180 23.5170 ;
        RECT 2.5840 22.4235 2.6100 23.5170 ;
        RECT 2.4760 22.4235 2.5020 23.5170 ;
        RECT 2.3680 22.4235 2.3940 23.5170 ;
        RECT 2.2600 22.4235 2.2860 23.5170 ;
        RECT 2.1520 22.4235 2.1780 23.5170 ;
        RECT 2.0440 22.4235 2.0700 23.5170 ;
        RECT 1.9360 22.4235 1.9620 23.5170 ;
        RECT 1.8280 22.4235 1.8540 23.5170 ;
        RECT 1.7200 22.4235 1.7460 23.5170 ;
        RECT 1.6120 22.4235 1.6380 23.5170 ;
        RECT 1.5040 22.4235 1.5300 23.5170 ;
        RECT 1.3960 22.4235 1.4220 23.5170 ;
        RECT 1.2880 22.4235 1.3140 23.5170 ;
        RECT 1.1800 22.4235 1.2060 23.5170 ;
        RECT 1.0720 22.4235 1.0980 23.5170 ;
        RECT 0.9640 22.4235 0.9900 23.5170 ;
        RECT 0.8560 22.4235 0.8820 23.5170 ;
        RECT 0.7480 22.4235 0.7740 23.5170 ;
        RECT 0.6400 22.4235 0.6660 23.5170 ;
        RECT 0.5320 22.4235 0.5580 23.5170 ;
        RECT 0.4240 22.4235 0.4500 23.5170 ;
        RECT 0.3160 22.4235 0.3420 23.5170 ;
        RECT 0.2080 22.4235 0.2340 23.5170 ;
        RECT 0.0050 22.4235 0.0900 23.5170 ;
        RECT 8.6410 23.5035 8.7690 24.5970 ;
        RECT 8.6270 24.1690 8.7690 24.4915 ;
        RECT 8.4790 23.8960 8.5410 24.5970 ;
        RECT 8.4650 24.2055 8.5410 24.3590 ;
        RECT 8.4790 23.5035 8.5050 24.5970 ;
        RECT 8.4790 23.6245 8.5190 23.8640 ;
        RECT 8.4790 23.5035 8.5410 23.5925 ;
        RECT 8.1820 23.9540 8.3880 24.5970 ;
        RECT 8.3620 23.5035 8.3880 24.5970 ;
        RECT 8.1820 24.2310 8.4020 24.4890 ;
        RECT 8.1820 23.5035 8.2800 24.5970 ;
        RECT 7.7650 23.5035 7.8480 24.5970 ;
        RECT 7.7650 23.5920 7.8620 24.5275 ;
        RECT 16.4440 23.5035 16.5290 24.5970 ;
        RECT 16.3000 23.5035 16.3260 24.5970 ;
        RECT 16.1920 23.5035 16.2180 24.5970 ;
        RECT 16.0840 23.5035 16.1100 24.5970 ;
        RECT 15.9760 23.5035 16.0020 24.5970 ;
        RECT 15.8680 23.5035 15.8940 24.5970 ;
        RECT 15.7600 23.5035 15.7860 24.5970 ;
        RECT 15.6520 23.5035 15.6780 24.5970 ;
        RECT 15.5440 23.5035 15.5700 24.5970 ;
        RECT 15.4360 23.5035 15.4620 24.5970 ;
        RECT 15.3280 23.5035 15.3540 24.5970 ;
        RECT 15.2200 23.5035 15.2460 24.5970 ;
        RECT 15.1120 23.5035 15.1380 24.5970 ;
        RECT 15.0040 23.5035 15.0300 24.5970 ;
        RECT 14.8960 23.5035 14.9220 24.5970 ;
        RECT 14.7880 23.5035 14.8140 24.5970 ;
        RECT 14.6800 23.5035 14.7060 24.5970 ;
        RECT 14.5720 23.5035 14.5980 24.5970 ;
        RECT 14.4640 23.5035 14.4900 24.5970 ;
        RECT 14.3560 23.5035 14.3820 24.5970 ;
        RECT 14.2480 23.5035 14.2740 24.5970 ;
        RECT 14.1400 23.5035 14.1660 24.5970 ;
        RECT 14.0320 23.5035 14.0580 24.5970 ;
        RECT 13.9240 23.5035 13.9500 24.5970 ;
        RECT 13.8160 23.5035 13.8420 24.5970 ;
        RECT 13.7080 23.5035 13.7340 24.5970 ;
        RECT 13.6000 23.5035 13.6260 24.5970 ;
        RECT 13.4920 23.5035 13.5180 24.5970 ;
        RECT 13.3840 23.5035 13.4100 24.5970 ;
        RECT 13.2760 23.5035 13.3020 24.5970 ;
        RECT 13.1680 23.5035 13.1940 24.5970 ;
        RECT 13.0600 23.5035 13.0860 24.5970 ;
        RECT 12.9520 23.5035 12.9780 24.5970 ;
        RECT 12.8440 23.5035 12.8700 24.5970 ;
        RECT 12.7360 23.5035 12.7620 24.5970 ;
        RECT 12.6280 23.5035 12.6540 24.5970 ;
        RECT 12.5200 23.5035 12.5460 24.5970 ;
        RECT 12.4120 23.5035 12.4380 24.5970 ;
        RECT 12.3040 23.5035 12.3300 24.5970 ;
        RECT 12.1960 23.5035 12.2220 24.5970 ;
        RECT 12.0880 23.5035 12.1140 24.5970 ;
        RECT 11.9800 23.5035 12.0060 24.5970 ;
        RECT 11.8720 23.5035 11.8980 24.5970 ;
        RECT 11.7640 23.5035 11.7900 24.5970 ;
        RECT 11.6560 23.5035 11.6820 24.5970 ;
        RECT 11.5480 23.5035 11.5740 24.5970 ;
        RECT 11.4400 23.5035 11.4660 24.5970 ;
        RECT 11.3320 23.5035 11.3580 24.5970 ;
        RECT 11.2240 23.5035 11.2500 24.5970 ;
        RECT 11.1160 23.5035 11.1420 24.5970 ;
        RECT 11.0080 23.5035 11.0340 24.5970 ;
        RECT 10.9000 23.5035 10.9260 24.5970 ;
        RECT 10.7920 23.5035 10.8180 24.5970 ;
        RECT 10.6840 23.5035 10.7100 24.5970 ;
        RECT 10.5760 23.5035 10.6020 24.5970 ;
        RECT 10.4680 23.5035 10.4940 24.5970 ;
        RECT 10.3600 23.5035 10.3860 24.5970 ;
        RECT 10.2520 23.5035 10.2780 24.5970 ;
        RECT 10.1440 23.5035 10.1700 24.5970 ;
        RECT 10.0360 23.5035 10.0620 24.5970 ;
        RECT 9.9280 23.5035 9.9540 24.5970 ;
        RECT 9.8200 23.5035 9.8460 24.5970 ;
        RECT 9.7120 23.5035 9.7380 24.5970 ;
        RECT 9.6040 23.5035 9.6300 24.5970 ;
        RECT 9.4960 23.5035 9.5220 24.5970 ;
        RECT 9.3880 23.5035 9.4140 24.5970 ;
        RECT 9.1750 23.5035 9.2520 24.5970 ;
        RECT 7.2820 23.5035 7.3590 24.5970 ;
        RECT 7.1200 23.5035 7.1460 24.5970 ;
        RECT 7.0120 23.5035 7.0380 24.5970 ;
        RECT 6.9040 23.5035 6.9300 24.5970 ;
        RECT 6.7960 23.5035 6.8220 24.5970 ;
        RECT 6.6880 23.5035 6.7140 24.5970 ;
        RECT 6.5800 23.5035 6.6060 24.5970 ;
        RECT 6.4720 23.5035 6.4980 24.5970 ;
        RECT 6.3640 23.5035 6.3900 24.5970 ;
        RECT 6.2560 23.5035 6.2820 24.5970 ;
        RECT 6.1480 23.5035 6.1740 24.5970 ;
        RECT 6.0400 23.5035 6.0660 24.5970 ;
        RECT 5.9320 23.5035 5.9580 24.5970 ;
        RECT 5.8240 23.5035 5.8500 24.5970 ;
        RECT 5.7160 23.5035 5.7420 24.5970 ;
        RECT 5.6080 23.5035 5.6340 24.5970 ;
        RECT 5.5000 23.5035 5.5260 24.5970 ;
        RECT 5.3920 23.5035 5.4180 24.5970 ;
        RECT 5.2840 23.5035 5.3100 24.5970 ;
        RECT 5.1760 23.5035 5.2020 24.5970 ;
        RECT 5.0680 23.5035 5.0940 24.5970 ;
        RECT 4.9600 23.5035 4.9860 24.5970 ;
        RECT 4.8520 23.5035 4.8780 24.5970 ;
        RECT 4.7440 23.5035 4.7700 24.5970 ;
        RECT 4.6360 23.5035 4.6620 24.5970 ;
        RECT 4.5280 23.5035 4.5540 24.5970 ;
        RECT 4.4200 23.5035 4.4460 24.5970 ;
        RECT 4.3120 23.5035 4.3380 24.5970 ;
        RECT 4.2040 23.5035 4.2300 24.5970 ;
        RECT 4.0960 23.5035 4.1220 24.5970 ;
        RECT 3.9880 23.5035 4.0140 24.5970 ;
        RECT 3.8800 23.5035 3.9060 24.5970 ;
        RECT 3.7720 23.5035 3.7980 24.5970 ;
        RECT 3.6640 23.5035 3.6900 24.5970 ;
        RECT 3.5560 23.5035 3.5820 24.5970 ;
        RECT 3.4480 23.5035 3.4740 24.5970 ;
        RECT 3.3400 23.5035 3.3660 24.5970 ;
        RECT 3.2320 23.5035 3.2580 24.5970 ;
        RECT 3.1240 23.5035 3.1500 24.5970 ;
        RECT 3.0160 23.5035 3.0420 24.5970 ;
        RECT 2.9080 23.5035 2.9340 24.5970 ;
        RECT 2.8000 23.5035 2.8260 24.5970 ;
        RECT 2.6920 23.5035 2.7180 24.5970 ;
        RECT 2.5840 23.5035 2.6100 24.5970 ;
        RECT 2.4760 23.5035 2.5020 24.5970 ;
        RECT 2.3680 23.5035 2.3940 24.5970 ;
        RECT 2.2600 23.5035 2.2860 24.5970 ;
        RECT 2.1520 23.5035 2.1780 24.5970 ;
        RECT 2.0440 23.5035 2.0700 24.5970 ;
        RECT 1.9360 23.5035 1.9620 24.5970 ;
        RECT 1.8280 23.5035 1.8540 24.5970 ;
        RECT 1.7200 23.5035 1.7460 24.5970 ;
        RECT 1.6120 23.5035 1.6380 24.5970 ;
        RECT 1.5040 23.5035 1.5300 24.5970 ;
        RECT 1.3960 23.5035 1.4220 24.5970 ;
        RECT 1.2880 23.5035 1.3140 24.5970 ;
        RECT 1.1800 23.5035 1.2060 24.5970 ;
        RECT 1.0720 23.5035 1.0980 24.5970 ;
        RECT 0.9640 23.5035 0.9900 24.5970 ;
        RECT 0.8560 23.5035 0.8820 24.5970 ;
        RECT 0.7480 23.5035 0.7740 24.5970 ;
        RECT 0.6400 23.5035 0.6660 24.5970 ;
        RECT 0.5320 23.5035 0.5580 24.5970 ;
        RECT 0.4240 23.5035 0.4500 24.5970 ;
        RECT 0.3160 23.5035 0.3420 24.5970 ;
        RECT 0.2080 23.5035 0.2340 24.5970 ;
        RECT 0.0050 23.5035 0.0900 24.5970 ;
        RECT 8.6410 24.5835 8.7690 25.6770 ;
        RECT 8.6270 25.2490 8.7690 25.5715 ;
        RECT 8.4790 24.9760 8.5410 25.6770 ;
        RECT 8.4650 25.2855 8.5410 25.4390 ;
        RECT 8.4790 24.5835 8.5050 25.6770 ;
        RECT 8.4790 24.7045 8.5190 24.9440 ;
        RECT 8.4790 24.5835 8.5410 24.6725 ;
        RECT 8.1820 25.0340 8.3880 25.6770 ;
        RECT 8.3620 24.5835 8.3880 25.6770 ;
        RECT 8.1820 25.3110 8.4020 25.5690 ;
        RECT 8.1820 24.5835 8.2800 25.6770 ;
        RECT 7.7650 24.5835 7.8480 25.6770 ;
        RECT 7.7650 24.6720 7.8620 25.6075 ;
        RECT 16.4440 24.5835 16.5290 25.6770 ;
        RECT 16.3000 24.5835 16.3260 25.6770 ;
        RECT 16.1920 24.5835 16.2180 25.6770 ;
        RECT 16.0840 24.5835 16.1100 25.6770 ;
        RECT 15.9760 24.5835 16.0020 25.6770 ;
        RECT 15.8680 24.5835 15.8940 25.6770 ;
        RECT 15.7600 24.5835 15.7860 25.6770 ;
        RECT 15.6520 24.5835 15.6780 25.6770 ;
        RECT 15.5440 24.5835 15.5700 25.6770 ;
        RECT 15.4360 24.5835 15.4620 25.6770 ;
        RECT 15.3280 24.5835 15.3540 25.6770 ;
        RECT 15.2200 24.5835 15.2460 25.6770 ;
        RECT 15.1120 24.5835 15.1380 25.6770 ;
        RECT 15.0040 24.5835 15.0300 25.6770 ;
        RECT 14.8960 24.5835 14.9220 25.6770 ;
        RECT 14.7880 24.5835 14.8140 25.6770 ;
        RECT 14.6800 24.5835 14.7060 25.6770 ;
        RECT 14.5720 24.5835 14.5980 25.6770 ;
        RECT 14.4640 24.5835 14.4900 25.6770 ;
        RECT 14.3560 24.5835 14.3820 25.6770 ;
        RECT 14.2480 24.5835 14.2740 25.6770 ;
        RECT 14.1400 24.5835 14.1660 25.6770 ;
        RECT 14.0320 24.5835 14.0580 25.6770 ;
        RECT 13.9240 24.5835 13.9500 25.6770 ;
        RECT 13.8160 24.5835 13.8420 25.6770 ;
        RECT 13.7080 24.5835 13.7340 25.6770 ;
        RECT 13.6000 24.5835 13.6260 25.6770 ;
        RECT 13.4920 24.5835 13.5180 25.6770 ;
        RECT 13.3840 24.5835 13.4100 25.6770 ;
        RECT 13.2760 24.5835 13.3020 25.6770 ;
        RECT 13.1680 24.5835 13.1940 25.6770 ;
        RECT 13.0600 24.5835 13.0860 25.6770 ;
        RECT 12.9520 24.5835 12.9780 25.6770 ;
        RECT 12.8440 24.5835 12.8700 25.6770 ;
        RECT 12.7360 24.5835 12.7620 25.6770 ;
        RECT 12.6280 24.5835 12.6540 25.6770 ;
        RECT 12.5200 24.5835 12.5460 25.6770 ;
        RECT 12.4120 24.5835 12.4380 25.6770 ;
        RECT 12.3040 24.5835 12.3300 25.6770 ;
        RECT 12.1960 24.5835 12.2220 25.6770 ;
        RECT 12.0880 24.5835 12.1140 25.6770 ;
        RECT 11.9800 24.5835 12.0060 25.6770 ;
        RECT 11.8720 24.5835 11.8980 25.6770 ;
        RECT 11.7640 24.5835 11.7900 25.6770 ;
        RECT 11.6560 24.5835 11.6820 25.6770 ;
        RECT 11.5480 24.5835 11.5740 25.6770 ;
        RECT 11.4400 24.5835 11.4660 25.6770 ;
        RECT 11.3320 24.5835 11.3580 25.6770 ;
        RECT 11.2240 24.5835 11.2500 25.6770 ;
        RECT 11.1160 24.5835 11.1420 25.6770 ;
        RECT 11.0080 24.5835 11.0340 25.6770 ;
        RECT 10.9000 24.5835 10.9260 25.6770 ;
        RECT 10.7920 24.5835 10.8180 25.6770 ;
        RECT 10.6840 24.5835 10.7100 25.6770 ;
        RECT 10.5760 24.5835 10.6020 25.6770 ;
        RECT 10.4680 24.5835 10.4940 25.6770 ;
        RECT 10.3600 24.5835 10.3860 25.6770 ;
        RECT 10.2520 24.5835 10.2780 25.6770 ;
        RECT 10.1440 24.5835 10.1700 25.6770 ;
        RECT 10.0360 24.5835 10.0620 25.6770 ;
        RECT 9.9280 24.5835 9.9540 25.6770 ;
        RECT 9.8200 24.5835 9.8460 25.6770 ;
        RECT 9.7120 24.5835 9.7380 25.6770 ;
        RECT 9.6040 24.5835 9.6300 25.6770 ;
        RECT 9.4960 24.5835 9.5220 25.6770 ;
        RECT 9.3880 24.5835 9.4140 25.6770 ;
        RECT 9.1750 24.5835 9.2520 25.6770 ;
        RECT 7.2820 24.5835 7.3590 25.6770 ;
        RECT 7.1200 24.5835 7.1460 25.6770 ;
        RECT 7.0120 24.5835 7.0380 25.6770 ;
        RECT 6.9040 24.5835 6.9300 25.6770 ;
        RECT 6.7960 24.5835 6.8220 25.6770 ;
        RECT 6.6880 24.5835 6.7140 25.6770 ;
        RECT 6.5800 24.5835 6.6060 25.6770 ;
        RECT 6.4720 24.5835 6.4980 25.6770 ;
        RECT 6.3640 24.5835 6.3900 25.6770 ;
        RECT 6.2560 24.5835 6.2820 25.6770 ;
        RECT 6.1480 24.5835 6.1740 25.6770 ;
        RECT 6.0400 24.5835 6.0660 25.6770 ;
        RECT 5.9320 24.5835 5.9580 25.6770 ;
        RECT 5.8240 24.5835 5.8500 25.6770 ;
        RECT 5.7160 24.5835 5.7420 25.6770 ;
        RECT 5.6080 24.5835 5.6340 25.6770 ;
        RECT 5.5000 24.5835 5.5260 25.6770 ;
        RECT 5.3920 24.5835 5.4180 25.6770 ;
        RECT 5.2840 24.5835 5.3100 25.6770 ;
        RECT 5.1760 24.5835 5.2020 25.6770 ;
        RECT 5.0680 24.5835 5.0940 25.6770 ;
        RECT 4.9600 24.5835 4.9860 25.6770 ;
        RECT 4.8520 24.5835 4.8780 25.6770 ;
        RECT 4.7440 24.5835 4.7700 25.6770 ;
        RECT 4.6360 24.5835 4.6620 25.6770 ;
        RECT 4.5280 24.5835 4.5540 25.6770 ;
        RECT 4.4200 24.5835 4.4460 25.6770 ;
        RECT 4.3120 24.5835 4.3380 25.6770 ;
        RECT 4.2040 24.5835 4.2300 25.6770 ;
        RECT 4.0960 24.5835 4.1220 25.6770 ;
        RECT 3.9880 24.5835 4.0140 25.6770 ;
        RECT 3.8800 24.5835 3.9060 25.6770 ;
        RECT 3.7720 24.5835 3.7980 25.6770 ;
        RECT 3.6640 24.5835 3.6900 25.6770 ;
        RECT 3.5560 24.5835 3.5820 25.6770 ;
        RECT 3.4480 24.5835 3.4740 25.6770 ;
        RECT 3.3400 24.5835 3.3660 25.6770 ;
        RECT 3.2320 24.5835 3.2580 25.6770 ;
        RECT 3.1240 24.5835 3.1500 25.6770 ;
        RECT 3.0160 24.5835 3.0420 25.6770 ;
        RECT 2.9080 24.5835 2.9340 25.6770 ;
        RECT 2.8000 24.5835 2.8260 25.6770 ;
        RECT 2.6920 24.5835 2.7180 25.6770 ;
        RECT 2.5840 24.5835 2.6100 25.6770 ;
        RECT 2.4760 24.5835 2.5020 25.6770 ;
        RECT 2.3680 24.5835 2.3940 25.6770 ;
        RECT 2.2600 24.5835 2.2860 25.6770 ;
        RECT 2.1520 24.5835 2.1780 25.6770 ;
        RECT 2.0440 24.5835 2.0700 25.6770 ;
        RECT 1.9360 24.5835 1.9620 25.6770 ;
        RECT 1.8280 24.5835 1.8540 25.6770 ;
        RECT 1.7200 24.5835 1.7460 25.6770 ;
        RECT 1.6120 24.5835 1.6380 25.6770 ;
        RECT 1.5040 24.5835 1.5300 25.6770 ;
        RECT 1.3960 24.5835 1.4220 25.6770 ;
        RECT 1.2880 24.5835 1.3140 25.6770 ;
        RECT 1.1800 24.5835 1.2060 25.6770 ;
        RECT 1.0720 24.5835 1.0980 25.6770 ;
        RECT 0.9640 24.5835 0.9900 25.6770 ;
        RECT 0.8560 24.5835 0.8820 25.6770 ;
        RECT 0.7480 24.5835 0.7740 25.6770 ;
        RECT 0.6400 24.5835 0.6660 25.6770 ;
        RECT 0.5320 24.5835 0.5580 25.6770 ;
        RECT 0.4240 24.5835 0.4500 25.6770 ;
        RECT 0.3160 24.5835 0.3420 25.6770 ;
        RECT 0.2080 24.5835 0.2340 25.6770 ;
        RECT 0.0050 24.5835 0.0900 25.6770 ;
        RECT 8.6410 25.6635 8.7690 26.7570 ;
        RECT 8.6270 26.3290 8.7690 26.6515 ;
        RECT 8.4790 26.0560 8.5410 26.7570 ;
        RECT 8.4650 26.3655 8.5410 26.5190 ;
        RECT 8.4790 25.6635 8.5050 26.7570 ;
        RECT 8.4790 25.7845 8.5190 26.0240 ;
        RECT 8.4790 25.6635 8.5410 25.7525 ;
        RECT 8.1820 26.1140 8.3880 26.7570 ;
        RECT 8.3620 25.6635 8.3880 26.7570 ;
        RECT 8.1820 26.3910 8.4020 26.6490 ;
        RECT 8.1820 25.6635 8.2800 26.7570 ;
        RECT 7.7650 25.6635 7.8480 26.7570 ;
        RECT 7.7650 25.7520 7.8620 26.6875 ;
        RECT 16.4440 25.6635 16.5290 26.7570 ;
        RECT 16.3000 25.6635 16.3260 26.7570 ;
        RECT 16.1920 25.6635 16.2180 26.7570 ;
        RECT 16.0840 25.6635 16.1100 26.7570 ;
        RECT 15.9760 25.6635 16.0020 26.7570 ;
        RECT 15.8680 25.6635 15.8940 26.7570 ;
        RECT 15.7600 25.6635 15.7860 26.7570 ;
        RECT 15.6520 25.6635 15.6780 26.7570 ;
        RECT 15.5440 25.6635 15.5700 26.7570 ;
        RECT 15.4360 25.6635 15.4620 26.7570 ;
        RECT 15.3280 25.6635 15.3540 26.7570 ;
        RECT 15.2200 25.6635 15.2460 26.7570 ;
        RECT 15.1120 25.6635 15.1380 26.7570 ;
        RECT 15.0040 25.6635 15.0300 26.7570 ;
        RECT 14.8960 25.6635 14.9220 26.7570 ;
        RECT 14.7880 25.6635 14.8140 26.7570 ;
        RECT 14.6800 25.6635 14.7060 26.7570 ;
        RECT 14.5720 25.6635 14.5980 26.7570 ;
        RECT 14.4640 25.6635 14.4900 26.7570 ;
        RECT 14.3560 25.6635 14.3820 26.7570 ;
        RECT 14.2480 25.6635 14.2740 26.7570 ;
        RECT 14.1400 25.6635 14.1660 26.7570 ;
        RECT 14.0320 25.6635 14.0580 26.7570 ;
        RECT 13.9240 25.6635 13.9500 26.7570 ;
        RECT 13.8160 25.6635 13.8420 26.7570 ;
        RECT 13.7080 25.6635 13.7340 26.7570 ;
        RECT 13.6000 25.6635 13.6260 26.7570 ;
        RECT 13.4920 25.6635 13.5180 26.7570 ;
        RECT 13.3840 25.6635 13.4100 26.7570 ;
        RECT 13.2760 25.6635 13.3020 26.7570 ;
        RECT 13.1680 25.6635 13.1940 26.7570 ;
        RECT 13.0600 25.6635 13.0860 26.7570 ;
        RECT 12.9520 25.6635 12.9780 26.7570 ;
        RECT 12.8440 25.6635 12.8700 26.7570 ;
        RECT 12.7360 25.6635 12.7620 26.7570 ;
        RECT 12.6280 25.6635 12.6540 26.7570 ;
        RECT 12.5200 25.6635 12.5460 26.7570 ;
        RECT 12.4120 25.6635 12.4380 26.7570 ;
        RECT 12.3040 25.6635 12.3300 26.7570 ;
        RECT 12.1960 25.6635 12.2220 26.7570 ;
        RECT 12.0880 25.6635 12.1140 26.7570 ;
        RECT 11.9800 25.6635 12.0060 26.7570 ;
        RECT 11.8720 25.6635 11.8980 26.7570 ;
        RECT 11.7640 25.6635 11.7900 26.7570 ;
        RECT 11.6560 25.6635 11.6820 26.7570 ;
        RECT 11.5480 25.6635 11.5740 26.7570 ;
        RECT 11.4400 25.6635 11.4660 26.7570 ;
        RECT 11.3320 25.6635 11.3580 26.7570 ;
        RECT 11.2240 25.6635 11.2500 26.7570 ;
        RECT 11.1160 25.6635 11.1420 26.7570 ;
        RECT 11.0080 25.6635 11.0340 26.7570 ;
        RECT 10.9000 25.6635 10.9260 26.7570 ;
        RECT 10.7920 25.6635 10.8180 26.7570 ;
        RECT 10.6840 25.6635 10.7100 26.7570 ;
        RECT 10.5760 25.6635 10.6020 26.7570 ;
        RECT 10.4680 25.6635 10.4940 26.7570 ;
        RECT 10.3600 25.6635 10.3860 26.7570 ;
        RECT 10.2520 25.6635 10.2780 26.7570 ;
        RECT 10.1440 25.6635 10.1700 26.7570 ;
        RECT 10.0360 25.6635 10.0620 26.7570 ;
        RECT 9.9280 25.6635 9.9540 26.7570 ;
        RECT 9.8200 25.6635 9.8460 26.7570 ;
        RECT 9.7120 25.6635 9.7380 26.7570 ;
        RECT 9.6040 25.6635 9.6300 26.7570 ;
        RECT 9.4960 25.6635 9.5220 26.7570 ;
        RECT 9.3880 25.6635 9.4140 26.7570 ;
        RECT 9.1750 25.6635 9.2520 26.7570 ;
        RECT 7.2820 25.6635 7.3590 26.7570 ;
        RECT 7.1200 25.6635 7.1460 26.7570 ;
        RECT 7.0120 25.6635 7.0380 26.7570 ;
        RECT 6.9040 25.6635 6.9300 26.7570 ;
        RECT 6.7960 25.6635 6.8220 26.7570 ;
        RECT 6.6880 25.6635 6.7140 26.7570 ;
        RECT 6.5800 25.6635 6.6060 26.7570 ;
        RECT 6.4720 25.6635 6.4980 26.7570 ;
        RECT 6.3640 25.6635 6.3900 26.7570 ;
        RECT 6.2560 25.6635 6.2820 26.7570 ;
        RECT 6.1480 25.6635 6.1740 26.7570 ;
        RECT 6.0400 25.6635 6.0660 26.7570 ;
        RECT 5.9320 25.6635 5.9580 26.7570 ;
        RECT 5.8240 25.6635 5.8500 26.7570 ;
        RECT 5.7160 25.6635 5.7420 26.7570 ;
        RECT 5.6080 25.6635 5.6340 26.7570 ;
        RECT 5.5000 25.6635 5.5260 26.7570 ;
        RECT 5.3920 25.6635 5.4180 26.7570 ;
        RECT 5.2840 25.6635 5.3100 26.7570 ;
        RECT 5.1760 25.6635 5.2020 26.7570 ;
        RECT 5.0680 25.6635 5.0940 26.7570 ;
        RECT 4.9600 25.6635 4.9860 26.7570 ;
        RECT 4.8520 25.6635 4.8780 26.7570 ;
        RECT 4.7440 25.6635 4.7700 26.7570 ;
        RECT 4.6360 25.6635 4.6620 26.7570 ;
        RECT 4.5280 25.6635 4.5540 26.7570 ;
        RECT 4.4200 25.6635 4.4460 26.7570 ;
        RECT 4.3120 25.6635 4.3380 26.7570 ;
        RECT 4.2040 25.6635 4.2300 26.7570 ;
        RECT 4.0960 25.6635 4.1220 26.7570 ;
        RECT 3.9880 25.6635 4.0140 26.7570 ;
        RECT 3.8800 25.6635 3.9060 26.7570 ;
        RECT 3.7720 25.6635 3.7980 26.7570 ;
        RECT 3.6640 25.6635 3.6900 26.7570 ;
        RECT 3.5560 25.6635 3.5820 26.7570 ;
        RECT 3.4480 25.6635 3.4740 26.7570 ;
        RECT 3.3400 25.6635 3.3660 26.7570 ;
        RECT 3.2320 25.6635 3.2580 26.7570 ;
        RECT 3.1240 25.6635 3.1500 26.7570 ;
        RECT 3.0160 25.6635 3.0420 26.7570 ;
        RECT 2.9080 25.6635 2.9340 26.7570 ;
        RECT 2.8000 25.6635 2.8260 26.7570 ;
        RECT 2.6920 25.6635 2.7180 26.7570 ;
        RECT 2.5840 25.6635 2.6100 26.7570 ;
        RECT 2.4760 25.6635 2.5020 26.7570 ;
        RECT 2.3680 25.6635 2.3940 26.7570 ;
        RECT 2.2600 25.6635 2.2860 26.7570 ;
        RECT 2.1520 25.6635 2.1780 26.7570 ;
        RECT 2.0440 25.6635 2.0700 26.7570 ;
        RECT 1.9360 25.6635 1.9620 26.7570 ;
        RECT 1.8280 25.6635 1.8540 26.7570 ;
        RECT 1.7200 25.6635 1.7460 26.7570 ;
        RECT 1.6120 25.6635 1.6380 26.7570 ;
        RECT 1.5040 25.6635 1.5300 26.7570 ;
        RECT 1.3960 25.6635 1.4220 26.7570 ;
        RECT 1.2880 25.6635 1.3140 26.7570 ;
        RECT 1.1800 25.6635 1.2060 26.7570 ;
        RECT 1.0720 25.6635 1.0980 26.7570 ;
        RECT 0.9640 25.6635 0.9900 26.7570 ;
        RECT 0.8560 25.6635 0.8820 26.7570 ;
        RECT 0.7480 25.6635 0.7740 26.7570 ;
        RECT 0.6400 25.6635 0.6660 26.7570 ;
        RECT 0.5320 25.6635 0.5580 26.7570 ;
        RECT 0.4240 25.6635 0.4500 26.7570 ;
        RECT 0.3160 25.6635 0.3420 26.7570 ;
        RECT 0.2080 25.6635 0.2340 26.7570 ;
        RECT 0.0050 25.6635 0.0900 26.7570 ;
        RECT 8.6410 26.7435 8.7690 27.8370 ;
        RECT 8.6270 27.4090 8.7690 27.7315 ;
        RECT 8.4790 27.1360 8.5410 27.8370 ;
        RECT 8.4650 27.4455 8.5410 27.5990 ;
        RECT 8.4790 26.7435 8.5050 27.8370 ;
        RECT 8.4790 26.8645 8.5190 27.1040 ;
        RECT 8.4790 26.7435 8.5410 26.8325 ;
        RECT 8.1820 27.1940 8.3880 27.8370 ;
        RECT 8.3620 26.7435 8.3880 27.8370 ;
        RECT 8.1820 27.4710 8.4020 27.7290 ;
        RECT 8.1820 26.7435 8.2800 27.8370 ;
        RECT 7.7650 26.7435 7.8480 27.8370 ;
        RECT 7.7650 26.8320 7.8620 27.7675 ;
        RECT 16.4440 26.7435 16.5290 27.8370 ;
        RECT 16.3000 26.7435 16.3260 27.8370 ;
        RECT 16.1920 26.7435 16.2180 27.8370 ;
        RECT 16.0840 26.7435 16.1100 27.8370 ;
        RECT 15.9760 26.7435 16.0020 27.8370 ;
        RECT 15.8680 26.7435 15.8940 27.8370 ;
        RECT 15.7600 26.7435 15.7860 27.8370 ;
        RECT 15.6520 26.7435 15.6780 27.8370 ;
        RECT 15.5440 26.7435 15.5700 27.8370 ;
        RECT 15.4360 26.7435 15.4620 27.8370 ;
        RECT 15.3280 26.7435 15.3540 27.8370 ;
        RECT 15.2200 26.7435 15.2460 27.8370 ;
        RECT 15.1120 26.7435 15.1380 27.8370 ;
        RECT 15.0040 26.7435 15.0300 27.8370 ;
        RECT 14.8960 26.7435 14.9220 27.8370 ;
        RECT 14.7880 26.7435 14.8140 27.8370 ;
        RECT 14.6800 26.7435 14.7060 27.8370 ;
        RECT 14.5720 26.7435 14.5980 27.8370 ;
        RECT 14.4640 26.7435 14.4900 27.8370 ;
        RECT 14.3560 26.7435 14.3820 27.8370 ;
        RECT 14.2480 26.7435 14.2740 27.8370 ;
        RECT 14.1400 26.7435 14.1660 27.8370 ;
        RECT 14.0320 26.7435 14.0580 27.8370 ;
        RECT 13.9240 26.7435 13.9500 27.8370 ;
        RECT 13.8160 26.7435 13.8420 27.8370 ;
        RECT 13.7080 26.7435 13.7340 27.8370 ;
        RECT 13.6000 26.7435 13.6260 27.8370 ;
        RECT 13.4920 26.7435 13.5180 27.8370 ;
        RECT 13.3840 26.7435 13.4100 27.8370 ;
        RECT 13.2760 26.7435 13.3020 27.8370 ;
        RECT 13.1680 26.7435 13.1940 27.8370 ;
        RECT 13.0600 26.7435 13.0860 27.8370 ;
        RECT 12.9520 26.7435 12.9780 27.8370 ;
        RECT 12.8440 26.7435 12.8700 27.8370 ;
        RECT 12.7360 26.7435 12.7620 27.8370 ;
        RECT 12.6280 26.7435 12.6540 27.8370 ;
        RECT 12.5200 26.7435 12.5460 27.8370 ;
        RECT 12.4120 26.7435 12.4380 27.8370 ;
        RECT 12.3040 26.7435 12.3300 27.8370 ;
        RECT 12.1960 26.7435 12.2220 27.8370 ;
        RECT 12.0880 26.7435 12.1140 27.8370 ;
        RECT 11.9800 26.7435 12.0060 27.8370 ;
        RECT 11.8720 26.7435 11.8980 27.8370 ;
        RECT 11.7640 26.7435 11.7900 27.8370 ;
        RECT 11.6560 26.7435 11.6820 27.8370 ;
        RECT 11.5480 26.7435 11.5740 27.8370 ;
        RECT 11.4400 26.7435 11.4660 27.8370 ;
        RECT 11.3320 26.7435 11.3580 27.8370 ;
        RECT 11.2240 26.7435 11.2500 27.8370 ;
        RECT 11.1160 26.7435 11.1420 27.8370 ;
        RECT 11.0080 26.7435 11.0340 27.8370 ;
        RECT 10.9000 26.7435 10.9260 27.8370 ;
        RECT 10.7920 26.7435 10.8180 27.8370 ;
        RECT 10.6840 26.7435 10.7100 27.8370 ;
        RECT 10.5760 26.7435 10.6020 27.8370 ;
        RECT 10.4680 26.7435 10.4940 27.8370 ;
        RECT 10.3600 26.7435 10.3860 27.8370 ;
        RECT 10.2520 26.7435 10.2780 27.8370 ;
        RECT 10.1440 26.7435 10.1700 27.8370 ;
        RECT 10.0360 26.7435 10.0620 27.8370 ;
        RECT 9.9280 26.7435 9.9540 27.8370 ;
        RECT 9.8200 26.7435 9.8460 27.8370 ;
        RECT 9.7120 26.7435 9.7380 27.8370 ;
        RECT 9.6040 26.7435 9.6300 27.8370 ;
        RECT 9.4960 26.7435 9.5220 27.8370 ;
        RECT 9.3880 26.7435 9.4140 27.8370 ;
        RECT 9.1750 26.7435 9.2520 27.8370 ;
        RECT 7.2820 26.7435 7.3590 27.8370 ;
        RECT 7.1200 26.7435 7.1460 27.8370 ;
        RECT 7.0120 26.7435 7.0380 27.8370 ;
        RECT 6.9040 26.7435 6.9300 27.8370 ;
        RECT 6.7960 26.7435 6.8220 27.8370 ;
        RECT 6.6880 26.7435 6.7140 27.8370 ;
        RECT 6.5800 26.7435 6.6060 27.8370 ;
        RECT 6.4720 26.7435 6.4980 27.8370 ;
        RECT 6.3640 26.7435 6.3900 27.8370 ;
        RECT 6.2560 26.7435 6.2820 27.8370 ;
        RECT 6.1480 26.7435 6.1740 27.8370 ;
        RECT 6.0400 26.7435 6.0660 27.8370 ;
        RECT 5.9320 26.7435 5.9580 27.8370 ;
        RECT 5.8240 26.7435 5.8500 27.8370 ;
        RECT 5.7160 26.7435 5.7420 27.8370 ;
        RECT 5.6080 26.7435 5.6340 27.8370 ;
        RECT 5.5000 26.7435 5.5260 27.8370 ;
        RECT 5.3920 26.7435 5.4180 27.8370 ;
        RECT 5.2840 26.7435 5.3100 27.8370 ;
        RECT 5.1760 26.7435 5.2020 27.8370 ;
        RECT 5.0680 26.7435 5.0940 27.8370 ;
        RECT 4.9600 26.7435 4.9860 27.8370 ;
        RECT 4.8520 26.7435 4.8780 27.8370 ;
        RECT 4.7440 26.7435 4.7700 27.8370 ;
        RECT 4.6360 26.7435 4.6620 27.8370 ;
        RECT 4.5280 26.7435 4.5540 27.8370 ;
        RECT 4.4200 26.7435 4.4460 27.8370 ;
        RECT 4.3120 26.7435 4.3380 27.8370 ;
        RECT 4.2040 26.7435 4.2300 27.8370 ;
        RECT 4.0960 26.7435 4.1220 27.8370 ;
        RECT 3.9880 26.7435 4.0140 27.8370 ;
        RECT 3.8800 26.7435 3.9060 27.8370 ;
        RECT 3.7720 26.7435 3.7980 27.8370 ;
        RECT 3.6640 26.7435 3.6900 27.8370 ;
        RECT 3.5560 26.7435 3.5820 27.8370 ;
        RECT 3.4480 26.7435 3.4740 27.8370 ;
        RECT 3.3400 26.7435 3.3660 27.8370 ;
        RECT 3.2320 26.7435 3.2580 27.8370 ;
        RECT 3.1240 26.7435 3.1500 27.8370 ;
        RECT 3.0160 26.7435 3.0420 27.8370 ;
        RECT 2.9080 26.7435 2.9340 27.8370 ;
        RECT 2.8000 26.7435 2.8260 27.8370 ;
        RECT 2.6920 26.7435 2.7180 27.8370 ;
        RECT 2.5840 26.7435 2.6100 27.8370 ;
        RECT 2.4760 26.7435 2.5020 27.8370 ;
        RECT 2.3680 26.7435 2.3940 27.8370 ;
        RECT 2.2600 26.7435 2.2860 27.8370 ;
        RECT 2.1520 26.7435 2.1780 27.8370 ;
        RECT 2.0440 26.7435 2.0700 27.8370 ;
        RECT 1.9360 26.7435 1.9620 27.8370 ;
        RECT 1.8280 26.7435 1.8540 27.8370 ;
        RECT 1.7200 26.7435 1.7460 27.8370 ;
        RECT 1.6120 26.7435 1.6380 27.8370 ;
        RECT 1.5040 26.7435 1.5300 27.8370 ;
        RECT 1.3960 26.7435 1.4220 27.8370 ;
        RECT 1.2880 26.7435 1.3140 27.8370 ;
        RECT 1.1800 26.7435 1.2060 27.8370 ;
        RECT 1.0720 26.7435 1.0980 27.8370 ;
        RECT 0.9640 26.7435 0.9900 27.8370 ;
        RECT 0.8560 26.7435 0.8820 27.8370 ;
        RECT 0.7480 26.7435 0.7740 27.8370 ;
        RECT 0.6400 26.7435 0.6660 27.8370 ;
        RECT 0.5320 26.7435 0.5580 27.8370 ;
        RECT 0.4240 26.7435 0.4500 27.8370 ;
        RECT 0.3160 26.7435 0.3420 27.8370 ;
        RECT 0.2080 26.7435 0.2340 27.8370 ;
        RECT 0.0050 26.7435 0.0900 27.8370 ;
  LAYER V3 SPACING 0.018  ;
      RECT 0.0050 1.2200 16.5290 1.3500 ;
      RECT 16.4120 0.2565 16.5290 1.3500 ;
      RECT 9.3020 1.1240 16.3940 1.3500 ;
      RECT 7.9700 1.1240 9.2840 1.3500 ;
      RECT 7.2500 0.2565 7.8800 1.3500 ;
      RECT 0.1400 1.1240 7.2320 1.3500 ;
      RECT 0.0050 0.2565 0.1220 1.3500 ;
      RECT 16.3760 0.2565 16.5290 1.1720 ;
      RECT 9.3560 0.2565 16.3580 1.3500 ;
      RECT 8.6090 0.2565 9.3380 1.1720 ;
      RECT 8.4470 0.4520 8.5730 1.3500 ;
      RECT 7.1960 0.3560 8.4200 1.1720 ;
      RECT 0.1760 0.2565 7.1780 1.3500 ;
      RECT 0.0050 0.2565 0.1580 1.1720 ;
      RECT 8.5550 0.2565 16.5290 1.0760 ;
      RECT 0.0050 0.3560 8.5370 1.0760 ;
      RECT 8.3300 0.2565 16.5290 0.4280 ;
      RECT 0.0050 0.2565 8.3120 1.0760 ;
      RECT 0.0050 0.2565 16.5290 0.3320 ;
      RECT 0.0050 2.3000 16.5290 2.4300 ;
      RECT 16.4120 1.3365 16.5290 2.4300 ;
      RECT 9.3020 2.2040 16.3940 2.4300 ;
      RECT 7.9700 2.2040 9.2840 2.4300 ;
      RECT 7.2500 1.3365 7.8800 2.4300 ;
      RECT 0.1400 2.2040 7.2320 2.4300 ;
      RECT 0.0050 1.3365 0.1220 2.4300 ;
      RECT 16.3760 1.3365 16.5290 2.2520 ;
      RECT 9.3560 1.3365 16.3580 2.4300 ;
      RECT 8.6090 1.3365 9.3380 2.2520 ;
      RECT 8.4470 1.5320 8.5730 2.4300 ;
      RECT 7.1960 1.4360 8.4200 2.2520 ;
      RECT 0.1760 1.3365 7.1780 2.4300 ;
      RECT 0.0050 1.3365 0.1580 2.2520 ;
      RECT 8.5550 1.3365 16.5290 2.1560 ;
      RECT 0.0050 1.4360 8.5370 2.1560 ;
      RECT 8.3300 1.3365 16.5290 1.5080 ;
      RECT 0.0050 1.3365 8.3120 2.1560 ;
      RECT 0.0050 1.3365 16.5290 1.4120 ;
      RECT 0.0050 3.3800 16.5290 3.5100 ;
      RECT 16.4120 2.4165 16.5290 3.5100 ;
      RECT 9.3020 3.2840 16.3940 3.5100 ;
      RECT 7.9700 3.2840 9.2840 3.5100 ;
      RECT 7.2500 2.4165 7.8800 3.5100 ;
      RECT 0.1400 3.2840 7.2320 3.5100 ;
      RECT 0.0050 2.4165 0.1220 3.5100 ;
      RECT 16.3760 2.4165 16.5290 3.3320 ;
      RECT 9.3560 2.4165 16.3580 3.5100 ;
      RECT 8.6090 2.4165 9.3380 3.3320 ;
      RECT 8.4470 2.6120 8.5730 3.5100 ;
      RECT 7.1960 2.5160 8.4200 3.3320 ;
      RECT 0.1760 2.4165 7.1780 3.5100 ;
      RECT 0.0050 2.4165 0.1580 3.3320 ;
      RECT 8.5550 2.4165 16.5290 3.2360 ;
      RECT 0.0050 2.5160 8.5370 3.2360 ;
      RECT 8.3300 2.4165 16.5290 2.5880 ;
      RECT 0.0050 2.4165 8.3120 3.2360 ;
      RECT 0.0050 2.4165 16.5290 2.4920 ;
      RECT 0.0050 4.4600 16.5290 4.5900 ;
      RECT 16.4120 3.4965 16.5290 4.5900 ;
      RECT 9.3020 4.3640 16.3940 4.5900 ;
      RECT 7.9700 4.3640 9.2840 4.5900 ;
      RECT 7.2500 3.4965 7.8800 4.5900 ;
      RECT 0.1400 4.3640 7.2320 4.5900 ;
      RECT 0.0050 3.4965 0.1220 4.5900 ;
      RECT 16.3760 3.4965 16.5290 4.4120 ;
      RECT 9.3560 3.4965 16.3580 4.5900 ;
      RECT 8.6090 3.4965 9.3380 4.4120 ;
      RECT 8.4470 3.6920 8.5730 4.5900 ;
      RECT 7.1960 3.5960 8.4200 4.4120 ;
      RECT 0.1760 3.4965 7.1780 4.5900 ;
      RECT 0.0050 3.4965 0.1580 4.4120 ;
      RECT 8.5550 3.4965 16.5290 4.3160 ;
      RECT 0.0050 3.5960 8.5370 4.3160 ;
      RECT 8.3300 3.4965 16.5290 3.6680 ;
      RECT 0.0050 3.4965 8.3120 4.3160 ;
      RECT 0.0050 3.4965 16.5290 3.5720 ;
      RECT 0.0050 5.5400 16.5290 5.6700 ;
      RECT 16.4120 4.5765 16.5290 5.6700 ;
      RECT 9.3020 5.4440 16.3940 5.6700 ;
      RECT 7.9700 5.4440 9.2840 5.6700 ;
      RECT 7.2500 4.5765 7.8800 5.6700 ;
      RECT 0.1400 5.4440 7.2320 5.6700 ;
      RECT 0.0050 4.5765 0.1220 5.6700 ;
      RECT 16.3760 4.5765 16.5290 5.4920 ;
      RECT 9.3560 4.5765 16.3580 5.6700 ;
      RECT 8.6090 4.5765 9.3380 5.4920 ;
      RECT 8.4470 4.7720 8.5730 5.6700 ;
      RECT 7.1960 4.6760 8.4200 5.4920 ;
      RECT 0.1760 4.5765 7.1780 5.6700 ;
      RECT 0.0050 4.5765 0.1580 5.4920 ;
      RECT 8.5550 4.5765 16.5290 5.3960 ;
      RECT 0.0050 4.6760 8.5370 5.3960 ;
      RECT 8.3300 4.5765 16.5290 4.7480 ;
      RECT 0.0050 4.5765 8.3120 5.3960 ;
      RECT 0.0050 4.5765 16.5290 4.6520 ;
      RECT 0.0050 6.6200 16.5290 6.7500 ;
      RECT 16.4120 5.6565 16.5290 6.7500 ;
      RECT 9.3020 6.5240 16.3940 6.7500 ;
      RECT 7.9700 6.5240 9.2840 6.7500 ;
      RECT 7.2500 5.6565 7.8800 6.7500 ;
      RECT 0.1400 6.5240 7.2320 6.7500 ;
      RECT 0.0050 5.6565 0.1220 6.7500 ;
      RECT 16.3760 5.6565 16.5290 6.5720 ;
      RECT 9.3560 5.6565 16.3580 6.7500 ;
      RECT 8.6090 5.6565 9.3380 6.5720 ;
      RECT 8.4470 5.8520 8.5730 6.7500 ;
      RECT 7.1960 5.7560 8.4200 6.5720 ;
      RECT 0.1760 5.6565 7.1780 6.7500 ;
      RECT 0.0050 5.6565 0.1580 6.5720 ;
      RECT 8.5550 5.6565 16.5290 6.4760 ;
      RECT 0.0050 5.7560 8.5370 6.4760 ;
      RECT 8.3300 5.6565 16.5290 5.8280 ;
      RECT 0.0050 5.6565 8.3120 6.4760 ;
      RECT 0.0050 5.6565 16.5290 5.7320 ;
      RECT 0.0050 7.7000 16.5290 7.8300 ;
      RECT 16.4120 6.7365 16.5290 7.8300 ;
      RECT 9.3020 7.6040 16.3940 7.8300 ;
      RECT 7.9700 7.6040 9.2840 7.8300 ;
      RECT 7.2500 6.7365 7.8800 7.8300 ;
      RECT 0.1400 7.6040 7.2320 7.8300 ;
      RECT 0.0050 6.7365 0.1220 7.8300 ;
      RECT 16.3760 6.7365 16.5290 7.6520 ;
      RECT 9.3560 6.7365 16.3580 7.8300 ;
      RECT 8.6090 6.7365 9.3380 7.6520 ;
      RECT 8.4470 6.9320 8.5730 7.8300 ;
      RECT 7.1960 6.8360 8.4200 7.6520 ;
      RECT 0.1760 6.7365 7.1780 7.8300 ;
      RECT 0.0050 6.7365 0.1580 7.6520 ;
      RECT 8.5550 6.7365 16.5290 7.5560 ;
      RECT 0.0050 6.8360 8.5370 7.5560 ;
      RECT 8.3300 6.7365 16.5290 6.9080 ;
      RECT 0.0050 6.7365 8.3120 7.5560 ;
      RECT 0.0050 6.7365 16.5290 6.8120 ;
      RECT 0.0050 8.7800 16.5290 8.9100 ;
      RECT 16.4120 7.8165 16.5290 8.9100 ;
      RECT 9.3020 8.6840 16.3940 8.9100 ;
      RECT 7.9700 8.6840 9.2840 8.9100 ;
      RECT 7.2500 7.8165 7.8800 8.9100 ;
      RECT 0.1400 8.6840 7.2320 8.9100 ;
      RECT 0.0050 7.8165 0.1220 8.9100 ;
      RECT 16.3760 7.8165 16.5290 8.7320 ;
      RECT 9.3560 7.8165 16.3580 8.9100 ;
      RECT 8.6090 7.8165 9.3380 8.7320 ;
      RECT 8.4470 8.0120 8.5730 8.9100 ;
      RECT 7.1960 7.9160 8.4200 8.7320 ;
      RECT 0.1760 7.8165 7.1780 8.9100 ;
      RECT 0.0050 7.8165 0.1580 8.7320 ;
      RECT 8.5550 7.8165 16.5290 8.6360 ;
      RECT 0.0050 7.9160 8.5370 8.6360 ;
      RECT 8.3300 7.8165 16.5290 7.9880 ;
      RECT 0.0050 7.8165 8.3120 8.6360 ;
      RECT 0.0050 7.8165 16.5290 7.8920 ;
      RECT 0.0050 9.8600 16.5290 9.9900 ;
      RECT 16.4120 8.8965 16.5290 9.9900 ;
      RECT 9.3020 9.7640 16.3940 9.9900 ;
      RECT 7.9700 9.7640 9.2840 9.9900 ;
      RECT 7.2500 8.8965 7.8800 9.9900 ;
      RECT 0.1400 9.7640 7.2320 9.9900 ;
      RECT 0.0050 8.8965 0.1220 9.9900 ;
      RECT 16.3760 8.8965 16.5290 9.8120 ;
      RECT 9.3560 8.8965 16.3580 9.9900 ;
      RECT 8.6090 8.8965 9.3380 9.8120 ;
      RECT 8.4470 9.0920 8.5730 9.9900 ;
      RECT 7.1960 8.9960 8.4200 9.8120 ;
      RECT 0.1760 8.8965 7.1780 9.9900 ;
      RECT 0.0050 8.8965 0.1580 9.8120 ;
      RECT 8.5550 8.8965 16.5290 9.7160 ;
      RECT 0.0050 8.9960 8.5370 9.7160 ;
      RECT 8.3300 8.8965 16.5290 9.0680 ;
      RECT 0.0050 8.8965 8.3120 9.7160 ;
      RECT 0.0050 8.8965 16.5290 8.9720 ;
      RECT 0.0000 17.2770 16.5240 18.6105 ;
      RECT 10.8090 9.9570 16.5240 18.6105 ;
      RECT 8.6090 13.8210 16.5240 18.6105 ;
      RECT 9.5130 11.2290 16.5240 18.6105 ;
      RECT 8.5570 9.9570 8.5910 18.6105 ;
      RECT 8.5050 9.9570 8.5390 18.6105 ;
      RECT 8.4530 9.9570 8.4870 18.6105 ;
      RECT 8.4010 9.9570 8.4350 18.6105 ;
      RECT 0.0000 16.8450 8.3830 18.6105 ;
      RECT 8.1410 14.1090 16.5240 17.0610 ;
      RECT 8.0890 9.9570 8.1230 18.6105 ;
      RECT 8.0370 9.9570 8.0710 18.6105 ;
      RECT 7.9850 9.9570 8.0190 18.6105 ;
      RECT 7.9330 9.9570 7.9670 18.6105 ;
      RECT 0.0000 11.5170 7.9150 18.6105 ;
      RECT 0.0000 13.6770 8.3830 16.6290 ;
      RECT 8.1410 10.9410 9.2790 13.8930 ;
      RECT 9.3150 11.4210 16.5240 18.6105 ;
      RECT 0.0000 13.6770 9.2970 13.8930 ;
      RECT 8.1410 11.4210 16.5240 13.7970 ;
      RECT 7.4610 10.5090 8.2350 13.4610 ;
      RECT 7.2450 10.6530 7.9150 18.6105 ;
      RECT 0.0000 11.2290 7.2270 18.6105 ;
      RECT 6.8130 9.9570 7.2630 11.4930 ;
      RECT 0.0000 11.3250 9.4950 11.4930 ;
      RECT 9.2970 11.2290 16.5240 11.3970 ;
      RECT 10.5930 9.9570 10.7910 18.6105 ;
      RECT 6.8130 11.0370 10.5750 11.3010 ;
      RECT 5.9490 10.6530 6.7950 18.6105 ;
      RECT 0.0000 9.9570 5.9310 18.6105 ;
      RECT 10.3770 9.9570 16.5240 11.2050 ;
      RECT 10.1610 10.6530 16.5240 11.2050 ;
      RECT 0.0000 10.9415 10.1430 11.2050 ;
      RECT 9.9450 9.9570 10.3590 11.0130 ;
      RECT 9.3510 10.6530 16.5240 11.0130 ;
      RECT 8.6090 10.6530 9.3330 11.3010 ;
      RECT 8.1410 10.6050 8.3830 18.6105 ;
      RECT 8.2530 9.9570 8.6310 10.7250 ;
      RECT 8.6490 10.6050 9.9270 10.7255 ;
      RECT 6.5970 10.6050 7.4430 11.2050 ;
      RECT 6.1650 10.6050 6.5790 18.6105 ;
      RECT 0.0000 9.9570 6.1470 11.2050 ;
      RECT 9.7290 9.9570 16.5240 10.6290 ;
      RECT 8.2530 10.0370 9.7110 10.6290 ;
      RECT 7.2810 10.5090 8.2350 10.6290 ;
      RECT 6.3810 9.9570 7.2630 10.6290 ;
      RECT 0.0000 9.9570 6.3630 10.6290 ;
      RECT 9.2970 9.9570 16.5240 10.5810 ;
      RECT 8.1410 10.0370 16.5240 10.5810 ;
      RECT 0.0000 9.9570 7.9150 10.5810 ;
      RECT 0.0000 9.9570 9.2790 10.2930 ;
      RECT 0.0000 9.9570 16.5240 10.0130 ;
        RECT 0.0050 19.0670 16.5290 19.1970 ;
        RECT 16.4120 18.1035 16.5290 19.1970 ;
        RECT 9.3020 18.9710 16.3940 19.1970 ;
        RECT 7.9700 18.9710 9.2840 19.1970 ;
        RECT 7.2500 18.1035 7.8800 19.1970 ;
        RECT 0.1400 18.9710 7.2320 19.1970 ;
        RECT 0.0050 18.1035 0.1220 19.1970 ;
        RECT 16.3760 18.1035 16.5290 19.0190 ;
        RECT 9.3560 18.1035 16.3580 19.1970 ;
        RECT 8.6090 18.1035 9.3380 19.0190 ;
        RECT 8.4470 18.2990 8.5730 19.1970 ;
        RECT 7.1960 18.2030 8.4200 19.0190 ;
        RECT 0.1760 18.1035 7.1780 19.1970 ;
        RECT 0.0050 18.1035 0.1580 19.0190 ;
        RECT 8.5550 18.1035 16.5290 18.9230 ;
        RECT 0.0050 18.2030 8.5370 18.9230 ;
        RECT 8.3300 18.1035 16.5290 18.2750 ;
        RECT 0.0050 18.1035 8.3120 18.9230 ;
        RECT 0.0050 18.1035 16.5290 18.1790 ;
        RECT 0.0050 20.1470 16.5290 20.2770 ;
        RECT 16.4120 19.1835 16.5290 20.2770 ;
        RECT 9.3020 20.0510 16.3940 20.2770 ;
        RECT 7.9700 20.0510 9.2840 20.2770 ;
        RECT 7.2500 19.1835 7.8800 20.2770 ;
        RECT 0.1400 20.0510 7.2320 20.2770 ;
        RECT 0.0050 19.1835 0.1220 20.2770 ;
        RECT 16.3760 19.1835 16.5290 20.0990 ;
        RECT 9.3560 19.1835 16.3580 20.2770 ;
        RECT 8.6090 19.1835 9.3380 20.0990 ;
        RECT 8.4470 19.3790 8.5730 20.2770 ;
        RECT 7.1960 19.2830 8.4200 20.0990 ;
        RECT 0.1760 19.1835 7.1780 20.2770 ;
        RECT 0.0050 19.1835 0.1580 20.0990 ;
        RECT 8.5550 19.1835 16.5290 20.0030 ;
        RECT 0.0050 19.2830 8.5370 20.0030 ;
        RECT 8.3300 19.1835 16.5290 19.3550 ;
        RECT 0.0050 19.1835 8.3120 20.0030 ;
        RECT 0.0050 19.1835 16.5290 19.2590 ;
        RECT 0.0050 21.2270 16.5290 21.3570 ;
        RECT 16.4120 20.2635 16.5290 21.3570 ;
        RECT 9.3020 21.1310 16.3940 21.3570 ;
        RECT 7.9700 21.1310 9.2840 21.3570 ;
        RECT 7.2500 20.2635 7.8800 21.3570 ;
        RECT 0.1400 21.1310 7.2320 21.3570 ;
        RECT 0.0050 20.2635 0.1220 21.3570 ;
        RECT 16.3760 20.2635 16.5290 21.1790 ;
        RECT 9.3560 20.2635 16.3580 21.3570 ;
        RECT 8.6090 20.2635 9.3380 21.1790 ;
        RECT 8.4470 20.4590 8.5730 21.3570 ;
        RECT 7.1960 20.3630 8.4200 21.1790 ;
        RECT 0.1760 20.2635 7.1780 21.3570 ;
        RECT 0.0050 20.2635 0.1580 21.1790 ;
        RECT 8.5550 20.2635 16.5290 21.0830 ;
        RECT 0.0050 20.3630 8.5370 21.0830 ;
        RECT 8.3300 20.2635 16.5290 20.4350 ;
        RECT 0.0050 20.2635 8.3120 21.0830 ;
        RECT 0.0050 20.2635 16.5290 20.3390 ;
        RECT 0.0050 22.3070 16.5290 22.4370 ;
        RECT 16.4120 21.3435 16.5290 22.4370 ;
        RECT 9.3020 22.2110 16.3940 22.4370 ;
        RECT 7.9700 22.2110 9.2840 22.4370 ;
        RECT 7.2500 21.3435 7.8800 22.4370 ;
        RECT 0.1400 22.2110 7.2320 22.4370 ;
        RECT 0.0050 21.3435 0.1220 22.4370 ;
        RECT 16.3760 21.3435 16.5290 22.2590 ;
        RECT 9.3560 21.3435 16.3580 22.4370 ;
        RECT 8.6090 21.3435 9.3380 22.2590 ;
        RECT 8.4470 21.5390 8.5730 22.4370 ;
        RECT 7.1960 21.4430 8.4200 22.2590 ;
        RECT 0.1760 21.3435 7.1780 22.4370 ;
        RECT 0.0050 21.3435 0.1580 22.2590 ;
        RECT 8.5550 21.3435 16.5290 22.1630 ;
        RECT 0.0050 21.4430 8.5370 22.1630 ;
        RECT 8.3300 21.3435 16.5290 21.5150 ;
        RECT 0.0050 21.3435 8.3120 22.1630 ;
        RECT 0.0050 21.3435 16.5290 21.4190 ;
        RECT 0.0050 23.3870 16.5290 23.5170 ;
        RECT 16.4120 22.4235 16.5290 23.5170 ;
        RECT 9.3020 23.2910 16.3940 23.5170 ;
        RECT 7.9700 23.2910 9.2840 23.5170 ;
        RECT 7.2500 22.4235 7.8800 23.5170 ;
        RECT 0.1400 23.2910 7.2320 23.5170 ;
        RECT 0.0050 22.4235 0.1220 23.5170 ;
        RECT 16.3760 22.4235 16.5290 23.3390 ;
        RECT 9.3560 22.4235 16.3580 23.5170 ;
        RECT 8.6090 22.4235 9.3380 23.3390 ;
        RECT 8.4470 22.6190 8.5730 23.5170 ;
        RECT 7.1960 22.5230 8.4200 23.3390 ;
        RECT 0.1760 22.4235 7.1780 23.5170 ;
        RECT 0.0050 22.4235 0.1580 23.3390 ;
        RECT 8.5550 22.4235 16.5290 23.2430 ;
        RECT 0.0050 22.5230 8.5370 23.2430 ;
        RECT 8.3300 22.4235 16.5290 22.5950 ;
        RECT 0.0050 22.4235 8.3120 23.2430 ;
        RECT 0.0050 22.4235 16.5290 22.4990 ;
        RECT 0.0050 24.4670 16.5290 24.5970 ;
        RECT 16.4120 23.5035 16.5290 24.5970 ;
        RECT 9.3020 24.3710 16.3940 24.5970 ;
        RECT 7.9700 24.3710 9.2840 24.5970 ;
        RECT 7.2500 23.5035 7.8800 24.5970 ;
        RECT 0.1400 24.3710 7.2320 24.5970 ;
        RECT 0.0050 23.5035 0.1220 24.5970 ;
        RECT 16.3760 23.5035 16.5290 24.4190 ;
        RECT 9.3560 23.5035 16.3580 24.5970 ;
        RECT 8.6090 23.5035 9.3380 24.4190 ;
        RECT 8.4470 23.6990 8.5730 24.5970 ;
        RECT 7.1960 23.6030 8.4200 24.4190 ;
        RECT 0.1760 23.5035 7.1780 24.5970 ;
        RECT 0.0050 23.5035 0.1580 24.4190 ;
        RECT 8.5550 23.5035 16.5290 24.3230 ;
        RECT 0.0050 23.6030 8.5370 24.3230 ;
        RECT 8.3300 23.5035 16.5290 23.6750 ;
        RECT 0.0050 23.5035 8.3120 24.3230 ;
        RECT 0.0050 23.5035 16.5290 23.5790 ;
        RECT 0.0050 25.5470 16.5290 25.6770 ;
        RECT 16.4120 24.5835 16.5290 25.6770 ;
        RECT 9.3020 25.4510 16.3940 25.6770 ;
        RECT 7.9700 25.4510 9.2840 25.6770 ;
        RECT 7.2500 24.5835 7.8800 25.6770 ;
        RECT 0.1400 25.4510 7.2320 25.6770 ;
        RECT 0.0050 24.5835 0.1220 25.6770 ;
        RECT 16.3760 24.5835 16.5290 25.4990 ;
        RECT 9.3560 24.5835 16.3580 25.6770 ;
        RECT 8.6090 24.5835 9.3380 25.4990 ;
        RECT 8.4470 24.7790 8.5730 25.6770 ;
        RECT 7.1960 24.6830 8.4200 25.4990 ;
        RECT 0.1760 24.5835 7.1780 25.6770 ;
        RECT 0.0050 24.5835 0.1580 25.4990 ;
        RECT 8.5550 24.5835 16.5290 25.4030 ;
        RECT 0.0050 24.6830 8.5370 25.4030 ;
        RECT 8.3300 24.5835 16.5290 24.7550 ;
        RECT 0.0050 24.5835 8.3120 25.4030 ;
        RECT 0.0050 24.5835 16.5290 24.6590 ;
        RECT 0.0050 26.6270 16.5290 26.7570 ;
        RECT 16.4120 25.6635 16.5290 26.7570 ;
        RECT 9.3020 26.5310 16.3940 26.7570 ;
        RECT 7.9700 26.5310 9.2840 26.7570 ;
        RECT 7.2500 25.6635 7.8800 26.7570 ;
        RECT 0.1400 26.5310 7.2320 26.7570 ;
        RECT 0.0050 25.6635 0.1220 26.7570 ;
        RECT 16.3760 25.6635 16.5290 26.5790 ;
        RECT 9.3560 25.6635 16.3580 26.7570 ;
        RECT 8.6090 25.6635 9.3380 26.5790 ;
        RECT 8.4470 25.8590 8.5730 26.7570 ;
        RECT 7.1960 25.7630 8.4200 26.5790 ;
        RECT 0.1760 25.6635 7.1780 26.7570 ;
        RECT 0.0050 25.6635 0.1580 26.5790 ;
        RECT 8.5550 25.6635 16.5290 26.4830 ;
        RECT 0.0050 25.7630 8.5370 26.4830 ;
        RECT 8.3300 25.6635 16.5290 25.8350 ;
        RECT 0.0050 25.6635 8.3120 26.4830 ;
        RECT 0.0050 25.6635 16.5290 25.7390 ;
        RECT 0.0050 27.7070 16.5290 27.8370 ;
        RECT 16.4120 26.7435 16.5290 27.8370 ;
        RECT 9.3020 27.6110 16.3940 27.8370 ;
        RECT 7.9700 27.6110 9.2840 27.8370 ;
        RECT 7.2500 26.7435 7.8800 27.8370 ;
        RECT 0.1400 27.6110 7.2320 27.8370 ;
        RECT 0.0050 26.7435 0.1220 27.8370 ;
        RECT 16.3760 26.7435 16.5290 27.6590 ;
        RECT 9.3560 26.7435 16.3580 27.8370 ;
        RECT 8.6090 26.7435 9.3380 27.6590 ;
        RECT 8.4470 26.9390 8.5730 27.8370 ;
        RECT 7.1960 26.8430 8.4200 27.6590 ;
        RECT 0.1760 26.7435 7.1780 27.8370 ;
        RECT 0.0050 26.7435 0.1580 27.6590 ;
        RECT 8.5550 26.7435 16.5290 27.5630 ;
        RECT 0.0050 26.8430 8.5370 27.5630 ;
        RECT 8.3300 26.7435 16.5290 26.9150 ;
        RECT 0.0050 26.7435 8.3120 27.5630 ;
        RECT 0.0050 26.7435 16.5290 26.8190 ;
  LAYER M4  ;
      RECT 1.5690 11.6700 15.0095 11.6940 ;
      RECT 1.5690 11.9580 15.0095 11.9820 ;
      RECT 1.5690 12.3420 15.0095 12.3660 ;
      RECT 1.5690 12.4380 15.0095 12.4620 ;
      RECT 1.5690 12.7740 15.0095 12.7980 ;
      RECT 1.5690 13.1580 15.0095 13.1820 ;
      RECT 10.9550 10.6290 11.0390 10.6530 ;
      RECT 10.7670 11.0610 10.8970 11.0850 ;
      RECT 10.7750 11.7185 10.8920 11.7425 ;
      RECT 10.7750 12.0060 10.8920 12.0300 ;
      RECT 10.1360 11.0610 10.7070 11.0850 ;
      RECT 10.1960 11.8380 10.3040 11.8620 ;
      RECT 8.8630 12.2130 9.9560 12.2370 ;
      RECT 9.5510 11.7810 9.6350 11.8050 ;
      RECT 8.7670 12.9810 9.6350 13.0050 ;
      RECT 9.5510 13.0770 9.6350 13.1010 ;
      RECT 9.3730 11.3010 9.4570 11.3250 ;
      RECT 9.3350 12.6450 9.4190 12.6690 ;
      RECT 9.3350 13.3650 9.4190 13.3890 ;
      RECT 9.1570 11.2050 9.2410 11.2290 ;
      RECT 8.9430 9.9170 9.2060 9.9410 ;
      RECT 8.9430 18.5410 9.2060 18.5650 ;
      RECT 8.9590 12.6930 9.2030 12.7170 ;
      RECT 9.1190 12.8370 9.2030 12.8610 ;
      RECT 7.6630 13.0770 9.2030 13.1010 ;
      RECT 9.1190 13.3650 9.2030 13.3890 ;
      RECT 8.8850 18.4450 9.1480 18.4690 ;
      RECT 8.8840 9.8210 9.1470 9.8450 ;
      RECT 8.8460 9.7250 9.1090 9.7490 ;
      RECT 8.8460 18.2530 9.1090 18.2770 ;
      RECT 9.0110 13.7970 9.0950 13.8210 ;
      RECT 8.2390 14.1810 9.0950 14.2050 ;
      RECT 8.6230 16.4370 9.0950 16.4610 ;
      RECT 9.0110 16.5330 9.0950 16.5570 ;
      RECT 8.7980 9.6290 9.0610 9.6530 ;
      RECT 8.7980 18.1570 9.0610 18.1810 ;
      RECT 8.5750 15.5250 9.0200 15.5490 ;
      RECT 8.7540 9.5330 9.0170 9.5570 ;
      RECT 8.7540 18.4930 9.0170 18.5170 ;
      RECT 8.7050 9.8690 8.9680 9.8930 ;
      RECT 8.7050 18.3970 8.9680 18.4210 ;
      RECT 8.8360 12.8370 8.9570 12.8610 ;
      RECT 8.8150 14.9490 8.9480 14.9730 ;
      RECT 8.6580 9.7730 8.9210 9.7970 ;
      RECT 8.6580 18.3010 8.9210 18.3250 ;
      RECT 8.6230 9.4850 8.8860 9.5090 ;
      RECT 8.6230 18.2050 8.8860 18.2290 ;
      RECT 7.8070 16.5330 8.8760 16.5570 ;
      RECT 8.7920 17.6850 8.8760 17.7090 ;
      RECT 8.5670 9.3410 8.8300 9.3650 ;
      RECT 8.5670 18.1090 8.8300 18.1330 ;
      RECT 8.7190 13.7970 8.8040 13.8210 ;
      RECT 7.6150 14.3730 8.7320 14.3970 ;
      RECT 8.2600 12.2130 8.7170 12.2370 ;
      RECT 8.0870 10.0610 8.3540 10.0850 ;
      RECT 8.0870 17.9650 8.3540 17.9890 ;
      RECT 8.2240 13.7490 8.3330 13.7730 ;
      RECT 8.0640 9.9650 8.3060 9.9890 ;
      RECT 8.0640 18.5890 8.3060 18.6130 ;
      RECT 8.0080 9.4850 8.2500 9.5090 ;
      RECT 8.0370 18.6850 8.2500 18.7090 ;
      RECT 8.1530 13.3650 8.2370 13.3890 ;
      RECT 7.9540 9.5810 8.2020 9.6050 ;
      RECT 7.9540 18.5410 8.2020 18.5650 ;
      RECT 7.7200 15.9570 8.1410 15.9810 ;
      RECT 7.6880 9.9170 7.9550 9.9410 ;
      RECT 7.6880 18.6850 7.9550 18.7090 ;
      RECT 7.8280 14.5170 7.9490 14.5410 ;
      RECT 7.8200 17.6850 7.9040 17.7090 ;
      RECT 7.6540 9.8210 7.9010 9.8450 ;
      RECT 7.5870 18.2530 7.9010 18.2770 ;
      RECT 7.6280 9.7250 7.8580 9.7490 ;
      RECT 7.6160 18.5890 7.8580 18.6130 ;
      RECT 7.5750 9.6290 7.8050 9.6530 ;
      RECT 7.7210 16.1010 7.8050 16.1250 ;
      RECT 7.5250 18.1570 7.8050 18.1810 ;
      RECT 7.5300 9.5330 7.7600 9.5570 ;
      RECT 7.5300 18.4930 7.7600 18.5170 ;
      RECT 6.5680 13.3650 7.7570 13.3890 ;
      RECT 7.4920 9.7730 7.7220 9.7970 ;
      RECT 7.4920 18.3970 7.7220 18.4210 ;
      RECT 7.4740 9.6770 7.6670 9.7010 ;
      RECT 7.4740 18.3010 7.6670 18.3250 ;
      RECT 7.4250 9.5810 7.6180 9.6050 ;
      RECT 7.4250 18.2050 7.6180 18.2290 ;
      RECT 7.4290 14.2770 7.6130 14.3010 ;
      RECT 7.3730 9.4850 7.5660 9.5090 ;
      RECT 7.3730 18.1090 7.5660 18.1330 ;
      RECT 6.8890 11.5890 7.5650 11.6130 ;
      RECT 7.4290 14.3730 7.5130 14.3970 ;
      RECT 7.1600 10.0130 7.4230 10.0370 ;
      RECT 7.1925 13.7970 7.3260 13.8210 ;
      RECT 6.8510 11.7810 6.9350 11.8050 ;
  LAYER V4  ;
      RECT 11.0040 10.6290 11.0280 10.6530 ;
      RECT 11.0040 11.6700 11.0280 11.6940 ;
      RECT 10.8360 11.0610 10.8600 11.0850 ;
      RECT 10.8360 11.7185 10.8600 11.7425 ;
      RECT 10.8360 12.0060 10.8600 12.0300 ;
      RECT 10.2120 11.0610 10.2360 11.0850 ;
      RECT 10.2120 11.8380 10.2360 11.8620 ;
      RECT 9.6000 11.7810 9.6240 11.8050 ;
      RECT 9.6000 11.9580 9.6240 11.9820 ;
      RECT 9.6000 12.9810 9.6240 13.0050 ;
      RECT 9.6000 13.0770 9.6240 13.1010 ;
      RECT 9.3840 11.3010 9.4080 11.3250 ;
      RECT 9.3840 12.3420 9.4080 12.3660 ;
      RECT 9.3840 12.6450 9.4080 12.6690 ;
      RECT 9.3840 12.7740 9.4080 12.7980 ;
      RECT 9.3840 13.1580 9.4080 13.1820 ;
      RECT 9.3840 13.3650 9.4080 13.3890 ;
      RECT 9.1680 11.2050 9.1920 11.2290 ;
      RECT 9.1680 12.4380 9.1920 12.4620 ;
      RECT 9.1680 12.6930 9.1920 12.7170 ;
      RECT 9.1680 12.8370 9.1920 12.8610 ;
      RECT 9.1680 13.0770 9.1920 13.1010 ;
      RECT 9.1680 13.3650 9.1920 13.3890 ;
      RECT 9.0600 13.7970 9.0840 13.8210 ;
      RECT 9.0600 14.1810 9.0840 14.2050 ;
      RECT 9.0600 16.4370 9.0840 16.4610 ;
      RECT 9.0600 16.5330 9.0840 16.5570 ;
      RECT 8.9700 9.9170 8.9940 9.9410 ;
      RECT 8.9700 12.6930 8.9940 12.7170 ;
      RECT 8.9700 18.5410 8.9940 18.5650 ;
      RECT 8.9220 9.8210 8.9460 9.8450 ;
      RECT 8.9220 12.8370 8.9460 12.8610 ;
      RECT 8.9220 18.4450 8.9460 18.4690 ;
      RECT 8.8740 9.7250 8.8980 9.7490 ;
      RECT 8.8740 12.2130 8.8980 12.2370 ;
      RECT 8.8740 18.2530 8.8980 18.2770 ;
      RECT 8.8260 9.6290 8.8500 9.6530 ;
      RECT 8.8260 14.9490 8.8500 14.9730 ;
      RECT 8.8260 17.6850 8.8500 17.7090 ;
      RECT 8.8260 18.1570 8.8500 18.1810 ;
      RECT 8.7780 9.5330 8.8020 9.5570 ;
      RECT 8.7780 12.9810 8.8020 13.0050 ;
      RECT 8.7780 18.4930 8.8020 18.5170 ;
      RECT 8.7300 9.8690 8.7540 9.8930 ;
      RECT 8.7300 13.7970 8.7540 13.8210 ;
      RECT 8.7300 18.3970 8.7540 18.4210 ;
      RECT 8.6820 9.7730 8.7060 9.7970 ;
      RECT 8.6820 12.2130 8.7060 12.2370 ;
      RECT 8.6820 18.3010 8.7060 18.3250 ;
      RECT 8.6340 9.4850 8.6580 9.5090 ;
      RECT 8.6340 16.4370 8.6580 16.4610 ;
      RECT 8.6340 18.2050 8.6580 18.2290 ;
      RECT 8.5860 9.3410 8.6100 9.3650 ;
      RECT 8.5860 15.5250 8.6100 15.5490 ;
      RECT 8.5860 18.1090 8.6100 18.1330 ;
      RECT 8.2980 10.0610 8.3220 10.0850 ;
      RECT 8.2980 13.7490 8.3220 13.7730 ;
      RECT 8.2980 17.9650 8.3220 17.9890 ;
      RECT 8.2500 9.9650 8.2740 9.9890 ;
      RECT 8.2500 14.1810 8.2740 14.2050 ;
      RECT 8.2500 18.5890 8.2740 18.6130 ;
      RECT 8.2020 9.4850 8.2260 9.5090 ;
      RECT 8.2020 13.3650 8.2260 13.3890 ;
      RECT 8.2020 18.6850 8.2260 18.7090 ;
      RECT 8.1060 9.5810 8.1300 9.6050 ;
      RECT 8.1060 15.9570 8.1300 15.9810 ;
      RECT 8.1060 18.5410 8.1300 18.5650 ;
      RECT 7.9140 9.9170 7.9380 9.9410 ;
      RECT 7.9140 14.5170 7.9380 14.5410 ;
      RECT 7.9140 18.6850 7.9380 18.7090 ;
      RECT 7.8660 9.8210 7.8900 9.8450 ;
      RECT 7.8660 17.6850 7.8900 17.7090 ;
      RECT 7.8660 18.2530 7.8900 18.2770 ;
      RECT 7.8180 9.7250 7.8420 9.7490 ;
      RECT 7.8180 16.5330 7.8420 16.5570 ;
      RECT 7.8180 18.5890 7.8420 18.6130 ;
      RECT 7.7700 9.6290 7.7940 9.6530 ;
      RECT 7.7700 16.1010 7.7940 16.1250 ;
      RECT 7.7700 18.1570 7.7940 18.1810 ;
      RECT 7.7220 9.5330 7.7460 9.5570 ;
      RECT 7.7220 13.3650 7.7460 13.3890 ;
      RECT 7.7220 18.4930 7.7460 18.5170 ;
      RECT 7.6740 9.7730 7.6980 9.7970 ;
      RECT 7.6740 13.0770 7.6980 13.1010 ;
      RECT 7.6740 18.3970 7.6980 18.4210 ;
      RECT 7.6260 9.6770 7.6500 9.7010 ;
      RECT 7.6260 14.3730 7.6500 14.3970 ;
      RECT 7.6260 18.3010 7.6500 18.3250 ;
      RECT 7.5780 9.5810 7.6020 9.6050 ;
      RECT 7.5780 14.2770 7.6020 14.3010 ;
      RECT 7.5780 18.2050 7.6020 18.2290 ;
      RECT 7.5300 9.4850 7.5540 9.5090 ;
      RECT 7.5300 11.5890 7.5540 11.6130 ;
      RECT 7.5300 18.1090 7.5540 18.1330 ;
      RECT 7.4400 14.2770 7.4640 14.3010 ;
      RECT 7.4400 14.3730 7.4640 14.3970 ;
      RECT 7.2720 10.0130 7.2960 10.0370 ;
      RECT 7.2720 13.7970 7.2960 13.8210 ;
      RECT 6.9000 11.5890 6.9240 11.6130 ;
      RECT 6.9000 11.7810 6.9240 11.8050 ;
  LAYER M5  ;
      RECT 11.0040 10.6180 11.0280 11.7050 ;
      RECT 10.8360 11.0330 10.8600 12.0935 ;
      RECT 10.2120 11.0415 10.2360 11.8740 ;
      RECT 9.6000 11.7700 9.6240 11.9930 ;
      RECT 9.6000 12.9700 9.6240 13.1120 ;
      RECT 9.3840 11.2900 9.4080 12.3770 ;
      RECT 9.3840 12.6340 9.4080 12.8090 ;
      RECT 9.3840 13.1470 9.4080 13.4000 ;
      RECT 9.1680 11.1940 9.1920 12.4730 ;
      RECT 9.1680 12.6820 9.1920 12.8720 ;
      RECT 9.1680 13.0660 9.1920 13.4000 ;
      RECT 9.0600 13.7860 9.0840 14.2160 ;
      RECT 9.0600 16.4260 9.0840 16.5680 ;
      RECT 8.9700 10.2540 8.9940 17.8370 ;
      RECT 8.9220 10.2540 8.9460 17.8370 ;
      RECT 8.8740 10.2540 8.8980 17.8370 ;
      RECT 8.8260 10.2540 8.8500 17.8370 ;
      RECT 8.7780 10.2540 8.8020 17.8370 ;
      RECT 8.7300 10.2540 8.7540 17.8370 ;
      RECT 8.6820 10.2540 8.7060 17.8370 ;
      RECT 8.6340 10.2540 8.6580 17.8370 ;
      RECT 8.5860 10.2540 8.6100 17.8370 ;
      RECT 8.2980 10.2540 8.3220 17.8370 ;
      RECT 8.2500 10.2540 8.2740 17.8370 ;
      RECT 8.2020 10.2540 8.2260 17.8370 ;
      RECT 8.1060 10.2540 8.1300 17.8370 ;
      RECT 7.9140 10.2540 7.9380 17.8370 ;
      RECT 7.8660 10.2540 7.8900 17.8370 ;
      RECT 7.8180 10.2540 7.8420 17.8370 ;
      RECT 7.7700 10.2540 7.7940 17.8370 ;
      RECT 7.7220 10.2540 7.7460 17.8370 ;
      RECT 7.6740 10.2540 7.6980 17.8370 ;
      RECT 7.6260 9.4120 7.6500 18.4670 ;
      RECT 7.5780 9.3750 7.6020 18.4210 ;
      RECT 7.5300 9.3210 7.5540 18.3670 ;
      RECT 7.4400 14.2660 7.4640 14.4080 ;
      RECT 7.2720 9.9950 7.2960 13.8390 ;
      RECT 6.9000 11.5780 6.9240 11.8160 ;
  LAYER M2  ;
    RECT 0.108 0.036 15.8920 28.0440 ;
  LAYER M1  ;
    RECT 0.108 0.036 15.8920 28.0440 ;
  END
END srambank_128x4x18_6t122 
