VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_64x4x34_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_64x4x34_6t122 0 0 ; 
  SIZE 38.448 BY 181.44 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.688 38.036 4.88 ; 
        RECT 0.404 9.008 38.036 9.2 ; 
        RECT 0.404 13.328 38.036 13.52 ; 
        RECT 0.404 17.648 38.036 17.84 ; 
        RECT 0.404 21.968 38.036 22.16 ; 
        RECT 0.404 26.288 38.036 26.48 ; 
        RECT 0.404 30.608 38.036 30.8 ; 
        RECT 0.404 34.928 38.036 35.12 ; 
        RECT 0.404 39.248 38.036 39.44 ; 
        RECT 0.404 43.568 38.036 43.76 ; 
        RECT 0.404 47.888 38.036 48.08 ; 
        RECT 0.404 52.208 38.036 52.4 ; 
        RECT 0.404 56.528 38.036 56.72 ; 
        RECT 0.404 60.848 38.036 61.04 ; 
        RECT 0.404 65.168 38.036 65.36 ; 
        RECT 0.404 69.488 38.036 69.68 ; 
        RECT 0.404 73.808 38.036 74 ; 
        RECT 0.432 75.756 38.016 76.62 ; 
        RECT 22.44 74.636 23.492 74.732 ; 
        RECT 22.964 89.772 23.412 89.868 ; 
        RECT 15.768 88.428 22.68 89.292 ; 
        RECT 15.768 101.1 22.68 101.964 ; 
        RECT 0.404 110.636 38.036 110.828 ; 
        RECT 0.404 114.956 38.036 115.148 ; 
        RECT 0.404 119.276 38.036 119.468 ; 
        RECT 0.404 123.596 38.036 123.788 ; 
        RECT 0.404 127.916 38.036 128.108 ; 
        RECT 0.404 132.236 38.036 132.428 ; 
        RECT 0.404 136.556 38.036 136.748 ; 
        RECT 0.404 140.876 38.036 141.068 ; 
        RECT 0.404 145.196 38.036 145.388 ; 
        RECT 0.404 149.516 38.036 149.708 ; 
        RECT 0.404 153.836 38.036 154.028 ; 
        RECT 0.404 158.156 38.036 158.348 ; 
        RECT 0.404 162.476 38.036 162.668 ; 
        RECT 0.404 166.796 38.036 166.988 ; 
        RECT 0.404 171.116 38.036 171.308 ; 
        RECT 0.404 175.436 38.036 175.628 ; 
        RECT 0.404 179.756 38.036 179.948 ; 
      LAYER M3 ; 
        RECT 37.908 0.866 37.98 5.506 ; 
        RECT 23.292 0.868 23.364 5.504 ; 
        RECT 17.676 1.012 18.036 5.468 ; 
        RECT 15.084 0.868 15.156 5.504 ; 
        RECT 0.468 0.866 0.54 5.506 ; 
        RECT 37.908 5.186 37.98 9.826 ; 
        RECT 23.292 5.188 23.364 9.824 ; 
        RECT 17.676 5.332 18.036 9.788 ; 
        RECT 15.084 5.188 15.156 9.824 ; 
        RECT 0.468 5.186 0.54 9.826 ; 
        RECT 37.908 9.506 37.98 14.146 ; 
        RECT 23.292 9.508 23.364 14.144 ; 
        RECT 17.676 9.652 18.036 14.108 ; 
        RECT 15.084 9.508 15.156 14.144 ; 
        RECT 0.468 9.506 0.54 14.146 ; 
        RECT 37.908 13.826 37.98 18.466 ; 
        RECT 23.292 13.828 23.364 18.464 ; 
        RECT 17.676 13.972 18.036 18.428 ; 
        RECT 15.084 13.828 15.156 18.464 ; 
        RECT 0.468 13.826 0.54 18.466 ; 
        RECT 37.908 18.146 37.98 22.786 ; 
        RECT 23.292 18.148 23.364 22.784 ; 
        RECT 17.676 18.292 18.036 22.748 ; 
        RECT 15.084 18.148 15.156 22.784 ; 
        RECT 0.468 18.146 0.54 22.786 ; 
        RECT 37.908 22.466 37.98 27.106 ; 
        RECT 23.292 22.468 23.364 27.104 ; 
        RECT 17.676 22.612 18.036 27.068 ; 
        RECT 15.084 22.468 15.156 27.104 ; 
        RECT 0.468 22.466 0.54 27.106 ; 
        RECT 37.908 26.786 37.98 31.426 ; 
        RECT 23.292 26.788 23.364 31.424 ; 
        RECT 17.676 26.932 18.036 31.388 ; 
        RECT 15.084 26.788 15.156 31.424 ; 
        RECT 0.468 26.786 0.54 31.426 ; 
        RECT 37.908 31.106 37.98 35.746 ; 
        RECT 23.292 31.108 23.364 35.744 ; 
        RECT 17.676 31.252 18.036 35.708 ; 
        RECT 15.084 31.108 15.156 35.744 ; 
        RECT 0.468 31.106 0.54 35.746 ; 
        RECT 37.908 35.426 37.98 40.066 ; 
        RECT 23.292 35.428 23.364 40.064 ; 
        RECT 17.676 35.572 18.036 40.028 ; 
        RECT 15.084 35.428 15.156 40.064 ; 
        RECT 0.468 35.426 0.54 40.066 ; 
        RECT 37.908 39.746 37.98 44.386 ; 
        RECT 23.292 39.748 23.364 44.384 ; 
        RECT 17.676 39.892 18.036 44.348 ; 
        RECT 15.084 39.748 15.156 44.384 ; 
        RECT 0.468 39.746 0.54 44.386 ; 
        RECT 37.908 44.066 37.98 48.706 ; 
        RECT 23.292 44.068 23.364 48.704 ; 
        RECT 17.676 44.212 18.036 48.668 ; 
        RECT 15.084 44.068 15.156 48.704 ; 
        RECT 0.468 44.066 0.54 48.706 ; 
        RECT 37.908 48.386 37.98 53.026 ; 
        RECT 23.292 48.388 23.364 53.024 ; 
        RECT 17.676 48.532 18.036 52.988 ; 
        RECT 15.084 48.388 15.156 53.024 ; 
        RECT 0.468 48.386 0.54 53.026 ; 
        RECT 37.908 52.706 37.98 57.346 ; 
        RECT 23.292 52.708 23.364 57.344 ; 
        RECT 17.676 52.852 18.036 57.308 ; 
        RECT 15.084 52.708 15.156 57.344 ; 
        RECT 0.468 52.706 0.54 57.346 ; 
        RECT 37.908 57.026 37.98 61.666 ; 
        RECT 23.292 57.028 23.364 61.664 ; 
        RECT 17.676 57.172 18.036 61.628 ; 
        RECT 15.084 57.028 15.156 61.664 ; 
        RECT 0.468 57.026 0.54 61.666 ; 
        RECT 37.908 61.346 37.98 65.986 ; 
        RECT 23.292 61.348 23.364 65.984 ; 
        RECT 17.676 61.492 18.036 65.948 ; 
        RECT 15.084 61.348 15.156 65.984 ; 
        RECT 0.468 61.346 0.54 65.986 ; 
        RECT 37.908 65.666 37.98 70.306 ; 
        RECT 23.292 65.668 23.364 70.304 ; 
        RECT 17.676 65.812 18.036 70.268 ; 
        RECT 15.084 65.668 15.156 70.304 ; 
        RECT 0.468 65.666 0.54 70.306 ; 
        RECT 37.908 69.986 37.98 74.626 ; 
        RECT 23.292 69.988 23.364 74.624 ; 
        RECT 17.676 70.132 18.036 74.588 ; 
        RECT 15.084 69.988 15.156 74.624 ; 
        RECT 0.468 69.986 0.54 74.626 ; 
        RECT 37.908 74.306 37.98 107.134 ; 
        RECT 23.292 74.624 23.364 74.99 ; 
        RECT 23.292 89.584 23.364 107.024 ; 
        RECT 17.82 75.6 18.756 105.932 ; 
        RECT 17.676 105.588 18.036 107.728 ; 
        RECT 17.676 74.48 18.036 76.62 ; 
        RECT 0.468 74.306 0.54 107.134 ; 
        RECT 37.908 106.814 37.98 111.454 ; 
        RECT 23.292 106.816 23.364 111.452 ; 
        RECT 17.676 106.96 18.036 111.416 ; 
        RECT 15.084 106.816 15.156 111.452 ; 
        RECT 0.468 106.814 0.54 111.454 ; 
        RECT 37.908 111.134 37.98 115.774 ; 
        RECT 23.292 111.136 23.364 115.772 ; 
        RECT 17.676 111.28 18.036 115.736 ; 
        RECT 15.084 111.136 15.156 115.772 ; 
        RECT 0.468 111.134 0.54 115.774 ; 
        RECT 37.908 115.454 37.98 120.094 ; 
        RECT 23.292 115.456 23.364 120.092 ; 
        RECT 17.676 115.6 18.036 120.056 ; 
        RECT 15.084 115.456 15.156 120.092 ; 
        RECT 0.468 115.454 0.54 120.094 ; 
        RECT 37.908 119.774 37.98 124.414 ; 
        RECT 23.292 119.776 23.364 124.412 ; 
        RECT 17.676 119.92 18.036 124.376 ; 
        RECT 15.084 119.776 15.156 124.412 ; 
        RECT 0.468 119.774 0.54 124.414 ; 
        RECT 37.908 124.094 37.98 128.734 ; 
        RECT 23.292 124.096 23.364 128.732 ; 
        RECT 17.676 124.24 18.036 128.696 ; 
        RECT 15.084 124.096 15.156 128.732 ; 
        RECT 0.468 124.094 0.54 128.734 ; 
        RECT 37.908 128.414 37.98 133.054 ; 
        RECT 23.292 128.416 23.364 133.052 ; 
        RECT 17.676 128.56 18.036 133.016 ; 
        RECT 15.084 128.416 15.156 133.052 ; 
        RECT 0.468 128.414 0.54 133.054 ; 
        RECT 37.908 132.734 37.98 137.374 ; 
        RECT 23.292 132.736 23.364 137.372 ; 
        RECT 17.676 132.88 18.036 137.336 ; 
        RECT 15.084 132.736 15.156 137.372 ; 
        RECT 0.468 132.734 0.54 137.374 ; 
        RECT 37.908 137.054 37.98 141.694 ; 
        RECT 23.292 137.056 23.364 141.692 ; 
        RECT 17.676 137.2 18.036 141.656 ; 
        RECT 15.084 137.056 15.156 141.692 ; 
        RECT 0.468 137.054 0.54 141.694 ; 
        RECT 37.908 141.374 37.98 146.014 ; 
        RECT 23.292 141.376 23.364 146.012 ; 
        RECT 17.676 141.52 18.036 145.976 ; 
        RECT 15.084 141.376 15.156 146.012 ; 
        RECT 0.468 141.374 0.54 146.014 ; 
        RECT 37.908 145.694 37.98 150.334 ; 
        RECT 23.292 145.696 23.364 150.332 ; 
        RECT 17.676 145.84 18.036 150.296 ; 
        RECT 15.084 145.696 15.156 150.332 ; 
        RECT 0.468 145.694 0.54 150.334 ; 
        RECT 37.908 150.014 37.98 154.654 ; 
        RECT 23.292 150.016 23.364 154.652 ; 
        RECT 17.676 150.16 18.036 154.616 ; 
        RECT 15.084 150.016 15.156 154.652 ; 
        RECT 0.468 150.014 0.54 154.654 ; 
        RECT 37.908 154.334 37.98 158.974 ; 
        RECT 23.292 154.336 23.364 158.972 ; 
        RECT 17.676 154.48 18.036 158.936 ; 
        RECT 15.084 154.336 15.156 158.972 ; 
        RECT 0.468 154.334 0.54 158.974 ; 
        RECT 37.908 158.654 37.98 163.294 ; 
        RECT 23.292 158.656 23.364 163.292 ; 
        RECT 17.676 158.8 18.036 163.256 ; 
        RECT 15.084 158.656 15.156 163.292 ; 
        RECT 0.468 158.654 0.54 163.294 ; 
        RECT 37.908 162.974 37.98 167.614 ; 
        RECT 23.292 162.976 23.364 167.612 ; 
        RECT 17.676 163.12 18.036 167.576 ; 
        RECT 15.084 162.976 15.156 167.612 ; 
        RECT 0.468 162.974 0.54 167.614 ; 
        RECT 37.908 167.294 37.98 171.934 ; 
        RECT 23.292 167.296 23.364 171.932 ; 
        RECT 17.676 167.44 18.036 171.896 ; 
        RECT 15.084 167.296 15.156 171.932 ; 
        RECT 0.468 167.294 0.54 171.934 ; 
        RECT 37.908 171.614 37.98 176.254 ; 
        RECT 23.292 171.616 23.364 176.252 ; 
        RECT 17.676 171.76 18.036 176.216 ; 
        RECT 15.084 171.616 15.156 176.252 ; 
        RECT 0.468 171.614 0.54 176.254 ; 
        RECT 37.908 175.934 37.98 180.574 ; 
        RECT 23.292 175.936 23.364 180.572 ; 
        RECT 17.676 176.08 18.036 180.536 ; 
        RECT 15.084 175.936 15.156 180.572 ; 
        RECT 0.468 175.934 0.54 180.574 ; 
      LAYER V3 ; 
        RECT 0.468 4.688 0.54 4.88 ; 
        RECT 15.084 4.688 15.156 4.88 ; 
        RECT 17.676 4.688 18.036 4.88 ; 
        RECT 23.292 4.688 23.364 4.88 ; 
        RECT 37.908 4.688 37.98 4.88 ; 
        RECT 0.468 9.008 0.54 9.2 ; 
        RECT 15.084 9.008 15.156 9.2 ; 
        RECT 17.676 9.008 18.036 9.2 ; 
        RECT 23.292 9.008 23.364 9.2 ; 
        RECT 37.908 9.008 37.98 9.2 ; 
        RECT 0.468 13.328 0.54 13.52 ; 
        RECT 15.084 13.328 15.156 13.52 ; 
        RECT 17.676 13.328 18.036 13.52 ; 
        RECT 23.292 13.328 23.364 13.52 ; 
        RECT 37.908 13.328 37.98 13.52 ; 
        RECT 0.468 17.648 0.54 17.84 ; 
        RECT 15.084 17.648 15.156 17.84 ; 
        RECT 17.676 17.648 18.036 17.84 ; 
        RECT 23.292 17.648 23.364 17.84 ; 
        RECT 37.908 17.648 37.98 17.84 ; 
        RECT 0.468 21.968 0.54 22.16 ; 
        RECT 15.084 21.968 15.156 22.16 ; 
        RECT 17.676 21.968 18.036 22.16 ; 
        RECT 23.292 21.968 23.364 22.16 ; 
        RECT 37.908 21.968 37.98 22.16 ; 
        RECT 0.468 26.288 0.54 26.48 ; 
        RECT 15.084 26.288 15.156 26.48 ; 
        RECT 17.676 26.288 18.036 26.48 ; 
        RECT 23.292 26.288 23.364 26.48 ; 
        RECT 37.908 26.288 37.98 26.48 ; 
        RECT 0.468 30.608 0.54 30.8 ; 
        RECT 15.084 30.608 15.156 30.8 ; 
        RECT 17.676 30.608 18.036 30.8 ; 
        RECT 23.292 30.608 23.364 30.8 ; 
        RECT 37.908 30.608 37.98 30.8 ; 
        RECT 0.468 34.928 0.54 35.12 ; 
        RECT 15.084 34.928 15.156 35.12 ; 
        RECT 17.676 34.928 18.036 35.12 ; 
        RECT 23.292 34.928 23.364 35.12 ; 
        RECT 37.908 34.928 37.98 35.12 ; 
        RECT 0.468 39.248 0.54 39.44 ; 
        RECT 15.084 39.248 15.156 39.44 ; 
        RECT 17.676 39.248 18.036 39.44 ; 
        RECT 23.292 39.248 23.364 39.44 ; 
        RECT 37.908 39.248 37.98 39.44 ; 
        RECT 0.468 43.568 0.54 43.76 ; 
        RECT 15.084 43.568 15.156 43.76 ; 
        RECT 17.676 43.568 18.036 43.76 ; 
        RECT 23.292 43.568 23.364 43.76 ; 
        RECT 37.908 43.568 37.98 43.76 ; 
        RECT 0.468 47.888 0.54 48.08 ; 
        RECT 15.084 47.888 15.156 48.08 ; 
        RECT 17.676 47.888 18.036 48.08 ; 
        RECT 23.292 47.888 23.364 48.08 ; 
        RECT 37.908 47.888 37.98 48.08 ; 
        RECT 0.468 52.208 0.54 52.4 ; 
        RECT 15.084 52.208 15.156 52.4 ; 
        RECT 17.676 52.208 18.036 52.4 ; 
        RECT 23.292 52.208 23.364 52.4 ; 
        RECT 37.908 52.208 37.98 52.4 ; 
        RECT 0.468 56.528 0.54 56.72 ; 
        RECT 15.084 56.528 15.156 56.72 ; 
        RECT 17.676 56.528 18.036 56.72 ; 
        RECT 23.292 56.528 23.364 56.72 ; 
        RECT 37.908 56.528 37.98 56.72 ; 
        RECT 0.468 60.848 0.54 61.04 ; 
        RECT 15.084 60.848 15.156 61.04 ; 
        RECT 17.676 60.848 18.036 61.04 ; 
        RECT 23.292 60.848 23.364 61.04 ; 
        RECT 37.908 60.848 37.98 61.04 ; 
        RECT 0.468 65.168 0.54 65.36 ; 
        RECT 15.084 65.168 15.156 65.36 ; 
        RECT 17.676 65.168 18.036 65.36 ; 
        RECT 23.292 65.168 23.364 65.36 ; 
        RECT 37.908 65.168 37.98 65.36 ; 
        RECT 0.468 69.488 0.54 69.68 ; 
        RECT 15.084 69.488 15.156 69.68 ; 
        RECT 17.676 69.488 18.036 69.68 ; 
        RECT 23.292 69.488 23.364 69.68 ; 
        RECT 37.908 69.488 37.98 69.68 ; 
        RECT 0.468 73.808 0.54 74 ; 
        RECT 15.084 73.808 15.156 74 ; 
        RECT 17.676 73.808 18.036 74 ; 
        RECT 23.292 73.808 23.364 74 ; 
        RECT 37.908 73.808 37.98 74 ; 
        RECT 0.468 75.756 0.54 76.62 ; 
        RECT 17.836 101.1 17.908 101.964 ; 
        RECT 17.836 88.428 17.908 89.292 ; 
        RECT 17.836 75.756 17.908 76.62 ; 
        RECT 18.044 101.1 18.116 101.964 ; 
        RECT 18.044 88.428 18.116 89.292 ; 
        RECT 18.044 75.756 18.116 76.62 ; 
        RECT 18.252 101.1 18.324 101.964 ; 
        RECT 18.252 88.428 18.324 89.292 ; 
        RECT 18.252 75.756 18.324 76.62 ; 
        RECT 18.46 101.1 18.532 101.964 ; 
        RECT 18.46 88.428 18.532 89.292 ; 
        RECT 18.46 75.756 18.532 76.62 ; 
        RECT 18.668 101.1 18.74 101.964 ; 
        RECT 18.668 88.428 18.74 89.292 ; 
        RECT 18.668 75.756 18.74 76.62 ; 
        RECT 23.292 89.772 23.364 89.868 ; 
        RECT 23.292 74.636 23.364 74.732 ; 
        RECT 0.468 110.636 0.54 110.828 ; 
        RECT 15.084 110.636 15.156 110.828 ; 
        RECT 17.676 110.636 18.036 110.828 ; 
        RECT 23.292 110.636 23.364 110.828 ; 
        RECT 37.908 110.636 37.98 110.828 ; 
        RECT 0.468 114.956 0.54 115.148 ; 
        RECT 15.084 114.956 15.156 115.148 ; 
        RECT 17.676 114.956 18.036 115.148 ; 
        RECT 23.292 114.956 23.364 115.148 ; 
        RECT 37.908 114.956 37.98 115.148 ; 
        RECT 0.468 119.276 0.54 119.468 ; 
        RECT 15.084 119.276 15.156 119.468 ; 
        RECT 17.676 119.276 18.036 119.468 ; 
        RECT 23.292 119.276 23.364 119.468 ; 
        RECT 37.908 119.276 37.98 119.468 ; 
        RECT 0.468 123.596 0.54 123.788 ; 
        RECT 15.084 123.596 15.156 123.788 ; 
        RECT 17.676 123.596 18.036 123.788 ; 
        RECT 23.292 123.596 23.364 123.788 ; 
        RECT 37.908 123.596 37.98 123.788 ; 
        RECT 0.468 127.916 0.54 128.108 ; 
        RECT 15.084 127.916 15.156 128.108 ; 
        RECT 17.676 127.916 18.036 128.108 ; 
        RECT 23.292 127.916 23.364 128.108 ; 
        RECT 37.908 127.916 37.98 128.108 ; 
        RECT 0.468 132.236 0.54 132.428 ; 
        RECT 15.084 132.236 15.156 132.428 ; 
        RECT 17.676 132.236 18.036 132.428 ; 
        RECT 23.292 132.236 23.364 132.428 ; 
        RECT 37.908 132.236 37.98 132.428 ; 
        RECT 0.468 136.556 0.54 136.748 ; 
        RECT 15.084 136.556 15.156 136.748 ; 
        RECT 17.676 136.556 18.036 136.748 ; 
        RECT 23.292 136.556 23.364 136.748 ; 
        RECT 37.908 136.556 37.98 136.748 ; 
        RECT 0.468 140.876 0.54 141.068 ; 
        RECT 15.084 140.876 15.156 141.068 ; 
        RECT 17.676 140.876 18.036 141.068 ; 
        RECT 23.292 140.876 23.364 141.068 ; 
        RECT 37.908 140.876 37.98 141.068 ; 
        RECT 0.468 145.196 0.54 145.388 ; 
        RECT 15.084 145.196 15.156 145.388 ; 
        RECT 17.676 145.196 18.036 145.388 ; 
        RECT 23.292 145.196 23.364 145.388 ; 
        RECT 37.908 145.196 37.98 145.388 ; 
        RECT 0.468 149.516 0.54 149.708 ; 
        RECT 15.084 149.516 15.156 149.708 ; 
        RECT 17.676 149.516 18.036 149.708 ; 
        RECT 23.292 149.516 23.364 149.708 ; 
        RECT 37.908 149.516 37.98 149.708 ; 
        RECT 0.468 153.836 0.54 154.028 ; 
        RECT 15.084 153.836 15.156 154.028 ; 
        RECT 17.676 153.836 18.036 154.028 ; 
        RECT 23.292 153.836 23.364 154.028 ; 
        RECT 37.908 153.836 37.98 154.028 ; 
        RECT 0.468 158.156 0.54 158.348 ; 
        RECT 15.084 158.156 15.156 158.348 ; 
        RECT 17.676 158.156 18.036 158.348 ; 
        RECT 23.292 158.156 23.364 158.348 ; 
        RECT 37.908 158.156 37.98 158.348 ; 
        RECT 0.468 162.476 0.54 162.668 ; 
        RECT 15.084 162.476 15.156 162.668 ; 
        RECT 17.676 162.476 18.036 162.668 ; 
        RECT 23.292 162.476 23.364 162.668 ; 
        RECT 37.908 162.476 37.98 162.668 ; 
        RECT 0.468 166.796 0.54 166.988 ; 
        RECT 15.084 166.796 15.156 166.988 ; 
        RECT 17.676 166.796 18.036 166.988 ; 
        RECT 23.292 166.796 23.364 166.988 ; 
        RECT 37.908 166.796 37.98 166.988 ; 
        RECT 0.468 171.116 0.54 171.308 ; 
        RECT 15.084 171.116 15.156 171.308 ; 
        RECT 17.676 171.116 18.036 171.308 ; 
        RECT 23.292 171.116 23.364 171.308 ; 
        RECT 37.908 171.116 37.98 171.308 ; 
        RECT 0.468 175.436 0.54 175.628 ; 
        RECT 15.084 175.436 15.156 175.628 ; 
        RECT 17.676 175.436 18.036 175.628 ; 
        RECT 23.292 175.436 23.364 175.628 ; 
        RECT 37.908 175.436 37.98 175.628 ; 
        RECT 0.468 179.756 0.54 179.948 ; 
        RECT 15.084 179.756 15.156 179.948 ; 
        RECT 17.676 179.756 18.036 179.948 ; 
        RECT 23.292 179.756 23.364 179.948 ; 
        RECT 37.908 179.756 37.98 179.948 ; 
      LAYER M5 ; 
        RECT 23.036 74.564 23.132 89.94 ; 
      LAYER V4 ; 
        RECT 23.036 89.772 23.132 89.868 ; 
        RECT 23.036 74.636 23.132 74.732 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.404 4.304 38.016 4.496 ; 
        RECT 0.404 8.624 38.016 8.816 ; 
        RECT 0.404 12.944 38.016 13.136 ; 
        RECT 0.404 17.264 38.016 17.456 ; 
        RECT 0.404 21.584 38.016 21.776 ; 
        RECT 0.404 25.904 38.016 26.096 ; 
        RECT 0.404 30.224 38.016 30.416 ; 
        RECT 0.404 34.544 38.016 34.736 ; 
        RECT 0.404 38.864 38.016 39.056 ; 
        RECT 0.404 43.184 38.016 43.376 ; 
        RECT 0.404 47.504 38.016 47.696 ; 
        RECT 0.404 51.824 38.016 52.016 ; 
        RECT 0.404 56.144 38.016 56.336 ; 
        RECT 0.404 60.464 38.016 60.656 ; 
        RECT 0.404 64.784 38.016 64.976 ; 
        RECT 0.404 69.104 38.016 69.296 ; 
        RECT 0.404 73.424 38.016 73.616 ; 
        RECT 0.432 77.484 38.016 78.348 ; 
        RECT 15.768 90.156 22.68 91.02 ; 
        RECT 15.768 102.828 22.68 103.692 ; 
        RECT 0.404 110.252 38.016 110.444 ; 
        RECT 0.404 114.572 38.016 114.764 ; 
        RECT 0.404 118.892 38.016 119.084 ; 
        RECT 0.404 123.212 38.016 123.404 ; 
        RECT 0.404 127.532 38.016 127.724 ; 
        RECT 0.404 131.852 38.016 132.044 ; 
        RECT 0.404 136.172 38.016 136.364 ; 
        RECT 0.404 140.492 38.016 140.684 ; 
        RECT 0.404 144.812 38.016 145.004 ; 
        RECT 0.404 149.132 38.016 149.324 ; 
        RECT 0.404 153.452 38.016 153.644 ; 
        RECT 0.404 157.772 38.016 157.964 ; 
        RECT 0.404 162.092 38.016 162.284 ; 
        RECT 0.404 166.412 38.016 166.604 ; 
        RECT 0.404 170.732 38.016 170.924 ; 
        RECT 0.404 175.052 38.016 175.244 ; 
        RECT 0.404 179.372 38.016 179.564 ; 
      LAYER M3 ; 
        RECT 37.764 0.866 37.836 5.506 ; 
        RECT 23.508 0.866 23.58 5.506 ; 
        RECT 20.448 1.012 20.592 5.468 ; 
        RECT 19.836 1.012 19.944 5.468 ; 
        RECT 14.868 0.866 14.94 5.506 ; 
        RECT 0.612 0.866 0.684 5.506 ; 
        RECT 37.764 5.186 37.836 9.826 ; 
        RECT 23.508 5.186 23.58 9.826 ; 
        RECT 20.448 5.332 20.592 9.788 ; 
        RECT 19.836 5.332 19.944 9.788 ; 
        RECT 14.868 5.186 14.94 9.826 ; 
        RECT 0.612 5.186 0.684 9.826 ; 
        RECT 37.764 9.506 37.836 14.146 ; 
        RECT 23.508 9.506 23.58 14.146 ; 
        RECT 20.448 9.652 20.592 14.108 ; 
        RECT 19.836 9.652 19.944 14.108 ; 
        RECT 14.868 9.506 14.94 14.146 ; 
        RECT 0.612 9.506 0.684 14.146 ; 
        RECT 37.764 13.826 37.836 18.466 ; 
        RECT 23.508 13.826 23.58 18.466 ; 
        RECT 20.448 13.972 20.592 18.428 ; 
        RECT 19.836 13.972 19.944 18.428 ; 
        RECT 14.868 13.826 14.94 18.466 ; 
        RECT 0.612 13.826 0.684 18.466 ; 
        RECT 37.764 18.146 37.836 22.786 ; 
        RECT 23.508 18.146 23.58 22.786 ; 
        RECT 20.448 18.292 20.592 22.748 ; 
        RECT 19.836 18.292 19.944 22.748 ; 
        RECT 14.868 18.146 14.94 22.786 ; 
        RECT 0.612 18.146 0.684 22.786 ; 
        RECT 37.764 22.466 37.836 27.106 ; 
        RECT 23.508 22.466 23.58 27.106 ; 
        RECT 20.448 22.612 20.592 27.068 ; 
        RECT 19.836 22.612 19.944 27.068 ; 
        RECT 14.868 22.466 14.94 27.106 ; 
        RECT 0.612 22.466 0.684 27.106 ; 
        RECT 37.764 26.786 37.836 31.426 ; 
        RECT 23.508 26.786 23.58 31.426 ; 
        RECT 20.448 26.932 20.592 31.388 ; 
        RECT 19.836 26.932 19.944 31.388 ; 
        RECT 14.868 26.786 14.94 31.426 ; 
        RECT 0.612 26.786 0.684 31.426 ; 
        RECT 37.764 31.106 37.836 35.746 ; 
        RECT 23.508 31.106 23.58 35.746 ; 
        RECT 20.448 31.252 20.592 35.708 ; 
        RECT 19.836 31.252 19.944 35.708 ; 
        RECT 14.868 31.106 14.94 35.746 ; 
        RECT 0.612 31.106 0.684 35.746 ; 
        RECT 37.764 35.426 37.836 40.066 ; 
        RECT 23.508 35.426 23.58 40.066 ; 
        RECT 20.448 35.572 20.592 40.028 ; 
        RECT 19.836 35.572 19.944 40.028 ; 
        RECT 14.868 35.426 14.94 40.066 ; 
        RECT 0.612 35.426 0.684 40.066 ; 
        RECT 37.764 39.746 37.836 44.386 ; 
        RECT 23.508 39.746 23.58 44.386 ; 
        RECT 20.448 39.892 20.592 44.348 ; 
        RECT 19.836 39.892 19.944 44.348 ; 
        RECT 14.868 39.746 14.94 44.386 ; 
        RECT 0.612 39.746 0.684 44.386 ; 
        RECT 37.764 44.066 37.836 48.706 ; 
        RECT 23.508 44.066 23.58 48.706 ; 
        RECT 20.448 44.212 20.592 48.668 ; 
        RECT 19.836 44.212 19.944 48.668 ; 
        RECT 14.868 44.066 14.94 48.706 ; 
        RECT 0.612 44.066 0.684 48.706 ; 
        RECT 37.764 48.386 37.836 53.026 ; 
        RECT 23.508 48.386 23.58 53.026 ; 
        RECT 20.448 48.532 20.592 52.988 ; 
        RECT 19.836 48.532 19.944 52.988 ; 
        RECT 14.868 48.386 14.94 53.026 ; 
        RECT 0.612 48.386 0.684 53.026 ; 
        RECT 37.764 52.706 37.836 57.346 ; 
        RECT 23.508 52.706 23.58 57.346 ; 
        RECT 20.448 52.852 20.592 57.308 ; 
        RECT 19.836 52.852 19.944 57.308 ; 
        RECT 14.868 52.706 14.94 57.346 ; 
        RECT 0.612 52.706 0.684 57.346 ; 
        RECT 37.764 57.026 37.836 61.666 ; 
        RECT 23.508 57.026 23.58 61.666 ; 
        RECT 20.448 57.172 20.592 61.628 ; 
        RECT 19.836 57.172 19.944 61.628 ; 
        RECT 14.868 57.026 14.94 61.666 ; 
        RECT 0.612 57.026 0.684 61.666 ; 
        RECT 37.764 61.346 37.836 65.986 ; 
        RECT 23.508 61.346 23.58 65.986 ; 
        RECT 20.448 61.492 20.592 65.948 ; 
        RECT 19.836 61.492 19.944 65.948 ; 
        RECT 14.868 61.346 14.94 65.986 ; 
        RECT 0.612 61.346 0.684 65.986 ; 
        RECT 37.764 65.666 37.836 70.306 ; 
        RECT 23.508 65.666 23.58 70.306 ; 
        RECT 20.448 65.812 20.592 70.268 ; 
        RECT 19.836 65.812 19.944 70.268 ; 
        RECT 14.868 65.666 14.94 70.306 ; 
        RECT 0.612 65.666 0.684 70.306 ; 
        RECT 37.764 69.986 37.836 74.626 ; 
        RECT 23.508 69.986 23.58 74.626 ; 
        RECT 20.448 70.132 20.592 74.588 ; 
        RECT 19.836 70.132 19.944 74.588 ; 
        RECT 14.868 69.986 14.94 74.626 ; 
        RECT 0.612 69.986 0.684 74.626 ; 
        RECT 37.764 74.306 37.836 107.134 ; 
        RECT 23.508 74.306 23.58 107.134 ; 
        RECT 19.692 75.2 20.628 105.932 ; 
        RECT 20.448 74.48 20.592 107.028 ; 
        RECT 19.836 74.48 19.944 107.016 ; 
        RECT 14.868 74.306 14.94 107.134 ; 
        RECT 0.612 74.306 0.684 107.134 ; 
        RECT 37.764 106.814 37.836 111.454 ; 
        RECT 23.508 106.814 23.58 111.454 ; 
        RECT 20.448 106.96 20.592 111.416 ; 
        RECT 19.836 106.96 19.944 111.416 ; 
        RECT 14.868 106.814 14.94 111.454 ; 
        RECT 0.612 106.814 0.684 111.454 ; 
        RECT 37.764 111.134 37.836 115.774 ; 
        RECT 23.508 111.134 23.58 115.774 ; 
        RECT 20.448 111.28 20.592 115.736 ; 
        RECT 19.836 111.28 19.944 115.736 ; 
        RECT 14.868 111.134 14.94 115.774 ; 
        RECT 0.612 111.134 0.684 115.774 ; 
        RECT 37.764 115.454 37.836 120.094 ; 
        RECT 23.508 115.454 23.58 120.094 ; 
        RECT 20.448 115.6 20.592 120.056 ; 
        RECT 19.836 115.6 19.944 120.056 ; 
        RECT 14.868 115.454 14.94 120.094 ; 
        RECT 0.612 115.454 0.684 120.094 ; 
        RECT 37.764 119.774 37.836 124.414 ; 
        RECT 23.508 119.774 23.58 124.414 ; 
        RECT 20.448 119.92 20.592 124.376 ; 
        RECT 19.836 119.92 19.944 124.376 ; 
        RECT 14.868 119.774 14.94 124.414 ; 
        RECT 0.612 119.774 0.684 124.414 ; 
        RECT 37.764 124.094 37.836 128.734 ; 
        RECT 23.508 124.094 23.58 128.734 ; 
        RECT 20.448 124.24 20.592 128.696 ; 
        RECT 19.836 124.24 19.944 128.696 ; 
        RECT 14.868 124.094 14.94 128.734 ; 
        RECT 0.612 124.094 0.684 128.734 ; 
        RECT 37.764 128.414 37.836 133.054 ; 
        RECT 23.508 128.414 23.58 133.054 ; 
        RECT 20.448 128.56 20.592 133.016 ; 
        RECT 19.836 128.56 19.944 133.016 ; 
        RECT 14.868 128.414 14.94 133.054 ; 
        RECT 0.612 128.414 0.684 133.054 ; 
        RECT 37.764 132.734 37.836 137.374 ; 
        RECT 23.508 132.734 23.58 137.374 ; 
        RECT 20.448 132.88 20.592 137.336 ; 
        RECT 19.836 132.88 19.944 137.336 ; 
        RECT 14.868 132.734 14.94 137.374 ; 
        RECT 0.612 132.734 0.684 137.374 ; 
        RECT 37.764 137.054 37.836 141.694 ; 
        RECT 23.508 137.054 23.58 141.694 ; 
        RECT 20.448 137.2 20.592 141.656 ; 
        RECT 19.836 137.2 19.944 141.656 ; 
        RECT 14.868 137.054 14.94 141.694 ; 
        RECT 0.612 137.054 0.684 141.694 ; 
        RECT 37.764 141.374 37.836 146.014 ; 
        RECT 23.508 141.374 23.58 146.014 ; 
        RECT 20.448 141.52 20.592 145.976 ; 
        RECT 19.836 141.52 19.944 145.976 ; 
        RECT 14.868 141.374 14.94 146.014 ; 
        RECT 0.612 141.374 0.684 146.014 ; 
        RECT 37.764 145.694 37.836 150.334 ; 
        RECT 23.508 145.694 23.58 150.334 ; 
        RECT 20.448 145.84 20.592 150.296 ; 
        RECT 19.836 145.84 19.944 150.296 ; 
        RECT 14.868 145.694 14.94 150.334 ; 
        RECT 0.612 145.694 0.684 150.334 ; 
        RECT 37.764 150.014 37.836 154.654 ; 
        RECT 23.508 150.014 23.58 154.654 ; 
        RECT 20.448 150.16 20.592 154.616 ; 
        RECT 19.836 150.16 19.944 154.616 ; 
        RECT 14.868 150.014 14.94 154.654 ; 
        RECT 0.612 150.014 0.684 154.654 ; 
        RECT 37.764 154.334 37.836 158.974 ; 
        RECT 23.508 154.334 23.58 158.974 ; 
        RECT 20.448 154.48 20.592 158.936 ; 
        RECT 19.836 154.48 19.944 158.936 ; 
        RECT 14.868 154.334 14.94 158.974 ; 
        RECT 0.612 154.334 0.684 158.974 ; 
        RECT 37.764 158.654 37.836 163.294 ; 
        RECT 23.508 158.654 23.58 163.294 ; 
        RECT 20.448 158.8 20.592 163.256 ; 
        RECT 19.836 158.8 19.944 163.256 ; 
        RECT 14.868 158.654 14.94 163.294 ; 
        RECT 0.612 158.654 0.684 163.294 ; 
        RECT 37.764 162.974 37.836 167.614 ; 
        RECT 23.508 162.974 23.58 167.614 ; 
        RECT 20.448 163.12 20.592 167.576 ; 
        RECT 19.836 163.12 19.944 167.576 ; 
        RECT 14.868 162.974 14.94 167.614 ; 
        RECT 0.612 162.974 0.684 167.614 ; 
        RECT 37.764 167.294 37.836 171.934 ; 
        RECT 23.508 167.294 23.58 171.934 ; 
        RECT 20.448 167.44 20.592 171.896 ; 
        RECT 19.836 167.44 19.944 171.896 ; 
        RECT 14.868 167.294 14.94 171.934 ; 
        RECT 0.612 167.294 0.684 171.934 ; 
        RECT 37.764 171.614 37.836 176.254 ; 
        RECT 23.508 171.614 23.58 176.254 ; 
        RECT 20.448 171.76 20.592 176.216 ; 
        RECT 19.836 171.76 19.944 176.216 ; 
        RECT 14.868 171.614 14.94 176.254 ; 
        RECT 0.612 171.614 0.684 176.254 ; 
        RECT 37.764 175.934 37.836 180.574 ; 
        RECT 23.508 175.934 23.58 180.574 ; 
        RECT 20.448 176.08 20.592 180.536 ; 
        RECT 19.836 176.08 19.944 180.536 ; 
        RECT 14.868 175.934 14.94 180.574 ; 
        RECT 0.612 175.934 0.684 180.574 ; 
      LAYER V3 ; 
        RECT 0.612 4.304 0.684 4.496 ; 
        RECT 14.868 4.304 14.94 4.496 ; 
        RECT 19.836 4.304 19.944 4.496 ; 
        RECT 20.448 4.304 20.592 4.496 ; 
        RECT 23.508 4.304 23.58 4.496 ; 
        RECT 37.764 4.304 37.836 4.496 ; 
        RECT 0.612 8.624 0.684 8.816 ; 
        RECT 14.868 8.624 14.94 8.816 ; 
        RECT 19.836 8.624 19.944 8.816 ; 
        RECT 20.448 8.624 20.592 8.816 ; 
        RECT 23.508 8.624 23.58 8.816 ; 
        RECT 37.764 8.624 37.836 8.816 ; 
        RECT 0.612 12.944 0.684 13.136 ; 
        RECT 14.868 12.944 14.94 13.136 ; 
        RECT 19.836 12.944 19.944 13.136 ; 
        RECT 20.448 12.944 20.592 13.136 ; 
        RECT 23.508 12.944 23.58 13.136 ; 
        RECT 37.764 12.944 37.836 13.136 ; 
        RECT 0.612 17.264 0.684 17.456 ; 
        RECT 14.868 17.264 14.94 17.456 ; 
        RECT 19.836 17.264 19.944 17.456 ; 
        RECT 20.448 17.264 20.592 17.456 ; 
        RECT 23.508 17.264 23.58 17.456 ; 
        RECT 37.764 17.264 37.836 17.456 ; 
        RECT 0.612 21.584 0.684 21.776 ; 
        RECT 14.868 21.584 14.94 21.776 ; 
        RECT 19.836 21.584 19.944 21.776 ; 
        RECT 20.448 21.584 20.592 21.776 ; 
        RECT 23.508 21.584 23.58 21.776 ; 
        RECT 37.764 21.584 37.836 21.776 ; 
        RECT 0.612 25.904 0.684 26.096 ; 
        RECT 14.868 25.904 14.94 26.096 ; 
        RECT 19.836 25.904 19.944 26.096 ; 
        RECT 20.448 25.904 20.592 26.096 ; 
        RECT 23.508 25.904 23.58 26.096 ; 
        RECT 37.764 25.904 37.836 26.096 ; 
        RECT 0.612 30.224 0.684 30.416 ; 
        RECT 14.868 30.224 14.94 30.416 ; 
        RECT 19.836 30.224 19.944 30.416 ; 
        RECT 20.448 30.224 20.592 30.416 ; 
        RECT 23.508 30.224 23.58 30.416 ; 
        RECT 37.764 30.224 37.836 30.416 ; 
        RECT 0.612 34.544 0.684 34.736 ; 
        RECT 14.868 34.544 14.94 34.736 ; 
        RECT 19.836 34.544 19.944 34.736 ; 
        RECT 20.448 34.544 20.592 34.736 ; 
        RECT 23.508 34.544 23.58 34.736 ; 
        RECT 37.764 34.544 37.836 34.736 ; 
        RECT 0.612 38.864 0.684 39.056 ; 
        RECT 14.868 38.864 14.94 39.056 ; 
        RECT 19.836 38.864 19.944 39.056 ; 
        RECT 20.448 38.864 20.592 39.056 ; 
        RECT 23.508 38.864 23.58 39.056 ; 
        RECT 37.764 38.864 37.836 39.056 ; 
        RECT 0.612 43.184 0.684 43.376 ; 
        RECT 14.868 43.184 14.94 43.376 ; 
        RECT 19.836 43.184 19.944 43.376 ; 
        RECT 20.448 43.184 20.592 43.376 ; 
        RECT 23.508 43.184 23.58 43.376 ; 
        RECT 37.764 43.184 37.836 43.376 ; 
        RECT 0.612 47.504 0.684 47.696 ; 
        RECT 14.868 47.504 14.94 47.696 ; 
        RECT 19.836 47.504 19.944 47.696 ; 
        RECT 20.448 47.504 20.592 47.696 ; 
        RECT 23.508 47.504 23.58 47.696 ; 
        RECT 37.764 47.504 37.836 47.696 ; 
        RECT 0.612 51.824 0.684 52.016 ; 
        RECT 14.868 51.824 14.94 52.016 ; 
        RECT 19.836 51.824 19.944 52.016 ; 
        RECT 20.448 51.824 20.592 52.016 ; 
        RECT 23.508 51.824 23.58 52.016 ; 
        RECT 37.764 51.824 37.836 52.016 ; 
        RECT 0.612 56.144 0.684 56.336 ; 
        RECT 14.868 56.144 14.94 56.336 ; 
        RECT 19.836 56.144 19.944 56.336 ; 
        RECT 20.448 56.144 20.592 56.336 ; 
        RECT 23.508 56.144 23.58 56.336 ; 
        RECT 37.764 56.144 37.836 56.336 ; 
        RECT 0.612 60.464 0.684 60.656 ; 
        RECT 14.868 60.464 14.94 60.656 ; 
        RECT 19.836 60.464 19.944 60.656 ; 
        RECT 20.448 60.464 20.592 60.656 ; 
        RECT 23.508 60.464 23.58 60.656 ; 
        RECT 37.764 60.464 37.836 60.656 ; 
        RECT 0.612 64.784 0.684 64.976 ; 
        RECT 14.868 64.784 14.94 64.976 ; 
        RECT 19.836 64.784 19.944 64.976 ; 
        RECT 20.448 64.784 20.592 64.976 ; 
        RECT 23.508 64.784 23.58 64.976 ; 
        RECT 37.764 64.784 37.836 64.976 ; 
        RECT 0.612 69.104 0.684 69.296 ; 
        RECT 14.868 69.104 14.94 69.296 ; 
        RECT 19.836 69.104 19.944 69.296 ; 
        RECT 20.448 69.104 20.592 69.296 ; 
        RECT 23.508 69.104 23.58 69.296 ; 
        RECT 37.764 69.104 37.836 69.296 ; 
        RECT 0.612 73.424 0.684 73.616 ; 
        RECT 14.868 73.424 14.94 73.616 ; 
        RECT 19.836 73.424 19.944 73.616 ; 
        RECT 20.448 73.424 20.592 73.616 ; 
        RECT 23.508 73.424 23.58 73.616 ; 
        RECT 37.764 73.424 37.836 73.616 ; 
        RECT 0.612 77.484 0.684 78.348 ; 
        RECT 19.708 102.828 19.78 103.692 ; 
        RECT 19.708 90.156 19.78 91.02 ; 
        RECT 19.708 77.484 19.78 78.348 ; 
        RECT 19.916 102.828 19.988 103.692 ; 
        RECT 19.916 90.156 19.988 91.02 ; 
        RECT 19.916 77.484 19.988 78.348 ; 
        RECT 20.124 102.828 20.196 103.692 ; 
        RECT 20.124 90.156 20.196 91.02 ; 
        RECT 20.124 77.484 20.196 78.348 ; 
        RECT 20.332 102.828 20.404 103.692 ; 
        RECT 20.332 90.156 20.404 91.02 ; 
        RECT 20.332 77.484 20.404 78.348 ; 
        RECT 20.54 102.828 20.612 103.692 ; 
        RECT 20.54 90.156 20.612 91.02 ; 
        RECT 20.54 77.484 20.612 78.348 ; 
        RECT 0.612 110.252 0.684 110.444 ; 
        RECT 14.868 110.252 14.94 110.444 ; 
        RECT 19.836 110.252 19.944 110.444 ; 
        RECT 20.448 110.252 20.592 110.444 ; 
        RECT 23.508 110.252 23.58 110.444 ; 
        RECT 37.764 110.252 37.836 110.444 ; 
        RECT 0.612 114.572 0.684 114.764 ; 
        RECT 14.868 114.572 14.94 114.764 ; 
        RECT 19.836 114.572 19.944 114.764 ; 
        RECT 20.448 114.572 20.592 114.764 ; 
        RECT 23.508 114.572 23.58 114.764 ; 
        RECT 37.764 114.572 37.836 114.764 ; 
        RECT 0.612 118.892 0.684 119.084 ; 
        RECT 14.868 118.892 14.94 119.084 ; 
        RECT 19.836 118.892 19.944 119.084 ; 
        RECT 20.448 118.892 20.592 119.084 ; 
        RECT 23.508 118.892 23.58 119.084 ; 
        RECT 37.764 118.892 37.836 119.084 ; 
        RECT 0.612 123.212 0.684 123.404 ; 
        RECT 14.868 123.212 14.94 123.404 ; 
        RECT 19.836 123.212 19.944 123.404 ; 
        RECT 20.448 123.212 20.592 123.404 ; 
        RECT 23.508 123.212 23.58 123.404 ; 
        RECT 37.764 123.212 37.836 123.404 ; 
        RECT 0.612 127.532 0.684 127.724 ; 
        RECT 14.868 127.532 14.94 127.724 ; 
        RECT 19.836 127.532 19.944 127.724 ; 
        RECT 20.448 127.532 20.592 127.724 ; 
        RECT 23.508 127.532 23.58 127.724 ; 
        RECT 37.764 127.532 37.836 127.724 ; 
        RECT 0.612 131.852 0.684 132.044 ; 
        RECT 14.868 131.852 14.94 132.044 ; 
        RECT 19.836 131.852 19.944 132.044 ; 
        RECT 20.448 131.852 20.592 132.044 ; 
        RECT 23.508 131.852 23.58 132.044 ; 
        RECT 37.764 131.852 37.836 132.044 ; 
        RECT 0.612 136.172 0.684 136.364 ; 
        RECT 14.868 136.172 14.94 136.364 ; 
        RECT 19.836 136.172 19.944 136.364 ; 
        RECT 20.448 136.172 20.592 136.364 ; 
        RECT 23.508 136.172 23.58 136.364 ; 
        RECT 37.764 136.172 37.836 136.364 ; 
        RECT 0.612 140.492 0.684 140.684 ; 
        RECT 14.868 140.492 14.94 140.684 ; 
        RECT 19.836 140.492 19.944 140.684 ; 
        RECT 20.448 140.492 20.592 140.684 ; 
        RECT 23.508 140.492 23.58 140.684 ; 
        RECT 37.764 140.492 37.836 140.684 ; 
        RECT 0.612 144.812 0.684 145.004 ; 
        RECT 14.868 144.812 14.94 145.004 ; 
        RECT 19.836 144.812 19.944 145.004 ; 
        RECT 20.448 144.812 20.592 145.004 ; 
        RECT 23.508 144.812 23.58 145.004 ; 
        RECT 37.764 144.812 37.836 145.004 ; 
        RECT 0.612 149.132 0.684 149.324 ; 
        RECT 14.868 149.132 14.94 149.324 ; 
        RECT 19.836 149.132 19.944 149.324 ; 
        RECT 20.448 149.132 20.592 149.324 ; 
        RECT 23.508 149.132 23.58 149.324 ; 
        RECT 37.764 149.132 37.836 149.324 ; 
        RECT 0.612 153.452 0.684 153.644 ; 
        RECT 14.868 153.452 14.94 153.644 ; 
        RECT 19.836 153.452 19.944 153.644 ; 
        RECT 20.448 153.452 20.592 153.644 ; 
        RECT 23.508 153.452 23.58 153.644 ; 
        RECT 37.764 153.452 37.836 153.644 ; 
        RECT 0.612 157.772 0.684 157.964 ; 
        RECT 14.868 157.772 14.94 157.964 ; 
        RECT 19.836 157.772 19.944 157.964 ; 
        RECT 20.448 157.772 20.592 157.964 ; 
        RECT 23.508 157.772 23.58 157.964 ; 
        RECT 37.764 157.772 37.836 157.964 ; 
        RECT 0.612 162.092 0.684 162.284 ; 
        RECT 14.868 162.092 14.94 162.284 ; 
        RECT 19.836 162.092 19.944 162.284 ; 
        RECT 20.448 162.092 20.592 162.284 ; 
        RECT 23.508 162.092 23.58 162.284 ; 
        RECT 37.764 162.092 37.836 162.284 ; 
        RECT 0.612 166.412 0.684 166.604 ; 
        RECT 14.868 166.412 14.94 166.604 ; 
        RECT 19.836 166.412 19.944 166.604 ; 
        RECT 20.448 166.412 20.592 166.604 ; 
        RECT 23.508 166.412 23.58 166.604 ; 
        RECT 37.764 166.412 37.836 166.604 ; 
        RECT 0.612 170.732 0.684 170.924 ; 
        RECT 14.868 170.732 14.94 170.924 ; 
        RECT 19.836 170.732 19.944 170.924 ; 
        RECT 20.448 170.732 20.592 170.924 ; 
        RECT 23.508 170.732 23.58 170.924 ; 
        RECT 37.764 170.732 37.836 170.924 ; 
        RECT 0.612 175.052 0.684 175.244 ; 
        RECT 14.868 175.052 14.94 175.244 ; 
        RECT 19.836 175.052 19.944 175.244 ; 
        RECT 20.448 175.052 20.592 175.244 ; 
        RECT 23.508 175.052 23.58 175.244 ; 
        RECT 37.764 175.052 37.836 175.244 ; 
        RECT 0.612 179.372 0.684 179.564 ; 
        RECT 14.868 179.372 14.94 179.564 ; 
        RECT 19.836 179.372 19.944 179.564 ; 
        RECT 20.448 179.372 20.592 179.564 ; 
        RECT 23.508 179.372 23.58 179.564 ; 
        RECT 37.764 179.372 37.836 179.564 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 29.34 79.372 29.412 79.52 ; 
      LAYER M4 ; 
        RECT 29.132 79.404 29.468 79.5 ; 
      LAYER M5 ; 
        RECT 29.328 75.6 29.424 88.56 ; 
      LAYER V3 ; 
        RECT 29.34 79.404 29.412 79.5 ; 
      LAYER V4 ; 
        RECT 29.328 79.404 29.424 79.5 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 28.476 79.384 28.548 79.532 ; 
      LAYER M4 ; 
        RECT 28.268 79.404 28.604 79.5 ; 
      LAYER M5 ; 
        RECT 28.464 75.6 28.56 88.56 ; 
      LAYER V3 ; 
        RECT 28.476 79.404 28.548 79.5 ; 
      LAYER V4 ; 
        RECT 28.464 79.404 28.56 79.5 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 27.612 77.068 27.684 77.216 ; 
      LAYER M4 ; 
        RECT 27.404 77.1 27.74 77.196 ; 
      LAYER M5 ; 
        RECT 27.6 75.6 27.696 88.56 ; 
      LAYER V3 ; 
        RECT 27.612 77.1 27.684 77.196 ; 
      LAYER V4 ; 
        RECT 27.6 77.1 27.696 77.196 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 26.748 78.028 26.82 78.752 ; 
      LAYER M4 ; 
        RECT 26.54 78.636 26.876 78.732 ; 
      LAYER M5 ; 
        RECT 26.736 75.6 26.832 88.56 ; 
      LAYER V3 ; 
        RECT 26.748 78.636 26.82 78.732 ; 
      LAYER V4 ; 
        RECT 26.736 78.636 26.832 78.732 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.884 77.08 25.956 77.348 ; 
      LAYER M4 ; 
        RECT 25.676 77.1 26.012 77.196 ; 
      LAYER M5 ; 
        RECT 25.872 75.6 25.968 88.56 ; 
      LAYER V3 ; 
        RECT 25.884 77.1 25.956 77.196 ; 
      LAYER V4 ; 
        RECT 25.872 77.1 25.968 77.196 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 25.02 76.012 25.092 77.024 ; 
      LAYER M4 ; 
        RECT 24.812 76.908 25.148 77.004 ; 
      LAYER M5 ; 
        RECT 25.008 75.6 25.104 88.56 ; 
      LAYER V3 ; 
        RECT 25.02 76.908 25.092 77.004 ; 
      LAYER V4 ; 
        RECT 25.008 76.908 25.104 77.004 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 24.156 80.152 24.228 80.3 ; 
      LAYER M4 ; 
        RECT 23.948 80.172 24.284 80.268 ; 
      LAYER M5 ; 
        RECT 24.144 75.6 24.24 88.56 ; 
      LAYER V3 ; 
        RECT 24.156 80.172 24.228 80.268 ; 
      LAYER V4 ; 
        RECT 24.144 80.172 24.24 80.268 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 20.7 77.08 20.772 77.348 ; 
      LAYER M4 ; 
        RECT 19.564 77.1 20.816 77.196 ; 
      LAYER M5 ; 
        RECT 19.608 75.6 19.704 88.56 ; 
      LAYER V3 ; 
        RECT 20.7 77.1 20.772 77.196 ; 
      LAYER V4 ; 
        RECT 19.608 77.1 19.704 77.196 ; 
    END 
  END ADDRESS[7] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 19.116 76.012 19.188 77.024 ; 
      LAYER M4 ; 
        RECT 18.268 76.908 19.232 77.004 ; 
      LAYER M5 ; 
        RECT 18.312 75.6 18.408 88.56 ; 
      LAYER V3 ; 
        RECT 19.116 76.908 19.188 77.004 ; 
      LAYER V4 ; 
        RECT 18.312 76.908 18.408 77.004 ; 
    END 
  END banksel 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.948 77.08 16.02 77.348 ; 
      LAYER M4 ; 
        RECT 15.74 77.1 16.076 77.196 ; 
      LAYER M5 ; 
        RECT 15.936 75.6 16.032 88.56 ; 
      LAYER V3 ; 
        RECT 15.948 77.1 16.02 77.196 ; 
      LAYER V4 ; 
        RECT 15.936 77.1 16.032 77.196 ; 
    END 
  END write 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.084 80.536 15.156 80.732 ; 
      LAYER M4 ; 
        RECT 14.876 80.556 15.212 80.652 ; 
      LAYER M5 ; 
        RECT 15.072 75.6 15.168 88.56 ; 
      LAYER V3 ; 
        RECT 15.084 80.556 15.156 80.652 ; 
      LAYER V4 ; 
        RECT 15.072 80.556 15.168 80.652 ; 
    END 
  END clk 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 15.228 76.012 15.3 77.024 ; 
      LAYER M4 ; 
        RECT 14.164 76.908 15.344 77.004 ; 
      LAYER M5 ; 
        RECT 14.208 75.6 14.304 88.56 ; 
      LAYER V3 ; 
        RECT 15.228 76.908 15.3 77.004 ; 
      LAYER V4 ; 
        RECT 14.208 76.908 14.304 77.004 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 13.356 79.372 13.428 79.52 ; 
      LAYER M4 ; 
        RECT 13.148 79.404 13.484 79.5 ; 
      LAYER M5 ; 
        RECT 13.344 75.6 13.44 88.56 ; 
      LAYER V3 ; 
        RECT 13.356 79.404 13.428 79.5 ; 
      LAYER V4 ; 
        RECT 13.344 79.404 13.44 79.5 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 12.492 77.08 12.564 77.996 ; 
      LAYER M4 ; 
        RECT 12.284 77.1 12.62 77.196 ; 
      LAYER M5 ; 
        RECT 12.48 75.6 12.576 88.56 ; 
      LAYER V3 ; 
        RECT 12.492 77.1 12.564 77.196 ; 
      LAYER V4 ; 
        RECT 12.48 77.1 12.576 77.196 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 11.628 76.012 11.7 77.024 ; 
      LAYER M4 ; 
        RECT 11.42 76.908 11.756 77.004 ; 
      LAYER M5 ; 
        RECT 11.616 75.6 11.712 88.56 ; 
      LAYER V3 ; 
        RECT 11.628 76.908 11.7 77.004 ; 
      LAYER V4 ; 
        RECT 11.616 76.908 11.712 77.004 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 10.764 77.068 10.836 77.216 ; 
      LAYER M4 ; 
        RECT 10.556 77.1 10.892 77.196 ; 
      LAYER M5 ; 
        RECT 10.752 75.6 10.848 88.56 ; 
      LAYER V3 ; 
        RECT 10.764 77.1 10.836 77.196 ; 
      LAYER V4 ; 
        RECT 10.752 77.1 10.848 77.196 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 9.9 79.372 9.972 79.52 ; 
      LAYER M4 ; 
        RECT 9.692 79.404 10.028 79.5 ; 
      LAYER M5 ; 
        RECT 9.888 75.6 9.984 88.56 ; 
      LAYER V3 ; 
        RECT 9.9 79.404 9.972 79.5 ; 
      LAYER V4 ; 
        RECT 9.888 79.404 9.984 79.5 ; 
    END 
  END sdel[4] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.712 20.544 1.808 ; 
      LAYER M3 ; 
        RECT 20.304 1.51 20.376 2.468 ; 
      LAYER V3 ; 
        RECT 20.304 1.712 20.376 1.808 ; 
    END 
  END dataout[0] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 1.328 20.816 1.424 ; 
      LAYER M3 ; 
        RECT 19.404 1.08 19.476 2.7 ; 
      LAYER V3 ; 
        RECT 19.404 1.328 19.476 1.424 ; 
    END 
  END wd[0] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 6.032 20.544 6.128 ; 
      LAYER M3 ; 
        RECT 20.304 5.83 20.376 6.788 ; 
      LAYER V3 ; 
        RECT 20.304 6.032 20.376 6.128 ; 
    END 
  END dataout[1] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 5.648 20.816 5.744 ; 
      LAYER M3 ; 
        RECT 19.404 5.4 19.476 7.02 ; 
      LAYER V3 ; 
        RECT 19.404 5.648 19.476 5.744 ; 
    END 
  END wd[1] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 10.352 20.544 10.448 ; 
      LAYER M3 ; 
        RECT 20.304 10.15 20.376 11.108 ; 
      LAYER V3 ; 
        RECT 20.304 10.352 20.376 10.448 ; 
    END 
  END dataout[2] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 9.968 20.816 10.064 ; 
      LAYER M3 ; 
        RECT 19.404 9.72 19.476 11.34 ; 
      LAYER V3 ; 
        RECT 19.404 9.968 19.476 10.064 ; 
    END 
  END wd[2] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.672 20.544 14.768 ; 
      LAYER M3 ; 
        RECT 20.304 14.47 20.376 15.428 ; 
      LAYER V3 ; 
        RECT 20.304 14.672 20.376 14.768 ; 
    END 
  END dataout[3] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 14.288 20.816 14.384 ; 
      LAYER M3 ; 
        RECT 19.404 14.04 19.476 15.66 ; 
      LAYER V3 ; 
        RECT 19.404 14.288 19.476 14.384 ; 
    END 
  END wd[3] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.992 20.544 19.088 ; 
      LAYER M3 ; 
        RECT 20.304 18.79 20.376 19.748 ; 
      LAYER V3 ; 
        RECT 20.304 18.992 20.376 19.088 ; 
    END 
  END dataout[4] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 18.608 20.816 18.704 ; 
      LAYER M3 ; 
        RECT 19.404 18.36 19.476 19.98 ; 
      LAYER V3 ; 
        RECT 19.404 18.608 19.476 18.704 ; 
    END 
  END wd[4] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 23.312 20.544 23.408 ; 
      LAYER M3 ; 
        RECT 20.304 23.11 20.376 24.068 ; 
      LAYER V3 ; 
        RECT 20.304 23.312 20.376 23.408 ; 
    END 
  END dataout[5] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 22.928 20.816 23.024 ; 
      LAYER M3 ; 
        RECT 19.404 22.68 19.476 24.3 ; 
      LAYER V3 ; 
        RECT 19.404 22.928 19.476 23.024 ; 
    END 
  END wd[5] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.632 20.544 27.728 ; 
      LAYER M3 ; 
        RECT 20.304 27.43 20.376 28.388 ; 
      LAYER V3 ; 
        RECT 20.304 27.632 20.376 27.728 ; 
    END 
  END dataout[6] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 27.248 20.816 27.344 ; 
      LAYER M3 ; 
        RECT 19.404 27 19.476 28.62 ; 
      LAYER V3 ; 
        RECT 19.404 27.248 19.476 27.344 ; 
    END 
  END wd[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.952 20.544 32.048 ; 
      LAYER M3 ; 
        RECT 20.304 31.75 20.376 32.708 ; 
      LAYER V3 ; 
        RECT 20.304 31.952 20.376 32.048 ; 
    END 
  END dataout[7] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 31.568 20.816 31.664 ; 
      LAYER M3 ; 
        RECT 19.404 31.32 19.476 32.94 ; 
      LAYER V3 ; 
        RECT 19.404 31.568 19.476 31.664 ; 
    END 
  END wd[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 36.272 20.544 36.368 ; 
      LAYER M3 ; 
        RECT 20.304 36.07 20.376 37.028 ; 
      LAYER V3 ; 
        RECT 20.304 36.272 20.376 36.368 ; 
    END 
  END dataout[8] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 35.888 20.816 35.984 ; 
      LAYER M3 ; 
        RECT 19.404 35.64 19.476 37.26 ; 
      LAYER V3 ; 
        RECT 19.404 35.888 19.476 35.984 ; 
    END 
  END wd[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 40.592 20.544 40.688 ; 
      LAYER M3 ; 
        RECT 20.304 40.39 20.376 41.348 ; 
      LAYER V3 ; 
        RECT 20.304 40.592 20.376 40.688 ; 
    END 
  END dataout[9] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 40.208 20.816 40.304 ; 
      LAYER M3 ; 
        RECT 19.404 39.96 19.476 41.58 ; 
      LAYER V3 ; 
        RECT 19.404 40.208 19.476 40.304 ; 
    END 
  END wd[9] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 44.912 20.544 45.008 ; 
      LAYER M3 ; 
        RECT 20.304 44.71 20.376 45.668 ; 
      LAYER V3 ; 
        RECT 20.304 44.912 20.376 45.008 ; 
    END 
  END dataout[10] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 44.528 20.816 44.624 ; 
      LAYER M3 ; 
        RECT 19.404 44.28 19.476 45.9 ; 
      LAYER V3 ; 
        RECT 19.404 44.528 19.476 44.624 ; 
    END 
  END wd[10] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 49.232 20.544 49.328 ; 
      LAYER M3 ; 
        RECT 20.304 49.03 20.376 49.988 ; 
      LAYER V3 ; 
        RECT 20.304 49.232 20.376 49.328 ; 
    END 
  END dataout[11] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 48.848 20.816 48.944 ; 
      LAYER M3 ; 
        RECT 19.404 48.6 19.476 50.22 ; 
      LAYER V3 ; 
        RECT 19.404 48.848 19.476 48.944 ; 
    END 
  END wd[11] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 53.552 20.544 53.648 ; 
      LAYER M3 ; 
        RECT 20.304 53.35 20.376 54.308 ; 
      LAYER V3 ; 
        RECT 20.304 53.552 20.376 53.648 ; 
    END 
  END dataout[12] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 53.168 20.816 53.264 ; 
      LAYER M3 ; 
        RECT 19.404 52.92 19.476 54.54 ; 
      LAYER V3 ; 
        RECT 19.404 53.168 19.476 53.264 ; 
    END 
  END wd[12] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 57.872 20.544 57.968 ; 
      LAYER M3 ; 
        RECT 20.304 57.67 20.376 58.628 ; 
      LAYER V3 ; 
        RECT 20.304 57.872 20.376 57.968 ; 
    END 
  END dataout[13] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 57.488 20.816 57.584 ; 
      LAYER M3 ; 
        RECT 19.404 57.24 19.476 58.86 ; 
      LAYER V3 ; 
        RECT 19.404 57.488 19.476 57.584 ; 
    END 
  END wd[13] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 62.192 20.544 62.288 ; 
      LAYER M3 ; 
        RECT 20.304 61.99 20.376 62.948 ; 
      LAYER V3 ; 
        RECT 20.304 62.192 20.376 62.288 ; 
    END 
  END dataout[14] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 61.808 20.816 61.904 ; 
      LAYER M3 ; 
        RECT 19.404 61.56 19.476 63.18 ; 
      LAYER V3 ; 
        RECT 19.404 61.808 19.476 61.904 ; 
    END 
  END wd[14] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 66.512 20.544 66.608 ; 
      LAYER M3 ; 
        RECT 20.304 66.31 20.376 67.268 ; 
      LAYER V3 ; 
        RECT 20.304 66.512 20.376 66.608 ; 
    END 
  END dataout[15] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 66.128 20.816 66.224 ; 
      LAYER M3 ; 
        RECT 19.404 65.88 19.476 67.5 ; 
      LAYER V3 ; 
        RECT 19.404 66.128 19.476 66.224 ; 
    END 
  END wd[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 70.832 20.544 70.928 ; 
      LAYER M3 ; 
        RECT 20.304 70.63 20.376 71.588 ; 
      LAYER V3 ; 
        RECT 20.304 70.832 20.376 70.928 ; 
    END 
  END dataout[16] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 70.448 20.816 70.544 ; 
      LAYER M3 ; 
        RECT 19.404 70.2 19.476 71.82 ; 
      LAYER V3 ; 
        RECT 19.404 70.448 19.476 70.544 ; 
    END 
  END wd[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 107.66 20.544 107.756 ; 
      LAYER M3 ; 
        RECT 20.304 107.458 20.376 108.416 ; 
      LAYER V3 ; 
        RECT 20.304 107.66 20.376 107.756 ; 
    END 
  END dataout[17] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 107.276 20.816 107.372 ; 
      LAYER M3 ; 
        RECT 19.404 107.028 19.476 108.648 ; 
      LAYER V3 ; 
        RECT 19.404 107.276 19.476 107.372 ; 
    END 
  END wd[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 111.98 20.544 112.076 ; 
      LAYER M3 ; 
        RECT 20.304 111.778 20.376 112.736 ; 
      LAYER V3 ; 
        RECT 20.304 111.98 20.376 112.076 ; 
    END 
  END dataout[18] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 111.596 20.816 111.692 ; 
      LAYER M3 ; 
        RECT 19.404 111.348 19.476 112.968 ; 
      LAYER V3 ; 
        RECT 19.404 111.596 19.476 111.692 ; 
    END 
  END wd[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 116.3 20.544 116.396 ; 
      LAYER M3 ; 
        RECT 20.304 116.098 20.376 117.056 ; 
      LAYER V3 ; 
        RECT 20.304 116.3 20.376 116.396 ; 
    END 
  END dataout[19] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 115.916 20.816 116.012 ; 
      LAYER M3 ; 
        RECT 19.404 115.668 19.476 117.288 ; 
      LAYER V3 ; 
        RECT 19.404 115.916 19.476 116.012 ; 
    END 
  END wd[19] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 120.62 20.544 120.716 ; 
      LAYER M3 ; 
        RECT 20.304 120.418 20.376 121.376 ; 
      LAYER V3 ; 
        RECT 20.304 120.62 20.376 120.716 ; 
    END 
  END dataout[20] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 120.236 20.816 120.332 ; 
      LAYER M3 ; 
        RECT 19.404 119.988 19.476 121.608 ; 
      LAYER V3 ; 
        RECT 19.404 120.236 19.476 120.332 ; 
    END 
  END wd[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 124.94 20.544 125.036 ; 
      LAYER M3 ; 
        RECT 20.304 124.738 20.376 125.696 ; 
      LAYER V3 ; 
        RECT 20.304 124.94 20.376 125.036 ; 
    END 
  END dataout[21] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 124.556 20.816 124.652 ; 
      LAYER M3 ; 
        RECT 19.404 124.308 19.476 125.928 ; 
      LAYER V3 ; 
        RECT 19.404 124.556 19.476 124.652 ; 
    END 
  END wd[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 129.26 20.544 129.356 ; 
      LAYER M3 ; 
        RECT 20.304 129.058 20.376 130.016 ; 
      LAYER V3 ; 
        RECT 20.304 129.26 20.376 129.356 ; 
    END 
  END dataout[22] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 128.876 20.816 128.972 ; 
      LAYER M3 ; 
        RECT 19.404 128.628 19.476 130.248 ; 
      LAYER V3 ; 
        RECT 19.404 128.876 19.476 128.972 ; 
    END 
  END wd[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 133.58 20.544 133.676 ; 
      LAYER M3 ; 
        RECT 20.304 133.378 20.376 134.336 ; 
      LAYER V3 ; 
        RECT 20.304 133.58 20.376 133.676 ; 
    END 
  END dataout[23] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 133.196 20.816 133.292 ; 
      LAYER M3 ; 
        RECT 19.404 132.948 19.476 134.568 ; 
      LAYER V3 ; 
        RECT 19.404 133.196 19.476 133.292 ; 
    END 
  END wd[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 137.9 20.544 137.996 ; 
      LAYER M3 ; 
        RECT 20.304 137.698 20.376 138.656 ; 
      LAYER V3 ; 
        RECT 20.304 137.9 20.376 137.996 ; 
    END 
  END dataout[24] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 137.516 20.816 137.612 ; 
      LAYER M3 ; 
        RECT 19.404 137.268 19.476 138.888 ; 
      LAYER V3 ; 
        RECT 19.404 137.516 19.476 137.612 ; 
    END 
  END wd[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 142.22 20.544 142.316 ; 
      LAYER M3 ; 
        RECT 20.304 142.018 20.376 142.976 ; 
      LAYER V3 ; 
        RECT 20.304 142.22 20.376 142.316 ; 
    END 
  END dataout[25] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 141.836 20.816 141.932 ; 
      LAYER M3 ; 
        RECT 19.404 141.588 19.476 143.208 ; 
      LAYER V3 ; 
        RECT 19.404 141.836 19.476 141.932 ; 
    END 
  END wd[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 146.54 20.544 146.636 ; 
      LAYER M3 ; 
        RECT 20.304 146.338 20.376 147.296 ; 
      LAYER V3 ; 
        RECT 20.304 146.54 20.376 146.636 ; 
    END 
  END dataout[26] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 146.156 20.816 146.252 ; 
      LAYER M3 ; 
        RECT 19.404 145.908 19.476 147.528 ; 
      LAYER V3 ; 
        RECT 19.404 146.156 19.476 146.252 ; 
    END 
  END wd[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 150.86 20.544 150.956 ; 
      LAYER M3 ; 
        RECT 20.304 150.658 20.376 151.616 ; 
      LAYER V3 ; 
        RECT 20.304 150.86 20.376 150.956 ; 
    END 
  END dataout[27] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 150.476 20.816 150.572 ; 
      LAYER M3 ; 
        RECT 19.404 150.228 19.476 151.848 ; 
      LAYER V3 ; 
        RECT 19.404 150.476 19.476 150.572 ; 
    END 
  END wd[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 155.18 20.544 155.276 ; 
      LAYER M3 ; 
        RECT 20.304 154.978 20.376 155.936 ; 
      LAYER V3 ; 
        RECT 20.304 155.18 20.376 155.276 ; 
    END 
  END dataout[28] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 154.796 20.816 154.892 ; 
      LAYER M3 ; 
        RECT 19.404 154.548 19.476 156.168 ; 
      LAYER V3 ; 
        RECT 19.404 154.796 19.476 154.892 ; 
    END 
  END wd[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 159.5 20.544 159.596 ; 
      LAYER M3 ; 
        RECT 20.304 159.298 20.376 160.256 ; 
      LAYER V3 ; 
        RECT 20.304 159.5 20.376 159.596 ; 
    END 
  END dataout[29] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 159.116 20.816 159.212 ; 
      LAYER M3 ; 
        RECT 19.404 158.868 19.476 160.488 ; 
      LAYER V3 ; 
        RECT 19.404 159.116 19.476 159.212 ; 
    END 
  END wd[29] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 163.82 20.544 163.916 ; 
      LAYER M3 ; 
        RECT 20.304 163.618 20.376 164.576 ; 
      LAYER V3 ; 
        RECT 20.304 163.82 20.376 163.916 ; 
    END 
  END dataout[30] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 163.436 20.816 163.532 ; 
      LAYER M3 ; 
        RECT 19.404 163.188 19.476 164.808 ; 
      LAYER V3 ; 
        RECT 19.404 163.436 19.476 163.532 ; 
    END 
  END wd[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 168.14 20.544 168.236 ; 
      LAYER M3 ; 
        RECT 20.304 167.938 20.376 168.896 ; 
      LAYER V3 ; 
        RECT 20.304 168.14 20.376 168.236 ; 
    END 
  END dataout[31] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 167.756 20.816 167.852 ; 
      LAYER M3 ; 
        RECT 19.404 167.508 19.476 169.128 ; 
      LAYER V3 ; 
        RECT 19.404 167.756 19.476 167.852 ; 
    END 
  END wd[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 172.46 20.544 172.556 ; 
      LAYER M3 ; 
        RECT 20.304 172.258 20.376 173.216 ; 
      LAYER V3 ; 
        RECT 20.304 172.46 20.376 172.556 ; 
    END 
  END dataout[32] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 172.076 20.816 172.172 ; 
      LAYER M3 ; 
        RECT 19.404 171.828 19.476 173.448 ; 
      LAYER V3 ; 
        RECT 19.404 172.076 19.476 172.172 ; 
    END 
  END wd[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 176.78 20.544 176.876 ; 
      LAYER M3 ; 
        RECT 20.304 176.578 20.376 177.536 ; 
      LAYER V3 ; 
        RECT 20.304 176.78 20.376 176.876 ; 
    END 
  END dataout[33] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M4 ; 
        RECT 17.952 176.396 20.816 176.492 ; 
      LAYER M3 ; 
        RECT 19.404 176.148 19.476 177.768 ; 
      LAYER V3 ; 
        RECT 19.404 176.396 19.476 176.492 ; 
    END 
  END wd[33] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.412 38.448 109.026 ; 
        RECT 0 106.974 38.448 111.348 ; 
        RECT 0 111.294 38.448 115.668 ; 
        RECT 0 115.614 38.448 119.988 ; 
        RECT 0 119.934 38.448 124.308 ; 
        RECT 0 124.254 38.448 128.628 ; 
        RECT 0 128.574 38.448 132.948 ; 
        RECT 0 132.894 38.448 137.268 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.412 38.448 109.026 ; 
        RECT 0 106.974 38.448 111.348 ; 
        RECT 0 111.294 38.448 115.668 ; 
        RECT 0 115.614 38.448 119.988 ; 
        RECT 0 119.934 38.448 124.308 ; 
        RECT 0 124.254 38.448 128.628 ; 
        RECT 0 128.574 38.448 132.948 ; 
        RECT 0 132.894 38.448 137.268 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
  LAYER V1 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.412 38.448 109.026 ; 
        RECT 0 106.974 38.448 111.348 ; 
        RECT 0 111.294 38.448 115.668 ; 
        RECT 0 115.614 38.448 119.988 ; 
        RECT 0 119.934 38.448 124.308 ; 
        RECT 0 124.254 38.448 128.628 ; 
        RECT 0 128.574 38.448 132.948 ; 
        RECT 0 132.894 38.448 137.268 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
  LAYER V2 ; 
      RECT 0 1.026 38.448 5.4 ; 
      RECT 0 5.346 38.448 9.72 ; 
      RECT 0 9.666 38.448 14.04 ; 
      RECT 0 13.986 38.448 18.36 ; 
      RECT 0 18.306 38.448 22.68 ; 
      RECT 0 22.626 38.448 27 ; 
      RECT 0 26.946 38.448 31.32 ; 
      RECT 0 31.266 38.448 35.64 ; 
      RECT 0 35.586 38.448 39.96 ; 
      RECT 0 39.906 38.448 44.28 ; 
      RECT 0 44.226 38.448 48.6 ; 
      RECT 0 48.546 38.448 52.92 ; 
      RECT 0 52.866 38.448 57.24 ; 
      RECT 0 57.186 38.448 61.56 ; 
      RECT 0 61.506 38.448 65.88 ; 
      RECT 0 65.826 38.448 70.2 ; 
      RECT 0 70.146 38.448 74.52 ; 
      RECT 0 74.412 38.448 109.026 ; 
        RECT 0 106.974 38.448 111.348 ; 
        RECT 0 111.294 38.448 115.668 ; 
        RECT 0 115.614 38.448 119.988 ; 
        RECT 0 119.934 38.448 124.308 ; 
        RECT 0 124.254 38.448 128.628 ; 
        RECT 0 128.574 38.448 132.948 ; 
        RECT 0 132.894 38.448 137.268 ; 
        RECT 0 137.214 38.448 141.588 ; 
        RECT 0 141.534 38.448 145.908 ; 
        RECT 0 145.854 38.448 150.228 ; 
        RECT 0 150.174 38.448 154.548 ; 
        RECT 0 154.494 38.448 158.868 ; 
        RECT 0 158.814 38.448 163.188 ; 
        RECT 0 163.134 38.448 167.508 ; 
        RECT 0 167.454 38.448 171.828 ; 
        RECT 0 171.774 38.448 176.148 ; 
        RECT 0 176.094 38.448 180.468 ; 
  LAYER M3 ; 
      RECT 20.952 1.38 21.024 5.122 ; 
      RECT 20.808 1.38 20.88 5.122 ; 
      RECT 20.664 3.688 20.736 4.978 ; 
      RECT 20.196 4.476 20.268 4.914 ; 
      RECT 20.16 1.51 20.232 2.468 ; 
      RECT 20.016 3.834 20.088 4.448 ; 
      RECT 19.692 3.936 19.764 4.968 ; 
      RECT 17.532 1.38 17.604 5.122 ; 
      RECT 17.388 1.38 17.46 5.122 ; 
      RECT 17.244 2.104 17.316 4.376 ; 
      RECT 20.952 5.7 21.024 9.442 ; 
      RECT 20.808 5.7 20.88 9.442 ; 
      RECT 20.664 8.008 20.736 9.298 ; 
      RECT 20.196 8.796 20.268 9.234 ; 
      RECT 20.16 5.83 20.232 6.788 ; 
      RECT 20.016 8.154 20.088 8.768 ; 
      RECT 19.692 8.256 19.764 9.288 ; 
      RECT 17.532 5.7 17.604 9.442 ; 
      RECT 17.388 5.7 17.46 9.442 ; 
      RECT 17.244 6.424 17.316 8.696 ; 
      RECT 20.952 10.02 21.024 13.762 ; 
      RECT 20.808 10.02 20.88 13.762 ; 
      RECT 20.664 12.328 20.736 13.618 ; 
      RECT 20.196 13.116 20.268 13.554 ; 
      RECT 20.16 10.15 20.232 11.108 ; 
      RECT 20.016 12.474 20.088 13.088 ; 
      RECT 19.692 12.576 19.764 13.608 ; 
      RECT 17.532 10.02 17.604 13.762 ; 
      RECT 17.388 10.02 17.46 13.762 ; 
      RECT 17.244 10.744 17.316 13.016 ; 
      RECT 20.952 14.34 21.024 18.082 ; 
      RECT 20.808 14.34 20.88 18.082 ; 
      RECT 20.664 16.648 20.736 17.938 ; 
      RECT 20.196 17.436 20.268 17.874 ; 
      RECT 20.16 14.47 20.232 15.428 ; 
      RECT 20.016 16.794 20.088 17.408 ; 
      RECT 19.692 16.896 19.764 17.928 ; 
      RECT 17.532 14.34 17.604 18.082 ; 
      RECT 17.388 14.34 17.46 18.082 ; 
      RECT 17.244 15.064 17.316 17.336 ; 
      RECT 20.952 18.66 21.024 22.402 ; 
      RECT 20.808 18.66 20.88 22.402 ; 
      RECT 20.664 20.968 20.736 22.258 ; 
      RECT 20.196 21.756 20.268 22.194 ; 
      RECT 20.16 18.79 20.232 19.748 ; 
      RECT 20.016 21.114 20.088 21.728 ; 
      RECT 19.692 21.216 19.764 22.248 ; 
      RECT 17.532 18.66 17.604 22.402 ; 
      RECT 17.388 18.66 17.46 22.402 ; 
      RECT 17.244 19.384 17.316 21.656 ; 
      RECT 20.952 22.98 21.024 26.722 ; 
      RECT 20.808 22.98 20.88 26.722 ; 
      RECT 20.664 25.288 20.736 26.578 ; 
      RECT 20.196 26.076 20.268 26.514 ; 
      RECT 20.16 23.11 20.232 24.068 ; 
      RECT 20.016 25.434 20.088 26.048 ; 
      RECT 19.692 25.536 19.764 26.568 ; 
      RECT 17.532 22.98 17.604 26.722 ; 
      RECT 17.388 22.98 17.46 26.722 ; 
      RECT 17.244 23.704 17.316 25.976 ; 
      RECT 20.952 27.3 21.024 31.042 ; 
      RECT 20.808 27.3 20.88 31.042 ; 
      RECT 20.664 29.608 20.736 30.898 ; 
      RECT 20.196 30.396 20.268 30.834 ; 
      RECT 20.16 27.43 20.232 28.388 ; 
      RECT 20.016 29.754 20.088 30.368 ; 
      RECT 19.692 29.856 19.764 30.888 ; 
      RECT 17.532 27.3 17.604 31.042 ; 
      RECT 17.388 27.3 17.46 31.042 ; 
      RECT 17.244 28.024 17.316 30.296 ; 
      RECT 20.952 31.62 21.024 35.362 ; 
      RECT 20.808 31.62 20.88 35.362 ; 
      RECT 20.664 33.928 20.736 35.218 ; 
      RECT 20.196 34.716 20.268 35.154 ; 
      RECT 20.16 31.75 20.232 32.708 ; 
      RECT 20.016 34.074 20.088 34.688 ; 
      RECT 19.692 34.176 19.764 35.208 ; 
      RECT 17.532 31.62 17.604 35.362 ; 
      RECT 17.388 31.62 17.46 35.362 ; 
      RECT 17.244 32.344 17.316 34.616 ; 
      RECT 20.952 35.94 21.024 39.682 ; 
      RECT 20.808 35.94 20.88 39.682 ; 
      RECT 20.664 38.248 20.736 39.538 ; 
      RECT 20.196 39.036 20.268 39.474 ; 
      RECT 20.16 36.07 20.232 37.028 ; 
      RECT 20.016 38.394 20.088 39.008 ; 
      RECT 19.692 38.496 19.764 39.528 ; 
      RECT 17.532 35.94 17.604 39.682 ; 
      RECT 17.388 35.94 17.46 39.682 ; 
      RECT 17.244 36.664 17.316 38.936 ; 
      RECT 20.952 40.26 21.024 44.002 ; 
      RECT 20.808 40.26 20.88 44.002 ; 
      RECT 20.664 42.568 20.736 43.858 ; 
      RECT 20.196 43.356 20.268 43.794 ; 
      RECT 20.16 40.39 20.232 41.348 ; 
      RECT 20.016 42.714 20.088 43.328 ; 
      RECT 19.692 42.816 19.764 43.848 ; 
      RECT 17.532 40.26 17.604 44.002 ; 
      RECT 17.388 40.26 17.46 44.002 ; 
      RECT 17.244 40.984 17.316 43.256 ; 
      RECT 20.952 44.58 21.024 48.322 ; 
      RECT 20.808 44.58 20.88 48.322 ; 
      RECT 20.664 46.888 20.736 48.178 ; 
      RECT 20.196 47.676 20.268 48.114 ; 
      RECT 20.16 44.71 20.232 45.668 ; 
      RECT 20.016 47.034 20.088 47.648 ; 
      RECT 19.692 47.136 19.764 48.168 ; 
      RECT 17.532 44.58 17.604 48.322 ; 
      RECT 17.388 44.58 17.46 48.322 ; 
      RECT 17.244 45.304 17.316 47.576 ; 
      RECT 20.952 48.9 21.024 52.642 ; 
      RECT 20.808 48.9 20.88 52.642 ; 
      RECT 20.664 51.208 20.736 52.498 ; 
      RECT 20.196 51.996 20.268 52.434 ; 
      RECT 20.16 49.03 20.232 49.988 ; 
      RECT 20.016 51.354 20.088 51.968 ; 
      RECT 19.692 51.456 19.764 52.488 ; 
      RECT 17.532 48.9 17.604 52.642 ; 
      RECT 17.388 48.9 17.46 52.642 ; 
      RECT 17.244 49.624 17.316 51.896 ; 
      RECT 20.952 53.22 21.024 56.962 ; 
      RECT 20.808 53.22 20.88 56.962 ; 
      RECT 20.664 55.528 20.736 56.818 ; 
      RECT 20.196 56.316 20.268 56.754 ; 
      RECT 20.16 53.35 20.232 54.308 ; 
      RECT 20.016 55.674 20.088 56.288 ; 
      RECT 19.692 55.776 19.764 56.808 ; 
      RECT 17.532 53.22 17.604 56.962 ; 
      RECT 17.388 53.22 17.46 56.962 ; 
      RECT 17.244 53.944 17.316 56.216 ; 
      RECT 20.952 57.54 21.024 61.282 ; 
      RECT 20.808 57.54 20.88 61.282 ; 
      RECT 20.664 59.848 20.736 61.138 ; 
      RECT 20.196 60.636 20.268 61.074 ; 
      RECT 20.16 57.67 20.232 58.628 ; 
      RECT 20.016 59.994 20.088 60.608 ; 
      RECT 19.692 60.096 19.764 61.128 ; 
      RECT 17.532 57.54 17.604 61.282 ; 
      RECT 17.388 57.54 17.46 61.282 ; 
      RECT 17.244 58.264 17.316 60.536 ; 
      RECT 20.952 61.86 21.024 65.602 ; 
      RECT 20.808 61.86 20.88 65.602 ; 
      RECT 20.664 64.168 20.736 65.458 ; 
      RECT 20.196 64.956 20.268 65.394 ; 
      RECT 20.16 61.99 20.232 62.948 ; 
      RECT 20.016 64.314 20.088 64.928 ; 
      RECT 19.692 64.416 19.764 65.448 ; 
      RECT 17.532 61.86 17.604 65.602 ; 
      RECT 17.388 61.86 17.46 65.602 ; 
      RECT 17.244 62.584 17.316 64.856 ; 
      RECT 20.952 66.18 21.024 69.922 ; 
      RECT 20.808 66.18 20.88 69.922 ; 
      RECT 20.664 68.488 20.736 69.778 ; 
      RECT 20.196 69.276 20.268 69.714 ; 
      RECT 20.16 66.31 20.232 67.268 ; 
      RECT 20.016 68.634 20.088 69.248 ; 
      RECT 19.692 68.736 19.764 69.768 ; 
      RECT 17.532 66.18 17.604 69.922 ; 
      RECT 17.388 66.18 17.46 69.922 ; 
      RECT 17.244 66.904 17.316 69.176 ; 
      RECT 20.952 70.5 21.024 74.242 ; 
      RECT 20.808 70.5 20.88 74.242 ; 
      RECT 20.664 72.808 20.736 74.098 ; 
      RECT 20.196 73.596 20.268 74.034 ; 
      RECT 20.16 70.63 20.232 71.588 ; 
      RECT 20.016 72.954 20.088 73.568 ; 
      RECT 19.692 73.056 19.764 74.088 ; 
      RECT 17.532 70.5 17.604 74.242 ; 
      RECT 17.388 70.5 17.46 74.242 ; 
      RECT 17.244 71.224 17.316 73.496 ; 
      RECT 37.62 89.584 37.692 107.006 ; 
      RECT 37.476 84.324 37.548 84.6 ; 
      RECT 37.476 91.556 37.548 93.414 ; 
      RECT 37.332 74.306 37.404 107.134 ; 
      RECT 37.188 89.384 37.26 92.474 ; 
      RECT 37.188 92.6788 37.26 94.644 ; 
      RECT 37.188 94.844 37.26 96.33 ; 
      RECT 37.188 96.582 37.26 99.828 ; 
      RECT 37.044 89.726 37.116 92.294 ; 
      RECT 37.044 95.004 37.116 97.132 ; 
      RECT 36.9 74.306 36.972 75.706 ; 
      RECT 36.468 74.306 36.54 75.706 ; 
      RECT 36.036 74.306 36.108 75.706 ; 
      RECT 35.604 74.306 35.676 75.706 ; 
      RECT 35.172 74.306 35.244 75.706 ; 
      RECT 34.74 74.306 34.812 75.706 ; 
      RECT 34.308 74.306 34.38 75.706 ; 
      RECT 33.876 74.306 33.948 75.706 ; 
      RECT 33.444 74.306 33.516 75.706 ; 
      RECT 33.012 74.306 33.084 75.706 ; 
      RECT 32.58 74.306 32.652 75.706 ; 
      RECT 32.148 74.306 32.22 75.706 ; 
      RECT 31.716 74.306 31.788 75.706 ; 
      RECT 31.284 74.306 31.356 75.706 ; 
      RECT 30.852 74.306 30.924 75.706 ; 
      RECT 30.42 74.306 30.492 75.706 ; 
      RECT 29.988 74.306 30.06 75.706 ; 
      RECT 29.556 74.306 29.628 75.706 ; 
      RECT 29.124 74.306 29.196 75.706 ; 
      RECT 28.692 74.306 28.764 75.706 ; 
      RECT 28.26 74.306 28.332 75.706 ; 
      RECT 27.828 74.306 27.9 75.706 ; 
      RECT 27.396 74.306 27.468 75.706 ; 
      RECT 26.964 74.306 27.036 75.706 ; 
      RECT 26.532 74.306 26.604 75.706 ; 
      RECT 26.1 74.306 26.172 75.706 ; 
      RECT 25.668 74.306 25.74 75.706 ; 
      RECT 25.236 74.306 25.308 75.706 ; 
      RECT 24.804 74.306 24.876 75.706 ; 
      RECT 24.372 74.306 24.444 75.706 ; 
      RECT 24.228 89.46 24.3 92.2788 ; 
      RECT 24.228 95.248 24.3 99.972 ; 
      RECT 24.156 76.948 24.228 79.652 ; 
      RECT 24.156 82.636 24.228 83.828 ; 
      RECT 24.084 89.714 24.156 92.474 ; 
      RECT 24.084 92.678 24.156 96.644 ; 
      RECT 24.084 96.764 24.156 99.9 ; 
      RECT 23.94 74.306 24.012 107.134 ; 
      RECT 23.796 90.804 23.868 91.136 ; 
      RECT 23.724 77.38 23.796 79.904 ; 
      RECT 23.724 81.556 23.796 82.316 ; 
      RECT 23.724 85.084 23.796 85.28 ; 
      RECT 23.652 89.584 23.724 107.024 ; 
      RECT 23.292 75.868 23.364 79.076 ; 
      RECT 23.292 81.268 23.364 83.54 ; 
      RECT 23.148 81.556 23.22 83.036 ; 
      RECT 23.004 78.964 23.076 79.508 ; 
      RECT 23.004 82.924 23.076 83.828 ; 
      RECT 23.004 87.892 23.076 88.148 ; 
      RECT 22.86 79.372 22.932 79.52 ; 
      RECT 22.86 85.876 22.932 86.048 ; 
      RECT 22.86 88.012 22.932 88.16 ; 
      RECT 22.716 80.62 22.788 82.604 ; 
      RECT 22.716 82.78 22.788 83.54 ; 
      RECT 22.716 86.62 22.788 87.86 ; 
      RECT 22.572 95.74 22.644 98.66 ; 
      RECT 22.572 100.06 22.644 102.98 ; 
      RECT 21.276 79.108 21.348 80.3 ; 
      RECT 21.276 83.86 21.348 84.116 ; 
      RECT 21.276 84.94 21.348 86.78 ; 
      RECT 21.276 89.74 21.348 89.888 ; 
      RECT 21.276 97.9 21.348 99.092 ; 
      RECT 21.132 79.396 21.204 81.416 ; 
      RECT 21.132 82.492 21.204 85.7 ; 
      RECT 21.132 89.872 21.204 90.956 ; 
      RECT 21.132 91.276 21.204 92.18 ; 
      RECT 20.988 79.108 21.06 81.812 ; 
      RECT 20.988 82.204 21.06 83.54 ; 
      RECT 20.988 84.364 21.06 84.908 ; 
      RECT 20.988 87.1 21.06 90.308 ; 
      RECT 20.988 92.044 21.06 92.192 ; 
      RECT 20.988 100.708 21.06 102.044 ; 
      RECT 20.844 80.044 20.916 80.588 ; 
      RECT 20.844 87.604 20.916 91.532 ; 
      RECT 20.844 93.292 20.916 94.484 ; 
      RECT 20.844 100.06 20.916 101.108 ; 
      RECT 20.7 76.3 20.772 76.916 ; 
      RECT 20.7 79.54 20.772 86.684 ; 
      RECT 20.7 90.844 20.772 100.172 ; 
      RECT 20.7 100.996 20.772 105.428 ; 
      RECT 19.548 77.38 19.62 78.428 ; 
      RECT 19.548 78.964 19.62 79.22 ; 
      RECT 19.548 79.54 19.62 80.444 ; 
      RECT 19.548 80.62 19.62 81.38 ; 
      RECT 19.548 81.7 19.62 92.18 ; 
      RECT 19.548 92.356 19.62 97.58 ; 
      RECT 19.548 101.932 19.62 102.98 ; 
      RECT 19.404 81.376 19.476 82.46 ; 
      RECT 19.404 82.78 19.476 86.132 ; 
      RECT 19.404 86.812 19.476 90.164 ; 
      RECT 19.404 90.34 19.476 95.42 ; 
      RECT 19.404 96.244 19.476 96.932 ; 
      RECT 19.404 99.772 19.476 104.06 ; 
      RECT 19.26 81.7 19.332 82.784 ; 
      RECT 19.26 83.404 19.332 83.552 ; 
      RECT 19.26 86.524 19.332 90.452 ; 
      RECT 19.26 91.42 19.332 93.26 ; 
      RECT 19.26 94.66 19.332 97.616 ; 
      RECT 19.116 78.172 19.188 82.46 ; 
      RECT 19.116 88.828 19.188 89.696 ; 
      RECT 19.116 94.372 19.188 95.564 ; 
      RECT 18.972 80.764 19.044 82.604 ; 
      RECT 18.972 87.1 19.044 87.86 ; 
      RECT 18.972 88.024 19.044 88.172 ; 
      RECT 18.972 89.116 19.044 90.452 ; 
      RECT 18.972 90.988 19.044 96.356 ; 
      RECT 18.972 96.784 19.044 101.252 ; 
      RECT 18.828 78.46 18.9 79.22 ; 
      RECT 18.828 80.044 18.9 80.588 ; 
      RECT 18.828 81.7 18.9 94.34 ; 
      RECT 18.828 94.66 18.9 96.5 ; 
      RECT 18.828 98.98 18.9 100.82 ; 
      RECT 18.828 104.236 18.9 105.14 ; 
      RECT 18.684 74.412 18.756 75.028 ; 
      RECT 18.684 106.456 18.756 107.072 ; 
      RECT 18.54 74.412 18.612 74.612 ; 
      RECT 18.252 74.412 18.324 74.698 ; 
      RECT 18.252 106.734 18.324 107.134 ; 
      RECT 17.676 80.476 17.748 81.236 ; 
      RECT 17.676 83.428 17.748 84.908 ; 
      RECT 17.676 91.276 17.748 92.18 ; 
      RECT 17.676 93.436 17.748 98.012 ; 
      RECT 17.676 101.14 17.748 102.98 ; 
      RECT 17.676 105.292 17.748 105.44 ; 
      RECT 17.532 76.3 17.604 78.284 ; 
      RECT 17.532 92.62 17.604 92.768 ; 
      RECT 17.532 96.928 17.604 100.172 ; 
      RECT 17.388 78.172 17.46 79.22 ; 
      RECT 17.388 80.332 17.46 81.668 ; 
      RECT 17.388 82.492 17.46 82.892 ; 
      RECT 17.388 86.02 17.46 97.076 ; 
      RECT 17.388 97.612 17.46 98.516 ; 
      RECT 17.244 76.804 17.316 81.38 ; 
      RECT 17.244 95.74 17.316 96.5 ; 
      RECT 17.244 98.956 17.316 99.104 ; 
      RECT 17.244 100.06 17.316 103.268 ; 
      RECT 17.1 80.62 17.172 84.62 ; 
      RECT 17.1 98.38 17.172 98.528 ; 
      RECT 16.956 77.38 17.028 77.492 ; 
      RECT 15.66 78.964 15.732 80.588 ; 
      RECT 15.372 79.108 15.444 81.524 ; 
      RECT 15.228 78.46 15.3 78.716 ; 
      RECT 15.084 74.624 15.156 74.828 ; 
      RECT 15.084 87.1 15.156 87.86 ; 
      RECT 15.084 89.584 15.156 107.024 ; 
      RECT 14.724 89.584 14.796 107.024 ; 
      RECT 14.652 76.3 14.724 77.06 ; 
      RECT 14.652 79.396 14.724 88.436 ; 
      RECT 14.58 90.804 14.652 91.136 ; 
      RECT 14.436 74.306 14.508 107.134 ; 
      RECT 14.292 89.714 14.364 92.474 ; 
      RECT 14.292 92.678 14.364 96.644 ; 
      RECT 14.292 96.764 14.364 99.9 ; 
      RECT 14.22 76.3 14.292 78.284 ; 
      RECT 14.22 81.412 14.292 83.684 ; 
      RECT 14.22 84.94 14.292 87.86 ; 
      RECT 14.148 89.46 14.22 92.2788 ; 
      RECT 14.148 95.248 14.22 99.972 ; 
      RECT 14.004 74.306 14.076 75.706 ; 
      RECT 13.572 74.306 13.644 75.706 ; 
      RECT 13.14 74.306 13.212 75.706 ; 
      RECT 12.708 74.306 12.78 75.706 ; 
      RECT 12.276 74.306 12.348 75.706 ; 
      RECT 11.844 74.306 11.916 75.706 ; 
      RECT 11.412 74.306 11.484 75.706 ; 
      RECT 10.98 74.306 11.052 75.706 ; 
      RECT 10.548 74.306 10.62 75.706 ; 
      RECT 10.116 74.306 10.188 75.706 ; 
      RECT 9.684 74.306 9.756 75.706 ; 
      RECT 9.252 74.306 9.324 75.706 ; 
      RECT 8.82 74.306 8.892 75.706 ; 
      RECT 8.388 74.306 8.46 75.706 ; 
      RECT 7.956 74.306 8.028 75.706 ; 
      RECT 7.524 74.306 7.596 75.706 ; 
      RECT 7.092 74.306 7.164 75.706 ; 
      RECT 6.66 74.306 6.732 75.706 ; 
      RECT 6.228 74.306 6.3 75.706 ; 
      RECT 5.796 74.306 5.868 75.706 ; 
      RECT 5.364 74.306 5.436 75.706 ; 
      RECT 4.932 74.306 5.004 75.706 ; 
      RECT 4.5 74.306 4.572 75.706 ; 
      RECT 4.068 74.306 4.14 75.706 ; 
      RECT 3.636 74.306 3.708 75.706 ; 
      RECT 3.204 74.306 3.276 75.706 ; 
      RECT 2.772 74.306 2.844 75.706 ; 
      RECT 2.34 74.306 2.412 75.706 ; 
      RECT 1.908 74.306 1.98 75.706 ; 
      RECT 1.476 74.306 1.548 75.706 ; 
      RECT 1.332 89.726 1.404 92.294 ; 
      RECT 1.332 95.004 1.404 97.132 ; 
      RECT 1.26 78.46 1.332 79.364 ; 
      RECT 1.188 89.384 1.26 92.474 ; 
      RECT 1.188 92.6788 1.26 94.644 ; 
      RECT 1.188 94.844 1.26 96.33 ; 
      RECT 1.188 96.582 1.26 99.828 ; 
      RECT 1.044 74.306 1.116 107.134 ; 
      RECT 0.9 84.324 0.972 84.6 ; 
      RECT 0.9 91.556 0.972 93.414 ; 
      RECT 0.756 89.584 0.828 107.006 ; 
        RECT 20.952 107.328 21.024 111.07 ; 
        RECT 20.808 107.328 20.88 111.07 ; 
        RECT 20.664 109.636 20.736 110.926 ; 
        RECT 20.196 110.424 20.268 110.862 ; 
        RECT 20.16 107.458 20.232 108.416 ; 
        RECT 20.016 109.782 20.088 110.396 ; 
        RECT 19.692 109.884 19.764 110.916 ; 
        RECT 17.532 107.328 17.604 111.07 ; 
        RECT 17.388 107.328 17.46 111.07 ; 
        RECT 17.244 108.052 17.316 110.324 ; 
        RECT 20.952 111.648 21.024 115.39 ; 
        RECT 20.808 111.648 20.88 115.39 ; 
        RECT 20.664 113.956 20.736 115.246 ; 
        RECT 20.196 114.744 20.268 115.182 ; 
        RECT 20.16 111.778 20.232 112.736 ; 
        RECT 20.016 114.102 20.088 114.716 ; 
        RECT 19.692 114.204 19.764 115.236 ; 
        RECT 17.532 111.648 17.604 115.39 ; 
        RECT 17.388 111.648 17.46 115.39 ; 
        RECT 17.244 112.372 17.316 114.644 ; 
        RECT 20.952 115.968 21.024 119.71 ; 
        RECT 20.808 115.968 20.88 119.71 ; 
        RECT 20.664 118.276 20.736 119.566 ; 
        RECT 20.196 119.064 20.268 119.502 ; 
        RECT 20.16 116.098 20.232 117.056 ; 
        RECT 20.016 118.422 20.088 119.036 ; 
        RECT 19.692 118.524 19.764 119.556 ; 
        RECT 17.532 115.968 17.604 119.71 ; 
        RECT 17.388 115.968 17.46 119.71 ; 
        RECT 17.244 116.692 17.316 118.964 ; 
        RECT 20.952 120.288 21.024 124.03 ; 
        RECT 20.808 120.288 20.88 124.03 ; 
        RECT 20.664 122.596 20.736 123.886 ; 
        RECT 20.196 123.384 20.268 123.822 ; 
        RECT 20.16 120.418 20.232 121.376 ; 
        RECT 20.016 122.742 20.088 123.356 ; 
        RECT 19.692 122.844 19.764 123.876 ; 
        RECT 17.532 120.288 17.604 124.03 ; 
        RECT 17.388 120.288 17.46 124.03 ; 
        RECT 17.244 121.012 17.316 123.284 ; 
        RECT 20.952 124.608 21.024 128.35 ; 
        RECT 20.808 124.608 20.88 128.35 ; 
        RECT 20.664 126.916 20.736 128.206 ; 
        RECT 20.196 127.704 20.268 128.142 ; 
        RECT 20.16 124.738 20.232 125.696 ; 
        RECT 20.016 127.062 20.088 127.676 ; 
        RECT 19.692 127.164 19.764 128.196 ; 
        RECT 17.532 124.608 17.604 128.35 ; 
        RECT 17.388 124.608 17.46 128.35 ; 
        RECT 17.244 125.332 17.316 127.604 ; 
        RECT 20.952 128.928 21.024 132.67 ; 
        RECT 20.808 128.928 20.88 132.67 ; 
        RECT 20.664 131.236 20.736 132.526 ; 
        RECT 20.196 132.024 20.268 132.462 ; 
        RECT 20.16 129.058 20.232 130.016 ; 
        RECT 20.016 131.382 20.088 131.996 ; 
        RECT 19.692 131.484 19.764 132.516 ; 
        RECT 17.532 128.928 17.604 132.67 ; 
        RECT 17.388 128.928 17.46 132.67 ; 
        RECT 17.244 129.652 17.316 131.924 ; 
        RECT 20.952 133.248 21.024 136.99 ; 
        RECT 20.808 133.248 20.88 136.99 ; 
        RECT 20.664 135.556 20.736 136.846 ; 
        RECT 20.196 136.344 20.268 136.782 ; 
        RECT 20.16 133.378 20.232 134.336 ; 
        RECT 20.016 135.702 20.088 136.316 ; 
        RECT 19.692 135.804 19.764 136.836 ; 
        RECT 17.532 133.248 17.604 136.99 ; 
        RECT 17.388 133.248 17.46 136.99 ; 
        RECT 17.244 133.972 17.316 136.244 ; 
        RECT 20.952 137.568 21.024 141.31 ; 
        RECT 20.808 137.568 20.88 141.31 ; 
        RECT 20.664 139.876 20.736 141.166 ; 
        RECT 20.196 140.664 20.268 141.102 ; 
        RECT 20.16 137.698 20.232 138.656 ; 
        RECT 20.016 140.022 20.088 140.636 ; 
        RECT 19.692 140.124 19.764 141.156 ; 
        RECT 17.532 137.568 17.604 141.31 ; 
        RECT 17.388 137.568 17.46 141.31 ; 
        RECT 17.244 138.292 17.316 140.564 ; 
        RECT 20.952 141.888 21.024 145.63 ; 
        RECT 20.808 141.888 20.88 145.63 ; 
        RECT 20.664 144.196 20.736 145.486 ; 
        RECT 20.196 144.984 20.268 145.422 ; 
        RECT 20.16 142.018 20.232 142.976 ; 
        RECT 20.016 144.342 20.088 144.956 ; 
        RECT 19.692 144.444 19.764 145.476 ; 
        RECT 17.532 141.888 17.604 145.63 ; 
        RECT 17.388 141.888 17.46 145.63 ; 
        RECT 17.244 142.612 17.316 144.884 ; 
        RECT 20.952 146.208 21.024 149.95 ; 
        RECT 20.808 146.208 20.88 149.95 ; 
        RECT 20.664 148.516 20.736 149.806 ; 
        RECT 20.196 149.304 20.268 149.742 ; 
        RECT 20.16 146.338 20.232 147.296 ; 
        RECT 20.016 148.662 20.088 149.276 ; 
        RECT 19.692 148.764 19.764 149.796 ; 
        RECT 17.532 146.208 17.604 149.95 ; 
        RECT 17.388 146.208 17.46 149.95 ; 
        RECT 17.244 146.932 17.316 149.204 ; 
        RECT 20.952 150.528 21.024 154.27 ; 
        RECT 20.808 150.528 20.88 154.27 ; 
        RECT 20.664 152.836 20.736 154.126 ; 
        RECT 20.196 153.624 20.268 154.062 ; 
        RECT 20.16 150.658 20.232 151.616 ; 
        RECT 20.016 152.982 20.088 153.596 ; 
        RECT 19.692 153.084 19.764 154.116 ; 
        RECT 17.532 150.528 17.604 154.27 ; 
        RECT 17.388 150.528 17.46 154.27 ; 
        RECT 17.244 151.252 17.316 153.524 ; 
        RECT 20.952 154.848 21.024 158.59 ; 
        RECT 20.808 154.848 20.88 158.59 ; 
        RECT 20.664 157.156 20.736 158.446 ; 
        RECT 20.196 157.944 20.268 158.382 ; 
        RECT 20.16 154.978 20.232 155.936 ; 
        RECT 20.016 157.302 20.088 157.916 ; 
        RECT 19.692 157.404 19.764 158.436 ; 
        RECT 17.532 154.848 17.604 158.59 ; 
        RECT 17.388 154.848 17.46 158.59 ; 
        RECT 17.244 155.572 17.316 157.844 ; 
        RECT 20.952 159.168 21.024 162.91 ; 
        RECT 20.808 159.168 20.88 162.91 ; 
        RECT 20.664 161.476 20.736 162.766 ; 
        RECT 20.196 162.264 20.268 162.702 ; 
        RECT 20.16 159.298 20.232 160.256 ; 
        RECT 20.016 161.622 20.088 162.236 ; 
        RECT 19.692 161.724 19.764 162.756 ; 
        RECT 17.532 159.168 17.604 162.91 ; 
        RECT 17.388 159.168 17.46 162.91 ; 
        RECT 17.244 159.892 17.316 162.164 ; 
        RECT 20.952 163.488 21.024 167.23 ; 
        RECT 20.808 163.488 20.88 167.23 ; 
        RECT 20.664 165.796 20.736 167.086 ; 
        RECT 20.196 166.584 20.268 167.022 ; 
        RECT 20.16 163.618 20.232 164.576 ; 
        RECT 20.016 165.942 20.088 166.556 ; 
        RECT 19.692 166.044 19.764 167.076 ; 
        RECT 17.532 163.488 17.604 167.23 ; 
        RECT 17.388 163.488 17.46 167.23 ; 
        RECT 17.244 164.212 17.316 166.484 ; 
        RECT 20.952 167.808 21.024 171.55 ; 
        RECT 20.808 167.808 20.88 171.55 ; 
        RECT 20.664 170.116 20.736 171.406 ; 
        RECT 20.196 170.904 20.268 171.342 ; 
        RECT 20.16 167.938 20.232 168.896 ; 
        RECT 20.016 170.262 20.088 170.876 ; 
        RECT 19.692 170.364 19.764 171.396 ; 
        RECT 17.532 167.808 17.604 171.55 ; 
        RECT 17.388 167.808 17.46 171.55 ; 
        RECT 17.244 168.532 17.316 170.804 ; 
        RECT 20.952 172.128 21.024 175.87 ; 
        RECT 20.808 172.128 20.88 175.87 ; 
        RECT 20.664 174.436 20.736 175.726 ; 
        RECT 20.196 175.224 20.268 175.662 ; 
        RECT 20.16 172.258 20.232 173.216 ; 
        RECT 20.016 174.582 20.088 175.196 ; 
        RECT 19.692 174.684 19.764 175.716 ; 
        RECT 17.532 172.128 17.604 175.87 ; 
        RECT 17.388 172.128 17.46 175.87 ; 
        RECT 17.244 172.852 17.316 175.124 ; 
        RECT 20.952 176.448 21.024 180.19 ; 
        RECT 20.808 176.448 20.88 180.19 ; 
        RECT 20.664 178.756 20.736 180.046 ; 
        RECT 20.196 179.544 20.268 179.982 ; 
        RECT 20.16 176.578 20.232 177.536 ; 
        RECT 20.016 178.902 20.088 179.516 ; 
        RECT 19.692 179.004 19.764 180.036 ; 
        RECT 17.532 176.448 17.604 180.19 ; 
        RECT 17.388 176.448 17.46 180.19 ; 
        RECT 17.244 177.172 17.316 179.444 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 20.72 1.026 21.232 5.4 ; 
      RECT 20.664 3.688 21.232 4.978 ; 
      RECT 20.072 2.596 20.32 5.4 ; 
      RECT 20.016 3.834 20.32 4.448 ; 
      RECT 20.072 1.026 20.176 5.4 ; 
      RECT 20.072 1.51 20.232 2.468 ; 
      RECT 20.072 1.026 20.32 1.382 ; 
      RECT 18.884 2.828 19.708 5.4 ; 
      RECT 19.604 1.026 19.708 5.4 ; 
      RECT 18.884 3.936 19.764 4.968 ; 
      RECT 18.884 1.026 19.276 5.4 ; 
      RECT 17.216 1.026 17.548 5.4 ; 
      RECT 17.216 1.38 17.604 5.122 ; 
      RECT 38.108 1.026 38.448 5.4 ; 
      RECT 37.532 1.026 37.636 5.4 ; 
      RECT 37.1 1.026 37.204 5.4 ; 
      RECT 36.668 1.026 36.772 5.4 ; 
      RECT 36.236 1.026 36.34 5.4 ; 
      RECT 35.804 1.026 35.908 5.4 ; 
      RECT 35.372 1.026 35.476 5.4 ; 
      RECT 34.94 1.026 35.044 5.4 ; 
      RECT 34.508 1.026 34.612 5.4 ; 
      RECT 34.076 1.026 34.18 5.4 ; 
      RECT 33.644 1.026 33.748 5.4 ; 
      RECT 33.212 1.026 33.316 5.4 ; 
      RECT 32.78 1.026 32.884 5.4 ; 
      RECT 32.348 1.026 32.452 5.4 ; 
      RECT 31.916 1.026 32.02 5.4 ; 
      RECT 31.484 1.026 31.588 5.4 ; 
      RECT 31.052 1.026 31.156 5.4 ; 
      RECT 30.62 1.026 30.724 5.4 ; 
      RECT 30.188 1.026 30.292 5.4 ; 
      RECT 29.756 1.026 29.86 5.4 ; 
      RECT 29.324 1.026 29.428 5.4 ; 
      RECT 28.892 1.026 28.996 5.4 ; 
      RECT 28.46 1.026 28.564 5.4 ; 
      RECT 28.028 1.026 28.132 5.4 ; 
      RECT 27.596 1.026 27.7 5.4 ; 
      RECT 27.164 1.026 27.268 5.4 ; 
      RECT 26.732 1.026 26.836 5.4 ; 
      RECT 26.3 1.026 26.404 5.4 ; 
      RECT 25.868 1.026 25.972 5.4 ; 
      RECT 25.436 1.026 25.54 5.4 ; 
      RECT 25.004 1.026 25.108 5.4 ; 
      RECT 24.572 1.026 24.676 5.4 ; 
      RECT 24.14 1.026 24.244 5.4 ; 
      RECT 23.708 1.026 23.812 5.4 ; 
      RECT 22.856 1.026 23.164 5.4 ; 
      RECT 15.284 1.026 15.592 5.4 ; 
      RECT 14.636 1.026 14.74 5.4 ; 
      RECT 14.204 1.026 14.308 5.4 ; 
      RECT 13.772 1.026 13.876 5.4 ; 
      RECT 13.34 1.026 13.444 5.4 ; 
      RECT 12.908 1.026 13.012 5.4 ; 
      RECT 12.476 1.026 12.58 5.4 ; 
      RECT 12.044 1.026 12.148 5.4 ; 
      RECT 11.612 1.026 11.716 5.4 ; 
      RECT 11.18 1.026 11.284 5.4 ; 
      RECT 10.748 1.026 10.852 5.4 ; 
      RECT 10.316 1.026 10.42 5.4 ; 
      RECT 9.884 1.026 9.988 5.4 ; 
      RECT 9.452 1.026 9.556 5.4 ; 
      RECT 9.02 1.026 9.124 5.4 ; 
      RECT 8.588 1.026 8.692 5.4 ; 
      RECT 8.156 1.026 8.26 5.4 ; 
      RECT 7.724 1.026 7.828 5.4 ; 
      RECT 7.292 1.026 7.396 5.4 ; 
      RECT 6.86 1.026 6.964 5.4 ; 
      RECT 6.428 1.026 6.532 5.4 ; 
      RECT 5.996 1.026 6.1 5.4 ; 
      RECT 5.564 1.026 5.668 5.4 ; 
      RECT 5.132 1.026 5.236 5.4 ; 
      RECT 4.7 1.026 4.804 5.4 ; 
      RECT 4.268 1.026 4.372 5.4 ; 
      RECT 3.836 1.026 3.94 5.4 ; 
      RECT 3.404 1.026 3.508 5.4 ; 
      RECT 2.972 1.026 3.076 5.4 ; 
      RECT 2.54 1.026 2.644 5.4 ; 
      RECT 2.108 1.026 2.212 5.4 ; 
      RECT 1.676 1.026 1.78 5.4 ; 
      RECT 1.244 1.026 1.348 5.4 ; 
      RECT 0.812 1.026 0.916 5.4 ; 
      RECT 0 1.026 0.34 5.4 ; 
      RECT 20.72 5.346 21.232 9.72 ; 
      RECT 20.664 8.008 21.232 9.298 ; 
      RECT 20.072 6.916 20.32 9.72 ; 
      RECT 20.016 8.154 20.32 8.768 ; 
      RECT 20.072 5.346 20.176 9.72 ; 
      RECT 20.072 5.83 20.232 6.788 ; 
      RECT 20.072 5.346 20.32 5.702 ; 
      RECT 18.884 7.148 19.708 9.72 ; 
      RECT 19.604 5.346 19.708 9.72 ; 
      RECT 18.884 8.256 19.764 9.288 ; 
      RECT 18.884 5.346 19.276 9.72 ; 
      RECT 17.216 5.346 17.548 9.72 ; 
      RECT 17.216 5.7 17.604 9.442 ; 
      RECT 38.108 5.346 38.448 9.72 ; 
      RECT 37.532 5.346 37.636 9.72 ; 
      RECT 37.1 5.346 37.204 9.72 ; 
      RECT 36.668 5.346 36.772 9.72 ; 
      RECT 36.236 5.346 36.34 9.72 ; 
      RECT 35.804 5.346 35.908 9.72 ; 
      RECT 35.372 5.346 35.476 9.72 ; 
      RECT 34.94 5.346 35.044 9.72 ; 
      RECT 34.508 5.346 34.612 9.72 ; 
      RECT 34.076 5.346 34.18 9.72 ; 
      RECT 33.644 5.346 33.748 9.72 ; 
      RECT 33.212 5.346 33.316 9.72 ; 
      RECT 32.78 5.346 32.884 9.72 ; 
      RECT 32.348 5.346 32.452 9.72 ; 
      RECT 31.916 5.346 32.02 9.72 ; 
      RECT 31.484 5.346 31.588 9.72 ; 
      RECT 31.052 5.346 31.156 9.72 ; 
      RECT 30.62 5.346 30.724 9.72 ; 
      RECT 30.188 5.346 30.292 9.72 ; 
      RECT 29.756 5.346 29.86 9.72 ; 
      RECT 29.324 5.346 29.428 9.72 ; 
      RECT 28.892 5.346 28.996 9.72 ; 
      RECT 28.46 5.346 28.564 9.72 ; 
      RECT 28.028 5.346 28.132 9.72 ; 
      RECT 27.596 5.346 27.7 9.72 ; 
      RECT 27.164 5.346 27.268 9.72 ; 
      RECT 26.732 5.346 26.836 9.72 ; 
      RECT 26.3 5.346 26.404 9.72 ; 
      RECT 25.868 5.346 25.972 9.72 ; 
      RECT 25.436 5.346 25.54 9.72 ; 
      RECT 25.004 5.346 25.108 9.72 ; 
      RECT 24.572 5.346 24.676 9.72 ; 
      RECT 24.14 5.346 24.244 9.72 ; 
      RECT 23.708 5.346 23.812 9.72 ; 
      RECT 22.856 5.346 23.164 9.72 ; 
      RECT 15.284 5.346 15.592 9.72 ; 
      RECT 14.636 5.346 14.74 9.72 ; 
      RECT 14.204 5.346 14.308 9.72 ; 
      RECT 13.772 5.346 13.876 9.72 ; 
      RECT 13.34 5.346 13.444 9.72 ; 
      RECT 12.908 5.346 13.012 9.72 ; 
      RECT 12.476 5.346 12.58 9.72 ; 
      RECT 12.044 5.346 12.148 9.72 ; 
      RECT 11.612 5.346 11.716 9.72 ; 
      RECT 11.18 5.346 11.284 9.72 ; 
      RECT 10.748 5.346 10.852 9.72 ; 
      RECT 10.316 5.346 10.42 9.72 ; 
      RECT 9.884 5.346 9.988 9.72 ; 
      RECT 9.452 5.346 9.556 9.72 ; 
      RECT 9.02 5.346 9.124 9.72 ; 
      RECT 8.588 5.346 8.692 9.72 ; 
      RECT 8.156 5.346 8.26 9.72 ; 
      RECT 7.724 5.346 7.828 9.72 ; 
      RECT 7.292 5.346 7.396 9.72 ; 
      RECT 6.86 5.346 6.964 9.72 ; 
      RECT 6.428 5.346 6.532 9.72 ; 
      RECT 5.996 5.346 6.1 9.72 ; 
      RECT 5.564 5.346 5.668 9.72 ; 
      RECT 5.132 5.346 5.236 9.72 ; 
      RECT 4.7 5.346 4.804 9.72 ; 
      RECT 4.268 5.346 4.372 9.72 ; 
      RECT 3.836 5.346 3.94 9.72 ; 
      RECT 3.404 5.346 3.508 9.72 ; 
      RECT 2.972 5.346 3.076 9.72 ; 
      RECT 2.54 5.346 2.644 9.72 ; 
      RECT 2.108 5.346 2.212 9.72 ; 
      RECT 1.676 5.346 1.78 9.72 ; 
      RECT 1.244 5.346 1.348 9.72 ; 
      RECT 0.812 5.346 0.916 9.72 ; 
      RECT 0 5.346 0.34 9.72 ; 
      RECT 20.72 9.666 21.232 14.04 ; 
      RECT 20.664 12.328 21.232 13.618 ; 
      RECT 20.072 11.236 20.32 14.04 ; 
      RECT 20.016 12.474 20.32 13.088 ; 
      RECT 20.072 9.666 20.176 14.04 ; 
      RECT 20.072 10.15 20.232 11.108 ; 
      RECT 20.072 9.666 20.32 10.022 ; 
      RECT 18.884 11.468 19.708 14.04 ; 
      RECT 19.604 9.666 19.708 14.04 ; 
      RECT 18.884 12.576 19.764 13.608 ; 
      RECT 18.884 9.666 19.276 14.04 ; 
      RECT 17.216 9.666 17.548 14.04 ; 
      RECT 17.216 10.02 17.604 13.762 ; 
      RECT 38.108 9.666 38.448 14.04 ; 
      RECT 37.532 9.666 37.636 14.04 ; 
      RECT 37.1 9.666 37.204 14.04 ; 
      RECT 36.668 9.666 36.772 14.04 ; 
      RECT 36.236 9.666 36.34 14.04 ; 
      RECT 35.804 9.666 35.908 14.04 ; 
      RECT 35.372 9.666 35.476 14.04 ; 
      RECT 34.94 9.666 35.044 14.04 ; 
      RECT 34.508 9.666 34.612 14.04 ; 
      RECT 34.076 9.666 34.18 14.04 ; 
      RECT 33.644 9.666 33.748 14.04 ; 
      RECT 33.212 9.666 33.316 14.04 ; 
      RECT 32.78 9.666 32.884 14.04 ; 
      RECT 32.348 9.666 32.452 14.04 ; 
      RECT 31.916 9.666 32.02 14.04 ; 
      RECT 31.484 9.666 31.588 14.04 ; 
      RECT 31.052 9.666 31.156 14.04 ; 
      RECT 30.62 9.666 30.724 14.04 ; 
      RECT 30.188 9.666 30.292 14.04 ; 
      RECT 29.756 9.666 29.86 14.04 ; 
      RECT 29.324 9.666 29.428 14.04 ; 
      RECT 28.892 9.666 28.996 14.04 ; 
      RECT 28.46 9.666 28.564 14.04 ; 
      RECT 28.028 9.666 28.132 14.04 ; 
      RECT 27.596 9.666 27.7 14.04 ; 
      RECT 27.164 9.666 27.268 14.04 ; 
      RECT 26.732 9.666 26.836 14.04 ; 
      RECT 26.3 9.666 26.404 14.04 ; 
      RECT 25.868 9.666 25.972 14.04 ; 
      RECT 25.436 9.666 25.54 14.04 ; 
      RECT 25.004 9.666 25.108 14.04 ; 
      RECT 24.572 9.666 24.676 14.04 ; 
      RECT 24.14 9.666 24.244 14.04 ; 
      RECT 23.708 9.666 23.812 14.04 ; 
      RECT 22.856 9.666 23.164 14.04 ; 
      RECT 15.284 9.666 15.592 14.04 ; 
      RECT 14.636 9.666 14.74 14.04 ; 
      RECT 14.204 9.666 14.308 14.04 ; 
      RECT 13.772 9.666 13.876 14.04 ; 
      RECT 13.34 9.666 13.444 14.04 ; 
      RECT 12.908 9.666 13.012 14.04 ; 
      RECT 12.476 9.666 12.58 14.04 ; 
      RECT 12.044 9.666 12.148 14.04 ; 
      RECT 11.612 9.666 11.716 14.04 ; 
      RECT 11.18 9.666 11.284 14.04 ; 
      RECT 10.748 9.666 10.852 14.04 ; 
      RECT 10.316 9.666 10.42 14.04 ; 
      RECT 9.884 9.666 9.988 14.04 ; 
      RECT 9.452 9.666 9.556 14.04 ; 
      RECT 9.02 9.666 9.124 14.04 ; 
      RECT 8.588 9.666 8.692 14.04 ; 
      RECT 8.156 9.666 8.26 14.04 ; 
      RECT 7.724 9.666 7.828 14.04 ; 
      RECT 7.292 9.666 7.396 14.04 ; 
      RECT 6.86 9.666 6.964 14.04 ; 
      RECT 6.428 9.666 6.532 14.04 ; 
      RECT 5.996 9.666 6.1 14.04 ; 
      RECT 5.564 9.666 5.668 14.04 ; 
      RECT 5.132 9.666 5.236 14.04 ; 
      RECT 4.7 9.666 4.804 14.04 ; 
      RECT 4.268 9.666 4.372 14.04 ; 
      RECT 3.836 9.666 3.94 14.04 ; 
      RECT 3.404 9.666 3.508 14.04 ; 
      RECT 2.972 9.666 3.076 14.04 ; 
      RECT 2.54 9.666 2.644 14.04 ; 
      RECT 2.108 9.666 2.212 14.04 ; 
      RECT 1.676 9.666 1.78 14.04 ; 
      RECT 1.244 9.666 1.348 14.04 ; 
      RECT 0.812 9.666 0.916 14.04 ; 
      RECT 0 9.666 0.34 14.04 ; 
      RECT 20.72 13.986 21.232 18.36 ; 
      RECT 20.664 16.648 21.232 17.938 ; 
      RECT 20.072 15.556 20.32 18.36 ; 
      RECT 20.016 16.794 20.32 17.408 ; 
      RECT 20.072 13.986 20.176 18.36 ; 
      RECT 20.072 14.47 20.232 15.428 ; 
      RECT 20.072 13.986 20.32 14.342 ; 
      RECT 18.884 15.788 19.708 18.36 ; 
      RECT 19.604 13.986 19.708 18.36 ; 
      RECT 18.884 16.896 19.764 17.928 ; 
      RECT 18.884 13.986 19.276 18.36 ; 
      RECT 17.216 13.986 17.548 18.36 ; 
      RECT 17.216 14.34 17.604 18.082 ; 
      RECT 38.108 13.986 38.448 18.36 ; 
      RECT 37.532 13.986 37.636 18.36 ; 
      RECT 37.1 13.986 37.204 18.36 ; 
      RECT 36.668 13.986 36.772 18.36 ; 
      RECT 36.236 13.986 36.34 18.36 ; 
      RECT 35.804 13.986 35.908 18.36 ; 
      RECT 35.372 13.986 35.476 18.36 ; 
      RECT 34.94 13.986 35.044 18.36 ; 
      RECT 34.508 13.986 34.612 18.36 ; 
      RECT 34.076 13.986 34.18 18.36 ; 
      RECT 33.644 13.986 33.748 18.36 ; 
      RECT 33.212 13.986 33.316 18.36 ; 
      RECT 32.78 13.986 32.884 18.36 ; 
      RECT 32.348 13.986 32.452 18.36 ; 
      RECT 31.916 13.986 32.02 18.36 ; 
      RECT 31.484 13.986 31.588 18.36 ; 
      RECT 31.052 13.986 31.156 18.36 ; 
      RECT 30.62 13.986 30.724 18.36 ; 
      RECT 30.188 13.986 30.292 18.36 ; 
      RECT 29.756 13.986 29.86 18.36 ; 
      RECT 29.324 13.986 29.428 18.36 ; 
      RECT 28.892 13.986 28.996 18.36 ; 
      RECT 28.46 13.986 28.564 18.36 ; 
      RECT 28.028 13.986 28.132 18.36 ; 
      RECT 27.596 13.986 27.7 18.36 ; 
      RECT 27.164 13.986 27.268 18.36 ; 
      RECT 26.732 13.986 26.836 18.36 ; 
      RECT 26.3 13.986 26.404 18.36 ; 
      RECT 25.868 13.986 25.972 18.36 ; 
      RECT 25.436 13.986 25.54 18.36 ; 
      RECT 25.004 13.986 25.108 18.36 ; 
      RECT 24.572 13.986 24.676 18.36 ; 
      RECT 24.14 13.986 24.244 18.36 ; 
      RECT 23.708 13.986 23.812 18.36 ; 
      RECT 22.856 13.986 23.164 18.36 ; 
      RECT 15.284 13.986 15.592 18.36 ; 
      RECT 14.636 13.986 14.74 18.36 ; 
      RECT 14.204 13.986 14.308 18.36 ; 
      RECT 13.772 13.986 13.876 18.36 ; 
      RECT 13.34 13.986 13.444 18.36 ; 
      RECT 12.908 13.986 13.012 18.36 ; 
      RECT 12.476 13.986 12.58 18.36 ; 
      RECT 12.044 13.986 12.148 18.36 ; 
      RECT 11.612 13.986 11.716 18.36 ; 
      RECT 11.18 13.986 11.284 18.36 ; 
      RECT 10.748 13.986 10.852 18.36 ; 
      RECT 10.316 13.986 10.42 18.36 ; 
      RECT 9.884 13.986 9.988 18.36 ; 
      RECT 9.452 13.986 9.556 18.36 ; 
      RECT 9.02 13.986 9.124 18.36 ; 
      RECT 8.588 13.986 8.692 18.36 ; 
      RECT 8.156 13.986 8.26 18.36 ; 
      RECT 7.724 13.986 7.828 18.36 ; 
      RECT 7.292 13.986 7.396 18.36 ; 
      RECT 6.86 13.986 6.964 18.36 ; 
      RECT 6.428 13.986 6.532 18.36 ; 
      RECT 5.996 13.986 6.1 18.36 ; 
      RECT 5.564 13.986 5.668 18.36 ; 
      RECT 5.132 13.986 5.236 18.36 ; 
      RECT 4.7 13.986 4.804 18.36 ; 
      RECT 4.268 13.986 4.372 18.36 ; 
      RECT 3.836 13.986 3.94 18.36 ; 
      RECT 3.404 13.986 3.508 18.36 ; 
      RECT 2.972 13.986 3.076 18.36 ; 
      RECT 2.54 13.986 2.644 18.36 ; 
      RECT 2.108 13.986 2.212 18.36 ; 
      RECT 1.676 13.986 1.78 18.36 ; 
      RECT 1.244 13.986 1.348 18.36 ; 
      RECT 0.812 13.986 0.916 18.36 ; 
      RECT 0 13.986 0.34 18.36 ; 
      RECT 20.72 18.306 21.232 22.68 ; 
      RECT 20.664 20.968 21.232 22.258 ; 
      RECT 20.072 19.876 20.32 22.68 ; 
      RECT 20.016 21.114 20.32 21.728 ; 
      RECT 20.072 18.306 20.176 22.68 ; 
      RECT 20.072 18.79 20.232 19.748 ; 
      RECT 20.072 18.306 20.32 18.662 ; 
      RECT 18.884 20.108 19.708 22.68 ; 
      RECT 19.604 18.306 19.708 22.68 ; 
      RECT 18.884 21.216 19.764 22.248 ; 
      RECT 18.884 18.306 19.276 22.68 ; 
      RECT 17.216 18.306 17.548 22.68 ; 
      RECT 17.216 18.66 17.604 22.402 ; 
      RECT 38.108 18.306 38.448 22.68 ; 
      RECT 37.532 18.306 37.636 22.68 ; 
      RECT 37.1 18.306 37.204 22.68 ; 
      RECT 36.668 18.306 36.772 22.68 ; 
      RECT 36.236 18.306 36.34 22.68 ; 
      RECT 35.804 18.306 35.908 22.68 ; 
      RECT 35.372 18.306 35.476 22.68 ; 
      RECT 34.94 18.306 35.044 22.68 ; 
      RECT 34.508 18.306 34.612 22.68 ; 
      RECT 34.076 18.306 34.18 22.68 ; 
      RECT 33.644 18.306 33.748 22.68 ; 
      RECT 33.212 18.306 33.316 22.68 ; 
      RECT 32.78 18.306 32.884 22.68 ; 
      RECT 32.348 18.306 32.452 22.68 ; 
      RECT 31.916 18.306 32.02 22.68 ; 
      RECT 31.484 18.306 31.588 22.68 ; 
      RECT 31.052 18.306 31.156 22.68 ; 
      RECT 30.62 18.306 30.724 22.68 ; 
      RECT 30.188 18.306 30.292 22.68 ; 
      RECT 29.756 18.306 29.86 22.68 ; 
      RECT 29.324 18.306 29.428 22.68 ; 
      RECT 28.892 18.306 28.996 22.68 ; 
      RECT 28.46 18.306 28.564 22.68 ; 
      RECT 28.028 18.306 28.132 22.68 ; 
      RECT 27.596 18.306 27.7 22.68 ; 
      RECT 27.164 18.306 27.268 22.68 ; 
      RECT 26.732 18.306 26.836 22.68 ; 
      RECT 26.3 18.306 26.404 22.68 ; 
      RECT 25.868 18.306 25.972 22.68 ; 
      RECT 25.436 18.306 25.54 22.68 ; 
      RECT 25.004 18.306 25.108 22.68 ; 
      RECT 24.572 18.306 24.676 22.68 ; 
      RECT 24.14 18.306 24.244 22.68 ; 
      RECT 23.708 18.306 23.812 22.68 ; 
      RECT 22.856 18.306 23.164 22.68 ; 
      RECT 15.284 18.306 15.592 22.68 ; 
      RECT 14.636 18.306 14.74 22.68 ; 
      RECT 14.204 18.306 14.308 22.68 ; 
      RECT 13.772 18.306 13.876 22.68 ; 
      RECT 13.34 18.306 13.444 22.68 ; 
      RECT 12.908 18.306 13.012 22.68 ; 
      RECT 12.476 18.306 12.58 22.68 ; 
      RECT 12.044 18.306 12.148 22.68 ; 
      RECT 11.612 18.306 11.716 22.68 ; 
      RECT 11.18 18.306 11.284 22.68 ; 
      RECT 10.748 18.306 10.852 22.68 ; 
      RECT 10.316 18.306 10.42 22.68 ; 
      RECT 9.884 18.306 9.988 22.68 ; 
      RECT 9.452 18.306 9.556 22.68 ; 
      RECT 9.02 18.306 9.124 22.68 ; 
      RECT 8.588 18.306 8.692 22.68 ; 
      RECT 8.156 18.306 8.26 22.68 ; 
      RECT 7.724 18.306 7.828 22.68 ; 
      RECT 7.292 18.306 7.396 22.68 ; 
      RECT 6.86 18.306 6.964 22.68 ; 
      RECT 6.428 18.306 6.532 22.68 ; 
      RECT 5.996 18.306 6.1 22.68 ; 
      RECT 5.564 18.306 5.668 22.68 ; 
      RECT 5.132 18.306 5.236 22.68 ; 
      RECT 4.7 18.306 4.804 22.68 ; 
      RECT 4.268 18.306 4.372 22.68 ; 
      RECT 3.836 18.306 3.94 22.68 ; 
      RECT 3.404 18.306 3.508 22.68 ; 
      RECT 2.972 18.306 3.076 22.68 ; 
      RECT 2.54 18.306 2.644 22.68 ; 
      RECT 2.108 18.306 2.212 22.68 ; 
      RECT 1.676 18.306 1.78 22.68 ; 
      RECT 1.244 18.306 1.348 22.68 ; 
      RECT 0.812 18.306 0.916 22.68 ; 
      RECT 0 18.306 0.34 22.68 ; 
      RECT 20.72 22.626 21.232 27 ; 
      RECT 20.664 25.288 21.232 26.578 ; 
      RECT 20.072 24.196 20.32 27 ; 
      RECT 20.016 25.434 20.32 26.048 ; 
      RECT 20.072 22.626 20.176 27 ; 
      RECT 20.072 23.11 20.232 24.068 ; 
      RECT 20.072 22.626 20.32 22.982 ; 
      RECT 18.884 24.428 19.708 27 ; 
      RECT 19.604 22.626 19.708 27 ; 
      RECT 18.884 25.536 19.764 26.568 ; 
      RECT 18.884 22.626 19.276 27 ; 
      RECT 17.216 22.626 17.548 27 ; 
      RECT 17.216 22.98 17.604 26.722 ; 
      RECT 38.108 22.626 38.448 27 ; 
      RECT 37.532 22.626 37.636 27 ; 
      RECT 37.1 22.626 37.204 27 ; 
      RECT 36.668 22.626 36.772 27 ; 
      RECT 36.236 22.626 36.34 27 ; 
      RECT 35.804 22.626 35.908 27 ; 
      RECT 35.372 22.626 35.476 27 ; 
      RECT 34.94 22.626 35.044 27 ; 
      RECT 34.508 22.626 34.612 27 ; 
      RECT 34.076 22.626 34.18 27 ; 
      RECT 33.644 22.626 33.748 27 ; 
      RECT 33.212 22.626 33.316 27 ; 
      RECT 32.78 22.626 32.884 27 ; 
      RECT 32.348 22.626 32.452 27 ; 
      RECT 31.916 22.626 32.02 27 ; 
      RECT 31.484 22.626 31.588 27 ; 
      RECT 31.052 22.626 31.156 27 ; 
      RECT 30.62 22.626 30.724 27 ; 
      RECT 30.188 22.626 30.292 27 ; 
      RECT 29.756 22.626 29.86 27 ; 
      RECT 29.324 22.626 29.428 27 ; 
      RECT 28.892 22.626 28.996 27 ; 
      RECT 28.46 22.626 28.564 27 ; 
      RECT 28.028 22.626 28.132 27 ; 
      RECT 27.596 22.626 27.7 27 ; 
      RECT 27.164 22.626 27.268 27 ; 
      RECT 26.732 22.626 26.836 27 ; 
      RECT 26.3 22.626 26.404 27 ; 
      RECT 25.868 22.626 25.972 27 ; 
      RECT 25.436 22.626 25.54 27 ; 
      RECT 25.004 22.626 25.108 27 ; 
      RECT 24.572 22.626 24.676 27 ; 
      RECT 24.14 22.626 24.244 27 ; 
      RECT 23.708 22.626 23.812 27 ; 
      RECT 22.856 22.626 23.164 27 ; 
      RECT 15.284 22.626 15.592 27 ; 
      RECT 14.636 22.626 14.74 27 ; 
      RECT 14.204 22.626 14.308 27 ; 
      RECT 13.772 22.626 13.876 27 ; 
      RECT 13.34 22.626 13.444 27 ; 
      RECT 12.908 22.626 13.012 27 ; 
      RECT 12.476 22.626 12.58 27 ; 
      RECT 12.044 22.626 12.148 27 ; 
      RECT 11.612 22.626 11.716 27 ; 
      RECT 11.18 22.626 11.284 27 ; 
      RECT 10.748 22.626 10.852 27 ; 
      RECT 10.316 22.626 10.42 27 ; 
      RECT 9.884 22.626 9.988 27 ; 
      RECT 9.452 22.626 9.556 27 ; 
      RECT 9.02 22.626 9.124 27 ; 
      RECT 8.588 22.626 8.692 27 ; 
      RECT 8.156 22.626 8.26 27 ; 
      RECT 7.724 22.626 7.828 27 ; 
      RECT 7.292 22.626 7.396 27 ; 
      RECT 6.86 22.626 6.964 27 ; 
      RECT 6.428 22.626 6.532 27 ; 
      RECT 5.996 22.626 6.1 27 ; 
      RECT 5.564 22.626 5.668 27 ; 
      RECT 5.132 22.626 5.236 27 ; 
      RECT 4.7 22.626 4.804 27 ; 
      RECT 4.268 22.626 4.372 27 ; 
      RECT 3.836 22.626 3.94 27 ; 
      RECT 3.404 22.626 3.508 27 ; 
      RECT 2.972 22.626 3.076 27 ; 
      RECT 2.54 22.626 2.644 27 ; 
      RECT 2.108 22.626 2.212 27 ; 
      RECT 1.676 22.626 1.78 27 ; 
      RECT 1.244 22.626 1.348 27 ; 
      RECT 0.812 22.626 0.916 27 ; 
      RECT 0 22.626 0.34 27 ; 
      RECT 20.72 26.946 21.232 31.32 ; 
      RECT 20.664 29.608 21.232 30.898 ; 
      RECT 20.072 28.516 20.32 31.32 ; 
      RECT 20.016 29.754 20.32 30.368 ; 
      RECT 20.072 26.946 20.176 31.32 ; 
      RECT 20.072 27.43 20.232 28.388 ; 
      RECT 20.072 26.946 20.32 27.302 ; 
      RECT 18.884 28.748 19.708 31.32 ; 
      RECT 19.604 26.946 19.708 31.32 ; 
      RECT 18.884 29.856 19.764 30.888 ; 
      RECT 18.884 26.946 19.276 31.32 ; 
      RECT 17.216 26.946 17.548 31.32 ; 
      RECT 17.216 27.3 17.604 31.042 ; 
      RECT 38.108 26.946 38.448 31.32 ; 
      RECT 37.532 26.946 37.636 31.32 ; 
      RECT 37.1 26.946 37.204 31.32 ; 
      RECT 36.668 26.946 36.772 31.32 ; 
      RECT 36.236 26.946 36.34 31.32 ; 
      RECT 35.804 26.946 35.908 31.32 ; 
      RECT 35.372 26.946 35.476 31.32 ; 
      RECT 34.94 26.946 35.044 31.32 ; 
      RECT 34.508 26.946 34.612 31.32 ; 
      RECT 34.076 26.946 34.18 31.32 ; 
      RECT 33.644 26.946 33.748 31.32 ; 
      RECT 33.212 26.946 33.316 31.32 ; 
      RECT 32.78 26.946 32.884 31.32 ; 
      RECT 32.348 26.946 32.452 31.32 ; 
      RECT 31.916 26.946 32.02 31.32 ; 
      RECT 31.484 26.946 31.588 31.32 ; 
      RECT 31.052 26.946 31.156 31.32 ; 
      RECT 30.62 26.946 30.724 31.32 ; 
      RECT 30.188 26.946 30.292 31.32 ; 
      RECT 29.756 26.946 29.86 31.32 ; 
      RECT 29.324 26.946 29.428 31.32 ; 
      RECT 28.892 26.946 28.996 31.32 ; 
      RECT 28.46 26.946 28.564 31.32 ; 
      RECT 28.028 26.946 28.132 31.32 ; 
      RECT 27.596 26.946 27.7 31.32 ; 
      RECT 27.164 26.946 27.268 31.32 ; 
      RECT 26.732 26.946 26.836 31.32 ; 
      RECT 26.3 26.946 26.404 31.32 ; 
      RECT 25.868 26.946 25.972 31.32 ; 
      RECT 25.436 26.946 25.54 31.32 ; 
      RECT 25.004 26.946 25.108 31.32 ; 
      RECT 24.572 26.946 24.676 31.32 ; 
      RECT 24.14 26.946 24.244 31.32 ; 
      RECT 23.708 26.946 23.812 31.32 ; 
      RECT 22.856 26.946 23.164 31.32 ; 
      RECT 15.284 26.946 15.592 31.32 ; 
      RECT 14.636 26.946 14.74 31.32 ; 
      RECT 14.204 26.946 14.308 31.32 ; 
      RECT 13.772 26.946 13.876 31.32 ; 
      RECT 13.34 26.946 13.444 31.32 ; 
      RECT 12.908 26.946 13.012 31.32 ; 
      RECT 12.476 26.946 12.58 31.32 ; 
      RECT 12.044 26.946 12.148 31.32 ; 
      RECT 11.612 26.946 11.716 31.32 ; 
      RECT 11.18 26.946 11.284 31.32 ; 
      RECT 10.748 26.946 10.852 31.32 ; 
      RECT 10.316 26.946 10.42 31.32 ; 
      RECT 9.884 26.946 9.988 31.32 ; 
      RECT 9.452 26.946 9.556 31.32 ; 
      RECT 9.02 26.946 9.124 31.32 ; 
      RECT 8.588 26.946 8.692 31.32 ; 
      RECT 8.156 26.946 8.26 31.32 ; 
      RECT 7.724 26.946 7.828 31.32 ; 
      RECT 7.292 26.946 7.396 31.32 ; 
      RECT 6.86 26.946 6.964 31.32 ; 
      RECT 6.428 26.946 6.532 31.32 ; 
      RECT 5.996 26.946 6.1 31.32 ; 
      RECT 5.564 26.946 5.668 31.32 ; 
      RECT 5.132 26.946 5.236 31.32 ; 
      RECT 4.7 26.946 4.804 31.32 ; 
      RECT 4.268 26.946 4.372 31.32 ; 
      RECT 3.836 26.946 3.94 31.32 ; 
      RECT 3.404 26.946 3.508 31.32 ; 
      RECT 2.972 26.946 3.076 31.32 ; 
      RECT 2.54 26.946 2.644 31.32 ; 
      RECT 2.108 26.946 2.212 31.32 ; 
      RECT 1.676 26.946 1.78 31.32 ; 
      RECT 1.244 26.946 1.348 31.32 ; 
      RECT 0.812 26.946 0.916 31.32 ; 
      RECT 0 26.946 0.34 31.32 ; 
      RECT 20.72 31.266 21.232 35.64 ; 
      RECT 20.664 33.928 21.232 35.218 ; 
      RECT 20.072 32.836 20.32 35.64 ; 
      RECT 20.016 34.074 20.32 34.688 ; 
      RECT 20.072 31.266 20.176 35.64 ; 
      RECT 20.072 31.75 20.232 32.708 ; 
      RECT 20.072 31.266 20.32 31.622 ; 
      RECT 18.884 33.068 19.708 35.64 ; 
      RECT 19.604 31.266 19.708 35.64 ; 
      RECT 18.884 34.176 19.764 35.208 ; 
      RECT 18.884 31.266 19.276 35.64 ; 
      RECT 17.216 31.266 17.548 35.64 ; 
      RECT 17.216 31.62 17.604 35.362 ; 
      RECT 38.108 31.266 38.448 35.64 ; 
      RECT 37.532 31.266 37.636 35.64 ; 
      RECT 37.1 31.266 37.204 35.64 ; 
      RECT 36.668 31.266 36.772 35.64 ; 
      RECT 36.236 31.266 36.34 35.64 ; 
      RECT 35.804 31.266 35.908 35.64 ; 
      RECT 35.372 31.266 35.476 35.64 ; 
      RECT 34.94 31.266 35.044 35.64 ; 
      RECT 34.508 31.266 34.612 35.64 ; 
      RECT 34.076 31.266 34.18 35.64 ; 
      RECT 33.644 31.266 33.748 35.64 ; 
      RECT 33.212 31.266 33.316 35.64 ; 
      RECT 32.78 31.266 32.884 35.64 ; 
      RECT 32.348 31.266 32.452 35.64 ; 
      RECT 31.916 31.266 32.02 35.64 ; 
      RECT 31.484 31.266 31.588 35.64 ; 
      RECT 31.052 31.266 31.156 35.64 ; 
      RECT 30.62 31.266 30.724 35.64 ; 
      RECT 30.188 31.266 30.292 35.64 ; 
      RECT 29.756 31.266 29.86 35.64 ; 
      RECT 29.324 31.266 29.428 35.64 ; 
      RECT 28.892 31.266 28.996 35.64 ; 
      RECT 28.46 31.266 28.564 35.64 ; 
      RECT 28.028 31.266 28.132 35.64 ; 
      RECT 27.596 31.266 27.7 35.64 ; 
      RECT 27.164 31.266 27.268 35.64 ; 
      RECT 26.732 31.266 26.836 35.64 ; 
      RECT 26.3 31.266 26.404 35.64 ; 
      RECT 25.868 31.266 25.972 35.64 ; 
      RECT 25.436 31.266 25.54 35.64 ; 
      RECT 25.004 31.266 25.108 35.64 ; 
      RECT 24.572 31.266 24.676 35.64 ; 
      RECT 24.14 31.266 24.244 35.64 ; 
      RECT 23.708 31.266 23.812 35.64 ; 
      RECT 22.856 31.266 23.164 35.64 ; 
      RECT 15.284 31.266 15.592 35.64 ; 
      RECT 14.636 31.266 14.74 35.64 ; 
      RECT 14.204 31.266 14.308 35.64 ; 
      RECT 13.772 31.266 13.876 35.64 ; 
      RECT 13.34 31.266 13.444 35.64 ; 
      RECT 12.908 31.266 13.012 35.64 ; 
      RECT 12.476 31.266 12.58 35.64 ; 
      RECT 12.044 31.266 12.148 35.64 ; 
      RECT 11.612 31.266 11.716 35.64 ; 
      RECT 11.18 31.266 11.284 35.64 ; 
      RECT 10.748 31.266 10.852 35.64 ; 
      RECT 10.316 31.266 10.42 35.64 ; 
      RECT 9.884 31.266 9.988 35.64 ; 
      RECT 9.452 31.266 9.556 35.64 ; 
      RECT 9.02 31.266 9.124 35.64 ; 
      RECT 8.588 31.266 8.692 35.64 ; 
      RECT 8.156 31.266 8.26 35.64 ; 
      RECT 7.724 31.266 7.828 35.64 ; 
      RECT 7.292 31.266 7.396 35.64 ; 
      RECT 6.86 31.266 6.964 35.64 ; 
      RECT 6.428 31.266 6.532 35.64 ; 
      RECT 5.996 31.266 6.1 35.64 ; 
      RECT 5.564 31.266 5.668 35.64 ; 
      RECT 5.132 31.266 5.236 35.64 ; 
      RECT 4.7 31.266 4.804 35.64 ; 
      RECT 4.268 31.266 4.372 35.64 ; 
      RECT 3.836 31.266 3.94 35.64 ; 
      RECT 3.404 31.266 3.508 35.64 ; 
      RECT 2.972 31.266 3.076 35.64 ; 
      RECT 2.54 31.266 2.644 35.64 ; 
      RECT 2.108 31.266 2.212 35.64 ; 
      RECT 1.676 31.266 1.78 35.64 ; 
      RECT 1.244 31.266 1.348 35.64 ; 
      RECT 0.812 31.266 0.916 35.64 ; 
      RECT 0 31.266 0.34 35.64 ; 
      RECT 20.72 35.586 21.232 39.96 ; 
      RECT 20.664 38.248 21.232 39.538 ; 
      RECT 20.072 37.156 20.32 39.96 ; 
      RECT 20.016 38.394 20.32 39.008 ; 
      RECT 20.072 35.586 20.176 39.96 ; 
      RECT 20.072 36.07 20.232 37.028 ; 
      RECT 20.072 35.586 20.32 35.942 ; 
      RECT 18.884 37.388 19.708 39.96 ; 
      RECT 19.604 35.586 19.708 39.96 ; 
      RECT 18.884 38.496 19.764 39.528 ; 
      RECT 18.884 35.586 19.276 39.96 ; 
      RECT 17.216 35.586 17.548 39.96 ; 
      RECT 17.216 35.94 17.604 39.682 ; 
      RECT 38.108 35.586 38.448 39.96 ; 
      RECT 37.532 35.586 37.636 39.96 ; 
      RECT 37.1 35.586 37.204 39.96 ; 
      RECT 36.668 35.586 36.772 39.96 ; 
      RECT 36.236 35.586 36.34 39.96 ; 
      RECT 35.804 35.586 35.908 39.96 ; 
      RECT 35.372 35.586 35.476 39.96 ; 
      RECT 34.94 35.586 35.044 39.96 ; 
      RECT 34.508 35.586 34.612 39.96 ; 
      RECT 34.076 35.586 34.18 39.96 ; 
      RECT 33.644 35.586 33.748 39.96 ; 
      RECT 33.212 35.586 33.316 39.96 ; 
      RECT 32.78 35.586 32.884 39.96 ; 
      RECT 32.348 35.586 32.452 39.96 ; 
      RECT 31.916 35.586 32.02 39.96 ; 
      RECT 31.484 35.586 31.588 39.96 ; 
      RECT 31.052 35.586 31.156 39.96 ; 
      RECT 30.62 35.586 30.724 39.96 ; 
      RECT 30.188 35.586 30.292 39.96 ; 
      RECT 29.756 35.586 29.86 39.96 ; 
      RECT 29.324 35.586 29.428 39.96 ; 
      RECT 28.892 35.586 28.996 39.96 ; 
      RECT 28.46 35.586 28.564 39.96 ; 
      RECT 28.028 35.586 28.132 39.96 ; 
      RECT 27.596 35.586 27.7 39.96 ; 
      RECT 27.164 35.586 27.268 39.96 ; 
      RECT 26.732 35.586 26.836 39.96 ; 
      RECT 26.3 35.586 26.404 39.96 ; 
      RECT 25.868 35.586 25.972 39.96 ; 
      RECT 25.436 35.586 25.54 39.96 ; 
      RECT 25.004 35.586 25.108 39.96 ; 
      RECT 24.572 35.586 24.676 39.96 ; 
      RECT 24.14 35.586 24.244 39.96 ; 
      RECT 23.708 35.586 23.812 39.96 ; 
      RECT 22.856 35.586 23.164 39.96 ; 
      RECT 15.284 35.586 15.592 39.96 ; 
      RECT 14.636 35.586 14.74 39.96 ; 
      RECT 14.204 35.586 14.308 39.96 ; 
      RECT 13.772 35.586 13.876 39.96 ; 
      RECT 13.34 35.586 13.444 39.96 ; 
      RECT 12.908 35.586 13.012 39.96 ; 
      RECT 12.476 35.586 12.58 39.96 ; 
      RECT 12.044 35.586 12.148 39.96 ; 
      RECT 11.612 35.586 11.716 39.96 ; 
      RECT 11.18 35.586 11.284 39.96 ; 
      RECT 10.748 35.586 10.852 39.96 ; 
      RECT 10.316 35.586 10.42 39.96 ; 
      RECT 9.884 35.586 9.988 39.96 ; 
      RECT 9.452 35.586 9.556 39.96 ; 
      RECT 9.02 35.586 9.124 39.96 ; 
      RECT 8.588 35.586 8.692 39.96 ; 
      RECT 8.156 35.586 8.26 39.96 ; 
      RECT 7.724 35.586 7.828 39.96 ; 
      RECT 7.292 35.586 7.396 39.96 ; 
      RECT 6.86 35.586 6.964 39.96 ; 
      RECT 6.428 35.586 6.532 39.96 ; 
      RECT 5.996 35.586 6.1 39.96 ; 
      RECT 5.564 35.586 5.668 39.96 ; 
      RECT 5.132 35.586 5.236 39.96 ; 
      RECT 4.7 35.586 4.804 39.96 ; 
      RECT 4.268 35.586 4.372 39.96 ; 
      RECT 3.836 35.586 3.94 39.96 ; 
      RECT 3.404 35.586 3.508 39.96 ; 
      RECT 2.972 35.586 3.076 39.96 ; 
      RECT 2.54 35.586 2.644 39.96 ; 
      RECT 2.108 35.586 2.212 39.96 ; 
      RECT 1.676 35.586 1.78 39.96 ; 
      RECT 1.244 35.586 1.348 39.96 ; 
      RECT 0.812 35.586 0.916 39.96 ; 
      RECT 0 35.586 0.34 39.96 ; 
      RECT 20.72 39.906 21.232 44.28 ; 
      RECT 20.664 42.568 21.232 43.858 ; 
      RECT 20.072 41.476 20.32 44.28 ; 
      RECT 20.016 42.714 20.32 43.328 ; 
      RECT 20.072 39.906 20.176 44.28 ; 
      RECT 20.072 40.39 20.232 41.348 ; 
      RECT 20.072 39.906 20.32 40.262 ; 
      RECT 18.884 41.708 19.708 44.28 ; 
      RECT 19.604 39.906 19.708 44.28 ; 
      RECT 18.884 42.816 19.764 43.848 ; 
      RECT 18.884 39.906 19.276 44.28 ; 
      RECT 17.216 39.906 17.548 44.28 ; 
      RECT 17.216 40.26 17.604 44.002 ; 
      RECT 38.108 39.906 38.448 44.28 ; 
      RECT 37.532 39.906 37.636 44.28 ; 
      RECT 37.1 39.906 37.204 44.28 ; 
      RECT 36.668 39.906 36.772 44.28 ; 
      RECT 36.236 39.906 36.34 44.28 ; 
      RECT 35.804 39.906 35.908 44.28 ; 
      RECT 35.372 39.906 35.476 44.28 ; 
      RECT 34.94 39.906 35.044 44.28 ; 
      RECT 34.508 39.906 34.612 44.28 ; 
      RECT 34.076 39.906 34.18 44.28 ; 
      RECT 33.644 39.906 33.748 44.28 ; 
      RECT 33.212 39.906 33.316 44.28 ; 
      RECT 32.78 39.906 32.884 44.28 ; 
      RECT 32.348 39.906 32.452 44.28 ; 
      RECT 31.916 39.906 32.02 44.28 ; 
      RECT 31.484 39.906 31.588 44.28 ; 
      RECT 31.052 39.906 31.156 44.28 ; 
      RECT 30.62 39.906 30.724 44.28 ; 
      RECT 30.188 39.906 30.292 44.28 ; 
      RECT 29.756 39.906 29.86 44.28 ; 
      RECT 29.324 39.906 29.428 44.28 ; 
      RECT 28.892 39.906 28.996 44.28 ; 
      RECT 28.46 39.906 28.564 44.28 ; 
      RECT 28.028 39.906 28.132 44.28 ; 
      RECT 27.596 39.906 27.7 44.28 ; 
      RECT 27.164 39.906 27.268 44.28 ; 
      RECT 26.732 39.906 26.836 44.28 ; 
      RECT 26.3 39.906 26.404 44.28 ; 
      RECT 25.868 39.906 25.972 44.28 ; 
      RECT 25.436 39.906 25.54 44.28 ; 
      RECT 25.004 39.906 25.108 44.28 ; 
      RECT 24.572 39.906 24.676 44.28 ; 
      RECT 24.14 39.906 24.244 44.28 ; 
      RECT 23.708 39.906 23.812 44.28 ; 
      RECT 22.856 39.906 23.164 44.28 ; 
      RECT 15.284 39.906 15.592 44.28 ; 
      RECT 14.636 39.906 14.74 44.28 ; 
      RECT 14.204 39.906 14.308 44.28 ; 
      RECT 13.772 39.906 13.876 44.28 ; 
      RECT 13.34 39.906 13.444 44.28 ; 
      RECT 12.908 39.906 13.012 44.28 ; 
      RECT 12.476 39.906 12.58 44.28 ; 
      RECT 12.044 39.906 12.148 44.28 ; 
      RECT 11.612 39.906 11.716 44.28 ; 
      RECT 11.18 39.906 11.284 44.28 ; 
      RECT 10.748 39.906 10.852 44.28 ; 
      RECT 10.316 39.906 10.42 44.28 ; 
      RECT 9.884 39.906 9.988 44.28 ; 
      RECT 9.452 39.906 9.556 44.28 ; 
      RECT 9.02 39.906 9.124 44.28 ; 
      RECT 8.588 39.906 8.692 44.28 ; 
      RECT 8.156 39.906 8.26 44.28 ; 
      RECT 7.724 39.906 7.828 44.28 ; 
      RECT 7.292 39.906 7.396 44.28 ; 
      RECT 6.86 39.906 6.964 44.28 ; 
      RECT 6.428 39.906 6.532 44.28 ; 
      RECT 5.996 39.906 6.1 44.28 ; 
      RECT 5.564 39.906 5.668 44.28 ; 
      RECT 5.132 39.906 5.236 44.28 ; 
      RECT 4.7 39.906 4.804 44.28 ; 
      RECT 4.268 39.906 4.372 44.28 ; 
      RECT 3.836 39.906 3.94 44.28 ; 
      RECT 3.404 39.906 3.508 44.28 ; 
      RECT 2.972 39.906 3.076 44.28 ; 
      RECT 2.54 39.906 2.644 44.28 ; 
      RECT 2.108 39.906 2.212 44.28 ; 
      RECT 1.676 39.906 1.78 44.28 ; 
      RECT 1.244 39.906 1.348 44.28 ; 
      RECT 0.812 39.906 0.916 44.28 ; 
      RECT 0 39.906 0.34 44.28 ; 
      RECT 20.72 44.226 21.232 48.6 ; 
      RECT 20.664 46.888 21.232 48.178 ; 
      RECT 20.072 45.796 20.32 48.6 ; 
      RECT 20.016 47.034 20.32 47.648 ; 
      RECT 20.072 44.226 20.176 48.6 ; 
      RECT 20.072 44.71 20.232 45.668 ; 
      RECT 20.072 44.226 20.32 44.582 ; 
      RECT 18.884 46.028 19.708 48.6 ; 
      RECT 19.604 44.226 19.708 48.6 ; 
      RECT 18.884 47.136 19.764 48.168 ; 
      RECT 18.884 44.226 19.276 48.6 ; 
      RECT 17.216 44.226 17.548 48.6 ; 
      RECT 17.216 44.58 17.604 48.322 ; 
      RECT 38.108 44.226 38.448 48.6 ; 
      RECT 37.532 44.226 37.636 48.6 ; 
      RECT 37.1 44.226 37.204 48.6 ; 
      RECT 36.668 44.226 36.772 48.6 ; 
      RECT 36.236 44.226 36.34 48.6 ; 
      RECT 35.804 44.226 35.908 48.6 ; 
      RECT 35.372 44.226 35.476 48.6 ; 
      RECT 34.94 44.226 35.044 48.6 ; 
      RECT 34.508 44.226 34.612 48.6 ; 
      RECT 34.076 44.226 34.18 48.6 ; 
      RECT 33.644 44.226 33.748 48.6 ; 
      RECT 33.212 44.226 33.316 48.6 ; 
      RECT 32.78 44.226 32.884 48.6 ; 
      RECT 32.348 44.226 32.452 48.6 ; 
      RECT 31.916 44.226 32.02 48.6 ; 
      RECT 31.484 44.226 31.588 48.6 ; 
      RECT 31.052 44.226 31.156 48.6 ; 
      RECT 30.62 44.226 30.724 48.6 ; 
      RECT 30.188 44.226 30.292 48.6 ; 
      RECT 29.756 44.226 29.86 48.6 ; 
      RECT 29.324 44.226 29.428 48.6 ; 
      RECT 28.892 44.226 28.996 48.6 ; 
      RECT 28.46 44.226 28.564 48.6 ; 
      RECT 28.028 44.226 28.132 48.6 ; 
      RECT 27.596 44.226 27.7 48.6 ; 
      RECT 27.164 44.226 27.268 48.6 ; 
      RECT 26.732 44.226 26.836 48.6 ; 
      RECT 26.3 44.226 26.404 48.6 ; 
      RECT 25.868 44.226 25.972 48.6 ; 
      RECT 25.436 44.226 25.54 48.6 ; 
      RECT 25.004 44.226 25.108 48.6 ; 
      RECT 24.572 44.226 24.676 48.6 ; 
      RECT 24.14 44.226 24.244 48.6 ; 
      RECT 23.708 44.226 23.812 48.6 ; 
      RECT 22.856 44.226 23.164 48.6 ; 
      RECT 15.284 44.226 15.592 48.6 ; 
      RECT 14.636 44.226 14.74 48.6 ; 
      RECT 14.204 44.226 14.308 48.6 ; 
      RECT 13.772 44.226 13.876 48.6 ; 
      RECT 13.34 44.226 13.444 48.6 ; 
      RECT 12.908 44.226 13.012 48.6 ; 
      RECT 12.476 44.226 12.58 48.6 ; 
      RECT 12.044 44.226 12.148 48.6 ; 
      RECT 11.612 44.226 11.716 48.6 ; 
      RECT 11.18 44.226 11.284 48.6 ; 
      RECT 10.748 44.226 10.852 48.6 ; 
      RECT 10.316 44.226 10.42 48.6 ; 
      RECT 9.884 44.226 9.988 48.6 ; 
      RECT 9.452 44.226 9.556 48.6 ; 
      RECT 9.02 44.226 9.124 48.6 ; 
      RECT 8.588 44.226 8.692 48.6 ; 
      RECT 8.156 44.226 8.26 48.6 ; 
      RECT 7.724 44.226 7.828 48.6 ; 
      RECT 7.292 44.226 7.396 48.6 ; 
      RECT 6.86 44.226 6.964 48.6 ; 
      RECT 6.428 44.226 6.532 48.6 ; 
      RECT 5.996 44.226 6.1 48.6 ; 
      RECT 5.564 44.226 5.668 48.6 ; 
      RECT 5.132 44.226 5.236 48.6 ; 
      RECT 4.7 44.226 4.804 48.6 ; 
      RECT 4.268 44.226 4.372 48.6 ; 
      RECT 3.836 44.226 3.94 48.6 ; 
      RECT 3.404 44.226 3.508 48.6 ; 
      RECT 2.972 44.226 3.076 48.6 ; 
      RECT 2.54 44.226 2.644 48.6 ; 
      RECT 2.108 44.226 2.212 48.6 ; 
      RECT 1.676 44.226 1.78 48.6 ; 
      RECT 1.244 44.226 1.348 48.6 ; 
      RECT 0.812 44.226 0.916 48.6 ; 
      RECT 0 44.226 0.34 48.6 ; 
      RECT 20.72 48.546 21.232 52.92 ; 
      RECT 20.664 51.208 21.232 52.498 ; 
      RECT 20.072 50.116 20.32 52.92 ; 
      RECT 20.016 51.354 20.32 51.968 ; 
      RECT 20.072 48.546 20.176 52.92 ; 
      RECT 20.072 49.03 20.232 49.988 ; 
      RECT 20.072 48.546 20.32 48.902 ; 
      RECT 18.884 50.348 19.708 52.92 ; 
      RECT 19.604 48.546 19.708 52.92 ; 
      RECT 18.884 51.456 19.764 52.488 ; 
      RECT 18.884 48.546 19.276 52.92 ; 
      RECT 17.216 48.546 17.548 52.92 ; 
      RECT 17.216 48.9 17.604 52.642 ; 
      RECT 38.108 48.546 38.448 52.92 ; 
      RECT 37.532 48.546 37.636 52.92 ; 
      RECT 37.1 48.546 37.204 52.92 ; 
      RECT 36.668 48.546 36.772 52.92 ; 
      RECT 36.236 48.546 36.34 52.92 ; 
      RECT 35.804 48.546 35.908 52.92 ; 
      RECT 35.372 48.546 35.476 52.92 ; 
      RECT 34.94 48.546 35.044 52.92 ; 
      RECT 34.508 48.546 34.612 52.92 ; 
      RECT 34.076 48.546 34.18 52.92 ; 
      RECT 33.644 48.546 33.748 52.92 ; 
      RECT 33.212 48.546 33.316 52.92 ; 
      RECT 32.78 48.546 32.884 52.92 ; 
      RECT 32.348 48.546 32.452 52.92 ; 
      RECT 31.916 48.546 32.02 52.92 ; 
      RECT 31.484 48.546 31.588 52.92 ; 
      RECT 31.052 48.546 31.156 52.92 ; 
      RECT 30.62 48.546 30.724 52.92 ; 
      RECT 30.188 48.546 30.292 52.92 ; 
      RECT 29.756 48.546 29.86 52.92 ; 
      RECT 29.324 48.546 29.428 52.92 ; 
      RECT 28.892 48.546 28.996 52.92 ; 
      RECT 28.46 48.546 28.564 52.92 ; 
      RECT 28.028 48.546 28.132 52.92 ; 
      RECT 27.596 48.546 27.7 52.92 ; 
      RECT 27.164 48.546 27.268 52.92 ; 
      RECT 26.732 48.546 26.836 52.92 ; 
      RECT 26.3 48.546 26.404 52.92 ; 
      RECT 25.868 48.546 25.972 52.92 ; 
      RECT 25.436 48.546 25.54 52.92 ; 
      RECT 25.004 48.546 25.108 52.92 ; 
      RECT 24.572 48.546 24.676 52.92 ; 
      RECT 24.14 48.546 24.244 52.92 ; 
      RECT 23.708 48.546 23.812 52.92 ; 
      RECT 22.856 48.546 23.164 52.92 ; 
      RECT 15.284 48.546 15.592 52.92 ; 
      RECT 14.636 48.546 14.74 52.92 ; 
      RECT 14.204 48.546 14.308 52.92 ; 
      RECT 13.772 48.546 13.876 52.92 ; 
      RECT 13.34 48.546 13.444 52.92 ; 
      RECT 12.908 48.546 13.012 52.92 ; 
      RECT 12.476 48.546 12.58 52.92 ; 
      RECT 12.044 48.546 12.148 52.92 ; 
      RECT 11.612 48.546 11.716 52.92 ; 
      RECT 11.18 48.546 11.284 52.92 ; 
      RECT 10.748 48.546 10.852 52.92 ; 
      RECT 10.316 48.546 10.42 52.92 ; 
      RECT 9.884 48.546 9.988 52.92 ; 
      RECT 9.452 48.546 9.556 52.92 ; 
      RECT 9.02 48.546 9.124 52.92 ; 
      RECT 8.588 48.546 8.692 52.92 ; 
      RECT 8.156 48.546 8.26 52.92 ; 
      RECT 7.724 48.546 7.828 52.92 ; 
      RECT 7.292 48.546 7.396 52.92 ; 
      RECT 6.86 48.546 6.964 52.92 ; 
      RECT 6.428 48.546 6.532 52.92 ; 
      RECT 5.996 48.546 6.1 52.92 ; 
      RECT 5.564 48.546 5.668 52.92 ; 
      RECT 5.132 48.546 5.236 52.92 ; 
      RECT 4.7 48.546 4.804 52.92 ; 
      RECT 4.268 48.546 4.372 52.92 ; 
      RECT 3.836 48.546 3.94 52.92 ; 
      RECT 3.404 48.546 3.508 52.92 ; 
      RECT 2.972 48.546 3.076 52.92 ; 
      RECT 2.54 48.546 2.644 52.92 ; 
      RECT 2.108 48.546 2.212 52.92 ; 
      RECT 1.676 48.546 1.78 52.92 ; 
      RECT 1.244 48.546 1.348 52.92 ; 
      RECT 0.812 48.546 0.916 52.92 ; 
      RECT 0 48.546 0.34 52.92 ; 
      RECT 20.72 52.866 21.232 57.24 ; 
      RECT 20.664 55.528 21.232 56.818 ; 
      RECT 20.072 54.436 20.32 57.24 ; 
      RECT 20.016 55.674 20.32 56.288 ; 
      RECT 20.072 52.866 20.176 57.24 ; 
      RECT 20.072 53.35 20.232 54.308 ; 
      RECT 20.072 52.866 20.32 53.222 ; 
      RECT 18.884 54.668 19.708 57.24 ; 
      RECT 19.604 52.866 19.708 57.24 ; 
      RECT 18.884 55.776 19.764 56.808 ; 
      RECT 18.884 52.866 19.276 57.24 ; 
      RECT 17.216 52.866 17.548 57.24 ; 
      RECT 17.216 53.22 17.604 56.962 ; 
      RECT 38.108 52.866 38.448 57.24 ; 
      RECT 37.532 52.866 37.636 57.24 ; 
      RECT 37.1 52.866 37.204 57.24 ; 
      RECT 36.668 52.866 36.772 57.24 ; 
      RECT 36.236 52.866 36.34 57.24 ; 
      RECT 35.804 52.866 35.908 57.24 ; 
      RECT 35.372 52.866 35.476 57.24 ; 
      RECT 34.94 52.866 35.044 57.24 ; 
      RECT 34.508 52.866 34.612 57.24 ; 
      RECT 34.076 52.866 34.18 57.24 ; 
      RECT 33.644 52.866 33.748 57.24 ; 
      RECT 33.212 52.866 33.316 57.24 ; 
      RECT 32.78 52.866 32.884 57.24 ; 
      RECT 32.348 52.866 32.452 57.24 ; 
      RECT 31.916 52.866 32.02 57.24 ; 
      RECT 31.484 52.866 31.588 57.24 ; 
      RECT 31.052 52.866 31.156 57.24 ; 
      RECT 30.62 52.866 30.724 57.24 ; 
      RECT 30.188 52.866 30.292 57.24 ; 
      RECT 29.756 52.866 29.86 57.24 ; 
      RECT 29.324 52.866 29.428 57.24 ; 
      RECT 28.892 52.866 28.996 57.24 ; 
      RECT 28.46 52.866 28.564 57.24 ; 
      RECT 28.028 52.866 28.132 57.24 ; 
      RECT 27.596 52.866 27.7 57.24 ; 
      RECT 27.164 52.866 27.268 57.24 ; 
      RECT 26.732 52.866 26.836 57.24 ; 
      RECT 26.3 52.866 26.404 57.24 ; 
      RECT 25.868 52.866 25.972 57.24 ; 
      RECT 25.436 52.866 25.54 57.24 ; 
      RECT 25.004 52.866 25.108 57.24 ; 
      RECT 24.572 52.866 24.676 57.24 ; 
      RECT 24.14 52.866 24.244 57.24 ; 
      RECT 23.708 52.866 23.812 57.24 ; 
      RECT 22.856 52.866 23.164 57.24 ; 
      RECT 15.284 52.866 15.592 57.24 ; 
      RECT 14.636 52.866 14.74 57.24 ; 
      RECT 14.204 52.866 14.308 57.24 ; 
      RECT 13.772 52.866 13.876 57.24 ; 
      RECT 13.34 52.866 13.444 57.24 ; 
      RECT 12.908 52.866 13.012 57.24 ; 
      RECT 12.476 52.866 12.58 57.24 ; 
      RECT 12.044 52.866 12.148 57.24 ; 
      RECT 11.612 52.866 11.716 57.24 ; 
      RECT 11.18 52.866 11.284 57.24 ; 
      RECT 10.748 52.866 10.852 57.24 ; 
      RECT 10.316 52.866 10.42 57.24 ; 
      RECT 9.884 52.866 9.988 57.24 ; 
      RECT 9.452 52.866 9.556 57.24 ; 
      RECT 9.02 52.866 9.124 57.24 ; 
      RECT 8.588 52.866 8.692 57.24 ; 
      RECT 8.156 52.866 8.26 57.24 ; 
      RECT 7.724 52.866 7.828 57.24 ; 
      RECT 7.292 52.866 7.396 57.24 ; 
      RECT 6.86 52.866 6.964 57.24 ; 
      RECT 6.428 52.866 6.532 57.24 ; 
      RECT 5.996 52.866 6.1 57.24 ; 
      RECT 5.564 52.866 5.668 57.24 ; 
      RECT 5.132 52.866 5.236 57.24 ; 
      RECT 4.7 52.866 4.804 57.24 ; 
      RECT 4.268 52.866 4.372 57.24 ; 
      RECT 3.836 52.866 3.94 57.24 ; 
      RECT 3.404 52.866 3.508 57.24 ; 
      RECT 2.972 52.866 3.076 57.24 ; 
      RECT 2.54 52.866 2.644 57.24 ; 
      RECT 2.108 52.866 2.212 57.24 ; 
      RECT 1.676 52.866 1.78 57.24 ; 
      RECT 1.244 52.866 1.348 57.24 ; 
      RECT 0.812 52.866 0.916 57.24 ; 
      RECT 0 52.866 0.34 57.24 ; 
      RECT 20.72 57.186 21.232 61.56 ; 
      RECT 20.664 59.848 21.232 61.138 ; 
      RECT 20.072 58.756 20.32 61.56 ; 
      RECT 20.016 59.994 20.32 60.608 ; 
      RECT 20.072 57.186 20.176 61.56 ; 
      RECT 20.072 57.67 20.232 58.628 ; 
      RECT 20.072 57.186 20.32 57.542 ; 
      RECT 18.884 58.988 19.708 61.56 ; 
      RECT 19.604 57.186 19.708 61.56 ; 
      RECT 18.884 60.096 19.764 61.128 ; 
      RECT 18.884 57.186 19.276 61.56 ; 
      RECT 17.216 57.186 17.548 61.56 ; 
      RECT 17.216 57.54 17.604 61.282 ; 
      RECT 38.108 57.186 38.448 61.56 ; 
      RECT 37.532 57.186 37.636 61.56 ; 
      RECT 37.1 57.186 37.204 61.56 ; 
      RECT 36.668 57.186 36.772 61.56 ; 
      RECT 36.236 57.186 36.34 61.56 ; 
      RECT 35.804 57.186 35.908 61.56 ; 
      RECT 35.372 57.186 35.476 61.56 ; 
      RECT 34.94 57.186 35.044 61.56 ; 
      RECT 34.508 57.186 34.612 61.56 ; 
      RECT 34.076 57.186 34.18 61.56 ; 
      RECT 33.644 57.186 33.748 61.56 ; 
      RECT 33.212 57.186 33.316 61.56 ; 
      RECT 32.78 57.186 32.884 61.56 ; 
      RECT 32.348 57.186 32.452 61.56 ; 
      RECT 31.916 57.186 32.02 61.56 ; 
      RECT 31.484 57.186 31.588 61.56 ; 
      RECT 31.052 57.186 31.156 61.56 ; 
      RECT 30.62 57.186 30.724 61.56 ; 
      RECT 30.188 57.186 30.292 61.56 ; 
      RECT 29.756 57.186 29.86 61.56 ; 
      RECT 29.324 57.186 29.428 61.56 ; 
      RECT 28.892 57.186 28.996 61.56 ; 
      RECT 28.46 57.186 28.564 61.56 ; 
      RECT 28.028 57.186 28.132 61.56 ; 
      RECT 27.596 57.186 27.7 61.56 ; 
      RECT 27.164 57.186 27.268 61.56 ; 
      RECT 26.732 57.186 26.836 61.56 ; 
      RECT 26.3 57.186 26.404 61.56 ; 
      RECT 25.868 57.186 25.972 61.56 ; 
      RECT 25.436 57.186 25.54 61.56 ; 
      RECT 25.004 57.186 25.108 61.56 ; 
      RECT 24.572 57.186 24.676 61.56 ; 
      RECT 24.14 57.186 24.244 61.56 ; 
      RECT 23.708 57.186 23.812 61.56 ; 
      RECT 22.856 57.186 23.164 61.56 ; 
      RECT 15.284 57.186 15.592 61.56 ; 
      RECT 14.636 57.186 14.74 61.56 ; 
      RECT 14.204 57.186 14.308 61.56 ; 
      RECT 13.772 57.186 13.876 61.56 ; 
      RECT 13.34 57.186 13.444 61.56 ; 
      RECT 12.908 57.186 13.012 61.56 ; 
      RECT 12.476 57.186 12.58 61.56 ; 
      RECT 12.044 57.186 12.148 61.56 ; 
      RECT 11.612 57.186 11.716 61.56 ; 
      RECT 11.18 57.186 11.284 61.56 ; 
      RECT 10.748 57.186 10.852 61.56 ; 
      RECT 10.316 57.186 10.42 61.56 ; 
      RECT 9.884 57.186 9.988 61.56 ; 
      RECT 9.452 57.186 9.556 61.56 ; 
      RECT 9.02 57.186 9.124 61.56 ; 
      RECT 8.588 57.186 8.692 61.56 ; 
      RECT 8.156 57.186 8.26 61.56 ; 
      RECT 7.724 57.186 7.828 61.56 ; 
      RECT 7.292 57.186 7.396 61.56 ; 
      RECT 6.86 57.186 6.964 61.56 ; 
      RECT 6.428 57.186 6.532 61.56 ; 
      RECT 5.996 57.186 6.1 61.56 ; 
      RECT 5.564 57.186 5.668 61.56 ; 
      RECT 5.132 57.186 5.236 61.56 ; 
      RECT 4.7 57.186 4.804 61.56 ; 
      RECT 4.268 57.186 4.372 61.56 ; 
      RECT 3.836 57.186 3.94 61.56 ; 
      RECT 3.404 57.186 3.508 61.56 ; 
      RECT 2.972 57.186 3.076 61.56 ; 
      RECT 2.54 57.186 2.644 61.56 ; 
      RECT 2.108 57.186 2.212 61.56 ; 
      RECT 1.676 57.186 1.78 61.56 ; 
      RECT 1.244 57.186 1.348 61.56 ; 
      RECT 0.812 57.186 0.916 61.56 ; 
      RECT 0 57.186 0.34 61.56 ; 
      RECT 20.72 61.506 21.232 65.88 ; 
      RECT 20.664 64.168 21.232 65.458 ; 
      RECT 20.072 63.076 20.32 65.88 ; 
      RECT 20.016 64.314 20.32 64.928 ; 
      RECT 20.072 61.506 20.176 65.88 ; 
      RECT 20.072 61.99 20.232 62.948 ; 
      RECT 20.072 61.506 20.32 61.862 ; 
      RECT 18.884 63.308 19.708 65.88 ; 
      RECT 19.604 61.506 19.708 65.88 ; 
      RECT 18.884 64.416 19.764 65.448 ; 
      RECT 18.884 61.506 19.276 65.88 ; 
      RECT 17.216 61.506 17.548 65.88 ; 
      RECT 17.216 61.86 17.604 65.602 ; 
      RECT 38.108 61.506 38.448 65.88 ; 
      RECT 37.532 61.506 37.636 65.88 ; 
      RECT 37.1 61.506 37.204 65.88 ; 
      RECT 36.668 61.506 36.772 65.88 ; 
      RECT 36.236 61.506 36.34 65.88 ; 
      RECT 35.804 61.506 35.908 65.88 ; 
      RECT 35.372 61.506 35.476 65.88 ; 
      RECT 34.94 61.506 35.044 65.88 ; 
      RECT 34.508 61.506 34.612 65.88 ; 
      RECT 34.076 61.506 34.18 65.88 ; 
      RECT 33.644 61.506 33.748 65.88 ; 
      RECT 33.212 61.506 33.316 65.88 ; 
      RECT 32.78 61.506 32.884 65.88 ; 
      RECT 32.348 61.506 32.452 65.88 ; 
      RECT 31.916 61.506 32.02 65.88 ; 
      RECT 31.484 61.506 31.588 65.88 ; 
      RECT 31.052 61.506 31.156 65.88 ; 
      RECT 30.62 61.506 30.724 65.88 ; 
      RECT 30.188 61.506 30.292 65.88 ; 
      RECT 29.756 61.506 29.86 65.88 ; 
      RECT 29.324 61.506 29.428 65.88 ; 
      RECT 28.892 61.506 28.996 65.88 ; 
      RECT 28.46 61.506 28.564 65.88 ; 
      RECT 28.028 61.506 28.132 65.88 ; 
      RECT 27.596 61.506 27.7 65.88 ; 
      RECT 27.164 61.506 27.268 65.88 ; 
      RECT 26.732 61.506 26.836 65.88 ; 
      RECT 26.3 61.506 26.404 65.88 ; 
      RECT 25.868 61.506 25.972 65.88 ; 
      RECT 25.436 61.506 25.54 65.88 ; 
      RECT 25.004 61.506 25.108 65.88 ; 
      RECT 24.572 61.506 24.676 65.88 ; 
      RECT 24.14 61.506 24.244 65.88 ; 
      RECT 23.708 61.506 23.812 65.88 ; 
      RECT 22.856 61.506 23.164 65.88 ; 
      RECT 15.284 61.506 15.592 65.88 ; 
      RECT 14.636 61.506 14.74 65.88 ; 
      RECT 14.204 61.506 14.308 65.88 ; 
      RECT 13.772 61.506 13.876 65.88 ; 
      RECT 13.34 61.506 13.444 65.88 ; 
      RECT 12.908 61.506 13.012 65.88 ; 
      RECT 12.476 61.506 12.58 65.88 ; 
      RECT 12.044 61.506 12.148 65.88 ; 
      RECT 11.612 61.506 11.716 65.88 ; 
      RECT 11.18 61.506 11.284 65.88 ; 
      RECT 10.748 61.506 10.852 65.88 ; 
      RECT 10.316 61.506 10.42 65.88 ; 
      RECT 9.884 61.506 9.988 65.88 ; 
      RECT 9.452 61.506 9.556 65.88 ; 
      RECT 9.02 61.506 9.124 65.88 ; 
      RECT 8.588 61.506 8.692 65.88 ; 
      RECT 8.156 61.506 8.26 65.88 ; 
      RECT 7.724 61.506 7.828 65.88 ; 
      RECT 7.292 61.506 7.396 65.88 ; 
      RECT 6.86 61.506 6.964 65.88 ; 
      RECT 6.428 61.506 6.532 65.88 ; 
      RECT 5.996 61.506 6.1 65.88 ; 
      RECT 5.564 61.506 5.668 65.88 ; 
      RECT 5.132 61.506 5.236 65.88 ; 
      RECT 4.7 61.506 4.804 65.88 ; 
      RECT 4.268 61.506 4.372 65.88 ; 
      RECT 3.836 61.506 3.94 65.88 ; 
      RECT 3.404 61.506 3.508 65.88 ; 
      RECT 2.972 61.506 3.076 65.88 ; 
      RECT 2.54 61.506 2.644 65.88 ; 
      RECT 2.108 61.506 2.212 65.88 ; 
      RECT 1.676 61.506 1.78 65.88 ; 
      RECT 1.244 61.506 1.348 65.88 ; 
      RECT 0.812 61.506 0.916 65.88 ; 
      RECT 0 61.506 0.34 65.88 ; 
      RECT 20.72 65.826 21.232 70.2 ; 
      RECT 20.664 68.488 21.232 69.778 ; 
      RECT 20.072 67.396 20.32 70.2 ; 
      RECT 20.016 68.634 20.32 69.248 ; 
      RECT 20.072 65.826 20.176 70.2 ; 
      RECT 20.072 66.31 20.232 67.268 ; 
      RECT 20.072 65.826 20.32 66.182 ; 
      RECT 18.884 67.628 19.708 70.2 ; 
      RECT 19.604 65.826 19.708 70.2 ; 
      RECT 18.884 68.736 19.764 69.768 ; 
      RECT 18.884 65.826 19.276 70.2 ; 
      RECT 17.216 65.826 17.548 70.2 ; 
      RECT 17.216 66.18 17.604 69.922 ; 
      RECT 38.108 65.826 38.448 70.2 ; 
      RECT 37.532 65.826 37.636 70.2 ; 
      RECT 37.1 65.826 37.204 70.2 ; 
      RECT 36.668 65.826 36.772 70.2 ; 
      RECT 36.236 65.826 36.34 70.2 ; 
      RECT 35.804 65.826 35.908 70.2 ; 
      RECT 35.372 65.826 35.476 70.2 ; 
      RECT 34.94 65.826 35.044 70.2 ; 
      RECT 34.508 65.826 34.612 70.2 ; 
      RECT 34.076 65.826 34.18 70.2 ; 
      RECT 33.644 65.826 33.748 70.2 ; 
      RECT 33.212 65.826 33.316 70.2 ; 
      RECT 32.78 65.826 32.884 70.2 ; 
      RECT 32.348 65.826 32.452 70.2 ; 
      RECT 31.916 65.826 32.02 70.2 ; 
      RECT 31.484 65.826 31.588 70.2 ; 
      RECT 31.052 65.826 31.156 70.2 ; 
      RECT 30.62 65.826 30.724 70.2 ; 
      RECT 30.188 65.826 30.292 70.2 ; 
      RECT 29.756 65.826 29.86 70.2 ; 
      RECT 29.324 65.826 29.428 70.2 ; 
      RECT 28.892 65.826 28.996 70.2 ; 
      RECT 28.46 65.826 28.564 70.2 ; 
      RECT 28.028 65.826 28.132 70.2 ; 
      RECT 27.596 65.826 27.7 70.2 ; 
      RECT 27.164 65.826 27.268 70.2 ; 
      RECT 26.732 65.826 26.836 70.2 ; 
      RECT 26.3 65.826 26.404 70.2 ; 
      RECT 25.868 65.826 25.972 70.2 ; 
      RECT 25.436 65.826 25.54 70.2 ; 
      RECT 25.004 65.826 25.108 70.2 ; 
      RECT 24.572 65.826 24.676 70.2 ; 
      RECT 24.14 65.826 24.244 70.2 ; 
      RECT 23.708 65.826 23.812 70.2 ; 
      RECT 22.856 65.826 23.164 70.2 ; 
      RECT 15.284 65.826 15.592 70.2 ; 
      RECT 14.636 65.826 14.74 70.2 ; 
      RECT 14.204 65.826 14.308 70.2 ; 
      RECT 13.772 65.826 13.876 70.2 ; 
      RECT 13.34 65.826 13.444 70.2 ; 
      RECT 12.908 65.826 13.012 70.2 ; 
      RECT 12.476 65.826 12.58 70.2 ; 
      RECT 12.044 65.826 12.148 70.2 ; 
      RECT 11.612 65.826 11.716 70.2 ; 
      RECT 11.18 65.826 11.284 70.2 ; 
      RECT 10.748 65.826 10.852 70.2 ; 
      RECT 10.316 65.826 10.42 70.2 ; 
      RECT 9.884 65.826 9.988 70.2 ; 
      RECT 9.452 65.826 9.556 70.2 ; 
      RECT 9.02 65.826 9.124 70.2 ; 
      RECT 8.588 65.826 8.692 70.2 ; 
      RECT 8.156 65.826 8.26 70.2 ; 
      RECT 7.724 65.826 7.828 70.2 ; 
      RECT 7.292 65.826 7.396 70.2 ; 
      RECT 6.86 65.826 6.964 70.2 ; 
      RECT 6.428 65.826 6.532 70.2 ; 
      RECT 5.996 65.826 6.1 70.2 ; 
      RECT 5.564 65.826 5.668 70.2 ; 
      RECT 5.132 65.826 5.236 70.2 ; 
      RECT 4.7 65.826 4.804 70.2 ; 
      RECT 4.268 65.826 4.372 70.2 ; 
      RECT 3.836 65.826 3.94 70.2 ; 
      RECT 3.404 65.826 3.508 70.2 ; 
      RECT 2.972 65.826 3.076 70.2 ; 
      RECT 2.54 65.826 2.644 70.2 ; 
      RECT 2.108 65.826 2.212 70.2 ; 
      RECT 1.676 65.826 1.78 70.2 ; 
      RECT 1.244 65.826 1.348 70.2 ; 
      RECT 0.812 65.826 0.916 70.2 ; 
      RECT 0 65.826 0.34 70.2 ; 
      RECT 20.72 70.146 21.232 74.52 ; 
      RECT 20.664 72.808 21.232 74.098 ; 
      RECT 20.072 71.716 20.32 74.52 ; 
      RECT 20.016 72.954 20.32 73.568 ; 
      RECT 20.072 70.146 20.176 74.52 ; 
      RECT 20.072 70.63 20.232 71.588 ; 
      RECT 20.072 70.146 20.32 70.502 ; 
      RECT 18.884 71.948 19.708 74.52 ; 
      RECT 19.604 70.146 19.708 74.52 ; 
      RECT 18.884 73.056 19.764 74.088 ; 
      RECT 18.884 70.146 19.276 74.52 ; 
      RECT 17.216 70.146 17.548 74.52 ; 
      RECT 17.216 70.5 17.604 74.242 ; 
      RECT 38.108 70.146 38.448 74.52 ; 
      RECT 37.532 70.146 37.636 74.52 ; 
      RECT 37.1 70.146 37.204 74.52 ; 
      RECT 36.668 70.146 36.772 74.52 ; 
      RECT 36.236 70.146 36.34 74.52 ; 
      RECT 35.804 70.146 35.908 74.52 ; 
      RECT 35.372 70.146 35.476 74.52 ; 
      RECT 34.94 70.146 35.044 74.52 ; 
      RECT 34.508 70.146 34.612 74.52 ; 
      RECT 34.076 70.146 34.18 74.52 ; 
      RECT 33.644 70.146 33.748 74.52 ; 
      RECT 33.212 70.146 33.316 74.52 ; 
      RECT 32.78 70.146 32.884 74.52 ; 
      RECT 32.348 70.146 32.452 74.52 ; 
      RECT 31.916 70.146 32.02 74.52 ; 
      RECT 31.484 70.146 31.588 74.52 ; 
      RECT 31.052 70.146 31.156 74.52 ; 
      RECT 30.62 70.146 30.724 74.52 ; 
      RECT 30.188 70.146 30.292 74.52 ; 
      RECT 29.756 70.146 29.86 74.52 ; 
      RECT 29.324 70.146 29.428 74.52 ; 
      RECT 28.892 70.146 28.996 74.52 ; 
      RECT 28.46 70.146 28.564 74.52 ; 
      RECT 28.028 70.146 28.132 74.52 ; 
      RECT 27.596 70.146 27.7 74.52 ; 
      RECT 27.164 70.146 27.268 74.52 ; 
      RECT 26.732 70.146 26.836 74.52 ; 
      RECT 26.3 70.146 26.404 74.52 ; 
      RECT 25.868 70.146 25.972 74.52 ; 
      RECT 25.436 70.146 25.54 74.52 ; 
      RECT 25.004 70.146 25.108 74.52 ; 
      RECT 24.572 70.146 24.676 74.52 ; 
      RECT 24.14 70.146 24.244 74.52 ; 
      RECT 23.708 70.146 23.812 74.52 ; 
      RECT 22.856 70.146 23.164 74.52 ; 
      RECT 15.284 70.146 15.592 74.52 ; 
      RECT 14.636 70.146 14.74 74.52 ; 
      RECT 14.204 70.146 14.308 74.52 ; 
      RECT 13.772 70.146 13.876 74.52 ; 
      RECT 13.34 70.146 13.444 74.52 ; 
      RECT 12.908 70.146 13.012 74.52 ; 
      RECT 12.476 70.146 12.58 74.52 ; 
      RECT 12.044 70.146 12.148 74.52 ; 
      RECT 11.612 70.146 11.716 74.52 ; 
      RECT 11.18 70.146 11.284 74.52 ; 
      RECT 10.748 70.146 10.852 74.52 ; 
      RECT 10.316 70.146 10.42 74.52 ; 
      RECT 9.884 70.146 9.988 74.52 ; 
      RECT 9.452 70.146 9.556 74.52 ; 
      RECT 9.02 70.146 9.124 74.52 ; 
      RECT 8.588 70.146 8.692 74.52 ; 
      RECT 8.156 70.146 8.26 74.52 ; 
      RECT 7.724 70.146 7.828 74.52 ; 
      RECT 7.292 70.146 7.396 74.52 ; 
      RECT 6.86 70.146 6.964 74.52 ; 
      RECT 6.428 70.146 6.532 74.52 ; 
      RECT 5.996 70.146 6.1 74.52 ; 
      RECT 5.564 70.146 5.668 74.52 ; 
      RECT 5.132 70.146 5.236 74.52 ; 
      RECT 4.7 70.146 4.804 74.52 ; 
      RECT 4.268 70.146 4.372 74.52 ; 
      RECT 3.836 70.146 3.94 74.52 ; 
      RECT 3.404 70.146 3.508 74.52 ; 
      RECT 2.972 70.146 3.076 74.52 ; 
      RECT 2.54 70.146 2.644 74.52 ; 
      RECT 2.108 70.146 2.212 74.52 ; 
      RECT 1.676 70.146 1.78 74.52 ; 
      RECT 1.244 70.146 1.348 74.52 ; 
      RECT 0.812 70.146 0.916 74.52 ; 
      RECT 0 70.146 0.34 74.52 ; 
      RECT 0 107.856 38.448 109.026 ; 
      RECT 38.108 74.412 38.448 109.026 ; 
      RECT 18.164 107.262 38.448 109.026 ; 
      RECT 0 107.262 17.548 109.026 ; 
      RECT 23.708 80.428 37.636 109.026 ; 
      RECT 29.54 74.412 37.636 109.026 ; 
      RECT 18.164 107.156 23.38 109.026 ; 
      RECT 20.72 107.152 23.38 109.026 ; 
      RECT 15.068 80.86 17.548 109.026 ; 
      RECT 15.284 77.476 17.548 109.026 ; 
      RECT 0.812 79.648 14.74 109.026 ; 
      RECT 13.556 74.412 14.74 109.026 ; 
      RECT 0 74.412 0.34 109.026 ; 
      RECT 18.164 107.144 20.32 109.026 ; 
      RECT 20.072 106.06 20.32 109.026 ; 
      RECT 20.72 106.06 23.164 109.026 ; 
      RECT 18.164 106.06 19.708 109.026 ; 
      RECT 23.652 89.584 37.636 107.024 ; 
      RECT 0.812 89.584 14.796 107.024 ; 
      RECT 23.652 89.584 37.692 107.006 ; 
      RECT 0.756 89.584 14.796 107.006 ; 
      RECT 20.756 77.476 23.164 109.026 ; 
      RECT 18.884 77.152 19.564 109.026 ; 
      RECT 19.316 74.412 19.564 109.026 ; 
      RECT 16.148 76.748 17.692 105.46 ; 
      RECT 15.068 105.292 17.748 105.44 ; 
      RECT 20.7 100.996 23.164 105.428 ; 
      RECT 18.828 104.236 19.564 105.14 ; 
      RECT 18.884 101.932 19.62 102.98 ; 
      RECT 15.068 101.14 17.748 102.98 ; 
      RECT 18.828 98.98 19.564 100.82 ; 
      RECT 20.7 90.844 23.164 100.172 ; 
      RECT 15.068 93.436 17.748 98.012 ; 
      RECT 18.884 92.356 19.62 97.58 ; 
      RECT 18.828 94.66 19.62 96.5 ; 
      RECT 18.828 81.7 19.564 94.34 ; 
      RECT 18.828 81.7 19.62 92.18 ; 
      RECT 15.068 91.276 17.748 92.18 ; 
      RECT 20.9 75.118 23.38 89.456 ; 
      RECT 20.7 79.54 23.38 86.684 ; 
      RECT 15.068 83.428 17.748 84.908 ; 
      RECT 18.884 80.62 19.62 81.38 ; 
      RECT 15.284 80.476 17.748 81.236 ; 
      RECT 18.828 80.044 19.564 80.588 ; 
      RECT 18.884 79.54 19.62 80.444 ; 
      RECT 24.356 79.66 37.636 109.026 ; 
      RECT 28.676 79.648 37.636 109.026 ; 
      RECT 23.708 74.412 24.028 109.026 ; 
      RECT 15.068 77.152 15.82 80.408 ; 
      RECT 23.708 74.412 24.892 80.024 ; 
      RECT 23.708 78.88 28.348 80.024 ; 
      RECT 28.676 74.412 29.212 109.026 ; 
      RECT 10.1 78.124 13.228 109.026 ; 
      RECT 0.812 74.412 9.772 109.026 ; 
      RECT 23.708 78.88 29.212 79.256 ; 
      RECT 27.812 74.412 37.636 79.244 ; 
      RECT 12.692 74.412 14.74 79.244 ; 
      RECT 18.828 78.964 19.62 79.22 ; 
      RECT 18.828 78.46 19.564 79.22 ; 
      RECT 26.948 77.344 37.636 79.244 ; 
      RECT 23.708 77.476 26.62 80.024 ; 
      RECT 18.884 77.38 19.62 78.428 ; 
      RECT 0.812 77.344 12.364 79.244 ; 
      RECT 11.828 74.412 12.364 109.026 ; 
      RECT 26.084 74.412 27.484 77.9 ; 
      RECT 23.708 77.152 25.756 80.024 ; 
      RECT 25.22 74.412 25.756 109.026 ; 
      RECT 10.964 77.152 12.364 109.026 ; 
      RECT 0.812 74.412 10.636 79.244 ; 
      RECT 18.884 74.412 18.988 109.026 ; 
      RECT 15.428 74.412 15.82 109.026 ; 
      RECT 10.964 74.412 11.5 109.026 ; 
      RECT 25.22 74.412 27.484 76.952 ; 
      RECT 20.756 74.412 23.164 76.952 ; 
      RECT 15.428 74.412 17.548 76.952 ; 
      RECT 11.828 74.412 14.74 76.952 ; 
      RECT 25.22 74.412 37.636 76.94 ; 
      RECT 0.812 74.412 11.5 76.94 ; 
      RECT 20.7 76.3 23.38 76.916 ; 
      RECT 15.428 76.3 17.604 76.952 ; 
      RECT 23.708 74.412 37.636 75.884 ; 
      RECT 18.884 74.412 19.564 75.884 ; 
      RECT 15.068 74.412 17.548 75.884 ; 
      RECT 0.812 74.412 14.74 75.884 ; 
      RECT 18.164 74.412 19.564 75.472 ; 
      RECT 20.72 74.412 23.164 75.072 ; 
      RECT 18.164 74.412 19.708 75.072 ; 
      RECT 20.72 74.412 23.38 74.496 ; 
      RECT 25.236 74.306 25.308 109.026 ; 
      RECT 24.804 74.306 24.876 109.026 ; 
      RECT 11.844 74.306 11.916 109.026 ; 
      RECT 11.412 74.306 11.484 109.026 ; 
      RECT 20.072 74.412 20.32 75.072 ; 
        RECT 20.72 106.974 21.232 111.348 ; 
        RECT 20.664 109.636 21.232 110.926 ; 
        RECT 20.072 108.544 20.32 111.348 ; 
        RECT 20.016 109.782 20.32 110.396 ; 
        RECT 20.072 106.974 20.176 111.348 ; 
        RECT 20.072 107.458 20.232 108.416 ; 
        RECT 20.072 106.974 20.32 107.33 ; 
        RECT 18.884 108.776 19.708 111.348 ; 
        RECT 19.604 106.974 19.708 111.348 ; 
        RECT 18.884 109.884 19.764 110.916 ; 
        RECT 18.884 106.974 19.276 111.348 ; 
        RECT 17.216 106.974 17.548 111.348 ; 
        RECT 17.216 107.328 17.604 111.07 ; 
        RECT 38.108 106.974 38.448 111.348 ; 
        RECT 37.532 106.974 37.636 111.348 ; 
        RECT 37.1 106.974 37.204 111.348 ; 
        RECT 36.668 106.974 36.772 111.348 ; 
        RECT 36.236 106.974 36.34 111.348 ; 
        RECT 35.804 106.974 35.908 111.348 ; 
        RECT 35.372 106.974 35.476 111.348 ; 
        RECT 34.94 106.974 35.044 111.348 ; 
        RECT 34.508 106.974 34.612 111.348 ; 
        RECT 34.076 106.974 34.18 111.348 ; 
        RECT 33.644 106.974 33.748 111.348 ; 
        RECT 33.212 106.974 33.316 111.348 ; 
        RECT 32.78 106.974 32.884 111.348 ; 
        RECT 32.348 106.974 32.452 111.348 ; 
        RECT 31.916 106.974 32.02 111.348 ; 
        RECT 31.484 106.974 31.588 111.348 ; 
        RECT 31.052 106.974 31.156 111.348 ; 
        RECT 30.62 106.974 30.724 111.348 ; 
        RECT 30.188 106.974 30.292 111.348 ; 
        RECT 29.756 106.974 29.86 111.348 ; 
        RECT 29.324 106.974 29.428 111.348 ; 
        RECT 28.892 106.974 28.996 111.348 ; 
        RECT 28.46 106.974 28.564 111.348 ; 
        RECT 28.028 106.974 28.132 111.348 ; 
        RECT 27.596 106.974 27.7 111.348 ; 
        RECT 27.164 106.974 27.268 111.348 ; 
        RECT 26.732 106.974 26.836 111.348 ; 
        RECT 26.3 106.974 26.404 111.348 ; 
        RECT 25.868 106.974 25.972 111.348 ; 
        RECT 25.436 106.974 25.54 111.348 ; 
        RECT 25.004 106.974 25.108 111.348 ; 
        RECT 24.572 106.974 24.676 111.348 ; 
        RECT 24.14 106.974 24.244 111.348 ; 
        RECT 23.708 106.974 23.812 111.348 ; 
        RECT 22.856 106.974 23.164 111.348 ; 
        RECT 15.284 106.974 15.592 111.348 ; 
        RECT 14.636 106.974 14.74 111.348 ; 
        RECT 14.204 106.974 14.308 111.348 ; 
        RECT 13.772 106.974 13.876 111.348 ; 
        RECT 13.34 106.974 13.444 111.348 ; 
        RECT 12.908 106.974 13.012 111.348 ; 
        RECT 12.476 106.974 12.58 111.348 ; 
        RECT 12.044 106.974 12.148 111.348 ; 
        RECT 11.612 106.974 11.716 111.348 ; 
        RECT 11.18 106.974 11.284 111.348 ; 
        RECT 10.748 106.974 10.852 111.348 ; 
        RECT 10.316 106.974 10.42 111.348 ; 
        RECT 9.884 106.974 9.988 111.348 ; 
        RECT 9.452 106.974 9.556 111.348 ; 
        RECT 9.02 106.974 9.124 111.348 ; 
        RECT 8.588 106.974 8.692 111.348 ; 
        RECT 8.156 106.974 8.26 111.348 ; 
        RECT 7.724 106.974 7.828 111.348 ; 
        RECT 7.292 106.974 7.396 111.348 ; 
        RECT 6.86 106.974 6.964 111.348 ; 
        RECT 6.428 106.974 6.532 111.348 ; 
        RECT 5.996 106.974 6.1 111.348 ; 
        RECT 5.564 106.974 5.668 111.348 ; 
        RECT 5.132 106.974 5.236 111.348 ; 
        RECT 4.7 106.974 4.804 111.348 ; 
        RECT 4.268 106.974 4.372 111.348 ; 
        RECT 3.836 106.974 3.94 111.348 ; 
        RECT 3.404 106.974 3.508 111.348 ; 
        RECT 2.972 106.974 3.076 111.348 ; 
        RECT 2.54 106.974 2.644 111.348 ; 
        RECT 2.108 106.974 2.212 111.348 ; 
        RECT 1.676 106.974 1.78 111.348 ; 
        RECT 1.244 106.974 1.348 111.348 ; 
        RECT 0.812 106.974 0.916 111.348 ; 
        RECT 0 106.974 0.34 111.348 ; 
        RECT 20.72 111.294 21.232 115.668 ; 
        RECT 20.664 113.956 21.232 115.246 ; 
        RECT 20.072 112.864 20.32 115.668 ; 
        RECT 20.016 114.102 20.32 114.716 ; 
        RECT 20.072 111.294 20.176 115.668 ; 
        RECT 20.072 111.778 20.232 112.736 ; 
        RECT 20.072 111.294 20.32 111.65 ; 
        RECT 18.884 113.096 19.708 115.668 ; 
        RECT 19.604 111.294 19.708 115.668 ; 
        RECT 18.884 114.204 19.764 115.236 ; 
        RECT 18.884 111.294 19.276 115.668 ; 
        RECT 17.216 111.294 17.548 115.668 ; 
        RECT 17.216 111.648 17.604 115.39 ; 
        RECT 38.108 111.294 38.448 115.668 ; 
        RECT 37.532 111.294 37.636 115.668 ; 
        RECT 37.1 111.294 37.204 115.668 ; 
        RECT 36.668 111.294 36.772 115.668 ; 
        RECT 36.236 111.294 36.34 115.668 ; 
        RECT 35.804 111.294 35.908 115.668 ; 
        RECT 35.372 111.294 35.476 115.668 ; 
        RECT 34.94 111.294 35.044 115.668 ; 
        RECT 34.508 111.294 34.612 115.668 ; 
        RECT 34.076 111.294 34.18 115.668 ; 
        RECT 33.644 111.294 33.748 115.668 ; 
        RECT 33.212 111.294 33.316 115.668 ; 
        RECT 32.78 111.294 32.884 115.668 ; 
        RECT 32.348 111.294 32.452 115.668 ; 
        RECT 31.916 111.294 32.02 115.668 ; 
        RECT 31.484 111.294 31.588 115.668 ; 
        RECT 31.052 111.294 31.156 115.668 ; 
        RECT 30.62 111.294 30.724 115.668 ; 
        RECT 30.188 111.294 30.292 115.668 ; 
        RECT 29.756 111.294 29.86 115.668 ; 
        RECT 29.324 111.294 29.428 115.668 ; 
        RECT 28.892 111.294 28.996 115.668 ; 
        RECT 28.46 111.294 28.564 115.668 ; 
        RECT 28.028 111.294 28.132 115.668 ; 
        RECT 27.596 111.294 27.7 115.668 ; 
        RECT 27.164 111.294 27.268 115.668 ; 
        RECT 26.732 111.294 26.836 115.668 ; 
        RECT 26.3 111.294 26.404 115.668 ; 
        RECT 25.868 111.294 25.972 115.668 ; 
        RECT 25.436 111.294 25.54 115.668 ; 
        RECT 25.004 111.294 25.108 115.668 ; 
        RECT 24.572 111.294 24.676 115.668 ; 
        RECT 24.14 111.294 24.244 115.668 ; 
        RECT 23.708 111.294 23.812 115.668 ; 
        RECT 22.856 111.294 23.164 115.668 ; 
        RECT 15.284 111.294 15.592 115.668 ; 
        RECT 14.636 111.294 14.74 115.668 ; 
        RECT 14.204 111.294 14.308 115.668 ; 
        RECT 13.772 111.294 13.876 115.668 ; 
        RECT 13.34 111.294 13.444 115.668 ; 
        RECT 12.908 111.294 13.012 115.668 ; 
        RECT 12.476 111.294 12.58 115.668 ; 
        RECT 12.044 111.294 12.148 115.668 ; 
        RECT 11.612 111.294 11.716 115.668 ; 
        RECT 11.18 111.294 11.284 115.668 ; 
        RECT 10.748 111.294 10.852 115.668 ; 
        RECT 10.316 111.294 10.42 115.668 ; 
        RECT 9.884 111.294 9.988 115.668 ; 
        RECT 9.452 111.294 9.556 115.668 ; 
        RECT 9.02 111.294 9.124 115.668 ; 
        RECT 8.588 111.294 8.692 115.668 ; 
        RECT 8.156 111.294 8.26 115.668 ; 
        RECT 7.724 111.294 7.828 115.668 ; 
        RECT 7.292 111.294 7.396 115.668 ; 
        RECT 6.86 111.294 6.964 115.668 ; 
        RECT 6.428 111.294 6.532 115.668 ; 
        RECT 5.996 111.294 6.1 115.668 ; 
        RECT 5.564 111.294 5.668 115.668 ; 
        RECT 5.132 111.294 5.236 115.668 ; 
        RECT 4.7 111.294 4.804 115.668 ; 
        RECT 4.268 111.294 4.372 115.668 ; 
        RECT 3.836 111.294 3.94 115.668 ; 
        RECT 3.404 111.294 3.508 115.668 ; 
        RECT 2.972 111.294 3.076 115.668 ; 
        RECT 2.54 111.294 2.644 115.668 ; 
        RECT 2.108 111.294 2.212 115.668 ; 
        RECT 1.676 111.294 1.78 115.668 ; 
        RECT 1.244 111.294 1.348 115.668 ; 
        RECT 0.812 111.294 0.916 115.668 ; 
        RECT 0 111.294 0.34 115.668 ; 
        RECT 20.72 115.614 21.232 119.988 ; 
        RECT 20.664 118.276 21.232 119.566 ; 
        RECT 20.072 117.184 20.32 119.988 ; 
        RECT 20.016 118.422 20.32 119.036 ; 
        RECT 20.072 115.614 20.176 119.988 ; 
        RECT 20.072 116.098 20.232 117.056 ; 
        RECT 20.072 115.614 20.32 115.97 ; 
        RECT 18.884 117.416 19.708 119.988 ; 
        RECT 19.604 115.614 19.708 119.988 ; 
        RECT 18.884 118.524 19.764 119.556 ; 
        RECT 18.884 115.614 19.276 119.988 ; 
        RECT 17.216 115.614 17.548 119.988 ; 
        RECT 17.216 115.968 17.604 119.71 ; 
        RECT 38.108 115.614 38.448 119.988 ; 
        RECT 37.532 115.614 37.636 119.988 ; 
        RECT 37.1 115.614 37.204 119.988 ; 
        RECT 36.668 115.614 36.772 119.988 ; 
        RECT 36.236 115.614 36.34 119.988 ; 
        RECT 35.804 115.614 35.908 119.988 ; 
        RECT 35.372 115.614 35.476 119.988 ; 
        RECT 34.94 115.614 35.044 119.988 ; 
        RECT 34.508 115.614 34.612 119.988 ; 
        RECT 34.076 115.614 34.18 119.988 ; 
        RECT 33.644 115.614 33.748 119.988 ; 
        RECT 33.212 115.614 33.316 119.988 ; 
        RECT 32.78 115.614 32.884 119.988 ; 
        RECT 32.348 115.614 32.452 119.988 ; 
        RECT 31.916 115.614 32.02 119.988 ; 
        RECT 31.484 115.614 31.588 119.988 ; 
        RECT 31.052 115.614 31.156 119.988 ; 
        RECT 30.62 115.614 30.724 119.988 ; 
        RECT 30.188 115.614 30.292 119.988 ; 
        RECT 29.756 115.614 29.86 119.988 ; 
        RECT 29.324 115.614 29.428 119.988 ; 
        RECT 28.892 115.614 28.996 119.988 ; 
        RECT 28.46 115.614 28.564 119.988 ; 
        RECT 28.028 115.614 28.132 119.988 ; 
        RECT 27.596 115.614 27.7 119.988 ; 
        RECT 27.164 115.614 27.268 119.988 ; 
        RECT 26.732 115.614 26.836 119.988 ; 
        RECT 26.3 115.614 26.404 119.988 ; 
        RECT 25.868 115.614 25.972 119.988 ; 
        RECT 25.436 115.614 25.54 119.988 ; 
        RECT 25.004 115.614 25.108 119.988 ; 
        RECT 24.572 115.614 24.676 119.988 ; 
        RECT 24.14 115.614 24.244 119.988 ; 
        RECT 23.708 115.614 23.812 119.988 ; 
        RECT 22.856 115.614 23.164 119.988 ; 
        RECT 15.284 115.614 15.592 119.988 ; 
        RECT 14.636 115.614 14.74 119.988 ; 
        RECT 14.204 115.614 14.308 119.988 ; 
        RECT 13.772 115.614 13.876 119.988 ; 
        RECT 13.34 115.614 13.444 119.988 ; 
        RECT 12.908 115.614 13.012 119.988 ; 
        RECT 12.476 115.614 12.58 119.988 ; 
        RECT 12.044 115.614 12.148 119.988 ; 
        RECT 11.612 115.614 11.716 119.988 ; 
        RECT 11.18 115.614 11.284 119.988 ; 
        RECT 10.748 115.614 10.852 119.988 ; 
        RECT 10.316 115.614 10.42 119.988 ; 
        RECT 9.884 115.614 9.988 119.988 ; 
        RECT 9.452 115.614 9.556 119.988 ; 
        RECT 9.02 115.614 9.124 119.988 ; 
        RECT 8.588 115.614 8.692 119.988 ; 
        RECT 8.156 115.614 8.26 119.988 ; 
        RECT 7.724 115.614 7.828 119.988 ; 
        RECT 7.292 115.614 7.396 119.988 ; 
        RECT 6.86 115.614 6.964 119.988 ; 
        RECT 6.428 115.614 6.532 119.988 ; 
        RECT 5.996 115.614 6.1 119.988 ; 
        RECT 5.564 115.614 5.668 119.988 ; 
        RECT 5.132 115.614 5.236 119.988 ; 
        RECT 4.7 115.614 4.804 119.988 ; 
        RECT 4.268 115.614 4.372 119.988 ; 
        RECT 3.836 115.614 3.94 119.988 ; 
        RECT 3.404 115.614 3.508 119.988 ; 
        RECT 2.972 115.614 3.076 119.988 ; 
        RECT 2.54 115.614 2.644 119.988 ; 
        RECT 2.108 115.614 2.212 119.988 ; 
        RECT 1.676 115.614 1.78 119.988 ; 
        RECT 1.244 115.614 1.348 119.988 ; 
        RECT 0.812 115.614 0.916 119.988 ; 
        RECT 0 115.614 0.34 119.988 ; 
        RECT 20.72 119.934 21.232 124.308 ; 
        RECT 20.664 122.596 21.232 123.886 ; 
        RECT 20.072 121.504 20.32 124.308 ; 
        RECT 20.016 122.742 20.32 123.356 ; 
        RECT 20.072 119.934 20.176 124.308 ; 
        RECT 20.072 120.418 20.232 121.376 ; 
        RECT 20.072 119.934 20.32 120.29 ; 
        RECT 18.884 121.736 19.708 124.308 ; 
        RECT 19.604 119.934 19.708 124.308 ; 
        RECT 18.884 122.844 19.764 123.876 ; 
        RECT 18.884 119.934 19.276 124.308 ; 
        RECT 17.216 119.934 17.548 124.308 ; 
        RECT 17.216 120.288 17.604 124.03 ; 
        RECT 38.108 119.934 38.448 124.308 ; 
        RECT 37.532 119.934 37.636 124.308 ; 
        RECT 37.1 119.934 37.204 124.308 ; 
        RECT 36.668 119.934 36.772 124.308 ; 
        RECT 36.236 119.934 36.34 124.308 ; 
        RECT 35.804 119.934 35.908 124.308 ; 
        RECT 35.372 119.934 35.476 124.308 ; 
        RECT 34.94 119.934 35.044 124.308 ; 
        RECT 34.508 119.934 34.612 124.308 ; 
        RECT 34.076 119.934 34.18 124.308 ; 
        RECT 33.644 119.934 33.748 124.308 ; 
        RECT 33.212 119.934 33.316 124.308 ; 
        RECT 32.78 119.934 32.884 124.308 ; 
        RECT 32.348 119.934 32.452 124.308 ; 
        RECT 31.916 119.934 32.02 124.308 ; 
        RECT 31.484 119.934 31.588 124.308 ; 
        RECT 31.052 119.934 31.156 124.308 ; 
        RECT 30.62 119.934 30.724 124.308 ; 
        RECT 30.188 119.934 30.292 124.308 ; 
        RECT 29.756 119.934 29.86 124.308 ; 
        RECT 29.324 119.934 29.428 124.308 ; 
        RECT 28.892 119.934 28.996 124.308 ; 
        RECT 28.46 119.934 28.564 124.308 ; 
        RECT 28.028 119.934 28.132 124.308 ; 
        RECT 27.596 119.934 27.7 124.308 ; 
        RECT 27.164 119.934 27.268 124.308 ; 
        RECT 26.732 119.934 26.836 124.308 ; 
        RECT 26.3 119.934 26.404 124.308 ; 
        RECT 25.868 119.934 25.972 124.308 ; 
        RECT 25.436 119.934 25.54 124.308 ; 
        RECT 25.004 119.934 25.108 124.308 ; 
        RECT 24.572 119.934 24.676 124.308 ; 
        RECT 24.14 119.934 24.244 124.308 ; 
        RECT 23.708 119.934 23.812 124.308 ; 
        RECT 22.856 119.934 23.164 124.308 ; 
        RECT 15.284 119.934 15.592 124.308 ; 
        RECT 14.636 119.934 14.74 124.308 ; 
        RECT 14.204 119.934 14.308 124.308 ; 
        RECT 13.772 119.934 13.876 124.308 ; 
        RECT 13.34 119.934 13.444 124.308 ; 
        RECT 12.908 119.934 13.012 124.308 ; 
        RECT 12.476 119.934 12.58 124.308 ; 
        RECT 12.044 119.934 12.148 124.308 ; 
        RECT 11.612 119.934 11.716 124.308 ; 
        RECT 11.18 119.934 11.284 124.308 ; 
        RECT 10.748 119.934 10.852 124.308 ; 
        RECT 10.316 119.934 10.42 124.308 ; 
        RECT 9.884 119.934 9.988 124.308 ; 
        RECT 9.452 119.934 9.556 124.308 ; 
        RECT 9.02 119.934 9.124 124.308 ; 
        RECT 8.588 119.934 8.692 124.308 ; 
        RECT 8.156 119.934 8.26 124.308 ; 
        RECT 7.724 119.934 7.828 124.308 ; 
        RECT 7.292 119.934 7.396 124.308 ; 
        RECT 6.86 119.934 6.964 124.308 ; 
        RECT 6.428 119.934 6.532 124.308 ; 
        RECT 5.996 119.934 6.1 124.308 ; 
        RECT 5.564 119.934 5.668 124.308 ; 
        RECT 5.132 119.934 5.236 124.308 ; 
        RECT 4.7 119.934 4.804 124.308 ; 
        RECT 4.268 119.934 4.372 124.308 ; 
        RECT 3.836 119.934 3.94 124.308 ; 
        RECT 3.404 119.934 3.508 124.308 ; 
        RECT 2.972 119.934 3.076 124.308 ; 
        RECT 2.54 119.934 2.644 124.308 ; 
        RECT 2.108 119.934 2.212 124.308 ; 
        RECT 1.676 119.934 1.78 124.308 ; 
        RECT 1.244 119.934 1.348 124.308 ; 
        RECT 0.812 119.934 0.916 124.308 ; 
        RECT 0 119.934 0.34 124.308 ; 
        RECT 20.72 124.254 21.232 128.628 ; 
        RECT 20.664 126.916 21.232 128.206 ; 
        RECT 20.072 125.824 20.32 128.628 ; 
        RECT 20.016 127.062 20.32 127.676 ; 
        RECT 20.072 124.254 20.176 128.628 ; 
        RECT 20.072 124.738 20.232 125.696 ; 
        RECT 20.072 124.254 20.32 124.61 ; 
        RECT 18.884 126.056 19.708 128.628 ; 
        RECT 19.604 124.254 19.708 128.628 ; 
        RECT 18.884 127.164 19.764 128.196 ; 
        RECT 18.884 124.254 19.276 128.628 ; 
        RECT 17.216 124.254 17.548 128.628 ; 
        RECT 17.216 124.608 17.604 128.35 ; 
        RECT 38.108 124.254 38.448 128.628 ; 
        RECT 37.532 124.254 37.636 128.628 ; 
        RECT 37.1 124.254 37.204 128.628 ; 
        RECT 36.668 124.254 36.772 128.628 ; 
        RECT 36.236 124.254 36.34 128.628 ; 
        RECT 35.804 124.254 35.908 128.628 ; 
        RECT 35.372 124.254 35.476 128.628 ; 
        RECT 34.94 124.254 35.044 128.628 ; 
        RECT 34.508 124.254 34.612 128.628 ; 
        RECT 34.076 124.254 34.18 128.628 ; 
        RECT 33.644 124.254 33.748 128.628 ; 
        RECT 33.212 124.254 33.316 128.628 ; 
        RECT 32.78 124.254 32.884 128.628 ; 
        RECT 32.348 124.254 32.452 128.628 ; 
        RECT 31.916 124.254 32.02 128.628 ; 
        RECT 31.484 124.254 31.588 128.628 ; 
        RECT 31.052 124.254 31.156 128.628 ; 
        RECT 30.62 124.254 30.724 128.628 ; 
        RECT 30.188 124.254 30.292 128.628 ; 
        RECT 29.756 124.254 29.86 128.628 ; 
        RECT 29.324 124.254 29.428 128.628 ; 
        RECT 28.892 124.254 28.996 128.628 ; 
        RECT 28.46 124.254 28.564 128.628 ; 
        RECT 28.028 124.254 28.132 128.628 ; 
        RECT 27.596 124.254 27.7 128.628 ; 
        RECT 27.164 124.254 27.268 128.628 ; 
        RECT 26.732 124.254 26.836 128.628 ; 
        RECT 26.3 124.254 26.404 128.628 ; 
        RECT 25.868 124.254 25.972 128.628 ; 
        RECT 25.436 124.254 25.54 128.628 ; 
        RECT 25.004 124.254 25.108 128.628 ; 
        RECT 24.572 124.254 24.676 128.628 ; 
        RECT 24.14 124.254 24.244 128.628 ; 
        RECT 23.708 124.254 23.812 128.628 ; 
        RECT 22.856 124.254 23.164 128.628 ; 
        RECT 15.284 124.254 15.592 128.628 ; 
        RECT 14.636 124.254 14.74 128.628 ; 
        RECT 14.204 124.254 14.308 128.628 ; 
        RECT 13.772 124.254 13.876 128.628 ; 
        RECT 13.34 124.254 13.444 128.628 ; 
        RECT 12.908 124.254 13.012 128.628 ; 
        RECT 12.476 124.254 12.58 128.628 ; 
        RECT 12.044 124.254 12.148 128.628 ; 
        RECT 11.612 124.254 11.716 128.628 ; 
        RECT 11.18 124.254 11.284 128.628 ; 
        RECT 10.748 124.254 10.852 128.628 ; 
        RECT 10.316 124.254 10.42 128.628 ; 
        RECT 9.884 124.254 9.988 128.628 ; 
        RECT 9.452 124.254 9.556 128.628 ; 
        RECT 9.02 124.254 9.124 128.628 ; 
        RECT 8.588 124.254 8.692 128.628 ; 
        RECT 8.156 124.254 8.26 128.628 ; 
        RECT 7.724 124.254 7.828 128.628 ; 
        RECT 7.292 124.254 7.396 128.628 ; 
        RECT 6.86 124.254 6.964 128.628 ; 
        RECT 6.428 124.254 6.532 128.628 ; 
        RECT 5.996 124.254 6.1 128.628 ; 
        RECT 5.564 124.254 5.668 128.628 ; 
        RECT 5.132 124.254 5.236 128.628 ; 
        RECT 4.7 124.254 4.804 128.628 ; 
        RECT 4.268 124.254 4.372 128.628 ; 
        RECT 3.836 124.254 3.94 128.628 ; 
        RECT 3.404 124.254 3.508 128.628 ; 
        RECT 2.972 124.254 3.076 128.628 ; 
        RECT 2.54 124.254 2.644 128.628 ; 
        RECT 2.108 124.254 2.212 128.628 ; 
        RECT 1.676 124.254 1.78 128.628 ; 
        RECT 1.244 124.254 1.348 128.628 ; 
        RECT 0.812 124.254 0.916 128.628 ; 
        RECT 0 124.254 0.34 128.628 ; 
        RECT 20.72 128.574 21.232 132.948 ; 
        RECT 20.664 131.236 21.232 132.526 ; 
        RECT 20.072 130.144 20.32 132.948 ; 
        RECT 20.016 131.382 20.32 131.996 ; 
        RECT 20.072 128.574 20.176 132.948 ; 
        RECT 20.072 129.058 20.232 130.016 ; 
        RECT 20.072 128.574 20.32 128.93 ; 
        RECT 18.884 130.376 19.708 132.948 ; 
        RECT 19.604 128.574 19.708 132.948 ; 
        RECT 18.884 131.484 19.764 132.516 ; 
        RECT 18.884 128.574 19.276 132.948 ; 
        RECT 17.216 128.574 17.548 132.948 ; 
        RECT 17.216 128.928 17.604 132.67 ; 
        RECT 38.108 128.574 38.448 132.948 ; 
        RECT 37.532 128.574 37.636 132.948 ; 
        RECT 37.1 128.574 37.204 132.948 ; 
        RECT 36.668 128.574 36.772 132.948 ; 
        RECT 36.236 128.574 36.34 132.948 ; 
        RECT 35.804 128.574 35.908 132.948 ; 
        RECT 35.372 128.574 35.476 132.948 ; 
        RECT 34.94 128.574 35.044 132.948 ; 
        RECT 34.508 128.574 34.612 132.948 ; 
        RECT 34.076 128.574 34.18 132.948 ; 
        RECT 33.644 128.574 33.748 132.948 ; 
        RECT 33.212 128.574 33.316 132.948 ; 
        RECT 32.78 128.574 32.884 132.948 ; 
        RECT 32.348 128.574 32.452 132.948 ; 
        RECT 31.916 128.574 32.02 132.948 ; 
        RECT 31.484 128.574 31.588 132.948 ; 
        RECT 31.052 128.574 31.156 132.948 ; 
        RECT 30.62 128.574 30.724 132.948 ; 
        RECT 30.188 128.574 30.292 132.948 ; 
        RECT 29.756 128.574 29.86 132.948 ; 
        RECT 29.324 128.574 29.428 132.948 ; 
        RECT 28.892 128.574 28.996 132.948 ; 
        RECT 28.46 128.574 28.564 132.948 ; 
        RECT 28.028 128.574 28.132 132.948 ; 
        RECT 27.596 128.574 27.7 132.948 ; 
        RECT 27.164 128.574 27.268 132.948 ; 
        RECT 26.732 128.574 26.836 132.948 ; 
        RECT 26.3 128.574 26.404 132.948 ; 
        RECT 25.868 128.574 25.972 132.948 ; 
        RECT 25.436 128.574 25.54 132.948 ; 
        RECT 25.004 128.574 25.108 132.948 ; 
        RECT 24.572 128.574 24.676 132.948 ; 
        RECT 24.14 128.574 24.244 132.948 ; 
        RECT 23.708 128.574 23.812 132.948 ; 
        RECT 22.856 128.574 23.164 132.948 ; 
        RECT 15.284 128.574 15.592 132.948 ; 
        RECT 14.636 128.574 14.74 132.948 ; 
        RECT 14.204 128.574 14.308 132.948 ; 
        RECT 13.772 128.574 13.876 132.948 ; 
        RECT 13.34 128.574 13.444 132.948 ; 
        RECT 12.908 128.574 13.012 132.948 ; 
        RECT 12.476 128.574 12.58 132.948 ; 
        RECT 12.044 128.574 12.148 132.948 ; 
        RECT 11.612 128.574 11.716 132.948 ; 
        RECT 11.18 128.574 11.284 132.948 ; 
        RECT 10.748 128.574 10.852 132.948 ; 
        RECT 10.316 128.574 10.42 132.948 ; 
        RECT 9.884 128.574 9.988 132.948 ; 
        RECT 9.452 128.574 9.556 132.948 ; 
        RECT 9.02 128.574 9.124 132.948 ; 
        RECT 8.588 128.574 8.692 132.948 ; 
        RECT 8.156 128.574 8.26 132.948 ; 
        RECT 7.724 128.574 7.828 132.948 ; 
        RECT 7.292 128.574 7.396 132.948 ; 
        RECT 6.86 128.574 6.964 132.948 ; 
        RECT 6.428 128.574 6.532 132.948 ; 
        RECT 5.996 128.574 6.1 132.948 ; 
        RECT 5.564 128.574 5.668 132.948 ; 
        RECT 5.132 128.574 5.236 132.948 ; 
        RECT 4.7 128.574 4.804 132.948 ; 
        RECT 4.268 128.574 4.372 132.948 ; 
        RECT 3.836 128.574 3.94 132.948 ; 
        RECT 3.404 128.574 3.508 132.948 ; 
        RECT 2.972 128.574 3.076 132.948 ; 
        RECT 2.54 128.574 2.644 132.948 ; 
        RECT 2.108 128.574 2.212 132.948 ; 
        RECT 1.676 128.574 1.78 132.948 ; 
        RECT 1.244 128.574 1.348 132.948 ; 
        RECT 0.812 128.574 0.916 132.948 ; 
        RECT 0 128.574 0.34 132.948 ; 
        RECT 20.72 132.894 21.232 137.268 ; 
        RECT 20.664 135.556 21.232 136.846 ; 
        RECT 20.072 134.464 20.32 137.268 ; 
        RECT 20.016 135.702 20.32 136.316 ; 
        RECT 20.072 132.894 20.176 137.268 ; 
        RECT 20.072 133.378 20.232 134.336 ; 
        RECT 20.072 132.894 20.32 133.25 ; 
        RECT 18.884 134.696 19.708 137.268 ; 
        RECT 19.604 132.894 19.708 137.268 ; 
        RECT 18.884 135.804 19.764 136.836 ; 
        RECT 18.884 132.894 19.276 137.268 ; 
        RECT 17.216 132.894 17.548 137.268 ; 
        RECT 17.216 133.248 17.604 136.99 ; 
        RECT 38.108 132.894 38.448 137.268 ; 
        RECT 37.532 132.894 37.636 137.268 ; 
        RECT 37.1 132.894 37.204 137.268 ; 
        RECT 36.668 132.894 36.772 137.268 ; 
        RECT 36.236 132.894 36.34 137.268 ; 
        RECT 35.804 132.894 35.908 137.268 ; 
        RECT 35.372 132.894 35.476 137.268 ; 
        RECT 34.94 132.894 35.044 137.268 ; 
        RECT 34.508 132.894 34.612 137.268 ; 
        RECT 34.076 132.894 34.18 137.268 ; 
        RECT 33.644 132.894 33.748 137.268 ; 
        RECT 33.212 132.894 33.316 137.268 ; 
        RECT 32.78 132.894 32.884 137.268 ; 
        RECT 32.348 132.894 32.452 137.268 ; 
        RECT 31.916 132.894 32.02 137.268 ; 
        RECT 31.484 132.894 31.588 137.268 ; 
        RECT 31.052 132.894 31.156 137.268 ; 
        RECT 30.62 132.894 30.724 137.268 ; 
        RECT 30.188 132.894 30.292 137.268 ; 
        RECT 29.756 132.894 29.86 137.268 ; 
        RECT 29.324 132.894 29.428 137.268 ; 
        RECT 28.892 132.894 28.996 137.268 ; 
        RECT 28.46 132.894 28.564 137.268 ; 
        RECT 28.028 132.894 28.132 137.268 ; 
        RECT 27.596 132.894 27.7 137.268 ; 
        RECT 27.164 132.894 27.268 137.268 ; 
        RECT 26.732 132.894 26.836 137.268 ; 
        RECT 26.3 132.894 26.404 137.268 ; 
        RECT 25.868 132.894 25.972 137.268 ; 
        RECT 25.436 132.894 25.54 137.268 ; 
        RECT 25.004 132.894 25.108 137.268 ; 
        RECT 24.572 132.894 24.676 137.268 ; 
        RECT 24.14 132.894 24.244 137.268 ; 
        RECT 23.708 132.894 23.812 137.268 ; 
        RECT 22.856 132.894 23.164 137.268 ; 
        RECT 15.284 132.894 15.592 137.268 ; 
        RECT 14.636 132.894 14.74 137.268 ; 
        RECT 14.204 132.894 14.308 137.268 ; 
        RECT 13.772 132.894 13.876 137.268 ; 
        RECT 13.34 132.894 13.444 137.268 ; 
        RECT 12.908 132.894 13.012 137.268 ; 
        RECT 12.476 132.894 12.58 137.268 ; 
        RECT 12.044 132.894 12.148 137.268 ; 
        RECT 11.612 132.894 11.716 137.268 ; 
        RECT 11.18 132.894 11.284 137.268 ; 
        RECT 10.748 132.894 10.852 137.268 ; 
        RECT 10.316 132.894 10.42 137.268 ; 
        RECT 9.884 132.894 9.988 137.268 ; 
        RECT 9.452 132.894 9.556 137.268 ; 
        RECT 9.02 132.894 9.124 137.268 ; 
        RECT 8.588 132.894 8.692 137.268 ; 
        RECT 8.156 132.894 8.26 137.268 ; 
        RECT 7.724 132.894 7.828 137.268 ; 
        RECT 7.292 132.894 7.396 137.268 ; 
        RECT 6.86 132.894 6.964 137.268 ; 
        RECT 6.428 132.894 6.532 137.268 ; 
        RECT 5.996 132.894 6.1 137.268 ; 
        RECT 5.564 132.894 5.668 137.268 ; 
        RECT 5.132 132.894 5.236 137.268 ; 
        RECT 4.7 132.894 4.804 137.268 ; 
        RECT 4.268 132.894 4.372 137.268 ; 
        RECT 3.836 132.894 3.94 137.268 ; 
        RECT 3.404 132.894 3.508 137.268 ; 
        RECT 2.972 132.894 3.076 137.268 ; 
        RECT 2.54 132.894 2.644 137.268 ; 
        RECT 2.108 132.894 2.212 137.268 ; 
        RECT 1.676 132.894 1.78 137.268 ; 
        RECT 1.244 132.894 1.348 137.268 ; 
        RECT 0.812 132.894 0.916 137.268 ; 
        RECT 0 132.894 0.34 137.268 ; 
        RECT 20.72 137.214 21.232 141.588 ; 
        RECT 20.664 139.876 21.232 141.166 ; 
        RECT 20.072 138.784 20.32 141.588 ; 
        RECT 20.016 140.022 20.32 140.636 ; 
        RECT 20.072 137.214 20.176 141.588 ; 
        RECT 20.072 137.698 20.232 138.656 ; 
        RECT 20.072 137.214 20.32 137.57 ; 
        RECT 18.884 139.016 19.708 141.588 ; 
        RECT 19.604 137.214 19.708 141.588 ; 
        RECT 18.884 140.124 19.764 141.156 ; 
        RECT 18.884 137.214 19.276 141.588 ; 
        RECT 17.216 137.214 17.548 141.588 ; 
        RECT 17.216 137.568 17.604 141.31 ; 
        RECT 38.108 137.214 38.448 141.588 ; 
        RECT 37.532 137.214 37.636 141.588 ; 
        RECT 37.1 137.214 37.204 141.588 ; 
        RECT 36.668 137.214 36.772 141.588 ; 
        RECT 36.236 137.214 36.34 141.588 ; 
        RECT 35.804 137.214 35.908 141.588 ; 
        RECT 35.372 137.214 35.476 141.588 ; 
        RECT 34.94 137.214 35.044 141.588 ; 
        RECT 34.508 137.214 34.612 141.588 ; 
        RECT 34.076 137.214 34.18 141.588 ; 
        RECT 33.644 137.214 33.748 141.588 ; 
        RECT 33.212 137.214 33.316 141.588 ; 
        RECT 32.78 137.214 32.884 141.588 ; 
        RECT 32.348 137.214 32.452 141.588 ; 
        RECT 31.916 137.214 32.02 141.588 ; 
        RECT 31.484 137.214 31.588 141.588 ; 
        RECT 31.052 137.214 31.156 141.588 ; 
        RECT 30.62 137.214 30.724 141.588 ; 
        RECT 30.188 137.214 30.292 141.588 ; 
        RECT 29.756 137.214 29.86 141.588 ; 
        RECT 29.324 137.214 29.428 141.588 ; 
        RECT 28.892 137.214 28.996 141.588 ; 
        RECT 28.46 137.214 28.564 141.588 ; 
        RECT 28.028 137.214 28.132 141.588 ; 
        RECT 27.596 137.214 27.7 141.588 ; 
        RECT 27.164 137.214 27.268 141.588 ; 
        RECT 26.732 137.214 26.836 141.588 ; 
        RECT 26.3 137.214 26.404 141.588 ; 
        RECT 25.868 137.214 25.972 141.588 ; 
        RECT 25.436 137.214 25.54 141.588 ; 
        RECT 25.004 137.214 25.108 141.588 ; 
        RECT 24.572 137.214 24.676 141.588 ; 
        RECT 24.14 137.214 24.244 141.588 ; 
        RECT 23.708 137.214 23.812 141.588 ; 
        RECT 22.856 137.214 23.164 141.588 ; 
        RECT 15.284 137.214 15.592 141.588 ; 
        RECT 14.636 137.214 14.74 141.588 ; 
        RECT 14.204 137.214 14.308 141.588 ; 
        RECT 13.772 137.214 13.876 141.588 ; 
        RECT 13.34 137.214 13.444 141.588 ; 
        RECT 12.908 137.214 13.012 141.588 ; 
        RECT 12.476 137.214 12.58 141.588 ; 
        RECT 12.044 137.214 12.148 141.588 ; 
        RECT 11.612 137.214 11.716 141.588 ; 
        RECT 11.18 137.214 11.284 141.588 ; 
        RECT 10.748 137.214 10.852 141.588 ; 
        RECT 10.316 137.214 10.42 141.588 ; 
        RECT 9.884 137.214 9.988 141.588 ; 
        RECT 9.452 137.214 9.556 141.588 ; 
        RECT 9.02 137.214 9.124 141.588 ; 
        RECT 8.588 137.214 8.692 141.588 ; 
        RECT 8.156 137.214 8.26 141.588 ; 
        RECT 7.724 137.214 7.828 141.588 ; 
        RECT 7.292 137.214 7.396 141.588 ; 
        RECT 6.86 137.214 6.964 141.588 ; 
        RECT 6.428 137.214 6.532 141.588 ; 
        RECT 5.996 137.214 6.1 141.588 ; 
        RECT 5.564 137.214 5.668 141.588 ; 
        RECT 5.132 137.214 5.236 141.588 ; 
        RECT 4.7 137.214 4.804 141.588 ; 
        RECT 4.268 137.214 4.372 141.588 ; 
        RECT 3.836 137.214 3.94 141.588 ; 
        RECT 3.404 137.214 3.508 141.588 ; 
        RECT 2.972 137.214 3.076 141.588 ; 
        RECT 2.54 137.214 2.644 141.588 ; 
        RECT 2.108 137.214 2.212 141.588 ; 
        RECT 1.676 137.214 1.78 141.588 ; 
        RECT 1.244 137.214 1.348 141.588 ; 
        RECT 0.812 137.214 0.916 141.588 ; 
        RECT 0 137.214 0.34 141.588 ; 
        RECT 20.72 141.534 21.232 145.908 ; 
        RECT 20.664 144.196 21.232 145.486 ; 
        RECT 20.072 143.104 20.32 145.908 ; 
        RECT 20.016 144.342 20.32 144.956 ; 
        RECT 20.072 141.534 20.176 145.908 ; 
        RECT 20.072 142.018 20.232 142.976 ; 
        RECT 20.072 141.534 20.32 141.89 ; 
        RECT 18.884 143.336 19.708 145.908 ; 
        RECT 19.604 141.534 19.708 145.908 ; 
        RECT 18.884 144.444 19.764 145.476 ; 
        RECT 18.884 141.534 19.276 145.908 ; 
        RECT 17.216 141.534 17.548 145.908 ; 
        RECT 17.216 141.888 17.604 145.63 ; 
        RECT 38.108 141.534 38.448 145.908 ; 
        RECT 37.532 141.534 37.636 145.908 ; 
        RECT 37.1 141.534 37.204 145.908 ; 
        RECT 36.668 141.534 36.772 145.908 ; 
        RECT 36.236 141.534 36.34 145.908 ; 
        RECT 35.804 141.534 35.908 145.908 ; 
        RECT 35.372 141.534 35.476 145.908 ; 
        RECT 34.94 141.534 35.044 145.908 ; 
        RECT 34.508 141.534 34.612 145.908 ; 
        RECT 34.076 141.534 34.18 145.908 ; 
        RECT 33.644 141.534 33.748 145.908 ; 
        RECT 33.212 141.534 33.316 145.908 ; 
        RECT 32.78 141.534 32.884 145.908 ; 
        RECT 32.348 141.534 32.452 145.908 ; 
        RECT 31.916 141.534 32.02 145.908 ; 
        RECT 31.484 141.534 31.588 145.908 ; 
        RECT 31.052 141.534 31.156 145.908 ; 
        RECT 30.62 141.534 30.724 145.908 ; 
        RECT 30.188 141.534 30.292 145.908 ; 
        RECT 29.756 141.534 29.86 145.908 ; 
        RECT 29.324 141.534 29.428 145.908 ; 
        RECT 28.892 141.534 28.996 145.908 ; 
        RECT 28.46 141.534 28.564 145.908 ; 
        RECT 28.028 141.534 28.132 145.908 ; 
        RECT 27.596 141.534 27.7 145.908 ; 
        RECT 27.164 141.534 27.268 145.908 ; 
        RECT 26.732 141.534 26.836 145.908 ; 
        RECT 26.3 141.534 26.404 145.908 ; 
        RECT 25.868 141.534 25.972 145.908 ; 
        RECT 25.436 141.534 25.54 145.908 ; 
        RECT 25.004 141.534 25.108 145.908 ; 
        RECT 24.572 141.534 24.676 145.908 ; 
        RECT 24.14 141.534 24.244 145.908 ; 
        RECT 23.708 141.534 23.812 145.908 ; 
        RECT 22.856 141.534 23.164 145.908 ; 
        RECT 15.284 141.534 15.592 145.908 ; 
        RECT 14.636 141.534 14.74 145.908 ; 
        RECT 14.204 141.534 14.308 145.908 ; 
        RECT 13.772 141.534 13.876 145.908 ; 
        RECT 13.34 141.534 13.444 145.908 ; 
        RECT 12.908 141.534 13.012 145.908 ; 
        RECT 12.476 141.534 12.58 145.908 ; 
        RECT 12.044 141.534 12.148 145.908 ; 
        RECT 11.612 141.534 11.716 145.908 ; 
        RECT 11.18 141.534 11.284 145.908 ; 
        RECT 10.748 141.534 10.852 145.908 ; 
        RECT 10.316 141.534 10.42 145.908 ; 
        RECT 9.884 141.534 9.988 145.908 ; 
        RECT 9.452 141.534 9.556 145.908 ; 
        RECT 9.02 141.534 9.124 145.908 ; 
        RECT 8.588 141.534 8.692 145.908 ; 
        RECT 8.156 141.534 8.26 145.908 ; 
        RECT 7.724 141.534 7.828 145.908 ; 
        RECT 7.292 141.534 7.396 145.908 ; 
        RECT 6.86 141.534 6.964 145.908 ; 
        RECT 6.428 141.534 6.532 145.908 ; 
        RECT 5.996 141.534 6.1 145.908 ; 
        RECT 5.564 141.534 5.668 145.908 ; 
        RECT 5.132 141.534 5.236 145.908 ; 
        RECT 4.7 141.534 4.804 145.908 ; 
        RECT 4.268 141.534 4.372 145.908 ; 
        RECT 3.836 141.534 3.94 145.908 ; 
        RECT 3.404 141.534 3.508 145.908 ; 
        RECT 2.972 141.534 3.076 145.908 ; 
        RECT 2.54 141.534 2.644 145.908 ; 
        RECT 2.108 141.534 2.212 145.908 ; 
        RECT 1.676 141.534 1.78 145.908 ; 
        RECT 1.244 141.534 1.348 145.908 ; 
        RECT 0.812 141.534 0.916 145.908 ; 
        RECT 0 141.534 0.34 145.908 ; 
        RECT 20.72 145.854 21.232 150.228 ; 
        RECT 20.664 148.516 21.232 149.806 ; 
        RECT 20.072 147.424 20.32 150.228 ; 
        RECT 20.016 148.662 20.32 149.276 ; 
        RECT 20.072 145.854 20.176 150.228 ; 
        RECT 20.072 146.338 20.232 147.296 ; 
        RECT 20.072 145.854 20.32 146.21 ; 
        RECT 18.884 147.656 19.708 150.228 ; 
        RECT 19.604 145.854 19.708 150.228 ; 
        RECT 18.884 148.764 19.764 149.796 ; 
        RECT 18.884 145.854 19.276 150.228 ; 
        RECT 17.216 145.854 17.548 150.228 ; 
        RECT 17.216 146.208 17.604 149.95 ; 
        RECT 38.108 145.854 38.448 150.228 ; 
        RECT 37.532 145.854 37.636 150.228 ; 
        RECT 37.1 145.854 37.204 150.228 ; 
        RECT 36.668 145.854 36.772 150.228 ; 
        RECT 36.236 145.854 36.34 150.228 ; 
        RECT 35.804 145.854 35.908 150.228 ; 
        RECT 35.372 145.854 35.476 150.228 ; 
        RECT 34.94 145.854 35.044 150.228 ; 
        RECT 34.508 145.854 34.612 150.228 ; 
        RECT 34.076 145.854 34.18 150.228 ; 
        RECT 33.644 145.854 33.748 150.228 ; 
        RECT 33.212 145.854 33.316 150.228 ; 
        RECT 32.78 145.854 32.884 150.228 ; 
        RECT 32.348 145.854 32.452 150.228 ; 
        RECT 31.916 145.854 32.02 150.228 ; 
        RECT 31.484 145.854 31.588 150.228 ; 
        RECT 31.052 145.854 31.156 150.228 ; 
        RECT 30.62 145.854 30.724 150.228 ; 
        RECT 30.188 145.854 30.292 150.228 ; 
        RECT 29.756 145.854 29.86 150.228 ; 
        RECT 29.324 145.854 29.428 150.228 ; 
        RECT 28.892 145.854 28.996 150.228 ; 
        RECT 28.46 145.854 28.564 150.228 ; 
        RECT 28.028 145.854 28.132 150.228 ; 
        RECT 27.596 145.854 27.7 150.228 ; 
        RECT 27.164 145.854 27.268 150.228 ; 
        RECT 26.732 145.854 26.836 150.228 ; 
        RECT 26.3 145.854 26.404 150.228 ; 
        RECT 25.868 145.854 25.972 150.228 ; 
        RECT 25.436 145.854 25.54 150.228 ; 
        RECT 25.004 145.854 25.108 150.228 ; 
        RECT 24.572 145.854 24.676 150.228 ; 
        RECT 24.14 145.854 24.244 150.228 ; 
        RECT 23.708 145.854 23.812 150.228 ; 
        RECT 22.856 145.854 23.164 150.228 ; 
        RECT 15.284 145.854 15.592 150.228 ; 
        RECT 14.636 145.854 14.74 150.228 ; 
        RECT 14.204 145.854 14.308 150.228 ; 
        RECT 13.772 145.854 13.876 150.228 ; 
        RECT 13.34 145.854 13.444 150.228 ; 
        RECT 12.908 145.854 13.012 150.228 ; 
        RECT 12.476 145.854 12.58 150.228 ; 
        RECT 12.044 145.854 12.148 150.228 ; 
        RECT 11.612 145.854 11.716 150.228 ; 
        RECT 11.18 145.854 11.284 150.228 ; 
        RECT 10.748 145.854 10.852 150.228 ; 
        RECT 10.316 145.854 10.42 150.228 ; 
        RECT 9.884 145.854 9.988 150.228 ; 
        RECT 9.452 145.854 9.556 150.228 ; 
        RECT 9.02 145.854 9.124 150.228 ; 
        RECT 8.588 145.854 8.692 150.228 ; 
        RECT 8.156 145.854 8.26 150.228 ; 
        RECT 7.724 145.854 7.828 150.228 ; 
        RECT 7.292 145.854 7.396 150.228 ; 
        RECT 6.86 145.854 6.964 150.228 ; 
        RECT 6.428 145.854 6.532 150.228 ; 
        RECT 5.996 145.854 6.1 150.228 ; 
        RECT 5.564 145.854 5.668 150.228 ; 
        RECT 5.132 145.854 5.236 150.228 ; 
        RECT 4.7 145.854 4.804 150.228 ; 
        RECT 4.268 145.854 4.372 150.228 ; 
        RECT 3.836 145.854 3.94 150.228 ; 
        RECT 3.404 145.854 3.508 150.228 ; 
        RECT 2.972 145.854 3.076 150.228 ; 
        RECT 2.54 145.854 2.644 150.228 ; 
        RECT 2.108 145.854 2.212 150.228 ; 
        RECT 1.676 145.854 1.78 150.228 ; 
        RECT 1.244 145.854 1.348 150.228 ; 
        RECT 0.812 145.854 0.916 150.228 ; 
        RECT 0 145.854 0.34 150.228 ; 
        RECT 20.72 150.174 21.232 154.548 ; 
        RECT 20.664 152.836 21.232 154.126 ; 
        RECT 20.072 151.744 20.32 154.548 ; 
        RECT 20.016 152.982 20.32 153.596 ; 
        RECT 20.072 150.174 20.176 154.548 ; 
        RECT 20.072 150.658 20.232 151.616 ; 
        RECT 20.072 150.174 20.32 150.53 ; 
        RECT 18.884 151.976 19.708 154.548 ; 
        RECT 19.604 150.174 19.708 154.548 ; 
        RECT 18.884 153.084 19.764 154.116 ; 
        RECT 18.884 150.174 19.276 154.548 ; 
        RECT 17.216 150.174 17.548 154.548 ; 
        RECT 17.216 150.528 17.604 154.27 ; 
        RECT 38.108 150.174 38.448 154.548 ; 
        RECT 37.532 150.174 37.636 154.548 ; 
        RECT 37.1 150.174 37.204 154.548 ; 
        RECT 36.668 150.174 36.772 154.548 ; 
        RECT 36.236 150.174 36.34 154.548 ; 
        RECT 35.804 150.174 35.908 154.548 ; 
        RECT 35.372 150.174 35.476 154.548 ; 
        RECT 34.94 150.174 35.044 154.548 ; 
        RECT 34.508 150.174 34.612 154.548 ; 
        RECT 34.076 150.174 34.18 154.548 ; 
        RECT 33.644 150.174 33.748 154.548 ; 
        RECT 33.212 150.174 33.316 154.548 ; 
        RECT 32.78 150.174 32.884 154.548 ; 
        RECT 32.348 150.174 32.452 154.548 ; 
        RECT 31.916 150.174 32.02 154.548 ; 
        RECT 31.484 150.174 31.588 154.548 ; 
        RECT 31.052 150.174 31.156 154.548 ; 
        RECT 30.62 150.174 30.724 154.548 ; 
        RECT 30.188 150.174 30.292 154.548 ; 
        RECT 29.756 150.174 29.86 154.548 ; 
        RECT 29.324 150.174 29.428 154.548 ; 
        RECT 28.892 150.174 28.996 154.548 ; 
        RECT 28.46 150.174 28.564 154.548 ; 
        RECT 28.028 150.174 28.132 154.548 ; 
        RECT 27.596 150.174 27.7 154.548 ; 
        RECT 27.164 150.174 27.268 154.548 ; 
        RECT 26.732 150.174 26.836 154.548 ; 
        RECT 26.3 150.174 26.404 154.548 ; 
        RECT 25.868 150.174 25.972 154.548 ; 
        RECT 25.436 150.174 25.54 154.548 ; 
        RECT 25.004 150.174 25.108 154.548 ; 
        RECT 24.572 150.174 24.676 154.548 ; 
        RECT 24.14 150.174 24.244 154.548 ; 
        RECT 23.708 150.174 23.812 154.548 ; 
        RECT 22.856 150.174 23.164 154.548 ; 
        RECT 15.284 150.174 15.592 154.548 ; 
        RECT 14.636 150.174 14.74 154.548 ; 
        RECT 14.204 150.174 14.308 154.548 ; 
        RECT 13.772 150.174 13.876 154.548 ; 
        RECT 13.34 150.174 13.444 154.548 ; 
        RECT 12.908 150.174 13.012 154.548 ; 
        RECT 12.476 150.174 12.58 154.548 ; 
        RECT 12.044 150.174 12.148 154.548 ; 
        RECT 11.612 150.174 11.716 154.548 ; 
        RECT 11.18 150.174 11.284 154.548 ; 
        RECT 10.748 150.174 10.852 154.548 ; 
        RECT 10.316 150.174 10.42 154.548 ; 
        RECT 9.884 150.174 9.988 154.548 ; 
        RECT 9.452 150.174 9.556 154.548 ; 
        RECT 9.02 150.174 9.124 154.548 ; 
        RECT 8.588 150.174 8.692 154.548 ; 
        RECT 8.156 150.174 8.26 154.548 ; 
        RECT 7.724 150.174 7.828 154.548 ; 
        RECT 7.292 150.174 7.396 154.548 ; 
        RECT 6.86 150.174 6.964 154.548 ; 
        RECT 6.428 150.174 6.532 154.548 ; 
        RECT 5.996 150.174 6.1 154.548 ; 
        RECT 5.564 150.174 5.668 154.548 ; 
        RECT 5.132 150.174 5.236 154.548 ; 
        RECT 4.7 150.174 4.804 154.548 ; 
        RECT 4.268 150.174 4.372 154.548 ; 
        RECT 3.836 150.174 3.94 154.548 ; 
        RECT 3.404 150.174 3.508 154.548 ; 
        RECT 2.972 150.174 3.076 154.548 ; 
        RECT 2.54 150.174 2.644 154.548 ; 
        RECT 2.108 150.174 2.212 154.548 ; 
        RECT 1.676 150.174 1.78 154.548 ; 
        RECT 1.244 150.174 1.348 154.548 ; 
        RECT 0.812 150.174 0.916 154.548 ; 
        RECT 0 150.174 0.34 154.548 ; 
        RECT 20.72 154.494 21.232 158.868 ; 
        RECT 20.664 157.156 21.232 158.446 ; 
        RECT 20.072 156.064 20.32 158.868 ; 
        RECT 20.016 157.302 20.32 157.916 ; 
        RECT 20.072 154.494 20.176 158.868 ; 
        RECT 20.072 154.978 20.232 155.936 ; 
        RECT 20.072 154.494 20.32 154.85 ; 
        RECT 18.884 156.296 19.708 158.868 ; 
        RECT 19.604 154.494 19.708 158.868 ; 
        RECT 18.884 157.404 19.764 158.436 ; 
        RECT 18.884 154.494 19.276 158.868 ; 
        RECT 17.216 154.494 17.548 158.868 ; 
        RECT 17.216 154.848 17.604 158.59 ; 
        RECT 38.108 154.494 38.448 158.868 ; 
        RECT 37.532 154.494 37.636 158.868 ; 
        RECT 37.1 154.494 37.204 158.868 ; 
        RECT 36.668 154.494 36.772 158.868 ; 
        RECT 36.236 154.494 36.34 158.868 ; 
        RECT 35.804 154.494 35.908 158.868 ; 
        RECT 35.372 154.494 35.476 158.868 ; 
        RECT 34.94 154.494 35.044 158.868 ; 
        RECT 34.508 154.494 34.612 158.868 ; 
        RECT 34.076 154.494 34.18 158.868 ; 
        RECT 33.644 154.494 33.748 158.868 ; 
        RECT 33.212 154.494 33.316 158.868 ; 
        RECT 32.78 154.494 32.884 158.868 ; 
        RECT 32.348 154.494 32.452 158.868 ; 
        RECT 31.916 154.494 32.02 158.868 ; 
        RECT 31.484 154.494 31.588 158.868 ; 
        RECT 31.052 154.494 31.156 158.868 ; 
        RECT 30.62 154.494 30.724 158.868 ; 
        RECT 30.188 154.494 30.292 158.868 ; 
        RECT 29.756 154.494 29.86 158.868 ; 
        RECT 29.324 154.494 29.428 158.868 ; 
        RECT 28.892 154.494 28.996 158.868 ; 
        RECT 28.46 154.494 28.564 158.868 ; 
        RECT 28.028 154.494 28.132 158.868 ; 
        RECT 27.596 154.494 27.7 158.868 ; 
        RECT 27.164 154.494 27.268 158.868 ; 
        RECT 26.732 154.494 26.836 158.868 ; 
        RECT 26.3 154.494 26.404 158.868 ; 
        RECT 25.868 154.494 25.972 158.868 ; 
        RECT 25.436 154.494 25.54 158.868 ; 
        RECT 25.004 154.494 25.108 158.868 ; 
        RECT 24.572 154.494 24.676 158.868 ; 
        RECT 24.14 154.494 24.244 158.868 ; 
        RECT 23.708 154.494 23.812 158.868 ; 
        RECT 22.856 154.494 23.164 158.868 ; 
        RECT 15.284 154.494 15.592 158.868 ; 
        RECT 14.636 154.494 14.74 158.868 ; 
        RECT 14.204 154.494 14.308 158.868 ; 
        RECT 13.772 154.494 13.876 158.868 ; 
        RECT 13.34 154.494 13.444 158.868 ; 
        RECT 12.908 154.494 13.012 158.868 ; 
        RECT 12.476 154.494 12.58 158.868 ; 
        RECT 12.044 154.494 12.148 158.868 ; 
        RECT 11.612 154.494 11.716 158.868 ; 
        RECT 11.18 154.494 11.284 158.868 ; 
        RECT 10.748 154.494 10.852 158.868 ; 
        RECT 10.316 154.494 10.42 158.868 ; 
        RECT 9.884 154.494 9.988 158.868 ; 
        RECT 9.452 154.494 9.556 158.868 ; 
        RECT 9.02 154.494 9.124 158.868 ; 
        RECT 8.588 154.494 8.692 158.868 ; 
        RECT 8.156 154.494 8.26 158.868 ; 
        RECT 7.724 154.494 7.828 158.868 ; 
        RECT 7.292 154.494 7.396 158.868 ; 
        RECT 6.86 154.494 6.964 158.868 ; 
        RECT 6.428 154.494 6.532 158.868 ; 
        RECT 5.996 154.494 6.1 158.868 ; 
        RECT 5.564 154.494 5.668 158.868 ; 
        RECT 5.132 154.494 5.236 158.868 ; 
        RECT 4.7 154.494 4.804 158.868 ; 
        RECT 4.268 154.494 4.372 158.868 ; 
        RECT 3.836 154.494 3.94 158.868 ; 
        RECT 3.404 154.494 3.508 158.868 ; 
        RECT 2.972 154.494 3.076 158.868 ; 
        RECT 2.54 154.494 2.644 158.868 ; 
        RECT 2.108 154.494 2.212 158.868 ; 
        RECT 1.676 154.494 1.78 158.868 ; 
        RECT 1.244 154.494 1.348 158.868 ; 
        RECT 0.812 154.494 0.916 158.868 ; 
        RECT 0 154.494 0.34 158.868 ; 
        RECT 20.72 158.814 21.232 163.188 ; 
        RECT 20.664 161.476 21.232 162.766 ; 
        RECT 20.072 160.384 20.32 163.188 ; 
        RECT 20.016 161.622 20.32 162.236 ; 
        RECT 20.072 158.814 20.176 163.188 ; 
        RECT 20.072 159.298 20.232 160.256 ; 
        RECT 20.072 158.814 20.32 159.17 ; 
        RECT 18.884 160.616 19.708 163.188 ; 
        RECT 19.604 158.814 19.708 163.188 ; 
        RECT 18.884 161.724 19.764 162.756 ; 
        RECT 18.884 158.814 19.276 163.188 ; 
        RECT 17.216 158.814 17.548 163.188 ; 
        RECT 17.216 159.168 17.604 162.91 ; 
        RECT 38.108 158.814 38.448 163.188 ; 
        RECT 37.532 158.814 37.636 163.188 ; 
        RECT 37.1 158.814 37.204 163.188 ; 
        RECT 36.668 158.814 36.772 163.188 ; 
        RECT 36.236 158.814 36.34 163.188 ; 
        RECT 35.804 158.814 35.908 163.188 ; 
        RECT 35.372 158.814 35.476 163.188 ; 
        RECT 34.94 158.814 35.044 163.188 ; 
        RECT 34.508 158.814 34.612 163.188 ; 
        RECT 34.076 158.814 34.18 163.188 ; 
        RECT 33.644 158.814 33.748 163.188 ; 
        RECT 33.212 158.814 33.316 163.188 ; 
        RECT 32.78 158.814 32.884 163.188 ; 
        RECT 32.348 158.814 32.452 163.188 ; 
        RECT 31.916 158.814 32.02 163.188 ; 
        RECT 31.484 158.814 31.588 163.188 ; 
        RECT 31.052 158.814 31.156 163.188 ; 
        RECT 30.62 158.814 30.724 163.188 ; 
        RECT 30.188 158.814 30.292 163.188 ; 
        RECT 29.756 158.814 29.86 163.188 ; 
        RECT 29.324 158.814 29.428 163.188 ; 
        RECT 28.892 158.814 28.996 163.188 ; 
        RECT 28.46 158.814 28.564 163.188 ; 
        RECT 28.028 158.814 28.132 163.188 ; 
        RECT 27.596 158.814 27.7 163.188 ; 
        RECT 27.164 158.814 27.268 163.188 ; 
        RECT 26.732 158.814 26.836 163.188 ; 
        RECT 26.3 158.814 26.404 163.188 ; 
        RECT 25.868 158.814 25.972 163.188 ; 
        RECT 25.436 158.814 25.54 163.188 ; 
        RECT 25.004 158.814 25.108 163.188 ; 
        RECT 24.572 158.814 24.676 163.188 ; 
        RECT 24.14 158.814 24.244 163.188 ; 
        RECT 23.708 158.814 23.812 163.188 ; 
        RECT 22.856 158.814 23.164 163.188 ; 
        RECT 15.284 158.814 15.592 163.188 ; 
        RECT 14.636 158.814 14.74 163.188 ; 
        RECT 14.204 158.814 14.308 163.188 ; 
        RECT 13.772 158.814 13.876 163.188 ; 
        RECT 13.34 158.814 13.444 163.188 ; 
        RECT 12.908 158.814 13.012 163.188 ; 
        RECT 12.476 158.814 12.58 163.188 ; 
        RECT 12.044 158.814 12.148 163.188 ; 
        RECT 11.612 158.814 11.716 163.188 ; 
        RECT 11.18 158.814 11.284 163.188 ; 
        RECT 10.748 158.814 10.852 163.188 ; 
        RECT 10.316 158.814 10.42 163.188 ; 
        RECT 9.884 158.814 9.988 163.188 ; 
        RECT 9.452 158.814 9.556 163.188 ; 
        RECT 9.02 158.814 9.124 163.188 ; 
        RECT 8.588 158.814 8.692 163.188 ; 
        RECT 8.156 158.814 8.26 163.188 ; 
        RECT 7.724 158.814 7.828 163.188 ; 
        RECT 7.292 158.814 7.396 163.188 ; 
        RECT 6.86 158.814 6.964 163.188 ; 
        RECT 6.428 158.814 6.532 163.188 ; 
        RECT 5.996 158.814 6.1 163.188 ; 
        RECT 5.564 158.814 5.668 163.188 ; 
        RECT 5.132 158.814 5.236 163.188 ; 
        RECT 4.7 158.814 4.804 163.188 ; 
        RECT 4.268 158.814 4.372 163.188 ; 
        RECT 3.836 158.814 3.94 163.188 ; 
        RECT 3.404 158.814 3.508 163.188 ; 
        RECT 2.972 158.814 3.076 163.188 ; 
        RECT 2.54 158.814 2.644 163.188 ; 
        RECT 2.108 158.814 2.212 163.188 ; 
        RECT 1.676 158.814 1.78 163.188 ; 
        RECT 1.244 158.814 1.348 163.188 ; 
        RECT 0.812 158.814 0.916 163.188 ; 
        RECT 0 158.814 0.34 163.188 ; 
        RECT 20.72 163.134 21.232 167.508 ; 
        RECT 20.664 165.796 21.232 167.086 ; 
        RECT 20.072 164.704 20.32 167.508 ; 
        RECT 20.016 165.942 20.32 166.556 ; 
        RECT 20.072 163.134 20.176 167.508 ; 
        RECT 20.072 163.618 20.232 164.576 ; 
        RECT 20.072 163.134 20.32 163.49 ; 
        RECT 18.884 164.936 19.708 167.508 ; 
        RECT 19.604 163.134 19.708 167.508 ; 
        RECT 18.884 166.044 19.764 167.076 ; 
        RECT 18.884 163.134 19.276 167.508 ; 
        RECT 17.216 163.134 17.548 167.508 ; 
        RECT 17.216 163.488 17.604 167.23 ; 
        RECT 38.108 163.134 38.448 167.508 ; 
        RECT 37.532 163.134 37.636 167.508 ; 
        RECT 37.1 163.134 37.204 167.508 ; 
        RECT 36.668 163.134 36.772 167.508 ; 
        RECT 36.236 163.134 36.34 167.508 ; 
        RECT 35.804 163.134 35.908 167.508 ; 
        RECT 35.372 163.134 35.476 167.508 ; 
        RECT 34.94 163.134 35.044 167.508 ; 
        RECT 34.508 163.134 34.612 167.508 ; 
        RECT 34.076 163.134 34.18 167.508 ; 
        RECT 33.644 163.134 33.748 167.508 ; 
        RECT 33.212 163.134 33.316 167.508 ; 
        RECT 32.78 163.134 32.884 167.508 ; 
        RECT 32.348 163.134 32.452 167.508 ; 
        RECT 31.916 163.134 32.02 167.508 ; 
        RECT 31.484 163.134 31.588 167.508 ; 
        RECT 31.052 163.134 31.156 167.508 ; 
        RECT 30.62 163.134 30.724 167.508 ; 
        RECT 30.188 163.134 30.292 167.508 ; 
        RECT 29.756 163.134 29.86 167.508 ; 
        RECT 29.324 163.134 29.428 167.508 ; 
        RECT 28.892 163.134 28.996 167.508 ; 
        RECT 28.46 163.134 28.564 167.508 ; 
        RECT 28.028 163.134 28.132 167.508 ; 
        RECT 27.596 163.134 27.7 167.508 ; 
        RECT 27.164 163.134 27.268 167.508 ; 
        RECT 26.732 163.134 26.836 167.508 ; 
        RECT 26.3 163.134 26.404 167.508 ; 
        RECT 25.868 163.134 25.972 167.508 ; 
        RECT 25.436 163.134 25.54 167.508 ; 
        RECT 25.004 163.134 25.108 167.508 ; 
        RECT 24.572 163.134 24.676 167.508 ; 
        RECT 24.14 163.134 24.244 167.508 ; 
        RECT 23.708 163.134 23.812 167.508 ; 
        RECT 22.856 163.134 23.164 167.508 ; 
        RECT 15.284 163.134 15.592 167.508 ; 
        RECT 14.636 163.134 14.74 167.508 ; 
        RECT 14.204 163.134 14.308 167.508 ; 
        RECT 13.772 163.134 13.876 167.508 ; 
        RECT 13.34 163.134 13.444 167.508 ; 
        RECT 12.908 163.134 13.012 167.508 ; 
        RECT 12.476 163.134 12.58 167.508 ; 
        RECT 12.044 163.134 12.148 167.508 ; 
        RECT 11.612 163.134 11.716 167.508 ; 
        RECT 11.18 163.134 11.284 167.508 ; 
        RECT 10.748 163.134 10.852 167.508 ; 
        RECT 10.316 163.134 10.42 167.508 ; 
        RECT 9.884 163.134 9.988 167.508 ; 
        RECT 9.452 163.134 9.556 167.508 ; 
        RECT 9.02 163.134 9.124 167.508 ; 
        RECT 8.588 163.134 8.692 167.508 ; 
        RECT 8.156 163.134 8.26 167.508 ; 
        RECT 7.724 163.134 7.828 167.508 ; 
        RECT 7.292 163.134 7.396 167.508 ; 
        RECT 6.86 163.134 6.964 167.508 ; 
        RECT 6.428 163.134 6.532 167.508 ; 
        RECT 5.996 163.134 6.1 167.508 ; 
        RECT 5.564 163.134 5.668 167.508 ; 
        RECT 5.132 163.134 5.236 167.508 ; 
        RECT 4.7 163.134 4.804 167.508 ; 
        RECT 4.268 163.134 4.372 167.508 ; 
        RECT 3.836 163.134 3.94 167.508 ; 
        RECT 3.404 163.134 3.508 167.508 ; 
        RECT 2.972 163.134 3.076 167.508 ; 
        RECT 2.54 163.134 2.644 167.508 ; 
        RECT 2.108 163.134 2.212 167.508 ; 
        RECT 1.676 163.134 1.78 167.508 ; 
        RECT 1.244 163.134 1.348 167.508 ; 
        RECT 0.812 163.134 0.916 167.508 ; 
        RECT 0 163.134 0.34 167.508 ; 
        RECT 20.72 167.454 21.232 171.828 ; 
        RECT 20.664 170.116 21.232 171.406 ; 
        RECT 20.072 169.024 20.32 171.828 ; 
        RECT 20.016 170.262 20.32 170.876 ; 
        RECT 20.072 167.454 20.176 171.828 ; 
        RECT 20.072 167.938 20.232 168.896 ; 
        RECT 20.072 167.454 20.32 167.81 ; 
        RECT 18.884 169.256 19.708 171.828 ; 
        RECT 19.604 167.454 19.708 171.828 ; 
        RECT 18.884 170.364 19.764 171.396 ; 
        RECT 18.884 167.454 19.276 171.828 ; 
        RECT 17.216 167.454 17.548 171.828 ; 
        RECT 17.216 167.808 17.604 171.55 ; 
        RECT 38.108 167.454 38.448 171.828 ; 
        RECT 37.532 167.454 37.636 171.828 ; 
        RECT 37.1 167.454 37.204 171.828 ; 
        RECT 36.668 167.454 36.772 171.828 ; 
        RECT 36.236 167.454 36.34 171.828 ; 
        RECT 35.804 167.454 35.908 171.828 ; 
        RECT 35.372 167.454 35.476 171.828 ; 
        RECT 34.94 167.454 35.044 171.828 ; 
        RECT 34.508 167.454 34.612 171.828 ; 
        RECT 34.076 167.454 34.18 171.828 ; 
        RECT 33.644 167.454 33.748 171.828 ; 
        RECT 33.212 167.454 33.316 171.828 ; 
        RECT 32.78 167.454 32.884 171.828 ; 
        RECT 32.348 167.454 32.452 171.828 ; 
        RECT 31.916 167.454 32.02 171.828 ; 
        RECT 31.484 167.454 31.588 171.828 ; 
        RECT 31.052 167.454 31.156 171.828 ; 
        RECT 30.62 167.454 30.724 171.828 ; 
        RECT 30.188 167.454 30.292 171.828 ; 
        RECT 29.756 167.454 29.86 171.828 ; 
        RECT 29.324 167.454 29.428 171.828 ; 
        RECT 28.892 167.454 28.996 171.828 ; 
        RECT 28.46 167.454 28.564 171.828 ; 
        RECT 28.028 167.454 28.132 171.828 ; 
        RECT 27.596 167.454 27.7 171.828 ; 
        RECT 27.164 167.454 27.268 171.828 ; 
        RECT 26.732 167.454 26.836 171.828 ; 
        RECT 26.3 167.454 26.404 171.828 ; 
        RECT 25.868 167.454 25.972 171.828 ; 
        RECT 25.436 167.454 25.54 171.828 ; 
        RECT 25.004 167.454 25.108 171.828 ; 
        RECT 24.572 167.454 24.676 171.828 ; 
        RECT 24.14 167.454 24.244 171.828 ; 
        RECT 23.708 167.454 23.812 171.828 ; 
        RECT 22.856 167.454 23.164 171.828 ; 
        RECT 15.284 167.454 15.592 171.828 ; 
        RECT 14.636 167.454 14.74 171.828 ; 
        RECT 14.204 167.454 14.308 171.828 ; 
        RECT 13.772 167.454 13.876 171.828 ; 
        RECT 13.34 167.454 13.444 171.828 ; 
        RECT 12.908 167.454 13.012 171.828 ; 
        RECT 12.476 167.454 12.58 171.828 ; 
        RECT 12.044 167.454 12.148 171.828 ; 
        RECT 11.612 167.454 11.716 171.828 ; 
        RECT 11.18 167.454 11.284 171.828 ; 
        RECT 10.748 167.454 10.852 171.828 ; 
        RECT 10.316 167.454 10.42 171.828 ; 
        RECT 9.884 167.454 9.988 171.828 ; 
        RECT 9.452 167.454 9.556 171.828 ; 
        RECT 9.02 167.454 9.124 171.828 ; 
        RECT 8.588 167.454 8.692 171.828 ; 
        RECT 8.156 167.454 8.26 171.828 ; 
        RECT 7.724 167.454 7.828 171.828 ; 
        RECT 7.292 167.454 7.396 171.828 ; 
        RECT 6.86 167.454 6.964 171.828 ; 
        RECT 6.428 167.454 6.532 171.828 ; 
        RECT 5.996 167.454 6.1 171.828 ; 
        RECT 5.564 167.454 5.668 171.828 ; 
        RECT 5.132 167.454 5.236 171.828 ; 
        RECT 4.7 167.454 4.804 171.828 ; 
        RECT 4.268 167.454 4.372 171.828 ; 
        RECT 3.836 167.454 3.94 171.828 ; 
        RECT 3.404 167.454 3.508 171.828 ; 
        RECT 2.972 167.454 3.076 171.828 ; 
        RECT 2.54 167.454 2.644 171.828 ; 
        RECT 2.108 167.454 2.212 171.828 ; 
        RECT 1.676 167.454 1.78 171.828 ; 
        RECT 1.244 167.454 1.348 171.828 ; 
        RECT 0.812 167.454 0.916 171.828 ; 
        RECT 0 167.454 0.34 171.828 ; 
        RECT 20.72 171.774 21.232 176.148 ; 
        RECT 20.664 174.436 21.232 175.726 ; 
        RECT 20.072 173.344 20.32 176.148 ; 
        RECT 20.016 174.582 20.32 175.196 ; 
        RECT 20.072 171.774 20.176 176.148 ; 
        RECT 20.072 172.258 20.232 173.216 ; 
        RECT 20.072 171.774 20.32 172.13 ; 
        RECT 18.884 173.576 19.708 176.148 ; 
        RECT 19.604 171.774 19.708 176.148 ; 
        RECT 18.884 174.684 19.764 175.716 ; 
        RECT 18.884 171.774 19.276 176.148 ; 
        RECT 17.216 171.774 17.548 176.148 ; 
        RECT 17.216 172.128 17.604 175.87 ; 
        RECT 38.108 171.774 38.448 176.148 ; 
        RECT 37.532 171.774 37.636 176.148 ; 
        RECT 37.1 171.774 37.204 176.148 ; 
        RECT 36.668 171.774 36.772 176.148 ; 
        RECT 36.236 171.774 36.34 176.148 ; 
        RECT 35.804 171.774 35.908 176.148 ; 
        RECT 35.372 171.774 35.476 176.148 ; 
        RECT 34.94 171.774 35.044 176.148 ; 
        RECT 34.508 171.774 34.612 176.148 ; 
        RECT 34.076 171.774 34.18 176.148 ; 
        RECT 33.644 171.774 33.748 176.148 ; 
        RECT 33.212 171.774 33.316 176.148 ; 
        RECT 32.78 171.774 32.884 176.148 ; 
        RECT 32.348 171.774 32.452 176.148 ; 
        RECT 31.916 171.774 32.02 176.148 ; 
        RECT 31.484 171.774 31.588 176.148 ; 
        RECT 31.052 171.774 31.156 176.148 ; 
        RECT 30.62 171.774 30.724 176.148 ; 
        RECT 30.188 171.774 30.292 176.148 ; 
        RECT 29.756 171.774 29.86 176.148 ; 
        RECT 29.324 171.774 29.428 176.148 ; 
        RECT 28.892 171.774 28.996 176.148 ; 
        RECT 28.46 171.774 28.564 176.148 ; 
        RECT 28.028 171.774 28.132 176.148 ; 
        RECT 27.596 171.774 27.7 176.148 ; 
        RECT 27.164 171.774 27.268 176.148 ; 
        RECT 26.732 171.774 26.836 176.148 ; 
        RECT 26.3 171.774 26.404 176.148 ; 
        RECT 25.868 171.774 25.972 176.148 ; 
        RECT 25.436 171.774 25.54 176.148 ; 
        RECT 25.004 171.774 25.108 176.148 ; 
        RECT 24.572 171.774 24.676 176.148 ; 
        RECT 24.14 171.774 24.244 176.148 ; 
        RECT 23.708 171.774 23.812 176.148 ; 
        RECT 22.856 171.774 23.164 176.148 ; 
        RECT 15.284 171.774 15.592 176.148 ; 
        RECT 14.636 171.774 14.74 176.148 ; 
        RECT 14.204 171.774 14.308 176.148 ; 
        RECT 13.772 171.774 13.876 176.148 ; 
        RECT 13.34 171.774 13.444 176.148 ; 
        RECT 12.908 171.774 13.012 176.148 ; 
        RECT 12.476 171.774 12.58 176.148 ; 
        RECT 12.044 171.774 12.148 176.148 ; 
        RECT 11.612 171.774 11.716 176.148 ; 
        RECT 11.18 171.774 11.284 176.148 ; 
        RECT 10.748 171.774 10.852 176.148 ; 
        RECT 10.316 171.774 10.42 176.148 ; 
        RECT 9.884 171.774 9.988 176.148 ; 
        RECT 9.452 171.774 9.556 176.148 ; 
        RECT 9.02 171.774 9.124 176.148 ; 
        RECT 8.588 171.774 8.692 176.148 ; 
        RECT 8.156 171.774 8.26 176.148 ; 
        RECT 7.724 171.774 7.828 176.148 ; 
        RECT 7.292 171.774 7.396 176.148 ; 
        RECT 6.86 171.774 6.964 176.148 ; 
        RECT 6.428 171.774 6.532 176.148 ; 
        RECT 5.996 171.774 6.1 176.148 ; 
        RECT 5.564 171.774 5.668 176.148 ; 
        RECT 5.132 171.774 5.236 176.148 ; 
        RECT 4.7 171.774 4.804 176.148 ; 
        RECT 4.268 171.774 4.372 176.148 ; 
        RECT 3.836 171.774 3.94 176.148 ; 
        RECT 3.404 171.774 3.508 176.148 ; 
        RECT 2.972 171.774 3.076 176.148 ; 
        RECT 2.54 171.774 2.644 176.148 ; 
        RECT 2.108 171.774 2.212 176.148 ; 
        RECT 1.676 171.774 1.78 176.148 ; 
        RECT 1.244 171.774 1.348 176.148 ; 
        RECT 0.812 171.774 0.916 176.148 ; 
        RECT 0 171.774 0.34 176.148 ; 
        RECT 20.72 176.094 21.232 180.468 ; 
        RECT 20.664 178.756 21.232 180.046 ; 
        RECT 20.072 177.664 20.32 180.468 ; 
        RECT 20.016 178.902 20.32 179.516 ; 
        RECT 20.072 176.094 20.176 180.468 ; 
        RECT 20.072 176.578 20.232 177.536 ; 
        RECT 20.072 176.094 20.32 176.45 ; 
        RECT 18.884 177.896 19.708 180.468 ; 
        RECT 19.604 176.094 19.708 180.468 ; 
        RECT 18.884 179.004 19.764 180.036 ; 
        RECT 18.884 176.094 19.276 180.468 ; 
        RECT 17.216 176.094 17.548 180.468 ; 
        RECT 17.216 176.448 17.604 180.19 ; 
        RECT 38.108 176.094 38.448 180.468 ; 
        RECT 37.532 176.094 37.636 180.468 ; 
        RECT 37.1 176.094 37.204 180.468 ; 
        RECT 36.668 176.094 36.772 180.468 ; 
        RECT 36.236 176.094 36.34 180.468 ; 
        RECT 35.804 176.094 35.908 180.468 ; 
        RECT 35.372 176.094 35.476 180.468 ; 
        RECT 34.94 176.094 35.044 180.468 ; 
        RECT 34.508 176.094 34.612 180.468 ; 
        RECT 34.076 176.094 34.18 180.468 ; 
        RECT 33.644 176.094 33.748 180.468 ; 
        RECT 33.212 176.094 33.316 180.468 ; 
        RECT 32.78 176.094 32.884 180.468 ; 
        RECT 32.348 176.094 32.452 180.468 ; 
        RECT 31.916 176.094 32.02 180.468 ; 
        RECT 31.484 176.094 31.588 180.468 ; 
        RECT 31.052 176.094 31.156 180.468 ; 
        RECT 30.62 176.094 30.724 180.468 ; 
        RECT 30.188 176.094 30.292 180.468 ; 
        RECT 29.756 176.094 29.86 180.468 ; 
        RECT 29.324 176.094 29.428 180.468 ; 
        RECT 28.892 176.094 28.996 180.468 ; 
        RECT 28.46 176.094 28.564 180.468 ; 
        RECT 28.028 176.094 28.132 180.468 ; 
        RECT 27.596 176.094 27.7 180.468 ; 
        RECT 27.164 176.094 27.268 180.468 ; 
        RECT 26.732 176.094 26.836 180.468 ; 
        RECT 26.3 176.094 26.404 180.468 ; 
        RECT 25.868 176.094 25.972 180.468 ; 
        RECT 25.436 176.094 25.54 180.468 ; 
        RECT 25.004 176.094 25.108 180.468 ; 
        RECT 24.572 176.094 24.676 180.468 ; 
        RECT 24.14 176.094 24.244 180.468 ; 
        RECT 23.708 176.094 23.812 180.468 ; 
        RECT 22.856 176.094 23.164 180.468 ; 
        RECT 15.284 176.094 15.592 180.468 ; 
        RECT 14.636 176.094 14.74 180.468 ; 
        RECT 14.204 176.094 14.308 180.468 ; 
        RECT 13.772 176.094 13.876 180.468 ; 
        RECT 13.34 176.094 13.444 180.468 ; 
        RECT 12.908 176.094 13.012 180.468 ; 
        RECT 12.476 176.094 12.58 180.468 ; 
        RECT 12.044 176.094 12.148 180.468 ; 
        RECT 11.612 176.094 11.716 180.468 ; 
        RECT 11.18 176.094 11.284 180.468 ; 
        RECT 10.748 176.094 10.852 180.468 ; 
        RECT 10.316 176.094 10.42 180.468 ; 
        RECT 9.884 176.094 9.988 180.468 ; 
        RECT 9.452 176.094 9.556 180.468 ; 
        RECT 9.02 176.094 9.124 180.468 ; 
        RECT 8.588 176.094 8.692 180.468 ; 
        RECT 8.156 176.094 8.26 180.468 ; 
        RECT 7.724 176.094 7.828 180.468 ; 
        RECT 7.292 176.094 7.396 180.468 ; 
        RECT 6.86 176.094 6.964 180.468 ; 
        RECT 6.428 176.094 6.532 180.468 ; 
        RECT 5.996 176.094 6.1 180.468 ; 
        RECT 5.564 176.094 5.668 180.468 ; 
        RECT 5.132 176.094 5.236 180.468 ; 
        RECT 4.7 176.094 4.804 180.468 ; 
        RECT 4.268 176.094 4.372 180.468 ; 
        RECT 3.836 176.094 3.94 180.468 ; 
        RECT 3.404 176.094 3.508 180.468 ; 
        RECT 2.972 176.094 3.076 180.468 ; 
        RECT 2.54 176.094 2.644 180.468 ; 
        RECT 2.108 176.094 2.212 180.468 ; 
        RECT 1.676 176.094 1.78 180.468 ; 
        RECT 1.244 176.094 1.348 180.468 ; 
        RECT 0.812 176.094 0.916 180.468 ; 
        RECT 0 176.094 0.34 180.468 ; 
  LAYER V3 ; 
      RECT 0 4.88 38.448 5.4 ; 
      RECT 37.98 1.026 38.448 5.4 ; 
      RECT 23.364 4.496 37.908 5.4 ; 
      RECT 18.036 4.496 23.292 5.4 ; 
      RECT 15.156 1.026 17.676 5.4 ; 
      RECT 0.54 4.496 15.084 5.4 ; 
      RECT 0 1.026 0.468 5.4 ; 
      RECT 37.836 1.026 38.448 4.688 ; 
      RECT 23.58 1.026 37.764 5.4 ; 
      RECT 20.592 1.026 23.508 4.688 ; 
      RECT 19.944 1.808 20.448 5.4 ; 
      RECT 14.94 1.424 19.836 4.688 ; 
      RECT 0.684 1.026 14.868 5.4 ; 
      RECT 0 1.026 0.612 4.688 ; 
      RECT 20.376 1.026 38.448 4.304 ; 
      RECT 0 1.424 20.304 4.304 ; 
      RECT 19.476 1.026 38.448 1.712 ; 
      RECT 0 1.026 19.404 4.304 ; 
      RECT 0 1.026 38.448 1.328 ; 
      RECT 0 9.2 38.448 9.72 ; 
      RECT 37.98 5.346 38.448 9.72 ; 
      RECT 23.364 8.816 37.908 9.72 ; 
      RECT 18.036 8.816 23.292 9.72 ; 
      RECT 15.156 5.346 17.676 9.72 ; 
      RECT 0.54 8.816 15.084 9.72 ; 
      RECT 0 5.346 0.468 9.72 ; 
      RECT 37.836 5.346 38.448 9.008 ; 
      RECT 23.58 5.346 37.764 9.72 ; 
      RECT 20.592 5.346 23.508 9.008 ; 
      RECT 19.944 6.128 20.448 9.72 ; 
      RECT 14.94 5.744 19.836 9.008 ; 
      RECT 0.684 5.346 14.868 9.72 ; 
      RECT 0 5.346 0.612 9.008 ; 
      RECT 20.376 5.346 38.448 8.624 ; 
      RECT 0 5.744 20.304 8.624 ; 
      RECT 19.476 5.346 38.448 6.032 ; 
      RECT 0 5.346 19.404 8.624 ; 
      RECT 0 5.346 38.448 5.648 ; 
      RECT 0 13.52 38.448 14.04 ; 
      RECT 37.98 9.666 38.448 14.04 ; 
      RECT 23.364 13.136 37.908 14.04 ; 
      RECT 18.036 13.136 23.292 14.04 ; 
      RECT 15.156 9.666 17.676 14.04 ; 
      RECT 0.54 13.136 15.084 14.04 ; 
      RECT 0 9.666 0.468 14.04 ; 
      RECT 37.836 9.666 38.448 13.328 ; 
      RECT 23.58 9.666 37.764 14.04 ; 
      RECT 20.592 9.666 23.508 13.328 ; 
      RECT 19.944 10.448 20.448 14.04 ; 
      RECT 14.94 10.064 19.836 13.328 ; 
      RECT 0.684 9.666 14.868 14.04 ; 
      RECT 0 9.666 0.612 13.328 ; 
      RECT 20.376 9.666 38.448 12.944 ; 
      RECT 0 10.064 20.304 12.944 ; 
      RECT 19.476 9.666 38.448 10.352 ; 
      RECT 0 9.666 19.404 12.944 ; 
      RECT 0 9.666 38.448 9.968 ; 
      RECT 0 17.84 38.448 18.36 ; 
      RECT 37.98 13.986 38.448 18.36 ; 
      RECT 23.364 17.456 37.908 18.36 ; 
      RECT 18.036 17.456 23.292 18.36 ; 
      RECT 15.156 13.986 17.676 18.36 ; 
      RECT 0.54 17.456 15.084 18.36 ; 
      RECT 0 13.986 0.468 18.36 ; 
      RECT 37.836 13.986 38.448 17.648 ; 
      RECT 23.58 13.986 37.764 18.36 ; 
      RECT 20.592 13.986 23.508 17.648 ; 
      RECT 19.944 14.768 20.448 18.36 ; 
      RECT 14.94 14.384 19.836 17.648 ; 
      RECT 0.684 13.986 14.868 18.36 ; 
      RECT 0 13.986 0.612 17.648 ; 
      RECT 20.376 13.986 38.448 17.264 ; 
      RECT 0 14.384 20.304 17.264 ; 
      RECT 19.476 13.986 38.448 14.672 ; 
      RECT 0 13.986 19.404 17.264 ; 
      RECT 0 13.986 38.448 14.288 ; 
      RECT 0 22.16 38.448 22.68 ; 
      RECT 37.98 18.306 38.448 22.68 ; 
      RECT 23.364 21.776 37.908 22.68 ; 
      RECT 18.036 21.776 23.292 22.68 ; 
      RECT 15.156 18.306 17.676 22.68 ; 
      RECT 0.54 21.776 15.084 22.68 ; 
      RECT 0 18.306 0.468 22.68 ; 
      RECT 37.836 18.306 38.448 21.968 ; 
      RECT 23.58 18.306 37.764 22.68 ; 
      RECT 20.592 18.306 23.508 21.968 ; 
      RECT 19.944 19.088 20.448 22.68 ; 
      RECT 14.94 18.704 19.836 21.968 ; 
      RECT 0.684 18.306 14.868 22.68 ; 
      RECT 0 18.306 0.612 21.968 ; 
      RECT 20.376 18.306 38.448 21.584 ; 
      RECT 0 18.704 20.304 21.584 ; 
      RECT 19.476 18.306 38.448 18.992 ; 
      RECT 0 18.306 19.404 21.584 ; 
      RECT 0 18.306 38.448 18.608 ; 
      RECT 0 26.48 38.448 27 ; 
      RECT 37.98 22.626 38.448 27 ; 
      RECT 23.364 26.096 37.908 27 ; 
      RECT 18.036 26.096 23.292 27 ; 
      RECT 15.156 22.626 17.676 27 ; 
      RECT 0.54 26.096 15.084 27 ; 
      RECT 0 22.626 0.468 27 ; 
      RECT 37.836 22.626 38.448 26.288 ; 
      RECT 23.58 22.626 37.764 27 ; 
      RECT 20.592 22.626 23.508 26.288 ; 
      RECT 19.944 23.408 20.448 27 ; 
      RECT 14.94 23.024 19.836 26.288 ; 
      RECT 0.684 22.626 14.868 27 ; 
      RECT 0 22.626 0.612 26.288 ; 
      RECT 20.376 22.626 38.448 25.904 ; 
      RECT 0 23.024 20.304 25.904 ; 
      RECT 19.476 22.626 38.448 23.312 ; 
      RECT 0 22.626 19.404 25.904 ; 
      RECT 0 22.626 38.448 22.928 ; 
      RECT 0 30.8 38.448 31.32 ; 
      RECT 37.98 26.946 38.448 31.32 ; 
      RECT 23.364 30.416 37.908 31.32 ; 
      RECT 18.036 30.416 23.292 31.32 ; 
      RECT 15.156 26.946 17.676 31.32 ; 
      RECT 0.54 30.416 15.084 31.32 ; 
      RECT 0 26.946 0.468 31.32 ; 
      RECT 37.836 26.946 38.448 30.608 ; 
      RECT 23.58 26.946 37.764 31.32 ; 
      RECT 20.592 26.946 23.508 30.608 ; 
      RECT 19.944 27.728 20.448 31.32 ; 
      RECT 14.94 27.344 19.836 30.608 ; 
      RECT 0.684 26.946 14.868 31.32 ; 
      RECT 0 26.946 0.612 30.608 ; 
      RECT 20.376 26.946 38.448 30.224 ; 
      RECT 0 27.344 20.304 30.224 ; 
      RECT 19.476 26.946 38.448 27.632 ; 
      RECT 0 26.946 19.404 30.224 ; 
      RECT 0 26.946 38.448 27.248 ; 
      RECT 0 35.12 38.448 35.64 ; 
      RECT 37.98 31.266 38.448 35.64 ; 
      RECT 23.364 34.736 37.908 35.64 ; 
      RECT 18.036 34.736 23.292 35.64 ; 
      RECT 15.156 31.266 17.676 35.64 ; 
      RECT 0.54 34.736 15.084 35.64 ; 
      RECT 0 31.266 0.468 35.64 ; 
      RECT 37.836 31.266 38.448 34.928 ; 
      RECT 23.58 31.266 37.764 35.64 ; 
      RECT 20.592 31.266 23.508 34.928 ; 
      RECT 19.944 32.048 20.448 35.64 ; 
      RECT 14.94 31.664 19.836 34.928 ; 
      RECT 0.684 31.266 14.868 35.64 ; 
      RECT 0 31.266 0.612 34.928 ; 
      RECT 20.376 31.266 38.448 34.544 ; 
      RECT 0 31.664 20.304 34.544 ; 
      RECT 19.476 31.266 38.448 31.952 ; 
      RECT 0 31.266 19.404 34.544 ; 
      RECT 0 31.266 38.448 31.568 ; 
      RECT 0 39.44 38.448 39.96 ; 
      RECT 37.98 35.586 38.448 39.96 ; 
      RECT 23.364 39.056 37.908 39.96 ; 
      RECT 18.036 39.056 23.292 39.96 ; 
      RECT 15.156 35.586 17.676 39.96 ; 
      RECT 0.54 39.056 15.084 39.96 ; 
      RECT 0 35.586 0.468 39.96 ; 
      RECT 37.836 35.586 38.448 39.248 ; 
      RECT 23.58 35.586 37.764 39.96 ; 
      RECT 20.592 35.586 23.508 39.248 ; 
      RECT 19.944 36.368 20.448 39.96 ; 
      RECT 14.94 35.984 19.836 39.248 ; 
      RECT 0.684 35.586 14.868 39.96 ; 
      RECT 0 35.586 0.612 39.248 ; 
      RECT 20.376 35.586 38.448 38.864 ; 
      RECT 0 35.984 20.304 38.864 ; 
      RECT 19.476 35.586 38.448 36.272 ; 
      RECT 0 35.586 19.404 38.864 ; 
      RECT 0 35.586 38.448 35.888 ; 
      RECT 0 43.76 38.448 44.28 ; 
      RECT 37.98 39.906 38.448 44.28 ; 
      RECT 23.364 43.376 37.908 44.28 ; 
      RECT 18.036 43.376 23.292 44.28 ; 
      RECT 15.156 39.906 17.676 44.28 ; 
      RECT 0.54 43.376 15.084 44.28 ; 
      RECT 0 39.906 0.468 44.28 ; 
      RECT 37.836 39.906 38.448 43.568 ; 
      RECT 23.58 39.906 37.764 44.28 ; 
      RECT 20.592 39.906 23.508 43.568 ; 
      RECT 19.944 40.688 20.448 44.28 ; 
      RECT 14.94 40.304 19.836 43.568 ; 
      RECT 0.684 39.906 14.868 44.28 ; 
      RECT 0 39.906 0.612 43.568 ; 
      RECT 20.376 39.906 38.448 43.184 ; 
      RECT 0 40.304 20.304 43.184 ; 
      RECT 19.476 39.906 38.448 40.592 ; 
      RECT 0 39.906 19.404 43.184 ; 
      RECT 0 39.906 38.448 40.208 ; 
      RECT 0 48.08 38.448 48.6 ; 
      RECT 37.98 44.226 38.448 48.6 ; 
      RECT 23.364 47.696 37.908 48.6 ; 
      RECT 18.036 47.696 23.292 48.6 ; 
      RECT 15.156 44.226 17.676 48.6 ; 
      RECT 0.54 47.696 15.084 48.6 ; 
      RECT 0 44.226 0.468 48.6 ; 
      RECT 37.836 44.226 38.448 47.888 ; 
      RECT 23.58 44.226 37.764 48.6 ; 
      RECT 20.592 44.226 23.508 47.888 ; 
      RECT 19.944 45.008 20.448 48.6 ; 
      RECT 14.94 44.624 19.836 47.888 ; 
      RECT 0.684 44.226 14.868 48.6 ; 
      RECT 0 44.226 0.612 47.888 ; 
      RECT 20.376 44.226 38.448 47.504 ; 
      RECT 0 44.624 20.304 47.504 ; 
      RECT 19.476 44.226 38.448 44.912 ; 
      RECT 0 44.226 19.404 47.504 ; 
      RECT 0 44.226 38.448 44.528 ; 
      RECT 0 52.4 38.448 52.92 ; 
      RECT 37.98 48.546 38.448 52.92 ; 
      RECT 23.364 52.016 37.908 52.92 ; 
      RECT 18.036 52.016 23.292 52.92 ; 
      RECT 15.156 48.546 17.676 52.92 ; 
      RECT 0.54 52.016 15.084 52.92 ; 
      RECT 0 48.546 0.468 52.92 ; 
      RECT 37.836 48.546 38.448 52.208 ; 
      RECT 23.58 48.546 37.764 52.92 ; 
      RECT 20.592 48.546 23.508 52.208 ; 
      RECT 19.944 49.328 20.448 52.92 ; 
      RECT 14.94 48.944 19.836 52.208 ; 
      RECT 0.684 48.546 14.868 52.92 ; 
      RECT 0 48.546 0.612 52.208 ; 
      RECT 20.376 48.546 38.448 51.824 ; 
      RECT 0 48.944 20.304 51.824 ; 
      RECT 19.476 48.546 38.448 49.232 ; 
      RECT 0 48.546 19.404 51.824 ; 
      RECT 0 48.546 38.448 48.848 ; 
      RECT 0 56.72 38.448 57.24 ; 
      RECT 37.98 52.866 38.448 57.24 ; 
      RECT 23.364 56.336 37.908 57.24 ; 
      RECT 18.036 56.336 23.292 57.24 ; 
      RECT 15.156 52.866 17.676 57.24 ; 
      RECT 0.54 56.336 15.084 57.24 ; 
      RECT 0 52.866 0.468 57.24 ; 
      RECT 37.836 52.866 38.448 56.528 ; 
      RECT 23.58 52.866 37.764 57.24 ; 
      RECT 20.592 52.866 23.508 56.528 ; 
      RECT 19.944 53.648 20.448 57.24 ; 
      RECT 14.94 53.264 19.836 56.528 ; 
      RECT 0.684 52.866 14.868 57.24 ; 
      RECT 0 52.866 0.612 56.528 ; 
      RECT 20.376 52.866 38.448 56.144 ; 
      RECT 0 53.264 20.304 56.144 ; 
      RECT 19.476 52.866 38.448 53.552 ; 
      RECT 0 52.866 19.404 56.144 ; 
      RECT 0 52.866 38.448 53.168 ; 
      RECT 0 61.04 38.448 61.56 ; 
      RECT 37.98 57.186 38.448 61.56 ; 
      RECT 23.364 60.656 37.908 61.56 ; 
      RECT 18.036 60.656 23.292 61.56 ; 
      RECT 15.156 57.186 17.676 61.56 ; 
      RECT 0.54 60.656 15.084 61.56 ; 
      RECT 0 57.186 0.468 61.56 ; 
      RECT 37.836 57.186 38.448 60.848 ; 
      RECT 23.58 57.186 37.764 61.56 ; 
      RECT 20.592 57.186 23.508 60.848 ; 
      RECT 19.944 57.968 20.448 61.56 ; 
      RECT 14.94 57.584 19.836 60.848 ; 
      RECT 0.684 57.186 14.868 61.56 ; 
      RECT 0 57.186 0.612 60.848 ; 
      RECT 20.376 57.186 38.448 60.464 ; 
      RECT 0 57.584 20.304 60.464 ; 
      RECT 19.476 57.186 38.448 57.872 ; 
      RECT 0 57.186 19.404 60.464 ; 
      RECT 0 57.186 38.448 57.488 ; 
      RECT 0 65.36 38.448 65.88 ; 
      RECT 37.98 61.506 38.448 65.88 ; 
      RECT 23.364 64.976 37.908 65.88 ; 
      RECT 18.036 64.976 23.292 65.88 ; 
      RECT 15.156 61.506 17.676 65.88 ; 
      RECT 0.54 64.976 15.084 65.88 ; 
      RECT 0 61.506 0.468 65.88 ; 
      RECT 37.836 61.506 38.448 65.168 ; 
      RECT 23.58 61.506 37.764 65.88 ; 
      RECT 20.592 61.506 23.508 65.168 ; 
      RECT 19.944 62.288 20.448 65.88 ; 
      RECT 14.94 61.904 19.836 65.168 ; 
      RECT 0.684 61.506 14.868 65.88 ; 
      RECT 0 61.506 0.612 65.168 ; 
      RECT 20.376 61.506 38.448 64.784 ; 
      RECT 0 61.904 20.304 64.784 ; 
      RECT 19.476 61.506 38.448 62.192 ; 
      RECT 0 61.506 19.404 64.784 ; 
      RECT 0 61.506 38.448 61.808 ; 
      RECT 0 69.68 38.448 70.2 ; 
      RECT 37.98 65.826 38.448 70.2 ; 
      RECT 23.364 69.296 37.908 70.2 ; 
      RECT 18.036 69.296 23.292 70.2 ; 
      RECT 15.156 65.826 17.676 70.2 ; 
      RECT 0.54 69.296 15.084 70.2 ; 
      RECT 0 65.826 0.468 70.2 ; 
      RECT 37.836 65.826 38.448 69.488 ; 
      RECT 23.58 65.826 37.764 70.2 ; 
      RECT 20.592 65.826 23.508 69.488 ; 
      RECT 19.944 66.608 20.448 70.2 ; 
      RECT 14.94 66.224 19.836 69.488 ; 
      RECT 0.684 65.826 14.868 70.2 ; 
      RECT 0 65.826 0.612 69.488 ; 
      RECT 20.376 65.826 38.448 69.104 ; 
      RECT 0 66.224 20.304 69.104 ; 
      RECT 19.476 65.826 38.448 66.512 ; 
      RECT 0 65.826 19.404 69.104 ; 
      RECT 0 65.826 38.448 66.128 ; 
      RECT 0 74 38.448 74.52 ; 
      RECT 37.98 70.146 38.448 74.52 ; 
      RECT 23.364 73.616 37.908 74.52 ; 
      RECT 18.036 73.616 23.292 74.52 ; 
      RECT 15.156 70.146 17.676 74.52 ; 
      RECT 0.54 73.616 15.084 74.52 ; 
      RECT 0 70.146 0.468 74.52 ; 
      RECT 37.836 70.146 38.448 73.808 ; 
      RECT 23.58 70.146 37.764 74.52 ; 
      RECT 20.592 70.146 23.508 73.808 ; 
      RECT 19.944 70.928 20.448 74.52 ; 
      RECT 14.94 70.544 19.836 73.808 ; 
      RECT 0.684 70.146 14.868 74.52 ; 
      RECT 0 70.146 0.612 73.808 ; 
      RECT 20.376 70.146 38.448 73.424 ; 
      RECT 0 70.544 20.304 73.424 ; 
      RECT 19.476 70.146 38.448 70.832 ; 
      RECT 0 70.146 19.404 73.424 ; 
      RECT 0 70.146 38.448 70.448 ; 
      RECT 0 103.692 38.448 109.026 ; 
      RECT 29.412 74.412 38.448 109.026 ; 
      RECT 20.612 89.868 38.448 109.026 ; 
      RECT 24.228 79.5 38.448 109.026 ; 
      RECT 20.404 74.412 20.54 109.026 ; 
      RECT 20.196 74.412 20.332 109.026 ; 
      RECT 19.988 74.412 20.124 109.026 ; 
      RECT 19.78 74.412 19.916 109.026 ; 
      RECT 0 101.964 19.708 109.026 ; 
      RECT 18.74 91.02 38.448 102.828 ; 
      RECT 18.532 74.412 18.668 109.026 ; 
      RECT 18.324 74.412 18.46 109.026 ; 
      RECT 18.116 74.412 18.252 109.026 ; 
      RECT 17.908 74.412 18.044 109.026 ; 
      RECT 0 80.652 17.836 109.026 ; 
      RECT 0 89.292 19.708 101.1 ; 
      RECT 18.74 78.348 23.292 90.156 ; 
      RECT 23.364 80.268 38.448 109.026 ; 
      RECT 20.772 74.732 24.156 89.772 ; 
      RECT 16.02 76.62 19.116 88.428 ; 
      RECT 15.156 77.196 17.836 109.026 ; 
      RECT 0 79.5 15.084 109.026 ; 
      RECT 13.428 74.412 15.228 80.556 ; 
      RECT 28.548 74.412 29.34 109.026 ; 
      RECT 13.428 78.732 28.476 80.172 ; 
      RECT 9.972 77.196 13.356 109.026 ; 
      RECT 0 78.348 9.9 109.026 ; 
      RECT 27.684 74.412 38.448 79.404 ; 
      RECT 26.82 77.196 38.448 79.404 ; 
      RECT 0 78.348 26.748 79.404 ; 
      RECT 25.956 74.412 27.612 78.636 ; 
      RECT 20.612 77.196 38.448 78.636 ; 
      RECT 0.684 77.196 19.708 79.404 ; 
      RECT 18.74 77.004 19.708 109.026 ; 
      RECT 0 76.62 0.612 109.026 ; 
      RECT 19.188 74.412 20.7 77.484 ; 
      RECT 20.772 77.004 25.884 80.172 ; 
      RECT 12.564 77.004 15.948 79.404 ; 
      RECT 10.836 77.004 12.492 109.026 ; 
      RECT 0 76.62 10.764 77.484 ; 
      RECT 25.092 74.412 38.448 77.1 ; 
      RECT 19.188 74.732 25.02 77.1 ; 
      RECT 15.3 76.62 19.116 77.1 ; 
      RECT 11.7 74.412 15.228 77.1 ; 
      RECT 0 76.62 11.628 77.1 ; 
      RECT 23.364 74.412 38.448 76.908 ; 
      RECT 18.74 74.732 38.448 76.908 ; 
      RECT 0.54 74.412 17.836 76.908 ; 
      RECT 0 74.412 0.468 109.026 ; 
      RECT 0 74.412 23.292 75.756 ; 
      RECT 0 74.412 38.448 74.636 ; 
        RECT 0 110.828 38.448 111.348 ; 
        RECT 37.98 106.974 38.448 111.348 ; 
        RECT 23.364 110.444 37.908 111.348 ; 
        RECT 18.036 110.444 23.292 111.348 ; 
        RECT 15.156 106.974 17.676 111.348 ; 
        RECT 0.54 110.444 15.084 111.348 ; 
        RECT 0 106.974 0.468 111.348 ; 
        RECT 37.836 106.974 38.448 110.636 ; 
        RECT 23.58 106.974 37.764 111.348 ; 
        RECT 20.592 106.974 23.508 110.636 ; 
        RECT 19.944 107.756 20.448 111.348 ; 
        RECT 14.94 107.372 19.836 110.636 ; 
        RECT 0.684 106.974 14.868 111.348 ; 
        RECT 0 106.974 0.612 110.636 ; 
        RECT 20.376 106.974 38.448 110.252 ; 
        RECT 0 107.372 20.304 110.252 ; 
        RECT 19.476 106.974 38.448 107.66 ; 
        RECT 0 106.974 19.404 110.252 ; 
        RECT 0 106.974 38.448 107.276 ; 
        RECT 0 115.148 38.448 115.668 ; 
        RECT 37.98 111.294 38.448 115.668 ; 
        RECT 23.364 114.764 37.908 115.668 ; 
        RECT 18.036 114.764 23.292 115.668 ; 
        RECT 15.156 111.294 17.676 115.668 ; 
        RECT 0.54 114.764 15.084 115.668 ; 
        RECT 0 111.294 0.468 115.668 ; 
        RECT 37.836 111.294 38.448 114.956 ; 
        RECT 23.58 111.294 37.764 115.668 ; 
        RECT 20.592 111.294 23.508 114.956 ; 
        RECT 19.944 112.076 20.448 115.668 ; 
        RECT 14.94 111.692 19.836 114.956 ; 
        RECT 0.684 111.294 14.868 115.668 ; 
        RECT 0 111.294 0.612 114.956 ; 
        RECT 20.376 111.294 38.448 114.572 ; 
        RECT 0 111.692 20.304 114.572 ; 
        RECT 19.476 111.294 38.448 111.98 ; 
        RECT 0 111.294 19.404 114.572 ; 
        RECT 0 111.294 38.448 111.596 ; 
        RECT 0 119.468 38.448 119.988 ; 
        RECT 37.98 115.614 38.448 119.988 ; 
        RECT 23.364 119.084 37.908 119.988 ; 
        RECT 18.036 119.084 23.292 119.988 ; 
        RECT 15.156 115.614 17.676 119.988 ; 
        RECT 0.54 119.084 15.084 119.988 ; 
        RECT 0 115.614 0.468 119.988 ; 
        RECT 37.836 115.614 38.448 119.276 ; 
        RECT 23.58 115.614 37.764 119.988 ; 
        RECT 20.592 115.614 23.508 119.276 ; 
        RECT 19.944 116.396 20.448 119.988 ; 
        RECT 14.94 116.012 19.836 119.276 ; 
        RECT 0.684 115.614 14.868 119.988 ; 
        RECT 0 115.614 0.612 119.276 ; 
        RECT 20.376 115.614 38.448 118.892 ; 
        RECT 0 116.012 20.304 118.892 ; 
        RECT 19.476 115.614 38.448 116.3 ; 
        RECT 0 115.614 19.404 118.892 ; 
        RECT 0 115.614 38.448 115.916 ; 
        RECT 0 123.788 38.448 124.308 ; 
        RECT 37.98 119.934 38.448 124.308 ; 
        RECT 23.364 123.404 37.908 124.308 ; 
        RECT 18.036 123.404 23.292 124.308 ; 
        RECT 15.156 119.934 17.676 124.308 ; 
        RECT 0.54 123.404 15.084 124.308 ; 
        RECT 0 119.934 0.468 124.308 ; 
        RECT 37.836 119.934 38.448 123.596 ; 
        RECT 23.58 119.934 37.764 124.308 ; 
        RECT 20.592 119.934 23.508 123.596 ; 
        RECT 19.944 120.716 20.448 124.308 ; 
        RECT 14.94 120.332 19.836 123.596 ; 
        RECT 0.684 119.934 14.868 124.308 ; 
        RECT 0 119.934 0.612 123.596 ; 
        RECT 20.376 119.934 38.448 123.212 ; 
        RECT 0 120.332 20.304 123.212 ; 
        RECT 19.476 119.934 38.448 120.62 ; 
        RECT 0 119.934 19.404 123.212 ; 
        RECT 0 119.934 38.448 120.236 ; 
        RECT 0 128.108 38.448 128.628 ; 
        RECT 37.98 124.254 38.448 128.628 ; 
        RECT 23.364 127.724 37.908 128.628 ; 
        RECT 18.036 127.724 23.292 128.628 ; 
        RECT 15.156 124.254 17.676 128.628 ; 
        RECT 0.54 127.724 15.084 128.628 ; 
        RECT 0 124.254 0.468 128.628 ; 
        RECT 37.836 124.254 38.448 127.916 ; 
        RECT 23.58 124.254 37.764 128.628 ; 
        RECT 20.592 124.254 23.508 127.916 ; 
        RECT 19.944 125.036 20.448 128.628 ; 
        RECT 14.94 124.652 19.836 127.916 ; 
        RECT 0.684 124.254 14.868 128.628 ; 
        RECT 0 124.254 0.612 127.916 ; 
        RECT 20.376 124.254 38.448 127.532 ; 
        RECT 0 124.652 20.304 127.532 ; 
        RECT 19.476 124.254 38.448 124.94 ; 
        RECT 0 124.254 19.404 127.532 ; 
        RECT 0 124.254 38.448 124.556 ; 
        RECT 0 132.428 38.448 132.948 ; 
        RECT 37.98 128.574 38.448 132.948 ; 
        RECT 23.364 132.044 37.908 132.948 ; 
        RECT 18.036 132.044 23.292 132.948 ; 
        RECT 15.156 128.574 17.676 132.948 ; 
        RECT 0.54 132.044 15.084 132.948 ; 
        RECT 0 128.574 0.468 132.948 ; 
        RECT 37.836 128.574 38.448 132.236 ; 
        RECT 23.58 128.574 37.764 132.948 ; 
        RECT 20.592 128.574 23.508 132.236 ; 
        RECT 19.944 129.356 20.448 132.948 ; 
        RECT 14.94 128.972 19.836 132.236 ; 
        RECT 0.684 128.574 14.868 132.948 ; 
        RECT 0 128.574 0.612 132.236 ; 
        RECT 20.376 128.574 38.448 131.852 ; 
        RECT 0 128.972 20.304 131.852 ; 
        RECT 19.476 128.574 38.448 129.26 ; 
        RECT 0 128.574 19.404 131.852 ; 
        RECT 0 128.574 38.448 128.876 ; 
        RECT 0 136.748 38.448 137.268 ; 
        RECT 37.98 132.894 38.448 137.268 ; 
        RECT 23.364 136.364 37.908 137.268 ; 
        RECT 18.036 136.364 23.292 137.268 ; 
        RECT 15.156 132.894 17.676 137.268 ; 
        RECT 0.54 136.364 15.084 137.268 ; 
        RECT 0 132.894 0.468 137.268 ; 
        RECT 37.836 132.894 38.448 136.556 ; 
        RECT 23.58 132.894 37.764 137.268 ; 
        RECT 20.592 132.894 23.508 136.556 ; 
        RECT 19.944 133.676 20.448 137.268 ; 
        RECT 14.94 133.292 19.836 136.556 ; 
        RECT 0.684 132.894 14.868 137.268 ; 
        RECT 0 132.894 0.612 136.556 ; 
        RECT 20.376 132.894 38.448 136.172 ; 
        RECT 0 133.292 20.304 136.172 ; 
        RECT 19.476 132.894 38.448 133.58 ; 
        RECT 0 132.894 19.404 136.172 ; 
        RECT 0 132.894 38.448 133.196 ; 
        RECT 0 141.068 38.448 141.588 ; 
        RECT 37.98 137.214 38.448 141.588 ; 
        RECT 23.364 140.684 37.908 141.588 ; 
        RECT 18.036 140.684 23.292 141.588 ; 
        RECT 15.156 137.214 17.676 141.588 ; 
        RECT 0.54 140.684 15.084 141.588 ; 
        RECT 0 137.214 0.468 141.588 ; 
        RECT 37.836 137.214 38.448 140.876 ; 
        RECT 23.58 137.214 37.764 141.588 ; 
        RECT 20.592 137.214 23.508 140.876 ; 
        RECT 19.944 137.996 20.448 141.588 ; 
        RECT 14.94 137.612 19.836 140.876 ; 
        RECT 0.684 137.214 14.868 141.588 ; 
        RECT 0 137.214 0.612 140.876 ; 
        RECT 20.376 137.214 38.448 140.492 ; 
        RECT 0 137.612 20.304 140.492 ; 
        RECT 19.476 137.214 38.448 137.9 ; 
        RECT 0 137.214 19.404 140.492 ; 
        RECT 0 137.214 38.448 137.516 ; 
        RECT 0 145.388 38.448 145.908 ; 
        RECT 37.98 141.534 38.448 145.908 ; 
        RECT 23.364 145.004 37.908 145.908 ; 
        RECT 18.036 145.004 23.292 145.908 ; 
        RECT 15.156 141.534 17.676 145.908 ; 
        RECT 0.54 145.004 15.084 145.908 ; 
        RECT 0 141.534 0.468 145.908 ; 
        RECT 37.836 141.534 38.448 145.196 ; 
        RECT 23.58 141.534 37.764 145.908 ; 
        RECT 20.592 141.534 23.508 145.196 ; 
        RECT 19.944 142.316 20.448 145.908 ; 
        RECT 14.94 141.932 19.836 145.196 ; 
        RECT 0.684 141.534 14.868 145.908 ; 
        RECT 0 141.534 0.612 145.196 ; 
        RECT 20.376 141.534 38.448 144.812 ; 
        RECT 0 141.932 20.304 144.812 ; 
        RECT 19.476 141.534 38.448 142.22 ; 
        RECT 0 141.534 19.404 144.812 ; 
        RECT 0 141.534 38.448 141.836 ; 
        RECT 0 149.708 38.448 150.228 ; 
        RECT 37.98 145.854 38.448 150.228 ; 
        RECT 23.364 149.324 37.908 150.228 ; 
        RECT 18.036 149.324 23.292 150.228 ; 
        RECT 15.156 145.854 17.676 150.228 ; 
        RECT 0.54 149.324 15.084 150.228 ; 
        RECT 0 145.854 0.468 150.228 ; 
        RECT 37.836 145.854 38.448 149.516 ; 
        RECT 23.58 145.854 37.764 150.228 ; 
        RECT 20.592 145.854 23.508 149.516 ; 
        RECT 19.944 146.636 20.448 150.228 ; 
        RECT 14.94 146.252 19.836 149.516 ; 
        RECT 0.684 145.854 14.868 150.228 ; 
        RECT 0 145.854 0.612 149.516 ; 
        RECT 20.376 145.854 38.448 149.132 ; 
        RECT 0 146.252 20.304 149.132 ; 
        RECT 19.476 145.854 38.448 146.54 ; 
        RECT 0 145.854 19.404 149.132 ; 
        RECT 0 145.854 38.448 146.156 ; 
        RECT 0 154.028 38.448 154.548 ; 
        RECT 37.98 150.174 38.448 154.548 ; 
        RECT 23.364 153.644 37.908 154.548 ; 
        RECT 18.036 153.644 23.292 154.548 ; 
        RECT 15.156 150.174 17.676 154.548 ; 
        RECT 0.54 153.644 15.084 154.548 ; 
        RECT 0 150.174 0.468 154.548 ; 
        RECT 37.836 150.174 38.448 153.836 ; 
        RECT 23.58 150.174 37.764 154.548 ; 
        RECT 20.592 150.174 23.508 153.836 ; 
        RECT 19.944 150.956 20.448 154.548 ; 
        RECT 14.94 150.572 19.836 153.836 ; 
        RECT 0.684 150.174 14.868 154.548 ; 
        RECT 0 150.174 0.612 153.836 ; 
        RECT 20.376 150.174 38.448 153.452 ; 
        RECT 0 150.572 20.304 153.452 ; 
        RECT 19.476 150.174 38.448 150.86 ; 
        RECT 0 150.174 19.404 153.452 ; 
        RECT 0 150.174 38.448 150.476 ; 
        RECT 0 158.348 38.448 158.868 ; 
        RECT 37.98 154.494 38.448 158.868 ; 
        RECT 23.364 157.964 37.908 158.868 ; 
        RECT 18.036 157.964 23.292 158.868 ; 
        RECT 15.156 154.494 17.676 158.868 ; 
        RECT 0.54 157.964 15.084 158.868 ; 
        RECT 0 154.494 0.468 158.868 ; 
        RECT 37.836 154.494 38.448 158.156 ; 
        RECT 23.58 154.494 37.764 158.868 ; 
        RECT 20.592 154.494 23.508 158.156 ; 
        RECT 19.944 155.276 20.448 158.868 ; 
        RECT 14.94 154.892 19.836 158.156 ; 
        RECT 0.684 154.494 14.868 158.868 ; 
        RECT 0 154.494 0.612 158.156 ; 
        RECT 20.376 154.494 38.448 157.772 ; 
        RECT 0 154.892 20.304 157.772 ; 
        RECT 19.476 154.494 38.448 155.18 ; 
        RECT 0 154.494 19.404 157.772 ; 
        RECT 0 154.494 38.448 154.796 ; 
        RECT 0 162.668 38.448 163.188 ; 
        RECT 37.98 158.814 38.448 163.188 ; 
        RECT 23.364 162.284 37.908 163.188 ; 
        RECT 18.036 162.284 23.292 163.188 ; 
        RECT 15.156 158.814 17.676 163.188 ; 
        RECT 0.54 162.284 15.084 163.188 ; 
        RECT 0 158.814 0.468 163.188 ; 
        RECT 37.836 158.814 38.448 162.476 ; 
        RECT 23.58 158.814 37.764 163.188 ; 
        RECT 20.592 158.814 23.508 162.476 ; 
        RECT 19.944 159.596 20.448 163.188 ; 
        RECT 14.94 159.212 19.836 162.476 ; 
        RECT 0.684 158.814 14.868 163.188 ; 
        RECT 0 158.814 0.612 162.476 ; 
        RECT 20.376 158.814 38.448 162.092 ; 
        RECT 0 159.212 20.304 162.092 ; 
        RECT 19.476 158.814 38.448 159.5 ; 
        RECT 0 158.814 19.404 162.092 ; 
        RECT 0 158.814 38.448 159.116 ; 
        RECT 0 166.988 38.448 167.508 ; 
        RECT 37.98 163.134 38.448 167.508 ; 
        RECT 23.364 166.604 37.908 167.508 ; 
        RECT 18.036 166.604 23.292 167.508 ; 
        RECT 15.156 163.134 17.676 167.508 ; 
        RECT 0.54 166.604 15.084 167.508 ; 
        RECT 0 163.134 0.468 167.508 ; 
        RECT 37.836 163.134 38.448 166.796 ; 
        RECT 23.58 163.134 37.764 167.508 ; 
        RECT 20.592 163.134 23.508 166.796 ; 
        RECT 19.944 163.916 20.448 167.508 ; 
        RECT 14.94 163.532 19.836 166.796 ; 
        RECT 0.684 163.134 14.868 167.508 ; 
        RECT 0 163.134 0.612 166.796 ; 
        RECT 20.376 163.134 38.448 166.412 ; 
        RECT 0 163.532 20.304 166.412 ; 
        RECT 19.476 163.134 38.448 163.82 ; 
        RECT 0 163.134 19.404 166.412 ; 
        RECT 0 163.134 38.448 163.436 ; 
        RECT 0 171.308 38.448 171.828 ; 
        RECT 37.98 167.454 38.448 171.828 ; 
        RECT 23.364 170.924 37.908 171.828 ; 
        RECT 18.036 170.924 23.292 171.828 ; 
        RECT 15.156 167.454 17.676 171.828 ; 
        RECT 0.54 170.924 15.084 171.828 ; 
        RECT 0 167.454 0.468 171.828 ; 
        RECT 37.836 167.454 38.448 171.116 ; 
        RECT 23.58 167.454 37.764 171.828 ; 
        RECT 20.592 167.454 23.508 171.116 ; 
        RECT 19.944 168.236 20.448 171.828 ; 
        RECT 14.94 167.852 19.836 171.116 ; 
        RECT 0.684 167.454 14.868 171.828 ; 
        RECT 0 167.454 0.612 171.116 ; 
        RECT 20.376 167.454 38.448 170.732 ; 
        RECT 0 167.852 20.304 170.732 ; 
        RECT 19.476 167.454 38.448 168.14 ; 
        RECT 0 167.454 19.404 170.732 ; 
        RECT 0 167.454 38.448 167.756 ; 
        RECT 0 175.628 38.448 176.148 ; 
        RECT 37.98 171.774 38.448 176.148 ; 
        RECT 23.364 175.244 37.908 176.148 ; 
        RECT 18.036 175.244 23.292 176.148 ; 
        RECT 15.156 171.774 17.676 176.148 ; 
        RECT 0.54 175.244 15.084 176.148 ; 
        RECT 0 171.774 0.468 176.148 ; 
        RECT 37.836 171.774 38.448 175.436 ; 
        RECT 23.58 171.774 37.764 176.148 ; 
        RECT 20.592 171.774 23.508 175.436 ; 
        RECT 19.944 172.556 20.448 176.148 ; 
        RECT 14.94 172.172 19.836 175.436 ; 
        RECT 0.684 171.774 14.868 176.148 ; 
        RECT 0 171.774 0.612 175.436 ; 
        RECT 20.376 171.774 38.448 175.052 ; 
        RECT 0 172.172 20.304 175.052 ; 
        RECT 19.476 171.774 38.448 172.46 ; 
        RECT 0 171.774 19.404 175.052 ; 
        RECT 0 171.774 38.448 172.076 ; 
        RECT 0 179.948 38.448 180.468 ; 
        RECT 37.98 176.094 38.448 180.468 ; 
        RECT 23.364 179.564 37.908 180.468 ; 
        RECT 18.036 179.564 23.292 180.468 ; 
        RECT 15.156 176.094 17.676 180.468 ; 
        RECT 0.54 179.564 15.084 180.468 ; 
        RECT 0 176.094 0.468 180.468 ; 
        RECT 37.836 176.094 38.448 179.756 ; 
        RECT 23.58 176.094 37.764 180.468 ; 
        RECT 20.592 176.094 23.508 179.756 ; 
        RECT 19.944 176.876 20.448 180.468 ; 
        RECT 14.94 176.492 19.836 179.756 ; 
        RECT 0.684 176.094 14.868 180.468 ; 
        RECT 0 176.094 0.612 179.756 ; 
        RECT 20.376 176.094 38.448 179.372 ; 
        RECT 0 176.492 20.304 179.372 ; 
        RECT 19.476 176.094 38.448 176.78 ; 
        RECT 0 176.094 19.404 179.372 ; 
        RECT 0 176.094 38.448 176.396 ; 
  LAYER M4 ; 
      RECT 6.428 81.264 32.01 81.36 ; 
      RECT 6.428 82.416 32.01 82.512 ; 
      RECT 6.428 83.952 32.01 84.048 ; 
      RECT 6.428 84.336 32.01 84.432 ; 
      RECT 6.428 85.68 32.01 85.776 ; 
      RECT 29.996 77.1 30.332 77.196 ; 
      RECT 29.276 78.828 29.744 78.924 ; 
      RECT 29.276 81.456 29.744 81.552 ; 
      RECT 29.276 82.608 29.744 82.704 ; 
      RECT 26.714 78.828 28.992 78.924 ; 
      RECT 26.972 81.936 27.404 82.032 ; 
      RECT 21.628 83.436 26 83.532 ; 
      RECT 24.38 81.708 24.716 81.804 ; 
      RECT 21.244 86.508 24.716 86.604 ; 
      RECT 24.38 86.892 24.716 86.988 ; 
      RECT 23.668 79.788 24.004 79.884 ; 
      RECT 23.516 85.164 23.852 85.26 ; 
      RECT 22.804 79.404 23.14 79.5 ; 
      RECT 21.948 74.252 23 74.348 ; 
      RECT 21.948 108.812 23 108.908 ; 
      RECT 22.012 85.356 22.988 85.452 ; 
      RECT 22.652 85.932 22.988 86.028 ; 
      RECT 16.828 86.892 22.988 86.988 ; 
      RECT 22.652 88.044 22.988 88.14 ; 
      RECT 21.716 108.428 22.768 108.524 ; 
      RECT 21.712 73.868 22.764 73.964 ; 
      RECT 21.56 73.484 22.612 73.58 ; 
      RECT 21.56 107.66 22.612 107.756 ; 
      RECT 22.22 89.772 22.556 89.868 ; 
      RECT 19.132 91.308 22.556 91.404 ; 
      RECT 20.668 100.332 22.556 100.428 ; 
      RECT 22.22 100.716 22.556 100.812 ; 
      RECT 21.368 73.1 22.42 73.196 ; 
      RECT 21.368 107.276 22.42 107.372 ; 
      RECT 20.476 96.684 22.256 96.78 ; 
      RECT 21.192 72.716 22.244 72.812 ; 
      RECT 21.192 108.62 22.244 108.716 ; 
      RECT 20.996 74.06 22.048 74.156 ; 
      RECT 20.996 108.236 22.048 108.332 ; 
      RECT 21.52 85.932 22.004 86.028 ; 
      RECT 21.436 94.38 21.968 94.476 ; 
      RECT 20.808 73.676 21.86 73.772 ; 
      RECT 20.808 107.852 21.86 107.948 ; 
      RECT 20.668 72.524 21.72 72.62 ; 
      RECT 20.668 107.468 21.72 107.564 ; 
      RECT 17.404 100.716 21.68 100.812 ; 
      RECT 21.344 105.324 21.68 105.42 ; 
      RECT 20.444 71.948 21.496 72.044 ; 
      RECT 20.444 107.084 21.496 107.18 ; 
      RECT 21.052 89.772 21.392 89.868 ; 
      RECT 16.636 92.076 21.104 92.172 ; 
      RECT 19.216 83.436 21.044 83.532 ; 
      RECT 18.524 74.828 19.592 74.924 ; 
      RECT 18.524 106.508 19.592 106.604 ; 
      RECT 19.072 89.58 19.508 89.676 ; 
      RECT 18.432 74.444 19.4 74.54 ; 
      RECT 18.432 109.004 19.4 109.1 ; 
      RECT 18.208 72.524 19.176 72.62 ; 
      RECT 18.324 109.388 19.176 109.484 ; 
      RECT 18.788 88.044 19.124 88.14 ; 
      RECT 17.992 72.908 18.984 73.004 ; 
      RECT 17.992 108.812 18.984 108.908 ; 
      RECT 17.056 98.412 18.74 98.508 ; 
      RECT 16.928 74.252 17.996 74.348 ; 
      RECT 16.928 109.388 17.996 109.484 ; 
      RECT 17.488 92.652 17.972 92.748 ; 
      RECT 17.456 105.324 17.792 105.42 ; 
      RECT 16.792 73.868 17.78 73.964 ; 
      RECT 16.524 107.66 17.78 107.756 ; 
      RECT 16.688 73.484 17.608 73.58 ; 
      RECT 16.64 109.004 17.608 109.1 ; 
      RECT 16.476 73.1 17.396 73.196 ; 
      RECT 17.06 98.988 17.396 99.084 ; 
      RECT 16.276 107.276 17.396 107.372 ; 
      RECT 16.296 72.716 17.216 72.812 ; 
      RECT 16.296 108.62 17.216 108.716 ; 
      RECT 12.448 88.044 17.204 88.14 ; 
      RECT 16.144 73.676 17.064 73.772 ; 
      RECT 16.144 108.236 17.064 108.332 ; 
      RECT 16.072 73.292 16.844 73.388 ; 
      RECT 16.072 107.852 16.844 107.948 ; 
      RECT 15.876 72.908 16.648 73.004 ; 
      RECT 15.876 107.468 16.648 107.564 ; 
      RECT 15.892 91.692 16.628 91.788 ; 
      RECT 15.668 72.524 16.44 72.62 ; 
      RECT 15.668 107.084 16.44 107.18 ; 
      RECT 13.732 80.94 16.436 81.036 ; 
      RECT 15.892 92.076 16.228 92.172 ; 
      RECT 14.816 74.636 15.868 74.732 ; 
      RECT 15.032 89.772 15.48 89.868 ; 
      RECT 13.58 81.708 13.916 81.804 ; 
  LAYER V4 ; 
      RECT 30.192 77.1 30.288 77.196 ; 
      RECT 30.192 81.264 30.288 81.36 ; 
      RECT 29.52 78.828 29.616 78.924 ; 
      RECT 29.52 81.456 29.616 81.552 ; 
      RECT 29.52 82.608 29.616 82.704 ; 
      RECT 27.024 78.828 27.12 78.924 ; 
      RECT 27.024 81.936 27.12 82.032 ; 
      RECT 24.576 81.708 24.672 81.804 ; 
      RECT 24.576 82.416 24.672 82.512 ; 
      RECT 24.576 86.508 24.672 86.604 ; 
      RECT 24.576 86.892 24.672 86.988 ; 
      RECT 23.712 79.788 23.808 79.884 ; 
      RECT 23.712 83.952 23.808 84.048 ; 
      RECT 23.712 85.164 23.808 85.26 ; 
      RECT 23.712 85.68 23.808 85.776 ; 
      RECT 22.848 79.404 22.944 79.5 ; 
      RECT 22.848 84.336 22.944 84.432 ; 
      RECT 22.848 85.356 22.944 85.452 ; 
      RECT 22.848 85.932 22.944 86.028 ; 
      RECT 22.848 86.892 22.944 86.988 ; 
      RECT 22.848 88.044 22.944 88.14 ; 
      RECT 22.416 89.772 22.512 89.868 ; 
      RECT 22.416 91.308 22.512 91.404 ; 
      RECT 22.416 100.332 22.512 100.428 ; 
      RECT 22.416 100.716 22.512 100.812 ; 
      RECT 22.056 74.252 22.152 74.348 ; 
      RECT 22.056 85.356 22.152 85.452 ; 
      RECT 22.056 108.812 22.152 108.908 ; 
      RECT 21.864 73.868 21.96 73.964 ; 
      RECT 21.864 85.932 21.96 86.028 ; 
      RECT 21.864 108.428 21.96 108.524 ; 
      RECT 21.672 73.484 21.768 73.58 ; 
      RECT 21.672 83.436 21.768 83.532 ; 
      RECT 21.672 107.66 21.768 107.756 ; 
      RECT 21.48 73.1 21.576 73.196 ; 
      RECT 21.48 94.38 21.576 94.476 ; 
      RECT 21.48 105.324 21.576 105.42 ; 
      RECT 21.48 107.276 21.576 107.372 ; 
      RECT 21.288 72.716 21.384 72.812 ; 
      RECT 21.288 86.508 21.384 86.604 ; 
      RECT 21.288 108.62 21.384 108.716 ; 
      RECT 21.096 74.06 21.192 74.156 ; 
      RECT 21.096 89.772 21.192 89.868 ; 
      RECT 21.096 108.236 21.192 108.332 ; 
      RECT 20.904 73.676 21 73.772 ; 
      RECT 20.904 83.436 21 83.532 ; 
      RECT 20.904 107.852 21 107.948 ; 
      RECT 20.712 72.524 20.808 72.62 ; 
      RECT 20.712 100.332 20.808 100.428 ; 
      RECT 20.712 107.468 20.808 107.564 ; 
      RECT 20.52 71.948 20.616 72.044 ; 
      RECT 20.52 96.684 20.616 96.78 ; 
      RECT 20.52 107.084 20.616 107.18 ; 
      RECT 19.368 74.828 19.464 74.924 ; 
      RECT 19.368 89.58 19.464 89.676 ; 
      RECT 19.368 106.508 19.464 106.604 ; 
      RECT 19.176 74.444 19.272 74.54 ; 
      RECT 19.176 91.308 19.272 91.404 ; 
      RECT 19.176 109.004 19.272 109.1 ; 
      RECT 18.984 72.524 19.08 72.62 ; 
      RECT 18.984 88.044 19.08 88.14 ; 
      RECT 18.984 109.388 19.08 109.484 ; 
      RECT 18.6 72.908 18.696 73.004 ; 
      RECT 18.6 98.412 18.696 98.508 ; 
      RECT 18.6 108.812 18.696 108.908 ; 
      RECT 17.832 74.252 17.928 74.348 ; 
      RECT 17.832 92.652 17.928 92.748 ; 
      RECT 17.832 109.388 17.928 109.484 ; 
      RECT 17.64 73.868 17.736 73.964 ; 
      RECT 17.64 105.324 17.736 105.42 ; 
      RECT 17.64 107.66 17.736 107.756 ; 
      RECT 17.448 73.484 17.544 73.58 ; 
      RECT 17.448 100.716 17.544 100.812 ; 
      RECT 17.448 109.004 17.544 109.1 ; 
      RECT 17.256 73.1 17.352 73.196 ; 
      RECT 17.256 98.988 17.352 99.084 ; 
      RECT 17.256 107.276 17.352 107.372 ; 
      RECT 17.064 72.716 17.16 72.812 ; 
      RECT 17.064 88.044 17.16 88.14 ; 
      RECT 17.064 108.62 17.16 108.716 ; 
      RECT 16.872 73.676 16.968 73.772 ; 
      RECT 16.872 86.892 16.968 86.988 ; 
      RECT 16.872 108.236 16.968 108.332 ; 
      RECT 16.68 73.292 16.776 73.388 ; 
      RECT 16.68 92.076 16.776 92.172 ; 
      RECT 16.68 107.852 16.776 107.948 ; 
      RECT 16.488 72.908 16.584 73.004 ; 
      RECT 16.488 91.692 16.584 91.788 ; 
      RECT 16.488 107.468 16.584 107.564 ; 
      RECT 16.296 72.524 16.392 72.62 ; 
      RECT 16.296 80.94 16.392 81.036 ; 
      RECT 16.296 107.084 16.392 107.18 ; 
      RECT 15.936 91.692 16.032 91.788 ; 
      RECT 15.936 92.076 16.032 92.172 ; 
      RECT 15.268 74.636 15.364 74.732 ; 
      RECT 15.268 89.772 15.364 89.868 ; 
      RECT 13.776 80.94 13.872 81.036 ; 
      RECT 13.776 81.708 13.872 81.804 ; 
  LAYER M5 ; 
      RECT 30.192 77.056 30.288 81.404 ; 
      RECT 29.52 78.774 29.616 82.904 ; 
      RECT 27.024 78.75 27.12 82.08 ; 
      RECT 24.576 81.664 24.672 82.556 ; 
      RECT 24.576 86.464 24.672 87.032 ; 
      RECT 23.712 79.744 23.808 84.092 ; 
      RECT 23.712 85.12 23.808 85.82 ; 
      RECT 22.848 79.36 22.944 84.476 ; 
      RECT 22.848 85.312 22.944 86.072 ; 
      RECT 22.848 86.848 22.944 88.184 ; 
      RECT 22.416 89.728 22.512 91.448 ; 
      RECT 22.416 100.288 22.512 100.856 ; 
      RECT 22.056 75.6 22.152 105.932 ; 
      RECT 21.864 75.6 21.96 105.932 ; 
      RECT 21.672 75.6 21.768 105.932 ; 
      RECT 21.48 75.6 21.576 105.932 ; 
      RECT 21.288 75.6 21.384 105.932 ; 
      RECT 21.096 75.6 21.192 105.932 ; 
      RECT 20.904 75.6 21 105.932 ; 
      RECT 20.712 75.6 20.808 105.932 ; 
      RECT 20.52 75.6 20.616 105.932 ; 
      RECT 19.368 74.552 19.464 106.684 ; 
      RECT 19.176 72.468 19.272 109.784 ; 
      RECT 18.984 72.344 19.08 109.78 ; 
      RECT 18.6 72.528 18.696 109.784 ; 
      RECT 17.832 72.524 17.928 109.596 ; 
      RECT 17.64 72.524 17.736 109.596 ; 
      RECT 17.448 72.524 17.544 109.596 ; 
      RECT 17.256 72.524 17.352 109.596 ; 
      RECT 17.064 72.524 17.16 109.596 ; 
      RECT 16.872 72.408 16.968 109.596 ; 
      RECT 16.68 72.232 16.776 109.6 ; 
      RECT 16.488 72.084 16.584 109.604 ; 
      RECT 16.296 71.844 16.392 109.604 ; 
      RECT 15.936 91.648 16.032 92.216 ; 
      RECT 15.268 74.564 15.364 89.94 ; 
      RECT 13.776 80.896 13.872 81.848 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 38.016 181.296 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 38.016 181.296 ; 
  END 
END srambank_64x4x34_6t122 
