VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_128x4x48_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_128x4x48_6t122 0 0 ;
  SIZE 16.0 BY 60.480000000000004 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.1720 16.4420 1.2200 ;
        RECT 0.0940 2.2520 16.4420 2.3000 ;
        RECT 0.0940 3.3320 16.4420 3.3800 ;
        RECT 0.0940 4.4120 16.4420 4.4600 ;
        RECT 0.0940 5.4920 16.4420 5.5400 ;
        RECT 0.0940 6.5720 16.4420 6.6200 ;
        RECT 0.0940 7.6520 16.4420 7.7000 ;
        RECT 0.0940 8.7320 16.4420 8.7800 ;
        RECT 0.0940 9.8120 16.4420 9.8600 ;
        RECT 0.0940 10.8920 16.4420 10.9400 ;
        RECT 0.0940 11.9720 16.4420 12.0200 ;
        RECT 0.0940 13.0520 16.4420 13.1000 ;
        RECT 0.0940 14.1320 16.4420 14.1800 ;
        RECT 0.0940 15.2120 16.4420 15.2600 ;
        RECT 0.0940 16.2920 16.4420 16.3400 ;
        RECT 0.0940 17.3720 16.4420 17.4200 ;
        RECT 0.0940 18.4520 16.4420 18.5000 ;
        RECT 0.0940 19.5320 16.4420 19.5800 ;
        RECT 0.0940 20.6120 16.4420 20.6600 ;
        RECT 0.0940 21.6920 16.4420 21.7400 ;
        RECT 0.0940 22.7720 16.4420 22.8200 ;
        RECT 0.0940 23.8520 16.4420 23.9000 ;
        RECT 0.0940 24.9320 16.4420 24.9800 ;
        RECT 0.0940 26.0120 16.4420 26.0600 ;
        RECT 3.5640 26.4930 12.9600 26.7090 ;
        RECT 9.1970 29.9970 9.3380 30.0210 ;
        RECT 9.0660 26.2130 9.3290 26.2370 ;
        RECT 7.3980 29.6610 9.1260 29.8770 ;
        RECT 7.3980 32.8290 9.1260 33.0450 ;
        RECT 0.0940 35.2190 16.4420 35.2670 ;
        RECT 0.0940 36.2990 16.4420 36.3470 ;
        RECT 0.0940 37.3790 16.4420 37.4270 ;
        RECT 0.0940 38.4590 16.4420 38.5070 ;
        RECT 0.0940 39.5390 16.4420 39.5870 ;
        RECT 0.0940 40.6190 16.4420 40.6670 ;
        RECT 0.0940 41.6990 16.4420 41.7470 ;
        RECT 0.0940 42.7790 16.4420 42.8270 ;
        RECT 0.0940 43.8590 16.4420 43.9070 ;
        RECT 0.0940 44.9390 16.4420 44.9870 ;
        RECT 0.0940 46.0190 16.4420 46.0670 ;
        RECT 0.0940 47.0990 16.4420 47.1470 ;
        RECT 0.0940 48.1790 16.4420 48.2270 ;
        RECT 0.0940 49.2590 16.4420 49.3070 ;
        RECT 0.0940 50.3390 16.4420 50.3870 ;
        RECT 0.0940 51.4190 16.4420 51.4670 ;
        RECT 0.0940 52.4990 16.4420 52.5470 ;
        RECT 0.0940 53.5790 16.4420 53.6270 ;
        RECT 0.0940 54.6590 16.4420 54.7070 ;
        RECT 0.0940 55.7390 16.4420 55.7870 ;
        RECT 0.0940 56.8190 16.4420 56.8670 ;
        RECT 0.0940 57.8990 16.4420 57.9470 ;
        RECT 0.0940 58.9790 16.4420 59.0270 ;
        RECT 0.0940 60.0590 16.4420 60.1070 ;
      LAYER M3  ;
        RECT 16.3940 0.2165 16.4120 1.3765 ;
        RECT 9.2840 0.2170 9.3020 1.3760 ;
        RECT 7.8800 0.2570 7.9700 1.3710 ;
        RECT 7.2320 0.2170 7.2500 1.3760 ;
        RECT 0.1220 0.2165 0.1400 1.3765 ;
        RECT 16.3940 1.2965 16.4120 2.4565 ;
        RECT 9.2840 1.2970 9.3020 2.4560 ;
        RECT 7.8800 1.3370 7.9700 2.4510 ;
        RECT 7.2320 1.2970 7.2500 2.4560 ;
        RECT 0.1220 1.2965 0.1400 2.4565 ;
        RECT 16.3940 2.3765 16.4120 3.5365 ;
        RECT 9.2840 2.3770 9.3020 3.5360 ;
        RECT 7.8800 2.4170 7.9700 3.5310 ;
        RECT 7.2320 2.3770 7.2500 3.5360 ;
        RECT 0.1220 2.3765 0.1400 3.5365 ;
        RECT 16.3940 3.4565 16.4120 4.6165 ;
        RECT 9.2840 3.4570 9.3020 4.6160 ;
        RECT 7.8800 3.4970 7.9700 4.6110 ;
        RECT 7.2320 3.4570 7.2500 4.6160 ;
        RECT 0.1220 3.4565 0.1400 4.6165 ;
        RECT 16.3940 4.5365 16.4120 5.6965 ;
        RECT 9.2840 4.5370 9.3020 5.6960 ;
        RECT 7.8800 4.5770 7.9700 5.6910 ;
        RECT 7.2320 4.5370 7.2500 5.6960 ;
        RECT 0.1220 4.5365 0.1400 5.6965 ;
        RECT 16.3940 5.6165 16.4120 6.7765 ;
        RECT 9.2840 5.6170 9.3020 6.7760 ;
        RECT 7.8800 5.6570 7.9700 6.7710 ;
        RECT 7.2320 5.6170 7.2500 6.7760 ;
        RECT 0.1220 5.6165 0.1400 6.7765 ;
        RECT 16.3940 6.6965 16.4120 7.8565 ;
        RECT 9.2840 6.6970 9.3020 7.8560 ;
        RECT 7.8800 6.7370 7.9700 7.8510 ;
        RECT 7.2320 6.6970 7.2500 7.8560 ;
        RECT 0.1220 6.6965 0.1400 7.8565 ;
        RECT 16.3940 7.7765 16.4120 8.9365 ;
        RECT 9.2840 7.7770 9.3020 8.9360 ;
        RECT 7.8800 7.8170 7.9700 8.9310 ;
        RECT 7.2320 7.7770 7.2500 8.9360 ;
        RECT 0.1220 7.7765 0.1400 8.9365 ;
        RECT 16.3940 8.8565 16.4120 10.0165 ;
        RECT 9.2840 8.8570 9.3020 10.0160 ;
        RECT 7.8800 8.8970 7.9700 10.0110 ;
        RECT 7.2320 8.8570 7.2500 10.0160 ;
        RECT 0.1220 8.8565 0.1400 10.0165 ;
        RECT 16.3940 9.9365 16.4120 11.0965 ;
        RECT 9.2840 9.9370 9.3020 11.0960 ;
        RECT 7.8800 9.9770 7.9700 11.0910 ;
        RECT 7.2320 9.9370 7.2500 11.0960 ;
        RECT 0.1220 9.9365 0.1400 11.0965 ;
        RECT 16.3940 11.0165 16.4120 12.1765 ;
        RECT 9.2840 11.0170 9.3020 12.1760 ;
        RECT 7.8800 11.0570 7.9700 12.1710 ;
        RECT 7.2320 11.0170 7.2500 12.1760 ;
        RECT 0.1220 11.0165 0.1400 12.1765 ;
        RECT 16.3940 12.0965 16.4120 13.2565 ;
        RECT 9.2840 12.0970 9.3020 13.2560 ;
        RECT 7.8800 12.1370 7.9700 13.2510 ;
        RECT 7.2320 12.0970 7.2500 13.2560 ;
        RECT 0.1220 12.0965 0.1400 13.2565 ;
        RECT 16.3940 13.1765 16.4120 14.3365 ;
        RECT 9.2840 13.1770 9.3020 14.3360 ;
        RECT 7.8800 13.2170 7.9700 14.3310 ;
        RECT 7.2320 13.1770 7.2500 14.3360 ;
        RECT 0.1220 13.1765 0.1400 14.3365 ;
        RECT 16.3940 14.2565 16.4120 15.4165 ;
        RECT 9.2840 14.2570 9.3020 15.4160 ;
        RECT 7.8800 14.2970 7.9700 15.4110 ;
        RECT 7.2320 14.2570 7.2500 15.4160 ;
        RECT 0.1220 14.2565 0.1400 15.4165 ;
        RECT 16.3940 15.3365 16.4120 16.4965 ;
        RECT 9.2840 15.3370 9.3020 16.4960 ;
        RECT 7.8800 15.3770 7.9700 16.4910 ;
        RECT 7.2320 15.3370 7.2500 16.4960 ;
        RECT 0.1220 15.3365 0.1400 16.4965 ;
        RECT 16.3940 16.4165 16.4120 17.5765 ;
        RECT 9.2840 16.4170 9.3020 17.5760 ;
        RECT 7.8800 16.4570 7.9700 17.5710 ;
        RECT 7.2320 16.4170 7.2500 17.5760 ;
        RECT 0.1220 16.4165 0.1400 17.5765 ;
        RECT 16.3940 17.4965 16.4120 18.6565 ;
        RECT 9.2840 17.4970 9.3020 18.6560 ;
        RECT 7.8800 17.5370 7.9700 18.6510 ;
        RECT 7.2320 17.4970 7.2500 18.6560 ;
        RECT 0.1220 17.4965 0.1400 18.6565 ;
        RECT 16.3940 18.5765 16.4120 19.7365 ;
        RECT 9.2840 18.5770 9.3020 19.7360 ;
        RECT 7.8800 18.6170 7.9700 19.7310 ;
        RECT 7.2320 18.5770 7.2500 19.7360 ;
        RECT 0.1220 18.5765 0.1400 19.7365 ;
        RECT 16.3940 19.6565 16.4120 20.8165 ;
        RECT 9.2840 19.6570 9.3020 20.8160 ;
        RECT 7.8800 19.6970 7.9700 20.8110 ;
        RECT 7.2320 19.6570 7.2500 20.8160 ;
        RECT 0.1220 19.6565 0.1400 20.8165 ;
        RECT 16.3940 20.7365 16.4120 21.8965 ;
        RECT 9.2840 20.7370 9.3020 21.8960 ;
        RECT 7.8800 20.7770 7.9700 21.8910 ;
        RECT 7.2320 20.7370 7.2500 21.8960 ;
        RECT 0.1220 20.7365 0.1400 21.8965 ;
        RECT 16.3940 21.8165 16.4120 22.9765 ;
        RECT 9.2840 21.8170 9.3020 22.9760 ;
        RECT 7.8800 21.8570 7.9700 22.9710 ;
        RECT 7.2320 21.8170 7.2500 22.9760 ;
        RECT 0.1220 21.8165 0.1400 22.9765 ;
        RECT 16.3940 22.8965 16.4120 24.0565 ;
        RECT 9.2840 22.8970 9.3020 24.0560 ;
        RECT 7.8800 22.9370 7.9700 24.0510 ;
        RECT 7.2320 22.8970 7.2500 24.0560 ;
        RECT 0.1220 22.8965 0.1400 24.0565 ;
        RECT 16.3940 23.9765 16.4120 25.1365 ;
        RECT 9.2840 23.9770 9.3020 25.1360 ;
        RECT 7.8800 24.0170 7.9700 25.1310 ;
        RECT 7.2320 23.9770 7.2500 25.1360 ;
        RECT 0.1220 23.9765 0.1400 25.1365 ;
        RECT 16.3940 25.0565 16.4120 26.2165 ;
        RECT 9.2840 25.0570 9.3020 26.2160 ;
        RECT 7.8800 25.0970 7.9700 26.2110 ;
        RECT 7.2320 25.0570 7.2500 26.2160 ;
        RECT 0.1220 25.0565 0.1400 26.2165 ;
        RECT 16.3890 26.1305 16.4070 34.3375 ;
        RECT 9.2970 29.9500 9.3150 34.2985 ;
        RECT 9.2790 26.1635 9.2970 26.3015 ;
        RECT 7.9110 26.4540 8.1450 34.0370 ;
        RECT 7.8750 33.9540 7.9650 34.3300 ;
        RECT 7.8750 26.1700 7.9650 26.5460 ;
        RECT 0.1170 26.1305 0.1350 34.3375 ;
        RECT 16.3940 34.2635 16.4120 35.4235 ;
        RECT 9.2840 34.2640 9.3020 35.4230 ;
        RECT 7.8800 34.3040 7.9700 35.4180 ;
        RECT 7.2320 34.2640 7.2500 35.4230 ;
        RECT 0.1220 34.2635 0.1400 35.4235 ;
        RECT 16.3940 35.3435 16.4120 36.5035 ;
        RECT 9.2840 35.3440 9.3020 36.5030 ;
        RECT 7.8800 35.3840 7.9700 36.4980 ;
        RECT 7.2320 35.3440 7.2500 36.5030 ;
        RECT 0.1220 35.3435 0.1400 36.5035 ;
        RECT 16.3940 36.4235 16.4120 37.5835 ;
        RECT 9.2840 36.4240 9.3020 37.5830 ;
        RECT 7.8800 36.4640 7.9700 37.5780 ;
        RECT 7.2320 36.4240 7.2500 37.5830 ;
        RECT 0.1220 36.4235 0.1400 37.5835 ;
        RECT 16.3940 37.5035 16.4120 38.6635 ;
        RECT 9.2840 37.5040 9.3020 38.6630 ;
        RECT 7.8800 37.5440 7.9700 38.6580 ;
        RECT 7.2320 37.5040 7.2500 38.6630 ;
        RECT 0.1220 37.5035 0.1400 38.6635 ;
        RECT 16.3940 38.5835 16.4120 39.7435 ;
        RECT 9.2840 38.5840 9.3020 39.7430 ;
        RECT 7.8800 38.6240 7.9700 39.7380 ;
        RECT 7.2320 38.5840 7.2500 39.7430 ;
        RECT 0.1220 38.5835 0.1400 39.7435 ;
        RECT 16.3940 39.6635 16.4120 40.8235 ;
        RECT 9.2840 39.6640 9.3020 40.8230 ;
        RECT 7.8800 39.7040 7.9700 40.8180 ;
        RECT 7.2320 39.6640 7.2500 40.8230 ;
        RECT 0.1220 39.6635 0.1400 40.8235 ;
        RECT 16.3940 40.7435 16.4120 41.9035 ;
        RECT 9.2840 40.7440 9.3020 41.9030 ;
        RECT 7.8800 40.7840 7.9700 41.8980 ;
        RECT 7.2320 40.7440 7.2500 41.9030 ;
        RECT 0.1220 40.7435 0.1400 41.9035 ;
        RECT 16.3940 41.8235 16.4120 42.9835 ;
        RECT 9.2840 41.8240 9.3020 42.9830 ;
        RECT 7.8800 41.8640 7.9700 42.9780 ;
        RECT 7.2320 41.8240 7.2500 42.9830 ;
        RECT 0.1220 41.8235 0.1400 42.9835 ;
        RECT 16.3940 42.9035 16.4120 44.0635 ;
        RECT 9.2840 42.9040 9.3020 44.0630 ;
        RECT 7.8800 42.9440 7.9700 44.0580 ;
        RECT 7.2320 42.9040 7.2500 44.0630 ;
        RECT 0.1220 42.9035 0.1400 44.0635 ;
        RECT 16.3940 43.9835 16.4120 45.1435 ;
        RECT 9.2840 43.9840 9.3020 45.1430 ;
        RECT 7.8800 44.0240 7.9700 45.1380 ;
        RECT 7.2320 43.9840 7.2500 45.1430 ;
        RECT 0.1220 43.9835 0.1400 45.1435 ;
        RECT 16.3940 45.0635 16.4120 46.2235 ;
        RECT 9.2840 45.0640 9.3020 46.2230 ;
        RECT 7.8800 45.1040 7.9700 46.2180 ;
        RECT 7.2320 45.0640 7.2500 46.2230 ;
        RECT 0.1220 45.0635 0.1400 46.2235 ;
        RECT 16.3940 46.1435 16.4120 47.3035 ;
        RECT 9.2840 46.1440 9.3020 47.3030 ;
        RECT 7.8800 46.1840 7.9700 47.2980 ;
        RECT 7.2320 46.1440 7.2500 47.3030 ;
        RECT 0.1220 46.1435 0.1400 47.3035 ;
        RECT 16.3940 47.2235 16.4120 48.3835 ;
        RECT 9.2840 47.2240 9.3020 48.3830 ;
        RECT 7.8800 47.2640 7.9700 48.3780 ;
        RECT 7.2320 47.2240 7.2500 48.3830 ;
        RECT 0.1220 47.2235 0.1400 48.3835 ;
        RECT 16.3940 48.3035 16.4120 49.4635 ;
        RECT 9.2840 48.3040 9.3020 49.4630 ;
        RECT 7.8800 48.3440 7.9700 49.4580 ;
        RECT 7.2320 48.3040 7.2500 49.4630 ;
        RECT 0.1220 48.3035 0.1400 49.4635 ;
        RECT 16.3940 49.3835 16.4120 50.5435 ;
        RECT 9.2840 49.3840 9.3020 50.5430 ;
        RECT 7.8800 49.4240 7.9700 50.5380 ;
        RECT 7.2320 49.3840 7.2500 50.5430 ;
        RECT 0.1220 49.3835 0.1400 50.5435 ;
        RECT 16.3940 50.4635 16.4120 51.6235 ;
        RECT 9.2840 50.4640 9.3020 51.6230 ;
        RECT 7.8800 50.5040 7.9700 51.6180 ;
        RECT 7.2320 50.4640 7.2500 51.6230 ;
        RECT 0.1220 50.4635 0.1400 51.6235 ;
        RECT 16.3940 51.5435 16.4120 52.7035 ;
        RECT 9.2840 51.5440 9.3020 52.7030 ;
        RECT 7.8800 51.5840 7.9700 52.6980 ;
        RECT 7.2320 51.5440 7.2500 52.7030 ;
        RECT 0.1220 51.5435 0.1400 52.7035 ;
        RECT 16.3940 52.6235 16.4120 53.7835 ;
        RECT 9.2840 52.6240 9.3020 53.7830 ;
        RECT 7.8800 52.6640 7.9700 53.7780 ;
        RECT 7.2320 52.6240 7.2500 53.7830 ;
        RECT 0.1220 52.6235 0.1400 53.7835 ;
        RECT 16.3940 53.7035 16.4120 54.8635 ;
        RECT 9.2840 53.7040 9.3020 54.8630 ;
        RECT 7.8800 53.7440 7.9700 54.8580 ;
        RECT 7.2320 53.7040 7.2500 54.8630 ;
        RECT 0.1220 53.7035 0.1400 54.8635 ;
        RECT 16.3940 54.7835 16.4120 55.9435 ;
        RECT 9.2840 54.7840 9.3020 55.9430 ;
        RECT 7.8800 54.8240 7.9700 55.9380 ;
        RECT 7.2320 54.7840 7.2500 55.9430 ;
        RECT 0.1220 54.7835 0.1400 55.9435 ;
        RECT 16.3940 55.8635 16.4120 57.0235 ;
        RECT 9.2840 55.8640 9.3020 57.0230 ;
        RECT 7.8800 55.9040 7.9700 57.0180 ;
        RECT 7.2320 55.8640 7.2500 57.0230 ;
        RECT 0.1220 55.8635 0.1400 57.0235 ;
        RECT 16.3940 56.9435 16.4120 58.1035 ;
        RECT 9.2840 56.9440 9.3020 58.1030 ;
        RECT 7.8800 56.9840 7.9700 58.0980 ;
        RECT 7.2320 56.9440 7.2500 58.1030 ;
        RECT 0.1220 56.9435 0.1400 58.1035 ;
        RECT 16.3940 58.0235 16.4120 59.1835 ;
        RECT 9.2840 58.0240 9.3020 59.1830 ;
        RECT 7.8800 58.0640 7.9700 59.1780 ;
        RECT 7.2320 58.0240 7.2500 59.1830 ;
        RECT 0.1220 58.0235 0.1400 59.1835 ;
        RECT 16.3940 59.1035 16.4120 60.2635 ;
        RECT 9.2840 59.1040 9.3020 60.2630 ;
        RECT 7.8800 59.1440 7.9700 60.2580 ;
        RECT 7.2320 59.1040 7.2500 60.2630 ;
        RECT 0.1220 59.1035 0.1400 60.2635 ;
      LAYER V3  ;
        RECT 0.1220 1.1720 0.1400 1.2200 ;
        RECT 7.2320 1.1720 7.2500 1.2200 ;
        RECT 7.8800 1.1720 7.9700 1.2200 ;
        RECT 9.2840 1.1720 9.3020 1.2200 ;
        RECT 16.3940 1.1720 16.4120 1.2200 ;
        RECT 0.1220 2.2520 0.1400 2.3000 ;
        RECT 7.2320 2.2520 7.2500 2.3000 ;
        RECT 7.8800 2.2520 7.9700 2.3000 ;
        RECT 9.2840 2.2520 9.3020 2.3000 ;
        RECT 16.3940 2.2520 16.4120 2.3000 ;
        RECT 0.1220 3.3320 0.1400 3.3800 ;
        RECT 7.2320 3.3320 7.2500 3.3800 ;
        RECT 7.8800 3.3320 7.9700 3.3800 ;
        RECT 9.2840 3.3320 9.3020 3.3800 ;
        RECT 16.3940 3.3320 16.4120 3.3800 ;
        RECT 0.1220 4.4120 0.1400 4.4600 ;
        RECT 7.2320 4.4120 7.2500 4.4600 ;
        RECT 7.8800 4.4120 7.9700 4.4600 ;
        RECT 9.2840 4.4120 9.3020 4.4600 ;
        RECT 16.3940 4.4120 16.4120 4.4600 ;
        RECT 0.1220 5.4920 0.1400 5.5400 ;
        RECT 7.2320 5.4920 7.2500 5.5400 ;
        RECT 7.8800 5.4920 7.9700 5.5400 ;
        RECT 9.2840 5.4920 9.3020 5.5400 ;
        RECT 16.3940 5.4920 16.4120 5.5400 ;
        RECT 0.1220 6.5720 0.1400 6.6200 ;
        RECT 7.2320 6.5720 7.2500 6.6200 ;
        RECT 7.8800 6.5720 7.9700 6.6200 ;
        RECT 9.2840 6.5720 9.3020 6.6200 ;
        RECT 16.3940 6.5720 16.4120 6.6200 ;
        RECT 0.1220 7.6520 0.1400 7.7000 ;
        RECT 7.2320 7.6520 7.2500 7.7000 ;
        RECT 7.8800 7.6520 7.9700 7.7000 ;
        RECT 9.2840 7.6520 9.3020 7.7000 ;
        RECT 16.3940 7.6520 16.4120 7.7000 ;
        RECT 0.1220 8.7320 0.1400 8.7800 ;
        RECT 7.2320 8.7320 7.2500 8.7800 ;
        RECT 7.8800 8.7320 7.9700 8.7800 ;
        RECT 9.2840 8.7320 9.3020 8.7800 ;
        RECT 16.3940 8.7320 16.4120 8.7800 ;
        RECT 0.1220 9.8120 0.1400 9.8600 ;
        RECT 7.2320 9.8120 7.2500 9.8600 ;
        RECT 7.8800 9.8120 7.9700 9.8600 ;
        RECT 9.2840 9.8120 9.3020 9.8600 ;
        RECT 16.3940 9.8120 16.4120 9.8600 ;
        RECT 0.1220 10.8920 0.1400 10.9400 ;
        RECT 7.2320 10.8920 7.2500 10.9400 ;
        RECT 7.8800 10.8920 7.9700 10.9400 ;
        RECT 9.2840 10.8920 9.3020 10.9400 ;
        RECT 16.3940 10.8920 16.4120 10.9400 ;
        RECT 0.1220 11.9720 0.1400 12.0200 ;
        RECT 7.2320 11.9720 7.2500 12.0200 ;
        RECT 7.8800 11.9720 7.9700 12.0200 ;
        RECT 9.2840 11.9720 9.3020 12.0200 ;
        RECT 16.3940 11.9720 16.4120 12.0200 ;
        RECT 0.1220 13.0520 0.1400 13.1000 ;
        RECT 7.2320 13.0520 7.2500 13.1000 ;
        RECT 7.8800 13.0520 7.9700 13.1000 ;
        RECT 9.2840 13.0520 9.3020 13.1000 ;
        RECT 16.3940 13.0520 16.4120 13.1000 ;
        RECT 0.1220 14.1320 0.1400 14.1800 ;
        RECT 7.2320 14.1320 7.2500 14.1800 ;
        RECT 7.8800 14.1320 7.9700 14.1800 ;
        RECT 9.2840 14.1320 9.3020 14.1800 ;
        RECT 16.3940 14.1320 16.4120 14.1800 ;
        RECT 0.1220 15.2120 0.1400 15.2600 ;
        RECT 7.2320 15.2120 7.2500 15.2600 ;
        RECT 7.8800 15.2120 7.9700 15.2600 ;
        RECT 9.2840 15.2120 9.3020 15.2600 ;
        RECT 16.3940 15.2120 16.4120 15.2600 ;
        RECT 0.1220 16.2920 0.1400 16.3400 ;
        RECT 7.2320 16.2920 7.2500 16.3400 ;
        RECT 7.8800 16.2920 7.9700 16.3400 ;
        RECT 9.2840 16.2920 9.3020 16.3400 ;
        RECT 16.3940 16.2920 16.4120 16.3400 ;
        RECT 0.1220 17.3720 0.1400 17.4200 ;
        RECT 7.2320 17.3720 7.2500 17.4200 ;
        RECT 7.8800 17.3720 7.9700 17.4200 ;
        RECT 9.2840 17.3720 9.3020 17.4200 ;
        RECT 16.3940 17.3720 16.4120 17.4200 ;
        RECT 0.1220 18.4520 0.1400 18.5000 ;
        RECT 7.2320 18.4520 7.2500 18.5000 ;
        RECT 7.8800 18.4520 7.9700 18.5000 ;
        RECT 9.2840 18.4520 9.3020 18.5000 ;
        RECT 16.3940 18.4520 16.4120 18.5000 ;
        RECT 0.1220 19.5320 0.1400 19.5800 ;
        RECT 7.2320 19.5320 7.2500 19.5800 ;
        RECT 7.8800 19.5320 7.9700 19.5800 ;
        RECT 9.2840 19.5320 9.3020 19.5800 ;
        RECT 16.3940 19.5320 16.4120 19.5800 ;
        RECT 0.1220 20.6120 0.1400 20.6600 ;
        RECT 7.2320 20.6120 7.2500 20.6600 ;
        RECT 7.8800 20.6120 7.9700 20.6600 ;
        RECT 9.2840 20.6120 9.3020 20.6600 ;
        RECT 16.3940 20.6120 16.4120 20.6600 ;
        RECT 0.1220 21.6920 0.1400 21.7400 ;
        RECT 7.2320 21.6920 7.2500 21.7400 ;
        RECT 7.8800 21.6920 7.9700 21.7400 ;
        RECT 9.2840 21.6920 9.3020 21.7400 ;
        RECT 16.3940 21.6920 16.4120 21.7400 ;
        RECT 0.1220 22.7720 0.1400 22.8200 ;
        RECT 7.2320 22.7720 7.2500 22.8200 ;
        RECT 7.8800 22.7720 7.9700 22.8200 ;
        RECT 9.2840 22.7720 9.3020 22.8200 ;
        RECT 16.3940 22.7720 16.4120 22.8200 ;
        RECT 0.1220 23.8520 0.1400 23.9000 ;
        RECT 7.2320 23.8520 7.2500 23.9000 ;
        RECT 7.8800 23.8520 7.9700 23.9000 ;
        RECT 9.2840 23.8520 9.3020 23.9000 ;
        RECT 16.3940 23.8520 16.4120 23.9000 ;
        RECT 0.1220 24.9320 0.1400 24.9800 ;
        RECT 7.2320 24.9320 7.2500 24.9800 ;
        RECT 7.8800 24.9320 7.9700 24.9800 ;
        RECT 9.2840 24.9320 9.3020 24.9800 ;
        RECT 16.3940 24.9320 16.4120 24.9800 ;
        RECT 0.1220 26.0120 0.1400 26.0600 ;
        RECT 7.2320 26.0120 7.2500 26.0600 ;
        RECT 7.8800 26.0120 7.9700 26.0600 ;
        RECT 9.2840 26.0120 9.3020 26.0600 ;
        RECT 16.3940 26.0120 16.4120 26.0600 ;
        RECT 7.9150 32.8290 7.9330 33.0450 ;
        RECT 7.9150 29.6610 7.9330 29.8770 ;
        RECT 7.9150 26.4930 7.9330 26.7090 ;
        RECT 7.9670 32.8290 7.9850 33.0450 ;
        RECT 7.9670 29.6610 7.9850 29.8770 ;
        RECT 7.9670 26.4930 7.9850 26.7090 ;
        RECT 8.0190 32.8290 8.0370 33.0450 ;
        RECT 8.0190 29.6610 8.0370 29.8770 ;
        RECT 8.0190 26.4930 8.0370 26.7090 ;
        RECT 8.0710 32.8290 8.0890 33.0450 ;
        RECT 8.0710 29.6610 8.0890 29.8770 ;
        RECT 8.0710 26.4930 8.0890 26.7090 ;
        RECT 8.1230 32.8290 8.1410 33.0450 ;
        RECT 8.1230 29.6610 8.1410 29.8770 ;
        RECT 8.1230 26.4930 8.1410 26.7090 ;
        RECT 9.2790 26.2130 9.2970 26.2370 ;
        RECT 9.2970 29.9970 9.3150 30.0210 ;
        RECT 0.1220 35.2190 0.1400 35.2670 ;
        RECT 7.2320 35.2190 7.2500 35.2670 ;
        RECT 7.8800 35.2190 7.9700 35.2670 ;
        RECT 9.2840 35.2190 9.3020 35.2670 ;
        RECT 16.3940 35.2190 16.4120 35.2670 ;
        RECT 0.1220 36.2990 0.1400 36.3470 ;
        RECT 7.2320 36.2990 7.2500 36.3470 ;
        RECT 7.8800 36.2990 7.9700 36.3470 ;
        RECT 9.2840 36.2990 9.3020 36.3470 ;
        RECT 16.3940 36.2990 16.4120 36.3470 ;
        RECT 0.1220 37.3790 0.1400 37.4270 ;
        RECT 7.2320 37.3790 7.2500 37.4270 ;
        RECT 7.8800 37.3790 7.9700 37.4270 ;
        RECT 9.2840 37.3790 9.3020 37.4270 ;
        RECT 16.3940 37.3790 16.4120 37.4270 ;
        RECT 0.1220 38.4590 0.1400 38.5070 ;
        RECT 7.2320 38.4590 7.2500 38.5070 ;
        RECT 7.8800 38.4590 7.9700 38.5070 ;
        RECT 9.2840 38.4590 9.3020 38.5070 ;
        RECT 16.3940 38.4590 16.4120 38.5070 ;
        RECT 0.1220 39.5390 0.1400 39.5870 ;
        RECT 7.2320 39.5390 7.2500 39.5870 ;
        RECT 7.8800 39.5390 7.9700 39.5870 ;
        RECT 9.2840 39.5390 9.3020 39.5870 ;
        RECT 16.3940 39.5390 16.4120 39.5870 ;
        RECT 0.1220 40.6190 0.1400 40.6670 ;
        RECT 7.2320 40.6190 7.2500 40.6670 ;
        RECT 7.8800 40.6190 7.9700 40.6670 ;
        RECT 9.2840 40.6190 9.3020 40.6670 ;
        RECT 16.3940 40.6190 16.4120 40.6670 ;
        RECT 0.1220 41.6990 0.1400 41.7470 ;
        RECT 7.2320 41.6990 7.2500 41.7470 ;
        RECT 7.8800 41.6990 7.9700 41.7470 ;
        RECT 9.2840 41.6990 9.3020 41.7470 ;
        RECT 16.3940 41.6990 16.4120 41.7470 ;
        RECT 0.1220 42.7790 0.1400 42.8270 ;
        RECT 7.2320 42.7790 7.2500 42.8270 ;
        RECT 7.8800 42.7790 7.9700 42.8270 ;
        RECT 9.2840 42.7790 9.3020 42.8270 ;
        RECT 16.3940 42.7790 16.4120 42.8270 ;
        RECT 0.1220 43.8590 0.1400 43.9070 ;
        RECT 7.2320 43.8590 7.2500 43.9070 ;
        RECT 7.8800 43.8590 7.9700 43.9070 ;
        RECT 9.2840 43.8590 9.3020 43.9070 ;
        RECT 16.3940 43.8590 16.4120 43.9070 ;
        RECT 0.1220 44.9390 0.1400 44.9870 ;
        RECT 7.2320 44.9390 7.2500 44.9870 ;
        RECT 7.8800 44.9390 7.9700 44.9870 ;
        RECT 9.2840 44.9390 9.3020 44.9870 ;
        RECT 16.3940 44.9390 16.4120 44.9870 ;
        RECT 0.1220 46.0190 0.1400 46.0670 ;
        RECT 7.2320 46.0190 7.2500 46.0670 ;
        RECT 7.8800 46.0190 7.9700 46.0670 ;
        RECT 9.2840 46.0190 9.3020 46.0670 ;
        RECT 16.3940 46.0190 16.4120 46.0670 ;
        RECT 0.1220 47.0990 0.1400 47.1470 ;
        RECT 7.2320 47.0990 7.2500 47.1470 ;
        RECT 7.8800 47.0990 7.9700 47.1470 ;
        RECT 9.2840 47.0990 9.3020 47.1470 ;
        RECT 16.3940 47.0990 16.4120 47.1470 ;
        RECT 0.1220 48.1790 0.1400 48.2270 ;
        RECT 7.2320 48.1790 7.2500 48.2270 ;
        RECT 7.8800 48.1790 7.9700 48.2270 ;
        RECT 9.2840 48.1790 9.3020 48.2270 ;
        RECT 16.3940 48.1790 16.4120 48.2270 ;
        RECT 0.1220 49.2590 0.1400 49.3070 ;
        RECT 7.2320 49.2590 7.2500 49.3070 ;
        RECT 7.8800 49.2590 7.9700 49.3070 ;
        RECT 9.2840 49.2590 9.3020 49.3070 ;
        RECT 16.3940 49.2590 16.4120 49.3070 ;
        RECT 0.1220 50.3390 0.1400 50.3870 ;
        RECT 7.2320 50.3390 7.2500 50.3870 ;
        RECT 7.8800 50.3390 7.9700 50.3870 ;
        RECT 9.2840 50.3390 9.3020 50.3870 ;
        RECT 16.3940 50.3390 16.4120 50.3870 ;
        RECT 0.1220 51.4190 0.1400 51.4670 ;
        RECT 7.2320 51.4190 7.2500 51.4670 ;
        RECT 7.8800 51.4190 7.9700 51.4670 ;
        RECT 9.2840 51.4190 9.3020 51.4670 ;
        RECT 16.3940 51.4190 16.4120 51.4670 ;
        RECT 0.1220 52.4990 0.1400 52.5470 ;
        RECT 7.2320 52.4990 7.2500 52.5470 ;
        RECT 7.8800 52.4990 7.9700 52.5470 ;
        RECT 9.2840 52.4990 9.3020 52.5470 ;
        RECT 16.3940 52.4990 16.4120 52.5470 ;
        RECT 0.1220 53.5790 0.1400 53.6270 ;
        RECT 7.2320 53.5790 7.2500 53.6270 ;
        RECT 7.8800 53.5790 7.9700 53.6270 ;
        RECT 9.2840 53.5790 9.3020 53.6270 ;
        RECT 16.3940 53.5790 16.4120 53.6270 ;
        RECT 0.1220 54.6590 0.1400 54.7070 ;
        RECT 7.2320 54.6590 7.2500 54.7070 ;
        RECT 7.8800 54.6590 7.9700 54.7070 ;
        RECT 9.2840 54.6590 9.3020 54.7070 ;
        RECT 16.3940 54.6590 16.4120 54.7070 ;
        RECT 0.1220 55.7390 0.1400 55.7870 ;
        RECT 7.2320 55.7390 7.2500 55.7870 ;
        RECT 7.8800 55.7390 7.9700 55.7870 ;
        RECT 9.2840 55.7390 9.3020 55.7870 ;
        RECT 16.3940 55.7390 16.4120 55.7870 ;
        RECT 0.1220 56.8190 0.1400 56.8670 ;
        RECT 7.2320 56.8190 7.2500 56.8670 ;
        RECT 7.8800 56.8190 7.9700 56.8670 ;
        RECT 9.2840 56.8190 9.3020 56.8670 ;
        RECT 16.3940 56.8190 16.4120 56.8670 ;
        RECT 0.1220 57.8990 0.1400 57.9470 ;
        RECT 7.2320 57.8990 7.2500 57.9470 ;
        RECT 7.8800 57.8990 7.9700 57.9470 ;
        RECT 9.2840 57.8990 9.3020 57.9470 ;
        RECT 16.3940 57.8990 16.4120 57.9470 ;
        RECT 0.1220 58.9790 0.1400 59.0270 ;
        RECT 7.2320 58.9790 7.2500 59.0270 ;
        RECT 7.8800 58.9790 7.9700 59.0270 ;
        RECT 9.2840 58.9790 9.3020 59.0270 ;
        RECT 16.3940 58.9790 16.4120 59.0270 ;
        RECT 0.1220 60.0590 0.1400 60.1070 ;
        RECT 7.2320 60.0590 7.2500 60.1070 ;
        RECT 7.8800 60.0590 7.9700 60.1070 ;
        RECT 9.2840 60.0590 9.3020 60.1070 ;
        RECT 16.3940 60.0590 16.4120 60.1070 ;
      LAYER M5  ;
        RECT 9.2160 26.1950 9.2400 30.0390 ;
      LAYER V4  ;
        RECT 9.2160 29.9970 9.2400 30.0210 ;
        RECT 9.2160 26.4930 9.2400 26.7090 ;
        RECT 9.2160 26.2130 9.2400 26.2370 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.0940 1.0760 16.4370 1.1240 ;
        RECT 0.0940 2.1560 16.4370 2.2040 ;
        RECT 0.0940 3.2360 16.4370 3.2840 ;
        RECT 0.0940 4.3160 16.4370 4.3640 ;
        RECT 0.0940 5.3960 16.4370 5.4440 ;
        RECT 0.0940 6.4760 16.4370 6.5240 ;
        RECT 0.0940 7.5560 16.4370 7.6040 ;
        RECT 0.0940 8.6360 16.4370 8.6840 ;
        RECT 0.0940 9.7160 16.4370 9.7640 ;
        RECT 0.0940 10.7960 16.4370 10.8440 ;
        RECT 0.0940 11.8760 16.4370 11.9240 ;
        RECT 0.0940 12.9560 16.4370 13.0040 ;
        RECT 0.0940 14.0360 16.4370 14.0840 ;
        RECT 0.0940 15.1160 16.4370 15.1640 ;
        RECT 0.0940 16.1960 16.4370 16.2440 ;
        RECT 0.0940 17.2760 16.4370 17.3240 ;
        RECT 0.0940 18.3560 16.4370 18.4040 ;
        RECT 0.0940 19.4360 16.4370 19.4840 ;
        RECT 0.0940 20.5160 16.4370 20.5640 ;
        RECT 0.0940 21.5960 16.4370 21.6440 ;
        RECT 0.0940 22.6760 16.4370 22.7240 ;
        RECT 0.0940 23.7560 16.4370 23.8040 ;
        RECT 0.0940 24.8360 16.4370 24.8840 ;
        RECT 0.0940 25.9160 16.4370 25.9640 ;
        RECT 3.5640 26.9250 12.9600 27.1410 ;
        RECT 7.3980 30.0930 9.1260 30.3090 ;
        RECT 7.3980 33.2610 9.1260 33.4770 ;
        RECT 0.0940 35.1230 16.4370 35.1710 ;
        RECT 0.0940 36.2030 16.4370 36.2510 ;
        RECT 0.0940 37.2830 16.4370 37.3310 ;
        RECT 0.0940 38.3630 16.4370 38.4110 ;
        RECT 0.0940 39.4430 16.4370 39.4910 ;
        RECT 0.0940 40.5230 16.4370 40.5710 ;
        RECT 0.0940 41.6030 16.4370 41.6510 ;
        RECT 0.0940 42.6830 16.4370 42.7310 ;
        RECT 0.0940 43.7630 16.4370 43.8110 ;
        RECT 0.0940 44.8430 16.4370 44.8910 ;
        RECT 0.0940 45.9230 16.4370 45.9710 ;
        RECT 0.0940 47.0030 16.4370 47.0510 ;
        RECT 0.0940 48.0830 16.4370 48.1310 ;
        RECT 0.0940 49.1630 16.4370 49.2110 ;
        RECT 0.0940 50.2430 16.4370 50.2910 ;
        RECT 0.0940 51.3230 16.4370 51.3710 ;
        RECT 0.0940 52.4030 16.4370 52.4510 ;
        RECT 0.0940 53.4830 16.4370 53.5310 ;
        RECT 0.0940 54.5630 16.4370 54.6110 ;
        RECT 0.0940 55.6430 16.4370 55.6910 ;
        RECT 0.0940 56.7230 16.4370 56.7710 ;
        RECT 0.0940 57.8030 16.4370 57.8510 ;
        RECT 0.0940 58.8830 16.4370 58.9310 ;
        RECT 0.0940 59.9630 16.4370 60.0110 ;
      LAYER M3  ;
        RECT 16.3580 0.2165 16.3760 1.3765 ;
        RECT 9.3380 0.2165 9.3560 1.3765 ;
        RECT 8.5730 0.2530 8.6090 1.3670 ;
        RECT 8.4200 0.2530 8.4470 1.3670 ;
        RECT 7.1780 0.2165 7.1960 1.3765 ;
        RECT 0.1580 0.2165 0.1760 1.3765 ;
        RECT 16.3580 1.2965 16.3760 2.4565 ;
        RECT 9.3380 1.2965 9.3560 2.4565 ;
        RECT 8.5730 1.3330 8.6090 2.4470 ;
        RECT 8.4200 1.3330 8.4470 2.4470 ;
        RECT 7.1780 1.2965 7.1960 2.4565 ;
        RECT 0.1580 1.2965 0.1760 2.4565 ;
        RECT 16.3580 2.3765 16.3760 3.5365 ;
        RECT 9.3380 2.3765 9.3560 3.5365 ;
        RECT 8.5730 2.4130 8.6090 3.5270 ;
        RECT 8.4200 2.4130 8.4470 3.5270 ;
        RECT 7.1780 2.3765 7.1960 3.5365 ;
        RECT 0.1580 2.3765 0.1760 3.5365 ;
        RECT 16.3580 3.4565 16.3760 4.6165 ;
        RECT 9.3380 3.4565 9.3560 4.6165 ;
        RECT 8.5730 3.4930 8.6090 4.6070 ;
        RECT 8.4200 3.4930 8.4470 4.6070 ;
        RECT 7.1780 3.4565 7.1960 4.6165 ;
        RECT 0.1580 3.4565 0.1760 4.6165 ;
        RECT 16.3580 4.5365 16.3760 5.6965 ;
        RECT 9.3380 4.5365 9.3560 5.6965 ;
        RECT 8.5730 4.5730 8.6090 5.6870 ;
        RECT 8.4200 4.5730 8.4470 5.6870 ;
        RECT 7.1780 4.5365 7.1960 5.6965 ;
        RECT 0.1580 4.5365 0.1760 5.6965 ;
        RECT 16.3580 5.6165 16.3760 6.7765 ;
        RECT 9.3380 5.6165 9.3560 6.7765 ;
        RECT 8.5730 5.6530 8.6090 6.7670 ;
        RECT 8.4200 5.6530 8.4470 6.7670 ;
        RECT 7.1780 5.6165 7.1960 6.7765 ;
        RECT 0.1580 5.6165 0.1760 6.7765 ;
        RECT 16.3580 6.6965 16.3760 7.8565 ;
        RECT 9.3380 6.6965 9.3560 7.8565 ;
        RECT 8.5730 6.7330 8.6090 7.8470 ;
        RECT 8.4200 6.7330 8.4470 7.8470 ;
        RECT 7.1780 6.6965 7.1960 7.8565 ;
        RECT 0.1580 6.6965 0.1760 7.8565 ;
        RECT 16.3580 7.7765 16.3760 8.9365 ;
        RECT 9.3380 7.7765 9.3560 8.9365 ;
        RECT 8.5730 7.8130 8.6090 8.9270 ;
        RECT 8.4200 7.8130 8.4470 8.9270 ;
        RECT 7.1780 7.7765 7.1960 8.9365 ;
        RECT 0.1580 7.7765 0.1760 8.9365 ;
        RECT 16.3580 8.8565 16.3760 10.0165 ;
        RECT 9.3380 8.8565 9.3560 10.0165 ;
        RECT 8.5730 8.8930 8.6090 10.0070 ;
        RECT 8.4200 8.8930 8.4470 10.0070 ;
        RECT 7.1780 8.8565 7.1960 10.0165 ;
        RECT 0.1580 8.8565 0.1760 10.0165 ;
        RECT 16.3580 9.9365 16.3760 11.0965 ;
        RECT 9.3380 9.9365 9.3560 11.0965 ;
        RECT 8.5730 9.9730 8.6090 11.0870 ;
        RECT 8.4200 9.9730 8.4470 11.0870 ;
        RECT 7.1780 9.9365 7.1960 11.0965 ;
        RECT 0.1580 9.9365 0.1760 11.0965 ;
        RECT 16.3580 11.0165 16.3760 12.1765 ;
        RECT 9.3380 11.0165 9.3560 12.1765 ;
        RECT 8.5730 11.0530 8.6090 12.1670 ;
        RECT 8.4200 11.0530 8.4470 12.1670 ;
        RECT 7.1780 11.0165 7.1960 12.1765 ;
        RECT 0.1580 11.0165 0.1760 12.1765 ;
        RECT 16.3580 12.0965 16.3760 13.2565 ;
        RECT 9.3380 12.0965 9.3560 13.2565 ;
        RECT 8.5730 12.1330 8.6090 13.2470 ;
        RECT 8.4200 12.1330 8.4470 13.2470 ;
        RECT 7.1780 12.0965 7.1960 13.2565 ;
        RECT 0.1580 12.0965 0.1760 13.2565 ;
        RECT 16.3580 13.1765 16.3760 14.3365 ;
        RECT 9.3380 13.1765 9.3560 14.3365 ;
        RECT 8.5730 13.2130 8.6090 14.3270 ;
        RECT 8.4200 13.2130 8.4470 14.3270 ;
        RECT 7.1780 13.1765 7.1960 14.3365 ;
        RECT 0.1580 13.1765 0.1760 14.3365 ;
        RECT 16.3580 14.2565 16.3760 15.4165 ;
        RECT 9.3380 14.2565 9.3560 15.4165 ;
        RECT 8.5730 14.2930 8.6090 15.4070 ;
        RECT 8.4200 14.2930 8.4470 15.4070 ;
        RECT 7.1780 14.2565 7.1960 15.4165 ;
        RECT 0.1580 14.2565 0.1760 15.4165 ;
        RECT 16.3580 15.3365 16.3760 16.4965 ;
        RECT 9.3380 15.3365 9.3560 16.4965 ;
        RECT 8.5730 15.3730 8.6090 16.4870 ;
        RECT 8.4200 15.3730 8.4470 16.4870 ;
        RECT 7.1780 15.3365 7.1960 16.4965 ;
        RECT 0.1580 15.3365 0.1760 16.4965 ;
        RECT 16.3580 16.4165 16.3760 17.5765 ;
        RECT 9.3380 16.4165 9.3560 17.5765 ;
        RECT 8.5730 16.4530 8.6090 17.5670 ;
        RECT 8.4200 16.4530 8.4470 17.5670 ;
        RECT 7.1780 16.4165 7.1960 17.5765 ;
        RECT 0.1580 16.4165 0.1760 17.5765 ;
        RECT 16.3580 17.4965 16.3760 18.6565 ;
        RECT 9.3380 17.4965 9.3560 18.6565 ;
        RECT 8.5730 17.5330 8.6090 18.6470 ;
        RECT 8.4200 17.5330 8.4470 18.6470 ;
        RECT 7.1780 17.4965 7.1960 18.6565 ;
        RECT 0.1580 17.4965 0.1760 18.6565 ;
        RECT 16.3580 18.5765 16.3760 19.7365 ;
        RECT 9.3380 18.5765 9.3560 19.7365 ;
        RECT 8.5730 18.6130 8.6090 19.7270 ;
        RECT 8.4200 18.6130 8.4470 19.7270 ;
        RECT 7.1780 18.5765 7.1960 19.7365 ;
        RECT 0.1580 18.5765 0.1760 19.7365 ;
        RECT 16.3580 19.6565 16.3760 20.8165 ;
        RECT 9.3380 19.6565 9.3560 20.8165 ;
        RECT 8.5730 19.6930 8.6090 20.8070 ;
        RECT 8.4200 19.6930 8.4470 20.8070 ;
        RECT 7.1780 19.6565 7.1960 20.8165 ;
        RECT 0.1580 19.6565 0.1760 20.8165 ;
        RECT 16.3580 20.7365 16.3760 21.8965 ;
        RECT 9.3380 20.7365 9.3560 21.8965 ;
        RECT 8.5730 20.7730 8.6090 21.8870 ;
        RECT 8.4200 20.7730 8.4470 21.8870 ;
        RECT 7.1780 20.7365 7.1960 21.8965 ;
        RECT 0.1580 20.7365 0.1760 21.8965 ;
        RECT 16.3580 21.8165 16.3760 22.9765 ;
        RECT 9.3380 21.8165 9.3560 22.9765 ;
        RECT 8.5730 21.8530 8.6090 22.9670 ;
        RECT 8.4200 21.8530 8.4470 22.9670 ;
        RECT 7.1780 21.8165 7.1960 22.9765 ;
        RECT 0.1580 21.8165 0.1760 22.9765 ;
        RECT 16.3580 22.8965 16.3760 24.0565 ;
        RECT 9.3380 22.8965 9.3560 24.0565 ;
        RECT 8.5730 22.9330 8.6090 24.0470 ;
        RECT 8.4200 22.9330 8.4470 24.0470 ;
        RECT 7.1780 22.8965 7.1960 24.0565 ;
        RECT 0.1580 22.8965 0.1760 24.0565 ;
        RECT 16.3580 23.9765 16.3760 25.1365 ;
        RECT 9.3380 23.9765 9.3560 25.1365 ;
        RECT 8.5730 24.0130 8.6090 25.1270 ;
        RECT 8.4200 24.0130 8.4470 25.1270 ;
        RECT 7.1780 23.9765 7.1960 25.1365 ;
        RECT 0.1580 23.9765 0.1760 25.1365 ;
        RECT 16.3580 25.0565 16.3760 26.2165 ;
        RECT 9.3380 25.0565 9.3560 26.2165 ;
        RECT 8.5730 25.0930 8.6090 26.2070 ;
        RECT 8.4200 25.0930 8.4470 26.2070 ;
        RECT 7.1780 25.0565 7.1960 26.2165 ;
        RECT 0.1580 25.0565 0.1760 26.2165 ;
        RECT 16.3530 26.1305 16.3710 34.3375 ;
        RECT 9.3330 26.1305 9.3510 34.3375 ;
        RECT 8.3790 26.3540 8.6130 34.0370 ;
        RECT 8.5680 26.1745 8.6040 34.2940 ;
        RECT 8.4150 26.1740 8.4420 34.2940 ;
        RECT 7.1730 26.1305 7.1910 34.3375 ;
        RECT 0.1530 26.1305 0.1710 34.3375 ;
        RECT 16.3580 34.2635 16.3760 35.4235 ;
        RECT 9.3380 34.2635 9.3560 35.4235 ;
        RECT 8.5730 34.3000 8.6090 35.4140 ;
        RECT 8.4200 34.3000 8.4470 35.4140 ;
        RECT 7.1780 34.2635 7.1960 35.4235 ;
        RECT 0.1580 34.2635 0.1760 35.4235 ;
        RECT 16.3580 35.3435 16.3760 36.5035 ;
        RECT 9.3380 35.3435 9.3560 36.5035 ;
        RECT 8.5730 35.3800 8.6090 36.4940 ;
        RECT 8.4200 35.3800 8.4470 36.4940 ;
        RECT 7.1780 35.3435 7.1960 36.5035 ;
        RECT 0.1580 35.3435 0.1760 36.5035 ;
        RECT 16.3580 36.4235 16.3760 37.5835 ;
        RECT 9.3380 36.4235 9.3560 37.5835 ;
        RECT 8.5730 36.4600 8.6090 37.5740 ;
        RECT 8.4200 36.4600 8.4470 37.5740 ;
        RECT 7.1780 36.4235 7.1960 37.5835 ;
        RECT 0.1580 36.4235 0.1760 37.5835 ;
        RECT 16.3580 37.5035 16.3760 38.6635 ;
        RECT 9.3380 37.5035 9.3560 38.6635 ;
        RECT 8.5730 37.5400 8.6090 38.6540 ;
        RECT 8.4200 37.5400 8.4470 38.6540 ;
        RECT 7.1780 37.5035 7.1960 38.6635 ;
        RECT 0.1580 37.5035 0.1760 38.6635 ;
        RECT 16.3580 38.5835 16.3760 39.7435 ;
        RECT 9.3380 38.5835 9.3560 39.7435 ;
        RECT 8.5730 38.6200 8.6090 39.7340 ;
        RECT 8.4200 38.6200 8.4470 39.7340 ;
        RECT 7.1780 38.5835 7.1960 39.7435 ;
        RECT 0.1580 38.5835 0.1760 39.7435 ;
        RECT 16.3580 39.6635 16.3760 40.8235 ;
        RECT 9.3380 39.6635 9.3560 40.8235 ;
        RECT 8.5730 39.7000 8.6090 40.8140 ;
        RECT 8.4200 39.7000 8.4470 40.8140 ;
        RECT 7.1780 39.6635 7.1960 40.8235 ;
        RECT 0.1580 39.6635 0.1760 40.8235 ;
        RECT 16.3580 40.7435 16.3760 41.9035 ;
        RECT 9.3380 40.7435 9.3560 41.9035 ;
        RECT 8.5730 40.7800 8.6090 41.8940 ;
        RECT 8.4200 40.7800 8.4470 41.8940 ;
        RECT 7.1780 40.7435 7.1960 41.9035 ;
        RECT 0.1580 40.7435 0.1760 41.9035 ;
        RECT 16.3580 41.8235 16.3760 42.9835 ;
        RECT 9.3380 41.8235 9.3560 42.9835 ;
        RECT 8.5730 41.8600 8.6090 42.9740 ;
        RECT 8.4200 41.8600 8.4470 42.9740 ;
        RECT 7.1780 41.8235 7.1960 42.9835 ;
        RECT 0.1580 41.8235 0.1760 42.9835 ;
        RECT 16.3580 42.9035 16.3760 44.0635 ;
        RECT 9.3380 42.9035 9.3560 44.0635 ;
        RECT 8.5730 42.9400 8.6090 44.0540 ;
        RECT 8.4200 42.9400 8.4470 44.0540 ;
        RECT 7.1780 42.9035 7.1960 44.0635 ;
        RECT 0.1580 42.9035 0.1760 44.0635 ;
        RECT 16.3580 43.9835 16.3760 45.1435 ;
        RECT 9.3380 43.9835 9.3560 45.1435 ;
        RECT 8.5730 44.0200 8.6090 45.1340 ;
        RECT 8.4200 44.0200 8.4470 45.1340 ;
        RECT 7.1780 43.9835 7.1960 45.1435 ;
        RECT 0.1580 43.9835 0.1760 45.1435 ;
        RECT 16.3580 45.0635 16.3760 46.2235 ;
        RECT 9.3380 45.0635 9.3560 46.2235 ;
        RECT 8.5730 45.1000 8.6090 46.2140 ;
        RECT 8.4200 45.1000 8.4470 46.2140 ;
        RECT 7.1780 45.0635 7.1960 46.2235 ;
        RECT 0.1580 45.0635 0.1760 46.2235 ;
        RECT 16.3580 46.1435 16.3760 47.3035 ;
        RECT 9.3380 46.1435 9.3560 47.3035 ;
        RECT 8.5730 46.1800 8.6090 47.2940 ;
        RECT 8.4200 46.1800 8.4470 47.2940 ;
        RECT 7.1780 46.1435 7.1960 47.3035 ;
        RECT 0.1580 46.1435 0.1760 47.3035 ;
        RECT 16.3580 47.2235 16.3760 48.3835 ;
        RECT 9.3380 47.2235 9.3560 48.3835 ;
        RECT 8.5730 47.2600 8.6090 48.3740 ;
        RECT 8.4200 47.2600 8.4470 48.3740 ;
        RECT 7.1780 47.2235 7.1960 48.3835 ;
        RECT 0.1580 47.2235 0.1760 48.3835 ;
        RECT 16.3580 48.3035 16.3760 49.4635 ;
        RECT 9.3380 48.3035 9.3560 49.4635 ;
        RECT 8.5730 48.3400 8.6090 49.4540 ;
        RECT 8.4200 48.3400 8.4470 49.4540 ;
        RECT 7.1780 48.3035 7.1960 49.4635 ;
        RECT 0.1580 48.3035 0.1760 49.4635 ;
        RECT 16.3580 49.3835 16.3760 50.5435 ;
        RECT 9.3380 49.3835 9.3560 50.5435 ;
        RECT 8.5730 49.4200 8.6090 50.5340 ;
        RECT 8.4200 49.4200 8.4470 50.5340 ;
        RECT 7.1780 49.3835 7.1960 50.5435 ;
        RECT 0.1580 49.3835 0.1760 50.5435 ;
        RECT 16.3580 50.4635 16.3760 51.6235 ;
        RECT 9.3380 50.4635 9.3560 51.6235 ;
        RECT 8.5730 50.5000 8.6090 51.6140 ;
        RECT 8.4200 50.5000 8.4470 51.6140 ;
        RECT 7.1780 50.4635 7.1960 51.6235 ;
        RECT 0.1580 50.4635 0.1760 51.6235 ;
        RECT 16.3580 51.5435 16.3760 52.7035 ;
        RECT 9.3380 51.5435 9.3560 52.7035 ;
        RECT 8.5730 51.5800 8.6090 52.6940 ;
        RECT 8.4200 51.5800 8.4470 52.6940 ;
        RECT 7.1780 51.5435 7.1960 52.7035 ;
        RECT 0.1580 51.5435 0.1760 52.7035 ;
        RECT 16.3580 52.6235 16.3760 53.7835 ;
        RECT 9.3380 52.6235 9.3560 53.7835 ;
        RECT 8.5730 52.6600 8.6090 53.7740 ;
        RECT 8.4200 52.6600 8.4470 53.7740 ;
        RECT 7.1780 52.6235 7.1960 53.7835 ;
        RECT 0.1580 52.6235 0.1760 53.7835 ;
        RECT 16.3580 53.7035 16.3760 54.8635 ;
        RECT 9.3380 53.7035 9.3560 54.8635 ;
        RECT 8.5730 53.7400 8.6090 54.8540 ;
        RECT 8.4200 53.7400 8.4470 54.8540 ;
        RECT 7.1780 53.7035 7.1960 54.8635 ;
        RECT 0.1580 53.7035 0.1760 54.8635 ;
        RECT 16.3580 54.7835 16.3760 55.9435 ;
        RECT 9.3380 54.7835 9.3560 55.9435 ;
        RECT 8.5730 54.8200 8.6090 55.9340 ;
        RECT 8.4200 54.8200 8.4470 55.9340 ;
        RECT 7.1780 54.7835 7.1960 55.9435 ;
        RECT 0.1580 54.7835 0.1760 55.9435 ;
        RECT 16.3580 55.8635 16.3760 57.0235 ;
        RECT 9.3380 55.8635 9.3560 57.0235 ;
        RECT 8.5730 55.9000 8.6090 57.0140 ;
        RECT 8.4200 55.9000 8.4470 57.0140 ;
        RECT 7.1780 55.8635 7.1960 57.0235 ;
        RECT 0.1580 55.8635 0.1760 57.0235 ;
        RECT 16.3580 56.9435 16.3760 58.1035 ;
        RECT 9.3380 56.9435 9.3560 58.1035 ;
        RECT 8.5730 56.9800 8.6090 58.0940 ;
        RECT 8.4200 56.9800 8.4470 58.0940 ;
        RECT 7.1780 56.9435 7.1960 58.1035 ;
        RECT 0.1580 56.9435 0.1760 58.1035 ;
        RECT 16.3580 58.0235 16.3760 59.1835 ;
        RECT 9.3380 58.0235 9.3560 59.1835 ;
        RECT 8.5730 58.0600 8.6090 59.1740 ;
        RECT 8.4200 58.0600 8.4470 59.1740 ;
        RECT 7.1780 58.0235 7.1960 59.1835 ;
        RECT 0.1580 58.0235 0.1760 59.1835 ;
        RECT 16.3580 59.1035 16.3760 60.2635 ;
        RECT 9.3380 59.1035 9.3560 60.2635 ;
        RECT 8.5730 59.1400 8.6090 60.2540 ;
        RECT 8.4200 59.1400 8.4470 60.2540 ;
        RECT 7.1780 59.1035 7.1960 60.2635 ;
        RECT 0.1580 59.1035 0.1760 60.2635 ;
      LAYER V3  ;
        RECT 0.1580 1.0760 0.1760 1.1240 ;
        RECT 7.1780 1.0760 7.1960 1.1240 ;
        RECT 8.4200 1.0760 8.4470 1.1240 ;
        RECT 8.5730 1.0760 8.6090 1.1240 ;
        RECT 9.3380 1.0760 9.3560 1.1240 ;
        RECT 16.3580 1.0760 16.3760 1.1240 ;
        RECT 0.1580 2.1560 0.1760 2.2040 ;
        RECT 7.1780 2.1560 7.1960 2.2040 ;
        RECT 8.4200 2.1560 8.4470 2.2040 ;
        RECT 8.5730 2.1560 8.6090 2.2040 ;
        RECT 9.3380 2.1560 9.3560 2.2040 ;
        RECT 16.3580 2.1560 16.3760 2.2040 ;
        RECT 0.1580 3.2360 0.1760 3.2840 ;
        RECT 7.1780 3.2360 7.1960 3.2840 ;
        RECT 8.4200 3.2360 8.4470 3.2840 ;
        RECT 8.5730 3.2360 8.6090 3.2840 ;
        RECT 9.3380 3.2360 9.3560 3.2840 ;
        RECT 16.3580 3.2360 16.3760 3.2840 ;
        RECT 0.1580 4.3160 0.1760 4.3640 ;
        RECT 7.1780 4.3160 7.1960 4.3640 ;
        RECT 8.4200 4.3160 8.4470 4.3640 ;
        RECT 8.5730 4.3160 8.6090 4.3640 ;
        RECT 9.3380 4.3160 9.3560 4.3640 ;
        RECT 16.3580 4.3160 16.3760 4.3640 ;
        RECT 0.1580 5.3960 0.1760 5.4440 ;
        RECT 7.1780 5.3960 7.1960 5.4440 ;
        RECT 8.4200 5.3960 8.4470 5.4440 ;
        RECT 8.5730 5.3960 8.6090 5.4440 ;
        RECT 9.3380 5.3960 9.3560 5.4440 ;
        RECT 16.3580 5.3960 16.3760 5.4440 ;
        RECT 0.1580 6.4760 0.1760 6.5240 ;
        RECT 7.1780 6.4760 7.1960 6.5240 ;
        RECT 8.4200 6.4760 8.4470 6.5240 ;
        RECT 8.5730 6.4760 8.6090 6.5240 ;
        RECT 9.3380 6.4760 9.3560 6.5240 ;
        RECT 16.3580 6.4760 16.3760 6.5240 ;
        RECT 0.1580 7.5560 0.1760 7.6040 ;
        RECT 7.1780 7.5560 7.1960 7.6040 ;
        RECT 8.4200 7.5560 8.4470 7.6040 ;
        RECT 8.5730 7.5560 8.6090 7.6040 ;
        RECT 9.3380 7.5560 9.3560 7.6040 ;
        RECT 16.3580 7.5560 16.3760 7.6040 ;
        RECT 0.1580 8.6360 0.1760 8.6840 ;
        RECT 7.1780 8.6360 7.1960 8.6840 ;
        RECT 8.4200 8.6360 8.4470 8.6840 ;
        RECT 8.5730 8.6360 8.6090 8.6840 ;
        RECT 9.3380 8.6360 9.3560 8.6840 ;
        RECT 16.3580 8.6360 16.3760 8.6840 ;
        RECT 0.1580 9.7160 0.1760 9.7640 ;
        RECT 7.1780 9.7160 7.1960 9.7640 ;
        RECT 8.4200 9.7160 8.4470 9.7640 ;
        RECT 8.5730 9.7160 8.6090 9.7640 ;
        RECT 9.3380 9.7160 9.3560 9.7640 ;
        RECT 16.3580 9.7160 16.3760 9.7640 ;
        RECT 0.1580 10.7960 0.1760 10.8440 ;
        RECT 7.1780 10.7960 7.1960 10.8440 ;
        RECT 8.4200 10.7960 8.4470 10.8440 ;
        RECT 8.5730 10.7960 8.6090 10.8440 ;
        RECT 9.3380 10.7960 9.3560 10.8440 ;
        RECT 16.3580 10.7960 16.3760 10.8440 ;
        RECT 0.1580 11.8760 0.1760 11.9240 ;
        RECT 7.1780 11.8760 7.1960 11.9240 ;
        RECT 8.4200 11.8760 8.4470 11.9240 ;
        RECT 8.5730 11.8760 8.6090 11.9240 ;
        RECT 9.3380 11.8760 9.3560 11.9240 ;
        RECT 16.3580 11.8760 16.3760 11.9240 ;
        RECT 0.1580 12.9560 0.1760 13.0040 ;
        RECT 7.1780 12.9560 7.1960 13.0040 ;
        RECT 8.4200 12.9560 8.4470 13.0040 ;
        RECT 8.5730 12.9560 8.6090 13.0040 ;
        RECT 9.3380 12.9560 9.3560 13.0040 ;
        RECT 16.3580 12.9560 16.3760 13.0040 ;
        RECT 0.1580 14.0360 0.1760 14.0840 ;
        RECT 7.1780 14.0360 7.1960 14.0840 ;
        RECT 8.4200 14.0360 8.4470 14.0840 ;
        RECT 8.5730 14.0360 8.6090 14.0840 ;
        RECT 9.3380 14.0360 9.3560 14.0840 ;
        RECT 16.3580 14.0360 16.3760 14.0840 ;
        RECT 0.1580 15.1160 0.1760 15.1640 ;
        RECT 7.1780 15.1160 7.1960 15.1640 ;
        RECT 8.4200 15.1160 8.4470 15.1640 ;
        RECT 8.5730 15.1160 8.6090 15.1640 ;
        RECT 9.3380 15.1160 9.3560 15.1640 ;
        RECT 16.3580 15.1160 16.3760 15.1640 ;
        RECT 0.1580 16.1960 0.1760 16.2440 ;
        RECT 7.1780 16.1960 7.1960 16.2440 ;
        RECT 8.4200 16.1960 8.4470 16.2440 ;
        RECT 8.5730 16.1960 8.6090 16.2440 ;
        RECT 9.3380 16.1960 9.3560 16.2440 ;
        RECT 16.3580 16.1960 16.3760 16.2440 ;
        RECT 0.1580 17.2760 0.1760 17.3240 ;
        RECT 7.1780 17.2760 7.1960 17.3240 ;
        RECT 8.4200 17.2760 8.4470 17.3240 ;
        RECT 8.5730 17.2760 8.6090 17.3240 ;
        RECT 9.3380 17.2760 9.3560 17.3240 ;
        RECT 16.3580 17.2760 16.3760 17.3240 ;
        RECT 0.1580 18.3560 0.1760 18.4040 ;
        RECT 7.1780 18.3560 7.1960 18.4040 ;
        RECT 8.4200 18.3560 8.4470 18.4040 ;
        RECT 8.5730 18.3560 8.6090 18.4040 ;
        RECT 9.3380 18.3560 9.3560 18.4040 ;
        RECT 16.3580 18.3560 16.3760 18.4040 ;
        RECT 0.1580 19.4360 0.1760 19.4840 ;
        RECT 7.1780 19.4360 7.1960 19.4840 ;
        RECT 8.4200 19.4360 8.4470 19.4840 ;
        RECT 8.5730 19.4360 8.6090 19.4840 ;
        RECT 9.3380 19.4360 9.3560 19.4840 ;
        RECT 16.3580 19.4360 16.3760 19.4840 ;
        RECT 0.1580 20.5160 0.1760 20.5640 ;
        RECT 7.1780 20.5160 7.1960 20.5640 ;
        RECT 8.4200 20.5160 8.4470 20.5640 ;
        RECT 8.5730 20.5160 8.6090 20.5640 ;
        RECT 9.3380 20.5160 9.3560 20.5640 ;
        RECT 16.3580 20.5160 16.3760 20.5640 ;
        RECT 0.1580 21.5960 0.1760 21.6440 ;
        RECT 7.1780 21.5960 7.1960 21.6440 ;
        RECT 8.4200 21.5960 8.4470 21.6440 ;
        RECT 8.5730 21.5960 8.6090 21.6440 ;
        RECT 9.3380 21.5960 9.3560 21.6440 ;
        RECT 16.3580 21.5960 16.3760 21.6440 ;
        RECT 0.1580 22.6760 0.1760 22.7240 ;
        RECT 7.1780 22.6760 7.1960 22.7240 ;
        RECT 8.4200 22.6760 8.4470 22.7240 ;
        RECT 8.5730 22.6760 8.6090 22.7240 ;
        RECT 9.3380 22.6760 9.3560 22.7240 ;
        RECT 16.3580 22.6760 16.3760 22.7240 ;
        RECT 0.1580 23.7560 0.1760 23.8040 ;
        RECT 7.1780 23.7560 7.1960 23.8040 ;
        RECT 8.4200 23.7560 8.4470 23.8040 ;
        RECT 8.5730 23.7560 8.6090 23.8040 ;
        RECT 9.3380 23.7560 9.3560 23.8040 ;
        RECT 16.3580 23.7560 16.3760 23.8040 ;
        RECT 0.1580 24.8360 0.1760 24.8840 ;
        RECT 7.1780 24.8360 7.1960 24.8840 ;
        RECT 8.4200 24.8360 8.4470 24.8840 ;
        RECT 8.5730 24.8360 8.6090 24.8840 ;
        RECT 9.3380 24.8360 9.3560 24.8840 ;
        RECT 16.3580 24.8360 16.3760 24.8840 ;
        RECT 0.1580 25.9160 0.1760 25.9640 ;
        RECT 7.1780 25.9160 7.1960 25.9640 ;
        RECT 8.4200 25.9160 8.4470 25.9640 ;
        RECT 8.5730 25.9160 8.6090 25.9640 ;
        RECT 9.3380 25.9160 9.3560 25.9640 ;
        RECT 16.3580 25.9160 16.3760 25.9640 ;
        RECT 8.3830 33.2610 8.4010 33.4770 ;
        RECT 8.3830 30.0930 8.4010 30.3090 ;
        RECT 8.3830 26.9250 8.4010 27.1410 ;
        RECT 8.4350 33.2610 8.4530 33.4770 ;
        RECT 8.4350 30.0930 8.4530 30.3090 ;
        RECT 8.4350 26.9250 8.4530 27.1410 ;
        RECT 8.4870 33.2610 8.5050 33.4770 ;
        RECT 8.4870 30.0930 8.5050 30.3090 ;
        RECT 8.4870 26.9250 8.5050 27.1410 ;
        RECT 8.5390 33.2610 8.5570 33.4770 ;
        RECT 8.5390 30.0930 8.5570 30.3090 ;
        RECT 8.5390 26.9250 8.5570 27.1410 ;
        RECT 8.5910 33.2610 8.6090 33.4770 ;
        RECT 8.5910 30.0930 8.6090 30.3090 ;
        RECT 8.5910 26.9250 8.6090 27.1410 ;
        RECT 9.3330 26.9255 9.3510 27.1415 ;
        RECT 0.1580 35.1230 0.1760 35.1710 ;
        RECT 7.1780 35.1230 7.1960 35.1710 ;
        RECT 8.4200 35.1230 8.4470 35.1710 ;
        RECT 8.5730 35.1230 8.6090 35.1710 ;
        RECT 9.3380 35.1230 9.3560 35.1710 ;
        RECT 16.3580 35.1230 16.3760 35.1710 ;
        RECT 0.1580 36.2030 0.1760 36.2510 ;
        RECT 7.1780 36.2030 7.1960 36.2510 ;
        RECT 8.4200 36.2030 8.4470 36.2510 ;
        RECT 8.5730 36.2030 8.6090 36.2510 ;
        RECT 9.3380 36.2030 9.3560 36.2510 ;
        RECT 16.3580 36.2030 16.3760 36.2510 ;
        RECT 0.1580 37.2830 0.1760 37.3310 ;
        RECT 7.1780 37.2830 7.1960 37.3310 ;
        RECT 8.4200 37.2830 8.4470 37.3310 ;
        RECT 8.5730 37.2830 8.6090 37.3310 ;
        RECT 9.3380 37.2830 9.3560 37.3310 ;
        RECT 16.3580 37.2830 16.3760 37.3310 ;
        RECT 0.1580 38.3630 0.1760 38.4110 ;
        RECT 7.1780 38.3630 7.1960 38.4110 ;
        RECT 8.4200 38.3630 8.4470 38.4110 ;
        RECT 8.5730 38.3630 8.6090 38.4110 ;
        RECT 9.3380 38.3630 9.3560 38.4110 ;
        RECT 16.3580 38.3630 16.3760 38.4110 ;
        RECT 0.1580 39.4430 0.1760 39.4910 ;
        RECT 7.1780 39.4430 7.1960 39.4910 ;
        RECT 8.4200 39.4430 8.4470 39.4910 ;
        RECT 8.5730 39.4430 8.6090 39.4910 ;
        RECT 9.3380 39.4430 9.3560 39.4910 ;
        RECT 16.3580 39.4430 16.3760 39.4910 ;
        RECT 0.1580 40.5230 0.1760 40.5710 ;
        RECT 7.1780 40.5230 7.1960 40.5710 ;
        RECT 8.4200 40.5230 8.4470 40.5710 ;
        RECT 8.5730 40.5230 8.6090 40.5710 ;
        RECT 9.3380 40.5230 9.3560 40.5710 ;
        RECT 16.3580 40.5230 16.3760 40.5710 ;
        RECT 0.1580 41.6030 0.1760 41.6510 ;
        RECT 7.1780 41.6030 7.1960 41.6510 ;
        RECT 8.4200 41.6030 8.4470 41.6510 ;
        RECT 8.5730 41.6030 8.6090 41.6510 ;
        RECT 9.3380 41.6030 9.3560 41.6510 ;
        RECT 16.3580 41.6030 16.3760 41.6510 ;
        RECT 0.1580 42.6830 0.1760 42.7310 ;
        RECT 7.1780 42.6830 7.1960 42.7310 ;
        RECT 8.4200 42.6830 8.4470 42.7310 ;
        RECT 8.5730 42.6830 8.6090 42.7310 ;
        RECT 9.3380 42.6830 9.3560 42.7310 ;
        RECT 16.3580 42.6830 16.3760 42.7310 ;
        RECT 0.1580 43.7630 0.1760 43.8110 ;
        RECT 7.1780 43.7630 7.1960 43.8110 ;
        RECT 8.4200 43.7630 8.4470 43.8110 ;
        RECT 8.5730 43.7630 8.6090 43.8110 ;
        RECT 9.3380 43.7630 9.3560 43.8110 ;
        RECT 16.3580 43.7630 16.3760 43.8110 ;
        RECT 0.1580 44.8430 0.1760 44.8910 ;
        RECT 7.1780 44.8430 7.1960 44.8910 ;
        RECT 8.4200 44.8430 8.4470 44.8910 ;
        RECT 8.5730 44.8430 8.6090 44.8910 ;
        RECT 9.3380 44.8430 9.3560 44.8910 ;
        RECT 16.3580 44.8430 16.3760 44.8910 ;
        RECT 0.1580 45.9230 0.1760 45.9710 ;
        RECT 7.1780 45.9230 7.1960 45.9710 ;
        RECT 8.4200 45.9230 8.4470 45.9710 ;
        RECT 8.5730 45.9230 8.6090 45.9710 ;
        RECT 9.3380 45.9230 9.3560 45.9710 ;
        RECT 16.3580 45.9230 16.3760 45.9710 ;
        RECT 0.1580 47.0030 0.1760 47.0510 ;
        RECT 7.1780 47.0030 7.1960 47.0510 ;
        RECT 8.4200 47.0030 8.4470 47.0510 ;
        RECT 8.5730 47.0030 8.6090 47.0510 ;
        RECT 9.3380 47.0030 9.3560 47.0510 ;
        RECT 16.3580 47.0030 16.3760 47.0510 ;
        RECT 0.1580 48.0830 0.1760 48.1310 ;
        RECT 7.1780 48.0830 7.1960 48.1310 ;
        RECT 8.4200 48.0830 8.4470 48.1310 ;
        RECT 8.5730 48.0830 8.6090 48.1310 ;
        RECT 9.3380 48.0830 9.3560 48.1310 ;
        RECT 16.3580 48.0830 16.3760 48.1310 ;
        RECT 0.1580 49.1630 0.1760 49.2110 ;
        RECT 7.1780 49.1630 7.1960 49.2110 ;
        RECT 8.4200 49.1630 8.4470 49.2110 ;
        RECT 8.5730 49.1630 8.6090 49.2110 ;
        RECT 9.3380 49.1630 9.3560 49.2110 ;
        RECT 16.3580 49.1630 16.3760 49.2110 ;
        RECT 0.1580 50.2430 0.1760 50.2910 ;
        RECT 7.1780 50.2430 7.1960 50.2910 ;
        RECT 8.4200 50.2430 8.4470 50.2910 ;
        RECT 8.5730 50.2430 8.6090 50.2910 ;
        RECT 9.3380 50.2430 9.3560 50.2910 ;
        RECT 16.3580 50.2430 16.3760 50.2910 ;
        RECT 0.1580 51.3230 0.1760 51.3710 ;
        RECT 7.1780 51.3230 7.1960 51.3710 ;
        RECT 8.4200 51.3230 8.4470 51.3710 ;
        RECT 8.5730 51.3230 8.6090 51.3710 ;
        RECT 9.3380 51.3230 9.3560 51.3710 ;
        RECT 16.3580 51.3230 16.3760 51.3710 ;
        RECT 0.1580 52.4030 0.1760 52.4510 ;
        RECT 7.1780 52.4030 7.1960 52.4510 ;
        RECT 8.4200 52.4030 8.4470 52.4510 ;
        RECT 8.5730 52.4030 8.6090 52.4510 ;
        RECT 9.3380 52.4030 9.3560 52.4510 ;
        RECT 16.3580 52.4030 16.3760 52.4510 ;
        RECT 0.1580 53.4830 0.1760 53.5310 ;
        RECT 7.1780 53.4830 7.1960 53.5310 ;
        RECT 8.4200 53.4830 8.4470 53.5310 ;
        RECT 8.5730 53.4830 8.6090 53.5310 ;
        RECT 9.3380 53.4830 9.3560 53.5310 ;
        RECT 16.3580 53.4830 16.3760 53.5310 ;
        RECT 0.1580 54.5630 0.1760 54.6110 ;
        RECT 7.1780 54.5630 7.1960 54.6110 ;
        RECT 8.4200 54.5630 8.4470 54.6110 ;
        RECT 8.5730 54.5630 8.6090 54.6110 ;
        RECT 9.3380 54.5630 9.3560 54.6110 ;
        RECT 16.3580 54.5630 16.3760 54.6110 ;
        RECT 0.1580 55.6430 0.1760 55.6910 ;
        RECT 7.1780 55.6430 7.1960 55.6910 ;
        RECT 8.4200 55.6430 8.4470 55.6910 ;
        RECT 8.5730 55.6430 8.6090 55.6910 ;
        RECT 9.3380 55.6430 9.3560 55.6910 ;
        RECT 16.3580 55.6430 16.3760 55.6910 ;
        RECT 0.1580 56.7230 0.1760 56.7710 ;
        RECT 7.1780 56.7230 7.1960 56.7710 ;
        RECT 8.4200 56.7230 8.4470 56.7710 ;
        RECT 8.5730 56.7230 8.6090 56.7710 ;
        RECT 9.3380 56.7230 9.3560 56.7710 ;
        RECT 16.3580 56.7230 16.3760 56.7710 ;
        RECT 0.1580 57.8030 0.1760 57.8510 ;
        RECT 7.1780 57.8030 7.1960 57.8510 ;
        RECT 8.4200 57.8030 8.4470 57.8510 ;
        RECT 8.5730 57.8030 8.6090 57.8510 ;
        RECT 9.3380 57.8030 9.3560 57.8510 ;
        RECT 16.3580 57.8030 16.3760 57.8510 ;
        RECT 0.1580 58.8830 0.1760 58.9310 ;
        RECT 7.1780 58.8830 7.1960 58.9310 ;
        RECT 8.4200 58.8830 8.4470 58.9310 ;
        RECT 8.5730 58.8830 8.6090 58.9310 ;
        RECT 9.3380 58.8830 9.3560 58.9310 ;
        RECT 16.3580 58.8830 16.3760 58.9310 ;
        RECT 0.1580 59.9630 0.1760 60.0110 ;
        RECT 7.1780 59.9630 7.1960 60.0110 ;
        RECT 8.4200 59.9630 8.4470 60.0110 ;
        RECT 8.5730 59.9630 8.6090 60.0110 ;
        RECT 9.3380 59.9630 9.3560 60.0110 ;
        RECT 16.3580 59.9630 16.3760 60.0110 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.7910 27.3970 10.8090 27.4340 ;
      LAYER M4  ;
        RECT 10.7390 27.4050 10.8230 27.4290 ;
      LAYER M5  ;
        RECT 10.7880 26.4540 10.8120 29.6940 ;
      LAYER V3  ;
        RECT 10.7910 27.4050 10.8090 27.4290 ;
      LAYER V4  ;
        RECT 10.7880 27.4050 10.8120 27.4290 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.5750 27.4000 10.5930 27.4370 ;
      LAYER M4  ;
        RECT 10.5230 27.4050 10.6070 27.4290 ;
      LAYER M5  ;
        RECT 10.5720 26.4540 10.5960 29.6940 ;
      LAYER V3  ;
        RECT 10.5750 27.4050 10.5930 27.4290 ;
      LAYER V4  ;
        RECT 10.5720 27.4050 10.5960 27.4290 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.3590 26.8210 10.3770 26.8580 ;
      LAYER M4  ;
        RECT 10.3070 26.8290 10.3910 26.8530 ;
      LAYER M5  ;
        RECT 10.3560 26.4540 10.3800 29.6940 ;
      LAYER V3  ;
        RECT 10.3590 26.8290 10.3770 26.8530 ;
      LAYER V4  ;
        RECT 10.3560 26.8290 10.3800 26.8530 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 10.1430 27.0610 10.1610 27.2420 ;
      LAYER M4  ;
        RECT 10.0910 27.2130 10.1750 27.2370 ;
      LAYER M5  ;
        RECT 10.1400 26.4540 10.1640 29.6940 ;
      LAYER V3  ;
        RECT 10.1430 27.2130 10.1610 27.2370 ;
      LAYER V4  ;
        RECT 10.1400 27.2130 10.1640 27.2370 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.9270 26.8240 9.9450 26.8910 ;
      LAYER M4  ;
        RECT 9.8750 26.8290 9.9590 26.8530 ;
      LAYER M5  ;
        RECT 9.9240 26.4540 9.9480 29.6940 ;
      LAYER V3  ;
        RECT 9.9270 26.8290 9.9450 26.8530 ;
      LAYER V4  ;
        RECT 9.9240 26.8290 9.9480 26.8530 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.7110 26.5570 9.7290 26.8100 ;
      LAYER M4  ;
        RECT 9.6590 26.7810 9.7430 26.8050 ;
      LAYER M5  ;
        RECT 9.7080 26.4540 9.7320 29.6940 ;
      LAYER V3  ;
        RECT 9.7110 26.7810 9.7290 26.8050 ;
      LAYER V4  ;
        RECT 9.7080 26.7810 9.7320 26.8050 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.4950 27.5920 9.5130 27.6290 ;
      LAYER M4  ;
        RECT 9.4430 27.5970 9.5270 27.6210 ;
      LAYER M5  ;
        RECT 9.4920 26.4540 9.5160 29.6940 ;
      LAYER V3  ;
        RECT 9.4950 27.5970 9.5130 27.6210 ;
      LAYER V4  ;
        RECT 9.4920 27.5970 9.5160 27.6210 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 9.2790 27.4390 9.2970 27.5300 ;
      LAYER M4  ;
        RECT 9.2270 27.5010 9.3110 27.5250 ;
      LAYER M5  ;
        RECT 9.2760 26.4540 9.3000 29.6940 ;
      LAYER V3  ;
        RECT 9.2790 27.5010 9.2970 27.5250 ;
      LAYER V4  ;
        RECT 9.2760 27.5010 9.3000 27.5250 ;
    END
  END ADDRESS[7]
  PIN ADDRESS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.6310 26.8240 8.6490 26.8910 ;
      LAYER M4  ;
        RECT 8.3470 26.8290 8.6600 26.8530 ;
      LAYER M5  ;
        RECT 8.3580 26.4540 8.3820 29.6940 ;
      LAYER V3  ;
        RECT 8.6310 26.8290 8.6490 26.8530 ;
      LAYER V4  ;
        RECT 8.3580 26.8290 8.3820 26.8530 ;
    END
  END ADDRESS[8]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 8.2350 26.5570 8.2530 26.8100 ;
      LAYER M4  ;
        RECT 8.0230 26.7810 8.2640 26.8050 ;
      LAYER M5  ;
        RECT 8.0340 26.4540 8.0580 29.6940 ;
      LAYER V3  ;
        RECT 8.2350 26.7810 8.2530 26.8050 ;
      LAYER V4  ;
        RECT 8.0340 26.7810 8.0580 26.8050 ;
    END
  END banksel
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.4430 26.8240 7.4610 26.8910 ;
      LAYER M4  ;
        RECT 7.3910 26.8290 7.4750 26.8530 ;
      LAYER M5  ;
        RECT 7.4400 26.4540 7.4640 29.6940 ;
      LAYER V3  ;
        RECT 7.4430 26.8290 7.4610 26.8530 ;
      LAYER V4  ;
        RECT 7.4400 26.8290 7.4640 26.8530 ;
    END
  END write
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2270 27.6880 7.2450 27.7370 ;
      LAYER M4  ;
        RECT 7.1750 27.6930 7.2590 27.7170 ;
      LAYER M5  ;
        RECT 7.2240 26.4540 7.2480 29.6940 ;
      LAYER V3  ;
        RECT 7.2270 27.6930 7.2450 27.7170 ;
      LAYER V4  ;
        RECT 7.2240 27.6930 7.2480 27.7170 ;
    END
  END clk
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 7.2630 26.5570 7.2810 26.8100 ;
      LAYER M4  ;
        RECT 6.9970 26.7810 7.2920 26.8050 ;
      LAYER M5  ;
        RECT 7.0080 26.4540 7.0320 29.6940 ;
      LAYER V3  ;
        RECT 7.2630 26.7810 7.2810 26.8050 ;
      LAYER V4  ;
        RECT 7.0080 26.7810 7.0320 26.8050 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.7950 27.3970 6.8130 27.4340 ;
      LAYER M4  ;
        RECT 6.7430 27.4050 6.8270 27.4290 ;
      LAYER M5  ;
        RECT 6.7920 26.4540 6.8160 29.6940 ;
      LAYER V3  ;
        RECT 6.7950 27.4050 6.8130 27.4290 ;
      LAYER V4  ;
        RECT 6.7920 27.4050 6.8160 27.4290 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.5790 26.8240 6.5970 27.0530 ;
      LAYER M4  ;
        RECT 6.5270 26.8290 6.6110 26.8530 ;
      LAYER M5  ;
        RECT 6.5760 26.4540 6.6000 29.6940 ;
      LAYER V3  ;
        RECT 6.5790 26.8290 6.5970 26.8530 ;
      LAYER V4  ;
        RECT 6.5760 26.8290 6.6000 26.8530 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.3630 26.5570 6.3810 26.8100 ;
      LAYER M4  ;
        RECT 6.3110 26.7810 6.3950 26.8050 ;
      LAYER M5  ;
        RECT 6.3600 26.4540 6.3840 29.6940 ;
      LAYER V3  ;
        RECT 6.3630 26.7810 6.3810 26.8050 ;
      LAYER V4  ;
        RECT 6.3600 26.7810 6.3840 26.8050 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 6.1470 26.8210 6.1650 26.8580 ;
      LAYER M4  ;
        RECT 6.0950 26.8290 6.1790 26.8530 ;
      LAYER M5  ;
        RECT 6.1440 26.4540 6.1680 29.6940 ;
      LAYER V3  ;
        RECT 6.1470 26.8290 6.1650 26.8530 ;
      LAYER V4  ;
        RECT 6.1440 26.8290 6.1680 26.8530 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 5.9310 27.3970 5.9490 27.4340 ;
      LAYER M4  ;
        RECT 5.8790 27.4050 5.9630 27.4290 ;
      LAYER M5  ;
        RECT 5.9280 26.4540 5.9520 29.6940 ;
      LAYER V3  ;
        RECT 5.9310 27.4050 5.9490 27.4290 ;
      LAYER V4  ;
        RECT 5.9280 27.4050 5.9520 27.4290 ;
    END
  END sdel[4]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.4280 8.5970 0.4520 ;
      LAYER M3  ;
        RECT 8.5370 0.3775 8.5550 0.6170 ;
      LAYER V3  ;
        RECT 8.5370 0.4280 8.5550 0.4520 ;
    END
  END dataout[0]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 0.3320 8.6650 0.3560 ;
      LAYER M3  ;
        RECT 8.3120 0.2700 8.3300 0.6750 ;
      LAYER V3  ;
        RECT 8.3120 0.3320 8.3300 0.3560 ;
    END
  END wd[0]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.5080 8.5970 1.5320 ;
      LAYER M3  ;
        RECT 8.5370 1.4575 8.5550 1.6970 ;
      LAYER V3  ;
        RECT 8.5370 1.5080 8.5550 1.5320 ;
    END
  END dataout[1]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 1.4120 8.6650 1.4360 ;
      LAYER M3  ;
        RECT 8.3120 1.3500 8.3300 1.7550 ;
      LAYER V3  ;
        RECT 8.3120 1.4120 8.3300 1.4360 ;
    END
  END wd[1]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.5880 8.5970 2.6120 ;
      LAYER M3  ;
        RECT 8.5370 2.5375 8.5550 2.7770 ;
      LAYER V3  ;
        RECT 8.5370 2.5880 8.5550 2.6120 ;
    END
  END dataout[2]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 2.4920 8.6650 2.5160 ;
      LAYER M3  ;
        RECT 8.3120 2.4300 8.3300 2.8350 ;
      LAYER V3  ;
        RECT 8.3120 2.4920 8.3300 2.5160 ;
    END
  END wd[2]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.6680 8.5970 3.6920 ;
      LAYER M3  ;
        RECT 8.5370 3.6175 8.5550 3.8570 ;
      LAYER V3  ;
        RECT 8.5370 3.6680 8.5550 3.6920 ;
    END
  END dataout[3]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 3.5720 8.6650 3.5960 ;
      LAYER M3  ;
        RECT 8.3120 3.5100 8.3300 3.9150 ;
      LAYER V3  ;
        RECT 8.3120 3.5720 8.3300 3.5960 ;
    END
  END wd[3]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.7480 8.5970 4.7720 ;
      LAYER M3  ;
        RECT 8.5370 4.6975 8.5550 4.9370 ;
      LAYER V3  ;
        RECT 8.5370 4.7480 8.5550 4.7720 ;
    END
  END dataout[4]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 4.6520 8.6650 4.6760 ;
      LAYER M3  ;
        RECT 8.3120 4.5900 8.3300 4.9950 ;
      LAYER V3  ;
        RECT 8.3120 4.6520 8.3300 4.6760 ;
    END
  END wd[4]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.8280 8.5970 5.8520 ;
      LAYER M3  ;
        RECT 8.5370 5.7775 8.5550 6.0170 ;
      LAYER V3  ;
        RECT 8.5370 5.8280 8.5550 5.8520 ;
    END
  END dataout[5]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 5.7320 8.6650 5.7560 ;
      LAYER M3  ;
        RECT 8.3120 5.6700 8.3300 6.0750 ;
      LAYER V3  ;
        RECT 8.3120 5.7320 8.3300 5.7560 ;
    END
  END wd[5]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.9080 8.5970 6.9320 ;
      LAYER M3  ;
        RECT 8.5370 6.8575 8.5550 7.0970 ;
      LAYER V3  ;
        RECT 8.5370 6.9080 8.5550 6.9320 ;
    END
  END dataout[6]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 6.8120 8.6650 6.8360 ;
      LAYER M3  ;
        RECT 8.3120 6.7500 8.3300 7.1550 ;
      LAYER V3  ;
        RECT 8.3120 6.8120 8.3300 6.8360 ;
    END
  END wd[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.9880 8.5970 8.0120 ;
      LAYER M3  ;
        RECT 8.5370 7.9375 8.5550 8.1770 ;
      LAYER V3  ;
        RECT 8.5370 7.9880 8.5550 8.0120 ;
    END
  END dataout[7]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 7.8920 8.6650 7.9160 ;
      LAYER M3  ;
        RECT 8.3120 7.8300 8.3300 8.2350 ;
      LAYER V3  ;
        RECT 8.3120 7.8920 8.3300 7.9160 ;
    END
  END wd[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 9.0680 8.5970 9.0920 ;
      LAYER M3  ;
        RECT 8.5370 9.0175 8.5550 9.2570 ;
      LAYER V3  ;
        RECT 8.5370 9.0680 8.5550 9.0920 ;
    END
  END dataout[8]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 8.9720 8.6650 8.9960 ;
      LAYER M3  ;
        RECT 8.3120 8.9100 8.3300 9.3150 ;
      LAYER V3  ;
        RECT 8.3120 8.9720 8.3300 8.9960 ;
    END
  END wd[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 10.1480 8.5970 10.1720 ;
      LAYER M3  ;
        RECT 8.5370 10.0975 8.5550 10.3370 ;
      LAYER V3  ;
        RECT 8.5370 10.1480 8.5550 10.1720 ;
    END
  END dataout[9]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 10.0520 8.6650 10.0760 ;
      LAYER M3  ;
        RECT 8.3120 9.9900 8.3300 10.3950 ;
      LAYER V3  ;
        RECT 8.3120 10.0520 8.3300 10.0760 ;
    END
  END wd[9]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 11.2280 8.5970 11.2520 ;
      LAYER M3  ;
        RECT 8.5370 11.1775 8.5550 11.4170 ;
      LAYER V3  ;
        RECT 8.5370 11.2280 8.5550 11.2520 ;
    END
  END dataout[10]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 11.1320 8.6650 11.1560 ;
      LAYER M3  ;
        RECT 8.3120 11.0700 8.3300 11.4750 ;
      LAYER V3  ;
        RECT 8.3120 11.1320 8.3300 11.1560 ;
    END
  END wd[10]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 12.3080 8.5970 12.3320 ;
      LAYER M3  ;
        RECT 8.5370 12.2575 8.5550 12.4970 ;
      LAYER V3  ;
        RECT 8.5370 12.3080 8.5550 12.3320 ;
    END
  END dataout[11]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 12.2120 8.6650 12.2360 ;
      LAYER M3  ;
        RECT 8.3120 12.1500 8.3300 12.5550 ;
      LAYER V3  ;
        RECT 8.3120 12.2120 8.3300 12.2360 ;
    END
  END wd[11]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 13.3880 8.5970 13.4120 ;
      LAYER M3  ;
        RECT 8.5370 13.3375 8.5550 13.5770 ;
      LAYER V3  ;
        RECT 8.5370 13.3880 8.5550 13.4120 ;
    END
  END dataout[12]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 13.2920 8.6650 13.3160 ;
      LAYER M3  ;
        RECT 8.3120 13.2300 8.3300 13.6350 ;
      LAYER V3  ;
        RECT 8.3120 13.2920 8.3300 13.3160 ;
    END
  END wd[12]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 14.4680 8.5970 14.4920 ;
      LAYER M3  ;
        RECT 8.5370 14.4175 8.5550 14.6570 ;
      LAYER V3  ;
        RECT 8.5370 14.4680 8.5550 14.4920 ;
    END
  END dataout[13]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 14.3720 8.6650 14.3960 ;
      LAYER M3  ;
        RECT 8.3120 14.3100 8.3300 14.7150 ;
      LAYER V3  ;
        RECT 8.3120 14.3720 8.3300 14.3960 ;
    END
  END wd[13]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 15.5480 8.5970 15.5720 ;
      LAYER M3  ;
        RECT 8.5370 15.4975 8.5550 15.7370 ;
      LAYER V3  ;
        RECT 8.5370 15.5480 8.5550 15.5720 ;
    END
  END dataout[14]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 15.4520 8.6650 15.4760 ;
      LAYER M3  ;
        RECT 8.3120 15.3900 8.3300 15.7950 ;
      LAYER V3  ;
        RECT 8.3120 15.4520 8.3300 15.4760 ;
    END
  END wd[14]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 16.6280 8.5970 16.6520 ;
      LAYER M3  ;
        RECT 8.5370 16.5775 8.5550 16.8170 ;
      LAYER V3  ;
        RECT 8.5370 16.6280 8.5550 16.6520 ;
    END
  END dataout[15]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 16.5320 8.6650 16.5560 ;
      LAYER M3  ;
        RECT 8.3120 16.4700 8.3300 16.8750 ;
      LAYER V3  ;
        RECT 8.3120 16.5320 8.3300 16.5560 ;
    END
  END wd[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 17.7080 8.5970 17.7320 ;
      LAYER M3  ;
        RECT 8.5370 17.6575 8.5550 17.8970 ;
      LAYER V3  ;
        RECT 8.5370 17.7080 8.5550 17.7320 ;
    END
  END dataout[16]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 17.6120 8.6650 17.6360 ;
      LAYER M3  ;
        RECT 8.3120 17.5500 8.3300 17.9550 ;
      LAYER V3  ;
        RECT 8.3120 17.6120 8.3300 17.6360 ;
    END
  END wd[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 18.7880 8.5970 18.8120 ;
      LAYER M3  ;
        RECT 8.5370 18.7375 8.5550 18.9770 ;
      LAYER V3  ;
        RECT 8.5370 18.7880 8.5550 18.8120 ;
    END
  END dataout[17]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 18.6920 8.6650 18.7160 ;
      LAYER M3  ;
        RECT 8.3120 18.6300 8.3300 19.0350 ;
      LAYER V3  ;
        RECT 8.3120 18.6920 8.3300 18.7160 ;
    END
  END wd[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.8680 8.5970 19.8920 ;
      LAYER M3  ;
        RECT 8.5370 19.8175 8.5550 20.0570 ;
      LAYER V3  ;
        RECT 8.5370 19.8680 8.5550 19.8920 ;
    END
  END dataout[18]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 19.7720 8.6650 19.7960 ;
      LAYER M3  ;
        RECT 8.3120 19.7100 8.3300 20.1150 ;
      LAYER V3  ;
        RECT 8.3120 19.7720 8.3300 19.7960 ;
    END
  END wd[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.9480 8.5970 20.9720 ;
      LAYER M3  ;
        RECT 8.5370 20.8975 8.5550 21.1370 ;
      LAYER V3  ;
        RECT 8.5370 20.9480 8.5550 20.9720 ;
    END
  END dataout[19]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 20.8520 8.6650 20.8760 ;
      LAYER M3  ;
        RECT 8.3120 20.7900 8.3300 21.1950 ;
      LAYER V3  ;
        RECT 8.3120 20.8520 8.3300 20.8760 ;
    END
  END wd[19]
  PIN dataout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 22.0280 8.5970 22.0520 ;
      LAYER M3  ;
        RECT 8.5370 21.9775 8.5550 22.2170 ;
      LAYER V3  ;
        RECT 8.5370 22.0280 8.5550 22.0520 ;
    END
  END dataout[20]
  PIN wd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 21.9320 8.6650 21.9560 ;
      LAYER M3  ;
        RECT 8.3120 21.8700 8.3300 22.2750 ;
      LAYER V3  ;
        RECT 8.3120 21.9320 8.3300 21.9560 ;
    END
  END wd[20]
  PIN dataout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.1080 8.5970 23.1320 ;
      LAYER M3  ;
        RECT 8.5370 23.0575 8.5550 23.2970 ;
      LAYER V3  ;
        RECT 8.5370 23.1080 8.5550 23.1320 ;
    END
  END dataout[21]
  PIN wd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 23.0120 8.6650 23.0360 ;
      LAYER M3  ;
        RECT 8.3120 22.9500 8.3300 23.3550 ;
      LAYER V3  ;
        RECT 8.3120 23.0120 8.3300 23.0360 ;
    END
  END wd[21]
  PIN dataout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.1880 8.5970 24.2120 ;
      LAYER M3  ;
        RECT 8.5370 24.1375 8.5550 24.3770 ;
      LAYER V3  ;
        RECT 8.5370 24.1880 8.5550 24.2120 ;
    END
  END dataout[22]
  PIN wd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 24.0920 8.6650 24.1160 ;
      LAYER M3  ;
        RECT 8.3120 24.0300 8.3300 24.4350 ;
      LAYER V3  ;
        RECT 8.3120 24.0920 8.3300 24.1160 ;
    END
  END wd[22]
  PIN dataout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.2680 8.5970 25.2920 ;
      LAYER M3  ;
        RECT 8.5370 25.2175 8.5550 25.4570 ;
      LAYER V3  ;
        RECT 8.5370 25.2680 8.5550 25.2920 ;
    END
  END dataout[23]
  PIN wd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 25.1720 8.6650 25.1960 ;
      LAYER M3  ;
        RECT 8.3120 25.1100 8.3300 25.5150 ;
      LAYER V3  ;
        RECT 8.3120 25.1720 8.3300 25.1960 ;
    END
  END wd[23]
  PIN dataout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 34.4750 8.5970 34.4990 ;
      LAYER M3  ;
        RECT 8.5370 34.4245 8.5550 34.6640 ;
      LAYER V3  ;
        RECT 8.5370 34.4750 8.5550 34.4990 ;
    END
  END dataout[24]
  PIN wd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 34.3790 8.6650 34.4030 ;
      LAYER M3  ;
        RECT 8.3120 34.3170 8.3300 34.7220 ;
      LAYER V3  ;
        RECT 8.3120 34.3790 8.3300 34.4030 ;
    END
  END wd[24]
  PIN dataout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 35.5550 8.5970 35.5790 ;
      LAYER M3  ;
        RECT 8.5370 35.5045 8.5550 35.7440 ;
      LAYER V3  ;
        RECT 8.5370 35.5550 8.5550 35.5790 ;
    END
  END dataout[25]
  PIN wd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 35.4590 8.6650 35.4830 ;
      LAYER M3  ;
        RECT 8.3120 35.3970 8.3300 35.8020 ;
      LAYER V3  ;
        RECT 8.3120 35.4590 8.3300 35.4830 ;
    END
  END wd[25]
  PIN dataout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 36.6350 8.5970 36.6590 ;
      LAYER M3  ;
        RECT 8.5370 36.5845 8.5550 36.8240 ;
      LAYER V3  ;
        RECT 8.5370 36.6350 8.5550 36.6590 ;
    END
  END dataout[26]
  PIN wd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 36.5390 8.6650 36.5630 ;
      LAYER M3  ;
        RECT 8.3120 36.4770 8.3300 36.8820 ;
      LAYER V3  ;
        RECT 8.3120 36.5390 8.3300 36.5630 ;
    END
  END wd[26]
  PIN dataout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 37.7150 8.5970 37.7390 ;
      LAYER M3  ;
        RECT 8.5370 37.6645 8.5550 37.9040 ;
      LAYER V3  ;
        RECT 8.5370 37.7150 8.5550 37.7390 ;
    END
  END dataout[27]
  PIN wd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 37.6190 8.6650 37.6430 ;
      LAYER M3  ;
        RECT 8.3120 37.5570 8.3300 37.9620 ;
      LAYER V3  ;
        RECT 8.3120 37.6190 8.3300 37.6430 ;
    END
  END wd[27]
  PIN dataout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 38.7950 8.5970 38.8190 ;
      LAYER M3  ;
        RECT 8.5370 38.7445 8.5550 38.9840 ;
      LAYER V3  ;
        RECT 8.5370 38.7950 8.5550 38.8190 ;
    END
  END dataout[28]
  PIN wd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 38.6990 8.6650 38.7230 ;
      LAYER M3  ;
        RECT 8.3120 38.6370 8.3300 39.0420 ;
      LAYER V3  ;
        RECT 8.3120 38.6990 8.3300 38.7230 ;
    END
  END wd[28]
  PIN dataout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 39.8750 8.5970 39.8990 ;
      LAYER M3  ;
        RECT 8.5370 39.8245 8.5550 40.0640 ;
      LAYER V3  ;
        RECT 8.5370 39.8750 8.5550 39.8990 ;
    END
  END dataout[29]
  PIN wd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 39.7790 8.6650 39.8030 ;
      LAYER M3  ;
        RECT 8.3120 39.7170 8.3300 40.1220 ;
      LAYER V3  ;
        RECT 8.3120 39.7790 8.3300 39.8030 ;
    END
  END wd[29]
  PIN dataout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 40.9550 8.5970 40.9790 ;
      LAYER M3  ;
        RECT 8.5370 40.9045 8.5550 41.1440 ;
      LAYER V3  ;
        RECT 8.5370 40.9550 8.5550 40.9790 ;
    END
  END dataout[30]
  PIN wd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 40.8590 8.6650 40.8830 ;
      LAYER M3  ;
        RECT 8.3120 40.7970 8.3300 41.2020 ;
      LAYER V3  ;
        RECT 8.3120 40.8590 8.3300 40.8830 ;
    END
  END wd[30]
  PIN dataout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 42.0350 8.5970 42.0590 ;
      LAYER M3  ;
        RECT 8.5370 41.9845 8.5550 42.2240 ;
      LAYER V3  ;
        RECT 8.5370 42.0350 8.5550 42.0590 ;
    END
  END dataout[31]
  PIN wd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 41.9390 8.6650 41.9630 ;
      LAYER M3  ;
        RECT 8.3120 41.8770 8.3300 42.2820 ;
      LAYER V3  ;
        RECT 8.3120 41.9390 8.3300 41.9630 ;
    END
  END wd[31]
  PIN dataout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 43.1150 8.5970 43.1390 ;
      LAYER M3  ;
        RECT 8.5370 43.0645 8.5550 43.3040 ;
      LAYER V3  ;
        RECT 8.5370 43.1150 8.5550 43.1390 ;
    END
  END dataout[32]
  PIN wd[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 43.0190 8.6650 43.0430 ;
      LAYER M3  ;
        RECT 8.3120 42.9570 8.3300 43.3620 ;
      LAYER V3  ;
        RECT 8.3120 43.0190 8.3300 43.0430 ;
    END
  END wd[32]
  PIN dataout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 44.1950 8.5970 44.2190 ;
      LAYER M3  ;
        RECT 8.5370 44.1445 8.5550 44.3840 ;
      LAYER V3  ;
        RECT 8.5370 44.1950 8.5550 44.2190 ;
    END
  END dataout[33]
  PIN wd[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 44.0990 8.6650 44.1230 ;
      LAYER M3  ;
        RECT 8.3120 44.0370 8.3300 44.4420 ;
      LAYER V3  ;
        RECT 8.3120 44.0990 8.3300 44.1230 ;
    END
  END wd[33]
  PIN dataout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 45.2750 8.5970 45.2990 ;
      LAYER M3  ;
        RECT 8.5370 45.2245 8.5550 45.4640 ;
      LAYER V3  ;
        RECT 8.5370 45.2750 8.5550 45.2990 ;
    END
  END dataout[34]
  PIN wd[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 45.1790 8.6650 45.2030 ;
      LAYER M3  ;
        RECT 8.3120 45.1170 8.3300 45.5220 ;
      LAYER V3  ;
        RECT 8.3120 45.1790 8.3300 45.2030 ;
    END
  END wd[34]
  PIN dataout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 46.3550 8.5970 46.3790 ;
      LAYER M3  ;
        RECT 8.5370 46.3045 8.5550 46.5440 ;
      LAYER V3  ;
        RECT 8.5370 46.3550 8.5550 46.3790 ;
    END
  END dataout[35]
  PIN wd[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 46.2590 8.6650 46.2830 ;
      LAYER M3  ;
        RECT 8.3120 46.1970 8.3300 46.6020 ;
      LAYER V3  ;
        RECT 8.3120 46.2590 8.3300 46.2830 ;
    END
  END wd[35]
  PIN dataout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 47.4350 8.5970 47.4590 ;
      LAYER M3  ;
        RECT 8.5370 47.3845 8.5550 47.6240 ;
      LAYER V3  ;
        RECT 8.5370 47.4350 8.5550 47.4590 ;
    END
  END dataout[36]
  PIN wd[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 47.3390 8.6650 47.3630 ;
      LAYER M3  ;
        RECT 8.3120 47.2770 8.3300 47.6820 ;
      LAYER V3  ;
        RECT 8.3120 47.3390 8.3300 47.3630 ;
    END
  END wd[36]
  PIN dataout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 48.5150 8.5970 48.5390 ;
      LAYER M3  ;
        RECT 8.5370 48.4645 8.5550 48.7040 ;
      LAYER V3  ;
        RECT 8.5370 48.5150 8.5550 48.5390 ;
    END
  END dataout[37]
  PIN wd[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 48.4190 8.6650 48.4430 ;
      LAYER M3  ;
        RECT 8.3120 48.3570 8.3300 48.7620 ;
      LAYER V3  ;
        RECT 8.3120 48.4190 8.3300 48.4430 ;
    END
  END wd[37]
  PIN dataout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 49.5950 8.5970 49.6190 ;
      LAYER M3  ;
        RECT 8.5370 49.5445 8.5550 49.7840 ;
      LAYER V3  ;
        RECT 8.5370 49.5950 8.5550 49.6190 ;
    END
  END dataout[38]
  PIN wd[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 49.4990 8.6650 49.5230 ;
      LAYER M3  ;
        RECT 8.3120 49.4370 8.3300 49.8420 ;
      LAYER V3  ;
        RECT 8.3120 49.4990 8.3300 49.5230 ;
    END
  END wd[38]
  PIN dataout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 50.6750 8.5970 50.6990 ;
      LAYER M3  ;
        RECT 8.5370 50.6245 8.5550 50.8640 ;
      LAYER V3  ;
        RECT 8.5370 50.6750 8.5550 50.6990 ;
    END
  END dataout[39]
  PIN wd[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 50.5790 8.6650 50.6030 ;
      LAYER M3  ;
        RECT 8.3120 50.5170 8.3300 50.9220 ;
      LAYER V3  ;
        RECT 8.3120 50.5790 8.3300 50.6030 ;
    END
  END wd[39]
  PIN dataout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 51.7550 8.5970 51.7790 ;
      LAYER M3  ;
        RECT 8.5370 51.7045 8.5550 51.9440 ;
      LAYER V3  ;
        RECT 8.5370 51.7550 8.5550 51.7790 ;
    END
  END dataout[40]
  PIN wd[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 51.6590 8.6650 51.6830 ;
      LAYER M3  ;
        RECT 8.3120 51.5970 8.3300 52.0020 ;
      LAYER V3  ;
        RECT 8.3120 51.6590 8.3300 51.6830 ;
    END
  END wd[40]
  PIN dataout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 52.8350 8.5970 52.8590 ;
      LAYER M3  ;
        RECT 8.5370 52.7845 8.5550 53.0240 ;
      LAYER V3  ;
        RECT 8.5370 52.8350 8.5550 52.8590 ;
    END
  END dataout[41]
  PIN wd[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 52.7390 8.6650 52.7630 ;
      LAYER M3  ;
        RECT 8.3120 52.6770 8.3300 53.0820 ;
      LAYER V3  ;
        RECT 8.3120 52.7390 8.3300 52.7630 ;
    END
  END wd[41]
  PIN dataout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 53.9150 8.5970 53.9390 ;
      LAYER M3  ;
        RECT 8.5370 53.8645 8.5550 54.1040 ;
      LAYER V3  ;
        RECT 8.5370 53.9150 8.5550 53.9390 ;
    END
  END dataout[42]
  PIN wd[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 53.8190 8.6650 53.8430 ;
      LAYER M3  ;
        RECT 8.3120 53.7570 8.3300 54.1620 ;
      LAYER V3  ;
        RECT 8.3120 53.8190 8.3300 53.8430 ;
    END
  END wd[42]
  PIN dataout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 54.9950 8.5970 55.0190 ;
      LAYER M3  ;
        RECT 8.5370 54.9445 8.5550 55.1840 ;
      LAYER V3  ;
        RECT 8.5370 54.9950 8.5550 55.0190 ;
    END
  END dataout[43]
  PIN wd[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 54.8990 8.6650 54.9230 ;
      LAYER M3  ;
        RECT 8.3120 54.8370 8.3300 55.2420 ;
      LAYER V3  ;
        RECT 8.3120 54.8990 8.3300 54.9230 ;
    END
  END wd[43]
  PIN dataout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 56.0750 8.5970 56.0990 ;
      LAYER M3  ;
        RECT 8.5370 56.0245 8.5550 56.2640 ;
      LAYER V3  ;
        RECT 8.5370 56.0750 8.5550 56.0990 ;
    END
  END dataout[44]
  PIN wd[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 55.9790 8.6650 56.0030 ;
      LAYER M3  ;
        RECT 8.3120 55.9170 8.3300 56.3220 ;
      LAYER V3  ;
        RECT 8.3120 55.9790 8.3300 56.0030 ;
    END
  END wd[44]
  PIN dataout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 57.1550 8.5970 57.1790 ;
      LAYER M3  ;
        RECT 8.5370 57.1045 8.5550 57.3440 ;
      LAYER V3  ;
        RECT 8.5370 57.1550 8.5550 57.1790 ;
    END
  END dataout[45]
  PIN wd[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 57.0590 8.6650 57.0830 ;
      LAYER M3  ;
        RECT 8.3120 56.9970 8.3300 57.4020 ;
      LAYER V3  ;
        RECT 8.3120 57.0590 8.3300 57.0830 ;
    END
  END wd[45]
  PIN dataout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 58.2350 8.5970 58.2590 ;
      LAYER M3  ;
        RECT 8.5370 58.1845 8.5550 58.4240 ;
      LAYER V3  ;
        RECT 8.5370 58.2350 8.5550 58.2590 ;
    END
  END dataout[46]
  PIN wd[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 58.1390 8.6650 58.1630 ;
      LAYER M3  ;
        RECT 8.3120 58.0770 8.3300 58.4820 ;
      LAYER V3  ;
        RECT 8.3120 58.1390 8.3300 58.1630 ;
    END
  END wd[46]
  PIN dataout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 59.3150 8.5970 59.3390 ;
      LAYER M3  ;
        RECT 8.5370 59.2645 8.5550 59.5040 ;
      LAYER V3  ;
        RECT 8.5370 59.3150 8.5550 59.3390 ;
    END
  END dataout[47]
  PIN wd[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4  ;
        RECT 7.9490 59.2190 8.6650 59.2430 ;
      LAYER M3  ;
        RECT 8.3120 59.1570 8.3300 59.5620 ;
      LAYER V3  ;
        RECT 8.3120 59.2190 8.3300 59.2430 ;
    END
  END wd[47]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0000 26.1570 16.5240 34.8105 ;
        RECT 0.0050 34.3035 16.5290 35.3970 ;
        RECT 0.0050 35.3835 16.5290 36.4770 ;
        RECT 0.0050 36.4635 16.5290 37.5570 ;
        RECT 0.0050 37.5435 16.5290 38.6370 ;
        RECT 0.0050 38.6235 16.5290 39.7170 ;
        RECT 0.0050 39.7035 16.5290 40.7970 ;
        RECT 0.0050 40.7835 16.5290 41.8770 ;
        RECT 0.0050 41.8635 16.5290 42.9570 ;
        RECT 0.0050 42.9435 16.5290 44.0370 ;
        RECT 0.0050 44.0235 16.5290 45.1170 ;
        RECT 0.0050 45.1035 16.5290 46.1970 ;
        RECT 0.0050 46.1835 16.5290 47.2770 ;
        RECT 0.0050 47.2635 16.5290 48.3570 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0000 26.1570 16.5240 34.8105 ;
        RECT 0.0050 34.3035 16.5290 35.3970 ;
        RECT 0.0050 35.3835 16.5290 36.4770 ;
        RECT 0.0050 36.4635 16.5290 37.5570 ;
        RECT 0.0050 37.5435 16.5290 38.6370 ;
        RECT 0.0050 38.6235 16.5290 39.7170 ;
        RECT 0.0050 39.7035 16.5290 40.7970 ;
        RECT 0.0050 40.7835 16.5290 41.8770 ;
        RECT 0.0050 41.8635 16.5290 42.9570 ;
        RECT 0.0050 42.9435 16.5290 44.0370 ;
        RECT 0.0050 44.0235 16.5290 45.1170 ;
        RECT 0.0050 45.1035 16.5290 46.1970 ;
        RECT 0.0050 46.1835 16.5290 47.2770 ;
        RECT 0.0050 47.2635 16.5290 48.3570 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
  LAYER V1 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0000 26.1570 16.5240 34.8105 ;
        RECT 0.0050 34.3035 16.5290 35.3970 ;
        RECT 0.0050 35.3835 16.5290 36.4770 ;
        RECT 0.0050 36.4635 16.5290 37.5570 ;
        RECT 0.0050 37.5435 16.5290 38.6370 ;
        RECT 0.0050 38.6235 16.5290 39.7170 ;
        RECT 0.0050 39.7035 16.5290 40.7970 ;
        RECT 0.0050 40.7835 16.5290 41.8770 ;
        RECT 0.0050 41.8635 16.5290 42.9570 ;
        RECT 0.0050 42.9435 16.5290 44.0370 ;
        RECT 0.0050 44.0235 16.5290 45.1170 ;
        RECT 0.0050 45.1035 16.5290 46.1970 ;
        RECT 0.0050 46.1835 16.5290 47.2770 ;
        RECT 0.0050 47.2635 16.5290 48.3570 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
  LAYER V2 SPACING 0.018  ;
      RECT 0.0050 0.2565 16.5290 1.3500 ;
      RECT 0.0050 1.3365 16.5290 2.4300 ;
      RECT 0.0050 2.4165 16.5290 3.5100 ;
      RECT 0.0050 3.4965 16.5290 4.5900 ;
      RECT 0.0050 4.5765 16.5290 5.6700 ;
      RECT 0.0050 5.6565 16.5290 6.7500 ;
      RECT 0.0050 6.7365 16.5290 7.8300 ;
      RECT 0.0050 7.8165 16.5290 8.9100 ;
      RECT 0.0050 8.8965 16.5290 9.9900 ;
      RECT 0.0050 9.9765 16.5290 11.0700 ;
      RECT 0.0050 11.0565 16.5290 12.1500 ;
      RECT 0.0050 12.1365 16.5290 13.2300 ;
      RECT 0.0050 13.2165 16.5290 14.3100 ;
      RECT 0.0050 14.2965 16.5290 15.3900 ;
      RECT 0.0050 15.3765 16.5290 16.4700 ;
      RECT 0.0050 16.4565 16.5290 17.5500 ;
      RECT 0.0050 17.5365 16.5290 18.6300 ;
      RECT 0.0050 18.6165 16.5290 19.7100 ;
      RECT 0.0050 19.6965 16.5290 20.7900 ;
      RECT 0.0050 20.7765 16.5290 21.8700 ;
      RECT 0.0050 21.8565 16.5290 22.9500 ;
      RECT 0.0050 22.9365 16.5290 24.0300 ;
      RECT 0.0050 24.0165 16.5290 25.1100 ;
      RECT 0.0050 25.0965 16.5290 26.1900 ;
      RECT 0.0000 26.1570 16.5240 34.8105 ;
        RECT 0.0050 34.3035 16.5290 35.3970 ;
        RECT 0.0050 35.3835 16.5290 36.4770 ;
        RECT 0.0050 36.4635 16.5290 37.5570 ;
        RECT 0.0050 37.5435 16.5290 38.6370 ;
        RECT 0.0050 38.6235 16.5290 39.7170 ;
        RECT 0.0050 39.7035 16.5290 40.7970 ;
        RECT 0.0050 40.7835 16.5290 41.8770 ;
        RECT 0.0050 41.8635 16.5290 42.9570 ;
        RECT 0.0050 42.9435 16.5290 44.0370 ;
        RECT 0.0050 44.0235 16.5290 45.1170 ;
        RECT 0.0050 45.1035 16.5290 46.1970 ;
        RECT 0.0050 46.1835 16.5290 47.2770 ;
        RECT 0.0050 47.2635 16.5290 48.3570 ;
        RECT 0.0050 48.3435 16.5290 49.4370 ;
        RECT 0.0050 49.4235 16.5290 50.5170 ;
        RECT 0.0050 50.5035 16.5290 51.5970 ;
        RECT 0.0050 51.5835 16.5290 52.6770 ;
        RECT 0.0050 52.6635 16.5290 53.7570 ;
        RECT 0.0050 53.7435 16.5290 54.8370 ;
        RECT 0.0050 54.8235 16.5290 55.9170 ;
        RECT 0.0050 55.9035 16.5290 56.9970 ;
        RECT 0.0050 56.9835 16.5290 58.0770 ;
        RECT 0.0050 58.0635 16.5290 59.1570 ;
        RECT 0.0050 59.1435 16.5290 60.2370 ;
  LAYER M3  ;
      RECT 8.6990 0.3450 8.7170 1.2805 ;
      RECT 8.6630 0.3450 8.6810 1.2805 ;
      RECT 8.6270 0.9220 8.6450 1.2445 ;
      RECT 8.5100 1.1190 8.5280 1.2285 ;
      RECT 8.5010 0.3775 8.5190 0.6170 ;
      RECT 8.4650 0.9585 8.4830 1.1120 ;
      RECT 8.3840 0.9840 8.4020 1.2420 ;
      RECT 7.8440 0.3450 7.8620 1.2805 ;
      RECT 7.8080 0.3450 7.8260 1.2805 ;
      RECT 7.7720 0.5260 7.7900 1.0940 ;
      RECT 8.6990 1.4250 8.7170 2.3605 ;
      RECT 8.6630 1.4250 8.6810 2.3605 ;
      RECT 8.6270 2.0020 8.6450 2.3245 ;
      RECT 8.5100 2.1990 8.5280 2.3085 ;
      RECT 8.5010 1.4575 8.5190 1.6970 ;
      RECT 8.4650 2.0385 8.4830 2.1920 ;
      RECT 8.3840 2.0640 8.4020 2.3220 ;
      RECT 7.8440 1.4250 7.8620 2.3605 ;
      RECT 7.8080 1.4250 7.8260 2.3605 ;
      RECT 7.7720 1.6060 7.7900 2.1740 ;
      RECT 8.6990 2.5050 8.7170 3.4405 ;
      RECT 8.6630 2.5050 8.6810 3.4405 ;
      RECT 8.6270 3.0820 8.6450 3.4045 ;
      RECT 8.5100 3.2790 8.5280 3.3885 ;
      RECT 8.5010 2.5375 8.5190 2.7770 ;
      RECT 8.4650 3.1185 8.4830 3.2720 ;
      RECT 8.3840 3.1440 8.4020 3.4020 ;
      RECT 7.8440 2.5050 7.8620 3.4405 ;
      RECT 7.8080 2.5050 7.8260 3.4405 ;
      RECT 7.7720 2.6860 7.7900 3.2540 ;
      RECT 8.6990 3.5850 8.7170 4.5205 ;
      RECT 8.6630 3.5850 8.6810 4.5205 ;
      RECT 8.6270 4.1620 8.6450 4.4845 ;
      RECT 8.5100 4.3590 8.5280 4.4685 ;
      RECT 8.5010 3.6175 8.5190 3.8570 ;
      RECT 8.4650 4.1985 8.4830 4.3520 ;
      RECT 8.3840 4.2240 8.4020 4.4820 ;
      RECT 7.8440 3.5850 7.8620 4.5205 ;
      RECT 7.8080 3.5850 7.8260 4.5205 ;
      RECT 7.7720 3.7660 7.7900 4.3340 ;
      RECT 8.6990 4.6650 8.7170 5.6005 ;
      RECT 8.6630 4.6650 8.6810 5.6005 ;
      RECT 8.6270 5.2420 8.6450 5.5645 ;
      RECT 8.5100 5.4390 8.5280 5.5485 ;
      RECT 8.5010 4.6975 8.5190 4.9370 ;
      RECT 8.4650 5.2785 8.4830 5.4320 ;
      RECT 8.3840 5.3040 8.4020 5.5620 ;
      RECT 7.8440 4.6650 7.8620 5.6005 ;
      RECT 7.8080 4.6650 7.8260 5.6005 ;
      RECT 7.7720 4.8460 7.7900 5.4140 ;
      RECT 8.6990 5.7450 8.7170 6.6805 ;
      RECT 8.6630 5.7450 8.6810 6.6805 ;
      RECT 8.6270 6.3220 8.6450 6.6445 ;
      RECT 8.5100 6.5190 8.5280 6.6285 ;
      RECT 8.5010 5.7775 8.5190 6.0170 ;
      RECT 8.4650 6.3585 8.4830 6.5120 ;
      RECT 8.3840 6.3840 8.4020 6.6420 ;
      RECT 7.8440 5.7450 7.8620 6.6805 ;
      RECT 7.8080 5.7450 7.8260 6.6805 ;
      RECT 7.7720 5.9260 7.7900 6.4940 ;
      RECT 8.6990 6.8250 8.7170 7.7605 ;
      RECT 8.6630 6.8250 8.6810 7.7605 ;
      RECT 8.6270 7.4020 8.6450 7.7245 ;
      RECT 8.5100 7.5990 8.5280 7.7085 ;
      RECT 8.5010 6.8575 8.5190 7.0970 ;
      RECT 8.4650 7.4385 8.4830 7.5920 ;
      RECT 8.3840 7.4640 8.4020 7.7220 ;
      RECT 7.8440 6.8250 7.8620 7.7605 ;
      RECT 7.8080 6.8250 7.8260 7.7605 ;
      RECT 7.7720 7.0060 7.7900 7.5740 ;
      RECT 8.6990 7.9050 8.7170 8.8405 ;
      RECT 8.6630 7.9050 8.6810 8.8405 ;
      RECT 8.6270 8.4820 8.6450 8.8045 ;
      RECT 8.5100 8.6790 8.5280 8.7885 ;
      RECT 8.5010 7.9375 8.5190 8.1770 ;
      RECT 8.4650 8.5185 8.4830 8.6720 ;
      RECT 8.3840 8.5440 8.4020 8.8020 ;
      RECT 7.8440 7.9050 7.8620 8.8405 ;
      RECT 7.8080 7.9050 7.8260 8.8405 ;
      RECT 7.7720 8.0860 7.7900 8.6540 ;
      RECT 8.6990 8.9850 8.7170 9.9205 ;
      RECT 8.6630 8.9850 8.6810 9.9205 ;
      RECT 8.6270 9.5620 8.6450 9.8845 ;
      RECT 8.5100 9.7590 8.5280 9.8685 ;
      RECT 8.5010 9.0175 8.5190 9.2570 ;
      RECT 8.4650 9.5985 8.4830 9.7520 ;
      RECT 8.3840 9.6240 8.4020 9.8820 ;
      RECT 7.8440 8.9850 7.8620 9.9205 ;
      RECT 7.8080 8.9850 7.8260 9.9205 ;
      RECT 7.7720 9.1660 7.7900 9.7340 ;
      RECT 8.6990 10.0650 8.7170 11.0005 ;
      RECT 8.6630 10.0650 8.6810 11.0005 ;
      RECT 8.6270 10.6420 8.6450 10.9645 ;
      RECT 8.5100 10.8390 8.5280 10.9485 ;
      RECT 8.5010 10.0975 8.5190 10.3370 ;
      RECT 8.4650 10.6785 8.4830 10.8320 ;
      RECT 8.3840 10.7040 8.4020 10.9620 ;
      RECT 7.8440 10.0650 7.8620 11.0005 ;
      RECT 7.8080 10.0650 7.8260 11.0005 ;
      RECT 7.7720 10.2460 7.7900 10.8140 ;
      RECT 8.6990 11.1450 8.7170 12.0805 ;
      RECT 8.6630 11.1450 8.6810 12.0805 ;
      RECT 8.6270 11.7220 8.6450 12.0445 ;
      RECT 8.5100 11.9190 8.5280 12.0285 ;
      RECT 8.5010 11.1775 8.5190 11.4170 ;
      RECT 8.4650 11.7585 8.4830 11.9120 ;
      RECT 8.3840 11.7840 8.4020 12.0420 ;
      RECT 7.8440 11.1450 7.8620 12.0805 ;
      RECT 7.8080 11.1450 7.8260 12.0805 ;
      RECT 7.7720 11.3260 7.7900 11.8940 ;
      RECT 8.6990 12.2250 8.7170 13.1605 ;
      RECT 8.6630 12.2250 8.6810 13.1605 ;
      RECT 8.6270 12.8020 8.6450 13.1245 ;
      RECT 8.5100 12.9990 8.5280 13.1085 ;
      RECT 8.5010 12.2575 8.5190 12.4970 ;
      RECT 8.4650 12.8385 8.4830 12.9920 ;
      RECT 8.3840 12.8640 8.4020 13.1220 ;
      RECT 7.8440 12.2250 7.8620 13.1605 ;
      RECT 7.8080 12.2250 7.8260 13.1605 ;
      RECT 7.7720 12.4060 7.7900 12.9740 ;
      RECT 8.6990 13.3050 8.7170 14.2405 ;
      RECT 8.6630 13.3050 8.6810 14.2405 ;
      RECT 8.6270 13.8820 8.6450 14.2045 ;
      RECT 8.5100 14.0790 8.5280 14.1885 ;
      RECT 8.5010 13.3375 8.5190 13.5770 ;
      RECT 8.4650 13.9185 8.4830 14.0720 ;
      RECT 8.3840 13.9440 8.4020 14.2020 ;
      RECT 7.8440 13.3050 7.8620 14.2405 ;
      RECT 7.8080 13.3050 7.8260 14.2405 ;
      RECT 7.7720 13.4860 7.7900 14.0540 ;
      RECT 8.6990 14.3850 8.7170 15.3205 ;
      RECT 8.6630 14.3850 8.6810 15.3205 ;
      RECT 8.6270 14.9620 8.6450 15.2845 ;
      RECT 8.5100 15.1590 8.5280 15.2685 ;
      RECT 8.5010 14.4175 8.5190 14.6570 ;
      RECT 8.4650 14.9985 8.4830 15.1520 ;
      RECT 8.3840 15.0240 8.4020 15.2820 ;
      RECT 7.8440 14.3850 7.8620 15.3205 ;
      RECT 7.8080 14.3850 7.8260 15.3205 ;
      RECT 7.7720 14.5660 7.7900 15.1340 ;
      RECT 8.6990 15.4650 8.7170 16.4005 ;
      RECT 8.6630 15.4650 8.6810 16.4005 ;
      RECT 8.6270 16.0420 8.6450 16.3645 ;
      RECT 8.5100 16.2390 8.5280 16.3485 ;
      RECT 8.5010 15.4975 8.5190 15.7370 ;
      RECT 8.4650 16.0785 8.4830 16.2320 ;
      RECT 8.3840 16.1040 8.4020 16.3620 ;
      RECT 7.8440 15.4650 7.8620 16.4005 ;
      RECT 7.8080 15.4650 7.8260 16.4005 ;
      RECT 7.7720 15.6460 7.7900 16.2140 ;
      RECT 8.6990 16.5450 8.7170 17.4805 ;
      RECT 8.6630 16.5450 8.6810 17.4805 ;
      RECT 8.6270 17.1220 8.6450 17.4445 ;
      RECT 8.5100 17.3190 8.5280 17.4285 ;
      RECT 8.5010 16.5775 8.5190 16.8170 ;
      RECT 8.4650 17.1585 8.4830 17.3120 ;
      RECT 8.3840 17.1840 8.4020 17.4420 ;
      RECT 7.8440 16.5450 7.8620 17.4805 ;
      RECT 7.8080 16.5450 7.8260 17.4805 ;
      RECT 7.7720 16.7260 7.7900 17.2940 ;
      RECT 8.6990 17.6250 8.7170 18.5605 ;
      RECT 8.6630 17.6250 8.6810 18.5605 ;
      RECT 8.6270 18.2020 8.6450 18.5245 ;
      RECT 8.5100 18.3990 8.5280 18.5085 ;
      RECT 8.5010 17.6575 8.5190 17.8970 ;
      RECT 8.4650 18.2385 8.4830 18.3920 ;
      RECT 8.3840 18.2640 8.4020 18.5220 ;
      RECT 7.8440 17.6250 7.8620 18.5605 ;
      RECT 7.8080 17.6250 7.8260 18.5605 ;
      RECT 7.7720 17.8060 7.7900 18.3740 ;
      RECT 8.6990 18.7050 8.7170 19.6405 ;
      RECT 8.6630 18.7050 8.6810 19.6405 ;
      RECT 8.6270 19.2820 8.6450 19.6045 ;
      RECT 8.5100 19.4790 8.5280 19.5885 ;
      RECT 8.5010 18.7375 8.5190 18.9770 ;
      RECT 8.4650 19.3185 8.4830 19.4720 ;
      RECT 8.3840 19.3440 8.4020 19.6020 ;
      RECT 7.8440 18.7050 7.8620 19.6405 ;
      RECT 7.8080 18.7050 7.8260 19.6405 ;
      RECT 7.7720 18.8860 7.7900 19.4540 ;
      RECT 8.6990 19.7850 8.7170 20.7205 ;
      RECT 8.6630 19.7850 8.6810 20.7205 ;
      RECT 8.6270 20.3620 8.6450 20.6845 ;
      RECT 8.5100 20.5590 8.5280 20.6685 ;
      RECT 8.5010 19.8175 8.5190 20.0570 ;
      RECT 8.4650 20.3985 8.4830 20.5520 ;
      RECT 8.3840 20.4240 8.4020 20.6820 ;
      RECT 7.8440 19.7850 7.8620 20.7205 ;
      RECT 7.8080 19.7850 7.8260 20.7205 ;
      RECT 7.7720 19.9660 7.7900 20.5340 ;
      RECT 8.6990 20.8650 8.7170 21.8005 ;
      RECT 8.6630 20.8650 8.6810 21.8005 ;
      RECT 8.6270 21.4420 8.6450 21.7645 ;
      RECT 8.5100 21.6390 8.5280 21.7485 ;
      RECT 8.5010 20.8975 8.5190 21.1370 ;
      RECT 8.4650 21.4785 8.4830 21.6320 ;
      RECT 8.3840 21.5040 8.4020 21.7620 ;
      RECT 7.8440 20.8650 7.8620 21.8005 ;
      RECT 7.8080 20.8650 7.8260 21.8005 ;
      RECT 7.7720 21.0460 7.7900 21.6140 ;
      RECT 8.6990 21.9450 8.7170 22.8805 ;
      RECT 8.6630 21.9450 8.6810 22.8805 ;
      RECT 8.6270 22.5220 8.6450 22.8445 ;
      RECT 8.5100 22.7190 8.5280 22.8285 ;
      RECT 8.5010 21.9775 8.5190 22.2170 ;
      RECT 8.4650 22.5585 8.4830 22.7120 ;
      RECT 8.3840 22.5840 8.4020 22.8420 ;
      RECT 7.8440 21.9450 7.8620 22.8805 ;
      RECT 7.8080 21.9450 7.8260 22.8805 ;
      RECT 7.7720 22.1260 7.7900 22.6940 ;
      RECT 8.6990 23.0250 8.7170 23.9605 ;
      RECT 8.6630 23.0250 8.6810 23.9605 ;
      RECT 8.6270 23.6020 8.6450 23.9245 ;
      RECT 8.5100 23.7990 8.5280 23.9085 ;
      RECT 8.5010 23.0575 8.5190 23.2970 ;
      RECT 8.4650 23.6385 8.4830 23.7920 ;
      RECT 8.3840 23.6640 8.4020 23.9220 ;
      RECT 7.8440 23.0250 7.8620 23.9605 ;
      RECT 7.8080 23.0250 7.8260 23.9605 ;
      RECT 7.7720 23.2060 7.7900 23.7740 ;
      RECT 8.6990 24.1050 8.7170 25.0405 ;
      RECT 8.6630 24.1050 8.6810 25.0405 ;
      RECT 8.6270 24.6820 8.6450 25.0045 ;
      RECT 8.5100 24.8790 8.5280 24.9885 ;
      RECT 8.5010 24.1375 8.5190 24.3770 ;
      RECT 8.4650 24.7185 8.4830 24.8720 ;
      RECT 8.3840 24.7440 8.4020 25.0020 ;
      RECT 7.8440 24.1050 7.8620 25.0405 ;
      RECT 7.8080 24.1050 7.8260 25.0405 ;
      RECT 7.7720 24.2860 7.7900 24.8540 ;
      RECT 8.6990 25.1850 8.7170 26.1205 ;
      RECT 8.6630 25.1850 8.6810 26.1205 ;
      RECT 8.6270 25.7620 8.6450 26.0845 ;
      RECT 8.5100 25.9590 8.5280 26.0685 ;
      RECT 8.5010 25.2175 8.5190 25.4570 ;
      RECT 8.4650 25.7985 8.4830 25.9520 ;
      RECT 8.3840 25.8240 8.4020 26.0820 ;
      RECT 7.8440 25.1850 7.8620 26.1205 ;
      RECT 7.8080 25.1850 7.8260 26.1205 ;
      RECT 7.7720 25.3660 7.7900 25.9340 ;
      RECT 16.3170 29.9500 16.3350 34.3040 ;
      RECT 16.2810 28.6350 16.2990 28.7040 ;
      RECT 16.2810 30.2550 16.2990 30.3380 ;
      RECT 16.2450 26.1305 16.2630 34.3375 ;
      RECT 16.2090 29.9825 16.2270 30.6725 ;
      RECT 16.2090 30.7235 16.2270 31.7100 ;
      RECT 16.2090 31.7500 16.2270 32.3670 ;
      RECT 16.1730 29.9190 16.1910 30.6237 ;
      RECT 16.1730 31.3770 16.1910 32.5470 ;
      RECT 16.1370 26.1305 16.1550 29.7270 ;
      RECT 16.0290 26.1305 16.0470 29.7270 ;
      RECT 15.9210 26.1305 15.9390 29.7270 ;
      RECT 15.8130 26.1305 15.8310 29.7270 ;
      RECT 15.7050 26.1305 15.7230 29.7270 ;
      RECT 15.5970 26.1305 15.6150 29.7270 ;
      RECT 15.4890 26.1305 15.5070 29.7270 ;
      RECT 15.3810 26.1305 15.3990 29.7270 ;
      RECT 15.2730 26.1305 15.2910 29.7270 ;
      RECT 15.1650 26.1305 15.1830 29.7270 ;
      RECT 15.0570 26.1305 15.0750 29.7270 ;
      RECT 14.9490 26.1305 14.9670 29.7270 ;
      RECT 14.8410 26.1305 14.8590 29.7270 ;
      RECT 14.7330 26.1305 14.7510 29.7270 ;
      RECT 14.6250 26.1305 14.6430 29.7270 ;
      RECT 14.5170 26.1305 14.5350 29.7270 ;
      RECT 14.4090 26.1305 14.4270 29.7270 ;
      RECT 14.3010 26.1305 14.3190 29.7270 ;
      RECT 14.1930 26.1305 14.2110 29.7270 ;
      RECT 14.0850 26.1305 14.1030 29.7270 ;
      RECT 13.9770 26.1305 13.9950 29.7270 ;
      RECT 13.8690 26.1305 13.8870 29.7270 ;
      RECT 13.7610 26.1305 13.7790 29.7270 ;
      RECT 13.6530 26.1305 13.6710 29.7270 ;
      RECT 13.5450 26.1305 13.5630 29.7270 ;
      RECT 13.4370 26.1305 13.4550 29.7270 ;
      RECT 13.3290 26.1305 13.3470 29.7270 ;
      RECT 13.2210 26.1305 13.2390 29.7270 ;
      RECT 13.1130 26.1305 13.1310 29.7270 ;
      RECT 13.0050 26.1305 13.0230 29.7270 ;
      RECT 12.8970 26.1305 12.9150 29.7270 ;
      RECT 12.7890 26.1305 12.8070 29.7270 ;
      RECT 12.6810 26.1305 12.6990 29.7270 ;
      RECT 12.5730 26.1305 12.5910 29.7270 ;
      RECT 12.4650 26.1305 12.4830 29.7270 ;
      RECT 12.3570 26.1305 12.3750 29.7270 ;
      RECT 12.2490 26.1305 12.2670 29.7270 ;
      RECT 12.1410 26.1305 12.1590 29.7270 ;
      RECT 12.0330 26.1305 12.0510 29.7270 ;
      RECT 11.9250 26.1305 11.9430 29.7270 ;
      RECT 11.8170 26.1305 11.8350 29.7270 ;
      RECT 11.7090 26.1305 11.7270 29.7270 ;
      RECT 11.6010 26.1305 11.6190 29.7270 ;
      RECT 11.4930 26.1305 11.5110 29.7270 ;
      RECT 11.3850 26.1305 11.4030 29.7270 ;
      RECT 11.2770 26.1305 11.2950 29.7270 ;
      RECT 11.1690 26.1305 11.1870 29.7270 ;
      RECT 11.0610 26.1305 11.0790 29.7270 ;
      RECT 10.9530 26.1305 10.9710 29.7270 ;
      RECT 10.8450 26.1305 10.8630 29.7270 ;
      RECT 10.7370 26.1305 10.7550 29.7270 ;
      RECT 10.6290 26.1305 10.6470 29.7270 ;
      RECT 10.5210 26.1305 10.5390 29.7270 ;
      RECT 10.4130 26.1305 10.4310 29.7270 ;
      RECT 10.3050 26.1305 10.3230 29.7270 ;
      RECT 10.1970 26.1305 10.2150 29.7270 ;
      RECT 10.0890 26.1305 10.1070 29.7270 ;
      RECT 9.9810 26.1305 9.9990 29.7270 ;
      RECT 9.8730 26.1305 9.8910 29.7270 ;
      RECT 9.7650 26.1305 9.7830 29.7270 ;
      RECT 9.6570 26.1305 9.6750 29.7270 ;
      RECT 9.5490 26.1305 9.5670 29.7270 ;
      RECT 9.5130 29.9855 9.5310 30.6275 ;
      RECT 9.5130 31.3050 9.5310 31.8370 ;
      RECT 9.4950 26.7910 9.5130 27.4670 ;
      RECT 9.4950 28.2130 9.5130 28.5110 ;
      RECT 9.4950 29.3290 9.5130 29.5910 ;
      RECT 9.4770 29.9000 9.4950 30.6725 ;
      RECT 9.4770 30.7237 9.4950 31.2150 ;
      RECT 9.4770 31.2600 9.4950 31.6310 ;
      RECT 9.4770 31.7070 9.4950 32.3670 ;
      RECT 9.4410 26.1305 9.4590 34.3375 ;
      RECT 9.4050 30.4430 9.4230 30.9075 ;
      RECT 9.3870 26.8990 9.4050 27.5300 ;
      RECT 9.3870 27.9430 9.4050 28.1330 ;
      RECT 9.3870 28.8250 9.4050 28.8740 ;
      RECT 9.3870 29.5570 9.4050 29.5940 ;
      RECT 9.3690 29.9500 9.3870 34.2995 ;
      RECT 9.2790 26.5210 9.2970 27.3230 ;
      RECT 9.2790 27.8710 9.2970 28.4390 ;
      RECT 9.2430 27.9430 9.2610 28.3130 ;
      RECT 9.2070 27.2950 9.2250 27.4310 ;
      RECT 9.2070 28.2850 9.2250 28.5110 ;
      RECT 9.2070 29.5270 9.2250 29.5910 ;
      RECT 9.1710 27.3970 9.1890 27.4340 ;
      RECT 9.1710 29.0230 9.1890 29.0660 ;
      RECT 9.1710 29.5570 9.1890 29.5940 ;
      RECT 9.1350 27.7090 9.1530 28.2050 ;
      RECT 9.1350 28.2490 9.1530 28.4390 ;
      RECT 9.1350 29.2090 9.1530 29.5190 ;
      RECT 9.0990 27.6010 9.1170 28.8480 ;
      RECT 9.0990 31.4890 9.1170 32.2190 ;
      RECT 9.0990 32.5690 9.1170 33.2990 ;
      RECT 8.7750 27.3310 8.7930 27.6290 ;
      RECT 8.7750 28.5190 8.7930 28.5830 ;
      RECT 8.7750 28.7890 8.7930 29.2490 ;
      RECT 8.7750 29.9890 8.7930 30.0260 ;
      RECT 8.7750 32.0290 8.7930 32.3270 ;
      RECT 8.7390 27.4030 8.7570 27.9080 ;
      RECT 8.7390 28.1770 8.7570 28.9790 ;
      RECT 8.7390 30.0220 8.7570 30.2930 ;
      RECT 8.7390 30.3730 8.7570 30.5990 ;
      RECT 8.7030 27.3310 8.7210 28.0070 ;
      RECT 8.7030 28.1050 8.7210 28.4390 ;
      RECT 8.7030 28.6450 8.7210 28.7810 ;
      RECT 8.7030 29.3290 8.7210 30.1310 ;
      RECT 8.7030 30.5650 8.7210 30.6020 ;
      RECT 8.7030 32.7310 8.7210 33.0650 ;
      RECT 8.6670 27.5650 8.6850 27.7010 ;
      RECT 8.6670 29.4550 8.6850 30.4370 ;
      RECT 8.6670 30.8770 8.6850 31.1750 ;
      RECT 8.6670 32.5690 8.6850 32.8310 ;
      RECT 8.6310 26.6290 8.6490 26.7830 ;
      RECT 8.6310 27.4390 8.6490 29.2250 ;
      RECT 8.6310 30.2650 8.6490 32.5970 ;
      RECT 8.6310 32.8030 8.6490 33.9110 ;
      RECT 8.3430 26.8990 8.3610 27.1610 ;
      RECT 8.3430 27.2950 8.3610 27.3590 ;
      RECT 8.3430 27.4390 8.3610 27.6650 ;
      RECT 8.3430 27.7090 8.3610 27.8990 ;
      RECT 8.3430 27.9790 8.3610 30.5990 ;
      RECT 8.3430 30.6430 8.3610 31.9490 ;
      RECT 8.3430 33.0370 8.3610 33.2990 ;
      RECT 8.3070 27.8980 8.3250 28.1690 ;
      RECT 8.3070 28.2490 8.3250 29.0870 ;
      RECT 8.3070 29.2570 8.3250 30.0950 ;
      RECT 8.3070 30.1390 8.3250 31.4090 ;
      RECT 8.3070 31.6150 8.3250 31.7870 ;
      RECT 8.3070 32.4970 8.3250 33.5690 ;
      RECT 8.2710 27.9790 8.2890 28.2500 ;
      RECT 8.2710 28.4050 8.2890 28.4420 ;
      RECT 8.2710 29.1850 8.2890 30.1670 ;
      RECT 8.2710 30.4090 8.2890 30.8690 ;
      RECT 8.2710 31.2190 8.2890 31.9580 ;
      RECT 8.2350 27.0970 8.2530 28.1690 ;
      RECT 8.2350 29.7610 8.2530 29.9780 ;
      RECT 8.2350 31.1470 8.2530 31.4450 ;
      RECT 8.1990 27.7450 8.2170 28.2050 ;
      RECT 8.1990 29.3290 8.2170 29.5190 ;
      RECT 8.1990 29.5600 8.2170 29.5970 ;
      RECT 8.1990 29.8330 8.2170 30.1670 ;
      RECT 8.1990 30.3010 8.2170 31.6430 ;
      RECT 8.1990 31.7500 8.2170 32.8670 ;
      RECT 8.1630 27.1690 8.1810 27.3590 ;
      RECT 8.1630 27.5650 8.1810 27.7010 ;
      RECT 8.1630 27.9790 8.1810 31.1390 ;
      RECT 8.1630 31.2190 8.1810 31.6790 ;
      RECT 8.1630 32.2990 8.1810 32.7590 ;
      RECT 8.1630 33.6130 8.1810 33.8390 ;
      RECT 8.1270 26.1570 8.1450 26.3110 ;
      RECT 8.1270 34.1520 8.1450 34.3180 ;
      RECT 8.0910 26.1570 8.1090 26.2070 ;
      RECT 8.0190 26.1570 8.0370 26.2285 ;
      RECT 8.0190 34.2215 8.0370 34.3375 ;
      RECT 7.8750 27.6730 7.8930 27.8630 ;
      RECT 7.8750 28.4110 7.8930 28.7810 ;
      RECT 7.8750 30.3730 7.8930 30.5990 ;
      RECT 7.8750 30.9130 7.8930 32.0570 ;
      RECT 7.8750 32.8390 7.8930 33.2990 ;
      RECT 7.8750 33.8770 7.8930 33.9140 ;
      RECT 7.8390 26.6290 7.8570 27.1250 ;
      RECT 7.8390 30.7090 7.8570 30.7460 ;
      RECT 7.8390 31.7860 7.8570 32.5970 ;
      RECT 7.8030 27.0970 7.8210 27.3590 ;
      RECT 7.8030 27.6370 7.8210 27.9710 ;
      RECT 7.8030 28.1770 7.8210 28.2770 ;
      RECT 7.8030 29.0590 7.8210 31.8230 ;
      RECT 7.8030 31.9570 7.8210 32.1830 ;
      RECT 7.7670 26.7550 7.7850 27.8990 ;
      RECT 7.7670 31.4890 7.7850 31.6790 ;
      RECT 7.7670 32.2930 7.7850 32.3300 ;
      RECT 7.7670 32.5690 7.7850 33.3710 ;
      RECT 7.7310 27.7090 7.7490 28.7090 ;
      RECT 7.7310 32.1490 7.7490 32.1860 ;
      RECT 7.3710 27.2950 7.3890 27.7010 ;
      RECT 7.2990 27.3310 7.3170 27.9350 ;
      RECT 7.2630 27.1690 7.2810 27.2330 ;
      RECT 7.2270 26.2100 7.2450 26.2610 ;
      RECT 7.2270 29.3290 7.2450 29.5190 ;
      RECT 7.2090 29.9500 7.2270 34.2985 ;
      RECT 7.1370 29.9500 7.1550 34.2995 ;
      RECT 7.1190 26.6290 7.1370 26.8190 ;
      RECT 7.1190 27.4030 7.1370 29.6630 ;
      RECT 7.1010 30.4430 7.1190 30.9075 ;
      RECT 7.0650 26.1305 7.0830 34.3375 ;
      RECT 7.0290 29.9000 7.0470 30.6725 ;
      RECT 7.0290 30.7237 7.0470 31.2150 ;
      RECT 7.0290 31.2600 7.0470 31.6310 ;
      RECT 7.0290 31.7070 7.0470 32.3670 ;
      RECT 7.0110 26.6290 7.0290 27.1250 ;
      RECT 7.0110 27.9070 7.0290 28.4750 ;
      RECT 7.0110 28.7890 7.0290 29.5190 ;
      RECT 6.9930 29.9855 7.0110 30.6275 ;
      RECT 6.9930 31.3050 7.0110 31.8370 ;
      RECT 6.9570 26.1305 6.9750 29.7270 ;
      RECT 6.8490 26.1305 6.8670 29.7270 ;
      RECT 6.7410 26.1305 6.7590 29.7270 ;
      RECT 6.6330 26.1305 6.6510 29.7270 ;
      RECT 6.5250 26.1305 6.5430 29.7270 ;
      RECT 6.4170 26.1305 6.4350 29.7270 ;
      RECT 6.3090 26.1305 6.3270 29.7270 ;
      RECT 6.2010 26.1305 6.2190 29.7270 ;
      RECT 6.0930 26.1305 6.1110 29.7270 ;
      RECT 5.9850 26.1305 6.0030 29.7270 ;
      RECT 5.8770 26.1305 5.8950 29.7270 ;
      RECT 5.7690 26.1305 5.7870 29.7270 ;
      RECT 5.6610 26.1305 5.6790 29.7270 ;
      RECT 5.5530 26.1305 5.5710 29.7270 ;
      RECT 5.4450 26.1305 5.4630 29.7270 ;
      RECT 5.3370 26.1305 5.3550 29.7270 ;
      RECT 5.2290 26.1305 5.2470 29.7270 ;
      RECT 5.1210 26.1305 5.1390 29.7270 ;
      RECT 5.0130 26.1305 5.0310 29.7270 ;
      RECT 4.9050 26.1305 4.9230 29.7270 ;
      RECT 4.7970 26.1305 4.8150 29.7270 ;
      RECT 4.6890 26.1305 4.7070 29.7270 ;
      RECT 4.5810 26.1305 4.5990 29.7270 ;
      RECT 4.4730 26.1305 4.4910 29.7270 ;
      RECT 4.3650 26.1305 4.3830 29.7270 ;
      RECT 4.2570 26.1305 4.2750 29.7270 ;
      RECT 4.1490 26.1305 4.1670 29.7270 ;
      RECT 4.0410 26.1305 4.0590 29.7270 ;
      RECT 3.9330 26.1305 3.9510 29.7270 ;
      RECT 3.8250 26.1305 3.8430 29.7270 ;
      RECT 3.7170 26.1305 3.7350 29.7270 ;
      RECT 3.6090 26.1305 3.6270 29.7270 ;
      RECT 3.5010 26.1305 3.5190 29.7270 ;
      RECT 3.3930 26.1305 3.4110 29.7270 ;
      RECT 3.2850 26.1305 3.3030 29.7270 ;
      RECT 3.1770 26.1305 3.1950 29.7270 ;
      RECT 3.0690 26.1305 3.0870 29.7270 ;
      RECT 2.9610 26.1305 2.9790 29.7270 ;
      RECT 2.8530 26.1305 2.8710 29.7270 ;
      RECT 2.7450 26.1305 2.7630 29.7270 ;
      RECT 2.6370 26.1305 2.6550 29.7270 ;
      RECT 2.5290 26.1305 2.5470 29.7270 ;
      RECT 2.4210 26.1305 2.4390 29.7270 ;
      RECT 2.3130 26.1305 2.3310 29.7270 ;
      RECT 2.2050 26.1305 2.2230 29.7270 ;
      RECT 2.0970 26.1305 2.1150 29.7270 ;
      RECT 1.9890 26.1305 2.0070 29.7270 ;
      RECT 1.8810 26.1305 1.8990 29.7270 ;
      RECT 1.7730 26.1305 1.7910 29.7270 ;
      RECT 1.6650 26.1305 1.6830 29.7270 ;
      RECT 1.5570 26.1305 1.5750 29.7270 ;
      RECT 1.4490 26.1305 1.4670 29.7270 ;
      RECT 1.3410 26.1305 1.3590 29.7270 ;
      RECT 1.2330 26.1305 1.2510 29.7270 ;
      RECT 1.1250 26.1305 1.1430 29.7270 ;
      RECT 1.0170 26.1305 1.0350 29.7270 ;
      RECT 0.9090 26.1305 0.9270 29.7270 ;
      RECT 0.8010 26.1305 0.8190 29.7270 ;
      RECT 0.6930 26.1305 0.7110 29.7270 ;
      RECT 0.5850 26.1305 0.6030 29.7270 ;
      RECT 0.4770 26.1305 0.4950 29.7270 ;
      RECT 0.3690 26.1305 0.3870 29.7270 ;
      RECT 0.3330 29.9190 0.3510 30.6237 ;
      RECT 0.3330 31.3770 0.3510 32.5470 ;
      RECT 0.2970 29.9825 0.3150 30.6725 ;
      RECT 0.2970 30.7235 0.3150 31.7100 ;
      RECT 0.2970 31.7500 0.3150 32.3670 ;
      RECT 0.2610 26.1305 0.2790 34.3375 ;
      RECT 0.2250 28.6350 0.2430 28.7040 ;
      RECT 0.2250 30.2550 0.2430 30.3380 ;
      RECT 0.1890 29.9500 0.2070 34.3040 ;
        RECT 8.6990 34.3920 8.7170 35.3275 ;
        RECT 8.6630 34.3920 8.6810 35.3275 ;
        RECT 8.6270 34.9690 8.6450 35.2915 ;
        RECT 8.5100 35.1660 8.5280 35.2755 ;
        RECT 8.5010 34.4245 8.5190 34.6640 ;
        RECT 8.4650 35.0055 8.4830 35.1590 ;
        RECT 8.3840 35.0310 8.4020 35.2890 ;
        RECT 7.8440 34.3920 7.8620 35.3275 ;
        RECT 7.8080 34.3920 7.8260 35.3275 ;
        RECT 7.7720 34.5730 7.7900 35.1410 ;
        RECT 8.6990 35.4720 8.7170 36.4075 ;
        RECT 8.6630 35.4720 8.6810 36.4075 ;
        RECT 8.6270 36.0490 8.6450 36.3715 ;
        RECT 8.5100 36.2460 8.5280 36.3555 ;
        RECT 8.5010 35.5045 8.5190 35.7440 ;
        RECT 8.4650 36.0855 8.4830 36.2390 ;
        RECT 8.3840 36.1110 8.4020 36.3690 ;
        RECT 7.8440 35.4720 7.8620 36.4075 ;
        RECT 7.8080 35.4720 7.8260 36.4075 ;
        RECT 7.7720 35.6530 7.7900 36.2210 ;
        RECT 8.6990 36.5520 8.7170 37.4875 ;
        RECT 8.6630 36.5520 8.6810 37.4875 ;
        RECT 8.6270 37.1290 8.6450 37.4515 ;
        RECT 8.5100 37.3260 8.5280 37.4355 ;
        RECT 8.5010 36.5845 8.5190 36.8240 ;
        RECT 8.4650 37.1655 8.4830 37.3190 ;
        RECT 8.3840 37.1910 8.4020 37.4490 ;
        RECT 7.8440 36.5520 7.8620 37.4875 ;
        RECT 7.8080 36.5520 7.8260 37.4875 ;
        RECT 7.7720 36.7330 7.7900 37.3010 ;
        RECT 8.6990 37.6320 8.7170 38.5675 ;
        RECT 8.6630 37.6320 8.6810 38.5675 ;
        RECT 8.6270 38.2090 8.6450 38.5315 ;
        RECT 8.5100 38.4060 8.5280 38.5155 ;
        RECT 8.5010 37.6645 8.5190 37.9040 ;
        RECT 8.4650 38.2455 8.4830 38.3990 ;
        RECT 8.3840 38.2710 8.4020 38.5290 ;
        RECT 7.8440 37.6320 7.8620 38.5675 ;
        RECT 7.8080 37.6320 7.8260 38.5675 ;
        RECT 7.7720 37.8130 7.7900 38.3810 ;
        RECT 8.6990 38.7120 8.7170 39.6475 ;
        RECT 8.6630 38.7120 8.6810 39.6475 ;
        RECT 8.6270 39.2890 8.6450 39.6115 ;
        RECT 8.5100 39.4860 8.5280 39.5955 ;
        RECT 8.5010 38.7445 8.5190 38.9840 ;
        RECT 8.4650 39.3255 8.4830 39.4790 ;
        RECT 8.3840 39.3510 8.4020 39.6090 ;
        RECT 7.8440 38.7120 7.8620 39.6475 ;
        RECT 7.8080 38.7120 7.8260 39.6475 ;
        RECT 7.7720 38.8930 7.7900 39.4610 ;
        RECT 8.6990 39.7920 8.7170 40.7275 ;
        RECT 8.6630 39.7920 8.6810 40.7275 ;
        RECT 8.6270 40.3690 8.6450 40.6915 ;
        RECT 8.5100 40.5660 8.5280 40.6755 ;
        RECT 8.5010 39.8245 8.5190 40.0640 ;
        RECT 8.4650 40.4055 8.4830 40.5590 ;
        RECT 8.3840 40.4310 8.4020 40.6890 ;
        RECT 7.8440 39.7920 7.8620 40.7275 ;
        RECT 7.8080 39.7920 7.8260 40.7275 ;
        RECT 7.7720 39.9730 7.7900 40.5410 ;
        RECT 8.6990 40.8720 8.7170 41.8075 ;
        RECT 8.6630 40.8720 8.6810 41.8075 ;
        RECT 8.6270 41.4490 8.6450 41.7715 ;
        RECT 8.5100 41.6460 8.5280 41.7555 ;
        RECT 8.5010 40.9045 8.5190 41.1440 ;
        RECT 8.4650 41.4855 8.4830 41.6390 ;
        RECT 8.3840 41.5110 8.4020 41.7690 ;
        RECT 7.8440 40.8720 7.8620 41.8075 ;
        RECT 7.8080 40.8720 7.8260 41.8075 ;
        RECT 7.7720 41.0530 7.7900 41.6210 ;
        RECT 8.6990 41.9520 8.7170 42.8875 ;
        RECT 8.6630 41.9520 8.6810 42.8875 ;
        RECT 8.6270 42.5290 8.6450 42.8515 ;
        RECT 8.5100 42.7260 8.5280 42.8355 ;
        RECT 8.5010 41.9845 8.5190 42.2240 ;
        RECT 8.4650 42.5655 8.4830 42.7190 ;
        RECT 8.3840 42.5910 8.4020 42.8490 ;
        RECT 7.8440 41.9520 7.8620 42.8875 ;
        RECT 7.8080 41.9520 7.8260 42.8875 ;
        RECT 7.7720 42.1330 7.7900 42.7010 ;
        RECT 8.6990 43.0320 8.7170 43.9675 ;
        RECT 8.6630 43.0320 8.6810 43.9675 ;
        RECT 8.6270 43.6090 8.6450 43.9315 ;
        RECT 8.5100 43.8060 8.5280 43.9155 ;
        RECT 8.5010 43.0645 8.5190 43.3040 ;
        RECT 8.4650 43.6455 8.4830 43.7990 ;
        RECT 8.3840 43.6710 8.4020 43.9290 ;
        RECT 7.8440 43.0320 7.8620 43.9675 ;
        RECT 7.8080 43.0320 7.8260 43.9675 ;
        RECT 7.7720 43.2130 7.7900 43.7810 ;
        RECT 8.6990 44.1120 8.7170 45.0475 ;
        RECT 8.6630 44.1120 8.6810 45.0475 ;
        RECT 8.6270 44.6890 8.6450 45.0115 ;
        RECT 8.5100 44.8860 8.5280 44.9955 ;
        RECT 8.5010 44.1445 8.5190 44.3840 ;
        RECT 8.4650 44.7255 8.4830 44.8790 ;
        RECT 8.3840 44.7510 8.4020 45.0090 ;
        RECT 7.8440 44.1120 7.8620 45.0475 ;
        RECT 7.8080 44.1120 7.8260 45.0475 ;
        RECT 7.7720 44.2930 7.7900 44.8610 ;
        RECT 8.6990 45.1920 8.7170 46.1275 ;
        RECT 8.6630 45.1920 8.6810 46.1275 ;
        RECT 8.6270 45.7690 8.6450 46.0915 ;
        RECT 8.5100 45.9660 8.5280 46.0755 ;
        RECT 8.5010 45.2245 8.5190 45.4640 ;
        RECT 8.4650 45.8055 8.4830 45.9590 ;
        RECT 8.3840 45.8310 8.4020 46.0890 ;
        RECT 7.8440 45.1920 7.8620 46.1275 ;
        RECT 7.8080 45.1920 7.8260 46.1275 ;
        RECT 7.7720 45.3730 7.7900 45.9410 ;
        RECT 8.6990 46.2720 8.7170 47.2075 ;
        RECT 8.6630 46.2720 8.6810 47.2075 ;
        RECT 8.6270 46.8490 8.6450 47.1715 ;
        RECT 8.5100 47.0460 8.5280 47.1555 ;
        RECT 8.5010 46.3045 8.5190 46.5440 ;
        RECT 8.4650 46.8855 8.4830 47.0390 ;
        RECT 8.3840 46.9110 8.4020 47.1690 ;
        RECT 7.8440 46.2720 7.8620 47.2075 ;
        RECT 7.8080 46.2720 7.8260 47.2075 ;
        RECT 7.7720 46.4530 7.7900 47.0210 ;
        RECT 8.6990 47.3520 8.7170 48.2875 ;
        RECT 8.6630 47.3520 8.6810 48.2875 ;
        RECT 8.6270 47.9290 8.6450 48.2515 ;
        RECT 8.5100 48.1260 8.5280 48.2355 ;
        RECT 8.5010 47.3845 8.5190 47.6240 ;
        RECT 8.4650 47.9655 8.4830 48.1190 ;
        RECT 8.3840 47.9910 8.4020 48.2490 ;
        RECT 7.8440 47.3520 7.8620 48.2875 ;
        RECT 7.8080 47.3520 7.8260 48.2875 ;
        RECT 7.7720 47.5330 7.7900 48.1010 ;
        RECT 8.6990 48.4320 8.7170 49.3675 ;
        RECT 8.6630 48.4320 8.6810 49.3675 ;
        RECT 8.6270 49.0090 8.6450 49.3315 ;
        RECT 8.5100 49.2060 8.5280 49.3155 ;
        RECT 8.5010 48.4645 8.5190 48.7040 ;
        RECT 8.4650 49.0455 8.4830 49.1990 ;
        RECT 8.3840 49.0710 8.4020 49.3290 ;
        RECT 7.8440 48.4320 7.8620 49.3675 ;
        RECT 7.8080 48.4320 7.8260 49.3675 ;
        RECT 7.7720 48.6130 7.7900 49.1810 ;
        RECT 8.6990 49.5120 8.7170 50.4475 ;
        RECT 8.6630 49.5120 8.6810 50.4475 ;
        RECT 8.6270 50.0890 8.6450 50.4115 ;
        RECT 8.5100 50.2860 8.5280 50.3955 ;
        RECT 8.5010 49.5445 8.5190 49.7840 ;
        RECT 8.4650 50.1255 8.4830 50.2790 ;
        RECT 8.3840 50.1510 8.4020 50.4090 ;
        RECT 7.8440 49.5120 7.8620 50.4475 ;
        RECT 7.8080 49.5120 7.8260 50.4475 ;
        RECT 7.7720 49.6930 7.7900 50.2610 ;
        RECT 8.6990 50.5920 8.7170 51.5275 ;
        RECT 8.6630 50.5920 8.6810 51.5275 ;
        RECT 8.6270 51.1690 8.6450 51.4915 ;
        RECT 8.5100 51.3660 8.5280 51.4755 ;
        RECT 8.5010 50.6245 8.5190 50.8640 ;
        RECT 8.4650 51.2055 8.4830 51.3590 ;
        RECT 8.3840 51.2310 8.4020 51.4890 ;
        RECT 7.8440 50.5920 7.8620 51.5275 ;
        RECT 7.8080 50.5920 7.8260 51.5275 ;
        RECT 7.7720 50.7730 7.7900 51.3410 ;
        RECT 8.6990 51.6720 8.7170 52.6075 ;
        RECT 8.6630 51.6720 8.6810 52.6075 ;
        RECT 8.6270 52.2490 8.6450 52.5715 ;
        RECT 8.5100 52.4460 8.5280 52.5555 ;
        RECT 8.5010 51.7045 8.5190 51.9440 ;
        RECT 8.4650 52.2855 8.4830 52.4390 ;
        RECT 8.3840 52.3110 8.4020 52.5690 ;
        RECT 7.8440 51.6720 7.8620 52.6075 ;
        RECT 7.8080 51.6720 7.8260 52.6075 ;
        RECT 7.7720 51.8530 7.7900 52.4210 ;
        RECT 8.6990 52.7520 8.7170 53.6875 ;
        RECT 8.6630 52.7520 8.6810 53.6875 ;
        RECT 8.6270 53.3290 8.6450 53.6515 ;
        RECT 8.5100 53.5260 8.5280 53.6355 ;
        RECT 8.5010 52.7845 8.5190 53.0240 ;
        RECT 8.4650 53.3655 8.4830 53.5190 ;
        RECT 8.3840 53.3910 8.4020 53.6490 ;
        RECT 7.8440 52.7520 7.8620 53.6875 ;
        RECT 7.8080 52.7520 7.8260 53.6875 ;
        RECT 7.7720 52.9330 7.7900 53.5010 ;
        RECT 8.6990 53.8320 8.7170 54.7675 ;
        RECT 8.6630 53.8320 8.6810 54.7675 ;
        RECT 8.6270 54.4090 8.6450 54.7315 ;
        RECT 8.5100 54.6060 8.5280 54.7155 ;
        RECT 8.5010 53.8645 8.5190 54.1040 ;
        RECT 8.4650 54.4455 8.4830 54.5990 ;
        RECT 8.3840 54.4710 8.4020 54.7290 ;
        RECT 7.8440 53.8320 7.8620 54.7675 ;
        RECT 7.8080 53.8320 7.8260 54.7675 ;
        RECT 7.7720 54.0130 7.7900 54.5810 ;
        RECT 8.6990 54.9120 8.7170 55.8475 ;
        RECT 8.6630 54.9120 8.6810 55.8475 ;
        RECT 8.6270 55.4890 8.6450 55.8115 ;
        RECT 8.5100 55.6860 8.5280 55.7955 ;
        RECT 8.5010 54.9445 8.5190 55.1840 ;
        RECT 8.4650 55.5255 8.4830 55.6790 ;
        RECT 8.3840 55.5510 8.4020 55.8090 ;
        RECT 7.8440 54.9120 7.8620 55.8475 ;
        RECT 7.8080 54.9120 7.8260 55.8475 ;
        RECT 7.7720 55.0930 7.7900 55.6610 ;
        RECT 8.6990 55.9920 8.7170 56.9275 ;
        RECT 8.6630 55.9920 8.6810 56.9275 ;
        RECT 8.6270 56.5690 8.6450 56.8915 ;
        RECT 8.5100 56.7660 8.5280 56.8755 ;
        RECT 8.5010 56.0245 8.5190 56.2640 ;
        RECT 8.4650 56.6055 8.4830 56.7590 ;
        RECT 8.3840 56.6310 8.4020 56.8890 ;
        RECT 7.8440 55.9920 7.8620 56.9275 ;
        RECT 7.8080 55.9920 7.8260 56.9275 ;
        RECT 7.7720 56.1730 7.7900 56.7410 ;
        RECT 8.6990 57.0720 8.7170 58.0075 ;
        RECT 8.6630 57.0720 8.6810 58.0075 ;
        RECT 8.6270 57.6490 8.6450 57.9715 ;
        RECT 8.5100 57.8460 8.5280 57.9555 ;
        RECT 8.5010 57.1045 8.5190 57.3440 ;
        RECT 8.4650 57.6855 8.4830 57.8390 ;
        RECT 8.3840 57.7110 8.4020 57.9690 ;
        RECT 7.8440 57.0720 7.8620 58.0075 ;
        RECT 7.8080 57.0720 7.8260 58.0075 ;
        RECT 7.7720 57.2530 7.7900 57.8210 ;
        RECT 8.6990 58.1520 8.7170 59.0875 ;
        RECT 8.6630 58.1520 8.6810 59.0875 ;
        RECT 8.6270 58.7290 8.6450 59.0515 ;
        RECT 8.5100 58.9260 8.5280 59.0355 ;
        RECT 8.5010 58.1845 8.5190 58.4240 ;
        RECT 8.4650 58.7655 8.4830 58.9190 ;
        RECT 8.3840 58.7910 8.4020 59.0490 ;
        RECT 7.8440 58.1520 7.8620 59.0875 ;
        RECT 7.8080 58.1520 7.8260 59.0875 ;
        RECT 7.7720 58.3330 7.7900 58.9010 ;
        RECT 8.6990 59.2320 8.7170 60.1675 ;
        RECT 8.6630 59.2320 8.6810 60.1675 ;
        RECT 8.6270 59.8090 8.6450 60.1315 ;
        RECT 8.5100 60.0060 8.5280 60.1155 ;
        RECT 8.5010 59.2645 8.5190 59.5040 ;
        RECT 8.4650 59.8455 8.4830 59.9990 ;
        RECT 8.3840 59.8710 8.4020 60.1290 ;
        RECT 7.8440 59.2320 7.8620 60.1675 ;
        RECT 7.8080 59.2320 7.8260 60.1675 ;
        RECT 7.7720 59.4130 7.7900 59.9810 ;
  LAYER M3 SPACING 0.018  ;
      RECT 8.6410 0.2565 8.7690 1.3500 ;
      RECT 8.6270 0.9220 8.7690 1.2445 ;
      RECT 8.4790 0.6490 8.5410 1.3500 ;
      RECT 8.4650 0.9585 8.5410 1.1120 ;
      RECT 8.4790 0.2565 8.5050 1.3500 ;
      RECT 8.4790 0.3775 8.5190 0.6170 ;
      RECT 8.4790 0.2565 8.5410 0.3455 ;
      RECT 8.1820 0.7070 8.3880 1.3500 ;
      RECT 8.3620 0.2565 8.3880 1.3500 ;
      RECT 8.1820 0.9840 8.4020 1.2420 ;
      RECT 8.1820 0.2565 8.2800 1.3500 ;
      RECT 7.7650 0.2565 7.8480 1.3500 ;
      RECT 7.7650 0.3450 7.8620 1.2805 ;
      RECT 16.4440 0.2565 16.5290 1.3500 ;
      RECT 16.3000 0.2565 16.3260 1.3500 ;
      RECT 16.1920 0.2565 16.2180 1.3500 ;
      RECT 16.0840 0.2565 16.1100 1.3500 ;
      RECT 15.9760 0.2565 16.0020 1.3500 ;
      RECT 15.8680 0.2565 15.8940 1.3500 ;
      RECT 15.7600 0.2565 15.7860 1.3500 ;
      RECT 15.6520 0.2565 15.6780 1.3500 ;
      RECT 15.5440 0.2565 15.5700 1.3500 ;
      RECT 15.4360 0.2565 15.4620 1.3500 ;
      RECT 15.3280 0.2565 15.3540 1.3500 ;
      RECT 15.2200 0.2565 15.2460 1.3500 ;
      RECT 15.1120 0.2565 15.1380 1.3500 ;
      RECT 15.0040 0.2565 15.0300 1.3500 ;
      RECT 14.8960 0.2565 14.9220 1.3500 ;
      RECT 14.7880 0.2565 14.8140 1.3500 ;
      RECT 14.6800 0.2565 14.7060 1.3500 ;
      RECT 14.5720 0.2565 14.5980 1.3500 ;
      RECT 14.4640 0.2565 14.4900 1.3500 ;
      RECT 14.3560 0.2565 14.3820 1.3500 ;
      RECT 14.2480 0.2565 14.2740 1.3500 ;
      RECT 14.1400 0.2565 14.1660 1.3500 ;
      RECT 14.0320 0.2565 14.0580 1.3500 ;
      RECT 13.9240 0.2565 13.9500 1.3500 ;
      RECT 13.8160 0.2565 13.8420 1.3500 ;
      RECT 13.7080 0.2565 13.7340 1.3500 ;
      RECT 13.6000 0.2565 13.6260 1.3500 ;
      RECT 13.4920 0.2565 13.5180 1.3500 ;
      RECT 13.3840 0.2565 13.4100 1.3500 ;
      RECT 13.2760 0.2565 13.3020 1.3500 ;
      RECT 13.1680 0.2565 13.1940 1.3500 ;
      RECT 13.0600 0.2565 13.0860 1.3500 ;
      RECT 12.9520 0.2565 12.9780 1.3500 ;
      RECT 12.8440 0.2565 12.8700 1.3500 ;
      RECT 12.7360 0.2565 12.7620 1.3500 ;
      RECT 12.6280 0.2565 12.6540 1.3500 ;
      RECT 12.5200 0.2565 12.5460 1.3500 ;
      RECT 12.4120 0.2565 12.4380 1.3500 ;
      RECT 12.3040 0.2565 12.3300 1.3500 ;
      RECT 12.1960 0.2565 12.2220 1.3500 ;
      RECT 12.0880 0.2565 12.1140 1.3500 ;
      RECT 11.9800 0.2565 12.0060 1.3500 ;
      RECT 11.8720 0.2565 11.8980 1.3500 ;
      RECT 11.7640 0.2565 11.7900 1.3500 ;
      RECT 11.6560 0.2565 11.6820 1.3500 ;
      RECT 11.5480 0.2565 11.5740 1.3500 ;
      RECT 11.4400 0.2565 11.4660 1.3500 ;
      RECT 11.3320 0.2565 11.3580 1.3500 ;
      RECT 11.2240 0.2565 11.2500 1.3500 ;
      RECT 11.1160 0.2565 11.1420 1.3500 ;
      RECT 11.0080 0.2565 11.0340 1.3500 ;
      RECT 10.9000 0.2565 10.9260 1.3500 ;
      RECT 10.7920 0.2565 10.8180 1.3500 ;
      RECT 10.6840 0.2565 10.7100 1.3500 ;
      RECT 10.5760 0.2565 10.6020 1.3500 ;
      RECT 10.4680 0.2565 10.4940 1.3500 ;
      RECT 10.3600 0.2565 10.3860 1.3500 ;
      RECT 10.2520 0.2565 10.2780 1.3500 ;
      RECT 10.1440 0.2565 10.1700 1.3500 ;
      RECT 10.0360 0.2565 10.0620 1.3500 ;
      RECT 9.9280 0.2565 9.9540 1.3500 ;
      RECT 9.8200 0.2565 9.8460 1.3500 ;
      RECT 9.7120 0.2565 9.7380 1.3500 ;
      RECT 9.6040 0.2565 9.6300 1.3500 ;
      RECT 9.4960 0.2565 9.5220 1.3500 ;
      RECT 9.3880 0.2565 9.4140 1.3500 ;
      RECT 9.1750 0.2565 9.2520 1.3500 ;
      RECT 7.2820 0.2565 7.3590 1.3500 ;
      RECT 7.1200 0.2565 7.1460 1.3500 ;
      RECT 7.0120 0.2565 7.0380 1.3500 ;
      RECT 6.9040 0.2565 6.9300 1.3500 ;
      RECT 6.7960 0.2565 6.8220 1.3500 ;
      RECT 6.6880 0.2565 6.7140 1.3500 ;
      RECT 6.5800 0.2565 6.6060 1.3500 ;
      RECT 6.4720 0.2565 6.4980 1.3500 ;
      RECT 6.3640 0.2565 6.3900 1.3500 ;
      RECT 6.2560 0.2565 6.2820 1.3500 ;
      RECT 6.1480 0.2565 6.1740 1.3500 ;
      RECT 6.0400 0.2565 6.0660 1.3500 ;
      RECT 5.9320 0.2565 5.9580 1.3500 ;
      RECT 5.8240 0.2565 5.8500 1.3500 ;
      RECT 5.7160 0.2565 5.7420 1.3500 ;
      RECT 5.6080 0.2565 5.6340 1.3500 ;
      RECT 5.5000 0.2565 5.5260 1.3500 ;
      RECT 5.3920 0.2565 5.4180 1.3500 ;
      RECT 5.2840 0.2565 5.3100 1.3500 ;
      RECT 5.1760 0.2565 5.2020 1.3500 ;
      RECT 5.0680 0.2565 5.0940 1.3500 ;
      RECT 4.9600 0.2565 4.9860 1.3500 ;
      RECT 4.8520 0.2565 4.8780 1.3500 ;
      RECT 4.7440 0.2565 4.7700 1.3500 ;
      RECT 4.6360 0.2565 4.6620 1.3500 ;
      RECT 4.5280 0.2565 4.5540 1.3500 ;
      RECT 4.4200 0.2565 4.4460 1.3500 ;
      RECT 4.3120 0.2565 4.3380 1.3500 ;
      RECT 4.2040 0.2565 4.2300 1.3500 ;
      RECT 4.0960 0.2565 4.1220 1.3500 ;
      RECT 3.9880 0.2565 4.0140 1.3500 ;
      RECT 3.8800 0.2565 3.9060 1.3500 ;
      RECT 3.7720 0.2565 3.7980 1.3500 ;
      RECT 3.6640 0.2565 3.6900 1.3500 ;
      RECT 3.5560 0.2565 3.5820 1.3500 ;
      RECT 3.4480 0.2565 3.4740 1.3500 ;
      RECT 3.3400 0.2565 3.3660 1.3500 ;
      RECT 3.2320 0.2565 3.2580 1.3500 ;
      RECT 3.1240 0.2565 3.1500 1.3500 ;
      RECT 3.0160 0.2565 3.0420 1.3500 ;
      RECT 2.9080 0.2565 2.9340 1.3500 ;
      RECT 2.8000 0.2565 2.8260 1.3500 ;
      RECT 2.6920 0.2565 2.7180 1.3500 ;
      RECT 2.5840 0.2565 2.6100 1.3500 ;
      RECT 2.4760 0.2565 2.5020 1.3500 ;
      RECT 2.3680 0.2565 2.3940 1.3500 ;
      RECT 2.2600 0.2565 2.2860 1.3500 ;
      RECT 2.1520 0.2565 2.1780 1.3500 ;
      RECT 2.0440 0.2565 2.0700 1.3500 ;
      RECT 1.9360 0.2565 1.9620 1.3500 ;
      RECT 1.8280 0.2565 1.8540 1.3500 ;
      RECT 1.7200 0.2565 1.7460 1.3500 ;
      RECT 1.6120 0.2565 1.6380 1.3500 ;
      RECT 1.5040 0.2565 1.5300 1.3500 ;
      RECT 1.3960 0.2565 1.4220 1.3500 ;
      RECT 1.2880 0.2565 1.3140 1.3500 ;
      RECT 1.1800 0.2565 1.2060 1.3500 ;
      RECT 1.0720 0.2565 1.0980 1.3500 ;
      RECT 0.9640 0.2565 0.9900 1.3500 ;
      RECT 0.8560 0.2565 0.8820 1.3500 ;
      RECT 0.7480 0.2565 0.7740 1.3500 ;
      RECT 0.6400 0.2565 0.6660 1.3500 ;
      RECT 0.5320 0.2565 0.5580 1.3500 ;
      RECT 0.4240 0.2565 0.4500 1.3500 ;
      RECT 0.3160 0.2565 0.3420 1.3500 ;
      RECT 0.2080 0.2565 0.2340 1.3500 ;
      RECT 0.0050 0.2565 0.0900 1.3500 ;
      RECT 8.6410 1.3365 8.7690 2.4300 ;
      RECT 8.6270 2.0020 8.7690 2.3245 ;
      RECT 8.4790 1.7290 8.5410 2.4300 ;
      RECT 8.4650 2.0385 8.5410 2.1920 ;
      RECT 8.4790 1.3365 8.5050 2.4300 ;
      RECT 8.4790 1.4575 8.5190 1.6970 ;
      RECT 8.4790 1.3365 8.5410 1.4255 ;
      RECT 8.1820 1.7870 8.3880 2.4300 ;
      RECT 8.3620 1.3365 8.3880 2.4300 ;
      RECT 8.1820 2.0640 8.4020 2.3220 ;
      RECT 8.1820 1.3365 8.2800 2.4300 ;
      RECT 7.7650 1.3365 7.8480 2.4300 ;
      RECT 7.7650 1.4250 7.8620 2.3605 ;
      RECT 16.4440 1.3365 16.5290 2.4300 ;
      RECT 16.3000 1.3365 16.3260 2.4300 ;
      RECT 16.1920 1.3365 16.2180 2.4300 ;
      RECT 16.0840 1.3365 16.1100 2.4300 ;
      RECT 15.9760 1.3365 16.0020 2.4300 ;
      RECT 15.8680 1.3365 15.8940 2.4300 ;
      RECT 15.7600 1.3365 15.7860 2.4300 ;
      RECT 15.6520 1.3365 15.6780 2.4300 ;
      RECT 15.5440 1.3365 15.5700 2.4300 ;
      RECT 15.4360 1.3365 15.4620 2.4300 ;
      RECT 15.3280 1.3365 15.3540 2.4300 ;
      RECT 15.2200 1.3365 15.2460 2.4300 ;
      RECT 15.1120 1.3365 15.1380 2.4300 ;
      RECT 15.0040 1.3365 15.0300 2.4300 ;
      RECT 14.8960 1.3365 14.9220 2.4300 ;
      RECT 14.7880 1.3365 14.8140 2.4300 ;
      RECT 14.6800 1.3365 14.7060 2.4300 ;
      RECT 14.5720 1.3365 14.5980 2.4300 ;
      RECT 14.4640 1.3365 14.4900 2.4300 ;
      RECT 14.3560 1.3365 14.3820 2.4300 ;
      RECT 14.2480 1.3365 14.2740 2.4300 ;
      RECT 14.1400 1.3365 14.1660 2.4300 ;
      RECT 14.0320 1.3365 14.0580 2.4300 ;
      RECT 13.9240 1.3365 13.9500 2.4300 ;
      RECT 13.8160 1.3365 13.8420 2.4300 ;
      RECT 13.7080 1.3365 13.7340 2.4300 ;
      RECT 13.6000 1.3365 13.6260 2.4300 ;
      RECT 13.4920 1.3365 13.5180 2.4300 ;
      RECT 13.3840 1.3365 13.4100 2.4300 ;
      RECT 13.2760 1.3365 13.3020 2.4300 ;
      RECT 13.1680 1.3365 13.1940 2.4300 ;
      RECT 13.0600 1.3365 13.0860 2.4300 ;
      RECT 12.9520 1.3365 12.9780 2.4300 ;
      RECT 12.8440 1.3365 12.8700 2.4300 ;
      RECT 12.7360 1.3365 12.7620 2.4300 ;
      RECT 12.6280 1.3365 12.6540 2.4300 ;
      RECT 12.5200 1.3365 12.5460 2.4300 ;
      RECT 12.4120 1.3365 12.4380 2.4300 ;
      RECT 12.3040 1.3365 12.3300 2.4300 ;
      RECT 12.1960 1.3365 12.2220 2.4300 ;
      RECT 12.0880 1.3365 12.1140 2.4300 ;
      RECT 11.9800 1.3365 12.0060 2.4300 ;
      RECT 11.8720 1.3365 11.8980 2.4300 ;
      RECT 11.7640 1.3365 11.7900 2.4300 ;
      RECT 11.6560 1.3365 11.6820 2.4300 ;
      RECT 11.5480 1.3365 11.5740 2.4300 ;
      RECT 11.4400 1.3365 11.4660 2.4300 ;
      RECT 11.3320 1.3365 11.3580 2.4300 ;
      RECT 11.2240 1.3365 11.2500 2.4300 ;
      RECT 11.1160 1.3365 11.1420 2.4300 ;
      RECT 11.0080 1.3365 11.0340 2.4300 ;
      RECT 10.9000 1.3365 10.9260 2.4300 ;
      RECT 10.7920 1.3365 10.8180 2.4300 ;
      RECT 10.6840 1.3365 10.7100 2.4300 ;
      RECT 10.5760 1.3365 10.6020 2.4300 ;
      RECT 10.4680 1.3365 10.4940 2.4300 ;
      RECT 10.3600 1.3365 10.3860 2.4300 ;
      RECT 10.2520 1.3365 10.2780 2.4300 ;
      RECT 10.1440 1.3365 10.1700 2.4300 ;
      RECT 10.0360 1.3365 10.0620 2.4300 ;
      RECT 9.9280 1.3365 9.9540 2.4300 ;
      RECT 9.8200 1.3365 9.8460 2.4300 ;
      RECT 9.7120 1.3365 9.7380 2.4300 ;
      RECT 9.6040 1.3365 9.6300 2.4300 ;
      RECT 9.4960 1.3365 9.5220 2.4300 ;
      RECT 9.3880 1.3365 9.4140 2.4300 ;
      RECT 9.1750 1.3365 9.2520 2.4300 ;
      RECT 7.2820 1.3365 7.3590 2.4300 ;
      RECT 7.1200 1.3365 7.1460 2.4300 ;
      RECT 7.0120 1.3365 7.0380 2.4300 ;
      RECT 6.9040 1.3365 6.9300 2.4300 ;
      RECT 6.7960 1.3365 6.8220 2.4300 ;
      RECT 6.6880 1.3365 6.7140 2.4300 ;
      RECT 6.5800 1.3365 6.6060 2.4300 ;
      RECT 6.4720 1.3365 6.4980 2.4300 ;
      RECT 6.3640 1.3365 6.3900 2.4300 ;
      RECT 6.2560 1.3365 6.2820 2.4300 ;
      RECT 6.1480 1.3365 6.1740 2.4300 ;
      RECT 6.0400 1.3365 6.0660 2.4300 ;
      RECT 5.9320 1.3365 5.9580 2.4300 ;
      RECT 5.8240 1.3365 5.8500 2.4300 ;
      RECT 5.7160 1.3365 5.7420 2.4300 ;
      RECT 5.6080 1.3365 5.6340 2.4300 ;
      RECT 5.5000 1.3365 5.5260 2.4300 ;
      RECT 5.3920 1.3365 5.4180 2.4300 ;
      RECT 5.2840 1.3365 5.3100 2.4300 ;
      RECT 5.1760 1.3365 5.2020 2.4300 ;
      RECT 5.0680 1.3365 5.0940 2.4300 ;
      RECT 4.9600 1.3365 4.9860 2.4300 ;
      RECT 4.8520 1.3365 4.8780 2.4300 ;
      RECT 4.7440 1.3365 4.7700 2.4300 ;
      RECT 4.6360 1.3365 4.6620 2.4300 ;
      RECT 4.5280 1.3365 4.5540 2.4300 ;
      RECT 4.4200 1.3365 4.4460 2.4300 ;
      RECT 4.3120 1.3365 4.3380 2.4300 ;
      RECT 4.2040 1.3365 4.2300 2.4300 ;
      RECT 4.0960 1.3365 4.1220 2.4300 ;
      RECT 3.9880 1.3365 4.0140 2.4300 ;
      RECT 3.8800 1.3365 3.9060 2.4300 ;
      RECT 3.7720 1.3365 3.7980 2.4300 ;
      RECT 3.6640 1.3365 3.6900 2.4300 ;
      RECT 3.5560 1.3365 3.5820 2.4300 ;
      RECT 3.4480 1.3365 3.4740 2.4300 ;
      RECT 3.3400 1.3365 3.3660 2.4300 ;
      RECT 3.2320 1.3365 3.2580 2.4300 ;
      RECT 3.1240 1.3365 3.1500 2.4300 ;
      RECT 3.0160 1.3365 3.0420 2.4300 ;
      RECT 2.9080 1.3365 2.9340 2.4300 ;
      RECT 2.8000 1.3365 2.8260 2.4300 ;
      RECT 2.6920 1.3365 2.7180 2.4300 ;
      RECT 2.5840 1.3365 2.6100 2.4300 ;
      RECT 2.4760 1.3365 2.5020 2.4300 ;
      RECT 2.3680 1.3365 2.3940 2.4300 ;
      RECT 2.2600 1.3365 2.2860 2.4300 ;
      RECT 2.1520 1.3365 2.1780 2.4300 ;
      RECT 2.0440 1.3365 2.0700 2.4300 ;
      RECT 1.9360 1.3365 1.9620 2.4300 ;
      RECT 1.8280 1.3365 1.8540 2.4300 ;
      RECT 1.7200 1.3365 1.7460 2.4300 ;
      RECT 1.6120 1.3365 1.6380 2.4300 ;
      RECT 1.5040 1.3365 1.5300 2.4300 ;
      RECT 1.3960 1.3365 1.4220 2.4300 ;
      RECT 1.2880 1.3365 1.3140 2.4300 ;
      RECT 1.1800 1.3365 1.2060 2.4300 ;
      RECT 1.0720 1.3365 1.0980 2.4300 ;
      RECT 0.9640 1.3365 0.9900 2.4300 ;
      RECT 0.8560 1.3365 0.8820 2.4300 ;
      RECT 0.7480 1.3365 0.7740 2.4300 ;
      RECT 0.6400 1.3365 0.6660 2.4300 ;
      RECT 0.5320 1.3365 0.5580 2.4300 ;
      RECT 0.4240 1.3365 0.4500 2.4300 ;
      RECT 0.3160 1.3365 0.3420 2.4300 ;
      RECT 0.2080 1.3365 0.2340 2.4300 ;
      RECT 0.0050 1.3365 0.0900 2.4300 ;
      RECT 8.6410 2.4165 8.7690 3.5100 ;
      RECT 8.6270 3.0820 8.7690 3.4045 ;
      RECT 8.4790 2.8090 8.5410 3.5100 ;
      RECT 8.4650 3.1185 8.5410 3.2720 ;
      RECT 8.4790 2.4165 8.5050 3.5100 ;
      RECT 8.4790 2.5375 8.5190 2.7770 ;
      RECT 8.4790 2.4165 8.5410 2.5055 ;
      RECT 8.1820 2.8670 8.3880 3.5100 ;
      RECT 8.3620 2.4165 8.3880 3.5100 ;
      RECT 8.1820 3.1440 8.4020 3.4020 ;
      RECT 8.1820 2.4165 8.2800 3.5100 ;
      RECT 7.7650 2.4165 7.8480 3.5100 ;
      RECT 7.7650 2.5050 7.8620 3.4405 ;
      RECT 16.4440 2.4165 16.5290 3.5100 ;
      RECT 16.3000 2.4165 16.3260 3.5100 ;
      RECT 16.1920 2.4165 16.2180 3.5100 ;
      RECT 16.0840 2.4165 16.1100 3.5100 ;
      RECT 15.9760 2.4165 16.0020 3.5100 ;
      RECT 15.8680 2.4165 15.8940 3.5100 ;
      RECT 15.7600 2.4165 15.7860 3.5100 ;
      RECT 15.6520 2.4165 15.6780 3.5100 ;
      RECT 15.5440 2.4165 15.5700 3.5100 ;
      RECT 15.4360 2.4165 15.4620 3.5100 ;
      RECT 15.3280 2.4165 15.3540 3.5100 ;
      RECT 15.2200 2.4165 15.2460 3.5100 ;
      RECT 15.1120 2.4165 15.1380 3.5100 ;
      RECT 15.0040 2.4165 15.0300 3.5100 ;
      RECT 14.8960 2.4165 14.9220 3.5100 ;
      RECT 14.7880 2.4165 14.8140 3.5100 ;
      RECT 14.6800 2.4165 14.7060 3.5100 ;
      RECT 14.5720 2.4165 14.5980 3.5100 ;
      RECT 14.4640 2.4165 14.4900 3.5100 ;
      RECT 14.3560 2.4165 14.3820 3.5100 ;
      RECT 14.2480 2.4165 14.2740 3.5100 ;
      RECT 14.1400 2.4165 14.1660 3.5100 ;
      RECT 14.0320 2.4165 14.0580 3.5100 ;
      RECT 13.9240 2.4165 13.9500 3.5100 ;
      RECT 13.8160 2.4165 13.8420 3.5100 ;
      RECT 13.7080 2.4165 13.7340 3.5100 ;
      RECT 13.6000 2.4165 13.6260 3.5100 ;
      RECT 13.4920 2.4165 13.5180 3.5100 ;
      RECT 13.3840 2.4165 13.4100 3.5100 ;
      RECT 13.2760 2.4165 13.3020 3.5100 ;
      RECT 13.1680 2.4165 13.1940 3.5100 ;
      RECT 13.0600 2.4165 13.0860 3.5100 ;
      RECT 12.9520 2.4165 12.9780 3.5100 ;
      RECT 12.8440 2.4165 12.8700 3.5100 ;
      RECT 12.7360 2.4165 12.7620 3.5100 ;
      RECT 12.6280 2.4165 12.6540 3.5100 ;
      RECT 12.5200 2.4165 12.5460 3.5100 ;
      RECT 12.4120 2.4165 12.4380 3.5100 ;
      RECT 12.3040 2.4165 12.3300 3.5100 ;
      RECT 12.1960 2.4165 12.2220 3.5100 ;
      RECT 12.0880 2.4165 12.1140 3.5100 ;
      RECT 11.9800 2.4165 12.0060 3.5100 ;
      RECT 11.8720 2.4165 11.8980 3.5100 ;
      RECT 11.7640 2.4165 11.7900 3.5100 ;
      RECT 11.6560 2.4165 11.6820 3.5100 ;
      RECT 11.5480 2.4165 11.5740 3.5100 ;
      RECT 11.4400 2.4165 11.4660 3.5100 ;
      RECT 11.3320 2.4165 11.3580 3.5100 ;
      RECT 11.2240 2.4165 11.2500 3.5100 ;
      RECT 11.1160 2.4165 11.1420 3.5100 ;
      RECT 11.0080 2.4165 11.0340 3.5100 ;
      RECT 10.9000 2.4165 10.9260 3.5100 ;
      RECT 10.7920 2.4165 10.8180 3.5100 ;
      RECT 10.6840 2.4165 10.7100 3.5100 ;
      RECT 10.5760 2.4165 10.6020 3.5100 ;
      RECT 10.4680 2.4165 10.4940 3.5100 ;
      RECT 10.3600 2.4165 10.3860 3.5100 ;
      RECT 10.2520 2.4165 10.2780 3.5100 ;
      RECT 10.1440 2.4165 10.1700 3.5100 ;
      RECT 10.0360 2.4165 10.0620 3.5100 ;
      RECT 9.9280 2.4165 9.9540 3.5100 ;
      RECT 9.8200 2.4165 9.8460 3.5100 ;
      RECT 9.7120 2.4165 9.7380 3.5100 ;
      RECT 9.6040 2.4165 9.6300 3.5100 ;
      RECT 9.4960 2.4165 9.5220 3.5100 ;
      RECT 9.3880 2.4165 9.4140 3.5100 ;
      RECT 9.1750 2.4165 9.2520 3.5100 ;
      RECT 7.2820 2.4165 7.3590 3.5100 ;
      RECT 7.1200 2.4165 7.1460 3.5100 ;
      RECT 7.0120 2.4165 7.0380 3.5100 ;
      RECT 6.9040 2.4165 6.9300 3.5100 ;
      RECT 6.7960 2.4165 6.8220 3.5100 ;
      RECT 6.6880 2.4165 6.7140 3.5100 ;
      RECT 6.5800 2.4165 6.6060 3.5100 ;
      RECT 6.4720 2.4165 6.4980 3.5100 ;
      RECT 6.3640 2.4165 6.3900 3.5100 ;
      RECT 6.2560 2.4165 6.2820 3.5100 ;
      RECT 6.1480 2.4165 6.1740 3.5100 ;
      RECT 6.0400 2.4165 6.0660 3.5100 ;
      RECT 5.9320 2.4165 5.9580 3.5100 ;
      RECT 5.8240 2.4165 5.8500 3.5100 ;
      RECT 5.7160 2.4165 5.7420 3.5100 ;
      RECT 5.6080 2.4165 5.6340 3.5100 ;
      RECT 5.5000 2.4165 5.5260 3.5100 ;
      RECT 5.3920 2.4165 5.4180 3.5100 ;
      RECT 5.2840 2.4165 5.3100 3.5100 ;
      RECT 5.1760 2.4165 5.2020 3.5100 ;
      RECT 5.0680 2.4165 5.0940 3.5100 ;
      RECT 4.9600 2.4165 4.9860 3.5100 ;
      RECT 4.8520 2.4165 4.8780 3.5100 ;
      RECT 4.7440 2.4165 4.7700 3.5100 ;
      RECT 4.6360 2.4165 4.6620 3.5100 ;
      RECT 4.5280 2.4165 4.5540 3.5100 ;
      RECT 4.4200 2.4165 4.4460 3.5100 ;
      RECT 4.3120 2.4165 4.3380 3.5100 ;
      RECT 4.2040 2.4165 4.2300 3.5100 ;
      RECT 4.0960 2.4165 4.1220 3.5100 ;
      RECT 3.9880 2.4165 4.0140 3.5100 ;
      RECT 3.8800 2.4165 3.9060 3.5100 ;
      RECT 3.7720 2.4165 3.7980 3.5100 ;
      RECT 3.6640 2.4165 3.6900 3.5100 ;
      RECT 3.5560 2.4165 3.5820 3.5100 ;
      RECT 3.4480 2.4165 3.4740 3.5100 ;
      RECT 3.3400 2.4165 3.3660 3.5100 ;
      RECT 3.2320 2.4165 3.2580 3.5100 ;
      RECT 3.1240 2.4165 3.1500 3.5100 ;
      RECT 3.0160 2.4165 3.0420 3.5100 ;
      RECT 2.9080 2.4165 2.9340 3.5100 ;
      RECT 2.8000 2.4165 2.8260 3.5100 ;
      RECT 2.6920 2.4165 2.7180 3.5100 ;
      RECT 2.5840 2.4165 2.6100 3.5100 ;
      RECT 2.4760 2.4165 2.5020 3.5100 ;
      RECT 2.3680 2.4165 2.3940 3.5100 ;
      RECT 2.2600 2.4165 2.2860 3.5100 ;
      RECT 2.1520 2.4165 2.1780 3.5100 ;
      RECT 2.0440 2.4165 2.0700 3.5100 ;
      RECT 1.9360 2.4165 1.9620 3.5100 ;
      RECT 1.8280 2.4165 1.8540 3.5100 ;
      RECT 1.7200 2.4165 1.7460 3.5100 ;
      RECT 1.6120 2.4165 1.6380 3.5100 ;
      RECT 1.5040 2.4165 1.5300 3.5100 ;
      RECT 1.3960 2.4165 1.4220 3.5100 ;
      RECT 1.2880 2.4165 1.3140 3.5100 ;
      RECT 1.1800 2.4165 1.2060 3.5100 ;
      RECT 1.0720 2.4165 1.0980 3.5100 ;
      RECT 0.9640 2.4165 0.9900 3.5100 ;
      RECT 0.8560 2.4165 0.8820 3.5100 ;
      RECT 0.7480 2.4165 0.7740 3.5100 ;
      RECT 0.6400 2.4165 0.6660 3.5100 ;
      RECT 0.5320 2.4165 0.5580 3.5100 ;
      RECT 0.4240 2.4165 0.4500 3.5100 ;
      RECT 0.3160 2.4165 0.3420 3.5100 ;
      RECT 0.2080 2.4165 0.2340 3.5100 ;
      RECT 0.0050 2.4165 0.0900 3.5100 ;
      RECT 8.6410 3.4965 8.7690 4.5900 ;
      RECT 8.6270 4.1620 8.7690 4.4845 ;
      RECT 8.4790 3.8890 8.5410 4.5900 ;
      RECT 8.4650 4.1985 8.5410 4.3520 ;
      RECT 8.4790 3.4965 8.5050 4.5900 ;
      RECT 8.4790 3.6175 8.5190 3.8570 ;
      RECT 8.4790 3.4965 8.5410 3.5855 ;
      RECT 8.1820 3.9470 8.3880 4.5900 ;
      RECT 8.3620 3.4965 8.3880 4.5900 ;
      RECT 8.1820 4.2240 8.4020 4.4820 ;
      RECT 8.1820 3.4965 8.2800 4.5900 ;
      RECT 7.7650 3.4965 7.8480 4.5900 ;
      RECT 7.7650 3.5850 7.8620 4.5205 ;
      RECT 16.4440 3.4965 16.5290 4.5900 ;
      RECT 16.3000 3.4965 16.3260 4.5900 ;
      RECT 16.1920 3.4965 16.2180 4.5900 ;
      RECT 16.0840 3.4965 16.1100 4.5900 ;
      RECT 15.9760 3.4965 16.0020 4.5900 ;
      RECT 15.8680 3.4965 15.8940 4.5900 ;
      RECT 15.7600 3.4965 15.7860 4.5900 ;
      RECT 15.6520 3.4965 15.6780 4.5900 ;
      RECT 15.5440 3.4965 15.5700 4.5900 ;
      RECT 15.4360 3.4965 15.4620 4.5900 ;
      RECT 15.3280 3.4965 15.3540 4.5900 ;
      RECT 15.2200 3.4965 15.2460 4.5900 ;
      RECT 15.1120 3.4965 15.1380 4.5900 ;
      RECT 15.0040 3.4965 15.0300 4.5900 ;
      RECT 14.8960 3.4965 14.9220 4.5900 ;
      RECT 14.7880 3.4965 14.8140 4.5900 ;
      RECT 14.6800 3.4965 14.7060 4.5900 ;
      RECT 14.5720 3.4965 14.5980 4.5900 ;
      RECT 14.4640 3.4965 14.4900 4.5900 ;
      RECT 14.3560 3.4965 14.3820 4.5900 ;
      RECT 14.2480 3.4965 14.2740 4.5900 ;
      RECT 14.1400 3.4965 14.1660 4.5900 ;
      RECT 14.0320 3.4965 14.0580 4.5900 ;
      RECT 13.9240 3.4965 13.9500 4.5900 ;
      RECT 13.8160 3.4965 13.8420 4.5900 ;
      RECT 13.7080 3.4965 13.7340 4.5900 ;
      RECT 13.6000 3.4965 13.6260 4.5900 ;
      RECT 13.4920 3.4965 13.5180 4.5900 ;
      RECT 13.3840 3.4965 13.4100 4.5900 ;
      RECT 13.2760 3.4965 13.3020 4.5900 ;
      RECT 13.1680 3.4965 13.1940 4.5900 ;
      RECT 13.0600 3.4965 13.0860 4.5900 ;
      RECT 12.9520 3.4965 12.9780 4.5900 ;
      RECT 12.8440 3.4965 12.8700 4.5900 ;
      RECT 12.7360 3.4965 12.7620 4.5900 ;
      RECT 12.6280 3.4965 12.6540 4.5900 ;
      RECT 12.5200 3.4965 12.5460 4.5900 ;
      RECT 12.4120 3.4965 12.4380 4.5900 ;
      RECT 12.3040 3.4965 12.3300 4.5900 ;
      RECT 12.1960 3.4965 12.2220 4.5900 ;
      RECT 12.0880 3.4965 12.1140 4.5900 ;
      RECT 11.9800 3.4965 12.0060 4.5900 ;
      RECT 11.8720 3.4965 11.8980 4.5900 ;
      RECT 11.7640 3.4965 11.7900 4.5900 ;
      RECT 11.6560 3.4965 11.6820 4.5900 ;
      RECT 11.5480 3.4965 11.5740 4.5900 ;
      RECT 11.4400 3.4965 11.4660 4.5900 ;
      RECT 11.3320 3.4965 11.3580 4.5900 ;
      RECT 11.2240 3.4965 11.2500 4.5900 ;
      RECT 11.1160 3.4965 11.1420 4.5900 ;
      RECT 11.0080 3.4965 11.0340 4.5900 ;
      RECT 10.9000 3.4965 10.9260 4.5900 ;
      RECT 10.7920 3.4965 10.8180 4.5900 ;
      RECT 10.6840 3.4965 10.7100 4.5900 ;
      RECT 10.5760 3.4965 10.6020 4.5900 ;
      RECT 10.4680 3.4965 10.4940 4.5900 ;
      RECT 10.3600 3.4965 10.3860 4.5900 ;
      RECT 10.2520 3.4965 10.2780 4.5900 ;
      RECT 10.1440 3.4965 10.1700 4.5900 ;
      RECT 10.0360 3.4965 10.0620 4.5900 ;
      RECT 9.9280 3.4965 9.9540 4.5900 ;
      RECT 9.8200 3.4965 9.8460 4.5900 ;
      RECT 9.7120 3.4965 9.7380 4.5900 ;
      RECT 9.6040 3.4965 9.6300 4.5900 ;
      RECT 9.4960 3.4965 9.5220 4.5900 ;
      RECT 9.3880 3.4965 9.4140 4.5900 ;
      RECT 9.1750 3.4965 9.2520 4.5900 ;
      RECT 7.2820 3.4965 7.3590 4.5900 ;
      RECT 7.1200 3.4965 7.1460 4.5900 ;
      RECT 7.0120 3.4965 7.0380 4.5900 ;
      RECT 6.9040 3.4965 6.9300 4.5900 ;
      RECT 6.7960 3.4965 6.8220 4.5900 ;
      RECT 6.6880 3.4965 6.7140 4.5900 ;
      RECT 6.5800 3.4965 6.6060 4.5900 ;
      RECT 6.4720 3.4965 6.4980 4.5900 ;
      RECT 6.3640 3.4965 6.3900 4.5900 ;
      RECT 6.2560 3.4965 6.2820 4.5900 ;
      RECT 6.1480 3.4965 6.1740 4.5900 ;
      RECT 6.0400 3.4965 6.0660 4.5900 ;
      RECT 5.9320 3.4965 5.9580 4.5900 ;
      RECT 5.8240 3.4965 5.8500 4.5900 ;
      RECT 5.7160 3.4965 5.7420 4.5900 ;
      RECT 5.6080 3.4965 5.6340 4.5900 ;
      RECT 5.5000 3.4965 5.5260 4.5900 ;
      RECT 5.3920 3.4965 5.4180 4.5900 ;
      RECT 5.2840 3.4965 5.3100 4.5900 ;
      RECT 5.1760 3.4965 5.2020 4.5900 ;
      RECT 5.0680 3.4965 5.0940 4.5900 ;
      RECT 4.9600 3.4965 4.9860 4.5900 ;
      RECT 4.8520 3.4965 4.8780 4.5900 ;
      RECT 4.7440 3.4965 4.7700 4.5900 ;
      RECT 4.6360 3.4965 4.6620 4.5900 ;
      RECT 4.5280 3.4965 4.5540 4.5900 ;
      RECT 4.4200 3.4965 4.4460 4.5900 ;
      RECT 4.3120 3.4965 4.3380 4.5900 ;
      RECT 4.2040 3.4965 4.2300 4.5900 ;
      RECT 4.0960 3.4965 4.1220 4.5900 ;
      RECT 3.9880 3.4965 4.0140 4.5900 ;
      RECT 3.8800 3.4965 3.9060 4.5900 ;
      RECT 3.7720 3.4965 3.7980 4.5900 ;
      RECT 3.6640 3.4965 3.6900 4.5900 ;
      RECT 3.5560 3.4965 3.5820 4.5900 ;
      RECT 3.4480 3.4965 3.4740 4.5900 ;
      RECT 3.3400 3.4965 3.3660 4.5900 ;
      RECT 3.2320 3.4965 3.2580 4.5900 ;
      RECT 3.1240 3.4965 3.1500 4.5900 ;
      RECT 3.0160 3.4965 3.0420 4.5900 ;
      RECT 2.9080 3.4965 2.9340 4.5900 ;
      RECT 2.8000 3.4965 2.8260 4.5900 ;
      RECT 2.6920 3.4965 2.7180 4.5900 ;
      RECT 2.5840 3.4965 2.6100 4.5900 ;
      RECT 2.4760 3.4965 2.5020 4.5900 ;
      RECT 2.3680 3.4965 2.3940 4.5900 ;
      RECT 2.2600 3.4965 2.2860 4.5900 ;
      RECT 2.1520 3.4965 2.1780 4.5900 ;
      RECT 2.0440 3.4965 2.0700 4.5900 ;
      RECT 1.9360 3.4965 1.9620 4.5900 ;
      RECT 1.8280 3.4965 1.8540 4.5900 ;
      RECT 1.7200 3.4965 1.7460 4.5900 ;
      RECT 1.6120 3.4965 1.6380 4.5900 ;
      RECT 1.5040 3.4965 1.5300 4.5900 ;
      RECT 1.3960 3.4965 1.4220 4.5900 ;
      RECT 1.2880 3.4965 1.3140 4.5900 ;
      RECT 1.1800 3.4965 1.2060 4.5900 ;
      RECT 1.0720 3.4965 1.0980 4.5900 ;
      RECT 0.9640 3.4965 0.9900 4.5900 ;
      RECT 0.8560 3.4965 0.8820 4.5900 ;
      RECT 0.7480 3.4965 0.7740 4.5900 ;
      RECT 0.6400 3.4965 0.6660 4.5900 ;
      RECT 0.5320 3.4965 0.5580 4.5900 ;
      RECT 0.4240 3.4965 0.4500 4.5900 ;
      RECT 0.3160 3.4965 0.3420 4.5900 ;
      RECT 0.2080 3.4965 0.2340 4.5900 ;
      RECT 0.0050 3.4965 0.0900 4.5900 ;
      RECT 8.6410 4.5765 8.7690 5.6700 ;
      RECT 8.6270 5.2420 8.7690 5.5645 ;
      RECT 8.4790 4.9690 8.5410 5.6700 ;
      RECT 8.4650 5.2785 8.5410 5.4320 ;
      RECT 8.4790 4.5765 8.5050 5.6700 ;
      RECT 8.4790 4.6975 8.5190 4.9370 ;
      RECT 8.4790 4.5765 8.5410 4.6655 ;
      RECT 8.1820 5.0270 8.3880 5.6700 ;
      RECT 8.3620 4.5765 8.3880 5.6700 ;
      RECT 8.1820 5.3040 8.4020 5.5620 ;
      RECT 8.1820 4.5765 8.2800 5.6700 ;
      RECT 7.7650 4.5765 7.8480 5.6700 ;
      RECT 7.7650 4.6650 7.8620 5.6005 ;
      RECT 16.4440 4.5765 16.5290 5.6700 ;
      RECT 16.3000 4.5765 16.3260 5.6700 ;
      RECT 16.1920 4.5765 16.2180 5.6700 ;
      RECT 16.0840 4.5765 16.1100 5.6700 ;
      RECT 15.9760 4.5765 16.0020 5.6700 ;
      RECT 15.8680 4.5765 15.8940 5.6700 ;
      RECT 15.7600 4.5765 15.7860 5.6700 ;
      RECT 15.6520 4.5765 15.6780 5.6700 ;
      RECT 15.5440 4.5765 15.5700 5.6700 ;
      RECT 15.4360 4.5765 15.4620 5.6700 ;
      RECT 15.3280 4.5765 15.3540 5.6700 ;
      RECT 15.2200 4.5765 15.2460 5.6700 ;
      RECT 15.1120 4.5765 15.1380 5.6700 ;
      RECT 15.0040 4.5765 15.0300 5.6700 ;
      RECT 14.8960 4.5765 14.9220 5.6700 ;
      RECT 14.7880 4.5765 14.8140 5.6700 ;
      RECT 14.6800 4.5765 14.7060 5.6700 ;
      RECT 14.5720 4.5765 14.5980 5.6700 ;
      RECT 14.4640 4.5765 14.4900 5.6700 ;
      RECT 14.3560 4.5765 14.3820 5.6700 ;
      RECT 14.2480 4.5765 14.2740 5.6700 ;
      RECT 14.1400 4.5765 14.1660 5.6700 ;
      RECT 14.0320 4.5765 14.0580 5.6700 ;
      RECT 13.9240 4.5765 13.9500 5.6700 ;
      RECT 13.8160 4.5765 13.8420 5.6700 ;
      RECT 13.7080 4.5765 13.7340 5.6700 ;
      RECT 13.6000 4.5765 13.6260 5.6700 ;
      RECT 13.4920 4.5765 13.5180 5.6700 ;
      RECT 13.3840 4.5765 13.4100 5.6700 ;
      RECT 13.2760 4.5765 13.3020 5.6700 ;
      RECT 13.1680 4.5765 13.1940 5.6700 ;
      RECT 13.0600 4.5765 13.0860 5.6700 ;
      RECT 12.9520 4.5765 12.9780 5.6700 ;
      RECT 12.8440 4.5765 12.8700 5.6700 ;
      RECT 12.7360 4.5765 12.7620 5.6700 ;
      RECT 12.6280 4.5765 12.6540 5.6700 ;
      RECT 12.5200 4.5765 12.5460 5.6700 ;
      RECT 12.4120 4.5765 12.4380 5.6700 ;
      RECT 12.3040 4.5765 12.3300 5.6700 ;
      RECT 12.1960 4.5765 12.2220 5.6700 ;
      RECT 12.0880 4.5765 12.1140 5.6700 ;
      RECT 11.9800 4.5765 12.0060 5.6700 ;
      RECT 11.8720 4.5765 11.8980 5.6700 ;
      RECT 11.7640 4.5765 11.7900 5.6700 ;
      RECT 11.6560 4.5765 11.6820 5.6700 ;
      RECT 11.5480 4.5765 11.5740 5.6700 ;
      RECT 11.4400 4.5765 11.4660 5.6700 ;
      RECT 11.3320 4.5765 11.3580 5.6700 ;
      RECT 11.2240 4.5765 11.2500 5.6700 ;
      RECT 11.1160 4.5765 11.1420 5.6700 ;
      RECT 11.0080 4.5765 11.0340 5.6700 ;
      RECT 10.9000 4.5765 10.9260 5.6700 ;
      RECT 10.7920 4.5765 10.8180 5.6700 ;
      RECT 10.6840 4.5765 10.7100 5.6700 ;
      RECT 10.5760 4.5765 10.6020 5.6700 ;
      RECT 10.4680 4.5765 10.4940 5.6700 ;
      RECT 10.3600 4.5765 10.3860 5.6700 ;
      RECT 10.2520 4.5765 10.2780 5.6700 ;
      RECT 10.1440 4.5765 10.1700 5.6700 ;
      RECT 10.0360 4.5765 10.0620 5.6700 ;
      RECT 9.9280 4.5765 9.9540 5.6700 ;
      RECT 9.8200 4.5765 9.8460 5.6700 ;
      RECT 9.7120 4.5765 9.7380 5.6700 ;
      RECT 9.6040 4.5765 9.6300 5.6700 ;
      RECT 9.4960 4.5765 9.5220 5.6700 ;
      RECT 9.3880 4.5765 9.4140 5.6700 ;
      RECT 9.1750 4.5765 9.2520 5.6700 ;
      RECT 7.2820 4.5765 7.3590 5.6700 ;
      RECT 7.1200 4.5765 7.1460 5.6700 ;
      RECT 7.0120 4.5765 7.0380 5.6700 ;
      RECT 6.9040 4.5765 6.9300 5.6700 ;
      RECT 6.7960 4.5765 6.8220 5.6700 ;
      RECT 6.6880 4.5765 6.7140 5.6700 ;
      RECT 6.5800 4.5765 6.6060 5.6700 ;
      RECT 6.4720 4.5765 6.4980 5.6700 ;
      RECT 6.3640 4.5765 6.3900 5.6700 ;
      RECT 6.2560 4.5765 6.2820 5.6700 ;
      RECT 6.1480 4.5765 6.1740 5.6700 ;
      RECT 6.0400 4.5765 6.0660 5.6700 ;
      RECT 5.9320 4.5765 5.9580 5.6700 ;
      RECT 5.8240 4.5765 5.8500 5.6700 ;
      RECT 5.7160 4.5765 5.7420 5.6700 ;
      RECT 5.6080 4.5765 5.6340 5.6700 ;
      RECT 5.5000 4.5765 5.5260 5.6700 ;
      RECT 5.3920 4.5765 5.4180 5.6700 ;
      RECT 5.2840 4.5765 5.3100 5.6700 ;
      RECT 5.1760 4.5765 5.2020 5.6700 ;
      RECT 5.0680 4.5765 5.0940 5.6700 ;
      RECT 4.9600 4.5765 4.9860 5.6700 ;
      RECT 4.8520 4.5765 4.8780 5.6700 ;
      RECT 4.7440 4.5765 4.7700 5.6700 ;
      RECT 4.6360 4.5765 4.6620 5.6700 ;
      RECT 4.5280 4.5765 4.5540 5.6700 ;
      RECT 4.4200 4.5765 4.4460 5.6700 ;
      RECT 4.3120 4.5765 4.3380 5.6700 ;
      RECT 4.2040 4.5765 4.2300 5.6700 ;
      RECT 4.0960 4.5765 4.1220 5.6700 ;
      RECT 3.9880 4.5765 4.0140 5.6700 ;
      RECT 3.8800 4.5765 3.9060 5.6700 ;
      RECT 3.7720 4.5765 3.7980 5.6700 ;
      RECT 3.6640 4.5765 3.6900 5.6700 ;
      RECT 3.5560 4.5765 3.5820 5.6700 ;
      RECT 3.4480 4.5765 3.4740 5.6700 ;
      RECT 3.3400 4.5765 3.3660 5.6700 ;
      RECT 3.2320 4.5765 3.2580 5.6700 ;
      RECT 3.1240 4.5765 3.1500 5.6700 ;
      RECT 3.0160 4.5765 3.0420 5.6700 ;
      RECT 2.9080 4.5765 2.9340 5.6700 ;
      RECT 2.8000 4.5765 2.8260 5.6700 ;
      RECT 2.6920 4.5765 2.7180 5.6700 ;
      RECT 2.5840 4.5765 2.6100 5.6700 ;
      RECT 2.4760 4.5765 2.5020 5.6700 ;
      RECT 2.3680 4.5765 2.3940 5.6700 ;
      RECT 2.2600 4.5765 2.2860 5.6700 ;
      RECT 2.1520 4.5765 2.1780 5.6700 ;
      RECT 2.0440 4.5765 2.0700 5.6700 ;
      RECT 1.9360 4.5765 1.9620 5.6700 ;
      RECT 1.8280 4.5765 1.8540 5.6700 ;
      RECT 1.7200 4.5765 1.7460 5.6700 ;
      RECT 1.6120 4.5765 1.6380 5.6700 ;
      RECT 1.5040 4.5765 1.5300 5.6700 ;
      RECT 1.3960 4.5765 1.4220 5.6700 ;
      RECT 1.2880 4.5765 1.3140 5.6700 ;
      RECT 1.1800 4.5765 1.2060 5.6700 ;
      RECT 1.0720 4.5765 1.0980 5.6700 ;
      RECT 0.9640 4.5765 0.9900 5.6700 ;
      RECT 0.8560 4.5765 0.8820 5.6700 ;
      RECT 0.7480 4.5765 0.7740 5.6700 ;
      RECT 0.6400 4.5765 0.6660 5.6700 ;
      RECT 0.5320 4.5765 0.5580 5.6700 ;
      RECT 0.4240 4.5765 0.4500 5.6700 ;
      RECT 0.3160 4.5765 0.3420 5.6700 ;
      RECT 0.2080 4.5765 0.2340 5.6700 ;
      RECT 0.0050 4.5765 0.0900 5.6700 ;
      RECT 8.6410 5.6565 8.7690 6.7500 ;
      RECT 8.6270 6.3220 8.7690 6.6445 ;
      RECT 8.4790 6.0490 8.5410 6.7500 ;
      RECT 8.4650 6.3585 8.5410 6.5120 ;
      RECT 8.4790 5.6565 8.5050 6.7500 ;
      RECT 8.4790 5.7775 8.5190 6.0170 ;
      RECT 8.4790 5.6565 8.5410 5.7455 ;
      RECT 8.1820 6.1070 8.3880 6.7500 ;
      RECT 8.3620 5.6565 8.3880 6.7500 ;
      RECT 8.1820 6.3840 8.4020 6.6420 ;
      RECT 8.1820 5.6565 8.2800 6.7500 ;
      RECT 7.7650 5.6565 7.8480 6.7500 ;
      RECT 7.7650 5.7450 7.8620 6.6805 ;
      RECT 16.4440 5.6565 16.5290 6.7500 ;
      RECT 16.3000 5.6565 16.3260 6.7500 ;
      RECT 16.1920 5.6565 16.2180 6.7500 ;
      RECT 16.0840 5.6565 16.1100 6.7500 ;
      RECT 15.9760 5.6565 16.0020 6.7500 ;
      RECT 15.8680 5.6565 15.8940 6.7500 ;
      RECT 15.7600 5.6565 15.7860 6.7500 ;
      RECT 15.6520 5.6565 15.6780 6.7500 ;
      RECT 15.5440 5.6565 15.5700 6.7500 ;
      RECT 15.4360 5.6565 15.4620 6.7500 ;
      RECT 15.3280 5.6565 15.3540 6.7500 ;
      RECT 15.2200 5.6565 15.2460 6.7500 ;
      RECT 15.1120 5.6565 15.1380 6.7500 ;
      RECT 15.0040 5.6565 15.0300 6.7500 ;
      RECT 14.8960 5.6565 14.9220 6.7500 ;
      RECT 14.7880 5.6565 14.8140 6.7500 ;
      RECT 14.6800 5.6565 14.7060 6.7500 ;
      RECT 14.5720 5.6565 14.5980 6.7500 ;
      RECT 14.4640 5.6565 14.4900 6.7500 ;
      RECT 14.3560 5.6565 14.3820 6.7500 ;
      RECT 14.2480 5.6565 14.2740 6.7500 ;
      RECT 14.1400 5.6565 14.1660 6.7500 ;
      RECT 14.0320 5.6565 14.0580 6.7500 ;
      RECT 13.9240 5.6565 13.9500 6.7500 ;
      RECT 13.8160 5.6565 13.8420 6.7500 ;
      RECT 13.7080 5.6565 13.7340 6.7500 ;
      RECT 13.6000 5.6565 13.6260 6.7500 ;
      RECT 13.4920 5.6565 13.5180 6.7500 ;
      RECT 13.3840 5.6565 13.4100 6.7500 ;
      RECT 13.2760 5.6565 13.3020 6.7500 ;
      RECT 13.1680 5.6565 13.1940 6.7500 ;
      RECT 13.0600 5.6565 13.0860 6.7500 ;
      RECT 12.9520 5.6565 12.9780 6.7500 ;
      RECT 12.8440 5.6565 12.8700 6.7500 ;
      RECT 12.7360 5.6565 12.7620 6.7500 ;
      RECT 12.6280 5.6565 12.6540 6.7500 ;
      RECT 12.5200 5.6565 12.5460 6.7500 ;
      RECT 12.4120 5.6565 12.4380 6.7500 ;
      RECT 12.3040 5.6565 12.3300 6.7500 ;
      RECT 12.1960 5.6565 12.2220 6.7500 ;
      RECT 12.0880 5.6565 12.1140 6.7500 ;
      RECT 11.9800 5.6565 12.0060 6.7500 ;
      RECT 11.8720 5.6565 11.8980 6.7500 ;
      RECT 11.7640 5.6565 11.7900 6.7500 ;
      RECT 11.6560 5.6565 11.6820 6.7500 ;
      RECT 11.5480 5.6565 11.5740 6.7500 ;
      RECT 11.4400 5.6565 11.4660 6.7500 ;
      RECT 11.3320 5.6565 11.3580 6.7500 ;
      RECT 11.2240 5.6565 11.2500 6.7500 ;
      RECT 11.1160 5.6565 11.1420 6.7500 ;
      RECT 11.0080 5.6565 11.0340 6.7500 ;
      RECT 10.9000 5.6565 10.9260 6.7500 ;
      RECT 10.7920 5.6565 10.8180 6.7500 ;
      RECT 10.6840 5.6565 10.7100 6.7500 ;
      RECT 10.5760 5.6565 10.6020 6.7500 ;
      RECT 10.4680 5.6565 10.4940 6.7500 ;
      RECT 10.3600 5.6565 10.3860 6.7500 ;
      RECT 10.2520 5.6565 10.2780 6.7500 ;
      RECT 10.1440 5.6565 10.1700 6.7500 ;
      RECT 10.0360 5.6565 10.0620 6.7500 ;
      RECT 9.9280 5.6565 9.9540 6.7500 ;
      RECT 9.8200 5.6565 9.8460 6.7500 ;
      RECT 9.7120 5.6565 9.7380 6.7500 ;
      RECT 9.6040 5.6565 9.6300 6.7500 ;
      RECT 9.4960 5.6565 9.5220 6.7500 ;
      RECT 9.3880 5.6565 9.4140 6.7500 ;
      RECT 9.1750 5.6565 9.2520 6.7500 ;
      RECT 7.2820 5.6565 7.3590 6.7500 ;
      RECT 7.1200 5.6565 7.1460 6.7500 ;
      RECT 7.0120 5.6565 7.0380 6.7500 ;
      RECT 6.9040 5.6565 6.9300 6.7500 ;
      RECT 6.7960 5.6565 6.8220 6.7500 ;
      RECT 6.6880 5.6565 6.7140 6.7500 ;
      RECT 6.5800 5.6565 6.6060 6.7500 ;
      RECT 6.4720 5.6565 6.4980 6.7500 ;
      RECT 6.3640 5.6565 6.3900 6.7500 ;
      RECT 6.2560 5.6565 6.2820 6.7500 ;
      RECT 6.1480 5.6565 6.1740 6.7500 ;
      RECT 6.0400 5.6565 6.0660 6.7500 ;
      RECT 5.9320 5.6565 5.9580 6.7500 ;
      RECT 5.8240 5.6565 5.8500 6.7500 ;
      RECT 5.7160 5.6565 5.7420 6.7500 ;
      RECT 5.6080 5.6565 5.6340 6.7500 ;
      RECT 5.5000 5.6565 5.5260 6.7500 ;
      RECT 5.3920 5.6565 5.4180 6.7500 ;
      RECT 5.2840 5.6565 5.3100 6.7500 ;
      RECT 5.1760 5.6565 5.2020 6.7500 ;
      RECT 5.0680 5.6565 5.0940 6.7500 ;
      RECT 4.9600 5.6565 4.9860 6.7500 ;
      RECT 4.8520 5.6565 4.8780 6.7500 ;
      RECT 4.7440 5.6565 4.7700 6.7500 ;
      RECT 4.6360 5.6565 4.6620 6.7500 ;
      RECT 4.5280 5.6565 4.5540 6.7500 ;
      RECT 4.4200 5.6565 4.4460 6.7500 ;
      RECT 4.3120 5.6565 4.3380 6.7500 ;
      RECT 4.2040 5.6565 4.2300 6.7500 ;
      RECT 4.0960 5.6565 4.1220 6.7500 ;
      RECT 3.9880 5.6565 4.0140 6.7500 ;
      RECT 3.8800 5.6565 3.9060 6.7500 ;
      RECT 3.7720 5.6565 3.7980 6.7500 ;
      RECT 3.6640 5.6565 3.6900 6.7500 ;
      RECT 3.5560 5.6565 3.5820 6.7500 ;
      RECT 3.4480 5.6565 3.4740 6.7500 ;
      RECT 3.3400 5.6565 3.3660 6.7500 ;
      RECT 3.2320 5.6565 3.2580 6.7500 ;
      RECT 3.1240 5.6565 3.1500 6.7500 ;
      RECT 3.0160 5.6565 3.0420 6.7500 ;
      RECT 2.9080 5.6565 2.9340 6.7500 ;
      RECT 2.8000 5.6565 2.8260 6.7500 ;
      RECT 2.6920 5.6565 2.7180 6.7500 ;
      RECT 2.5840 5.6565 2.6100 6.7500 ;
      RECT 2.4760 5.6565 2.5020 6.7500 ;
      RECT 2.3680 5.6565 2.3940 6.7500 ;
      RECT 2.2600 5.6565 2.2860 6.7500 ;
      RECT 2.1520 5.6565 2.1780 6.7500 ;
      RECT 2.0440 5.6565 2.0700 6.7500 ;
      RECT 1.9360 5.6565 1.9620 6.7500 ;
      RECT 1.8280 5.6565 1.8540 6.7500 ;
      RECT 1.7200 5.6565 1.7460 6.7500 ;
      RECT 1.6120 5.6565 1.6380 6.7500 ;
      RECT 1.5040 5.6565 1.5300 6.7500 ;
      RECT 1.3960 5.6565 1.4220 6.7500 ;
      RECT 1.2880 5.6565 1.3140 6.7500 ;
      RECT 1.1800 5.6565 1.2060 6.7500 ;
      RECT 1.0720 5.6565 1.0980 6.7500 ;
      RECT 0.9640 5.6565 0.9900 6.7500 ;
      RECT 0.8560 5.6565 0.8820 6.7500 ;
      RECT 0.7480 5.6565 0.7740 6.7500 ;
      RECT 0.6400 5.6565 0.6660 6.7500 ;
      RECT 0.5320 5.6565 0.5580 6.7500 ;
      RECT 0.4240 5.6565 0.4500 6.7500 ;
      RECT 0.3160 5.6565 0.3420 6.7500 ;
      RECT 0.2080 5.6565 0.2340 6.7500 ;
      RECT 0.0050 5.6565 0.0900 6.7500 ;
      RECT 8.6410 6.7365 8.7690 7.8300 ;
      RECT 8.6270 7.4020 8.7690 7.7245 ;
      RECT 8.4790 7.1290 8.5410 7.8300 ;
      RECT 8.4650 7.4385 8.5410 7.5920 ;
      RECT 8.4790 6.7365 8.5050 7.8300 ;
      RECT 8.4790 6.8575 8.5190 7.0970 ;
      RECT 8.4790 6.7365 8.5410 6.8255 ;
      RECT 8.1820 7.1870 8.3880 7.8300 ;
      RECT 8.3620 6.7365 8.3880 7.8300 ;
      RECT 8.1820 7.4640 8.4020 7.7220 ;
      RECT 8.1820 6.7365 8.2800 7.8300 ;
      RECT 7.7650 6.7365 7.8480 7.8300 ;
      RECT 7.7650 6.8250 7.8620 7.7605 ;
      RECT 16.4440 6.7365 16.5290 7.8300 ;
      RECT 16.3000 6.7365 16.3260 7.8300 ;
      RECT 16.1920 6.7365 16.2180 7.8300 ;
      RECT 16.0840 6.7365 16.1100 7.8300 ;
      RECT 15.9760 6.7365 16.0020 7.8300 ;
      RECT 15.8680 6.7365 15.8940 7.8300 ;
      RECT 15.7600 6.7365 15.7860 7.8300 ;
      RECT 15.6520 6.7365 15.6780 7.8300 ;
      RECT 15.5440 6.7365 15.5700 7.8300 ;
      RECT 15.4360 6.7365 15.4620 7.8300 ;
      RECT 15.3280 6.7365 15.3540 7.8300 ;
      RECT 15.2200 6.7365 15.2460 7.8300 ;
      RECT 15.1120 6.7365 15.1380 7.8300 ;
      RECT 15.0040 6.7365 15.0300 7.8300 ;
      RECT 14.8960 6.7365 14.9220 7.8300 ;
      RECT 14.7880 6.7365 14.8140 7.8300 ;
      RECT 14.6800 6.7365 14.7060 7.8300 ;
      RECT 14.5720 6.7365 14.5980 7.8300 ;
      RECT 14.4640 6.7365 14.4900 7.8300 ;
      RECT 14.3560 6.7365 14.3820 7.8300 ;
      RECT 14.2480 6.7365 14.2740 7.8300 ;
      RECT 14.1400 6.7365 14.1660 7.8300 ;
      RECT 14.0320 6.7365 14.0580 7.8300 ;
      RECT 13.9240 6.7365 13.9500 7.8300 ;
      RECT 13.8160 6.7365 13.8420 7.8300 ;
      RECT 13.7080 6.7365 13.7340 7.8300 ;
      RECT 13.6000 6.7365 13.6260 7.8300 ;
      RECT 13.4920 6.7365 13.5180 7.8300 ;
      RECT 13.3840 6.7365 13.4100 7.8300 ;
      RECT 13.2760 6.7365 13.3020 7.8300 ;
      RECT 13.1680 6.7365 13.1940 7.8300 ;
      RECT 13.0600 6.7365 13.0860 7.8300 ;
      RECT 12.9520 6.7365 12.9780 7.8300 ;
      RECT 12.8440 6.7365 12.8700 7.8300 ;
      RECT 12.7360 6.7365 12.7620 7.8300 ;
      RECT 12.6280 6.7365 12.6540 7.8300 ;
      RECT 12.5200 6.7365 12.5460 7.8300 ;
      RECT 12.4120 6.7365 12.4380 7.8300 ;
      RECT 12.3040 6.7365 12.3300 7.8300 ;
      RECT 12.1960 6.7365 12.2220 7.8300 ;
      RECT 12.0880 6.7365 12.1140 7.8300 ;
      RECT 11.9800 6.7365 12.0060 7.8300 ;
      RECT 11.8720 6.7365 11.8980 7.8300 ;
      RECT 11.7640 6.7365 11.7900 7.8300 ;
      RECT 11.6560 6.7365 11.6820 7.8300 ;
      RECT 11.5480 6.7365 11.5740 7.8300 ;
      RECT 11.4400 6.7365 11.4660 7.8300 ;
      RECT 11.3320 6.7365 11.3580 7.8300 ;
      RECT 11.2240 6.7365 11.2500 7.8300 ;
      RECT 11.1160 6.7365 11.1420 7.8300 ;
      RECT 11.0080 6.7365 11.0340 7.8300 ;
      RECT 10.9000 6.7365 10.9260 7.8300 ;
      RECT 10.7920 6.7365 10.8180 7.8300 ;
      RECT 10.6840 6.7365 10.7100 7.8300 ;
      RECT 10.5760 6.7365 10.6020 7.8300 ;
      RECT 10.4680 6.7365 10.4940 7.8300 ;
      RECT 10.3600 6.7365 10.3860 7.8300 ;
      RECT 10.2520 6.7365 10.2780 7.8300 ;
      RECT 10.1440 6.7365 10.1700 7.8300 ;
      RECT 10.0360 6.7365 10.0620 7.8300 ;
      RECT 9.9280 6.7365 9.9540 7.8300 ;
      RECT 9.8200 6.7365 9.8460 7.8300 ;
      RECT 9.7120 6.7365 9.7380 7.8300 ;
      RECT 9.6040 6.7365 9.6300 7.8300 ;
      RECT 9.4960 6.7365 9.5220 7.8300 ;
      RECT 9.3880 6.7365 9.4140 7.8300 ;
      RECT 9.1750 6.7365 9.2520 7.8300 ;
      RECT 7.2820 6.7365 7.3590 7.8300 ;
      RECT 7.1200 6.7365 7.1460 7.8300 ;
      RECT 7.0120 6.7365 7.0380 7.8300 ;
      RECT 6.9040 6.7365 6.9300 7.8300 ;
      RECT 6.7960 6.7365 6.8220 7.8300 ;
      RECT 6.6880 6.7365 6.7140 7.8300 ;
      RECT 6.5800 6.7365 6.6060 7.8300 ;
      RECT 6.4720 6.7365 6.4980 7.8300 ;
      RECT 6.3640 6.7365 6.3900 7.8300 ;
      RECT 6.2560 6.7365 6.2820 7.8300 ;
      RECT 6.1480 6.7365 6.1740 7.8300 ;
      RECT 6.0400 6.7365 6.0660 7.8300 ;
      RECT 5.9320 6.7365 5.9580 7.8300 ;
      RECT 5.8240 6.7365 5.8500 7.8300 ;
      RECT 5.7160 6.7365 5.7420 7.8300 ;
      RECT 5.6080 6.7365 5.6340 7.8300 ;
      RECT 5.5000 6.7365 5.5260 7.8300 ;
      RECT 5.3920 6.7365 5.4180 7.8300 ;
      RECT 5.2840 6.7365 5.3100 7.8300 ;
      RECT 5.1760 6.7365 5.2020 7.8300 ;
      RECT 5.0680 6.7365 5.0940 7.8300 ;
      RECT 4.9600 6.7365 4.9860 7.8300 ;
      RECT 4.8520 6.7365 4.8780 7.8300 ;
      RECT 4.7440 6.7365 4.7700 7.8300 ;
      RECT 4.6360 6.7365 4.6620 7.8300 ;
      RECT 4.5280 6.7365 4.5540 7.8300 ;
      RECT 4.4200 6.7365 4.4460 7.8300 ;
      RECT 4.3120 6.7365 4.3380 7.8300 ;
      RECT 4.2040 6.7365 4.2300 7.8300 ;
      RECT 4.0960 6.7365 4.1220 7.8300 ;
      RECT 3.9880 6.7365 4.0140 7.8300 ;
      RECT 3.8800 6.7365 3.9060 7.8300 ;
      RECT 3.7720 6.7365 3.7980 7.8300 ;
      RECT 3.6640 6.7365 3.6900 7.8300 ;
      RECT 3.5560 6.7365 3.5820 7.8300 ;
      RECT 3.4480 6.7365 3.4740 7.8300 ;
      RECT 3.3400 6.7365 3.3660 7.8300 ;
      RECT 3.2320 6.7365 3.2580 7.8300 ;
      RECT 3.1240 6.7365 3.1500 7.8300 ;
      RECT 3.0160 6.7365 3.0420 7.8300 ;
      RECT 2.9080 6.7365 2.9340 7.8300 ;
      RECT 2.8000 6.7365 2.8260 7.8300 ;
      RECT 2.6920 6.7365 2.7180 7.8300 ;
      RECT 2.5840 6.7365 2.6100 7.8300 ;
      RECT 2.4760 6.7365 2.5020 7.8300 ;
      RECT 2.3680 6.7365 2.3940 7.8300 ;
      RECT 2.2600 6.7365 2.2860 7.8300 ;
      RECT 2.1520 6.7365 2.1780 7.8300 ;
      RECT 2.0440 6.7365 2.0700 7.8300 ;
      RECT 1.9360 6.7365 1.9620 7.8300 ;
      RECT 1.8280 6.7365 1.8540 7.8300 ;
      RECT 1.7200 6.7365 1.7460 7.8300 ;
      RECT 1.6120 6.7365 1.6380 7.8300 ;
      RECT 1.5040 6.7365 1.5300 7.8300 ;
      RECT 1.3960 6.7365 1.4220 7.8300 ;
      RECT 1.2880 6.7365 1.3140 7.8300 ;
      RECT 1.1800 6.7365 1.2060 7.8300 ;
      RECT 1.0720 6.7365 1.0980 7.8300 ;
      RECT 0.9640 6.7365 0.9900 7.8300 ;
      RECT 0.8560 6.7365 0.8820 7.8300 ;
      RECT 0.7480 6.7365 0.7740 7.8300 ;
      RECT 0.6400 6.7365 0.6660 7.8300 ;
      RECT 0.5320 6.7365 0.5580 7.8300 ;
      RECT 0.4240 6.7365 0.4500 7.8300 ;
      RECT 0.3160 6.7365 0.3420 7.8300 ;
      RECT 0.2080 6.7365 0.2340 7.8300 ;
      RECT 0.0050 6.7365 0.0900 7.8300 ;
      RECT 8.6410 7.8165 8.7690 8.9100 ;
      RECT 8.6270 8.4820 8.7690 8.8045 ;
      RECT 8.4790 8.2090 8.5410 8.9100 ;
      RECT 8.4650 8.5185 8.5410 8.6720 ;
      RECT 8.4790 7.8165 8.5050 8.9100 ;
      RECT 8.4790 7.9375 8.5190 8.1770 ;
      RECT 8.4790 7.8165 8.5410 7.9055 ;
      RECT 8.1820 8.2670 8.3880 8.9100 ;
      RECT 8.3620 7.8165 8.3880 8.9100 ;
      RECT 8.1820 8.5440 8.4020 8.8020 ;
      RECT 8.1820 7.8165 8.2800 8.9100 ;
      RECT 7.7650 7.8165 7.8480 8.9100 ;
      RECT 7.7650 7.9050 7.8620 8.8405 ;
      RECT 16.4440 7.8165 16.5290 8.9100 ;
      RECT 16.3000 7.8165 16.3260 8.9100 ;
      RECT 16.1920 7.8165 16.2180 8.9100 ;
      RECT 16.0840 7.8165 16.1100 8.9100 ;
      RECT 15.9760 7.8165 16.0020 8.9100 ;
      RECT 15.8680 7.8165 15.8940 8.9100 ;
      RECT 15.7600 7.8165 15.7860 8.9100 ;
      RECT 15.6520 7.8165 15.6780 8.9100 ;
      RECT 15.5440 7.8165 15.5700 8.9100 ;
      RECT 15.4360 7.8165 15.4620 8.9100 ;
      RECT 15.3280 7.8165 15.3540 8.9100 ;
      RECT 15.2200 7.8165 15.2460 8.9100 ;
      RECT 15.1120 7.8165 15.1380 8.9100 ;
      RECT 15.0040 7.8165 15.0300 8.9100 ;
      RECT 14.8960 7.8165 14.9220 8.9100 ;
      RECT 14.7880 7.8165 14.8140 8.9100 ;
      RECT 14.6800 7.8165 14.7060 8.9100 ;
      RECT 14.5720 7.8165 14.5980 8.9100 ;
      RECT 14.4640 7.8165 14.4900 8.9100 ;
      RECT 14.3560 7.8165 14.3820 8.9100 ;
      RECT 14.2480 7.8165 14.2740 8.9100 ;
      RECT 14.1400 7.8165 14.1660 8.9100 ;
      RECT 14.0320 7.8165 14.0580 8.9100 ;
      RECT 13.9240 7.8165 13.9500 8.9100 ;
      RECT 13.8160 7.8165 13.8420 8.9100 ;
      RECT 13.7080 7.8165 13.7340 8.9100 ;
      RECT 13.6000 7.8165 13.6260 8.9100 ;
      RECT 13.4920 7.8165 13.5180 8.9100 ;
      RECT 13.3840 7.8165 13.4100 8.9100 ;
      RECT 13.2760 7.8165 13.3020 8.9100 ;
      RECT 13.1680 7.8165 13.1940 8.9100 ;
      RECT 13.0600 7.8165 13.0860 8.9100 ;
      RECT 12.9520 7.8165 12.9780 8.9100 ;
      RECT 12.8440 7.8165 12.8700 8.9100 ;
      RECT 12.7360 7.8165 12.7620 8.9100 ;
      RECT 12.6280 7.8165 12.6540 8.9100 ;
      RECT 12.5200 7.8165 12.5460 8.9100 ;
      RECT 12.4120 7.8165 12.4380 8.9100 ;
      RECT 12.3040 7.8165 12.3300 8.9100 ;
      RECT 12.1960 7.8165 12.2220 8.9100 ;
      RECT 12.0880 7.8165 12.1140 8.9100 ;
      RECT 11.9800 7.8165 12.0060 8.9100 ;
      RECT 11.8720 7.8165 11.8980 8.9100 ;
      RECT 11.7640 7.8165 11.7900 8.9100 ;
      RECT 11.6560 7.8165 11.6820 8.9100 ;
      RECT 11.5480 7.8165 11.5740 8.9100 ;
      RECT 11.4400 7.8165 11.4660 8.9100 ;
      RECT 11.3320 7.8165 11.3580 8.9100 ;
      RECT 11.2240 7.8165 11.2500 8.9100 ;
      RECT 11.1160 7.8165 11.1420 8.9100 ;
      RECT 11.0080 7.8165 11.0340 8.9100 ;
      RECT 10.9000 7.8165 10.9260 8.9100 ;
      RECT 10.7920 7.8165 10.8180 8.9100 ;
      RECT 10.6840 7.8165 10.7100 8.9100 ;
      RECT 10.5760 7.8165 10.6020 8.9100 ;
      RECT 10.4680 7.8165 10.4940 8.9100 ;
      RECT 10.3600 7.8165 10.3860 8.9100 ;
      RECT 10.2520 7.8165 10.2780 8.9100 ;
      RECT 10.1440 7.8165 10.1700 8.9100 ;
      RECT 10.0360 7.8165 10.0620 8.9100 ;
      RECT 9.9280 7.8165 9.9540 8.9100 ;
      RECT 9.8200 7.8165 9.8460 8.9100 ;
      RECT 9.7120 7.8165 9.7380 8.9100 ;
      RECT 9.6040 7.8165 9.6300 8.9100 ;
      RECT 9.4960 7.8165 9.5220 8.9100 ;
      RECT 9.3880 7.8165 9.4140 8.9100 ;
      RECT 9.1750 7.8165 9.2520 8.9100 ;
      RECT 7.2820 7.8165 7.3590 8.9100 ;
      RECT 7.1200 7.8165 7.1460 8.9100 ;
      RECT 7.0120 7.8165 7.0380 8.9100 ;
      RECT 6.9040 7.8165 6.9300 8.9100 ;
      RECT 6.7960 7.8165 6.8220 8.9100 ;
      RECT 6.6880 7.8165 6.7140 8.9100 ;
      RECT 6.5800 7.8165 6.6060 8.9100 ;
      RECT 6.4720 7.8165 6.4980 8.9100 ;
      RECT 6.3640 7.8165 6.3900 8.9100 ;
      RECT 6.2560 7.8165 6.2820 8.9100 ;
      RECT 6.1480 7.8165 6.1740 8.9100 ;
      RECT 6.0400 7.8165 6.0660 8.9100 ;
      RECT 5.9320 7.8165 5.9580 8.9100 ;
      RECT 5.8240 7.8165 5.8500 8.9100 ;
      RECT 5.7160 7.8165 5.7420 8.9100 ;
      RECT 5.6080 7.8165 5.6340 8.9100 ;
      RECT 5.5000 7.8165 5.5260 8.9100 ;
      RECT 5.3920 7.8165 5.4180 8.9100 ;
      RECT 5.2840 7.8165 5.3100 8.9100 ;
      RECT 5.1760 7.8165 5.2020 8.9100 ;
      RECT 5.0680 7.8165 5.0940 8.9100 ;
      RECT 4.9600 7.8165 4.9860 8.9100 ;
      RECT 4.8520 7.8165 4.8780 8.9100 ;
      RECT 4.7440 7.8165 4.7700 8.9100 ;
      RECT 4.6360 7.8165 4.6620 8.9100 ;
      RECT 4.5280 7.8165 4.5540 8.9100 ;
      RECT 4.4200 7.8165 4.4460 8.9100 ;
      RECT 4.3120 7.8165 4.3380 8.9100 ;
      RECT 4.2040 7.8165 4.2300 8.9100 ;
      RECT 4.0960 7.8165 4.1220 8.9100 ;
      RECT 3.9880 7.8165 4.0140 8.9100 ;
      RECT 3.8800 7.8165 3.9060 8.9100 ;
      RECT 3.7720 7.8165 3.7980 8.9100 ;
      RECT 3.6640 7.8165 3.6900 8.9100 ;
      RECT 3.5560 7.8165 3.5820 8.9100 ;
      RECT 3.4480 7.8165 3.4740 8.9100 ;
      RECT 3.3400 7.8165 3.3660 8.9100 ;
      RECT 3.2320 7.8165 3.2580 8.9100 ;
      RECT 3.1240 7.8165 3.1500 8.9100 ;
      RECT 3.0160 7.8165 3.0420 8.9100 ;
      RECT 2.9080 7.8165 2.9340 8.9100 ;
      RECT 2.8000 7.8165 2.8260 8.9100 ;
      RECT 2.6920 7.8165 2.7180 8.9100 ;
      RECT 2.5840 7.8165 2.6100 8.9100 ;
      RECT 2.4760 7.8165 2.5020 8.9100 ;
      RECT 2.3680 7.8165 2.3940 8.9100 ;
      RECT 2.2600 7.8165 2.2860 8.9100 ;
      RECT 2.1520 7.8165 2.1780 8.9100 ;
      RECT 2.0440 7.8165 2.0700 8.9100 ;
      RECT 1.9360 7.8165 1.9620 8.9100 ;
      RECT 1.8280 7.8165 1.8540 8.9100 ;
      RECT 1.7200 7.8165 1.7460 8.9100 ;
      RECT 1.6120 7.8165 1.6380 8.9100 ;
      RECT 1.5040 7.8165 1.5300 8.9100 ;
      RECT 1.3960 7.8165 1.4220 8.9100 ;
      RECT 1.2880 7.8165 1.3140 8.9100 ;
      RECT 1.1800 7.8165 1.2060 8.9100 ;
      RECT 1.0720 7.8165 1.0980 8.9100 ;
      RECT 0.9640 7.8165 0.9900 8.9100 ;
      RECT 0.8560 7.8165 0.8820 8.9100 ;
      RECT 0.7480 7.8165 0.7740 8.9100 ;
      RECT 0.6400 7.8165 0.6660 8.9100 ;
      RECT 0.5320 7.8165 0.5580 8.9100 ;
      RECT 0.4240 7.8165 0.4500 8.9100 ;
      RECT 0.3160 7.8165 0.3420 8.9100 ;
      RECT 0.2080 7.8165 0.2340 8.9100 ;
      RECT 0.0050 7.8165 0.0900 8.9100 ;
      RECT 8.6410 8.8965 8.7690 9.9900 ;
      RECT 8.6270 9.5620 8.7690 9.8845 ;
      RECT 8.4790 9.2890 8.5410 9.9900 ;
      RECT 8.4650 9.5985 8.5410 9.7520 ;
      RECT 8.4790 8.8965 8.5050 9.9900 ;
      RECT 8.4790 9.0175 8.5190 9.2570 ;
      RECT 8.4790 8.8965 8.5410 8.9855 ;
      RECT 8.1820 9.3470 8.3880 9.9900 ;
      RECT 8.3620 8.8965 8.3880 9.9900 ;
      RECT 8.1820 9.6240 8.4020 9.8820 ;
      RECT 8.1820 8.8965 8.2800 9.9900 ;
      RECT 7.7650 8.8965 7.8480 9.9900 ;
      RECT 7.7650 8.9850 7.8620 9.9205 ;
      RECT 16.4440 8.8965 16.5290 9.9900 ;
      RECT 16.3000 8.8965 16.3260 9.9900 ;
      RECT 16.1920 8.8965 16.2180 9.9900 ;
      RECT 16.0840 8.8965 16.1100 9.9900 ;
      RECT 15.9760 8.8965 16.0020 9.9900 ;
      RECT 15.8680 8.8965 15.8940 9.9900 ;
      RECT 15.7600 8.8965 15.7860 9.9900 ;
      RECT 15.6520 8.8965 15.6780 9.9900 ;
      RECT 15.5440 8.8965 15.5700 9.9900 ;
      RECT 15.4360 8.8965 15.4620 9.9900 ;
      RECT 15.3280 8.8965 15.3540 9.9900 ;
      RECT 15.2200 8.8965 15.2460 9.9900 ;
      RECT 15.1120 8.8965 15.1380 9.9900 ;
      RECT 15.0040 8.8965 15.0300 9.9900 ;
      RECT 14.8960 8.8965 14.9220 9.9900 ;
      RECT 14.7880 8.8965 14.8140 9.9900 ;
      RECT 14.6800 8.8965 14.7060 9.9900 ;
      RECT 14.5720 8.8965 14.5980 9.9900 ;
      RECT 14.4640 8.8965 14.4900 9.9900 ;
      RECT 14.3560 8.8965 14.3820 9.9900 ;
      RECT 14.2480 8.8965 14.2740 9.9900 ;
      RECT 14.1400 8.8965 14.1660 9.9900 ;
      RECT 14.0320 8.8965 14.0580 9.9900 ;
      RECT 13.9240 8.8965 13.9500 9.9900 ;
      RECT 13.8160 8.8965 13.8420 9.9900 ;
      RECT 13.7080 8.8965 13.7340 9.9900 ;
      RECT 13.6000 8.8965 13.6260 9.9900 ;
      RECT 13.4920 8.8965 13.5180 9.9900 ;
      RECT 13.3840 8.8965 13.4100 9.9900 ;
      RECT 13.2760 8.8965 13.3020 9.9900 ;
      RECT 13.1680 8.8965 13.1940 9.9900 ;
      RECT 13.0600 8.8965 13.0860 9.9900 ;
      RECT 12.9520 8.8965 12.9780 9.9900 ;
      RECT 12.8440 8.8965 12.8700 9.9900 ;
      RECT 12.7360 8.8965 12.7620 9.9900 ;
      RECT 12.6280 8.8965 12.6540 9.9900 ;
      RECT 12.5200 8.8965 12.5460 9.9900 ;
      RECT 12.4120 8.8965 12.4380 9.9900 ;
      RECT 12.3040 8.8965 12.3300 9.9900 ;
      RECT 12.1960 8.8965 12.2220 9.9900 ;
      RECT 12.0880 8.8965 12.1140 9.9900 ;
      RECT 11.9800 8.8965 12.0060 9.9900 ;
      RECT 11.8720 8.8965 11.8980 9.9900 ;
      RECT 11.7640 8.8965 11.7900 9.9900 ;
      RECT 11.6560 8.8965 11.6820 9.9900 ;
      RECT 11.5480 8.8965 11.5740 9.9900 ;
      RECT 11.4400 8.8965 11.4660 9.9900 ;
      RECT 11.3320 8.8965 11.3580 9.9900 ;
      RECT 11.2240 8.8965 11.2500 9.9900 ;
      RECT 11.1160 8.8965 11.1420 9.9900 ;
      RECT 11.0080 8.8965 11.0340 9.9900 ;
      RECT 10.9000 8.8965 10.9260 9.9900 ;
      RECT 10.7920 8.8965 10.8180 9.9900 ;
      RECT 10.6840 8.8965 10.7100 9.9900 ;
      RECT 10.5760 8.8965 10.6020 9.9900 ;
      RECT 10.4680 8.8965 10.4940 9.9900 ;
      RECT 10.3600 8.8965 10.3860 9.9900 ;
      RECT 10.2520 8.8965 10.2780 9.9900 ;
      RECT 10.1440 8.8965 10.1700 9.9900 ;
      RECT 10.0360 8.8965 10.0620 9.9900 ;
      RECT 9.9280 8.8965 9.9540 9.9900 ;
      RECT 9.8200 8.8965 9.8460 9.9900 ;
      RECT 9.7120 8.8965 9.7380 9.9900 ;
      RECT 9.6040 8.8965 9.6300 9.9900 ;
      RECT 9.4960 8.8965 9.5220 9.9900 ;
      RECT 9.3880 8.8965 9.4140 9.9900 ;
      RECT 9.1750 8.8965 9.2520 9.9900 ;
      RECT 7.2820 8.8965 7.3590 9.9900 ;
      RECT 7.1200 8.8965 7.1460 9.9900 ;
      RECT 7.0120 8.8965 7.0380 9.9900 ;
      RECT 6.9040 8.8965 6.9300 9.9900 ;
      RECT 6.7960 8.8965 6.8220 9.9900 ;
      RECT 6.6880 8.8965 6.7140 9.9900 ;
      RECT 6.5800 8.8965 6.6060 9.9900 ;
      RECT 6.4720 8.8965 6.4980 9.9900 ;
      RECT 6.3640 8.8965 6.3900 9.9900 ;
      RECT 6.2560 8.8965 6.2820 9.9900 ;
      RECT 6.1480 8.8965 6.1740 9.9900 ;
      RECT 6.0400 8.8965 6.0660 9.9900 ;
      RECT 5.9320 8.8965 5.9580 9.9900 ;
      RECT 5.8240 8.8965 5.8500 9.9900 ;
      RECT 5.7160 8.8965 5.7420 9.9900 ;
      RECT 5.6080 8.8965 5.6340 9.9900 ;
      RECT 5.5000 8.8965 5.5260 9.9900 ;
      RECT 5.3920 8.8965 5.4180 9.9900 ;
      RECT 5.2840 8.8965 5.3100 9.9900 ;
      RECT 5.1760 8.8965 5.2020 9.9900 ;
      RECT 5.0680 8.8965 5.0940 9.9900 ;
      RECT 4.9600 8.8965 4.9860 9.9900 ;
      RECT 4.8520 8.8965 4.8780 9.9900 ;
      RECT 4.7440 8.8965 4.7700 9.9900 ;
      RECT 4.6360 8.8965 4.6620 9.9900 ;
      RECT 4.5280 8.8965 4.5540 9.9900 ;
      RECT 4.4200 8.8965 4.4460 9.9900 ;
      RECT 4.3120 8.8965 4.3380 9.9900 ;
      RECT 4.2040 8.8965 4.2300 9.9900 ;
      RECT 4.0960 8.8965 4.1220 9.9900 ;
      RECT 3.9880 8.8965 4.0140 9.9900 ;
      RECT 3.8800 8.8965 3.9060 9.9900 ;
      RECT 3.7720 8.8965 3.7980 9.9900 ;
      RECT 3.6640 8.8965 3.6900 9.9900 ;
      RECT 3.5560 8.8965 3.5820 9.9900 ;
      RECT 3.4480 8.8965 3.4740 9.9900 ;
      RECT 3.3400 8.8965 3.3660 9.9900 ;
      RECT 3.2320 8.8965 3.2580 9.9900 ;
      RECT 3.1240 8.8965 3.1500 9.9900 ;
      RECT 3.0160 8.8965 3.0420 9.9900 ;
      RECT 2.9080 8.8965 2.9340 9.9900 ;
      RECT 2.8000 8.8965 2.8260 9.9900 ;
      RECT 2.6920 8.8965 2.7180 9.9900 ;
      RECT 2.5840 8.8965 2.6100 9.9900 ;
      RECT 2.4760 8.8965 2.5020 9.9900 ;
      RECT 2.3680 8.8965 2.3940 9.9900 ;
      RECT 2.2600 8.8965 2.2860 9.9900 ;
      RECT 2.1520 8.8965 2.1780 9.9900 ;
      RECT 2.0440 8.8965 2.0700 9.9900 ;
      RECT 1.9360 8.8965 1.9620 9.9900 ;
      RECT 1.8280 8.8965 1.8540 9.9900 ;
      RECT 1.7200 8.8965 1.7460 9.9900 ;
      RECT 1.6120 8.8965 1.6380 9.9900 ;
      RECT 1.5040 8.8965 1.5300 9.9900 ;
      RECT 1.3960 8.8965 1.4220 9.9900 ;
      RECT 1.2880 8.8965 1.3140 9.9900 ;
      RECT 1.1800 8.8965 1.2060 9.9900 ;
      RECT 1.0720 8.8965 1.0980 9.9900 ;
      RECT 0.9640 8.8965 0.9900 9.9900 ;
      RECT 0.8560 8.8965 0.8820 9.9900 ;
      RECT 0.7480 8.8965 0.7740 9.9900 ;
      RECT 0.6400 8.8965 0.6660 9.9900 ;
      RECT 0.5320 8.8965 0.5580 9.9900 ;
      RECT 0.4240 8.8965 0.4500 9.9900 ;
      RECT 0.3160 8.8965 0.3420 9.9900 ;
      RECT 0.2080 8.8965 0.2340 9.9900 ;
      RECT 0.0050 8.8965 0.0900 9.9900 ;
      RECT 8.6410 9.9765 8.7690 11.0700 ;
      RECT 8.6270 10.6420 8.7690 10.9645 ;
      RECT 8.4790 10.3690 8.5410 11.0700 ;
      RECT 8.4650 10.6785 8.5410 10.8320 ;
      RECT 8.4790 9.9765 8.5050 11.0700 ;
      RECT 8.4790 10.0975 8.5190 10.3370 ;
      RECT 8.4790 9.9765 8.5410 10.0655 ;
      RECT 8.1820 10.4270 8.3880 11.0700 ;
      RECT 8.3620 9.9765 8.3880 11.0700 ;
      RECT 8.1820 10.7040 8.4020 10.9620 ;
      RECT 8.1820 9.9765 8.2800 11.0700 ;
      RECT 7.7650 9.9765 7.8480 11.0700 ;
      RECT 7.7650 10.0650 7.8620 11.0005 ;
      RECT 16.4440 9.9765 16.5290 11.0700 ;
      RECT 16.3000 9.9765 16.3260 11.0700 ;
      RECT 16.1920 9.9765 16.2180 11.0700 ;
      RECT 16.0840 9.9765 16.1100 11.0700 ;
      RECT 15.9760 9.9765 16.0020 11.0700 ;
      RECT 15.8680 9.9765 15.8940 11.0700 ;
      RECT 15.7600 9.9765 15.7860 11.0700 ;
      RECT 15.6520 9.9765 15.6780 11.0700 ;
      RECT 15.5440 9.9765 15.5700 11.0700 ;
      RECT 15.4360 9.9765 15.4620 11.0700 ;
      RECT 15.3280 9.9765 15.3540 11.0700 ;
      RECT 15.2200 9.9765 15.2460 11.0700 ;
      RECT 15.1120 9.9765 15.1380 11.0700 ;
      RECT 15.0040 9.9765 15.0300 11.0700 ;
      RECT 14.8960 9.9765 14.9220 11.0700 ;
      RECT 14.7880 9.9765 14.8140 11.0700 ;
      RECT 14.6800 9.9765 14.7060 11.0700 ;
      RECT 14.5720 9.9765 14.5980 11.0700 ;
      RECT 14.4640 9.9765 14.4900 11.0700 ;
      RECT 14.3560 9.9765 14.3820 11.0700 ;
      RECT 14.2480 9.9765 14.2740 11.0700 ;
      RECT 14.1400 9.9765 14.1660 11.0700 ;
      RECT 14.0320 9.9765 14.0580 11.0700 ;
      RECT 13.9240 9.9765 13.9500 11.0700 ;
      RECT 13.8160 9.9765 13.8420 11.0700 ;
      RECT 13.7080 9.9765 13.7340 11.0700 ;
      RECT 13.6000 9.9765 13.6260 11.0700 ;
      RECT 13.4920 9.9765 13.5180 11.0700 ;
      RECT 13.3840 9.9765 13.4100 11.0700 ;
      RECT 13.2760 9.9765 13.3020 11.0700 ;
      RECT 13.1680 9.9765 13.1940 11.0700 ;
      RECT 13.0600 9.9765 13.0860 11.0700 ;
      RECT 12.9520 9.9765 12.9780 11.0700 ;
      RECT 12.8440 9.9765 12.8700 11.0700 ;
      RECT 12.7360 9.9765 12.7620 11.0700 ;
      RECT 12.6280 9.9765 12.6540 11.0700 ;
      RECT 12.5200 9.9765 12.5460 11.0700 ;
      RECT 12.4120 9.9765 12.4380 11.0700 ;
      RECT 12.3040 9.9765 12.3300 11.0700 ;
      RECT 12.1960 9.9765 12.2220 11.0700 ;
      RECT 12.0880 9.9765 12.1140 11.0700 ;
      RECT 11.9800 9.9765 12.0060 11.0700 ;
      RECT 11.8720 9.9765 11.8980 11.0700 ;
      RECT 11.7640 9.9765 11.7900 11.0700 ;
      RECT 11.6560 9.9765 11.6820 11.0700 ;
      RECT 11.5480 9.9765 11.5740 11.0700 ;
      RECT 11.4400 9.9765 11.4660 11.0700 ;
      RECT 11.3320 9.9765 11.3580 11.0700 ;
      RECT 11.2240 9.9765 11.2500 11.0700 ;
      RECT 11.1160 9.9765 11.1420 11.0700 ;
      RECT 11.0080 9.9765 11.0340 11.0700 ;
      RECT 10.9000 9.9765 10.9260 11.0700 ;
      RECT 10.7920 9.9765 10.8180 11.0700 ;
      RECT 10.6840 9.9765 10.7100 11.0700 ;
      RECT 10.5760 9.9765 10.6020 11.0700 ;
      RECT 10.4680 9.9765 10.4940 11.0700 ;
      RECT 10.3600 9.9765 10.3860 11.0700 ;
      RECT 10.2520 9.9765 10.2780 11.0700 ;
      RECT 10.1440 9.9765 10.1700 11.0700 ;
      RECT 10.0360 9.9765 10.0620 11.0700 ;
      RECT 9.9280 9.9765 9.9540 11.0700 ;
      RECT 9.8200 9.9765 9.8460 11.0700 ;
      RECT 9.7120 9.9765 9.7380 11.0700 ;
      RECT 9.6040 9.9765 9.6300 11.0700 ;
      RECT 9.4960 9.9765 9.5220 11.0700 ;
      RECT 9.3880 9.9765 9.4140 11.0700 ;
      RECT 9.1750 9.9765 9.2520 11.0700 ;
      RECT 7.2820 9.9765 7.3590 11.0700 ;
      RECT 7.1200 9.9765 7.1460 11.0700 ;
      RECT 7.0120 9.9765 7.0380 11.0700 ;
      RECT 6.9040 9.9765 6.9300 11.0700 ;
      RECT 6.7960 9.9765 6.8220 11.0700 ;
      RECT 6.6880 9.9765 6.7140 11.0700 ;
      RECT 6.5800 9.9765 6.6060 11.0700 ;
      RECT 6.4720 9.9765 6.4980 11.0700 ;
      RECT 6.3640 9.9765 6.3900 11.0700 ;
      RECT 6.2560 9.9765 6.2820 11.0700 ;
      RECT 6.1480 9.9765 6.1740 11.0700 ;
      RECT 6.0400 9.9765 6.0660 11.0700 ;
      RECT 5.9320 9.9765 5.9580 11.0700 ;
      RECT 5.8240 9.9765 5.8500 11.0700 ;
      RECT 5.7160 9.9765 5.7420 11.0700 ;
      RECT 5.6080 9.9765 5.6340 11.0700 ;
      RECT 5.5000 9.9765 5.5260 11.0700 ;
      RECT 5.3920 9.9765 5.4180 11.0700 ;
      RECT 5.2840 9.9765 5.3100 11.0700 ;
      RECT 5.1760 9.9765 5.2020 11.0700 ;
      RECT 5.0680 9.9765 5.0940 11.0700 ;
      RECT 4.9600 9.9765 4.9860 11.0700 ;
      RECT 4.8520 9.9765 4.8780 11.0700 ;
      RECT 4.7440 9.9765 4.7700 11.0700 ;
      RECT 4.6360 9.9765 4.6620 11.0700 ;
      RECT 4.5280 9.9765 4.5540 11.0700 ;
      RECT 4.4200 9.9765 4.4460 11.0700 ;
      RECT 4.3120 9.9765 4.3380 11.0700 ;
      RECT 4.2040 9.9765 4.2300 11.0700 ;
      RECT 4.0960 9.9765 4.1220 11.0700 ;
      RECT 3.9880 9.9765 4.0140 11.0700 ;
      RECT 3.8800 9.9765 3.9060 11.0700 ;
      RECT 3.7720 9.9765 3.7980 11.0700 ;
      RECT 3.6640 9.9765 3.6900 11.0700 ;
      RECT 3.5560 9.9765 3.5820 11.0700 ;
      RECT 3.4480 9.9765 3.4740 11.0700 ;
      RECT 3.3400 9.9765 3.3660 11.0700 ;
      RECT 3.2320 9.9765 3.2580 11.0700 ;
      RECT 3.1240 9.9765 3.1500 11.0700 ;
      RECT 3.0160 9.9765 3.0420 11.0700 ;
      RECT 2.9080 9.9765 2.9340 11.0700 ;
      RECT 2.8000 9.9765 2.8260 11.0700 ;
      RECT 2.6920 9.9765 2.7180 11.0700 ;
      RECT 2.5840 9.9765 2.6100 11.0700 ;
      RECT 2.4760 9.9765 2.5020 11.0700 ;
      RECT 2.3680 9.9765 2.3940 11.0700 ;
      RECT 2.2600 9.9765 2.2860 11.0700 ;
      RECT 2.1520 9.9765 2.1780 11.0700 ;
      RECT 2.0440 9.9765 2.0700 11.0700 ;
      RECT 1.9360 9.9765 1.9620 11.0700 ;
      RECT 1.8280 9.9765 1.8540 11.0700 ;
      RECT 1.7200 9.9765 1.7460 11.0700 ;
      RECT 1.6120 9.9765 1.6380 11.0700 ;
      RECT 1.5040 9.9765 1.5300 11.0700 ;
      RECT 1.3960 9.9765 1.4220 11.0700 ;
      RECT 1.2880 9.9765 1.3140 11.0700 ;
      RECT 1.1800 9.9765 1.2060 11.0700 ;
      RECT 1.0720 9.9765 1.0980 11.0700 ;
      RECT 0.9640 9.9765 0.9900 11.0700 ;
      RECT 0.8560 9.9765 0.8820 11.0700 ;
      RECT 0.7480 9.9765 0.7740 11.0700 ;
      RECT 0.6400 9.9765 0.6660 11.0700 ;
      RECT 0.5320 9.9765 0.5580 11.0700 ;
      RECT 0.4240 9.9765 0.4500 11.0700 ;
      RECT 0.3160 9.9765 0.3420 11.0700 ;
      RECT 0.2080 9.9765 0.2340 11.0700 ;
      RECT 0.0050 9.9765 0.0900 11.0700 ;
      RECT 8.6410 11.0565 8.7690 12.1500 ;
      RECT 8.6270 11.7220 8.7690 12.0445 ;
      RECT 8.4790 11.4490 8.5410 12.1500 ;
      RECT 8.4650 11.7585 8.5410 11.9120 ;
      RECT 8.4790 11.0565 8.5050 12.1500 ;
      RECT 8.4790 11.1775 8.5190 11.4170 ;
      RECT 8.4790 11.0565 8.5410 11.1455 ;
      RECT 8.1820 11.5070 8.3880 12.1500 ;
      RECT 8.3620 11.0565 8.3880 12.1500 ;
      RECT 8.1820 11.7840 8.4020 12.0420 ;
      RECT 8.1820 11.0565 8.2800 12.1500 ;
      RECT 7.7650 11.0565 7.8480 12.1500 ;
      RECT 7.7650 11.1450 7.8620 12.0805 ;
      RECT 16.4440 11.0565 16.5290 12.1500 ;
      RECT 16.3000 11.0565 16.3260 12.1500 ;
      RECT 16.1920 11.0565 16.2180 12.1500 ;
      RECT 16.0840 11.0565 16.1100 12.1500 ;
      RECT 15.9760 11.0565 16.0020 12.1500 ;
      RECT 15.8680 11.0565 15.8940 12.1500 ;
      RECT 15.7600 11.0565 15.7860 12.1500 ;
      RECT 15.6520 11.0565 15.6780 12.1500 ;
      RECT 15.5440 11.0565 15.5700 12.1500 ;
      RECT 15.4360 11.0565 15.4620 12.1500 ;
      RECT 15.3280 11.0565 15.3540 12.1500 ;
      RECT 15.2200 11.0565 15.2460 12.1500 ;
      RECT 15.1120 11.0565 15.1380 12.1500 ;
      RECT 15.0040 11.0565 15.0300 12.1500 ;
      RECT 14.8960 11.0565 14.9220 12.1500 ;
      RECT 14.7880 11.0565 14.8140 12.1500 ;
      RECT 14.6800 11.0565 14.7060 12.1500 ;
      RECT 14.5720 11.0565 14.5980 12.1500 ;
      RECT 14.4640 11.0565 14.4900 12.1500 ;
      RECT 14.3560 11.0565 14.3820 12.1500 ;
      RECT 14.2480 11.0565 14.2740 12.1500 ;
      RECT 14.1400 11.0565 14.1660 12.1500 ;
      RECT 14.0320 11.0565 14.0580 12.1500 ;
      RECT 13.9240 11.0565 13.9500 12.1500 ;
      RECT 13.8160 11.0565 13.8420 12.1500 ;
      RECT 13.7080 11.0565 13.7340 12.1500 ;
      RECT 13.6000 11.0565 13.6260 12.1500 ;
      RECT 13.4920 11.0565 13.5180 12.1500 ;
      RECT 13.3840 11.0565 13.4100 12.1500 ;
      RECT 13.2760 11.0565 13.3020 12.1500 ;
      RECT 13.1680 11.0565 13.1940 12.1500 ;
      RECT 13.0600 11.0565 13.0860 12.1500 ;
      RECT 12.9520 11.0565 12.9780 12.1500 ;
      RECT 12.8440 11.0565 12.8700 12.1500 ;
      RECT 12.7360 11.0565 12.7620 12.1500 ;
      RECT 12.6280 11.0565 12.6540 12.1500 ;
      RECT 12.5200 11.0565 12.5460 12.1500 ;
      RECT 12.4120 11.0565 12.4380 12.1500 ;
      RECT 12.3040 11.0565 12.3300 12.1500 ;
      RECT 12.1960 11.0565 12.2220 12.1500 ;
      RECT 12.0880 11.0565 12.1140 12.1500 ;
      RECT 11.9800 11.0565 12.0060 12.1500 ;
      RECT 11.8720 11.0565 11.8980 12.1500 ;
      RECT 11.7640 11.0565 11.7900 12.1500 ;
      RECT 11.6560 11.0565 11.6820 12.1500 ;
      RECT 11.5480 11.0565 11.5740 12.1500 ;
      RECT 11.4400 11.0565 11.4660 12.1500 ;
      RECT 11.3320 11.0565 11.3580 12.1500 ;
      RECT 11.2240 11.0565 11.2500 12.1500 ;
      RECT 11.1160 11.0565 11.1420 12.1500 ;
      RECT 11.0080 11.0565 11.0340 12.1500 ;
      RECT 10.9000 11.0565 10.9260 12.1500 ;
      RECT 10.7920 11.0565 10.8180 12.1500 ;
      RECT 10.6840 11.0565 10.7100 12.1500 ;
      RECT 10.5760 11.0565 10.6020 12.1500 ;
      RECT 10.4680 11.0565 10.4940 12.1500 ;
      RECT 10.3600 11.0565 10.3860 12.1500 ;
      RECT 10.2520 11.0565 10.2780 12.1500 ;
      RECT 10.1440 11.0565 10.1700 12.1500 ;
      RECT 10.0360 11.0565 10.0620 12.1500 ;
      RECT 9.9280 11.0565 9.9540 12.1500 ;
      RECT 9.8200 11.0565 9.8460 12.1500 ;
      RECT 9.7120 11.0565 9.7380 12.1500 ;
      RECT 9.6040 11.0565 9.6300 12.1500 ;
      RECT 9.4960 11.0565 9.5220 12.1500 ;
      RECT 9.3880 11.0565 9.4140 12.1500 ;
      RECT 9.1750 11.0565 9.2520 12.1500 ;
      RECT 7.2820 11.0565 7.3590 12.1500 ;
      RECT 7.1200 11.0565 7.1460 12.1500 ;
      RECT 7.0120 11.0565 7.0380 12.1500 ;
      RECT 6.9040 11.0565 6.9300 12.1500 ;
      RECT 6.7960 11.0565 6.8220 12.1500 ;
      RECT 6.6880 11.0565 6.7140 12.1500 ;
      RECT 6.5800 11.0565 6.6060 12.1500 ;
      RECT 6.4720 11.0565 6.4980 12.1500 ;
      RECT 6.3640 11.0565 6.3900 12.1500 ;
      RECT 6.2560 11.0565 6.2820 12.1500 ;
      RECT 6.1480 11.0565 6.1740 12.1500 ;
      RECT 6.0400 11.0565 6.0660 12.1500 ;
      RECT 5.9320 11.0565 5.9580 12.1500 ;
      RECT 5.8240 11.0565 5.8500 12.1500 ;
      RECT 5.7160 11.0565 5.7420 12.1500 ;
      RECT 5.6080 11.0565 5.6340 12.1500 ;
      RECT 5.5000 11.0565 5.5260 12.1500 ;
      RECT 5.3920 11.0565 5.4180 12.1500 ;
      RECT 5.2840 11.0565 5.3100 12.1500 ;
      RECT 5.1760 11.0565 5.2020 12.1500 ;
      RECT 5.0680 11.0565 5.0940 12.1500 ;
      RECT 4.9600 11.0565 4.9860 12.1500 ;
      RECT 4.8520 11.0565 4.8780 12.1500 ;
      RECT 4.7440 11.0565 4.7700 12.1500 ;
      RECT 4.6360 11.0565 4.6620 12.1500 ;
      RECT 4.5280 11.0565 4.5540 12.1500 ;
      RECT 4.4200 11.0565 4.4460 12.1500 ;
      RECT 4.3120 11.0565 4.3380 12.1500 ;
      RECT 4.2040 11.0565 4.2300 12.1500 ;
      RECT 4.0960 11.0565 4.1220 12.1500 ;
      RECT 3.9880 11.0565 4.0140 12.1500 ;
      RECT 3.8800 11.0565 3.9060 12.1500 ;
      RECT 3.7720 11.0565 3.7980 12.1500 ;
      RECT 3.6640 11.0565 3.6900 12.1500 ;
      RECT 3.5560 11.0565 3.5820 12.1500 ;
      RECT 3.4480 11.0565 3.4740 12.1500 ;
      RECT 3.3400 11.0565 3.3660 12.1500 ;
      RECT 3.2320 11.0565 3.2580 12.1500 ;
      RECT 3.1240 11.0565 3.1500 12.1500 ;
      RECT 3.0160 11.0565 3.0420 12.1500 ;
      RECT 2.9080 11.0565 2.9340 12.1500 ;
      RECT 2.8000 11.0565 2.8260 12.1500 ;
      RECT 2.6920 11.0565 2.7180 12.1500 ;
      RECT 2.5840 11.0565 2.6100 12.1500 ;
      RECT 2.4760 11.0565 2.5020 12.1500 ;
      RECT 2.3680 11.0565 2.3940 12.1500 ;
      RECT 2.2600 11.0565 2.2860 12.1500 ;
      RECT 2.1520 11.0565 2.1780 12.1500 ;
      RECT 2.0440 11.0565 2.0700 12.1500 ;
      RECT 1.9360 11.0565 1.9620 12.1500 ;
      RECT 1.8280 11.0565 1.8540 12.1500 ;
      RECT 1.7200 11.0565 1.7460 12.1500 ;
      RECT 1.6120 11.0565 1.6380 12.1500 ;
      RECT 1.5040 11.0565 1.5300 12.1500 ;
      RECT 1.3960 11.0565 1.4220 12.1500 ;
      RECT 1.2880 11.0565 1.3140 12.1500 ;
      RECT 1.1800 11.0565 1.2060 12.1500 ;
      RECT 1.0720 11.0565 1.0980 12.1500 ;
      RECT 0.9640 11.0565 0.9900 12.1500 ;
      RECT 0.8560 11.0565 0.8820 12.1500 ;
      RECT 0.7480 11.0565 0.7740 12.1500 ;
      RECT 0.6400 11.0565 0.6660 12.1500 ;
      RECT 0.5320 11.0565 0.5580 12.1500 ;
      RECT 0.4240 11.0565 0.4500 12.1500 ;
      RECT 0.3160 11.0565 0.3420 12.1500 ;
      RECT 0.2080 11.0565 0.2340 12.1500 ;
      RECT 0.0050 11.0565 0.0900 12.1500 ;
      RECT 8.6410 12.1365 8.7690 13.2300 ;
      RECT 8.6270 12.8020 8.7690 13.1245 ;
      RECT 8.4790 12.5290 8.5410 13.2300 ;
      RECT 8.4650 12.8385 8.5410 12.9920 ;
      RECT 8.4790 12.1365 8.5050 13.2300 ;
      RECT 8.4790 12.2575 8.5190 12.4970 ;
      RECT 8.4790 12.1365 8.5410 12.2255 ;
      RECT 8.1820 12.5870 8.3880 13.2300 ;
      RECT 8.3620 12.1365 8.3880 13.2300 ;
      RECT 8.1820 12.8640 8.4020 13.1220 ;
      RECT 8.1820 12.1365 8.2800 13.2300 ;
      RECT 7.7650 12.1365 7.8480 13.2300 ;
      RECT 7.7650 12.2250 7.8620 13.1605 ;
      RECT 16.4440 12.1365 16.5290 13.2300 ;
      RECT 16.3000 12.1365 16.3260 13.2300 ;
      RECT 16.1920 12.1365 16.2180 13.2300 ;
      RECT 16.0840 12.1365 16.1100 13.2300 ;
      RECT 15.9760 12.1365 16.0020 13.2300 ;
      RECT 15.8680 12.1365 15.8940 13.2300 ;
      RECT 15.7600 12.1365 15.7860 13.2300 ;
      RECT 15.6520 12.1365 15.6780 13.2300 ;
      RECT 15.5440 12.1365 15.5700 13.2300 ;
      RECT 15.4360 12.1365 15.4620 13.2300 ;
      RECT 15.3280 12.1365 15.3540 13.2300 ;
      RECT 15.2200 12.1365 15.2460 13.2300 ;
      RECT 15.1120 12.1365 15.1380 13.2300 ;
      RECT 15.0040 12.1365 15.0300 13.2300 ;
      RECT 14.8960 12.1365 14.9220 13.2300 ;
      RECT 14.7880 12.1365 14.8140 13.2300 ;
      RECT 14.6800 12.1365 14.7060 13.2300 ;
      RECT 14.5720 12.1365 14.5980 13.2300 ;
      RECT 14.4640 12.1365 14.4900 13.2300 ;
      RECT 14.3560 12.1365 14.3820 13.2300 ;
      RECT 14.2480 12.1365 14.2740 13.2300 ;
      RECT 14.1400 12.1365 14.1660 13.2300 ;
      RECT 14.0320 12.1365 14.0580 13.2300 ;
      RECT 13.9240 12.1365 13.9500 13.2300 ;
      RECT 13.8160 12.1365 13.8420 13.2300 ;
      RECT 13.7080 12.1365 13.7340 13.2300 ;
      RECT 13.6000 12.1365 13.6260 13.2300 ;
      RECT 13.4920 12.1365 13.5180 13.2300 ;
      RECT 13.3840 12.1365 13.4100 13.2300 ;
      RECT 13.2760 12.1365 13.3020 13.2300 ;
      RECT 13.1680 12.1365 13.1940 13.2300 ;
      RECT 13.0600 12.1365 13.0860 13.2300 ;
      RECT 12.9520 12.1365 12.9780 13.2300 ;
      RECT 12.8440 12.1365 12.8700 13.2300 ;
      RECT 12.7360 12.1365 12.7620 13.2300 ;
      RECT 12.6280 12.1365 12.6540 13.2300 ;
      RECT 12.5200 12.1365 12.5460 13.2300 ;
      RECT 12.4120 12.1365 12.4380 13.2300 ;
      RECT 12.3040 12.1365 12.3300 13.2300 ;
      RECT 12.1960 12.1365 12.2220 13.2300 ;
      RECT 12.0880 12.1365 12.1140 13.2300 ;
      RECT 11.9800 12.1365 12.0060 13.2300 ;
      RECT 11.8720 12.1365 11.8980 13.2300 ;
      RECT 11.7640 12.1365 11.7900 13.2300 ;
      RECT 11.6560 12.1365 11.6820 13.2300 ;
      RECT 11.5480 12.1365 11.5740 13.2300 ;
      RECT 11.4400 12.1365 11.4660 13.2300 ;
      RECT 11.3320 12.1365 11.3580 13.2300 ;
      RECT 11.2240 12.1365 11.2500 13.2300 ;
      RECT 11.1160 12.1365 11.1420 13.2300 ;
      RECT 11.0080 12.1365 11.0340 13.2300 ;
      RECT 10.9000 12.1365 10.9260 13.2300 ;
      RECT 10.7920 12.1365 10.8180 13.2300 ;
      RECT 10.6840 12.1365 10.7100 13.2300 ;
      RECT 10.5760 12.1365 10.6020 13.2300 ;
      RECT 10.4680 12.1365 10.4940 13.2300 ;
      RECT 10.3600 12.1365 10.3860 13.2300 ;
      RECT 10.2520 12.1365 10.2780 13.2300 ;
      RECT 10.1440 12.1365 10.1700 13.2300 ;
      RECT 10.0360 12.1365 10.0620 13.2300 ;
      RECT 9.9280 12.1365 9.9540 13.2300 ;
      RECT 9.8200 12.1365 9.8460 13.2300 ;
      RECT 9.7120 12.1365 9.7380 13.2300 ;
      RECT 9.6040 12.1365 9.6300 13.2300 ;
      RECT 9.4960 12.1365 9.5220 13.2300 ;
      RECT 9.3880 12.1365 9.4140 13.2300 ;
      RECT 9.1750 12.1365 9.2520 13.2300 ;
      RECT 7.2820 12.1365 7.3590 13.2300 ;
      RECT 7.1200 12.1365 7.1460 13.2300 ;
      RECT 7.0120 12.1365 7.0380 13.2300 ;
      RECT 6.9040 12.1365 6.9300 13.2300 ;
      RECT 6.7960 12.1365 6.8220 13.2300 ;
      RECT 6.6880 12.1365 6.7140 13.2300 ;
      RECT 6.5800 12.1365 6.6060 13.2300 ;
      RECT 6.4720 12.1365 6.4980 13.2300 ;
      RECT 6.3640 12.1365 6.3900 13.2300 ;
      RECT 6.2560 12.1365 6.2820 13.2300 ;
      RECT 6.1480 12.1365 6.1740 13.2300 ;
      RECT 6.0400 12.1365 6.0660 13.2300 ;
      RECT 5.9320 12.1365 5.9580 13.2300 ;
      RECT 5.8240 12.1365 5.8500 13.2300 ;
      RECT 5.7160 12.1365 5.7420 13.2300 ;
      RECT 5.6080 12.1365 5.6340 13.2300 ;
      RECT 5.5000 12.1365 5.5260 13.2300 ;
      RECT 5.3920 12.1365 5.4180 13.2300 ;
      RECT 5.2840 12.1365 5.3100 13.2300 ;
      RECT 5.1760 12.1365 5.2020 13.2300 ;
      RECT 5.0680 12.1365 5.0940 13.2300 ;
      RECT 4.9600 12.1365 4.9860 13.2300 ;
      RECT 4.8520 12.1365 4.8780 13.2300 ;
      RECT 4.7440 12.1365 4.7700 13.2300 ;
      RECT 4.6360 12.1365 4.6620 13.2300 ;
      RECT 4.5280 12.1365 4.5540 13.2300 ;
      RECT 4.4200 12.1365 4.4460 13.2300 ;
      RECT 4.3120 12.1365 4.3380 13.2300 ;
      RECT 4.2040 12.1365 4.2300 13.2300 ;
      RECT 4.0960 12.1365 4.1220 13.2300 ;
      RECT 3.9880 12.1365 4.0140 13.2300 ;
      RECT 3.8800 12.1365 3.9060 13.2300 ;
      RECT 3.7720 12.1365 3.7980 13.2300 ;
      RECT 3.6640 12.1365 3.6900 13.2300 ;
      RECT 3.5560 12.1365 3.5820 13.2300 ;
      RECT 3.4480 12.1365 3.4740 13.2300 ;
      RECT 3.3400 12.1365 3.3660 13.2300 ;
      RECT 3.2320 12.1365 3.2580 13.2300 ;
      RECT 3.1240 12.1365 3.1500 13.2300 ;
      RECT 3.0160 12.1365 3.0420 13.2300 ;
      RECT 2.9080 12.1365 2.9340 13.2300 ;
      RECT 2.8000 12.1365 2.8260 13.2300 ;
      RECT 2.6920 12.1365 2.7180 13.2300 ;
      RECT 2.5840 12.1365 2.6100 13.2300 ;
      RECT 2.4760 12.1365 2.5020 13.2300 ;
      RECT 2.3680 12.1365 2.3940 13.2300 ;
      RECT 2.2600 12.1365 2.2860 13.2300 ;
      RECT 2.1520 12.1365 2.1780 13.2300 ;
      RECT 2.0440 12.1365 2.0700 13.2300 ;
      RECT 1.9360 12.1365 1.9620 13.2300 ;
      RECT 1.8280 12.1365 1.8540 13.2300 ;
      RECT 1.7200 12.1365 1.7460 13.2300 ;
      RECT 1.6120 12.1365 1.6380 13.2300 ;
      RECT 1.5040 12.1365 1.5300 13.2300 ;
      RECT 1.3960 12.1365 1.4220 13.2300 ;
      RECT 1.2880 12.1365 1.3140 13.2300 ;
      RECT 1.1800 12.1365 1.2060 13.2300 ;
      RECT 1.0720 12.1365 1.0980 13.2300 ;
      RECT 0.9640 12.1365 0.9900 13.2300 ;
      RECT 0.8560 12.1365 0.8820 13.2300 ;
      RECT 0.7480 12.1365 0.7740 13.2300 ;
      RECT 0.6400 12.1365 0.6660 13.2300 ;
      RECT 0.5320 12.1365 0.5580 13.2300 ;
      RECT 0.4240 12.1365 0.4500 13.2300 ;
      RECT 0.3160 12.1365 0.3420 13.2300 ;
      RECT 0.2080 12.1365 0.2340 13.2300 ;
      RECT 0.0050 12.1365 0.0900 13.2300 ;
      RECT 8.6410 13.2165 8.7690 14.3100 ;
      RECT 8.6270 13.8820 8.7690 14.2045 ;
      RECT 8.4790 13.6090 8.5410 14.3100 ;
      RECT 8.4650 13.9185 8.5410 14.0720 ;
      RECT 8.4790 13.2165 8.5050 14.3100 ;
      RECT 8.4790 13.3375 8.5190 13.5770 ;
      RECT 8.4790 13.2165 8.5410 13.3055 ;
      RECT 8.1820 13.6670 8.3880 14.3100 ;
      RECT 8.3620 13.2165 8.3880 14.3100 ;
      RECT 8.1820 13.9440 8.4020 14.2020 ;
      RECT 8.1820 13.2165 8.2800 14.3100 ;
      RECT 7.7650 13.2165 7.8480 14.3100 ;
      RECT 7.7650 13.3050 7.8620 14.2405 ;
      RECT 16.4440 13.2165 16.5290 14.3100 ;
      RECT 16.3000 13.2165 16.3260 14.3100 ;
      RECT 16.1920 13.2165 16.2180 14.3100 ;
      RECT 16.0840 13.2165 16.1100 14.3100 ;
      RECT 15.9760 13.2165 16.0020 14.3100 ;
      RECT 15.8680 13.2165 15.8940 14.3100 ;
      RECT 15.7600 13.2165 15.7860 14.3100 ;
      RECT 15.6520 13.2165 15.6780 14.3100 ;
      RECT 15.5440 13.2165 15.5700 14.3100 ;
      RECT 15.4360 13.2165 15.4620 14.3100 ;
      RECT 15.3280 13.2165 15.3540 14.3100 ;
      RECT 15.2200 13.2165 15.2460 14.3100 ;
      RECT 15.1120 13.2165 15.1380 14.3100 ;
      RECT 15.0040 13.2165 15.0300 14.3100 ;
      RECT 14.8960 13.2165 14.9220 14.3100 ;
      RECT 14.7880 13.2165 14.8140 14.3100 ;
      RECT 14.6800 13.2165 14.7060 14.3100 ;
      RECT 14.5720 13.2165 14.5980 14.3100 ;
      RECT 14.4640 13.2165 14.4900 14.3100 ;
      RECT 14.3560 13.2165 14.3820 14.3100 ;
      RECT 14.2480 13.2165 14.2740 14.3100 ;
      RECT 14.1400 13.2165 14.1660 14.3100 ;
      RECT 14.0320 13.2165 14.0580 14.3100 ;
      RECT 13.9240 13.2165 13.9500 14.3100 ;
      RECT 13.8160 13.2165 13.8420 14.3100 ;
      RECT 13.7080 13.2165 13.7340 14.3100 ;
      RECT 13.6000 13.2165 13.6260 14.3100 ;
      RECT 13.4920 13.2165 13.5180 14.3100 ;
      RECT 13.3840 13.2165 13.4100 14.3100 ;
      RECT 13.2760 13.2165 13.3020 14.3100 ;
      RECT 13.1680 13.2165 13.1940 14.3100 ;
      RECT 13.0600 13.2165 13.0860 14.3100 ;
      RECT 12.9520 13.2165 12.9780 14.3100 ;
      RECT 12.8440 13.2165 12.8700 14.3100 ;
      RECT 12.7360 13.2165 12.7620 14.3100 ;
      RECT 12.6280 13.2165 12.6540 14.3100 ;
      RECT 12.5200 13.2165 12.5460 14.3100 ;
      RECT 12.4120 13.2165 12.4380 14.3100 ;
      RECT 12.3040 13.2165 12.3300 14.3100 ;
      RECT 12.1960 13.2165 12.2220 14.3100 ;
      RECT 12.0880 13.2165 12.1140 14.3100 ;
      RECT 11.9800 13.2165 12.0060 14.3100 ;
      RECT 11.8720 13.2165 11.8980 14.3100 ;
      RECT 11.7640 13.2165 11.7900 14.3100 ;
      RECT 11.6560 13.2165 11.6820 14.3100 ;
      RECT 11.5480 13.2165 11.5740 14.3100 ;
      RECT 11.4400 13.2165 11.4660 14.3100 ;
      RECT 11.3320 13.2165 11.3580 14.3100 ;
      RECT 11.2240 13.2165 11.2500 14.3100 ;
      RECT 11.1160 13.2165 11.1420 14.3100 ;
      RECT 11.0080 13.2165 11.0340 14.3100 ;
      RECT 10.9000 13.2165 10.9260 14.3100 ;
      RECT 10.7920 13.2165 10.8180 14.3100 ;
      RECT 10.6840 13.2165 10.7100 14.3100 ;
      RECT 10.5760 13.2165 10.6020 14.3100 ;
      RECT 10.4680 13.2165 10.4940 14.3100 ;
      RECT 10.3600 13.2165 10.3860 14.3100 ;
      RECT 10.2520 13.2165 10.2780 14.3100 ;
      RECT 10.1440 13.2165 10.1700 14.3100 ;
      RECT 10.0360 13.2165 10.0620 14.3100 ;
      RECT 9.9280 13.2165 9.9540 14.3100 ;
      RECT 9.8200 13.2165 9.8460 14.3100 ;
      RECT 9.7120 13.2165 9.7380 14.3100 ;
      RECT 9.6040 13.2165 9.6300 14.3100 ;
      RECT 9.4960 13.2165 9.5220 14.3100 ;
      RECT 9.3880 13.2165 9.4140 14.3100 ;
      RECT 9.1750 13.2165 9.2520 14.3100 ;
      RECT 7.2820 13.2165 7.3590 14.3100 ;
      RECT 7.1200 13.2165 7.1460 14.3100 ;
      RECT 7.0120 13.2165 7.0380 14.3100 ;
      RECT 6.9040 13.2165 6.9300 14.3100 ;
      RECT 6.7960 13.2165 6.8220 14.3100 ;
      RECT 6.6880 13.2165 6.7140 14.3100 ;
      RECT 6.5800 13.2165 6.6060 14.3100 ;
      RECT 6.4720 13.2165 6.4980 14.3100 ;
      RECT 6.3640 13.2165 6.3900 14.3100 ;
      RECT 6.2560 13.2165 6.2820 14.3100 ;
      RECT 6.1480 13.2165 6.1740 14.3100 ;
      RECT 6.0400 13.2165 6.0660 14.3100 ;
      RECT 5.9320 13.2165 5.9580 14.3100 ;
      RECT 5.8240 13.2165 5.8500 14.3100 ;
      RECT 5.7160 13.2165 5.7420 14.3100 ;
      RECT 5.6080 13.2165 5.6340 14.3100 ;
      RECT 5.5000 13.2165 5.5260 14.3100 ;
      RECT 5.3920 13.2165 5.4180 14.3100 ;
      RECT 5.2840 13.2165 5.3100 14.3100 ;
      RECT 5.1760 13.2165 5.2020 14.3100 ;
      RECT 5.0680 13.2165 5.0940 14.3100 ;
      RECT 4.9600 13.2165 4.9860 14.3100 ;
      RECT 4.8520 13.2165 4.8780 14.3100 ;
      RECT 4.7440 13.2165 4.7700 14.3100 ;
      RECT 4.6360 13.2165 4.6620 14.3100 ;
      RECT 4.5280 13.2165 4.5540 14.3100 ;
      RECT 4.4200 13.2165 4.4460 14.3100 ;
      RECT 4.3120 13.2165 4.3380 14.3100 ;
      RECT 4.2040 13.2165 4.2300 14.3100 ;
      RECT 4.0960 13.2165 4.1220 14.3100 ;
      RECT 3.9880 13.2165 4.0140 14.3100 ;
      RECT 3.8800 13.2165 3.9060 14.3100 ;
      RECT 3.7720 13.2165 3.7980 14.3100 ;
      RECT 3.6640 13.2165 3.6900 14.3100 ;
      RECT 3.5560 13.2165 3.5820 14.3100 ;
      RECT 3.4480 13.2165 3.4740 14.3100 ;
      RECT 3.3400 13.2165 3.3660 14.3100 ;
      RECT 3.2320 13.2165 3.2580 14.3100 ;
      RECT 3.1240 13.2165 3.1500 14.3100 ;
      RECT 3.0160 13.2165 3.0420 14.3100 ;
      RECT 2.9080 13.2165 2.9340 14.3100 ;
      RECT 2.8000 13.2165 2.8260 14.3100 ;
      RECT 2.6920 13.2165 2.7180 14.3100 ;
      RECT 2.5840 13.2165 2.6100 14.3100 ;
      RECT 2.4760 13.2165 2.5020 14.3100 ;
      RECT 2.3680 13.2165 2.3940 14.3100 ;
      RECT 2.2600 13.2165 2.2860 14.3100 ;
      RECT 2.1520 13.2165 2.1780 14.3100 ;
      RECT 2.0440 13.2165 2.0700 14.3100 ;
      RECT 1.9360 13.2165 1.9620 14.3100 ;
      RECT 1.8280 13.2165 1.8540 14.3100 ;
      RECT 1.7200 13.2165 1.7460 14.3100 ;
      RECT 1.6120 13.2165 1.6380 14.3100 ;
      RECT 1.5040 13.2165 1.5300 14.3100 ;
      RECT 1.3960 13.2165 1.4220 14.3100 ;
      RECT 1.2880 13.2165 1.3140 14.3100 ;
      RECT 1.1800 13.2165 1.2060 14.3100 ;
      RECT 1.0720 13.2165 1.0980 14.3100 ;
      RECT 0.9640 13.2165 0.9900 14.3100 ;
      RECT 0.8560 13.2165 0.8820 14.3100 ;
      RECT 0.7480 13.2165 0.7740 14.3100 ;
      RECT 0.6400 13.2165 0.6660 14.3100 ;
      RECT 0.5320 13.2165 0.5580 14.3100 ;
      RECT 0.4240 13.2165 0.4500 14.3100 ;
      RECT 0.3160 13.2165 0.3420 14.3100 ;
      RECT 0.2080 13.2165 0.2340 14.3100 ;
      RECT 0.0050 13.2165 0.0900 14.3100 ;
      RECT 8.6410 14.2965 8.7690 15.3900 ;
      RECT 8.6270 14.9620 8.7690 15.2845 ;
      RECT 8.4790 14.6890 8.5410 15.3900 ;
      RECT 8.4650 14.9985 8.5410 15.1520 ;
      RECT 8.4790 14.2965 8.5050 15.3900 ;
      RECT 8.4790 14.4175 8.5190 14.6570 ;
      RECT 8.4790 14.2965 8.5410 14.3855 ;
      RECT 8.1820 14.7470 8.3880 15.3900 ;
      RECT 8.3620 14.2965 8.3880 15.3900 ;
      RECT 8.1820 15.0240 8.4020 15.2820 ;
      RECT 8.1820 14.2965 8.2800 15.3900 ;
      RECT 7.7650 14.2965 7.8480 15.3900 ;
      RECT 7.7650 14.3850 7.8620 15.3205 ;
      RECT 16.4440 14.2965 16.5290 15.3900 ;
      RECT 16.3000 14.2965 16.3260 15.3900 ;
      RECT 16.1920 14.2965 16.2180 15.3900 ;
      RECT 16.0840 14.2965 16.1100 15.3900 ;
      RECT 15.9760 14.2965 16.0020 15.3900 ;
      RECT 15.8680 14.2965 15.8940 15.3900 ;
      RECT 15.7600 14.2965 15.7860 15.3900 ;
      RECT 15.6520 14.2965 15.6780 15.3900 ;
      RECT 15.5440 14.2965 15.5700 15.3900 ;
      RECT 15.4360 14.2965 15.4620 15.3900 ;
      RECT 15.3280 14.2965 15.3540 15.3900 ;
      RECT 15.2200 14.2965 15.2460 15.3900 ;
      RECT 15.1120 14.2965 15.1380 15.3900 ;
      RECT 15.0040 14.2965 15.0300 15.3900 ;
      RECT 14.8960 14.2965 14.9220 15.3900 ;
      RECT 14.7880 14.2965 14.8140 15.3900 ;
      RECT 14.6800 14.2965 14.7060 15.3900 ;
      RECT 14.5720 14.2965 14.5980 15.3900 ;
      RECT 14.4640 14.2965 14.4900 15.3900 ;
      RECT 14.3560 14.2965 14.3820 15.3900 ;
      RECT 14.2480 14.2965 14.2740 15.3900 ;
      RECT 14.1400 14.2965 14.1660 15.3900 ;
      RECT 14.0320 14.2965 14.0580 15.3900 ;
      RECT 13.9240 14.2965 13.9500 15.3900 ;
      RECT 13.8160 14.2965 13.8420 15.3900 ;
      RECT 13.7080 14.2965 13.7340 15.3900 ;
      RECT 13.6000 14.2965 13.6260 15.3900 ;
      RECT 13.4920 14.2965 13.5180 15.3900 ;
      RECT 13.3840 14.2965 13.4100 15.3900 ;
      RECT 13.2760 14.2965 13.3020 15.3900 ;
      RECT 13.1680 14.2965 13.1940 15.3900 ;
      RECT 13.0600 14.2965 13.0860 15.3900 ;
      RECT 12.9520 14.2965 12.9780 15.3900 ;
      RECT 12.8440 14.2965 12.8700 15.3900 ;
      RECT 12.7360 14.2965 12.7620 15.3900 ;
      RECT 12.6280 14.2965 12.6540 15.3900 ;
      RECT 12.5200 14.2965 12.5460 15.3900 ;
      RECT 12.4120 14.2965 12.4380 15.3900 ;
      RECT 12.3040 14.2965 12.3300 15.3900 ;
      RECT 12.1960 14.2965 12.2220 15.3900 ;
      RECT 12.0880 14.2965 12.1140 15.3900 ;
      RECT 11.9800 14.2965 12.0060 15.3900 ;
      RECT 11.8720 14.2965 11.8980 15.3900 ;
      RECT 11.7640 14.2965 11.7900 15.3900 ;
      RECT 11.6560 14.2965 11.6820 15.3900 ;
      RECT 11.5480 14.2965 11.5740 15.3900 ;
      RECT 11.4400 14.2965 11.4660 15.3900 ;
      RECT 11.3320 14.2965 11.3580 15.3900 ;
      RECT 11.2240 14.2965 11.2500 15.3900 ;
      RECT 11.1160 14.2965 11.1420 15.3900 ;
      RECT 11.0080 14.2965 11.0340 15.3900 ;
      RECT 10.9000 14.2965 10.9260 15.3900 ;
      RECT 10.7920 14.2965 10.8180 15.3900 ;
      RECT 10.6840 14.2965 10.7100 15.3900 ;
      RECT 10.5760 14.2965 10.6020 15.3900 ;
      RECT 10.4680 14.2965 10.4940 15.3900 ;
      RECT 10.3600 14.2965 10.3860 15.3900 ;
      RECT 10.2520 14.2965 10.2780 15.3900 ;
      RECT 10.1440 14.2965 10.1700 15.3900 ;
      RECT 10.0360 14.2965 10.0620 15.3900 ;
      RECT 9.9280 14.2965 9.9540 15.3900 ;
      RECT 9.8200 14.2965 9.8460 15.3900 ;
      RECT 9.7120 14.2965 9.7380 15.3900 ;
      RECT 9.6040 14.2965 9.6300 15.3900 ;
      RECT 9.4960 14.2965 9.5220 15.3900 ;
      RECT 9.3880 14.2965 9.4140 15.3900 ;
      RECT 9.1750 14.2965 9.2520 15.3900 ;
      RECT 7.2820 14.2965 7.3590 15.3900 ;
      RECT 7.1200 14.2965 7.1460 15.3900 ;
      RECT 7.0120 14.2965 7.0380 15.3900 ;
      RECT 6.9040 14.2965 6.9300 15.3900 ;
      RECT 6.7960 14.2965 6.8220 15.3900 ;
      RECT 6.6880 14.2965 6.7140 15.3900 ;
      RECT 6.5800 14.2965 6.6060 15.3900 ;
      RECT 6.4720 14.2965 6.4980 15.3900 ;
      RECT 6.3640 14.2965 6.3900 15.3900 ;
      RECT 6.2560 14.2965 6.2820 15.3900 ;
      RECT 6.1480 14.2965 6.1740 15.3900 ;
      RECT 6.0400 14.2965 6.0660 15.3900 ;
      RECT 5.9320 14.2965 5.9580 15.3900 ;
      RECT 5.8240 14.2965 5.8500 15.3900 ;
      RECT 5.7160 14.2965 5.7420 15.3900 ;
      RECT 5.6080 14.2965 5.6340 15.3900 ;
      RECT 5.5000 14.2965 5.5260 15.3900 ;
      RECT 5.3920 14.2965 5.4180 15.3900 ;
      RECT 5.2840 14.2965 5.3100 15.3900 ;
      RECT 5.1760 14.2965 5.2020 15.3900 ;
      RECT 5.0680 14.2965 5.0940 15.3900 ;
      RECT 4.9600 14.2965 4.9860 15.3900 ;
      RECT 4.8520 14.2965 4.8780 15.3900 ;
      RECT 4.7440 14.2965 4.7700 15.3900 ;
      RECT 4.6360 14.2965 4.6620 15.3900 ;
      RECT 4.5280 14.2965 4.5540 15.3900 ;
      RECT 4.4200 14.2965 4.4460 15.3900 ;
      RECT 4.3120 14.2965 4.3380 15.3900 ;
      RECT 4.2040 14.2965 4.2300 15.3900 ;
      RECT 4.0960 14.2965 4.1220 15.3900 ;
      RECT 3.9880 14.2965 4.0140 15.3900 ;
      RECT 3.8800 14.2965 3.9060 15.3900 ;
      RECT 3.7720 14.2965 3.7980 15.3900 ;
      RECT 3.6640 14.2965 3.6900 15.3900 ;
      RECT 3.5560 14.2965 3.5820 15.3900 ;
      RECT 3.4480 14.2965 3.4740 15.3900 ;
      RECT 3.3400 14.2965 3.3660 15.3900 ;
      RECT 3.2320 14.2965 3.2580 15.3900 ;
      RECT 3.1240 14.2965 3.1500 15.3900 ;
      RECT 3.0160 14.2965 3.0420 15.3900 ;
      RECT 2.9080 14.2965 2.9340 15.3900 ;
      RECT 2.8000 14.2965 2.8260 15.3900 ;
      RECT 2.6920 14.2965 2.7180 15.3900 ;
      RECT 2.5840 14.2965 2.6100 15.3900 ;
      RECT 2.4760 14.2965 2.5020 15.3900 ;
      RECT 2.3680 14.2965 2.3940 15.3900 ;
      RECT 2.2600 14.2965 2.2860 15.3900 ;
      RECT 2.1520 14.2965 2.1780 15.3900 ;
      RECT 2.0440 14.2965 2.0700 15.3900 ;
      RECT 1.9360 14.2965 1.9620 15.3900 ;
      RECT 1.8280 14.2965 1.8540 15.3900 ;
      RECT 1.7200 14.2965 1.7460 15.3900 ;
      RECT 1.6120 14.2965 1.6380 15.3900 ;
      RECT 1.5040 14.2965 1.5300 15.3900 ;
      RECT 1.3960 14.2965 1.4220 15.3900 ;
      RECT 1.2880 14.2965 1.3140 15.3900 ;
      RECT 1.1800 14.2965 1.2060 15.3900 ;
      RECT 1.0720 14.2965 1.0980 15.3900 ;
      RECT 0.9640 14.2965 0.9900 15.3900 ;
      RECT 0.8560 14.2965 0.8820 15.3900 ;
      RECT 0.7480 14.2965 0.7740 15.3900 ;
      RECT 0.6400 14.2965 0.6660 15.3900 ;
      RECT 0.5320 14.2965 0.5580 15.3900 ;
      RECT 0.4240 14.2965 0.4500 15.3900 ;
      RECT 0.3160 14.2965 0.3420 15.3900 ;
      RECT 0.2080 14.2965 0.2340 15.3900 ;
      RECT 0.0050 14.2965 0.0900 15.3900 ;
      RECT 8.6410 15.3765 8.7690 16.4700 ;
      RECT 8.6270 16.0420 8.7690 16.3645 ;
      RECT 8.4790 15.7690 8.5410 16.4700 ;
      RECT 8.4650 16.0785 8.5410 16.2320 ;
      RECT 8.4790 15.3765 8.5050 16.4700 ;
      RECT 8.4790 15.4975 8.5190 15.7370 ;
      RECT 8.4790 15.3765 8.5410 15.4655 ;
      RECT 8.1820 15.8270 8.3880 16.4700 ;
      RECT 8.3620 15.3765 8.3880 16.4700 ;
      RECT 8.1820 16.1040 8.4020 16.3620 ;
      RECT 8.1820 15.3765 8.2800 16.4700 ;
      RECT 7.7650 15.3765 7.8480 16.4700 ;
      RECT 7.7650 15.4650 7.8620 16.4005 ;
      RECT 16.4440 15.3765 16.5290 16.4700 ;
      RECT 16.3000 15.3765 16.3260 16.4700 ;
      RECT 16.1920 15.3765 16.2180 16.4700 ;
      RECT 16.0840 15.3765 16.1100 16.4700 ;
      RECT 15.9760 15.3765 16.0020 16.4700 ;
      RECT 15.8680 15.3765 15.8940 16.4700 ;
      RECT 15.7600 15.3765 15.7860 16.4700 ;
      RECT 15.6520 15.3765 15.6780 16.4700 ;
      RECT 15.5440 15.3765 15.5700 16.4700 ;
      RECT 15.4360 15.3765 15.4620 16.4700 ;
      RECT 15.3280 15.3765 15.3540 16.4700 ;
      RECT 15.2200 15.3765 15.2460 16.4700 ;
      RECT 15.1120 15.3765 15.1380 16.4700 ;
      RECT 15.0040 15.3765 15.0300 16.4700 ;
      RECT 14.8960 15.3765 14.9220 16.4700 ;
      RECT 14.7880 15.3765 14.8140 16.4700 ;
      RECT 14.6800 15.3765 14.7060 16.4700 ;
      RECT 14.5720 15.3765 14.5980 16.4700 ;
      RECT 14.4640 15.3765 14.4900 16.4700 ;
      RECT 14.3560 15.3765 14.3820 16.4700 ;
      RECT 14.2480 15.3765 14.2740 16.4700 ;
      RECT 14.1400 15.3765 14.1660 16.4700 ;
      RECT 14.0320 15.3765 14.0580 16.4700 ;
      RECT 13.9240 15.3765 13.9500 16.4700 ;
      RECT 13.8160 15.3765 13.8420 16.4700 ;
      RECT 13.7080 15.3765 13.7340 16.4700 ;
      RECT 13.6000 15.3765 13.6260 16.4700 ;
      RECT 13.4920 15.3765 13.5180 16.4700 ;
      RECT 13.3840 15.3765 13.4100 16.4700 ;
      RECT 13.2760 15.3765 13.3020 16.4700 ;
      RECT 13.1680 15.3765 13.1940 16.4700 ;
      RECT 13.0600 15.3765 13.0860 16.4700 ;
      RECT 12.9520 15.3765 12.9780 16.4700 ;
      RECT 12.8440 15.3765 12.8700 16.4700 ;
      RECT 12.7360 15.3765 12.7620 16.4700 ;
      RECT 12.6280 15.3765 12.6540 16.4700 ;
      RECT 12.5200 15.3765 12.5460 16.4700 ;
      RECT 12.4120 15.3765 12.4380 16.4700 ;
      RECT 12.3040 15.3765 12.3300 16.4700 ;
      RECT 12.1960 15.3765 12.2220 16.4700 ;
      RECT 12.0880 15.3765 12.1140 16.4700 ;
      RECT 11.9800 15.3765 12.0060 16.4700 ;
      RECT 11.8720 15.3765 11.8980 16.4700 ;
      RECT 11.7640 15.3765 11.7900 16.4700 ;
      RECT 11.6560 15.3765 11.6820 16.4700 ;
      RECT 11.5480 15.3765 11.5740 16.4700 ;
      RECT 11.4400 15.3765 11.4660 16.4700 ;
      RECT 11.3320 15.3765 11.3580 16.4700 ;
      RECT 11.2240 15.3765 11.2500 16.4700 ;
      RECT 11.1160 15.3765 11.1420 16.4700 ;
      RECT 11.0080 15.3765 11.0340 16.4700 ;
      RECT 10.9000 15.3765 10.9260 16.4700 ;
      RECT 10.7920 15.3765 10.8180 16.4700 ;
      RECT 10.6840 15.3765 10.7100 16.4700 ;
      RECT 10.5760 15.3765 10.6020 16.4700 ;
      RECT 10.4680 15.3765 10.4940 16.4700 ;
      RECT 10.3600 15.3765 10.3860 16.4700 ;
      RECT 10.2520 15.3765 10.2780 16.4700 ;
      RECT 10.1440 15.3765 10.1700 16.4700 ;
      RECT 10.0360 15.3765 10.0620 16.4700 ;
      RECT 9.9280 15.3765 9.9540 16.4700 ;
      RECT 9.8200 15.3765 9.8460 16.4700 ;
      RECT 9.7120 15.3765 9.7380 16.4700 ;
      RECT 9.6040 15.3765 9.6300 16.4700 ;
      RECT 9.4960 15.3765 9.5220 16.4700 ;
      RECT 9.3880 15.3765 9.4140 16.4700 ;
      RECT 9.1750 15.3765 9.2520 16.4700 ;
      RECT 7.2820 15.3765 7.3590 16.4700 ;
      RECT 7.1200 15.3765 7.1460 16.4700 ;
      RECT 7.0120 15.3765 7.0380 16.4700 ;
      RECT 6.9040 15.3765 6.9300 16.4700 ;
      RECT 6.7960 15.3765 6.8220 16.4700 ;
      RECT 6.6880 15.3765 6.7140 16.4700 ;
      RECT 6.5800 15.3765 6.6060 16.4700 ;
      RECT 6.4720 15.3765 6.4980 16.4700 ;
      RECT 6.3640 15.3765 6.3900 16.4700 ;
      RECT 6.2560 15.3765 6.2820 16.4700 ;
      RECT 6.1480 15.3765 6.1740 16.4700 ;
      RECT 6.0400 15.3765 6.0660 16.4700 ;
      RECT 5.9320 15.3765 5.9580 16.4700 ;
      RECT 5.8240 15.3765 5.8500 16.4700 ;
      RECT 5.7160 15.3765 5.7420 16.4700 ;
      RECT 5.6080 15.3765 5.6340 16.4700 ;
      RECT 5.5000 15.3765 5.5260 16.4700 ;
      RECT 5.3920 15.3765 5.4180 16.4700 ;
      RECT 5.2840 15.3765 5.3100 16.4700 ;
      RECT 5.1760 15.3765 5.2020 16.4700 ;
      RECT 5.0680 15.3765 5.0940 16.4700 ;
      RECT 4.9600 15.3765 4.9860 16.4700 ;
      RECT 4.8520 15.3765 4.8780 16.4700 ;
      RECT 4.7440 15.3765 4.7700 16.4700 ;
      RECT 4.6360 15.3765 4.6620 16.4700 ;
      RECT 4.5280 15.3765 4.5540 16.4700 ;
      RECT 4.4200 15.3765 4.4460 16.4700 ;
      RECT 4.3120 15.3765 4.3380 16.4700 ;
      RECT 4.2040 15.3765 4.2300 16.4700 ;
      RECT 4.0960 15.3765 4.1220 16.4700 ;
      RECT 3.9880 15.3765 4.0140 16.4700 ;
      RECT 3.8800 15.3765 3.9060 16.4700 ;
      RECT 3.7720 15.3765 3.7980 16.4700 ;
      RECT 3.6640 15.3765 3.6900 16.4700 ;
      RECT 3.5560 15.3765 3.5820 16.4700 ;
      RECT 3.4480 15.3765 3.4740 16.4700 ;
      RECT 3.3400 15.3765 3.3660 16.4700 ;
      RECT 3.2320 15.3765 3.2580 16.4700 ;
      RECT 3.1240 15.3765 3.1500 16.4700 ;
      RECT 3.0160 15.3765 3.0420 16.4700 ;
      RECT 2.9080 15.3765 2.9340 16.4700 ;
      RECT 2.8000 15.3765 2.8260 16.4700 ;
      RECT 2.6920 15.3765 2.7180 16.4700 ;
      RECT 2.5840 15.3765 2.6100 16.4700 ;
      RECT 2.4760 15.3765 2.5020 16.4700 ;
      RECT 2.3680 15.3765 2.3940 16.4700 ;
      RECT 2.2600 15.3765 2.2860 16.4700 ;
      RECT 2.1520 15.3765 2.1780 16.4700 ;
      RECT 2.0440 15.3765 2.0700 16.4700 ;
      RECT 1.9360 15.3765 1.9620 16.4700 ;
      RECT 1.8280 15.3765 1.8540 16.4700 ;
      RECT 1.7200 15.3765 1.7460 16.4700 ;
      RECT 1.6120 15.3765 1.6380 16.4700 ;
      RECT 1.5040 15.3765 1.5300 16.4700 ;
      RECT 1.3960 15.3765 1.4220 16.4700 ;
      RECT 1.2880 15.3765 1.3140 16.4700 ;
      RECT 1.1800 15.3765 1.2060 16.4700 ;
      RECT 1.0720 15.3765 1.0980 16.4700 ;
      RECT 0.9640 15.3765 0.9900 16.4700 ;
      RECT 0.8560 15.3765 0.8820 16.4700 ;
      RECT 0.7480 15.3765 0.7740 16.4700 ;
      RECT 0.6400 15.3765 0.6660 16.4700 ;
      RECT 0.5320 15.3765 0.5580 16.4700 ;
      RECT 0.4240 15.3765 0.4500 16.4700 ;
      RECT 0.3160 15.3765 0.3420 16.4700 ;
      RECT 0.2080 15.3765 0.2340 16.4700 ;
      RECT 0.0050 15.3765 0.0900 16.4700 ;
      RECT 8.6410 16.4565 8.7690 17.5500 ;
      RECT 8.6270 17.1220 8.7690 17.4445 ;
      RECT 8.4790 16.8490 8.5410 17.5500 ;
      RECT 8.4650 17.1585 8.5410 17.3120 ;
      RECT 8.4790 16.4565 8.5050 17.5500 ;
      RECT 8.4790 16.5775 8.5190 16.8170 ;
      RECT 8.4790 16.4565 8.5410 16.5455 ;
      RECT 8.1820 16.9070 8.3880 17.5500 ;
      RECT 8.3620 16.4565 8.3880 17.5500 ;
      RECT 8.1820 17.1840 8.4020 17.4420 ;
      RECT 8.1820 16.4565 8.2800 17.5500 ;
      RECT 7.7650 16.4565 7.8480 17.5500 ;
      RECT 7.7650 16.5450 7.8620 17.4805 ;
      RECT 16.4440 16.4565 16.5290 17.5500 ;
      RECT 16.3000 16.4565 16.3260 17.5500 ;
      RECT 16.1920 16.4565 16.2180 17.5500 ;
      RECT 16.0840 16.4565 16.1100 17.5500 ;
      RECT 15.9760 16.4565 16.0020 17.5500 ;
      RECT 15.8680 16.4565 15.8940 17.5500 ;
      RECT 15.7600 16.4565 15.7860 17.5500 ;
      RECT 15.6520 16.4565 15.6780 17.5500 ;
      RECT 15.5440 16.4565 15.5700 17.5500 ;
      RECT 15.4360 16.4565 15.4620 17.5500 ;
      RECT 15.3280 16.4565 15.3540 17.5500 ;
      RECT 15.2200 16.4565 15.2460 17.5500 ;
      RECT 15.1120 16.4565 15.1380 17.5500 ;
      RECT 15.0040 16.4565 15.0300 17.5500 ;
      RECT 14.8960 16.4565 14.9220 17.5500 ;
      RECT 14.7880 16.4565 14.8140 17.5500 ;
      RECT 14.6800 16.4565 14.7060 17.5500 ;
      RECT 14.5720 16.4565 14.5980 17.5500 ;
      RECT 14.4640 16.4565 14.4900 17.5500 ;
      RECT 14.3560 16.4565 14.3820 17.5500 ;
      RECT 14.2480 16.4565 14.2740 17.5500 ;
      RECT 14.1400 16.4565 14.1660 17.5500 ;
      RECT 14.0320 16.4565 14.0580 17.5500 ;
      RECT 13.9240 16.4565 13.9500 17.5500 ;
      RECT 13.8160 16.4565 13.8420 17.5500 ;
      RECT 13.7080 16.4565 13.7340 17.5500 ;
      RECT 13.6000 16.4565 13.6260 17.5500 ;
      RECT 13.4920 16.4565 13.5180 17.5500 ;
      RECT 13.3840 16.4565 13.4100 17.5500 ;
      RECT 13.2760 16.4565 13.3020 17.5500 ;
      RECT 13.1680 16.4565 13.1940 17.5500 ;
      RECT 13.0600 16.4565 13.0860 17.5500 ;
      RECT 12.9520 16.4565 12.9780 17.5500 ;
      RECT 12.8440 16.4565 12.8700 17.5500 ;
      RECT 12.7360 16.4565 12.7620 17.5500 ;
      RECT 12.6280 16.4565 12.6540 17.5500 ;
      RECT 12.5200 16.4565 12.5460 17.5500 ;
      RECT 12.4120 16.4565 12.4380 17.5500 ;
      RECT 12.3040 16.4565 12.3300 17.5500 ;
      RECT 12.1960 16.4565 12.2220 17.5500 ;
      RECT 12.0880 16.4565 12.1140 17.5500 ;
      RECT 11.9800 16.4565 12.0060 17.5500 ;
      RECT 11.8720 16.4565 11.8980 17.5500 ;
      RECT 11.7640 16.4565 11.7900 17.5500 ;
      RECT 11.6560 16.4565 11.6820 17.5500 ;
      RECT 11.5480 16.4565 11.5740 17.5500 ;
      RECT 11.4400 16.4565 11.4660 17.5500 ;
      RECT 11.3320 16.4565 11.3580 17.5500 ;
      RECT 11.2240 16.4565 11.2500 17.5500 ;
      RECT 11.1160 16.4565 11.1420 17.5500 ;
      RECT 11.0080 16.4565 11.0340 17.5500 ;
      RECT 10.9000 16.4565 10.9260 17.5500 ;
      RECT 10.7920 16.4565 10.8180 17.5500 ;
      RECT 10.6840 16.4565 10.7100 17.5500 ;
      RECT 10.5760 16.4565 10.6020 17.5500 ;
      RECT 10.4680 16.4565 10.4940 17.5500 ;
      RECT 10.3600 16.4565 10.3860 17.5500 ;
      RECT 10.2520 16.4565 10.2780 17.5500 ;
      RECT 10.1440 16.4565 10.1700 17.5500 ;
      RECT 10.0360 16.4565 10.0620 17.5500 ;
      RECT 9.9280 16.4565 9.9540 17.5500 ;
      RECT 9.8200 16.4565 9.8460 17.5500 ;
      RECT 9.7120 16.4565 9.7380 17.5500 ;
      RECT 9.6040 16.4565 9.6300 17.5500 ;
      RECT 9.4960 16.4565 9.5220 17.5500 ;
      RECT 9.3880 16.4565 9.4140 17.5500 ;
      RECT 9.1750 16.4565 9.2520 17.5500 ;
      RECT 7.2820 16.4565 7.3590 17.5500 ;
      RECT 7.1200 16.4565 7.1460 17.5500 ;
      RECT 7.0120 16.4565 7.0380 17.5500 ;
      RECT 6.9040 16.4565 6.9300 17.5500 ;
      RECT 6.7960 16.4565 6.8220 17.5500 ;
      RECT 6.6880 16.4565 6.7140 17.5500 ;
      RECT 6.5800 16.4565 6.6060 17.5500 ;
      RECT 6.4720 16.4565 6.4980 17.5500 ;
      RECT 6.3640 16.4565 6.3900 17.5500 ;
      RECT 6.2560 16.4565 6.2820 17.5500 ;
      RECT 6.1480 16.4565 6.1740 17.5500 ;
      RECT 6.0400 16.4565 6.0660 17.5500 ;
      RECT 5.9320 16.4565 5.9580 17.5500 ;
      RECT 5.8240 16.4565 5.8500 17.5500 ;
      RECT 5.7160 16.4565 5.7420 17.5500 ;
      RECT 5.6080 16.4565 5.6340 17.5500 ;
      RECT 5.5000 16.4565 5.5260 17.5500 ;
      RECT 5.3920 16.4565 5.4180 17.5500 ;
      RECT 5.2840 16.4565 5.3100 17.5500 ;
      RECT 5.1760 16.4565 5.2020 17.5500 ;
      RECT 5.0680 16.4565 5.0940 17.5500 ;
      RECT 4.9600 16.4565 4.9860 17.5500 ;
      RECT 4.8520 16.4565 4.8780 17.5500 ;
      RECT 4.7440 16.4565 4.7700 17.5500 ;
      RECT 4.6360 16.4565 4.6620 17.5500 ;
      RECT 4.5280 16.4565 4.5540 17.5500 ;
      RECT 4.4200 16.4565 4.4460 17.5500 ;
      RECT 4.3120 16.4565 4.3380 17.5500 ;
      RECT 4.2040 16.4565 4.2300 17.5500 ;
      RECT 4.0960 16.4565 4.1220 17.5500 ;
      RECT 3.9880 16.4565 4.0140 17.5500 ;
      RECT 3.8800 16.4565 3.9060 17.5500 ;
      RECT 3.7720 16.4565 3.7980 17.5500 ;
      RECT 3.6640 16.4565 3.6900 17.5500 ;
      RECT 3.5560 16.4565 3.5820 17.5500 ;
      RECT 3.4480 16.4565 3.4740 17.5500 ;
      RECT 3.3400 16.4565 3.3660 17.5500 ;
      RECT 3.2320 16.4565 3.2580 17.5500 ;
      RECT 3.1240 16.4565 3.1500 17.5500 ;
      RECT 3.0160 16.4565 3.0420 17.5500 ;
      RECT 2.9080 16.4565 2.9340 17.5500 ;
      RECT 2.8000 16.4565 2.8260 17.5500 ;
      RECT 2.6920 16.4565 2.7180 17.5500 ;
      RECT 2.5840 16.4565 2.6100 17.5500 ;
      RECT 2.4760 16.4565 2.5020 17.5500 ;
      RECT 2.3680 16.4565 2.3940 17.5500 ;
      RECT 2.2600 16.4565 2.2860 17.5500 ;
      RECT 2.1520 16.4565 2.1780 17.5500 ;
      RECT 2.0440 16.4565 2.0700 17.5500 ;
      RECT 1.9360 16.4565 1.9620 17.5500 ;
      RECT 1.8280 16.4565 1.8540 17.5500 ;
      RECT 1.7200 16.4565 1.7460 17.5500 ;
      RECT 1.6120 16.4565 1.6380 17.5500 ;
      RECT 1.5040 16.4565 1.5300 17.5500 ;
      RECT 1.3960 16.4565 1.4220 17.5500 ;
      RECT 1.2880 16.4565 1.3140 17.5500 ;
      RECT 1.1800 16.4565 1.2060 17.5500 ;
      RECT 1.0720 16.4565 1.0980 17.5500 ;
      RECT 0.9640 16.4565 0.9900 17.5500 ;
      RECT 0.8560 16.4565 0.8820 17.5500 ;
      RECT 0.7480 16.4565 0.7740 17.5500 ;
      RECT 0.6400 16.4565 0.6660 17.5500 ;
      RECT 0.5320 16.4565 0.5580 17.5500 ;
      RECT 0.4240 16.4565 0.4500 17.5500 ;
      RECT 0.3160 16.4565 0.3420 17.5500 ;
      RECT 0.2080 16.4565 0.2340 17.5500 ;
      RECT 0.0050 16.4565 0.0900 17.5500 ;
      RECT 8.6410 17.5365 8.7690 18.6300 ;
      RECT 8.6270 18.2020 8.7690 18.5245 ;
      RECT 8.4790 17.9290 8.5410 18.6300 ;
      RECT 8.4650 18.2385 8.5410 18.3920 ;
      RECT 8.4790 17.5365 8.5050 18.6300 ;
      RECT 8.4790 17.6575 8.5190 17.8970 ;
      RECT 8.4790 17.5365 8.5410 17.6255 ;
      RECT 8.1820 17.9870 8.3880 18.6300 ;
      RECT 8.3620 17.5365 8.3880 18.6300 ;
      RECT 8.1820 18.2640 8.4020 18.5220 ;
      RECT 8.1820 17.5365 8.2800 18.6300 ;
      RECT 7.7650 17.5365 7.8480 18.6300 ;
      RECT 7.7650 17.6250 7.8620 18.5605 ;
      RECT 16.4440 17.5365 16.5290 18.6300 ;
      RECT 16.3000 17.5365 16.3260 18.6300 ;
      RECT 16.1920 17.5365 16.2180 18.6300 ;
      RECT 16.0840 17.5365 16.1100 18.6300 ;
      RECT 15.9760 17.5365 16.0020 18.6300 ;
      RECT 15.8680 17.5365 15.8940 18.6300 ;
      RECT 15.7600 17.5365 15.7860 18.6300 ;
      RECT 15.6520 17.5365 15.6780 18.6300 ;
      RECT 15.5440 17.5365 15.5700 18.6300 ;
      RECT 15.4360 17.5365 15.4620 18.6300 ;
      RECT 15.3280 17.5365 15.3540 18.6300 ;
      RECT 15.2200 17.5365 15.2460 18.6300 ;
      RECT 15.1120 17.5365 15.1380 18.6300 ;
      RECT 15.0040 17.5365 15.0300 18.6300 ;
      RECT 14.8960 17.5365 14.9220 18.6300 ;
      RECT 14.7880 17.5365 14.8140 18.6300 ;
      RECT 14.6800 17.5365 14.7060 18.6300 ;
      RECT 14.5720 17.5365 14.5980 18.6300 ;
      RECT 14.4640 17.5365 14.4900 18.6300 ;
      RECT 14.3560 17.5365 14.3820 18.6300 ;
      RECT 14.2480 17.5365 14.2740 18.6300 ;
      RECT 14.1400 17.5365 14.1660 18.6300 ;
      RECT 14.0320 17.5365 14.0580 18.6300 ;
      RECT 13.9240 17.5365 13.9500 18.6300 ;
      RECT 13.8160 17.5365 13.8420 18.6300 ;
      RECT 13.7080 17.5365 13.7340 18.6300 ;
      RECT 13.6000 17.5365 13.6260 18.6300 ;
      RECT 13.4920 17.5365 13.5180 18.6300 ;
      RECT 13.3840 17.5365 13.4100 18.6300 ;
      RECT 13.2760 17.5365 13.3020 18.6300 ;
      RECT 13.1680 17.5365 13.1940 18.6300 ;
      RECT 13.0600 17.5365 13.0860 18.6300 ;
      RECT 12.9520 17.5365 12.9780 18.6300 ;
      RECT 12.8440 17.5365 12.8700 18.6300 ;
      RECT 12.7360 17.5365 12.7620 18.6300 ;
      RECT 12.6280 17.5365 12.6540 18.6300 ;
      RECT 12.5200 17.5365 12.5460 18.6300 ;
      RECT 12.4120 17.5365 12.4380 18.6300 ;
      RECT 12.3040 17.5365 12.3300 18.6300 ;
      RECT 12.1960 17.5365 12.2220 18.6300 ;
      RECT 12.0880 17.5365 12.1140 18.6300 ;
      RECT 11.9800 17.5365 12.0060 18.6300 ;
      RECT 11.8720 17.5365 11.8980 18.6300 ;
      RECT 11.7640 17.5365 11.7900 18.6300 ;
      RECT 11.6560 17.5365 11.6820 18.6300 ;
      RECT 11.5480 17.5365 11.5740 18.6300 ;
      RECT 11.4400 17.5365 11.4660 18.6300 ;
      RECT 11.3320 17.5365 11.3580 18.6300 ;
      RECT 11.2240 17.5365 11.2500 18.6300 ;
      RECT 11.1160 17.5365 11.1420 18.6300 ;
      RECT 11.0080 17.5365 11.0340 18.6300 ;
      RECT 10.9000 17.5365 10.9260 18.6300 ;
      RECT 10.7920 17.5365 10.8180 18.6300 ;
      RECT 10.6840 17.5365 10.7100 18.6300 ;
      RECT 10.5760 17.5365 10.6020 18.6300 ;
      RECT 10.4680 17.5365 10.4940 18.6300 ;
      RECT 10.3600 17.5365 10.3860 18.6300 ;
      RECT 10.2520 17.5365 10.2780 18.6300 ;
      RECT 10.1440 17.5365 10.1700 18.6300 ;
      RECT 10.0360 17.5365 10.0620 18.6300 ;
      RECT 9.9280 17.5365 9.9540 18.6300 ;
      RECT 9.8200 17.5365 9.8460 18.6300 ;
      RECT 9.7120 17.5365 9.7380 18.6300 ;
      RECT 9.6040 17.5365 9.6300 18.6300 ;
      RECT 9.4960 17.5365 9.5220 18.6300 ;
      RECT 9.3880 17.5365 9.4140 18.6300 ;
      RECT 9.1750 17.5365 9.2520 18.6300 ;
      RECT 7.2820 17.5365 7.3590 18.6300 ;
      RECT 7.1200 17.5365 7.1460 18.6300 ;
      RECT 7.0120 17.5365 7.0380 18.6300 ;
      RECT 6.9040 17.5365 6.9300 18.6300 ;
      RECT 6.7960 17.5365 6.8220 18.6300 ;
      RECT 6.6880 17.5365 6.7140 18.6300 ;
      RECT 6.5800 17.5365 6.6060 18.6300 ;
      RECT 6.4720 17.5365 6.4980 18.6300 ;
      RECT 6.3640 17.5365 6.3900 18.6300 ;
      RECT 6.2560 17.5365 6.2820 18.6300 ;
      RECT 6.1480 17.5365 6.1740 18.6300 ;
      RECT 6.0400 17.5365 6.0660 18.6300 ;
      RECT 5.9320 17.5365 5.9580 18.6300 ;
      RECT 5.8240 17.5365 5.8500 18.6300 ;
      RECT 5.7160 17.5365 5.7420 18.6300 ;
      RECT 5.6080 17.5365 5.6340 18.6300 ;
      RECT 5.5000 17.5365 5.5260 18.6300 ;
      RECT 5.3920 17.5365 5.4180 18.6300 ;
      RECT 5.2840 17.5365 5.3100 18.6300 ;
      RECT 5.1760 17.5365 5.2020 18.6300 ;
      RECT 5.0680 17.5365 5.0940 18.6300 ;
      RECT 4.9600 17.5365 4.9860 18.6300 ;
      RECT 4.8520 17.5365 4.8780 18.6300 ;
      RECT 4.7440 17.5365 4.7700 18.6300 ;
      RECT 4.6360 17.5365 4.6620 18.6300 ;
      RECT 4.5280 17.5365 4.5540 18.6300 ;
      RECT 4.4200 17.5365 4.4460 18.6300 ;
      RECT 4.3120 17.5365 4.3380 18.6300 ;
      RECT 4.2040 17.5365 4.2300 18.6300 ;
      RECT 4.0960 17.5365 4.1220 18.6300 ;
      RECT 3.9880 17.5365 4.0140 18.6300 ;
      RECT 3.8800 17.5365 3.9060 18.6300 ;
      RECT 3.7720 17.5365 3.7980 18.6300 ;
      RECT 3.6640 17.5365 3.6900 18.6300 ;
      RECT 3.5560 17.5365 3.5820 18.6300 ;
      RECT 3.4480 17.5365 3.4740 18.6300 ;
      RECT 3.3400 17.5365 3.3660 18.6300 ;
      RECT 3.2320 17.5365 3.2580 18.6300 ;
      RECT 3.1240 17.5365 3.1500 18.6300 ;
      RECT 3.0160 17.5365 3.0420 18.6300 ;
      RECT 2.9080 17.5365 2.9340 18.6300 ;
      RECT 2.8000 17.5365 2.8260 18.6300 ;
      RECT 2.6920 17.5365 2.7180 18.6300 ;
      RECT 2.5840 17.5365 2.6100 18.6300 ;
      RECT 2.4760 17.5365 2.5020 18.6300 ;
      RECT 2.3680 17.5365 2.3940 18.6300 ;
      RECT 2.2600 17.5365 2.2860 18.6300 ;
      RECT 2.1520 17.5365 2.1780 18.6300 ;
      RECT 2.0440 17.5365 2.0700 18.6300 ;
      RECT 1.9360 17.5365 1.9620 18.6300 ;
      RECT 1.8280 17.5365 1.8540 18.6300 ;
      RECT 1.7200 17.5365 1.7460 18.6300 ;
      RECT 1.6120 17.5365 1.6380 18.6300 ;
      RECT 1.5040 17.5365 1.5300 18.6300 ;
      RECT 1.3960 17.5365 1.4220 18.6300 ;
      RECT 1.2880 17.5365 1.3140 18.6300 ;
      RECT 1.1800 17.5365 1.2060 18.6300 ;
      RECT 1.0720 17.5365 1.0980 18.6300 ;
      RECT 0.9640 17.5365 0.9900 18.6300 ;
      RECT 0.8560 17.5365 0.8820 18.6300 ;
      RECT 0.7480 17.5365 0.7740 18.6300 ;
      RECT 0.6400 17.5365 0.6660 18.6300 ;
      RECT 0.5320 17.5365 0.5580 18.6300 ;
      RECT 0.4240 17.5365 0.4500 18.6300 ;
      RECT 0.3160 17.5365 0.3420 18.6300 ;
      RECT 0.2080 17.5365 0.2340 18.6300 ;
      RECT 0.0050 17.5365 0.0900 18.6300 ;
      RECT 8.6410 18.6165 8.7690 19.7100 ;
      RECT 8.6270 19.2820 8.7690 19.6045 ;
      RECT 8.4790 19.0090 8.5410 19.7100 ;
      RECT 8.4650 19.3185 8.5410 19.4720 ;
      RECT 8.4790 18.6165 8.5050 19.7100 ;
      RECT 8.4790 18.7375 8.5190 18.9770 ;
      RECT 8.4790 18.6165 8.5410 18.7055 ;
      RECT 8.1820 19.0670 8.3880 19.7100 ;
      RECT 8.3620 18.6165 8.3880 19.7100 ;
      RECT 8.1820 19.3440 8.4020 19.6020 ;
      RECT 8.1820 18.6165 8.2800 19.7100 ;
      RECT 7.7650 18.6165 7.8480 19.7100 ;
      RECT 7.7650 18.7050 7.8620 19.6405 ;
      RECT 16.4440 18.6165 16.5290 19.7100 ;
      RECT 16.3000 18.6165 16.3260 19.7100 ;
      RECT 16.1920 18.6165 16.2180 19.7100 ;
      RECT 16.0840 18.6165 16.1100 19.7100 ;
      RECT 15.9760 18.6165 16.0020 19.7100 ;
      RECT 15.8680 18.6165 15.8940 19.7100 ;
      RECT 15.7600 18.6165 15.7860 19.7100 ;
      RECT 15.6520 18.6165 15.6780 19.7100 ;
      RECT 15.5440 18.6165 15.5700 19.7100 ;
      RECT 15.4360 18.6165 15.4620 19.7100 ;
      RECT 15.3280 18.6165 15.3540 19.7100 ;
      RECT 15.2200 18.6165 15.2460 19.7100 ;
      RECT 15.1120 18.6165 15.1380 19.7100 ;
      RECT 15.0040 18.6165 15.0300 19.7100 ;
      RECT 14.8960 18.6165 14.9220 19.7100 ;
      RECT 14.7880 18.6165 14.8140 19.7100 ;
      RECT 14.6800 18.6165 14.7060 19.7100 ;
      RECT 14.5720 18.6165 14.5980 19.7100 ;
      RECT 14.4640 18.6165 14.4900 19.7100 ;
      RECT 14.3560 18.6165 14.3820 19.7100 ;
      RECT 14.2480 18.6165 14.2740 19.7100 ;
      RECT 14.1400 18.6165 14.1660 19.7100 ;
      RECT 14.0320 18.6165 14.0580 19.7100 ;
      RECT 13.9240 18.6165 13.9500 19.7100 ;
      RECT 13.8160 18.6165 13.8420 19.7100 ;
      RECT 13.7080 18.6165 13.7340 19.7100 ;
      RECT 13.6000 18.6165 13.6260 19.7100 ;
      RECT 13.4920 18.6165 13.5180 19.7100 ;
      RECT 13.3840 18.6165 13.4100 19.7100 ;
      RECT 13.2760 18.6165 13.3020 19.7100 ;
      RECT 13.1680 18.6165 13.1940 19.7100 ;
      RECT 13.0600 18.6165 13.0860 19.7100 ;
      RECT 12.9520 18.6165 12.9780 19.7100 ;
      RECT 12.8440 18.6165 12.8700 19.7100 ;
      RECT 12.7360 18.6165 12.7620 19.7100 ;
      RECT 12.6280 18.6165 12.6540 19.7100 ;
      RECT 12.5200 18.6165 12.5460 19.7100 ;
      RECT 12.4120 18.6165 12.4380 19.7100 ;
      RECT 12.3040 18.6165 12.3300 19.7100 ;
      RECT 12.1960 18.6165 12.2220 19.7100 ;
      RECT 12.0880 18.6165 12.1140 19.7100 ;
      RECT 11.9800 18.6165 12.0060 19.7100 ;
      RECT 11.8720 18.6165 11.8980 19.7100 ;
      RECT 11.7640 18.6165 11.7900 19.7100 ;
      RECT 11.6560 18.6165 11.6820 19.7100 ;
      RECT 11.5480 18.6165 11.5740 19.7100 ;
      RECT 11.4400 18.6165 11.4660 19.7100 ;
      RECT 11.3320 18.6165 11.3580 19.7100 ;
      RECT 11.2240 18.6165 11.2500 19.7100 ;
      RECT 11.1160 18.6165 11.1420 19.7100 ;
      RECT 11.0080 18.6165 11.0340 19.7100 ;
      RECT 10.9000 18.6165 10.9260 19.7100 ;
      RECT 10.7920 18.6165 10.8180 19.7100 ;
      RECT 10.6840 18.6165 10.7100 19.7100 ;
      RECT 10.5760 18.6165 10.6020 19.7100 ;
      RECT 10.4680 18.6165 10.4940 19.7100 ;
      RECT 10.3600 18.6165 10.3860 19.7100 ;
      RECT 10.2520 18.6165 10.2780 19.7100 ;
      RECT 10.1440 18.6165 10.1700 19.7100 ;
      RECT 10.0360 18.6165 10.0620 19.7100 ;
      RECT 9.9280 18.6165 9.9540 19.7100 ;
      RECT 9.8200 18.6165 9.8460 19.7100 ;
      RECT 9.7120 18.6165 9.7380 19.7100 ;
      RECT 9.6040 18.6165 9.6300 19.7100 ;
      RECT 9.4960 18.6165 9.5220 19.7100 ;
      RECT 9.3880 18.6165 9.4140 19.7100 ;
      RECT 9.1750 18.6165 9.2520 19.7100 ;
      RECT 7.2820 18.6165 7.3590 19.7100 ;
      RECT 7.1200 18.6165 7.1460 19.7100 ;
      RECT 7.0120 18.6165 7.0380 19.7100 ;
      RECT 6.9040 18.6165 6.9300 19.7100 ;
      RECT 6.7960 18.6165 6.8220 19.7100 ;
      RECT 6.6880 18.6165 6.7140 19.7100 ;
      RECT 6.5800 18.6165 6.6060 19.7100 ;
      RECT 6.4720 18.6165 6.4980 19.7100 ;
      RECT 6.3640 18.6165 6.3900 19.7100 ;
      RECT 6.2560 18.6165 6.2820 19.7100 ;
      RECT 6.1480 18.6165 6.1740 19.7100 ;
      RECT 6.0400 18.6165 6.0660 19.7100 ;
      RECT 5.9320 18.6165 5.9580 19.7100 ;
      RECT 5.8240 18.6165 5.8500 19.7100 ;
      RECT 5.7160 18.6165 5.7420 19.7100 ;
      RECT 5.6080 18.6165 5.6340 19.7100 ;
      RECT 5.5000 18.6165 5.5260 19.7100 ;
      RECT 5.3920 18.6165 5.4180 19.7100 ;
      RECT 5.2840 18.6165 5.3100 19.7100 ;
      RECT 5.1760 18.6165 5.2020 19.7100 ;
      RECT 5.0680 18.6165 5.0940 19.7100 ;
      RECT 4.9600 18.6165 4.9860 19.7100 ;
      RECT 4.8520 18.6165 4.8780 19.7100 ;
      RECT 4.7440 18.6165 4.7700 19.7100 ;
      RECT 4.6360 18.6165 4.6620 19.7100 ;
      RECT 4.5280 18.6165 4.5540 19.7100 ;
      RECT 4.4200 18.6165 4.4460 19.7100 ;
      RECT 4.3120 18.6165 4.3380 19.7100 ;
      RECT 4.2040 18.6165 4.2300 19.7100 ;
      RECT 4.0960 18.6165 4.1220 19.7100 ;
      RECT 3.9880 18.6165 4.0140 19.7100 ;
      RECT 3.8800 18.6165 3.9060 19.7100 ;
      RECT 3.7720 18.6165 3.7980 19.7100 ;
      RECT 3.6640 18.6165 3.6900 19.7100 ;
      RECT 3.5560 18.6165 3.5820 19.7100 ;
      RECT 3.4480 18.6165 3.4740 19.7100 ;
      RECT 3.3400 18.6165 3.3660 19.7100 ;
      RECT 3.2320 18.6165 3.2580 19.7100 ;
      RECT 3.1240 18.6165 3.1500 19.7100 ;
      RECT 3.0160 18.6165 3.0420 19.7100 ;
      RECT 2.9080 18.6165 2.9340 19.7100 ;
      RECT 2.8000 18.6165 2.8260 19.7100 ;
      RECT 2.6920 18.6165 2.7180 19.7100 ;
      RECT 2.5840 18.6165 2.6100 19.7100 ;
      RECT 2.4760 18.6165 2.5020 19.7100 ;
      RECT 2.3680 18.6165 2.3940 19.7100 ;
      RECT 2.2600 18.6165 2.2860 19.7100 ;
      RECT 2.1520 18.6165 2.1780 19.7100 ;
      RECT 2.0440 18.6165 2.0700 19.7100 ;
      RECT 1.9360 18.6165 1.9620 19.7100 ;
      RECT 1.8280 18.6165 1.8540 19.7100 ;
      RECT 1.7200 18.6165 1.7460 19.7100 ;
      RECT 1.6120 18.6165 1.6380 19.7100 ;
      RECT 1.5040 18.6165 1.5300 19.7100 ;
      RECT 1.3960 18.6165 1.4220 19.7100 ;
      RECT 1.2880 18.6165 1.3140 19.7100 ;
      RECT 1.1800 18.6165 1.2060 19.7100 ;
      RECT 1.0720 18.6165 1.0980 19.7100 ;
      RECT 0.9640 18.6165 0.9900 19.7100 ;
      RECT 0.8560 18.6165 0.8820 19.7100 ;
      RECT 0.7480 18.6165 0.7740 19.7100 ;
      RECT 0.6400 18.6165 0.6660 19.7100 ;
      RECT 0.5320 18.6165 0.5580 19.7100 ;
      RECT 0.4240 18.6165 0.4500 19.7100 ;
      RECT 0.3160 18.6165 0.3420 19.7100 ;
      RECT 0.2080 18.6165 0.2340 19.7100 ;
      RECT 0.0050 18.6165 0.0900 19.7100 ;
      RECT 8.6410 19.6965 8.7690 20.7900 ;
      RECT 8.6270 20.3620 8.7690 20.6845 ;
      RECT 8.4790 20.0890 8.5410 20.7900 ;
      RECT 8.4650 20.3985 8.5410 20.5520 ;
      RECT 8.4790 19.6965 8.5050 20.7900 ;
      RECT 8.4790 19.8175 8.5190 20.0570 ;
      RECT 8.4790 19.6965 8.5410 19.7855 ;
      RECT 8.1820 20.1470 8.3880 20.7900 ;
      RECT 8.3620 19.6965 8.3880 20.7900 ;
      RECT 8.1820 20.4240 8.4020 20.6820 ;
      RECT 8.1820 19.6965 8.2800 20.7900 ;
      RECT 7.7650 19.6965 7.8480 20.7900 ;
      RECT 7.7650 19.7850 7.8620 20.7205 ;
      RECT 16.4440 19.6965 16.5290 20.7900 ;
      RECT 16.3000 19.6965 16.3260 20.7900 ;
      RECT 16.1920 19.6965 16.2180 20.7900 ;
      RECT 16.0840 19.6965 16.1100 20.7900 ;
      RECT 15.9760 19.6965 16.0020 20.7900 ;
      RECT 15.8680 19.6965 15.8940 20.7900 ;
      RECT 15.7600 19.6965 15.7860 20.7900 ;
      RECT 15.6520 19.6965 15.6780 20.7900 ;
      RECT 15.5440 19.6965 15.5700 20.7900 ;
      RECT 15.4360 19.6965 15.4620 20.7900 ;
      RECT 15.3280 19.6965 15.3540 20.7900 ;
      RECT 15.2200 19.6965 15.2460 20.7900 ;
      RECT 15.1120 19.6965 15.1380 20.7900 ;
      RECT 15.0040 19.6965 15.0300 20.7900 ;
      RECT 14.8960 19.6965 14.9220 20.7900 ;
      RECT 14.7880 19.6965 14.8140 20.7900 ;
      RECT 14.6800 19.6965 14.7060 20.7900 ;
      RECT 14.5720 19.6965 14.5980 20.7900 ;
      RECT 14.4640 19.6965 14.4900 20.7900 ;
      RECT 14.3560 19.6965 14.3820 20.7900 ;
      RECT 14.2480 19.6965 14.2740 20.7900 ;
      RECT 14.1400 19.6965 14.1660 20.7900 ;
      RECT 14.0320 19.6965 14.0580 20.7900 ;
      RECT 13.9240 19.6965 13.9500 20.7900 ;
      RECT 13.8160 19.6965 13.8420 20.7900 ;
      RECT 13.7080 19.6965 13.7340 20.7900 ;
      RECT 13.6000 19.6965 13.6260 20.7900 ;
      RECT 13.4920 19.6965 13.5180 20.7900 ;
      RECT 13.3840 19.6965 13.4100 20.7900 ;
      RECT 13.2760 19.6965 13.3020 20.7900 ;
      RECT 13.1680 19.6965 13.1940 20.7900 ;
      RECT 13.0600 19.6965 13.0860 20.7900 ;
      RECT 12.9520 19.6965 12.9780 20.7900 ;
      RECT 12.8440 19.6965 12.8700 20.7900 ;
      RECT 12.7360 19.6965 12.7620 20.7900 ;
      RECT 12.6280 19.6965 12.6540 20.7900 ;
      RECT 12.5200 19.6965 12.5460 20.7900 ;
      RECT 12.4120 19.6965 12.4380 20.7900 ;
      RECT 12.3040 19.6965 12.3300 20.7900 ;
      RECT 12.1960 19.6965 12.2220 20.7900 ;
      RECT 12.0880 19.6965 12.1140 20.7900 ;
      RECT 11.9800 19.6965 12.0060 20.7900 ;
      RECT 11.8720 19.6965 11.8980 20.7900 ;
      RECT 11.7640 19.6965 11.7900 20.7900 ;
      RECT 11.6560 19.6965 11.6820 20.7900 ;
      RECT 11.5480 19.6965 11.5740 20.7900 ;
      RECT 11.4400 19.6965 11.4660 20.7900 ;
      RECT 11.3320 19.6965 11.3580 20.7900 ;
      RECT 11.2240 19.6965 11.2500 20.7900 ;
      RECT 11.1160 19.6965 11.1420 20.7900 ;
      RECT 11.0080 19.6965 11.0340 20.7900 ;
      RECT 10.9000 19.6965 10.9260 20.7900 ;
      RECT 10.7920 19.6965 10.8180 20.7900 ;
      RECT 10.6840 19.6965 10.7100 20.7900 ;
      RECT 10.5760 19.6965 10.6020 20.7900 ;
      RECT 10.4680 19.6965 10.4940 20.7900 ;
      RECT 10.3600 19.6965 10.3860 20.7900 ;
      RECT 10.2520 19.6965 10.2780 20.7900 ;
      RECT 10.1440 19.6965 10.1700 20.7900 ;
      RECT 10.0360 19.6965 10.0620 20.7900 ;
      RECT 9.9280 19.6965 9.9540 20.7900 ;
      RECT 9.8200 19.6965 9.8460 20.7900 ;
      RECT 9.7120 19.6965 9.7380 20.7900 ;
      RECT 9.6040 19.6965 9.6300 20.7900 ;
      RECT 9.4960 19.6965 9.5220 20.7900 ;
      RECT 9.3880 19.6965 9.4140 20.7900 ;
      RECT 9.1750 19.6965 9.2520 20.7900 ;
      RECT 7.2820 19.6965 7.3590 20.7900 ;
      RECT 7.1200 19.6965 7.1460 20.7900 ;
      RECT 7.0120 19.6965 7.0380 20.7900 ;
      RECT 6.9040 19.6965 6.9300 20.7900 ;
      RECT 6.7960 19.6965 6.8220 20.7900 ;
      RECT 6.6880 19.6965 6.7140 20.7900 ;
      RECT 6.5800 19.6965 6.6060 20.7900 ;
      RECT 6.4720 19.6965 6.4980 20.7900 ;
      RECT 6.3640 19.6965 6.3900 20.7900 ;
      RECT 6.2560 19.6965 6.2820 20.7900 ;
      RECT 6.1480 19.6965 6.1740 20.7900 ;
      RECT 6.0400 19.6965 6.0660 20.7900 ;
      RECT 5.9320 19.6965 5.9580 20.7900 ;
      RECT 5.8240 19.6965 5.8500 20.7900 ;
      RECT 5.7160 19.6965 5.7420 20.7900 ;
      RECT 5.6080 19.6965 5.6340 20.7900 ;
      RECT 5.5000 19.6965 5.5260 20.7900 ;
      RECT 5.3920 19.6965 5.4180 20.7900 ;
      RECT 5.2840 19.6965 5.3100 20.7900 ;
      RECT 5.1760 19.6965 5.2020 20.7900 ;
      RECT 5.0680 19.6965 5.0940 20.7900 ;
      RECT 4.9600 19.6965 4.9860 20.7900 ;
      RECT 4.8520 19.6965 4.8780 20.7900 ;
      RECT 4.7440 19.6965 4.7700 20.7900 ;
      RECT 4.6360 19.6965 4.6620 20.7900 ;
      RECT 4.5280 19.6965 4.5540 20.7900 ;
      RECT 4.4200 19.6965 4.4460 20.7900 ;
      RECT 4.3120 19.6965 4.3380 20.7900 ;
      RECT 4.2040 19.6965 4.2300 20.7900 ;
      RECT 4.0960 19.6965 4.1220 20.7900 ;
      RECT 3.9880 19.6965 4.0140 20.7900 ;
      RECT 3.8800 19.6965 3.9060 20.7900 ;
      RECT 3.7720 19.6965 3.7980 20.7900 ;
      RECT 3.6640 19.6965 3.6900 20.7900 ;
      RECT 3.5560 19.6965 3.5820 20.7900 ;
      RECT 3.4480 19.6965 3.4740 20.7900 ;
      RECT 3.3400 19.6965 3.3660 20.7900 ;
      RECT 3.2320 19.6965 3.2580 20.7900 ;
      RECT 3.1240 19.6965 3.1500 20.7900 ;
      RECT 3.0160 19.6965 3.0420 20.7900 ;
      RECT 2.9080 19.6965 2.9340 20.7900 ;
      RECT 2.8000 19.6965 2.8260 20.7900 ;
      RECT 2.6920 19.6965 2.7180 20.7900 ;
      RECT 2.5840 19.6965 2.6100 20.7900 ;
      RECT 2.4760 19.6965 2.5020 20.7900 ;
      RECT 2.3680 19.6965 2.3940 20.7900 ;
      RECT 2.2600 19.6965 2.2860 20.7900 ;
      RECT 2.1520 19.6965 2.1780 20.7900 ;
      RECT 2.0440 19.6965 2.0700 20.7900 ;
      RECT 1.9360 19.6965 1.9620 20.7900 ;
      RECT 1.8280 19.6965 1.8540 20.7900 ;
      RECT 1.7200 19.6965 1.7460 20.7900 ;
      RECT 1.6120 19.6965 1.6380 20.7900 ;
      RECT 1.5040 19.6965 1.5300 20.7900 ;
      RECT 1.3960 19.6965 1.4220 20.7900 ;
      RECT 1.2880 19.6965 1.3140 20.7900 ;
      RECT 1.1800 19.6965 1.2060 20.7900 ;
      RECT 1.0720 19.6965 1.0980 20.7900 ;
      RECT 0.9640 19.6965 0.9900 20.7900 ;
      RECT 0.8560 19.6965 0.8820 20.7900 ;
      RECT 0.7480 19.6965 0.7740 20.7900 ;
      RECT 0.6400 19.6965 0.6660 20.7900 ;
      RECT 0.5320 19.6965 0.5580 20.7900 ;
      RECT 0.4240 19.6965 0.4500 20.7900 ;
      RECT 0.3160 19.6965 0.3420 20.7900 ;
      RECT 0.2080 19.6965 0.2340 20.7900 ;
      RECT 0.0050 19.6965 0.0900 20.7900 ;
      RECT 8.6410 20.7765 8.7690 21.8700 ;
      RECT 8.6270 21.4420 8.7690 21.7645 ;
      RECT 8.4790 21.1690 8.5410 21.8700 ;
      RECT 8.4650 21.4785 8.5410 21.6320 ;
      RECT 8.4790 20.7765 8.5050 21.8700 ;
      RECT 8.4790 20.8975 8.5190 21.1370 ;
      RECT 8.4790 20.7765 8.5410 20.8655 ;
      RECT 8.1820 21.2270 8.3880 21.8700 ;
      RECT 8.3620 20.7765 8.3880 21.8700 ;
      RECT 8.1820 21.5040 8.4020 21.7620 ;
      RECT 8.1820 20.7765 8.2800 21.8700 ;
      RECT 7.7650 20.7765 7.8480 21.8700 ;
      RECT 7.7650 20.8650 7.8620 21.8005 ;
      RECT 16.4440 20.7765 16.5290 21.8700 ;
      RECT 16.3000 20.7765 16.3260 21.8700 ;
      RECT 16.1920 20.7765 16.2180 21.8700 ;
      RECT 16.0840 20.7765 16.1100 21.8700 ;
      RECT 15.9760 20.7765 16.0020 21.8700 ;
      RECT 15.8680 20.7765 15.8940 21.8700 ;
      RECT 15.7600 20.7765 15.7860 21.8700 ;
      RECT 15.6520 20.7765 15.6780 21.8700 ;
      RECT 15.5440 20.7765 15.5700 21.8700 ;
      RECT 15.4360 20.7765 15.4620 21.8700 ;
      RECT 15.3280 20.7765 15.3540 21.8700 ;
      RECT 15.2200 20.7765 15.2460 21.8700 ;
      RECT 15.1120 20.7765 15.1380 21.8700 ;
      RECT 15.0040 20.7765 15.0300 21.8700 ;
      RECT 14.8960 20.7765 14.9220 21.8700 ;
      RECT 14.7880 20.7765 14.8140 21.8700 ;
      RECT 14.6800 20.7765 14.7060 21.8700 ;
      RECT 14.5720 20.7765 14.5980 21.8700 ;
      RECT 14.4640 20.7765 14.4900 21.8700 ;
      RECT 14.3560 20.7765 14.3820 21.8700 ;
      RECT 14.2480 20.7765 14.2740 21.8700 ;
      RECT 14.1400 20.7765 14.1660 21.8700 ;
      RECT 14.0320 20.7765 14.0580 21.8700 ;
      RECT 13.9240 20.7765 13.9500 21.8700 ;
      RECT 13.8160 20.7765 13.8420 21.8700 ;
      RECT 13.7080 20.7765 13.7340 21.8700 ;
      RECT 13.6000 20.7765 13.6260 21.8700 ;
      RECT 13.4920 20.7765 13.5180 21.8700 ;
      RECT 13.3840 20.7765 13.4100 21.8700 ;
      RECT 13.2760 20.7765 13.3020 21.8700 ;
      RECT 13.1680 20.7765 13.1940 21.8700 ;
      RECT 13.0600 20.7765 13.0860 21.8700 ;
      RECT 12.9520 20.7765 12.9780 21.8700 ;
      RECT 12.8440 20.7765 12.8700 21.8700 ;
      RECT 12.7360 20.7765 12.7620 21.8700 ;
      RECT 12.6280 20.7765 12.6540 21.8700 ;
      RECT 12.5200 20.7765 12.5460 21.8700 ;
      RECT 12.4120 20.7765 12.4380 21.8700 ;
      RECT 12.3040 20.7765 12.3300 21.8700 ;
      RECT 12.1960 20.7765 12.2220 21.8700 ;
      RECT 12.0880 20.7765 12.1140 21.8700 ;
      RECT 11.9800 20.7765 12.0060 21.8700 ;
      RECT 11.8720 20.7765 11.8980 21.8700 ;
      RECT 11.7640 20.7765 11.7900 21.8700 ;
      RECT 11.6560 20.7765 11.6820 21.8700 ;
      RECT 11.5480 20.7765 11.5740 21.8700 ;
      RECT 11.4400 20.7765 11.4660 21.8700 ;
      RECT 11.3320 20.7765 11.3580 21.8700 ;
      RECT 11.2240 20.7765 11.2500 21.8700 ;
      RECT 11.1160 20.7765 11.1420 21.8700 ;
      RECT 11.0080 20.7765 11.0340 21.8700 ;
      RECT 10.9000 20.7765 10.9260 21.8700 ;
      RECT 10.7920 20.7765 10.8180 21.8700 ;
      RECT 10.6840 20.7765 10.7100 21.8700 ;
      RECT 10.5760 20.7765 10.6020 21.8700 ;
      RECT 10.4680 20.7765 10.4940 21.8700 ;
      RECT 10.3600 20.7765 10.3860 21.8700 ;
      RECT 10.2520 20.7765 10.2780 21.8700 ;
      RECT 10.1440 20.7765 10.1700 21.8700 ;
      RECT 10.0360 20.7765 10.0620 21.8700 ;
      RECT 9.9280 20.7765 9.9540 21.8700 ;
      RECT 9.8200 20.7765 9.8460 21.8700 ;
      RECT 9.7120 20.7765 9.7380 21.8700 ;
      RECT 9.6040 20.7765 9.6300 21.8700 ;
      RECT 9.4960 20.7765 9.5220 21.8700 ;
      RECT 9.3880 20.7765 9.4140 21.8700 ;
      RECT 9.1750 20.7765 9.2520 21.8700 ;
      RECT 7.2820 20.7765 7.3590 21.8700 ;
      RECT 7.1200 20.7765 7.1460 21.8700 ;
      RECT 7.0120 20.7765 7.0380 21.8700 ;
      RECT 6.9040 20.7765 6.9300 21.8700 ;
      RECT 6.7960 20.7765 6.8220 21.8700 ;
      RECT 6.6880 20.7765 6.7140 21.8700 ;
      RECT 6.5800 20.7765 6.6060 21.8700 ;
      RECT 6.4720 20.7765 6.4980 21.8700 ;
      RECT 6.3640 20.7765 6.3900 21.8700 ;
      RECT 6.2560 20.7765 6.2820 21.8700 ;
      RECT 6.1480 20.7765 6.1740 21.8700 ;
      RECT 6.0400 20.7765 6.0660 21.8700 ;
      RECT 5.9320 20.7765 5.9580 21.8700 ;
      RECT 5.8240 20.7765 5.8500 21.8700 ;
      RECT 5.7160 20.7765 5.7420 21.8700 ;
      RECT 5.6080 20.7765 5.6340 21.8700 ;
      RECT 5.5000 20.7765 5.5260 21.8700 ;
      RECT 5.3920 20.7765 5.4180 21.8700 ;
      RECT 5.2840 20.7765 5.3100 21.8700 ;
      RECT 5.1760 20.7765 5.2020 21.8700 ;
      RECT 5.0680 20.7765 5.0940 21.8700 ;
      RECT 4.9600 20.7765 4.9860 21.8700 ;
      RECT 4.8520 20.7765 4.8780 21.8700 ;
      RECT 4.7440 20.7765 4.7700 21.8700 ;
      RECT 4.6360 20.7765 4.6620 21.8700 ;
      RECT 4.5280 20.7765 4.5540 21.8700 ;
      RECT 4.4200 20.7765 4.4460 21.8700 ;
      RECT 4.3120 20.7765 4.3380 21.8700 ;
      RECT 4.2040 20.7765 4.2300 21.8700 ;
      RECT 4.0960 20.7765 4.1220 21.8700 ;
      RECT 3.9880 20.7765 4.0140 21.8700 ;
      RECT 3.8800 20.7765 3.9060 21.8700 ;
      RECT 3.7720 20.7765 3.7980 21.8700 ;
      RECT 3.6640 20.7765 3.6900 21.8700 ;
      RECT 3.5560 20.7765 3.5820 21.8700 ;
      RECT 3.4480 20.7765 3.4740 21.8700 ;
      RECT 3.3400 20.7765 3.3660 21.8700 ;
      RECT 3.2320 20.7765 3.2580 21.8700 ;
      RECT 3.1240 20.7765 3.1500 21.8700 ;
      RECT 3.0160 20.7765 3.0420 21.8700 ;
      RECT 2.9080 20.7765 2.9340 21.8700 ;
      RECT 2.8000 20.7765 2.8260 21.8700 ;
      RECT 2.6920 20.7765 2.7180 21.8700 ;
      RECT 2.5840 20.7765 2.6100 21.8700 ;
      RECT 2.4760 20.7765 2.5020 21.8700 ;
      RECT 2.3680 20.7765 2.3940 21.8700 ;
      RECT 2.2600 20.7765 2.2860 21.8700 ;
      RECT 2.1520 20.7765 2.1780 21.8700 ;
      RECT 2.0440 20.7765 2.0700 21.8700 ;
      RECT 1.9360 20.7765 1.9620 21.8700 ;
      RECT 1.8280 20.7765 1.8540 21.8700 ;
      RECT 1.7200 20.7765 1.7460 21.8700 ;
      RECT 1.6120 20.7765 1.6380 21.8700 ;
      RECT 1.5040 20.7765 1.5300 21.8700 ;
      RECT 1.3960 20.7765 1.4220 21.8700 ;
      RECT 1.2880 20.7765 1.3140 21.8700 ;
      RECT 1.1800 20.7765 1.2060 21.8700 ;
      RECT 1.0720 20.7765 1.0980 21.8700 ;
      RECT 0.9640 20.7765 0.9900 21.8700 ;
      RECT 0.8560 20.7765 0.8820 21.8700 ;
      RECT 0.7480 20.7765 0.7740 21.8700 ;
      RECT 0.6400 20.7765 0.6660 21.8700 ;
      RECT 0.5320 20.7765 0.5580 21.8700 ;
      RECT 0.4240 20.7765 0.4500 21.8700 ;
      RECT 0.3160 20.7765 0.3420 21.8700 ;
      RECT 0.2080 20.7765 0.2340 21.8700 ;
      RECT 0.0050 20.7765 0.0900 21.8700 ;
      RECT 8.6410 21.8565 8.7690 22.9500 ;
      RECT 8.6270 22.5220 8.7690 22.8445 ;
      RECT 8.4790 22.2490 8.5410 22.9500 ;
      RECT 8.4650 22.5585 8.5410 22.7120 ;
      RECT 8.4790 21.8565 8.5050 22.9500 ;
      RECT 8.4790 21.9775 8.5190 22.2170 ;
      RECT 8.4790 21.8565 8.5410 21.9455 ;
      RECT 8.1820 22.3070 8.3880 22.9500 ;
      RECT 8.3620 21.8565 8.3880 22.9500 ;
      RECT 8.1820 22.5840 8.4020 22.8420 ;
      RECT 8.1820 21.8565 8.2800 22.9500 ;
      RECT 7.7650 21.8565 7.8480 22.9500 ;
      RECT 7.7650 21.9450 7.8620 22.8805 ;
      RECT 16.4440 21.8565 16.5290 22.9500 ;
      RECT 16.3000 21.8565 16.3260 22.9500 ;
      RECT 16.1920 21.8565 16.2180 22.9500 ;
      RECT 16.0840 21.8565 16.1100 22.9500 ;
      RECT 15.9760 21.8565 16.0020 22.9500 ;
      RECT 15.8680 21.8565 15.8940 22.9500 ;
      RECT 15.7600 21.8565 15.7860 22.9500 ;
      RECT 15.6520 21.8565 15.6780 22.9500 ;
      RECT 15.5440 21.8565 15.5700 22.9500 ;
      RECT 15.4360 21.8565 15.4620 22.9500 ;
      RECT 15.3280 21.8565 15.3540 22.9500 ;
      RECT 15.2200 21.8565 15.2460 22.9500 ;
      RECT 15.1120 21.8565 15.1380 22.9500 ;
      RECT 15.0040 21.8565 15.0300 22.9500 ;
      RECT 14.8960 21.8565 14.9220 22.9500 ;
      RECT 14.7880 21.8565 14.8140 22.9500 ;
      RECT 14.6800 21.8565 14.7060 22.9500 ;
      RECT 14.5720 21.8565 14.5980 22.9500 ;
      RECT 14.4640 21.8565 14.4900 22.9500 ;
      RECT 14.3560 21.8565 14.3820 22.9500 ;
      RECT 14.2480 21.8565 14.2740 22.9500 ;
      RECT 14.1400 21.8565 14.1660 22.9500 ;
      RECT 14.0320 21.8565 14.0580 22.9500 ;
      RECT 13.9240 21.8565 13.9500 22.9500 ;
      RECT 13.8160 21.8565 13.8420 22.9500 ;
      RECT 13.7080 21.8565 13.7340 22.9500 ;
      RECT 13.6000 21.8565 13.6260 22.9500 ;
      RECT 13.4920 21.8565 13.5180 22.9500 ;
      RECT 13.3840 21.8565 13.4100 22.9500 ;
      RECT 13.2760 21.8565 13.3020 22.9500 ;
      RECT 13.1680 21.8565 13.1940 22.9500 ;
      RECT 13.0600 21.8565 13.0860 22.9500 ;
      RECT 12.9520 21.8565 12.9780 22.9500 ;
      RECT 12.8440 21.8565 12.8700 22.9500 ;
      RECT 12.7360 21.8565 12.7620 22.9500 ;
      RECT 12.6280 21.8565 12.6540 22.9500 ;
      RECT 12.5200 21.8565 12.5460 22.9500 ;
      RECT 12.4120 21.8565 12.4380 22.9500 ;
      RECT 12.3040 21.8565 12.3300 22.9500 ;
      RECT 12.1960 21.8565 12.2220 22.9500 ;
      RECT 12.0880 21.8565 12.1140 22.9500 ;
      RECT 11.9800 21.8565 12.0060 22.9500 ;
      RECT 11.8720 21.8565 11.8980 22.9500 ;
      RECT 11.7640 21.8565 11.7900 22.9500 ;
      RECT 11.6560 21.8565 11.6820 22.9500 ;
      RECT 11.5480 21.8565 11.5740 22.9500 ;
      RECT 11.4400 21.8565 11.4660 22.9500 ;
      RECT 11.3320 21.8565 11.3580 22.9500 ;
      RECT 11.2240 21.8565 11.2500 22.9500 ;
      RECT 11.1160 21.8565 11.1420 22.9500 ;
      RECT 11.0080 21.8565 11.0340 22.9500 ;
      RECT 10.9000 21.8565 10.9260 22.9500 ;
      RECT 10.7920 21.8565 10.8180 22.9500 ;
      RECT 10.6840 21.8565 10.7100 22.9500 ;
      RECT 10.5760 21.8565 10.6020 22.9500 ;
      RECT 10.4680 21.8565 10.4940 22.9500 ;
      RECT 10.3600 21.8565 10.3860 22.9500 ;
      RECT 10.2520 21.8565 10.2780 22.9500 ;
      RECT 10.1440 21.8565 10.1700 22.9500 ;
      RECT 10.0360 21.8565 10.0620 22.9500 ;
      RECT 9.9280 21.8565 9.9540 22.9500 ;
      RECT 9.8200 21.8565 9.8460 22.9500 ;
      RECT 9.7120 21.8565 9.7380 22.9500 ;
      RECT 9.6040 21.8565 9.6300 22.9500 ;
      RECT 9.4960 21.8565 9.5220 22.9500 ;
      RECT 9.3880 21.8565 9.4140 22.9500 ;
      RECT 9.1750 21.8565 9.2520 22.9500 ;
      RECT 7.2820 21.8565 7.3590 22.9500 ;
      RECT 7.1200 21.8565 7.1460 22.9500 ;
      RECT 7.0120 21.8565 7.0380 22.9500 ;
      RECT 6.9040 21.8565 6.9300 22.9500 ;
      RECT 6.7960 21.8565 6.8220 22.9500 ;
      RECT 6.6880 21.8565 6.7140 22.9500 ;
      RECT 6.5800 21.8565 6.6060 22.9500 ;
      RECT 6.4720 21.8565 6.4980 22.9500 ;
      RECT 6.3640 21.8565 6.3900 22.9500 ;
      RECT 6.2560 21.8565 6.2820 22.9500 ;
      RECT 6.1480 21.8565 6.1740 22.9500 ;
      RECT 6.0400 21.8565 6.0660 22.9500 ;
      RECT 5.9320 21.8565 5.9580 22.9500 ;
      RECT 5.8240 21.8565 5.8500 22.9500 ;
      RECT 5.7160 21.8565 5.7420 22.9500 ;
      RECT 5.6080 21.8565 5.6340 22.9500 ;
      RECT 5.5000 21.8565 5.5260 22.9500 ;
      RECT 5.3920 21.8565 5.4180 22.9500 ;
      RECT 5.2840 21.8565 5.3100 22.9500 ;
      RECT 5.1760 21.8565 5.2020 22.9500 ;
      RECT 5.0680 21.8565 5.0940 22.9500 ;
      RECT 4.9600 21.8565 4.9860 22.9500 ;
      RECT 4.8520 21.8565 4.8780 22.9500 ;
      RECT 4.7440 21.8565 4.7700 22.9500 ;
      RECT 4.6360 21.8565 4.6620 22.9500 ;
      RECT 4.5280 21.8565 4.5540 22.9500 ;
      RECT 4.4200 21.8565 4.4460 22.9500 ;
      RECT 4.3120 21.8565 4.3380 22.9500 ;
      RECT 4.2040 21.8565 4.2300 22.9500 ;
      RECT 4.0960 21.8565 4.1220 22.9500 ;
      RECT 3.9880 21.8565 4.0140 22.9500 ;
      RECT 3.8800 21.8565 3.9060 22.9500 ;
      RECT 3.7720 21.8565 3.7980 22.9500 ;
      RECT 3.6640 21.8565 3.6900 22.9500 ;
      RECT 3.5560 21.8565 3.5820 22.9500 ;
      RECT 3.4480 21.8565 3.4740 22.9500 ;
      RECT 3.3400 21.8565 3.3660 22.9500 ;
      RECT 3.2320 21.8565 3.2580 22.9500 ;
      RECT 3.1240 21.8565 3.1500 22.9500 ;
      RECT 3.0160 21.8565 3.0420 22.9500 ;
      RECT 2.9080 21.8565 2.9340 22.9500 ;
      RECT 2.8000 21.8565 2.8260 22.9500 ;
      RECT 2.6920 21.8565 2.7180 22.9500 ;
      RECT 2.5840 21.8565 2.6100 22.9500 ;
      RECT 2.4760 21.8565 2.5020 22.9500 ;
      RECT 2.3680 21.8565 2.3940 22.9500 ;
      RECT 2.2600 21.8565 2.2860 22.9500 ;
      RECT 2.1520 21.8565 2.1780 22.9500 ;
      RECT 2.0440 21.8565 2.0700 22.9500 ;
      RECT 1.9360 21.8565 1.9620 22.9500 ;
      RECT 1.8280 21.8565 1.8540 22.9500 ;
      RECT 1.7200 21.8565 1.7460 22.9500 ;
      RECT 1.6120 21.8565 1.6380 22.9500 ;
      RECT 1.5040 21.8565 1.5300 22.9500 ;
      RECT 1.3960 21.8565 1.4220 22.9500 ;
      RECT 1.2880 21.8565 1.3140 22.9500 ;
      RECT 1.1800 21.8565 1.2060 22.9500 ;
      RECT 1.0720 21.8565 1.0980 22.9500 ;
      RECT 0.9640 21.8565 0.9900 22.9500 ;
      RECT 0.8560 21.8565 0.8820 22.9500 ;
      RECT 0.7480 21.8565 0.7740 22.9500 ;
      RECT 0.6400 21.8565 0.6660 22.9500 ;
      RECT 0.5320 21.8565 0.5580 22.9500 ;
      RECT 0.4240 21.8565 0.4500 22.9500 ;
      RECT 0.3160 21.8565 0.3420 22.9500 ;
      RECT 0.2080 21.8565 0.2340 22.9500 ;
      RECT 0.0050 21.8565 0.0900 22.9500 ;
      RECT 8.6410 22.9365 8.7690 24.0300 ;
      RECT 8.6270 23.6020 8.7690 23.9245 ;
      RECT 8.4790 23.3290 8.5410 24.0300 ;
      RECT 8.4650 23.6385 8.5410 23.7920 ;
      RECT 8.4790 22.9365 8.5050 24.0300 ;
      RECT 8.4790 23.0575 8.5190 23.2970 ;
      RECT 8.4790 22.9365 8.5410 23.0255 ;
      RECT 8.1820 23.3870 8.3880 24.0300 ;
      RECT 8.3620 22.9365 8.3880 24.0300 ;
      RECT 8.1820 23.6640 8.4020 23.9220 ;
      RECT 8.1820 22.9365 8.2800 24.0300 ;
      RECT 7.7650 22.9365 7.8480 24.0300 ;
      RECT 7.7650 23.0250 7.8620 23.9605 ;
      RECT 16.4440 22.9365 16.5290 24.0300 ;
      RECT 16.3000 22.9365 16.3260 24.0300 ;
      RECT 16.1920 22.9365 16.2180 24.0300 ;
      RECT 16.0840 22.9365 16.1100 24.0300 ;
      RECT 15.9760 22.9365 16.0020 24.0300 ;
      RECT 15.8680 22.9365 15.8940 24.0300 ;
      RECT 15.7600 22.9365 15.7860 24.0300 ;
      RECT 15.6520 22.9365 15.6780 24.0300 ;
      RECT 15.5440 22.9365 15.5700 24.0300 ;
      RECT 15.4360 22.9365 15.4620 24.0300 ;
      RECT 15.3280 22.9365 15.3540 24.0300 ;
      RECT 15.2200 22.9365 15.2460 24.0300 ;
      RECT 15.1120 22.9365 15.1380 24.0300 ;
      RECT 15.0040 22.9365 15.0300 24.0300 ;
      RECT 14.8960 22.9365 14.9220 24.0300 ;
      RECT 14.7880 22.9365 14.8140 24.0300 ;
      RECT 14.6800 22.9365 14.7060 24.0300 ;
      RECT 14.5720 22.9365 14.5980 24.0300 ;
      RECT 14.4640 22.9365 14.4900 24.0300 ;
      RECT 14.3560 22.9365 14.3820 24.0300 ;
      RECT 14.2480 22.9365 14.2740 24.0300 ;
      RECT 14.1400 22.9365 14.1660 24.0300 ;
      RECT 14.0320 22.9365 14.0580 24.0300 ;
      RECT 13.9240 22.9365 13.9500 24.0300 ;
      RECT 13.8160 22.9365 13.8420 24.0300 ;
      RECT 13.7080 22.9365 13.7340 24.0300 ;
      RECT 13.6000 22.9365 13.6260 24.0300 ;
      RECT 13.4920 22.9365 13.5180 24.0300 ;
      RECT 13.3840 22.9365 13.4100 24.0300 ;
      RECT 13.2760 22.9365 13.3020 24.0300 ;
      RECT 13.1680 22.9365 13.1940 24.0300 ;
      RECT 13.0600 22.9365 13.0860 24.0300 ;
      RECT 12.9520 22.9365 12.9780 24.0300 ;
      RECT 12.8440 22.9365 12.8700 24.0300 ;
      RECT 12.7360 22.9365 12.7620 24.0300 ;
      RECT 12.6280 22.9365 12.6540 24.0300 ;
      RECT 12.5200 22.9365 12.5460 24.0300 ;
      RECT 12.4120 22.9365 12.4380 24.0300 ;
      RECT 12.3040 22.9365 12.3300 24.0300 ;
      RECT 12.1960 22.9365 12.2220 24.0300 ;
      RECT 12.0880 22.9365 12.1140 24.0300 ;
      RECT 11.9800 22.9365 12.0060 24.0300 ;
      RECT 11.8720 22.9365 11.8980 24.0300 ;
      RECT 11.7640 22.9365 11.7900 24.0300 ;
      RECT 11.6560 22.9365 11.6820 24.0300 ;
      RECT 11.5480 22.9365 11.5740 24.0300 ;
      RECT 11.4400 22.9365 11.4660 24.0300 ;
      RECT 11.3320 22.9365 11.3580 24.0300 ;
      RECT 11.2240 22.9365 11.2500 24.0300 ;
      RECT 11.1160 22.9365 11.1420 24.0300 ;
      RECT 11.0080 22.9365 11.0340 24.0300 ;
      RECT 10.9000 22.9365 10.9260 24.0300 ;
      RECT 10.7920 22.9365 10.8180 24.0300 ;
      RECT 10.6840 22.9365 10.7100 24.0300 ;
      RECT 10.5760 22.9365 10.6020 24.0300 ;
      RECT 10.4680 22.9365 10.4940 24.0300 ;
      RECT 10.3600 22.9365 10.3860 24.0300 ;
      RECT 10.2520 22.9365 10.2780 24.0300 ;
      RECT 10.1440 22.9365 10.1700 24.0300 ;
      RECT 10.0360 22.9365 10.0620 24.0300 ;
      RECT 9.9280 22.9365 9.9540 24.0300 ;
      RECT 9.8200 22.9365 9.8460 24.0300 ;
      RECT 9.7120 22.9365 9.7380 24.0300 ;
      RECT 9.6040 22.9365 9.6300 24.0300 ;
      RECT 9.4960 22.9365 9.5220 24.0300 ;
      RECT 9.3880 22.9365 9.4140 24.0300 ;
      RECT 9.1750 22.9365 9.2520 24.0300 ;
      RECT 7.2820 22.9365 7.3590 24.0300 ;
      RECT 7.1200 22.9365 7.1460 24.0300 ;
      RECT 7.0120 22.9365 7.0380 24.0300 ;
      RECT 6.9040 22.9365 6.9300 24.0300 ;
      RECT 6.7960 22.9365 6.8220 24.0300 ;
      RECT 6.6880 22.9365 6.7140 24.0300 ;
      RECT 6.5800 22.9365 6.6060 24.0300 ;
      RECT 6.4720 22.9365 6.4980 24.0300 ;
      RECT 6.3640 22.9365 6.3900 24.0300 ;
      RECT 6.2560 22.9365 6.2820 24.0300 ;
      RECT 6.1480 22.9365 6.1740 24.0300 ;
      RECT 6.0400 22.9365 6.0660 24.0300 ;
      RECT 5.9320 22.9365 5.9580 24.0300 ;
      RECT 5.8240 22.9365 5.8500 24.0300 ;
      RECT 5.7160 22.9365 5.7420 24.0300 ;
      RECT 5.6080 22.9365 5.6340 24.0300 ;
      RECT 5.5000 22.9365 5.5260 24.0300 ;
      RECT 5.3920 22.9365 5.4180 24.0300 ;
      RECT 5.2840 22.9365 5.3100 24.0300 ;
      RECT 5.1760 22.9365 5.2020 24.0300 ;
      RECT 5.0680 22.9365 5.0940 24.0300 ;
      RECT 4.9600 22.9365 4.9860 24.0300 ;
      RECT 4.8520 22.9365 4.8780 24.0300 ;
      RECT 4.7440 22.9365 4.7700 24.0300 ;
      RECT 4.6360 22.9365 4.6620 24.0300 ;
      RECT 4.5280 22.9365 4.5540 24.0300 ;
      RECT 4.4200 22.9365 4.4460 24.0300 ;
      RECT 4.3120 22.9365 4.3380 24.0300 ;
      RECT 4.2040 22.9365 4.2300 24.0300 ;
      RECT 4.0960 22.9365 4.1220 24.0300 ;
      RECT 3.9880 22.9365 4.0140 24.0300 ;
      RECT 3.8800 22.9365 3.9060 24.0300 ;
      RECT 3.7720 22.9365 3.7980 24.0300 ;
      RECT 3.6640 22.9365 3.6900 24.0300 ;
      RECT 3.5560 22.9365 3.5820 24.0300 ;
      RECT 3.4480 22.9365 3.4740 24.0300 ;
      RECT 3.3400 22.9365 3.3660 24.0300 ;
      RECT 3.2320 22.9365 3.2580 24.0300 ;
      RECT 3.1240 22.9365 3.1500 24.0300 ;
      RECT 3.0160 22.9365 3.0420 24.0300 ;
      RECT 2.9080 22.9365 2.9340 24.0300 ;
      RECT 2.8000 22.9365 2.8260 24.0300 ;
      RECT 2.6920 22.9365 2.7180 24.0300 ;
      RECT 2.5840 22.9365 2.6100 24.0300 ;
      RECT 2.4760 22.9365 2.5020 24.0300 ;
      RECT 2.3680 22.9365 2.3940 24.0300 ;
      RECT 2.2600 22.9365 2.2860 24.0300 ;
      RECT 2.1520 22.9365 2.1780 24.0300 ;
      RECT 2.0440 22.9365 2.0700 24.0300 ;
      RECT 1.9360 22.9365 1.9620 24.0300 ;
      RECT 1.8280 22.9365 1.8540 24.0300 ;
      RECT 1.7200 22.9365 1.7460 24.0300 ;
      RECT 1.6120 22.9365 1.6380 24.0300 ;
      RECT 1.5040 22.9365 1.5300 24.0300 ;
      RECT 1.3960 22.9365 1.4220 24.0300 ;
      RECT 1.2880 22.9365 1.3140 24.0300 ;
      RECT 1.1800 22.9365 1.2060 24.0300 ;
      RECT 1.0720 22.9365 1.0980 24.0300 ;
      RECT 0.9640 22.9365 0.9900 24.0300 ;
      RECT 0.8560 22.9365 0.8820 24.0300 ;
      RECT 0.7480 22.9365 0.7740 24.0300 ;
      RECT 0.6400 22.9365 0.6660 24.0300 ;
      RECT 0.5320 22.9365 0.5580 24.0300 ;
      RECT 0.4240 22.9365 0.4500 24.0300 ;
      RECT 0.3160 22.9365 0.3420 24.0300 ;
      RECT 0.2080 22.9365 0.2340 24.0300 ;
      RECT 0.0050 22.9365 0.0900 24.0300 ;
      RECT 8.6410 24.0165 8.7690 25.1100 ;
      RECT 8.6270 24.6820 8.7690 25.0045 ;
      RECT 8.4790 24.4090 8.5410 25.1100 ;
      RECT 8.4650 24.7185 8.5410 24.8720 ;
      RECT 8.4790 24.0165 8.5050 25.1100 ;
      RECT 8.4790 24.1375 8.5190 24.3770 ;
      RECT 8.4790 24.0165 8.5410 24.1055 ;
      RECT 8.1820 24.4670 8.3880 25.1100 ;
      RECT 8.3620 24.0165 8.3880 25.1100 ;
      RECT 8.1820 24.7440 8.4020 25.0020 ;
      RECT 8.1820 24.0165 8.2800 25.1100 ;
      RECT 7.7650 24.0165 7.8480 25.1100 ;
      RECT 7.7650 24.1050 7.8620 25.0405 ;
      RECT 16.4440 24.0165 16.5290 25.1100 ;
      RECT 16.3000 24.0165 16.3260 25.1100 ;
      RECT 16.1920 24.0165 16.2180 25.1100 ;
      RECT 16.0840 24.0165 16.1100 25.1100 ;
      RECT 15.9760 24.0165 16.0020 25.1100 ;
      RECT 15.8680 24.0165 15.8940 25.1100 ;
      RECT 15.7600 24.0165 15.7860 25.1100 ;
      RECT 15.6520 24.0165 15.6780 25.1100 ;
      RECT 15.5440 24.0165 15.5700 25.1100 ;
      RECT 15.4360 24.0165 15.4620 25.1100 ;
      RECT 15.3280 24.0165 15.3540 25.1100 ;
      RECT 15.2200 24.0165 15.2460 25.1100 ;
      RECT 15.1120 24.0165 15.1380 25.1100 ;
      RECT 15.0040 24.0165 15.0300 25.1100 ;
      RECT 14.8960 24.0165 14.9220 25.1100 ;
      RECT 14.7880 24.0165 14.8140 25.1100 ;
      RECT 14.6800 24.0165 14.7060 25.1100 ;
      RECT 14.5720 24.0165 14.5980 25.1100 ;
      RECT 14.4640 24.0165 14.4900 25.1100 ;
      RECT 14.3560 24.0165 14.3820 25.1100 ;
      RECT 14.2480 24.0165 14.2740 25.1100 ;
      RECT 14.1400 24.0165 14.1660 25.1100 ;
      RECT 14.0320 24.0165 14.0580 25.1100 ;
      RECT 13.9240 24.0165 13.9500 25.1100 ;
      RECT 13.8160 24.0165 13.8420 25.1100 ;
      RECT 13.7080 24.0165 13.7340 25.1100 ;
      RECT 13.6000 24.0165 13.6260 25.1100 ;
      RECT 13.4920 24.0165 13.5180 25.1100 ;
      RECT 13.3840 24.0165 13.4100 25.1100 ;
      RECT 13.2760 24.0165 13.3020 25.1100 ;
      RECT 13.1680 24.0165 13.1940 25.1100 ;
      RECT 13.0600 24.0165 13.0860 25.1100 ;
      RECT 12.9520 24.0165 12.9780 25.1100 ;
      RECT 12.8440 24.0165 12.8700 25.1100 ;
      RECT 12.7360 24.0165 12.7620 25.1100 ;
      RECT 12.6280 24.0165 12.6540 25.1100 ;
      RECT 12.5200 24.0165 12.5460 25.1100 ;
      RECT 12.4120 24.0165 12.4380 25.1100 ;
      RECT 12.3040 24.0165 12.3300 25.1100 ;
      RECT 12.1960 24.0165 12.2220 25.1100 ;
      RECT 12.0880 24.0165 12.1140 25.1100 ;
      RECT 11.9800 24.0165 12.0060 25.1100 ;
      RECT 11.8720 24.0165 11.8980 25.1100 ;
      RECT 11.7640 24.0165 11.7900 25.1100 ;
      RECT 11.6560 24.0165 11.6820 25.1100 ;
      RECT 11.5480 24.0165 11.5740 25.1100 ;
      RECT 11.4400 24.0165 11.4660 25.1100 ;
      RECT 11.3320 24.0165 11.3580 25.1100 ;
      RECT 11.2240 24.0165 11.2500 25.1100 ;
      RECT 11.1160 24.0165 11.1420 25.1100 ;
      RECT 11.0080 24.0165 11.0340 25.1100 ;
      RECT 10.9000 24.0165 10.9260 25.1100 ;
      RECT 10.7920 24.0165 10.8180 25.1100 ;
      RECT 10.6840 24.0165 10.7100 25.1100 ;
      RECT 10.5760 24.0165 10.6020 25.1100 ;
      RECT 10.4680 24.0165 10.4940 25.1100 ;
      RECT 10.3600 24.0165 10.3860 25.1100 ;
      RECT 10.2520 24.0165 10.2780 25.1100 ;
      RECT 10.1440 24.0165 10.1700 25.1100 ;
      RECT 10.0360 24.0165 10.0620 25.1100 ;
      RECT 9.9280 24.0165 9.9540 25.1100 ;
      RECT 9.8200 24.0165 9.8460 25.1100 ;
      RECT 9.7120 24.0165 9.7380 25.1100 ;
      RECT 9.6040 24.0165 9.6300 25.1100 ;
      RECT 9.4960 24.0165 9.5220 25.1100 ;
      RECT 9.3880 24.0165 9.4140 25.1100 ;
      RECT 9.1750 24.0165 9.2520 25.1100 ;
      RECT 7.2820 24.0165 7.3590 25.1100 ;
      RECT 7.1200 24.0165 7.1460 25.1100 ;
      RECT 7.0120 24.0165 7.0380 25.1100 ;
      RECT 6.9040 24.0165 6.9300 25.1100 ;
      RECT 6.7960 24.0165 6.8220 25.1100 ;
      RECT 6.6880 24.0165 6.7140 25.1100 ;
      RECT 6.5800 24.0165 6.6060 25.1100 ;
      RECT 6.4720 24.0165 6.4980 25.1100 ;
      RECT 6.3640 24.0165 6.3900 25.1100 ;
      RECT 6.2560 24.0165 6.2820 25.1100 ;
      RECT 6.1480 24.0165 6.1740 25.1100 ;
      RECT 6.0400 24.0165 6.0660 25.1100 ;
      RECT 5.9320 24.0165 5.9580 25.1100 ;
      RECT 5.8240 24.0165 5.8500 25.1100 ;
      RECT 5.7160 24.0165 5.7420 25.1100 ;
      RECT 5.6080 24.0165 5.6340 25.1100 ;
      RECT 5.5000 24.0165 5.5260 25.1100 ;
      RECT 5.3920 24.0165 5.4180 25.1100 ;
      RECT 5.2840 24.0165 5.3100 25.1100 ;
      RECT 5.1760 24.0165 5.2020 25.1100 ;
      RECT 5.0680 24.0165 5.0940 25.1100 ;
      RECT 4.9600 24.0165 4.9860 25.1100 ;
      RECT 4.8520 24.0165 4.8780 25.1100 ;
      RECT 4.7440 24.0165 4.7700 25.1100 ;
      RECT 4.6360 24.0165 4.6620 25.1100 ;
      RECT 4.5280 24.0165 4.5540 25.1100 ;
      RECT 4.4200 24.0165 4.4460 25.1100 ;
      RECT 4.3120 24.0165 4.3380 25.1100 ;
      RECT 4.2040 24.0165 4.2300 25.1100 ;
      RECT 4.0960 24.0165 4.1220 25.1100 ;
      RECT 3.9880 24.0165 4.0140 25.1100 ;
      RECT 3.8800 24.0165 3.9060 25.1100 ;
      RECT 3.7720 24.0165 3.7980 25.1100 ;
      RECT 3.6640 24.0165 3.6900 25.1100 ;
      RECT 3.5560 24.0165 3.5820 25.1100 ;
      RECT 3.4480 24.0165 3.4740 25.1100 ;
      RECT 3.3400 24.0165 3.3660 25.1100 ;
      RECT 3.2320 24.0165 3.2580 25.1100 ;
      RECT 3.1240 24.0165 3.1500 25.1100 ;
      RECT 3.0160 24.0165 3.0420 25.1100 ;
      RECT 2.9080 24.0165 2.9340 25.1100 ;
      RECT 2.8000 24.0165 2.8260 25.1100 ;
      RECT 2.6920 24.0165 2.7180 25.1100 ;
      RECT 2.5840 24.0165 2.6100 25.1100 ;
      RECT 2.4760 24.0165 2.5020 25.1100 ;
      RECT 2.3680 24.0165 2.3940 25.1100 ;
      RECT 2.2600 24.0165 2.2860 25.1100 ;
      RECT 2.1520 24.0165 2.1780 25.1100 ;
      RECT 2.0440 24.0165 2.0700 25.1100 ;
      RECT 1.9360 24.0165 1.9620 25.1100 ;
      RECT 1.8280 24.0165 1.8540 25.1100 ;
      RECT 1.7200 24.0165 1.7460 25.1100 ;
      RECT 1.6120 24.0165 1.6380 25.1100 ;
      RECT 1.5040 24.0165 1.5300 25.1100 ;
      RECT 1.3960 24.0165 1.4220 25.1100 ;
      RECT 1.2880 24.0165 1.3140 25.1100 ;
      RECT 1.1800 24.0165 1.2060 25.1100 ;
      RECT 1.0720 24.0165 1.0980 25.1100 ;
      RECT 0.9640 24.0165 0.9900 25.1100 ;
      RECT 0.8560 24.0165 0.8820 25.1100 ;
      RECT 0.7480 24.0165 0.7740 25.1100 ;
      RECT 0.6400 24.0165 0.6660 25.1100 ;
      RECT 0.5320 24.0165 0.5580 25.1100 ;
      RECT 0.4240 24.0165 0.4500 25.1100 ;
      RECT 0.3160 24.0165 0.3420 25.1100 ;
      RECT 0.2080 24.0165 0.2340 25.1100 ;
      RECT 0.0050 24.0165 0.0900 25.1100 ;
      RECT 8.6410 25.0965 8.7690 26.1900 ;
      RECT 8.6270 25.7620 8.7690 26.0845 ;
      RECT 8.4790 25.4890 8.5410 26.1900 ;
      RECT 8.4650 25.7985 8.5410 25.9520 ;
      RECT 8.4790 25.0965 8.5050 26.1900 ;
      RECT 8.4790 25.2175 8.5190 25.4570 ;
      RECT 8.4790 25.0965 8.5410 25.1855 ;
      RECT 8.1820 25.5470 8.3880 26.1900 ;
      RECT 8.3620 25.0965 8.3880 26.1900 ;
      RECT 8.1820 25.8240 8.4020 26.0820 ;
      RECT 8.1820 25.0965 8.2800 26.1900 ;
      RECT 7.7650 25.0965 7.8480 26.1900 ;
      RECT 7.7650 25.1850 7.8620 26.1205 ;
      RECT 16.4440 25.0965 16.5290 26.1900 ;
      RECT 16.3000 25.0965 16.3260 26.1900 ;
      RECT 16.1920 25.0965 16.2180 26.1900 ;
      RECT 16.0840 25.0965 16.1100 26.1900 ;
      RECT 15.9760 25.0965 16.0020 26.1900 ;
      RECT 15.8680 25.0965 15.8940 26.1900 ;
      RECT 15.7600 25.0965 15.7860 26.1900 ;
      RECT 15.6520 25.0965 15.6780 26.1900 ;
      RECT 15.5440 25.0965 15.5700 26.1900 ;
      RECT 15.4360 25.0965 15.4620 26.1900 ;
      RECT 15.3280 25.0965 15.3540 26.1900 ;
      RECT 15.2200 25.0965 15.2460 26.1900 ;
      RECT 15.1120 25.0965 15.1380 26.1900 ;
      RECT 15.0040 25.0965 15.0300 26.1900 ;
      RECT 14.8960 25.0965 14.9220 26.1900 ;
      RECT 14.7880 25.0965 14.8140 26.1900 ;
      RECT 14.6800 25.0965 14.7060 26.1900 ;
      RECT 14.5720 25.0965 14.5980 26.1900 ;
      RECT 14.4640 25.0965 14.4900 26.1900 ;
      RECT 14.3560 25.0965 14.3820 26.1900 ;
      RECT 14.2480 25.0965 14.2740 26.1900 ;
      RECT 14.1400 25.0965 14.1660 26.1900 ;
      RECT 14.0320 25.0965 14.0580 26.1900 ;
      RECT 13.9240 25.0965 13.9500 26.1900 ;
      RECT 13.8160 25.0965 13.8420 26.1900 ;
      RECT 13.7080 25.0965 13.7340 26.1900 ;
      RECT 13.6000 25.0965 13.6260 26.1900 ;
      RECT 13.4920 25.0965 13.5180 26.1900 ;
      RECT 13.3840 25.0965 13.4100 26.1900 ;
      RECT 13.2760 25.0965 13.3020 26.1900 ;
      RECT 13.1680 25.0965 13.1940 26.1900 ;
      RECT 13.0600 25.0965 13.0860 26.1900 ;
      RECT 12.9520 25.0965 12.9780 26.1900 ;
      RECT 12.8440 25.0965 12.8700 26.1900 ;
      RECT 12.7360 25.0965 12.7620 26.1900 ;
      RECT 12.6280 25.0965 12.6540 26.1900 ;
      RECT 12.5200 25.0965 12.5460 26.1900 ;
      RECT 12.4120 25.0965 12.4380 26.1900 ;
      RECT 12.3040 25.0965 12.3300 26.1900 ;
      RECT 12.1960 25.0965 12.2220 26.1900 ;
      RECT 12.0880 25.0965 12.1140 26.1900 ;
      RECT 11.9800 25.0965 12.0060 26.1900 ;
      RECT 11.8720 25.0965 11.8980 26.1900 ;
      RECT 11.7640 25.0965 11.7900 26.1900 ;
      RECT 11.6560 25.0965 11.6820 26.1900 ;
      RECT 11.5480 25.0965 11.5740 26.1900 ;
      RECT 11.4400 25.0965 11.4660 26.1900 ;
      RECT 11.3320 25.0965 11.3580 26.1900 ;
      RECT 11.2240 25.0965 11.2500 26.1900 ;
      RECT 11.1160 25.0965 11.1420 26.1900 ;
      RECT 11.0080 25.0965 11.0340 26.1900 ;
      RECT 10.9000 25.0965 10.9260 26.1900 ;
      RECT 10.7920 25.0965 10.8180 26.1900 ;
      RECT 10.6840 25.0965 10.7100 26.1900 ;
      RECT 10.5760 25.0965 10.6020 26.1900 ;
      RECT 10.4680 25.0965 10.4940 26.1900 ;
      RECT 10.3600 25.0965 10.3860 26.1900 ;
      RECT 10.2520 25.0965 10.2780 26.1900 ;
      RECT 10.1440 25.0965 10.1700 26.1900 ;
      RECT 10.0360 25.0965 10.0620 26.1900 ;
      RECT 9.9280 25.0965 9.9540 26.1900 ;
      RECT 9.8200 25.0965 9.8460 26.1900 ;
      RECT 9.7120 25.0965 9.7380 26.1900 ;
      RECT 9.6040 25.0965 9.6300 26.1900 ;
      RECT 9.4960 25.0965 9.5220 26.1900 ;
      RECT 9.3880 25.0965 9.4140 26.1900 ;
      RECT 9.1750 25.0965 9.2520 26.1900 ;
      RECT 7.2820 25.0965 7.3590 26.1900 ;
      RECT 7.1200 25.0965 7.1460 26.1900 ;
      RECT 7.0120 25.0965 7.0380 26.1900 ;
      RECT 6.9040 25.0965 6.9300 26.1900 ;
      RECT 6.7960 25.0965 6.8220 26.1900 ;
      RECT 6.6880 25.0965 6.7140 26.1900 ;
      RECT 6.5800 25.0965 6.6060 26.1900 ;
      RECT 6.4720 25.0965 6.4980 26.1900 ;
      RECT 6.3640 25.0965 6.3900 26.1900 ;
      RECT 6.2560 25.0965 6.2820 26.1900 ;
      RECT 6.1480 25.0965 6.1740 26.1900 ;
      RECT 6.0400 25.0965 6.0660 26.1900 ;
      RECT 5.9320 25.0965 5.9580 26.1900 ;
      RECT 5.8240 25.0965 5.8500 26.1900 ;
      RECT 5.7160 25.0965 5.7420 26.1900 ;
      RECT 5.6080 25.0965 5.6340 26.1900 ;
      RECT 5.5000 25.0965 5.5260 26.1900 ;
      RECT 5.3920 25.0965 5.4180 26.1900 ;
      RECT 5.2840 25.0965 5.3100 26.1900 ;
      RECT 5.1760 25.0965 5.2020 26.1900 ;
      RECT 5.0680 25.0965 5.0940 26.1900 ;
      RECT 4.9600 25.0965 4.9860 26.1900 ;
      RECT 4.8520 25.0965 4.8780 26.1900 ;
      RECT 4.7440 25.0965 4.7700 26.1900 ;
      RECT 4.6360 25.0965 4.6620 26.1900 ;
      RECT 4.5280 25.0965 4.5540 26.1900 ;
      RECT 4.4200 25.0965 4.4460 26.1900 ;
      RECT 4.3120 25.0965 4.3380 26.1900 ;
      RECT 4.2040 25.0965 4.2300 26.1900 ;
      RECT 4.0960 25.0965 4.1220 26.1900 ;
      RECT 3.9880 25.0965 4.0140 26.1900 ;
      RECT 3.8800 25.0965 3.9060 26.1900 ;
      RECT 3.7720 25.0965 3.7980 26.1900 ;
      RECT 3.6640 25.0965 3.6900 26.1900 ;
      RECT 3.5560 25.0965 3.5820 26.1900 ;
      RECT 3.4480 25.0965 3.4740 26.1900 ;
      RECT 3.3400 25.0965 3.3660 26.1900 ;
      RECT 3.2320 25.0965 3.2580 26.1900 ;
      RECT 3.1240 25.0965 3.1500 26.1900 ;
      RECT 3.0160 25.0965 3.0420 26.1900 ;
      RECT 2.9080 25.0965 2.9340 26.1900 ;
      RECT 2.8000 25.0965 2.8260 26.1900 ;
      RECT 2.6920 25.0965 2.7180 26.1900 ;
      RECT 2.5840 25.0965 2.6100 26.1900 ;
      RECT 2.4760 25.0965 2.5020 26.1900 ;
      RECT 2.3680 25.0965 2.3940 26.1900 ;
      RECT 2.2600 25.0965 2.2860 26.1900 ;
      RECT 2.1520 25.0965 2.1780 26.1900 ;
      RECT 2.0440 25.0965 2.0700 26.1900 ;
      RECT 1.9360 25.0965 1.9620 26.1900 ;
      RECT 1.8280 25.0965 1.8540 26.1900 ;
      RECT 1.7200 25.0965 1.7460 26.1900 ;
      RECT 1.6120 25.0965 1.6380 26.1900 ;
      RECT 1.5040 25.0965 1.5300 26.1900 ;
      RECT 1.3960 25.0965 1.4220 26.1900 ;
      RECT 1.2880 25.0965 1.3140 26.1900 ;
      RECT 1.1800 25.0965 1.2060 26.1900 ;
      RECT 1.0720 25.0965 1.0980 26.1900 ;
      RECT 0.9640 25.0965 0.9900 26.1900 ;
      RECT 0.8560 25.0965 0.8820 26.1900 ;
      RECT 0.7480 25.0965 0.7740 26.1900 ;
      RECT 0.6400 25.0965 0.6660 26.1900 ;
      RECT 0.5320 25.0965 0.5580 26.1900 ;
      RECT 0.4240 25.0965 0.4500 26.1900 ;
      RECT 0.3160 25.0965 0.3420 26.1900 ;
      RECT 0.2080 25.0965 0.2340 26.1900 ;
      RECT 0.0050 25.0965 0.0900 26.1900 ;
      RECT 0.0000 34.3695 16.5240 34.8105 ;
      RECT 16.4390 26.1570 16.5240 34.8105 ;
      RECT 9.3830 27.6610 16.3210 34.8105 ;
      RECT 10.8410 26.1570 16.3210 34.8105 ;
      RECT 7.2230 34.3620 9.3010 34.8105 ;
      RECT 7.9970 34.3305 9.3010 34.8105 ;
      RECT 0.2030 27.4660 7.1410 34.8105 ;
      RECT 6.8450 26.1570 7.1410 34.8105 ;
      RECT 0.0000 26.1570 0.0850 34.8105 ;
      RECT 7.2230 27.7690 7.8430 34.8105 ;
      RECT 7.9970 34.3260 9.2650 34.8105 ;
      RECT 8.6450 27.5620 9.2650 34.8105 ;
      RECT 8.6360 34.0690 9.2650 34.8105 ;
      RECT 8.4740 34.0690 8.5360 34.8105 ;
      RECT 7.9970 34.0690 8.3830 34.8105 ;
      RECT 9.3830 29.9500 16.3350 34.3040 ;
      RECT 0.1890 29.9500 7.1410 34.3040 ;
      RECT 9.3690 29.9500 16.3350 34.2995 ;
      RECT 0.1890 29.9500 7.1550 34.2995 ;
      RECT 7.2090 29.9500 7.8430 34.2985 ;
      RECT 8.1770 26.8420 8.3470 34.8105 ;
      RECT 8.2850 26.1570 8.3470 34.8105 ;
      RECT 7.4930 26.5780 7.8790 33.9220 ;
      RECT 7.2090 33.8770 7.8930 33.9140 ;
      RECT 8.6310 32.8030 9.2650 33.9110 ;
      RECT 8.1630 33.6130 8.3470 33.8390 ;
      RECT 8.1770 33.0370 8.3610 33.2990 ;
      RECT 7.2090 32.8390 7.8930 33.2990 ;
      RECT 8.1630 32.2990 8.3470 32.7590 ;
      RECT 8.6310 30.2650 9.2650 32.5970 ;
      RECT 7.2090 30.9130 7.8930 32.0570 ;
      RECT 8.1770 30.6430 8.3610 31.9490 ;
      RECT 8.1630 31.2190 8.3610 31.6790 ;
      RECT 8.1630 27.9790 8.3470 31.1390 ;
      RECT 8.1630 27.9790 8.3610 30.5990 ;
      RECT 7.2090 30.3730 7.8930 30.5990 ;
      RECT 8.6450 27.5620 9.3010 29.9180 ;
      RECT 8.6310 27.4390 9.2470 29.2250 ;
      RECT 7.2230 28.4110 7.8930 28.7810 ;
      RECT 8.1770 27.7090 8.3610 27.8990 ;
      RECT 7.2770 27.6730 7.8930 27.8630 ;
      RECT 8.1630 27.5650 8.3470 27.7010 ;
      RECT 7.2770 26.9230 7.8790 33.9220 ;
      RECT 8.1770 27.4390 8.3610 27.6650 ;
      RECT 9.5450 27.4690 16.3210 34.8105 ;
      RECT 10.6250 27.4660 16.3210 34.8105 ;
      RECT 9.3830 26.1570 9.4630 34.8105 ;
      RECT 7.2230 26.8420 7.4110 27.6560 ;
      RECT 9.3830 26.1570 9.6790 27.5600 ;
      RECT 9.3830 27.2740 10.5430 27.5600 ;
      RECT 10.6250 26.1570 10.7590 34.8105 ;
      RECT 5.9810 27.0850 6.7630 34.8105 ;
      RECT 0.2030 26.1570 5.8990 34.8105 ;
      RECT 8.6450 26.9230 9.2470 34.8105 ;
      RECT 8.6810 26.3335 9.3010 27.4070 ;
      RECT 9.3830 27.2740 10.7590 27.3680 ;
      RECT 10.4090 26.1570 16.3210 27.3650 ;
      RECT 6.6290 26.1570 7.1410 27.3650 ;
      RECT 8.1630 27.2950 8.3610 27.3590 ;
      RECT 8.1630 27.1690 8.3470 27.3590 ;
      RECT 10.1930 26.8900 16.3210 27.3650 ;
      RECT 9.3830 26.9230 10.1110 27.5600 ;
      RECT 8.1770 26.8990 8.3610 27.1610 ;
      RECT 0.2030 26.8900 6.5470 27.3650 ;
      RECT 6.4130 26.1570 6.5470 34.8105 ;
      RECT 9.9770 26.1570 10.3270 27.0290 ;
      RECT 9.3830 26.8420 9.8950 27.5600 ;
      RECT 9.7610 26.1570 9.8950 34.8105 ;
      RECT 6.1970 26.8420 6.5470 34.8105 ;
      RECT 0.2030 26.1570 6.1150 27.3650 ;
      RECT 8.1770 26.1570 8.2030 34.8105 ;
      RECT 7.3130 26.1570 7.4110 34.8105 ;
      RECT 6.1970 26.1570 6.3310 34.8105 ;
      RECT 9.7610 26.1570 10.3270 26.7920 ;
      RECT 8.6450 26.1570 9.2470 26.7920 ;
      RECT 7.3130 26.1570 7.8430 26.7920 ;
      RECT 6.4130 26.1570 7.1410 26.7920 ;
      RECT 9.7610 26.1570 16.3210 26.7890 ;
      RECT 0.2030 26.1570 6.3310 26.7890 ;
      RECT 8.6310 26.6290 9.3010 26.7830 ;
      RECT 9.3830 26.1570 16.3210 26.5250 ;
      RECT 8.1770 26.1570 8.3470 26.5250 ;
      RECT 7.2230 26.1570 7.8430 26.5250 ;
      RECT 0.2030 26.1570 7.1410 26.5250 ;
      RECT 7.9970 26.1570 8.3470 26.4220 ;
      RECT 8.6360 26.1570 9.2470 26.3220 ;
      RECT 7.9970 26.1570 8.3830 26.3220 ;
      RECT 9.7650 26.1305 9.7830 34.8105 ;
      RECT 9.6570 26.1305 9.6750 34.8105 ;
      RECT 6.8490 26.1430 6.8670 34.8105 ;
      RECT 6.7410 26.1430 6.7590 34.8105 ;
      RECT 6.6330 26.1430 6.6510 34.8105 ;
      RECT 6.5250 26.1430 6.5430 34.8105 ;
      RECT 6.4170 26.1305 6.4350 34.8105 ;
      RECT 6.3090 26.1305 6.3270 34.8105 ;
      RECT 6.2010 26.1430 6.2190 34.8105 ;
      RECT 6.0930 26.1430 6.1110 34.8105 ;
      RECT 5.9850 26.1430 6.0030 34.8105 ;
      RECT 5.8770 26.1430 5.8950 34.8105 ;
      RECT 8.4740 26.1570 8.5360 26.3220 ;
        RECT 8.6410 34.3035 8.7690 35.3970 ;
        RECT 8.6270 34.9690 8.7690 35.2915 ;
        RECT 8.4790 34.6960 8.5410 35.3970 ;
        RECT 8.4650 35.0055 8.5410 35.1590 ;
        RECT 8.4790 34.3035 8.5050 35.3970 ;
        RECT 8.4790 34.4245 8.5190 34.6640 ;
        RECT 8.4790 34.3035 8.5410 34.3925 ;
        RECT 8.1820 34.7540 8.3880 35.3970 ;
        RECT 8.3620 34.3035 8.3880 35.3970 ;
        RECT 8.1820 35.0310 8.4020 35.2890 ;
        RECT 8.1820 34.3035 8.2800 35.3970 ;
        RECT 7.7650 34.3035 7.8480 35.3970 ;
        RECT 7.7650 34.3920 7.8620 35.3275 ;
        RECT 16.4440 34.3035 16.5290 35.3970 ;
        RECT 16.3000 34.3035 16.3260 35.3970 ;
        RECT 16.1920 34.3035 16.2180 35.3970 ;
        RECT 16.0840 34.3035 16.1100 35.3970 ;
        RECT 15.9760 34.3035 16.0020 35.3970 ;
        RECT 15.8680 34.3035 15.8940 35.3970 ;
        RECT 15.7600 34.3035 15.7860 35.3970 ;
        RECT 15.6520 34.3035 15.6780 35.3970 ;
        RECT 15.5440 34.3035 15.5700 35.3970 ;
        RECT 15.4360 34.3035 15.4620 35.3970 ;
        RECT 15.3280 34.3035 15.3540 35.3970 ;
        RECT 15.2200 34.3035 15.2460 35.3970 ;
        RECT 15.1120 34.3035 15.1380 35.3970 ;
        RECT 15.0040 34.3035 15.0300 35.3970 ;
        RECT 14.8960 34.3035 14.9220 35.3970 ;
        RECT 14.7880 34.3035 14.8140 35.3970 ;
        RECT 14.6800 34.3035 14.7060 35.3970 ;
        RECT 14.5720 34.3035 14.5980 35.3970 ;
        RECT 14.4640 34.3035 14.4900 35.3970 ;
        RECT 14.3560 34.3035 14.3820 35.3970 ;
        RECT 14.2480 34.3035 14.2740 35.3970 ;
        RECT 14.1400 34.3035 14.1660 35.3970 ;
        RECT 14.0320 34.3035 14.0580 35.3970 ;
        RECT 13.9240 34.3035 13.9500 35.3970 ;
        RECT 13.8160 34.3035 13.8420 35.3970 ;
        RECT 13.7080 34.3035 13.7340 35.3970 ;
        RECT 13.6000 34.3035 13.6260 35.3970 ;
        RECT 13.4920 34.3035 13.5180 35.3970 ;
        RECT 13.3840 34.3035 13.4100 35.3970 ;
        RECT 13.2760 34.3035 13.3020 35.3970 ;
        RECT 13.1680 34.3035 13.1940 35.3970 ;
        RECT 13.0600 34.3035 13.0860 35.3970 ;
        RECT 12.9520 34.3035 12.9780 35.3970 ;
        RECT 12.8440 34.3035 12.8700 35.3970 ;
        RECT 12.7360 34.3035 12.7620 35.3970 ;
        RECT 12.6280 34.3035 12.6540 35.3970 ;
        RECT 12.5200 34.3035 12.5460 35.3970 ;
        RECT 12.4120 34.3035 12.4380 35.3970 ;
        RECT 12.3040 34.3035 12.3300 35.3970 ;
        RECT 12.1960 34.3035 12.2220 35.3970 ;
        RECT 12.0880 34.3035 12.1140 35.3970 ;
        RECT 11.9800 34.3035 12.0060 35.3970 ;
        RECT 11.8720 34.3035 11.8980 35.3970 ;
        RECT 11.7640 34.3035 11.7900 35.3970 ;
        RECT 11.6560 34.3035 11.6820 35.3970 ;
        RECT 11.5480 34.3035 11.5740 35.3970 ;
        RECT 11.4400 34.3035 11.4660 35.3970 ;
        RECT 11.3320 34.3035 11.3580 35.3970 ;
        RECT 11.2240 34.3035 11.2500 35.3970 ;
        RECT 11.1160 34.3035 11.1420 35.3970 ;
        RECT 11.0080 34.3035 11.0340 35.3970 ;
        RECT 10.9000 34.3035 10.9260 35.3970 ;
        RECT 10.7920 34.3035 10.8180 35.3970 ;
        RECT 10.6840 34.3035 10.7100 35.3970 ;
        RECT 10.5760 34.3035 10.6020 35.3970 ;
        RECT 10.4680 34.3035 10.4940 35.3970 ;
        RECT 10.3600 34.3035 10.3860 35.3970 ;
        RECT 10.2520 34.3035 10.2780 35.3970 ;
        RECT 10.1440 34.3035 10.1700 35.3970 ;
        RECT 10.0360 34.3035 10.0620 35.3970 ;
        RECT 9.9280 34.3035 9.9540 35.3970 ;
        RECT 9.8200 34.3035 9.8460 35.3970 ;
        RECT 9.7120 34.3035 9.7380 35.3970 ;
        RECT 9.6040 34.3035 9.6300 35.3970 ;
        RECT 9.4960 34.3035 9.5220 35.3970 ;
        RECT 9.3880 34.3035 9.4140 35.3970 ;
        RECT 9.1750 34.3035 9.2520 35.3970 ;
        RECT 7.2820 34.3035 7.3590 35.3970 ;
        RECT 7.1200 34.3035 7.1460 35.3970 ;
        RECT 7.0120 34.3035 7.0380 35.3970 ;
        RECT 6.9040 34.3035 6.9300 35.3970 ;
        RECT 6.7960 34.3035 6.8220 35.3970 ;
        RECT 6.6880 34.3035 6.7140 35.3970 ;
        RECT 6.5800 34.3035 6.6060 35.3970 ;
        RECT 6.4720 34.3035 6.4980 35.3970 ;
        RECT 6.3640 34.3035 6.3900 35.3970 ;
        RECT 6.2560 34.3035 6.2820 35.3970 ;
        RECT 6.1480 34.3035 6.1740 35.3970 ;
        RECT 6.0400 34.3035 6.0660 35.3970 ;
        RECT 5.9320 34.3035 5.9580 35.3970 ;
        RECT 5.8240 34.3035 5.8500 35.3970 ;
        RECT 5.7160 34.3035 5.7420 35.3970 ;
        RECT 5.6080 34.3035 5.6340 35.3970 ;
        RECT 5.5000 34.3035 5.5260 35.3970 ;
        RECT 5.3920 34.3035 5.4180 35.3970 ;
        RECT 5.2840 34.3035 5.3100 35.3970 ;
        RECT 5.1760 34.3035 5.2020 35.3970 ;
        RECT 5.0680 34.3035 5.0940 35.3970 ;
        RECT 4.9600 34.3035 4.9860 35.3970 ;
        RECT 4.8520 34.3035 4.8780 35.3970 ;
        RECT 4.7440 34.3035 4.7700 35.3970 ;
        RECT 4.6360 34.3035 4.6620 35.3970 ;
        RECT 4.5280 34.3035 4.5540 35.3970 ;
        RECT 4.4200 34.3035 4.4460 35.3970 ;
        RECT 4.3120 34.3035 4.3380 35.3970 ;
        RECT 4.2040 34.3035 4.2300 35.3970 ;
        RECT 4.0960 34.3035 4.1220 35.3970 ;
        RECT 3.9880 34.3035 4.0140 35.3970 ;
        RECT 3.8800 34.3035 3.9060 35.3970 ;
        RECT 3.7720 34.3035 3.7980 35.3970 ;
        RECT 3.6640 34.3035 3.6900 35.3970 ;
        RECT 3.5560 34.3035 3.5820 35.3970 ;
        RECT 3.4480 34.3035 3.4740 35.3970 ;
        RECT 3.3400 34.3035 3.3660 35.3970 ;
        RECT 3.2320 34.3035 3.2580 35.3970 ;
        RECT 3.1240 34.3035 3.1500 35.3970 ;
        RECT 3.0160 34.3035 3.0420 35.3970 ;
        RECT 2.9080 34.3035 2.9340 35.3970 ;
        RECT 2.8000 34.3035 2.8260 35.3970 ;
        RECT 2.6920 34.3035 2.7180 35.3970 ;
        RECT 2.5840 34.3035 2.6100 35.3970 ;
        RECT 2.4760 34.3035 2.5020 35.3970 ;
        RECT 2.3680 34.3035 2.3940 35.3970 ;
        RECT 2.2600 34.3035 2.2860 35.3970 ;
        RECT 2.1520 34.3035 2.1780 35.3970 ;
        RECT 2.0440 34.3035 2.0700 35.3970 ;
        RECT 1.9360 34.3035 1.9620 35.3970 ;
        RECT 1.8280 34.3035 1.8540 35.3970 ;
        RECT 1.7200 34.3035 1.7460 35.3970 ;
        RECT 1.6120 34.3035 1.6380 35.3970 ;
        RECT 1.5040 34.3035 1.5300 35.3970 ;
        RECT 1.3960 34.3035 1.4220 35.3970 ;
        RECT 1.2880 34.3035 1.3140 35.3970 ;
        RECT 1.1800 34.3035 1.2060 35.3970 ;
        RECT 1.0720 34.3035 1.0980 35.3970 ;
        RECT 0.9640 34.3035 0.9900 35.3970 ;
        RECT 0.8560 34.3035 0.8820 35.3970 ;
        RECT 0.7480 34.3035 0.7740 35.3970 ;
        RECT 0.6400 34.3035 0.6660 35.3970 ;
        RECT 0.5320 34.3035 0.5580 35.3970 ;
        RECT 0.4240 34.3035 0.4500 35.3970 ;
        RECT 0.3160 34.3035 0.3420 35.3970 ;
        RECT 0.2080 34.3035 0.2340 35.3970 ;
        RECT 0.0050 34.3035 0.0900 35.3970 ;
        RECT 8.6410 35.3835 8.7690 36.4770 ;
        RECT 8.6270 36.0490 8.7690 36.3715 ;
        RECT 8.4790 35.7760 8.5410 36.4770 ;
        RECT 8.4650 36.0855 8.5410 36.2390 ;
        RECT 8.4790 35.3835 8.5050 36.4770 ;
        RECT 8.4790 35.5045 8.5190 35.7440 ;
        RECT 8.4790 35.3835 8.5410 35.4725 ;
        RECT 8.1820 35.8340 8.3880 36.4770 ;
        RECT 8.3620 35.3835 8.3880 36.4770 ;
        RECT 8.1820 36.1110 8.4020 36.3690 ;
        RECT 8.1820 35.3835 8.2800 36.4770 ;
        RECT 7.7650 35.3835 7.8480 36.4770 ;
        RECT 7.7650 35.4720 7.8620 36.4075 ;
        RECT 16.4440 35.3835 16.5290 36.4770 ;
        RECT 16.3000 35.3835 16.3260 36.4770 ;
        RECT 16.1920 35.3835 16.2180 36.4770 ;
        RECT 16.0840 35.3835 16.1100 36.4770 ;
        RECT 15.9760 35.3835 16.0020 36.4770 ;
        RECT 15.8680 35.3835 15.8940 36.4770 ;
        RECT 15.7600 35.3835 15.7860 36.4770 ;
        RECT 15.6520 35.3835 15.6780 36.4770 ;
        RECT 15.5440 35.3835 15.5700 36.4770 ;
        RECT 15.4360 35.3835 15.4620 36.4770 ;
        RECT 15.3280 35.3835 15.3540 36.4770 ;
        RECT 15.2200 35.3835 15.2460 36.4770 ;
        RECT 15.1120 35.3835 15.1380 36.4770 ;
        RECT 15.0040 35.3835 15.0300 36.4770 ;
        RECT 14.8960 35.3835 14.9220 36.4770 ;
        RECT 14.7880 35.3835 14.8140 36.4770 ;
        RECT 14.6800 35.3835 14.7060 36.4770 ;
        RECT 14.5720 35.3835 14.5980 36.4770 ;
        RECT 14.4640 35.3835 14.4900 36.4770 ;
        RECT 14.3560 35.3835 14.3820 36.4770 ;
        RECT 14.2480 35.3835 14.2740 36.4770 ;
        RECT 14.1400 35.3835 14.1660 36.4770 ;
        RECT 14.0320 35.3835 14.0580 36.4770 ;
        RECT 13.9240 35.3835 13.9500 36.4770 ;
        RECT 13.8160 35.3835 13.8420 36.4770 ;
        RECT 13.7080 35.3835 13.7340 36.4770 ;
        RECT 13.6000 35.3835 13.6260 36.4770 ;
        RECT 13.4920 35.3835 13.5180 36.4770 ;
        RECT 13.3840 35.3835 13.4100 36.4770 ;
        RECT 13.2760 35.3835 13.3020 36.4770 ;
        RECT 13.1680 35.3835 13.1940 36.4770 ;
        RECT 13.0600 35.3835 13.0860 36.4770 ;
        RECT 12.9520 35.3835 12.9780 36.4770 ;
        RECT 12.8440 35.3835 12.8700 36.4770 ;
        RECT 12.7360 35.3835 12.7620 36.4770 ;
        RECT 12.6280 35.3835 12.6540 36.4770 ;
        RECT 12.5200 35.3835 12.5460 36.4770 ;
        RECT 12.4120 35.3835 12.4380 36.4770 ;
        RECT 12.3040 35.3835 12.3300 36.4770 ;
        RECT 12.1960 35.3835 12.2220 36.4770 ;
        RECT 12.0880 35.3835 12.1140 36.4770 ;
        RECT 11.9800 35.3835 12.0060 36.4770 ;
        RECT 11.8720 35.3835 11.8980 36.4770 ;
        RECT 11.7640 35.3835 11.7900 36.4770 ;
        RECT 11.6560 35.3835 11.6820 36.4770 ;
        RECT 11.5480 35.3835 11.5740 36.4770 ;
        RECT 11.4400 35.3835 11.4660 36.4770 ;
        RECT 11.3320 35.3835 11.3580 36.4770 ;
        RECT 11.2240 35.3835 11.2500 36.4770 ;
        RECT 11.1160 35.3835 11.1420 36.4770 ;
        RECT 11.0080 35.3835 11.0340 36.4770 ;
        RECT 10.9000 35.3835 10.9260 36.4770 ;
        RECT 10.7920 35.3835 10.8180 36.4770 ;
        RECT 10.6840 35.3835 10.7100 36.4770 ;
        RECT 10.5760 35.3835 10.6020 36.4770 ;
        RECT 10.4680 35.3835 10.4940 36.4770 ;
        RECT 10.3600 35.3835 10.3860 36.4770 ;
        RECT 10.2520 35.3835 10.2780 36.4770 ;
        RECT 10.1440 35.3835 10.1700 36.4770 ;
        RECT 10.0360 35.3835 10.0620 36.4770 ;
        RECT 9.9280 35.3835 9.9540 36.4770 ;
        RECT 9.8200 35.3835 9.8460 36.4770 ;
        RECT 9.7120 35.3835 9.7380 36.4770 ;
        RECT 9.6040 35.3835 9.6300 36.4770 ;
        RECT 9.4960 35.3835 9.5220 36.4770 ;
        RECT 9.3880 35.3835 9.4140 36.4770 ;
        RECT 9.1750 35.3835 9.2520 36.4770 ;
        RECT 7.2820 35.3835 7.3590 36.4770 ;
        RECT 7.1200 35.3835 7.1460 36.4770 ;
        RECT 7.0120 35.3835 7.0380 36.4770 ;
        RECT 6.9040 35.3835 6.9300 36.4770 ;
        RECT 6.7960 35.3835 6.8220 36.4770 ;
        RECT 6.6880 35.3835 6.7140 36.4770 ;
        RECT 6.5800 35.3835 6.6060 36.4770 ;
        RECT 6.4720 35.3835 6.4980 36.4770 ;
        RECT 6.3640 35.3835 6.3900 36.4770 ;
        RECT 6.2560 35.3835 6.2820 36.4770 ;
        RECT 6.1480 35.3835 6.1740 36.4770 ;
        RECT 6.0400 35.3835 6.0660 36.4770 ;
        RECT 5.9320 35.3835 5.9580 36.4770 ;
        RECT 5.8240 35.3835 5.8500 36.4770 ;
        RECT 5.7160 35.3835 5.7420 36.4770 ;
        RECT 5.6080 35.3835 5.6340 36.4770 ;
        RECT 5.5000 35.3835 5.5260 36.4770 ;
        RECT 5.3920 35.3835 5.4180 36.4770 ;
        RECT 5.2840 35.3835 5.3100 36.4770 ;
        RECT 5.1760 35.3835 5.2020 36.4770 ;
        RECT 5.0680 35.3835 5.0940 36.4770 ;
        RECT 4.9600 35.3835 4.9860 36.4770 ;
        RECT 4.8520 35.3835 4.8780 36.4770 ;
        RECT 4.7440 35.3835 4.7700 36.4770 ;
        RECT 4.6360 35.3835 4.6620 36.4770 ;
        RECT 4.5280 35.3835 4.5540 36.4770 ;
        RECT 4.4200 35.3835 4.4460 36.4770 ;
        RECT 4.3120 35.3835 4.3380 36.4770 ;
        RECT 4.2040 35.3835 4.2300 36.4770 ;
        RECT 4.0960 35.3835 4.1220 36.4770 ;
        RECT 3.9880 35.3835 4.0140 36.4770 ;
        RECT 3.8800 35.3835 3.9060 36.4770 ;
        RECT 3.7720 35.3835 3.7980 36.4770 ;
        RECT 3.6640 35.3835 3.6900 36.4770 ;
        RECT 3.5560 35.3835 3.5820 36.4770 ;
        RECT 3.4480 35.3835 3.4740 36.4770 ;
        RECT 3.3400 35.3835 3.3660 36.4770 ;
        RECT 3.2320 35.3835 3.2580 36.4770 ;
        RECT 3.1240 35.3835 3.1500 36.4770 ;
        RECT 3.0160 35.3835 3.0420 36.4770 ;
        RECT 2.9080 35.3835 2.9340 36.4770 ;
        RECT 2.8000 35.3835 2.8260 36.4770 ;
        RECT 2.6920 35.3835 2.7180 36.4770 ;
        RECT 2.5840 35.3835 2.6100 36.4770 ;
        RECT 2.4760 35.3835 2.5020 36.4770 ;
        RECT 2.3680 35.3835 2.3940 36.4770 ;
        RECT 2.2600 35.3835 2.2860 36.4770 ;
        RECT 2.1520 35.3835 2.1780 36.4770 ;
        RECT 2.0440 35.3835 2.0700 36.4770 ;
        RECT 1.9360 35.3835 1.9620 36.4770 ;
        RECT 1.8280 35.3835 1.8540 36.4770 ;
        RECT 1.7200 35.3835 1.7460 36.4770 ;
        RECT 1.6120 35.3835 1.6380 36.4770 ;
        RECT 1.5040 35.3835 1.5300 36.4770 ;
        RECT 1.3960 35.3835 1.4220 36.4770 ;
        RECT 1.2880 35.3835 1.3140 36.4770 ;
        RECT 1.1800 35.3835 1.2060 36.4770 ;
        RECT 1.0720 35.3835 1.0980 36.4770 ;
        RECT 0.9640 35.3835 0.9900 36.4770 ;
        RECT 0.8560 35.3835 0.8820 36.4770 ;
        RECT 0.7480 35.3835 0.7740 36.4770 ;
        RECT 0.6400 35.3835 0.6660 36.4770 ;
        RECT 0.5320 35.3835 0.5580 36.4770 ;
        RECT 0.4240 35.3835 0.4500 36.4770 ;
        RECT 0.3160 35.3835 0.3420 36.4770 ;
        RECT 0.2080 35.3835 0.2340 36.4770 ;
        RECT 0.0050 35.3835 0.0900 36.4770 ;
        RECT 8.6410 36.4635 8.7690 37.5570 ;
        RECT 8.6270 37.1290 8.7690 37.4515 ;
        RECT 8.4790 36.8560 8.5410 37.5570 ;
        RECT 8.4650 37.1655 8.5410 37.3190 ;
        RECT 8.4790 36.4635 8.5050 37.5570 ;
        RECT 8.4790 36.5845 8.5190 36.8240 ;
        RECT 8.4790 36.4635 8.5410 36.5525 ;
        RECT 8.1820 36.9140 8.3880 37.5570 ;
        RECT 8.3620 36.4635 8.3880 37.5570 ;
        RECT 8.1820 37.1910 8.4020 37.4490 ;
        RECT 8.1820 36.4635 8.2800 37.5570 ;
        RECT 7.7650 36.4635 7.8480 37.5570 ;
        RECT 7.7650 36.5520 7.8620 37.4875 ;
        RECT 16.4440 36.4635 16.5290 37.5570 ;
        RECT 16.3000 36.4635 16.3260 37.5570 ;
        RECT 16.1920 36.4635 16.2180 37.5570 ;
        RECT 16.0840 36.4635 16.1100 37.5570 ;
        RECT 15.9760 36.4635 16.0020 37.5570 ;
        RECT 15.8680 36.4635 15.8940 37.5570 ;
        RECT 15.7600 36.4635 15.7860 37.5570 ;
        RECT 15.6520 36.4635 15.6780 37.5570 ;
        RECT 15.5440 36.4635 15.5700 37.5570 ;
        RECT 15.4360 36.4635 15.4620 37.5570 ;
        RECT 15.3280 36.4635 15.3540 37.5570 ;
        RECT 15.2200 36.4635 15.2460 37.5570 ;
        RECT 15.1120 36.4635 15.1380 37.5570 ;
        RECT 15.0040 36.4635 15.0300 37.5570 ;
        RECT 14.8960 36.4635 14.9220 37.5570 ;
        RECT 14.7880 36.4635 14.8140 37.5570 ;
        RECT 14.6800 36.4635 14.7060 37.5570 ;
        RECT 14.5720 36.4635 14.5980 37.5570 ;
        RECT 14.4640 36.4635 14.4900 37.5570 ;
        RECT 14.3560 36.4635 14.3820 37.5570 ;
        RECT 14.2480 36.4635 14.2740 37.5570 ;
        RECT 14.1400 36.4635 14.1660 37.5570 ;
        RECT 14.0320 36.4635 14.0580 37.5570 ;
        RECT 13.9240 36.4635 13.9500 37.5570 ;
        RECT 13.8160 36.4635 13.8420 37.5570 ;
        RECT 13.7080 36.4635 13.7340 37.5570 ;
        RECT 13.6000 36.4635 13.6260 37.5570 ;
        RECT 13.4920 36.4635 13.5180 37.5570 ;
        RECT 13.3840 36.4635 13.4100 37.5570 ;
        RECT 13.2760 36.4635 13.3020 37.5570 ;
        RECT 13.1680 36.4635 13.1940 37.5570 ;
        RECT 13.0600 36.4635 13.0860 37.5570 ;
        RECT 12.9520 36.4635 12.9780 37.5570 ;
        RECT 12.8440 36.4635 12.8700 37.5570 ;
        RECT 12.7360 36.4635 12.7620 37.5570 ;
        RECT 12.6280 36.4635 12.6540 37.5570 ;
        RECT 12.5200 36.4635 12.5460 37.5570 ;
        RECT 12.4120 36.4635 12.4380 37.5570 ;
        RECT 12.3040 36.4635 12.3300 37.5570 ;
        RECT 12.1960 36.4635 12.2220 37.5570 ;
        RECT 12.0880 36.4635 12.1140 37.5570 ;
        RECT 11.9800 36.4635 12.0060 37.5570 ;
        RECT 11.8720 36.4635 11.8980 37.5570 ;
        RECT 11.7640 36.4635 11.7900 37.5570 ;
        RECT 11.6560 36.4635 11.6820 37.5570 ;
        RECT 11.5480 36.4635 11.5740 37.5570 ;
        RECT 11.4400 36.4635 11.4660 37.5570 ;
        RECT 11.3320 36.4635 11.3580 37.5570 ;
        RECT 11.2240 36.4635 11.2500 37.5570 ;
        RECT 11.1160 36.4635 11.1420 37.5570 ;
        RECT 11.0080 36.4635 11.0340 37.5570 ;
        RECT 10.9000 36.4635 10.9260 37.5570 ;
        RECT 10.7920 36.4635 10.8180 37.5570 ;
        RECT 10.6840 36.4635 10.7100 37.5570 ;
        RECT 10.5760 36.4635 10.6020 37.5570 ;
        RECT 10.4680 36.4635 10.4940 37.5570 ;
        RECT 10.3600 36.4635 10.3860 37.5570 ;
        RECT 10.2520 36.4635 10.2780 37.5570 ;
        RECT 10.1440 36.4635 10.1700 37.5570 ;
        RECT 10.0360 36.4635 10.0620 37.5570 ;
        RECT 9.9280 36.4635 9.9540 37.5570 ;
        RECT 9.8200 36.4635 9.8460 37.5570 ;
        RECT 9.7120 36.4635 9.7380 37.5570 ;
        RECT 9.6040 36.4635 9.6300 37.5570 ;
        RECT 9.4960 36.4635 9.5220 37.5570 ;
        RECT 9.3880 36.4635 9.4140 37.5570 ;
        RECT 9.1750 36.4635 9.2520 37.5570 ;
        RECT 7.2820 36.4635 7.3590 37.5570 ;
        RECT 7.1200 36.4635 7.1460 37.5570 ;
        RECT 7.0120 36.4635 7.0380 37.5570 ;
        RECT 6.9040 36.4635 6.9300 37.5570 ;
        RECT 6.7960 36.4635 6.8220 37.5570 ;
        RECT 6.6880 36.4635 6.7140 37.5570 ;
        RECT 6.5800 36.4635 6.6060 37.5570 ;
        RECT 6.4720 36.4635 6.4980 37.5570 ;
        RECT 6.3640 36.4635 6.3900 37.5570 ;
        RECT 6.2560 36.4635 6.2820 37.5570 ;
        RECT 6.1480 36.4635 6.1740 37.5570 ;
        RECT 6.0400 36.4635 6.0660 37.5570 ;
        RECT 5.9320 36.4635 5.9580 37.5570 ;
        RECT 5.8240 36.4635 5.8500 37.5570 ;
        RECT 5.7160 36.4635 5.7420 37.5570 ;
        RECT 5.6080 36.4635 5.6340 37.5570 ;
        RECT 5.5000 36.4635 5.5260 37.5570 ;
        RECT 5.3920 36.4635 5.4180 37.5570 ;
        RECT 5.2840 36.4635 5.3100 37.5570 ;
        RECT 5.1760 36.4635 5.2020 37.5570 ;
        RECT 5.0680 36.4635 5.0940 37.5570 ;
        RECT 4.9600 36.4635 4.9860 37.5570 ;
        RECT 4.8520 36.4635 4.8780 37.5570 ;
        RECT 4.7440 36.4635 4.7700 37.5570 ;
        RECT 4.6360 36.4635 4.6620 37.5570 ;
        RECT 4.5280 36.4635 4.5540 37.5570 ;
        RECT 4.4200 36.4635 4.4460 37.5570 ;
        RECT 4.3120 36.4635 4.3380 37.5570 ;
        RECT 4.2040 36.4635 4.2300 37.5570 ;
        RECT 4.0960 36.4635 4.1220 37.5570 ;
        RECT 3.9880 36.4635 4.0140 37.5570 ;
        RECT 3.8800 36.4635 3.9060 37.5570 ;
        RECT 3.7720 36.4635 3.7980 37.5570 ;
        RECT 3.6640 36.4635 3.6900 37.5570 ;
        RECT 3.5560 36.4635 3.5820 37.5570 ;
        RECT 3.4480 36.4635 3.4740 37.5570 ;
        RECT 3.3400 36.4635 3.3660 37.5570 ;
        RECT 3.2320 36.4635 3.2580 37.5570 ;
        RECT 3.1240 36.4635 3.1500 37.5570 ;
        RECT 3.0160 36.4635 3.0420 37.5570 ;
        RECT 2.9080 36.4635 2.9340 37.5570 ;
        RECT 2.8000 36.4635 2.8260 37.5570 ;
        RECT 2.6920 36.4635 2.7180 37.5570 ;
        RECT 2.5840 36.4635 2.6100 37.5570 ;
        RECT 2.4760 36.4635 2.5020 37.5570 ;
        RECT 2.3680 36.4635 2.3940 37.5570 ;
        RECT 2.2600 36.4635 2.2860 37.5570 ;
        RECT 2.1520 36.4635 2.1780 37.5570 ;
        RECT 2.0440 36.4635 2.0700 37.5570 ;
        RECT 1.9360 36.4635 1.9620 37.5570 ;
        RECT 1.8280 36.4635 1.8540 37.5570 ;
        RECT 1.7200 36.4635 1.7460 37.5570 ;
        RECT 1.6120 36.4635 1.6380 37.5570 ;
        RECT 1.5040 36.4635 1.5300 37.5570 ;
        RECT 1.3960 36.4635 1.4220 37.5570 ;
        RECT 1.2880 36.4635 1.3140 37.5570 ;
        RECT 1.1800 36.4635 1.2060 37.5570 ;
        RECT 1.0720 36.4635 1.0980 37.5570 ;
        RECT 0.9640 36.4635 0.9900 37.5570 ;
        RECT 0.8560 36.4635 0.8820 37.5570 ;
        RECT 0.7480 36.4635 0.7740 37.5570 ;
        RECT 0.6400 36.4635 0.6660 37.5570 ;
        RECT 0.5320 36.4635 0.5580 37.5570 ;
        RECT 0.4240 36.4635 0.4500 37.5570 ;
        RECT 0.3160 36.4635 0.3420 37.5570 ;
        RECT 0.2080 36.4635 0.2340 37.5570 ;
        RECT 0.0050 36.4635 0.0900 37.5570 ;
        RECT 8.6410 37.5435 8.7690 38.6370 ;
        RECT 8.6270 38.2090 8.7690 38.5315 ;
        RECT 8.4790 37.9360 8.5410 38.6370 ;
        RECT 8.4650 38.2455 8.5410 38.3990 ;
        RECT 8.4790 37.5435 8.5050 38.6370 ;
        RECT 8.4790 37.6645 8.5190 37.9040 ;
        RECT 8.4790 37.5435 8.5410 37.6325 ;
        RECT 8.1820 37.9940 8.3880 38.6370 ;
        RECT 8.3620 37.5435 8.3880 38.6370 ;
        RECT 8.1820 38.2710 8.4020 38.5290 ;
        RECT 8.1820 37.5435 8.2800 38.6370 ;
        RECT 7.7650 37.5435 7.8480 38.6370 ;
        RECT 7.7650 37.6320 7.8620 38.5675 ;
        RECT 16.4440 37.5435 16.5290 38.6370 ;
        RECT 16.3000 37.5435 16.3260 38.6370 ;
        RECT 16.1920 37.5435 16.2180 38.6370 ;
        RECT 16.0840 37.5435 16.1100 38.6370 ;
        RECT 15.9760 37.5435 16.0020 38.6370 ;
        RECT 15.8680 37.5435 15.8940 38.6370 ;
        RECT 15.7600 37.5435 15.7860 38.6370 ;
        RECT 15.6520 37.5435 15.6780 38.6370 ;
        RECT 15.5440 37.5435 15.5700 38.6370 ;
        RECT 15.4360 37.5435 15.4620 38.6370 ;
        RECT 15.3280 37.5435 15.3540 38.6370 ;
        RECT 15.2200 37.5435 15.2460 38.6370 ;
        RECT 15.1120 37.5435 15.1380 38.6370 ;
        RECT 15.0040 37.5435 15.0300 38.6370 ;
        RECT 14.8960 37.5435 14.9220 38.6370 ;
        RECT 14.7880 37.5435 14.8140 38.6370 ;
        RECT 14.6800 37.5435 14.7060 38.6370 ;
        RECT 14.5720 37.5435 14.5980 38.6370 ;
        RECT 14.4640 37.5435 14.4900 38.6370 ;
        RECT 14.3560 37.5435 14.3820 38.6370 ;
        RECT 14.2480 37.5435 14.2740 38.6370 ;
        RECT 14.1400 37.5435 14.1660 38.6370 ;
        RECT 14.0320 37.5435 14.0580 38.6370 ;
        RECT 13.9240 37.5435 13.9500 38.6370 ;
        RECT 13.8160 37.5435 13.8420 38.6370 ;
        RECT 13.7080 37.5435 13.7340 38.6370 ;
        RECT 13.6000 37.5435 13.6260 38.6370 ;
        RECT 13.4920 37.5435 13.5180 38.6370 ;
        RECT 13.3840 37.5435 13.4100 38.6370 ;
        RECT 13.2760 37.5435 13.3020 38.6370 ;
        RECT 13.1680 37.5435 13.1940 38.6370 ;
        RECT 13.0600 37.5435 13.0860 38.6370 ;
        RECT 12.9520 37.5435 12.9780 38.6370 ;
        RECT 12.8440 37.5435 12.8700 38.6370 ;
        RECT 12.7360 37.5435 12.7620 38.6370 ;
        RECT 12.6280 37.5435 12.6540 38.6370 ;
        RECT 12.5200 37.5435 12.5460 38.6370 ;
        RECT 12.4120 37.5435 12.4380 38.6370 ;
        RECT 12.3040 37.5435 12.3300 38.6370 ;
        RECT 12.1960 37.5435 12.2220 38.6370 ;
        RECT 12.0880 37.5435 12.1140 38.6370 ;
        RECT 11.9800 37.5435 12.0060 38.6370 ;
        RECT 11.8720 37.5435 11.8980 38.6370 ;
        RECT 11.7640 37.5435 11.7900 38.6370 ;
        RECT 11.6560 37.5435 11.6820 38.6370 ;
        RECT 11.5480 37.5435 11.5740 38.6370 ;
        RECT 11.4400 37.5435 11.4660 38.6370 ;
        RECT 11.3320 37.5435 11.3580 38.6370 ;
        RECT 11.2240 37.5435 11.2500 38.6370 ;
        RECT 11.1160 37.5435 11.1420 38.6370 ;
        RECT 11.0080 37.5435 11.0340 38.6370 ;
        RECT 10.9000 37.5435 10.9260 38.6370 ;
        RECT 10.7920 37.5435 10.8180 38.6370 ;
        RECT 10.6840 37.5435 10.7100 38.6370 ;
        RECT 10.5760 37.5435 10.6020 38.6370 ;
        RECT 10.4680 37.5435 10.4940 38.6370 ;
        RECT 10.3600 37.5435 10.3860 38.6370 ;
        RECT 10.2520 37.5435 10.2780 38.6370 ;
        RECT 10.1440 37.5435 10.1700 38.6370 ;
        RECT 10.0360 37.5435 10.0620 38.6370 ;
        RECT 9.9280 37.5435 9.9540 38.6370 ;
        RECT 9.8200 37.5435 9.8460 38.6370 ;
        RECT 9.7120 37.5435 9.7380 38.6370 ;
        RECT 9.6040 37.5435 9.6300 38.6370 ;
        RECT 9.4960 37.5435 9.5220 38.6370 ;
        RECT 9.3880 37.5435 9.4140 38.6370 ;
        RECT 9.1750 37.5435 9.2520 38.6370 ;
        RECT 7.2820 37.5435 7.3590 38.6370 ;
        RECT 7.1200 37.5435 7.1460 38.6370 ;
        RECT 7.0120 37.5435 7.0380 38.6370 ;
        RECT 6.9040 37.5435 6.9300 38.6370 ;
        RECT 6.7960 37.5435 6.8220 38.6370 ;
        RECT 6.6880 37.5435 6.7140 38.6370 ;
        RECT 6.5800 37.5435 6.6060 38.6370 ;
        RECT 6.4720 37.5435 6.4980 38.6370 ;
        RECT 6.3640 37.5435 6.3900 38.6370 ;
        RECT 6.2560 37.5435 6.2820 38.6370 ;
        RECT 6.1480 37.5435 6.1740 38.6370 ;
        RECT 6.0400 37.5435 6.0660 38.6370 ;
        RECT 5.9320 37.5435 5.9580 38.6370 ;
        RECT 5.8240 37.5435 5.8500 38.6370 ;
        RECT 5.7160 37.5435 5.7420 38.6370 ;
        RECT 5.6080 37.5435 5.6340 38.6370 ;
        RECT 5.5000 37.5435 5.5260 38.6370 ;
        RECT 5.3920 37.5435 5.4180 38.6370 ;
        RECT 5.2840 37.5435 5.3100 38.6370 ;
        RECT 5.1760 37.5435 5.2020 38.6370 ;
        RECT 5.0680 37.5435 5.0940 38.6370 ;
        RECT 4.9600 37.5435 4.9860 38.6370 ;
        RECT 4.8520 37.5435 4.8780 38.6370 ;
        RECT 4.7440 37.5435 4.7700 38.6370 ;
        RECT 4.6360 37.5435 4.6620 38.6370 ;
        RECT 4.5280 37.5435 4.5540 38.6370 ;
        RECT 4.4200 37.5435 4.4460 38.6370 ;
        RECT 4.3120 37.5435 4.3380 38.6370 ;
        RECT 4.2040 37.5435 4.2300 38.6370 ;
        RECT 4.0960 37.5435 4.1220 38.6370 ;
        RECT 3.9880 37.5435 4.0140 38.6370 ;
        RECT 3.8800 37.5435 3.9060 38.6370 ;
        RECT 3.7720 37.5435 3.7980 38.6370 ;
        RECT 3.6640 37.5435 3.6900 38.6370 ;
        RECT 3.5560 37.5435 3.5820 38.6370 ;
        RECT 3.4480 37.5435 3.4740 38.6370 ;
        RECT 3.3400 37.5435 3.3660 38.6370 ;
        RECT 3.2320 37.5435 3.2580 38.6370 ;
        RECT 3.1240 37.5435 3.1500 38.6370 ;
        RECT 3.0160 37.5435 3.0420 38.6370 ;
        RECT 2.9080 37.5435 2.9340 38.6370 ;
        RECT 2.8000 37.5435 2.8260 38.6370 ;
        RECT 2.6920 37.5435 2.7180 38.6370 ;
        RECT 2.5840 37.5435 2.6100 38.6370 ;
        RECT 2.4760 37.5435 2.5020 38.6370 ;
        RECT 2.3680 37.5435 2.3940 38.6370 ;
        RECT 2.2600 37.5435 2.2860 38.6370 ;
        RECT 2.1520 37.5435 2.1780 38.6370 ;
        RECT 2.0440 37.5435 2.0700 38.6370 ;
        RECT 1.9360 37.5435 1.9620 38.6370 ;
        RECT 1.8280 37.5435 1.8540 38.6370 ;
        RECT 1.7200 37.5435 1.7460 38.6370 ;
        RECT 1.6120 37.5435 1.6380 38.6370 ;
        RECT 1.5040 37.5435 1.5300 38.6370 ;
        RECT 1.3960 37.5435 1.4220 38.6370 ;
        RECT 1.2880 37.5435 1.3140 38.6370 ;
        RECT 1.1800 37.5435 1.2060 38.6370 ;
        RECT 1.0720 37.5435 1.0980 38.6370 ;
        RECT 0.9640 37.5435 0.9900 38.6370 ;
        RECT 0.8560 37.5435 0.8820 38.6370 ;
        RECT 0.7480 37.5435 0.7740 38.6370 ;
        RECT 0.6400 37.5435 0.6660 38.6370 ;
        RECT 0.5320 37.5435 0.5580 38.6370 ;
        RECT 0.4240 37.5435 0.4500 38.6370 ;
        RECT 0.3160 37.5435 0.3420 38.6370 ;
        RECT 0.2080 37.5435 0.2340 38.6370 ;
        RECT 0.0050 37.5435 0.0900 38.6370 ;
        RECT 8.6410 38.6235 8.7690 39.7170 ;
        RECT 8.6270 39.2890 8.7690 39.6115 ;
        RECT 8.4790 39.0160 8.5410 39.7170 ;
        RECT 8.4650 39.3255 8.5410 39.4790 ;
        RECT 8.4790 38.6235 8.5050 39.7170 ;
        RECT 8.4790 38.7445 8.5190 38.9840 ;
        RECT 8.4790 38.6235 8.5410 38.7125 ;
        RECT 8.1820 39.0740 8.3880 39.7170 ;
        RECT 8.3620 38.6235 8.3880 39.7170 ;
        RECT 8.1820 39.3510 8.4020 39.6090 ;
        RECT 8.1820 38.6235 8.2800 39.7170 ;
        RECT 7.7650 38.6235 7.8480 39.7170 ;
        RECT 7.7650 38.7120 7.8620 39.6475 ;
        RECT 16.4440 38.6235 16.5290 39.7170 ;
        RECT 16.3000 38.6235 16.3260 39.7170 ;
        RECT 16.1920 38.6235 16.2180 39.7170 ;
        RECT 16.0840 38.6235 16.1100 39.7170 ;
        RECT 15.9760 38.6235 16.0020 39.7170 ;
        RECT 15.8680 38.6235 15.8940 39.7170 ;
        RECT 15.7600 38.6235 15.7860 39.7170 ;
        RECT 15.6520 38.6235 15.6780 39.7170 ;
        RECT 15.5440 38.6235 15.5700 39.7170 ;
        RECT 15.4360 38.6235 15.4620 39.7170 ;
        RECT 15.3280 38.6235 15.3540 39.7170 ;
        RECT 15.2200 38.6235 15.2460 39.7170 ;
        RECT 15.1120 38.6235 15.1380 39.7170 ;
        RECT 15.0040 38.6235 15.0300 39.7170 ;
        RECT 14.8960 38.6235 14.9220 39.7170 ;
        RECT 14.7880 38.6235 14.8140 39.7170 ;
        RECT 14.6800 38.6235 14.7060 39.7170 ;
        RECT 14.5720 38.6235 14.5980 39.7170 ;
        RECT 14.4640 38.6235 14.4900 39.7170 ;
        RECT 14.3560 38.6235 14.3820 39.7170 ;
        RECT 14.2480 38.6235 14.2740 39.7170 ;
        RECT 14.1400 38.6235 14.1660 39.7170 ;
        RECT 14.0320 38.6235 14.0580 39.7170 ;
        RECT 13.9240 38.6235 13.9500 39.7170 ;
        RECT 13.8160 38.6235 13.8420 39.7170 ;
        RECT 13.7080 38.6235 13.7340 39.7170 ;
        RECT 13.6000 38.6235 13.6260 39.7170 ;
        RECT 13.4920 38.6235 13.5180 39.7170 ;
        RECT 13.3840 38.6235 13.4100 39.7170 ;
        RECT 13.2760 38.6235 13.3020 39.7170 ;
        RECT 13.1680 38.6235 13.1940 39.7170 ;
        RECT 13.0600 38.6235 13.0860 39.7170 ;
        RECT 12.9520 38.6235 12.9780 39.7170 ;
        RECT 12.8440 38.6235 12.8700 39.7170 ;
        RECT 12.7360 38.6235 12.7620 39.7170 ;
        RECT 12.6280 38.6235 12.6540 39.7170 ;
        RECT 12.5200 38.6235 12.5460 39.7170 ;
        RECT 12.4120 38.6235 12.4380 39.7170 ;
        RECT 12.3040 38.6235 12.3300 39.7170 ;
        RECT 12.1960 38.6235 12.2220 39.7170 ;
        RECT 12.0880 38.6235 12.1140 39.7170 ;
        RECT 11.9800 38.6235 12.0060 39.7170 ;
        RECT 11.8720 38.6235 11.8980 39.7170 ;
        RECT 11.7640 38.6235 11.7900 39.7170 ;
        RECT 11.6560 38.6235 11.6820 39.7170 ;
        RECT 11.5480 38.6235 11.5740 39.7170 ;
        RECT 11.4400 38.6235 11.4660 39.7170 ;
        RECT 11.3320 38.6235 11.3580 39.7170 ;
        RECT 11.2240 38.6235 11.2500 39.7170 ;
        RECT 11.1160 38.6235 11.1420 39.7170 ;
        RECT 11.0080 38.6235 11.0340 39.7170 ;
        RECT 10.9000 38.6235 10.9260 39.7170 ;
        RECT 10.7920 38.6235 10.8180 39.7170 ;
        RECT 10.6840 38.6235 10.7100 39.7170 ;
        RECT 10.5760 38.6235 10.6020 39.7170 ;
        RECT 10.4680 38.6235 10.4940 39.7170 ;
        RECT 10.3600 38.6235 10.3860 39.7170 ;
        RECT 10.2520 38.6235 10.2780 39.7170 ;
        RECT 10.1440 38.6235 10.1700 39.7170 ;
        RECT 10.0360 38.6235 10.0620 39.7170 ;
        RECT 9.9280 38.6235 9.9540 39.7170 ;
        RECT 9.8200 38.6235 9.8460 39.7170 ;
        RECT 9.7120 38.6235 9.7380 39.7170 ;
        RECT 9.6040 38.6235 9.6300 39.7170 ;
        RECT 9.4960 38.6235 9.5220 39.7170 ;
        RECT 9.3880 38.6235 9.4140 39.7170 ;
        RECT 9.1750 38.6235 9.2520 39.7170 ;
        RECT 7.2820 38.6235 7.3590 39.7170 ;
        RECT 7.1200 38.6235 7.1460 39.7170 ;
        RECT 7.0120 38.6235 7.0380 39.7170 ;
        RECT 6.9040 38.6235 6.9300 39.7170 ;
        RECT 6.7960 38.6235 6.8220 39.7170 ;
        RECT 6.6880 38.6235 6.7140 39.7170 ;
        RECT 6.5800 38.6235 6.6060 39.7170 ;
        RECT 6.4720 38.6235 6.4980 39.7170 ;
        RECT 6.3640 38.6235 6.3900 39.7170 ;
        RECT 6.2560 38.6235 6.2820 39.7170 ;
        RECT 6.1480 38.6235 6.1740 39.7170 ;
        RECT 6.0400 38.6235 6.0660 39.7170 ;
        RECT 5.9320 38.6235 5.9580 39.7170 ;
        RECT 5.8240 38.6235 5.8500 39.7170 ;
        RECT 5.7160 38.6235 5.7420 39.7170 ;
        RECT 5.6080 38.6235 5.6340 39.7170 ;
        RECT 5.5000 38.6235 5.5260 39.7170 ;
        RECT 5.3920 38.6235 5.4180 39.7170 ;
        RECT 5.2840 38.6235 5.3100 39.7170 ;
        RECT 5.1760 38.6235 5.2020 39.7170 ;
        RECT 5.0680 38.6235 5.0940 39.7170 ;
        RECT 4.9600 38.6235 4.9860 39.7170 ;
        RECT 4.8520 38.6235 4.8780 39.7170 ;
        RECT 4.7440 38.6235 4.7700 39.7170 ;
        RECT 4.6360 38.6235 4.6620 39.7170 ;
        RECT 4.5280 38.6235 4.5540 39.7170 ;
        RECT 4.4200 38.6235 4.4460 39.7170 ;
        RECT 4.3120 38.6235 4.3380 39.7170 ;
        RECT 4.2040 38.6235 4.2300 39.7170 ;
        RECT 4.0960 38.6235 4.1220 39.7170 ;
        RECT 3.9880 38.6235 4.0140 39.7170 ;
        RECT 3.8800 38.6235 3.9060 39.7170 ;
        RECT 3.7720 38.6235 3.7980 39.7170 ;
        RECT 3.6640 38.6235 3.6900 39.7170 ;
        RECT 3.5560 38.6235 3.5820 39.7170 ;
        RECT 3.4480 38.6235 3.4740 39.7170 ;
        RECT 3.3400 38.6235 3.3660 39.7170 ;
        RECT 3.2320 38.6235 3.2580 39.7170 ;
        RECT 3.1240 38.6235 3.1500 39.7170 ;
        RECT 3.0160 38.6235 3.0420 39.7170 ;
        RECT 2.9080 38.6235 2.9340 39.7170 ;
        RECT 2.8000 38.6235 2.8260 39.7170 ;
        RECT 2.6920 38.6235 2.7180 39.7170 ;
        RECT 2.5840 38.6235 2.6100 39.7170 ;
        RECT 2.4760 38.6235 2.5020 39.7170 ;
        RECT 2.3680 38.6235 2.3940 39.7170 ;
        RECT 2.2600 38.6235 2.2860 39.7170 ;
        RECT 2.1520 38.6235 2.1780 39.7170 ;
        RECT 2.0440 38.6235 2.0700 39.7170 ;
        RECT 1.9360 38.6235 1.9620 39.7170 ;
        RECT 1.8280 38.6235 1.8540 39.7170 ;
        RECT 1.7200 38.6235 1.7460 39.7170 ;
        RECT 1.6120 38.6235 1.6380 39.7170 ;
        RECT 1.5040 38.6235 1.5300 39.7170 ;
        RECT 1.3960 38.6235 1.4220 39.7170 ;
        RECT 1.2880 38.6235 1.3140 39.7170 ;
        RECT 1.1800 38.6235 1.2060 39.7170 ;
        RECT 1.0720 38.6235 1.0980 39.7170 ;
        RECT 0.9640 38.6235 0.9900 39.7170 ;
        RECT 0.8560 38.6235 0.8820 39.7170 ;
        RECT 0.7480 38.6235 0.7740 39.7170 ;
        RECT 0.6400 38.6235 0.6660 39.7170 ;
        RECT 0.5320 38.6235 0.5580 39.7170 ;
        RECT 0.4240 38.6235 0.4500 39.7170 ;
        RECT 0.3160 38.6235 0.3420 39.7170 ;
        RECT 0.2080 38.6235 0.2340 39.7170 ;
        RECT 0.0050 38.6235 0.0900 39.7170 ;
        RECT 8.6410 39.7035 8.7690 40.7970 ;
        RECT 8.6270 40.3690 8.7690 40.6915 ;
        RECT 8.4790 40.0960 8.5410 40.7970 ;
        RECT 8.4650 40.4055 8.5410 40.5590 ;
        RECT 8.4790 39.7035 8.5050 40.7970 ;
        RECT 8.4790 39.8245 8.5190 40.0640 ;
        RECT 8.4790 39.7035 8.5410 39.7925 ;
        RECT 8.1820 40.1540 8.3880 40.7970 ;
        RECT 8.3620 39.7035 8.3880 40.7970 ;
        RECT 8.1820 40.4310 8.4020 40.6890 ;
        RECT 8.1820 39.7035 8.2800 40.7970 ;
        RECT 7.7650 39.7035 7.8480 40.7970 ;
        RECT 7.7650 39.7920 7.8620 40.7275 ;
        RECT 16.4440 39.7035 16.5290 40.7970 ;
        RECT 16.3000 39.7035 16.3260 40.7970 ;
        RECT 16.1920 39.7035 16.2180 40.7970 ;
        RECT 16.0840 39.7035 16.1100 40.7970 ;
        RECT 15.9760 39.7035 16.0020 40.7970 ;
        RECT 15.8680 39.7035 15.8940 40.7970 ;
        RECT 15.7600 39.7035 15.7860 40.7970 ;
        RECT 15.6520 39.7035 15.6780 40.7970 ;
        RECT 15.5440 39.7035 15.5700 40.7970 ;
        RECT 15.4360 39.7035 15.4620 40.7970 ;
        RECT 15.3280 39.7035 15.3540 40.7970 ;
        RECT 15.2200 39.7035 15.2460 40.7970 ;
        RECT 15.1120 39.7035 15.1380 40.7970 ;
        RECT 15.0040 39.7035 15.0300 40.7970 ;
        RECT 14.8960 39.7035 14.9220 40.7970 ;
        RECT 14.7880 39.7035 14.8140 40.7970 ;
        RECT 14.6800 39.7035 14.7060 40.7970 ;
        RECT 14.5720 39.7035 14.5980 40.7970 ;
        RECT 14.4640 39.7035 14.4900 40.7970 ;
        RECT 14.3560 39.7035 14.3820 40.7970 ;
        RECT 14.2480 39.7035 14.2740 40.7970 ;
        RECT 14.1400 39.7035 14.1660 40.7970 ;
        RECT 14.0320 39.7035 14.0580 40.7970 ;
        RECT 13.9240 39.7035 13.9500 40.7970 ;
        RECT 13.8160 39.7035 13.8420 40.7970 ;
        RECT 13.7080 39.7035 13.7340 40.7970 ;
        RECT 13.6000 39.7035 13.6260 40.7970 ;
        RECT 13.4920 39.7035 13.5180 40.7970 ;
        RECT 13.3840 39.7035 13.4100 40.7970 ;
        RECT 13.2760 39.7035 13.3020 40.7970 ;
        RECT 13.1680 39.7035 13.1940 40.7970 ;
        RECT 13.0600 39.7035 13.0860 40.7970 ;
        RECT 12.9520 39.7035 12.9780 40.7970 ;
        RECT 12.8440 39.7035 12.8700 40.7970 ;
        RECT 12.7360 39.7035 12.7620 40.7970 ;
        RECT 12.6280 39.7035 12.6540 40.7970 ;
        RECT 12.5200 39.7035 12.5460 40.7970 ;
        RECT 12.4120 39.7035 12.4380 40.7970 ;
        RECT 12.3040 39.7035 12.3300 40.7970 ;
        RECT 12.1960 39.7035 12.2220 40.7970 ;
        RECT 12.0880 39.7035 12.1140 40.7970 ;
        RECT 11.9800 39.7035 12.0060 40.7970 ;
        RECT 11.8720 39.7035 11.8980 40.7970 ;
        RECT 11.7640 39.7035 11.7900 40.7970 ;
        RECT 11.6560 39.7035 11.6820 40.7970 ;
        RECT 11.5480 39.7035 11.5740 40.7970 ;
        RECT 11.4400 39.7035 11.4660 40.7970 ;
        RECT 11.3320 39.7035 11.3580 40.7970 ;
        RECT 11.2240 39.7035 11.2500 40.7970 ;
        RECT 11.1160 39.7035 11.1420 40.7970 ;
        RECT 11.0080 39.7035 11.0340 40.7970 ;
        RECT 10.9000 39.7035 10.9260 40.7970 ;
        RECT 10.7920 39.7035 10.8180 40.7970 ;
        RECT 10.6840 39.7035 10.7100 40.7970 ;
        RECT 10.5760 39.7035 10.6020 40.7970 ;
        RECT 10.4680 39.7035 10.4940 40.7970 ;
        RECT 10.3600 39.7035 10.3860 40.7970 ;
        RECT 10.2520 39.7035 10.2780 40.7970 ;
        RECT 10.1440 39.7035 10.1700 40.7970 ;
        RECT 10.0360 39.7035 10.0620 40.7970 ;
        RECT 9.9280 39.7035 9.9540 40.7970 ;
        RECT 9.8200 39.7035 9.8460 40.7970 ;
        RECT 9.7120 39.7035 9.7380 40.7970 ;
        RECT 9.6040 39.7035 9.6300 40.7970 ;
        RECT 9.4960 39.7035 9.5220 40.7970 ;
        RECT 9.3880 39.7035 9.4140 40.7970 ;
        RECT 9.1750 39.7035 9.2520 40.7970 ;
        RECT 7.2820 39.7035 7.3590 40.7970 ;
        RECT 7.1200 39.7035 7.1460 40.7970 ;
        RECT 7.0120 39.7035 7.0380 40.7970 ;
        RECT 6.9040 39.7035 6.9300 40.7970 ;
        RECT 6.7960 39.7035 6.8220 40.7970 ;
        RECT 6.6880 39.7035 6.7140 40.7970 ;
        RECT 6.5800 39.7035 6.6060 40.7970 ;
        RECT 6.4720 39.7035 6.4980 40.7970 ;
        RECT 6.3640 39.7035 6.3900 40.7970 ;
        RECT 6.2560 39.7035 6.2820 40.7970 ;
        RECT 6.1480 39.7035 6.1740 40.7970 ;
        RECT 6.0400 39.7035 6.0660 40.7970 ;
        RECT 5.9320 39.7035 5.9580 40.7970 ;
        RECT 5.8240 39.7035 5.8500 40.7970 ;
        RECT 5.7160 39.7035 5.7420 40.7970 ;
        RECT 5.6080 39.7035 5.6340 40.7970 ;
        RECT 5.5000 39.7035 5.5260 40.7970 ;
        RECT 5.3920 39.7035 5.4180 40.7970 ;
        RECT 5.2840 39.7035 5.3100 40.7970 ;
        RECT 5.1760 39.7035 5.2020 40.7970 ;
        RECT 5.0680 39.7035 5.0940 40.7970 ;
        RECT 4.9600 39.7035 4.9860 40.7970 ;
        RECT 4.8520 39.7035 4.8780 40.7970 ;
        RECT 4.7440 39.7035 4.7700 40.7970 ;
        RECT 4.6360 39.7035 4.6620 40.7970 ;
        RECT 4.5280 39.7035 4.5540 40.7970 ;
        RECT 4.4200 39.7035 4.4460 40.7970 ;
        RECT 4.3120 39.7035 4.3380 40.7970 ;
        RECT 4.2040 39.7035 4.2300 40.7970 ;
        RECT 4.0960 39.7035 4.1220 40.7970 ;
        RECT 3.9880 39.7035 4.0140 40.7970 ;
        RECT 3.8800 39.7035 3.9060 40.7970 ;
        RECT 3.7720 39.7035 3.7980 40.7970 ;
        RECT 3.6640 39.7035 3.6900 40.7970 ;
        RECT 3.5560 39.7035 3.5820 40.7970 ;
        RECT 3.4480 39.7035 3.4740 40.7970 ;
        RECT 3.3400 39.7035 3.3660 40.7970 ;
        RECT 3.2320 39.7035 3.2580 40.7970 ;
        RECT 3.1240 39.7035 3.1500 40.7970 ;
        RECT 3.0160 39.7035 3.0420 40.7970 ;
        RECT 2.9080 39.7035 2.9340 40.7970 ;
        RECT 2.8000 39.7035 2.8260 40.7970 ;
        RECT 2.6920 39.7035 2.7180 40.7970 ;
        RECT 2.5840 39.7035 2.6100 40.7970 ;
        RECT 2.4760 39.7035 2.5020 40.7970 ;
        RECT 2.3680 39.7035 2.3940 40.7970 ;
        RECT 2.2600 39.7035 2.2860 40.7970 ;
        RECT 2.1520 39.7035 2.1780 40.7970 ;
        RECT 2.0440 39.7035 2.0700 40.7970 ;
        RECT 1.9360 39.7035 1.9620 40.7970 ;
        RECT 1.8280 39.7035 1.8540 40.7970 ;
        RECT 1.7200 39.7035 1.7460 40.7970 ;
        RECT 1.6120 39.7035 1.6380 40.7970 ;
        RECT 1.5040 39.7035 1.5300 40.7970 ;
        RECT 1.3960 39.7035 1.4220 40.7970 ;
        RECT 1.2880 39.7035 1.3140 40.7970 ;
        RECT 1.1800 39.7035 1.2060 40.7970 ;
        RECT 1.0720 39.7035 1.0980 40.7970 ;
        RECT 0.9640 39.7035 0.9900 40.7970 ;
        RECT 0.8560 39.7035 0.8820 40.7970 ;
        RECT 0.7480 39.7035 0.7740 40.7970 ;
        RECT 0.6400 39.7035 0.6660 40.7970 ;
        RECT 0.5320 39.7035 0.5580 40.7970 ;
        RECT 0.4240 39.7035 0.4500 40.7970 ;
        RECT 0.3160 39.7035 0.3420 40.7970 ;
        RECT 0.2080 39.7035 0.2340 40.7970 ;
        RECT 0.0050 39.7035 0.0900 40.7970 ;
        RECT 8.6410 40.7835 8.7690 41.8770 ;
        RECT 8.6270 41.4490 8.7690 41.7715 ;
        RECT 8.4790 41.1760 8.5410 41.8770 ;
        RECT 8.4650 41.4855 8.5410 41.6390 ;
        RECT 8.4790 40.7835 8.5050 41.8770 ;
        RECT 8.4790 40.9045 8.5190 41.1440 ;
        RECT 8.4790 40.7835 8.5410 40.8725 ;
        RECT 8.1820 41.2340 8.3880 41.8770 ;
        RECT 8.3620 40.7835 8.3880 41.8770 ;
        RECT 8.1820 41.5110 8.4020 41.7690 ;
        RECT 8.1820 40.7835 8.2800 41.8770 ;
        RECT 7.7650 40.7835 7.8480 41.8770 ;
        RECT 7.7650 40.8720 7.8620 41.8075 ;
        RECT 16.4440 40.7835 16.5290 41.8770 ;
        RECT 16.3000 40.7835 16.3260 41.8770 ;
        RECT 16.1920 40.7835 16.2180 41.8770 ;
        RECT 16.0840 40.7835 16.1100 41.8770 ;
        RECT 15.9760 40.7835 16.0020 41.8770 ;
        RECT 15.8680 40.7835 15.8940 41.8770 ;
        RECT 15.7600 40.7835 15.7860 41.8770 ;
        RECT 15.6520 40.7835 15.6780 41.8770 ;
        RECT 15.5440 40.7835 15.5700 41.8770 ;
        RECT 15.4360 40.7835 15.4620 41.8770 ;
        RECT 15.3280 40.7835 15.3540 41.8770 ;
        RECT 15.2200 40.7835 15.2460 41.8770 ;
        RECT 15.1120 40.7835 15.1380 41.8770 ;
        RECT 15.0040 40.7835 15.0300 41.8770 ;
        RECT 14.8960 40.7835 14.9220 41.8770 ;
        RECT 14.7880 40.7835 14.8140 41.8770 ;
        RECT 14.6800 40.7835 14.7060 41.8770 ;
        RECT 14.5720 40.7835 14.5980 41.8770 ;
        RECT 14.4640 40.7835 14.4900 41.8770 ;
        RECT 14.3560 40.7835 14.3820 41.8770 ;
        RECT 14.2480 40.7835 14.2740 41.8770 ;
        RECT 14.1400 40.7835 14.1660 41.8770 ;
        RECT 14.0320 40.7835 14.0580 41.8770 ;
        RECT 13.9240 40.7835 13.9500 41.8770 ;
        RECT 13.8160 40.7835 13.8420 41.8770 ;
        RECT 13.7080 40.7835 13.7340 41.8770 ;
        RECT 13.6000 40.7835 13.6260 41.8770 ;
        RECT 13.4920 40.7835 13.5180 41.8770 ;
        RECT 13.3840 40.7835 13.4100 41.8770 ;
        RECT 13.2760 40.7835 13.3020 41.8770 ;
        RECT 13.1680 40.7835 13.1940 41.8770 ;
        RECT 13.0600 40.7835 13.0860 41.8770 ;
        RECT 12.9520 40.7835 12.9780 41.8770 ;
        RECT 12.8440 40.7835 12.8700 41.8770 ;
        RECT 12.7360 40.7835 12.7620 41.8770 ;
        RECT 12.6280 40.7835 12.6540 41.8770 ;
        RECT 12.5200 40.7835 12.5460 41.8770 ;
        RECT 12.4120 40.7835 12.4380 41.8770 ;
        RECT 12.3040 40.7835 12.3300 41.8770 ;
        RECT 12.1960 40.7835 12.2220 41.8770 ;
        RECT 12.0880 40.7835 12.1140 41.8770 ;
        RECT 11.9800 40.7835 12.0060 41.8770 ;
        RECT 11.8720 40.7835 11.8980 41.8770 ;
        RECT 11.7640 40.7835 11.7900 41.8770 ;
        RECT 11.6560 40.7835 11.6820 41.8770 ;
        RECT 11.5480 40.7835 11.5740 41.8770 ;
        RECT 11.4400 40.7835 11.4660 41.8770 ;
        RECT 11.3320 40.7835 11.3580 41.8770 ;
        RECT 11.2240 40.7835 11.2500 41.8770 ;
        RECT 11.1160 40.7835 11.1420 41.8770 ;
        RECT 11.0080 40.7835 11.0340 41.8770 ;
        RECT 10.9000 40.7835 10.9260 41.8770 ;
        RECT 10.7920 40.7835 10.8180 41.8770 ;
        RECT 10.6840 40.7835 10.7100 41.8770 ;
        RECT 10.5760 40.7835 10.6020 41.8770 ;
        RECT 10.4680 40.7835 10.4940 41.8770 ;
        RECT 10.3600 40.7835 10.3860 41.8770 ;
        RECT 10.2520 40.7835 10.2780 41.8770 ;
        RECT 10.1440 40.7835 10.1700 41.8770 ;
        RECT 10.0360 40.7835 10.0620 41.8770 ;
        RECT 9.9280 40.7835 9.9540 41.8770 ;
        RECT 9.8200 40.7835 9.8460 41.8770 ;
        RECT 9.7120 40.7835 9.7380 41.8770 ;
        RECT 9.6040 40.7835 9.6300 41.8770 ;
        RECT 9.4960 40.7835 9.5220 41.8770 ;
        RECT 9.3880 40.7835 9.4140 41.8770 ;
        RECT 9.1750 40.7835 9.2520 41.8770 ;
        RECT 7.2820 40.7835 7.3590 41.8770 ;
        RECT 7.1200 40.7835 7.1460 41.8770 ;
        RECT 7.0120 40.7835 7.0380 41.8770 ;
        RECT 6.9040 40.7835 6.9300 41.8770 ;
        RECT 6.7960 40.7835 6.8220 41.8770 ;
        RECT 6.6880 40.7835 6.7140 41.8770 ;
        RECT 6.5800 40.7835 6.6060 41.8770 ;
        RECT 6.4720 40.7835 6.4980 41.8770 ;
        RECT 6.3640 40.7835 6.3900 41.8770 ;
        RECT 6.2560 40.7835 6.2820 41.8770 ;
        RECT 6.1480 40.7835 6.1740 41.8770 ;
        RECT 6.0400 40.7835 6.0660 41.8770 ;
        RECT 5.9320 40.7835 5.9580 41.8770 ;
        RECT 5.8240 40.7835 5.8500 41.8770 ;
        RECT 5.7160 40.7835 5.7420 41.8770 ;
        RECT 5.6080 40.7835 5.6340 41.8770 ;
        RECT 5.5000 40.7835 5.5260 41.8770 ;
        RECT 5.3920 40.7835 5.4180 41.8770 ;
        RECT 5.2840 40.7835 5.3100 41.8770 ;
        RECT 5.1760 40.7835 5.2020 41.8770 ;
        RECT 5.0680 40.7835 5.0940 41.8770 ;
        RECT 4.9600 40.7835 4.9860 41.8770 ;
        RECT 4.8520 40.7835 4.8780 41.8770 ;
        RECT 4.7440 40.7835 4.7700 41.8770 ;
        RECT 4.6360 40.7835 4.6620 41.8770 ;
        RECT 4.5280 40.7835 4.5540 41.8770 ;
        RECT 4.4200 40.7835 4.4460 41.8770 ;
        RECT 4.3120 40.7835 4.3380 41.8770 ;
        RECT 4.2040 40.7835 4.2300 41.8770 ;
        RECT 4.0960 40.7835 4.1220 41.8770 ;
        RECT 3.9880 40.7835 4.0140 41.8770 ;
        RECT 3.8800 40.7835 3.9060 41.8770 ;
        RECT 3.7720 40.7835 3.7980 41.8770 ;
        RECT 3.6640 40.7835 3.6900 41.8770 ;
        RECT 3.5560 40.7835 3.5820 41.8770 ;
        RECT 3.4480 40.7835 3.4740 41.8770 ;
        RECT 3.3400 40.7835 3.3660 41.8770 ;
        RECT 3.2320 40.7835 3.2580 41.8770 ;
        RECT 3.1240 40.7835 3.1500 41.8770 ;
        RECT 3.0160 40.7835 3.0420 41.8770 ;
        RECT 2.9080 40.7835 2.9340 41.8770 ;
        RECT 2.8000 40.7835 2.8260 41.8770 ;
        RECT 2.6920 40.7835 2.7180 41.8770 ;
        RECT 2.5840 40.7835 2.6100 41.8770 ;
        RECT 2.4760 40.7835 2.5020 41.8770 ;
        RECT 2.3680 40.7835 2.3940 41.8770 ;
        RECT 2.2600 40.7835 2.2860 41.8770 ;
        RECT 2.1520 40.7835 2.1780 41.8770 ;
        RECT 2.0440 40.7835 2.0700 41.8770 ;
        RECT 1.9360 40.7835 1.9620 41.8770 ;
        RECT 1.8280 40.7835 1.8540 41.8770 ;
        RECT 1.7200 40.7835 1.7460 41.8770 ;
        RECT 1.6120 40.7835 1.6380 41.8770 ;
        RECT 1.5040 40.7835 1.5300 41.8770 ;
        RECT 1.3960 40.7835 1.4220 41.8770 ;
        RECT 1.2880 40.7835 1.3140 41.8770 ;
        RECT 1.1800 40.7835 1.2060 41.8770 ;
        RECT 1.0720 40.7835 1.0980 41.8770 ;
        RECT 0.9640 40.7835 0.9900 41.8770 ;
        RECT 0.8560 40.7835 0.8820 41.8770 ;
        RECT 0.7480 40.7835 0.7740 41.8770 ;
        RECT 0.6400 40.7835 0.6660 41.8770 ;
        RECT 0.5320 40.7835 0.5580 41.8770 ;
        RECT 0.4240 40.7835 0.4500 41.8770 ;
        RECT 0.3160 40.7835 0.3420 41.8770 ;
        RECT 0.2080 40.7835 0.2340 41.8770 ;
        RECT 0.0050 40.7835 0.0900 41.8770 ;
        RECT 8.6410 41.8635 8.7690 42.9570 ;
        RECT 8.6270 42.5290 8.7690 42.8515 ;
        RECT 8.4790 42.2560 8.5410 42.9570 ;
        RECT 8.4650 42.5655 8.5410 42.7190 ;
        RECT 8.4790 41.8635 8.5050 42.9570 ;
        RECT 8.4790 41.9845 8.5190 42.2240 ;
        RECT 8.4790 41.8635 8.5410 41.9525 ;
        RECT 8.1820 42.3140 8.3880 42.9570 ;
        RECT 8.3620 41.8635 8.3880 42.9570 ;
        RECT 8.1820 42.5910 8.4020 42.8490 ;
        RECT 8.1820 41.8635 8.2800 42.9570 ;
        RECT 7.7650 41.8635 7.8480 42.9570 ;
        RECT 7.7650 41.9520 7.8620 42.8875 ;
        RECT 16.4440 41.8635 16.5290 42.9570 ;
        RECT 16.3000 41.8635 16.3260 42.9570 ;
        RECT 16.1920 41.8635 16.2180 42.9570 ;
        RECT 16.0840 41.8635 16.1100 42.9570 ;
        RECT 15.9760 41.8635 16.0020 42.9570 ;
        RECT 15.8680 41.8635 15.8940 42.9570 ;
        RECT 15.7600 41.8635 15.7860 42.9570 ;
        RECT 15.6520 41.8635 15.6780 42.9570 ;
        RECT 15.5440 41.8635 15.5700 42.9570 ;
        RECT 15.4360 41.8635 15.4620 42.9570 ;
        RECT 15.3280 41.8635 15.3540 42.9570 ;
        RECT 15.2200 41.8635 15.2460 42.9570 ;
        RECT 15.1120 41.8635 15.1380 42.9570 ;
        RECT 15.0040 41.8635 15.0300 42.9570 ;
        RECT 14.8960 41.8635 14.9220 42.9570 ;
        RECT 14.7880 41.8635 14.8140 42.9570 ;
        RECT 14.6800 41.8635 14.7060 42.9570 ;
        RECT 14.5720 41.8635 14.5980 42.9570 ;
        RECT 14.4640 41.8635 14.4900 42.9570 ;
        RECT 14.3560 41.8635 14.3820 42.9570 ;
        RECT 14.2480 41.8635 14.2740 42.9570 ;
        RECT 14.1400 41.8635 14.1660 42.9570 ;
        RECT 14.0320 41.8635 14.0580 42.9570 ;
        RECT 13.9240 41.8635 13.9500 42.9570 ;
        RECT 13.8160 41.8635 13.8420 42.9570 ;
        RECT 13.7080 41.8635 13.7340 42.9570 ;
        RECT 13.6000 41.8635 13.6260 42.9570 ;
        RECT 13.4920 41.8635 13.5180 42.9570 ;
        RECT 13.3840 41.8635 13.4100 42.9570 ;
        RECT 13.2760 41.8635 13.3020 42.9570 ;
        RECT 13.1680 41.8635 13.1940 42.9570 ;
        RECT 13.0600 41.8635 13.0860 42.9570 ;
        RECT 12.9520 41.8635 12.9780 42.9570 ;
        RECT 12.8440 41.8635 12.8700 42.9570 ;
        RECT 12.7360 41.8635 12.7620 42.9570 ;
        RECT 12.6280 41.8635 12.6540 42.9570 ;
        RECT 12.5200 41.8635 12.5460 42.9570 ;
        RECT 12.4120 41.8635 12.4380 42.9570 ;
        RECT 12.3040 41.8635 12.3300 42.9570 ;
        RECT 12.1960 41.8635 12.2220 42.9570 ;
        RECT 12.0880 41.8635 12.1140 42.9570 ;
        RECT 11.9800 41.8635 12.0060 42.9570 ;
        RECT 11.8720 41.8635 11.8980 42.9570 ;
        RECT 11.7640 41.8635 11.7900 42.9570 ;
        RECT 11.6560 41.8635 11.6820 42.9570 ;
        RECT 11.5480 41.8635 11.5740 42.9570 ;
        RECT 11.4400 41.8635 11.4660 42.9570 ;
        RECT 11.3320 41.8635 11.3580 42.9570 ;
        RECT 11.2240 41.8635 11.2500 42.9570 ;
        RECT 11.1160 41.8635 11.1420 42.9570 ;
        RECT 11.0080 41.8635 11.0340 42.9570 ;
        RECT 10.9000 41.8635 10.9260 42.9570 ;
        RECT 10.7920 41.8635 10.8180 42.9570 ;
        RECT 10.6840 41.8635 10.7100 42.9570 ;
        RECT 10.5760 41.8635 10.6020 42.9570 ;
        RECT 10.4680 41.8635 10.4940 42.9570 ;
        RECT 10.3600 41.8635 10.3860 42.9570 ;
        RECT 10.2520 41.8635 10.2780 42.9570 ;
        RECT 10.1440 41.8635 10.1700 42.9570 ;
        RECT 10.0360 41.8635 10.0620 42.9570 ;
        RECT 9.9280 41.8635 9.9540 42.9570 ;
        RECT 9.8200 41.8635 9.8460 42.9570 ;
        RECT 9.7120 41.8635 9.7380 42.9570 ;
        RECT 9.6040 41.8635 9.6300 42.9570 ;
        RECT 9.4960 41.8635 9.5220 42.9570 ;
        RECT 9.3880 41.8635 9.4140 42.9570 ;
        RECT 9.1750 41.8635 9.2520 42.9570 ;
        RECT 7.2820 41.8635 7.3590 42.9570 ;
        RECT 7.1200 41.8635 7.1460 42.9570 ;
        RECT 7.0120 41.8635 7.0380 42.9570 ;
        RECT 6.9040 41.8635 6.9300 42.9570 ;
        RECT 6.7960 41.8635 6.8220 42.9570 ;
        RECT 6.6880 41.8635 6.7140 42.9570 ;
        RECT 6.5800 41.8635 6.6060 42.9570 ;
        RECT 6.4720 41.8635 6.4980 42.9570 ;
        RECT 6.3640 41.8635 6.3900 42.9570 ;
        RECT 6.2560 41.8635 6.2820 42.9570 ;
        RECT 6.1480 41.8635 6.1740 42.9570 ;
        RECT 6.0400 41.8635 6.0660 42.9570 ;
        RECT 5.9320 41.8635 5.9580 42.9570 ;
        RECT 5.8240 41.8635 5.8500 42.9570 ;
        RECT 5.7160 41.8635 5.7420 42.9570 ;
        RECT 5.6080 41.8635 5.6340 42.9570 ;
        RECT 5.5000 41.8635 5.5260 42.9570 ;
        RECT 5.3920 41.8635 5.4180 42.9570 ;
        RECT 5.2840 41.8635 5.3100 42.9570 ;
        RECT 5.1760 41.8635 5.2020 42.9570 ;
        RECT 5.0680 41.8635 5.0940 42.9570 ;
        RECT 4.9600 41.8635 4.9860 42.9570 ;
        RECT 4.8520 41.8635 4.8780 42.9570 ;
        RECT 4.7440 41.8635 4.7700 42.9570 ;
        RECT 4.6360 41.8635 4.6620 42.9570 ;
        RECT 4.5280 41.8635 4.5540 42.9570 ;
        RECT 4.4200 41.8635 4.4460 42.9570 ;
        RECT 4.3120 41.8635 4.3380 42.9570 ;
        RECT 4.2040 41.8635 4.2300 42.9570 ;
        RECT 4.0960 41.8635 4.1220 42.9570 ;
        RECT 3.9880 41.8635 4.0140 42.9570 ;
        RECT 3.8800 41.8635 3.9060 42.9570 ;
        RECT 3.7720 41.8635 3.7980 42.9570 ;
        RECT 3.6640 41.8635 3.6900 42.9570 ;
        RECT 3.5560 41.8635 3.5820 42.9570 ;
        RECT 3.4480 41.8635 3.4740 42.9570 ;
        RECT 3.3400 41.8635 3.3660 42.9570 ;
        RECT 3.2320 41.8635 3.2580 42.9570 ;
        RECT 3.1240 41.8635 3.1500 42.9570 ;
        RECT 3.0160 41.8635 3.0420 42.9570 ;
        RECT 2.9080 41.8635 2.9340 42.9570 ;
        RECT 2.8000 41.8635 2.8260 42.9570 ;
        RECT 2.6920 41.8635 2.7180 42.9570 ;
        RECT 2.5840 41.8635 2.6100 42.9570 ;
        RECT 2.4760 41.8635 2.5020 42.9570 ;
        RECT 2.3680 41.8635 2.3940 42.9570 ;
        RECT 2.2600 41.8635 2.2860 42.9570 ;
        RECT 2.1520 41.8635 2.1780 42.9570 ;
        RECT 2.0440 41.8635 2.0700 42.9570 ;
        RECT 1.9360 41.8635 1.9620 42.9570 ;
        RECT 1.8280 41.8635 1.8540 42.9570 ;
        RECT 1.7200 41.8635 1.7460 42.9570 ;
        RECT 1.6120 41.8635 1.6380 42.9570 ;
        RECT 1.5040 41.8635 1.5300 42.9570 ;
        RECT 1.3960 41.8635 1.4220 42.9570 ;
        RECT 1.2880 41.8635 1.3140 42.9570 ;
        RECT 1.1800 41.8635 1.2060 42.9570 ;
        RECT 1.0720 41.8635 1.0980 42.9570 ;
        RECT 0.9640 41.8635 0.9900 42.9570 ;
        RECT 0.8560 41.8635 0.8820 42.9570 ;
        RECT 0.7480 41.8635 0.7740 42.9570 ;
        RECT 0.6400 41.8635 0.6660 42.9570 ;
        RECT 0.5320 41.8635 0.5580 42.9570 ;
        RECT 0.4240 41.8635 0.4500 42.9570 ;
        RECT 0.3160 41.8635 0.3420 42.9570 ;
        RECT 0.2080 41.8635 0.2340 42.9570 ;
        RECT 0.0050 41.8635 0.0900 42.9570 ;
        RECT 8.6410 42.9435 8.7690 44.0370 ;
        RECT 8.6270 43.6090 8.7690 43.9315 ;
        RECT 8.4790 43.3360 8.5410 44.0370 ;
        RECT 8.4650 43.6455 8.5410 43.7990 ;
        RECT 8.4790 42.9435 8.5050 44.0370 ;
        RECT 8.4790 43.0645 8.5190 43.3040 ;
        RECT 8.4790 42.9435 8.5410 43.0325 ;
        RECT 8.1820 43.3940 8.3880 44.0370 ;
        RECT 8.3620 42.9435 8.3880 44.0370 ;
        RECT 8.1820 43.6710 8.4020 43.9290 ;
        RECT 8.1820 42.9435 8.2800 44.0370 ;
        RECT 7.7650 42.9435 7.8480 44.0370 ;
        RECT 7.7650 43.0320 7.8620 43.9675 ;
        RECT 16.4440 42.9435 16.5290 44.0370 ;
        RECT 16.3000 42.9435 16.3260 44.0370 ;
        RECT 16.1920 42.9435 16.2180 44.0370 ;
        RECT 16.0840 42.9435 16.1100 44.0370 ;
        RECT 15.9760 42.9435 16.0020 44.0370 ;
        RECT 15.8680 42.9435 15.8940 44.0370 ;
        RECT 15.7600 42.9435 15.7860 44.0370 ;
        RECT 15.6520 42.9435 15.6780 44.0370 ;
        RECT 15.5440 42.9435 15.5700 44.0370 ;
        RECT 15.4360 42.9435 15.4620 44.0370 ;
        RECT 15.3280 42.9435 15.3540 44.0370 ;
        RECT 15.2200 42.9435 15.2460 44.0370 ;
        RECT 15.1120 42.9435 15.1380 44.0370 ;
        RECT 15.0040 42.9435 15.0300 44.0370 ;
        RECT 14.8960 42.9435 14.9220 44.0370 ;
        RECT 14.7880 42.9435 14.8140 44.0370 ;
        RECT 14.6800 42.9435 14.7060 44.0370 ;
        RECT 14.5720 42.9435 14.5980 44.0370 ;
        RECT 14.4640 42.9435 14.4900 44.0370 ;
        RECT 14.3560 42.9435 14.3820 44.0370 ;
        RECT 14.2480 42.9435 14.2740 44.0370 ;
        RECT 14.1400 42.9435 14.1660 44.0370 ;
        RECT 14.0320 42.9435 14.0580 44.0370 ;
        RECT 13.9240 42.9435 13.9500 44.0370 ;
        RECT 13.8160 42.9435 13.8420 44.0370 ;
        RECT 13.7080 42.9435 13.7340 44.0370 ;
        RECT 13.6000 42.9435 13.6260 44.0370 ;
        RECT 13.4920 42.9435 13.5180 44.0370 ;
        RECT 13.3840 42.9435 13.4100 44.0370 ;
        RECT 13.2760 42.9435 13.3020 44.0370 ;
        RECT 13.1680 42.9435 13.1940 44.0370 ;
        RECT 13.0600 42.9435 13.0860 44.0370 ;
        RECT 12.9520 42.9435 12.9780 44.0370 ;
        RECT 12.8440 42.9435 12.8700 44.0370 ;
        RECT 12.7360 42.9435 12.7620 44.0370 ;
        RECT 12.6280 42.9435 12.6540 44.0370 ;
        RECT 12.5200 42.9435 12.5460 44.0370 ;
        RECT 12.4120 42.9435 12.4380 44.0370 ;
        RECT 12.3040 42.9435 12.3300 44.0370 ;
        RECT 12.1960 42.9435 12.2220 44.0370 ;
        RECT 12.0880 42.9435 12.1140 44.0370 ;
        RECT 11.9800 42.9435 12.0060 44.0370 ;
        RECT 11.8720 42.9435 11.8980 44.0370 ;
        RECT 11.7640 42.9435 11.7900 44.0370 ;
        RECT 11.6560 42.9435 11.6820 44.0370 ;
        RECT 11.5480 42.9435 11.5740 44.0370 ;
        RECT 11.4400 42.9435 11.4660 44.0370 ;
        RECT 11.3320 42.9435 11.3580 44.0370 ;
        RECT 11.2240 42.9435 11.2500 44.0370 ;
        RECT 11.1160 42.9435 11.1420 44.0370 ;
        RECT 11.0080 42.9435 11.0340 44.0370 ;
        RECT 10.9000 42.9435 10.9260 44.0370 ;
        RECT 10.7920 42.9435 10.8180 44.0370 ;
        RECT 10.6840 42.9435 10.7100 44.0370 ;
        RECT 10.5760 42.9435 10.6020 44.0370 ;
        RECT 10.4680 42.9435 10.4940 44.0370 ;
        RECT 10.3600 42.9435 10.3860 44.0370 ;
        RECT 10.2520 42.9435 10.2780 44.0370 ;
        RECT 10.1440 42.9435 10.1700 44.0370 ;
        RECT 10.0360 42.9435 10.0620 44.0370 ;
        RECT 9.9280 42.9435 9.9540 44.0370 ;
        RECT 9.8200 42.9435 9.8460 44.0370 ;
        RECT 9.7120 42.9435 9.7380 44.0370 ;
        RECT 9.6040 42.9435 9.6300 44.0370 ;
        RECT 9.4960 42.9435 9.5220 44.0370 ;
        RECT 9.3880 42.9435 9.4140 44.0370 ;
        RECT 9.1750 42.9435 9.2520 44.0370 ;
        RECT 7.2820 42.9435 7.3590 44.0370 ;
        RECT 7.1200 42.9435 7.1460 44.0370 ;
        RECT 7.0120 42.9435 7.0380 44.0370 ;
        RECT 6.9040 42.9435 6.9300 44.0370 ;
        RECT 6.7960 42.9435 6.8220 44.0370 ;
        RECT 6.6880 42.9435 6.7140 44.0370 ;
        RECT 6.5800 42.9435 6.6060 44.0370 ;
        RECT 6.4720 42.9435 6.4980 44.0370 ;
        RECT 6.3640 42.9435 6.3900 44.0370 ;
        RECT 6.2560 42.9435 6.2820 44.0370 ;
        RECT 6.1480 42.9435 6.1740 44.0370 ;
        RECT 6.0400 42.9435 6.0660 44.0370 ;
        RECT 5.9320 42.9435 5.9580 44.0370 ;
        RECT 5.8240 42.9435 5.8500 44.0370 ;
        RECT 5.7160 42.9435 5.7420 44.0370 ;
        RECT 5.6080 42.9435 5.6340 44.0370 ;
        RECT 5.5000 42.9435 5.5260 44.0370 ;
        RECT 5.3920 42.9435 5.4180 44.0370 ;
        RECT 5.2840 42.9435 5.3100 44.0370 ;
        RECT 5.1760 42.9435 5.2020 44.0370 ;
        RECT 5.0680 42.9435 5.0940 44.0370 ;
        RECT 4.9600 42.9435 4.9860 44.0370 ;
        RECT 4.8520 42.9435 4.8780 44.0370 ;
        RECT 4.7440 42.9435 4.7700 44.0370 ;
        RECT 4.6360 42.9435 4.6620 44.0370 ;
        RECT 4.5280 42.9435 4.5540 44.0370 ;
        RECT 4.4200 42.9435 4.4460 44.0370 ;
        RECT 4.3120 42.9435 4.3380 44.0370 ;
        RECT 4.2040 42.9435 4.2300 44.0370 ;
        RECT 4.0960 42.9435 4.1220 44.0370 ;
        RECT 3.9880 42.9435 4.0140 44.0370 ;
        RECT 3.8800 42.9435 3.9060 44.0370 ;
        RECT 3.7720 42.9435 3.7980 44.0370 ;
        RECT 3.6640 42.9435 3.6900 44.0370 ;
        RECT 3.5560 42.9435 3.5820 44.0370 ;
        RECT 3.4480 42.9435 3.4740 44.0370 ;
        RECT 3.3400 42.9435 3.3660 44.0370 ;
        RECT 3.2320 42.9435 3.2580 44.0370 ;
        RECT 3.1240 42.9435 3.1500 44.0370 ;
        RECT 3.0160 42.9435 3.0420 44.0370 ;
        RECT 2.9080 42.9435 2.9340 44.0370 ;
        RECT 2.8000 42.9435 2.8260 44.0370 ;
        RECT 2.6920 42.9435 2.7180 44.0370 ;
        RECT 2.5840 42.9435 2.6100 44.0370 ;
        RECT 2.4760 42.9435 2.5020 44.0370 ;
        RECT 2.3680 42.9435 2.3940 44.0370 ;
        RECT 2.2600 42.9435 2.2860 44.0370 ;
        RECT 2.1520 42.9435 2.1780 44.0370 ;
        RECT 2.0440 42.9435 2.0700 44.0370 ;
        RECT 1.9360 42.9435 1.9620 44.0370 ;
        RECT 1.8280 42.9435 1.8540 44.0370 ;
        RECT 1.7200 42.9435 1.7460 44.0370 ;
        RECT 1.6120 42.9435 1.6380 44.0370 ;
        RECT 1.5040 42.9435 1.5300 44.0370 ;
        RECT 1.3960 42.9435 1.4220 44.0370 ;
        RECT 1.2880 42.9435 1.3140 44.0370 ;
        RECT 1.1800 42.9435 1.2060 44.0370 ;
        RECT 1.0720 42.9435 1.0980 44.0370 ;
        RECT 0.9640 42.9435 0.9900 44.0370 ;
        RECT 0.8560 42.9435 0.8820 44.0370 ;
        RECT 0.7480 42.9435 0.7740 44.0370 ;
        RECT 0.6400 42.9435 0.6660 44.0370 ;
        RECT 0.5320 42.9435 0.5580 44.0370 ;
        RECT 0.4240 42.9435 0.4500 44.0370 ;
        RECT 0.3160 42.9435 0.3420 44.0370 ;
        RECT 0.2080 42.9435 0.2340 44.0370 ;
        RECT 0.0050 42.9435 0.0900 44.0370 ;
        RECT 8.6410 44.0235 8.7690 45.1170 ;
        RECT 8.6270 44.6890 8.7690 45.0115 ;
        RECT 8.4790 44.4160 8.5410 45.1170 ;
        RECT 8.4650 44.7255 8.5410 44.8790 ;
        RECT 8.4790 44.0235 8.5050 45.1170 ;
        RECT 8.4790 44.1445 8.5190 44.3840 ;
        RECT 8.4790 44.0235 8.5410 44.1125 ;
        RECT 8.1820 44.4740 8.3880 45.1170 ;
        RECT 8.3620 44.0235 8.3880 45.1170 ;
        RECT 8.1820 44.7510 8.4020 45.0090 ;
        RECT 8.1820 44.0235 8.2800 45.1170 ;
        RECT 7.7650 44.0235 7.8480 45.1170 ;
        RECT 7.7650 44.1120 7.8620 45.0475 ;
        RECT 16.4440 44.0235 16.5290 45.1170 ;
        RECT 16.3000 44.0235 16.3260 45.1170 ;
        RECT 16.1920 44.0235 16.2180 45.1170 ;
        RECT 16.0840 44.0235 16.1100 45.1170 ;
        RECT 15.9760 44.0235 16.0020 45.1170 ;
        RECT 15.8680 44.0235 15.8940 45.1170 ;
        RECT 15.7600 44.0235 15.7860 45.1170 ;
        RECT 15.6520 44.0235 15.6780 45.1170 ;
        RECT 15.5440 44.0235 15.5700 45.1170 ;
        RECT 15.4360 44.0235 15.4620 45.1170 ;
        RECT 15.3280 44.0235 15.3540 45.1170 ;
        RECT 15.2200 44.0235 15.2460 45.1170 ;
        RECT 15.1120 44.0235 15.1380 45.1170 ;
        RECT 15.0040 44.0235 15.0300 45.1170 ;
        RECT 14.8960 44.0235 14.9220 45.1170 ;
        RECT 14.7880 44.0235 14.8140 45.1170 ;
        RECT 14.6800 44.0235 14.7060 45.1170 ;
        RECT 14.5720 44.0235 14.5980 45.1170 ;
        RECT 14.4640 44.0235 14.4900 45.1170 ;
        RECT 14.3560 44.0235 14.3820 45.1170 ;
        RECT 14.2480 44.0235 14.2740 45.1170 ;
        RECT 14.1400 44.0235 14.1660 45.1170 ;
        RECT 14.0320 44.0235 14.0580 45.1170 ;
        RECT 13.9240 44.0235 13.9500 45.1170 ;
        RECT 13.8160 44.0235 13.8420 45.1170 ;
        RECT 13.7080 44.0235 13.7340 45.1170 ;
        RECT 13.6000 44.0235 13.6260 45.1170 ;
        RECT 13.4920 44.0235 13.5180 45.1170 ;
        RECT 13.3840 44.0235 13.4100 45.1170 ;
        RECT 13.2760 44.0235 13.3020 45.1170 ;
        RECT 13.1680 44.0235 13.1940 45.1170 ;
        RECT 13.0600 44.0235 13.0860 45.1170 ;
        RECT 12.9520 44.0235 12.9780 45.1170 ;
        RECT 12.8440 44.0235 12.8700 45.1170 ;
        RECT 12.7360 44.0235 12.7620 45.1170 ;
        RECT 12.6280 44.0235 12.6540 45.1170 ;
        RECT 12.5200 44.0235 12.5460 45.1170 ;
        RECT 12.4120 44.0235 12.4380 45.1170 ;
        RECT 12.3040 44.0235 12.3300 45.1170 ;
        RECT 12.1960 44.0235 12.2220 45.1170 ;
        RECT 12.0880 44.0235 12.1140 45.1170 ;
        RECT 11.9800 44.0235 12.0060 45.1170 ;
        RECT 11.8720 44.0235 11.8980 45.1170 ;
        RECT 11.7640 44.0235 11.7900 45.1170 ;
        RECT 11.6560 44.0235 11.6820 45.1170 ;
        RECT 11.5480 44.0235 11.5740 45.1170 ;
        RECT 11.4400 44.0235 11.4660 45.1170 ;
        RECT 11.3320 44.0235 11.3580 45.1170 ;
        RECT 11.2240 44.0235 11.2500 45.1170 ;
        RECT 11.1160 44.0235 11.1420 45.1170 ;
        RECT 11.0080 44.0235 11.0340 45.1170 ;
        RECT 10.9000 44.0235 10.9260 45.1170 ;
        RECT 10.7920 44.0235 10.8180 45.1170 ;
        RECT 10.6840 44.0235 10.7100 45.1170 ;
        RECT 10.5760 44.0235 10.6020 45.1170 ;
        RECT 10.4680 44.0235 10.4940 45.1170 ;
        RECT 10.3600 44.0235 10.3860 45.1170 ;
        RECT 10.2520 44.0235 10.2780 45.1170 ;
        RECT 10.1440 44.0235 10.1700 45.1170 ;
        RECT 10.0360 44.0235 10.0620 45.1170 ;
        RECT 9.9280 44.0235 9.9540 45.1170 ;
        RECT 9.8200 44.0235 9.8460 45.1170 ;
        RECT 9.7120 44.0235 9.7380 45.1170 ;
        RECT 9.6040 44.0235 9.6300 45.1170 ;
        RECT 9.4960 44.0235 9.5220 45.1170 ;
        RECT 9.3880 44.0235 9.4140 45.1170 ;
        RECT 9.1750 44.0235 9.2520 45.1170 ;
        RECT 7.2820 44.0235 7.3590 45.1170 ;
        RECT 7.1200 44.0235 7.1460 45.1170 ;
        RECT 7.0120 44.0235 7.0380 45.1170 ;
        RECT 6.9040 44.0235 6.9300 45.1170 ;
        RECT 6.7960 44.0235 6.8220 45.1170 ;
        RECT 6.6880 44.0235 6.7140 45.1170 ;
        RECT 6.5800 44.0235 6.6060 45.1170 ;
        RECT 6.4720 44.0235 6.4980 45.1170 ;
        RECT 6.3640 44.0235 6.3900 45.1170 ;
        RECT 6.2560 44.0235 6.2820 45.1170 ;
        RECT 6.1480 44.0235 6.1740 45.1170 ;
        RECT 6.0400 44.0235 6.0660 45.1170 ;
        RECT 5.9320 44.0235 5.9580 45.1170 ;
        RECT 5.8240 44.0235 5.8500 45.1170 ;
        RECT 5.7160 44.0235 5.7420 45.1170 ;
        RECT 5.6080 44.0235 5.6340 45.1170 ;
        RECT 5.5000 44.0235 5.5260 45.1170 ;
        RECT 5.3920 44.0235 5.4180 45.1170 ;
        RECT 5.2840 44.0235 5.3100 45.1170 ;
        RECT 5.1760 44.0235 5.2020 45.1170 ;
        RECT 5.0680 44.0235 5.0940 45.1170 ;
        RECT 4.9600 44.0235 4.9860 45.1170 ;
        RECT 4.8520 44.0235 4.8780 45.1170 ;
        RECT 4.7440 44.0235 4.7700 45.1170 ;
        RECT 4.6360 44.0235 4.6620 45.1170 ;
        RECT 4.5280 44.0235 4.5540 45.1170 ;
        RECT 4.4200 44.0235 4.4460 45.1170 ;
        RECT 4.3120 44.0235 4.3380 45.1170 ;
        RECT 4.2040 44.0235 4.2300 45.1170 ;
        RECT 4.0960 44.0235 4.1220 45.1170 ;
        RECT 3.9880 44.0235 4.0140 45.1170 ;
        RECT 3.8800 44.0235 3.9060 45.1170 ;
        RECT 3.7720 44.0235 3.7980 45.1170 ;
        RECT 3.6640 44.0235 3.6900 45.1170 ;
        RECT 3.5560 44.0235 3.5820 45.1170 ;
        RECT 3.4480 44.0235 3.4740 45.1170 ;
        RECT 3.3400 44.0235 3.3660 45.1170 ;
        RECT 3.2320 44.0235 3.2580 45.1170 ;
        RECT 3.1240 44.0235 3.1500 45.1170 ;
        RECT 3.0160 44.0235 3.0420 45.1170 ;
        RECT 2.9080 44.0235 2.9340 45.1170 ;
        RECT 2.8000 44.0235 2.8260 45.1170 ;
        RECT 2.6920 44.0235 2.7180 45.1170 ;
        RECT 2.5840 44.0235 2.6100 45.1170 ;
        RECT 2.4760 44.0235 2.5020 45.1170 ;
        RECT 2.3680 44.0235 2.3940 45.1170 ;
        RECT 2.2600 44.0235 2.2860 45.1170 ;
        RECT 2.1520 44.0235 2.1780 45.1170 ;
        RECT 2.0440 44.0235 2.0700 45.1170 ;
        RECT 1.9360 44.0235 1.9620 45.1170 ;
        RECT 1.8280 44.0235 1.8540 45.1170 ;
        RECT 1.7200 44.0235 1.7460 45.1170 ;
        RECT 1.6120 44.0235 1.6380 45.1170 ;
        RECT 1.5040 44.0235 1.5300 45.1170 ;
        RECT 1.3960 44.0235 1.4220 45.1170 ;
        RECT 1.2880 44.0235 1.3140 45.1170 ;
        RECT 1.1800 44.0235 1.2060 45.1170 ;
        RECT 1.0720 44.0235 1.0980 45.1170 ;
        RECT 0.9640 44.0235 0.9900 45.1170 ;
        RECT 0.8560 44.0235 0.8820 45.1170 ;
        RECT 0.7480 44.0235 0.7740 45.1170 ;
        RECT 0.6400 44.0235 0.6660 45.1170 ;
        RECT 0.5320 44.0235 0.5580 45.1170 ;
        RECT 0.4240 44.0235 0.4500 45.1170 ;
        RECT 0.3160 44.0235 0.3420 45.1170 ;
        RECT 0.2080 44.0235 0.2340 45.1170 ;
        RECT 0.0050 44.0235 0.0900 45.1170 ;
        RECT 8.6410 45.1035 8.7690 46.1970 ;
        RECT 8.6270 45.7690 8.7690 46.0915 ;
        RECT 8.4790 45.4960 8.5410 46.1970 ;
        RECT 8.4650 45.8055 8.5410 45.9590 ;
        RECT 8.4790 45.1035 8.5050 46.1970 ;
        RECT 8.4790 45.2245 8.5190 45.4640 ;
        RECT 8.4790 45.1035 8.5410 45.1925 ;
        RECT 8.1820 45.5540 8.3880 46.1970 ;
        RECT 8.3620 45.1035 8.3880 46.1970 ;
        RECT 8.1820 45.8310 8.4020 46.0890 ;
        RECT 8.1820 45.1035 8.2800 46.1970 ;
        RECT 7.7650 45.1035 7.8480 46.1970 ;
        RECT 7.7650 45.1920 7.8620 46.1275 ;
        RECT 16.4440 45.1035 16.5290 46.1970 ;
        RECT 16.3000 45.1035 16.3260 46.1970 ;
        RECT 16.1920 45.1035 16.2180 46.1970 ;
        RECT 16.0840 45.1035 16.1100 46.1970 ;
        RECT 15.9760 45.1035 16.0020 46.1970 ;
        RECT 15.8680 45.1035 15.8940 46.1970 ;
        RECT 15.7600 45.1035 15.7860 46.1970 ;
        RECT 15.6520 45.1035 15.6780 46.1970 ;
        RECT 15.5440 45.1035 15.5700 46.1970 ;
        RECT 15.4360 45.1035 15.4620 46.1970 ;
        RECT 15.3280 45.1035 15.3540 46.1970 ;
        RECT 15.2200 45.1035 15.2460 46.1970 ;
        RECT 15.1120 45.1035 15.1380 46.1970 ;
        RECT 15.0040 45.1035 15.0300 46.1970 ;
        RECT 14.8960 45.1035 14.9220 46.1970 ;
        RECT 14.7880 45.1035 14.8140 46.1970 ;
        RECT 14.6800 45.1035 14.7060 46.1970 ;
        RECT 14.5720 45.1035 14.5980 46.1970 ;
        RECT 14.4640 45.1035 14.4900 46.1970 ;
        RECT 14.3560 45.1035 14.3820 46.1970 ;
        RECT 14.2480 45.1035 14.2740 46.1970 ;
        RECT 14.1400 45.1035 14.1660 46.1970 ;
        RECT 14.0320 45.1035 14.0580 46.1970 ;
        RECT 13.9240 45.1035 13.9500 46.1970 ;
        RECT 13.8160 45.1035 13.8420 46.1970 ;
        RECT 13.7080 45.1035 13.7340 46.1970 ;
        RECT 13.6000 45.1035 13.6260 46.1970 ;
        RECT 13.4920 45.1035 13.5180 46.1970 ;
        RECT 13.3840 45.1035 13.4100 46.1970 ;
        RECT 13.2760 45.1035 13.3020 46.1970 ;
        RECT 13.1680 45.1035 13.1940 46.1970 ;
        RECT 13.0600 45.1035 13.0860 46.1970 ;
        RECT 12.9520 45.1035 12.9780 46.1970 ;
        RECT 12.8440 45.1035 12.8700 46.1970 ;
        RECT 12.7360 45.1035 12.7620 46.1970 ;
        RECT 12.6280 45.1035 12.6540 46.1970 ;
        RECT 12.5200 45.1035 12.5460 46.1970 ;
        RECT 12.4120 45.1035 12.4380 46.1970 ;
        RECT 12.3040 45.1035 12.3300 46.1970 ;
        RECT 12.1960 45.1035 12.2220 46.1970 ;
        RECT 12.0880 45.1035 12.1140 46.1970 ;
        RECT 11.9800 45.1035 12.0060 46.1970 ;
        RECT 11.8720 45.1035 11.8980 46.1970 ;
        RECT 11.7640 45.1035 11.7900 46.1970 ;
        RECT 11.6560 45.1035 11.6820 46.1970 ;
        RECT 11.5480 45.1035 11.5740 46.1970 ;
        RECT 11.4400 45.1035 11.4660 46.1970 ;
        RECT 11.3320 45.1035 11.3580 46.1970 ;
        RECT 11.2240 45.1035 11.2500 46.1970 ;
        RECT 11.1160 45.1035 11.1420 46.1970 ;
        RECT 11.0080 45.1035 11.0340 46.1970 ;
        RECT 10.9000 45.1035 10.9260 46.1970 ;
        RECT 10.7920 45.1035 10.8180 46.1970 ;
        RECT 10.6840 45.1035 10.7100 46.1970 ;
        RECT 10.5760 45.1035 10.6020 46.1970 ;
        RECT 10.4680 45.1035 10.4940 46.1970 ;
        RECT 10.3600 45.1035 10.3860 46.1970 ;
        RECT 10.2520 45.1035 10.2780 46.1970 ;
        RECT 10.1440 45.1035 10.1700 46.1970 ;
        RECT 10.0360 45.1035 10.0620 46.1970 ;
        RECT 9.9280 45.1035 9.9540 46.1970 ;
        RECT 9.8200 45.1035 9.8460 46.1970 ;
        RECT 9.7120 45.1035 9.7380 46.1970 ;
        RECT 9.6040 45.1035 9.6300 46.1970 ;
        RECT 9.4960 45.1035 9.5220 46.1970 ;
        RECT 9.3880 45.1035 9.4140 46.1970 ;
        RECT 9.1750 45.1035 9.2520 46.1970 ;
        RECT 7.2820 45.1035 7.3590 46.1970 ;
        RECT 7.1200 45.1035 7.1460 46.1970 ;
        RECT 7.0120 45.1035 7.0380 46.1970 ;
        RECT 6.9040 45.1035 6.9300 46.1970 ;
        RECT 6.7960 45.1035 6.8220 46.1970 ;
        RECT 6.6880 45.1035 6.7140 46.1970 ;
        RECT 6.5800 45.1035 6.6060 46.1970 ;
        RECT 6.4720 45.1035 6.4980 46.1970 ;
        RECT 6.3640 45.1035 6.3900 46.1970 ;
        RECT 6.2560 45.1035 6.2820 46.1970 ;
        RECT 6.1480 45.1035 6.1740 46.1970 ;
        RECT 6.0400 45.1035 6.0660 46.1970 ;
        RECT 5.9320 45.1035 5.9580 46.1970 ;
        RECT 5.8240 45.1035 5.8500 46.1970 ;
        RECT 5.7160 45.1035 5.7420 46.1970 ;
        RECT 5.6080 45.1035 5.6340 46.1970 ;
        RECT 5.5000 45.1035 5.5260 46.1970 ;
        RECT 5.3920 45.1035 5.4180 46.1970 ;
        RECT 5.2840 45.1035 5.3100 46.1970 ;
        RECT 5.1760 45.1035 5.2020 46.1970 ;
        RECT 5.0680 45.1035 5.0940 46.1970 ;
        RECT 4.9600 45.1035 4.9860 46.1970 ;
        RECT 4.8520 45.1035 4.8780 46.1970 ;
        RECT 4.7440 45.1035 4.7700 46.1970 ;
        RECT 4.6360 45.1035 4.6620 46.1970 ;
        RECT 4.5280 45.1035 4.5540 46.1970 ;
        RECT 4.4200 45.1035 4.4460 46.1970 ;
        RECT 4.3120 45.1035 4.3380 46.1970 ;
        RECT 4.2040 45.1035 4.2300 46.1970 ;
        RECT 4.0960 45.1035 4.1220 46.1970 ;
        RECT 3.9880 45.1035 4.0140 46.1970 ;
        RECT 3.8800 45.1035 3.9060 46.1970 ;
        RECT 3.7720 45.1035 3.7980 46.1970 ;
        RECT 3.6640 45.1035 3.6900 46.1970 ;
        RECT 3.5560 45.1035 3.5820 46.1970 ;
        RECT 3.4480 45.1035 3.4740 46.1970 ;
        RECT 3.3400 45.1035 3.3660 46.1970 ;
        RECT 3.2320 45.1035 3.2580 46.1970 ;
        RECT 3.1240 45.1035 3.1500 46.1970 ;
        RECT 3.0160 45.1035 3.0420 46.1970 ;
        RECT 2.9080 45.1035 2.9340 46.1970 ;
        RECT 2.8000 45.1035 2.8260 46.1970 ;
        RECT 2.6920 45.1035 2.7180 46.1970 ;
        RECT 2.5840 45.1035 2.6100 46.1970 ;
        RECT 2.4760 45.1035 2.5020 46.1970 ;
        RECT 2.3680 45.1035 2.3940 46.1970 ;
        RECT 2.2600 45.1035 2.2860 46.1970 ;
        RECT 2.1520 45.1035 2.1780 46.1970 ;
        RECT 2.0440 45.1035 2.0700 46.1970 ;
        RECT 1.9360 45.1035 1.9620 46.1970 ;
        RECT 1.8280 45.1035 1.8540 46.1970 ;
        RECT 1.7200 45.1035 1.7460 46.1970 ;
        RECT 1.6120 45.1035 1.6380 46.1970 ;
        RECT 1.5040 45.1035 1.5300 46.1970 ;
        RECT 1.3960 45.1035 1.4220 46.1970 ;
        RECT 1.2880 45.1035 1.3140 46.1970 ;
        RECT 1.1800 45.1035 1.2060 46.1970 ;
        RECT 1.0720 45.1035 1.0980 46.1970 ;
        RECT 0.9640 45.1035 0.9900 46.1970 ;
        RECT 0.8560 45.1035 0.8820 46.1970 ;
        RECT 0.7480 45.1035 0.7740 46.1970 ;
        RECT 0.6400 45.1035 0.6660 46.1970 ;
        RECT 0.5320 45.1035 0.5580 46.1970 ;
        RECT 0.4240 45.1035 0.4500 46.1970 ;
        RECT 0.3160 45.1035 0.3420 46.1970 ;
        RECT 0.2080 45.1035 0.2340 46.1970 ;
        RECT 0.0050 45.1035 0.0900 46.1970 ;
        RECT 8.6410 46.1835 8.7690 47.2770 ;
        RECT 8.6270 46.8490 8.7690 47.1715 ;
        RECT 8.4790 46.5760 8.5410 47.2770 ;
        RECT 8.4650 46.8855 8.5410 47.0390 ;
        RECT 8.4790 46.1835 8.5050 47.2770 ;
        RECT 8.4790 46.3045 8.5190 46.5440 ;
        RECT 8.4790 46.1835 8.5410 46.2725 ;
        RECT 8.1820 46.6340 8.3880 47.2770 ;
        RECT 8.3620 46.1835 8.3880 47.2770 ;
        RECT 8.1820 46.9110 8.4020 47.1690 ;
        RECT 8.1820 46.1835 8.2800 47.2770 ;
        RECT 7.7650 46.1835 7.8480 47.2770 ;
        RECT 7.7650 46.2720 7.8620 47.2075 ;
        RECT 16.4440 46.1835 16.5290 47.2770 ;
        RECT 16.3000 46.1835 16.3260 47.2770 ;
        RECT 16.1920 46.1835 16.2180 47.2770 ;
        RECT 16.0840 46.1835 16.1100 47.2770 ;
        RECT 15.9760 46.1835 16.0020 47.2770 ;
        RECT 15.8680 46.1835 15.8940 47.2770 ;
        RECT 15.7600 46.1835 15.7860 47.2770 ;
        RECT 15.6520 46.1835 15.6780 47.2770 ;
        RECT 15.5440 46.1835 15.5700 47.2770 ;
        RECT 15.4360 46.1835 15.4620 47.2770 ;
        RECT 15.3280 46.1835 15.3540 47.2770 ;
        RECT 15.2200 46.1835 15.2460 47.2770 ;
        RECT 15.1120 46.1835 15.1380 47.2770 ;
        RECT 15.0040 46.1835 15.0300 47.2770 ;
        RECT 14.8960 46.1835 14.9220 47.2770 ;
        RECT 14.7880 46.1835 14.8140 47.2770 ;
        RECT 14.6800 46.1835 14.7060 47.2770 ;
        RECT 14.5720 46.1835 14.5980 47.2770 ;
        RECT 14.4640 46.1835 14.4900 47.2770 ;
        RECT 14.3560 46.1835 14.3820 47.2770 ;
        RECT 14.2480 46.1835 14.2740 47.2770 ;
        RECT 14.1400 46.1835 14.1660 47.2770 ;
        RECT 14.0320 46.1835 14.0580 47.2770 ;
        RECT 13.9240 46.1835 13.9500 47.2770 ;
        RECT 13.8160 46.1835 13.8420 47.2770 ;
        RECT 13.7080 46.1835 13.7340 47.2770 ;
        RECT 13.6000 46.1835 13.6260 47.2770 ;
        RECT 13.4920 46.1835 13.5180 47.2770 ;
        RECT 13.3840 46.1835 13.4100 47.2770 ;
        RECT 13.2760 46.1835 13.3020 47.2770 ;
        RECT 13.1680 46.1835 13.1940 47.2770 ;
        RECT 13.0600 46.1835 13.0860 47.2770 ;
        RECT 12.9520 46.1835 12.9780 47.2770 ;
        RECT 12.8440 46.1835 12.8700 47.2770 ;
        RECT 12.7360 46.1835 12.7620 47.2770 ;
        RECT 12.6280 46.1835 12.6540 47.2770 ;
        RECT 12.5200 46.1835 12.5460 47.2770 ;
        RECT 12.4120 46.1835 12.4380 47.2770 ;
        RECT 12.3040 46.1835 12.3300 47.2770 ;
        RECT 12.1960 46.1835 12.2220 47.2770 ;
        RECT 12.0880 46.1835 12.1140 47.2770 ;
        RECT 11.9800 46.1835 12.0060 47.2770 ;
        RECT 11.8720 46.1835 11.8980 47.2770 ;
        RECT 11.7640 46.1835 11.7900 47.2770 ;
        RECT 11.6560 46.1835 11.6820 47.2770 ;
        RECT 11.5480 46.1835 11.5740 47.2770 ;
        RECT 11.4400 46.1835 11.4660 47.2770 ;
        RECT 11.3320 46.1835 11.3580 47.2770 ;
        RECT 11.2240 46.1835 11.2500 47.2770 ;
        RECT 11.1160 46.1835 11.1420 47.2770 ;
        RECT 11.0080 46.1835 11.0340 47.2770 ;
        RECT 10.9000 46.1835 10.9260 47.2770 ;
        RECT 10.7920 46.1835 10.8180 47.2770 ;
        RECT 10.6840 46.1835 10.7100 47.2770 ;
        RECT 10.5760 46.1835 10.6020 47.2770 ;
        RECT 10.4680 46.1835 10.4940 47.2770 ;
        RECT 10.3600 46.1835 10.3860 47.2770 ;
        RECT 10.2520 46.1835 10.2780 47.2770 ;
        RECT 10.1440 46.1835 10.1700 47.2770 ;
        RECT 10.0360 46.1835 10.0620 47.2770 ;
        RECT 9.9280 46.1835 9.9540 47.2770 ;
        RECT 9.8200 46.1835 9.8460 47.2770 ;
        RECT 9.7120 46.1835 9.7380 47.2770 ;
        RECT 9.6040 46.1835 9.6300 47.2770 ;
        RECT 9.4960 46.1835 9.5220 47.2770 ;
        RECT 9.3880 46.1835 9.4140 47.2770 ;
        RECT 9.1750 46.1835 9.2520 47.2770 ;
        RECT 7.2820 46.1835 7.3590 47.2770 ;
        RECT 7.1200 46.1835 7.1460 47.2770 ;
        RECT 7.0120 46.1835 7.0380 47.2770 ;
        RECT 6.9040 46.1835 6.9300 47.2770 ;
        RECT 6.7960 46.1835 6.8220 47.2770 ;
        RECT 6.6880 46.1835 6.7140 47.2770 ;
        RECT 6.5800 46.1835 6.6060 47.2770 ;
        RECT 6.4720 46.1835 6.4980 47.2770 ;
        RECT 6.3640 46.1835 6.3900 47.2770 ;
        RECT 6.2560 46.1835 6.2820 47.2770 ;
        RECT 6.1480 46.1835 6.1740 47.2770 ;
        RECT 6.0400 46.1835 6.0660 47.2770 ;
        RECT 5.9320 46.1835 5.9580 47.2770 ;
        RECT 5.8240 46.1835 5.8500 47.2770 ;
        RECT 5.7160 46.1835 5.7420 47.2770 ;
        RECT 5.6080 46.1835 5.6340 47.2770 ;
        RECT 5.5000 46.1835 5.5260 47.2770 ;
        RECT 5.3920 46.1835 5.4180 47.2770 ;
        RECT 5.2840 46.1835 5.3100 47.2770 ;
        RECT 5.1760 46.1835 5.2020 47.2770 ;
        RECT 5.0680 46.1835 5.0940 47.2770 ;
        RECT 4.9600 46.1835 4.9860 47.2770 ;
        RECT 4.8520 46.1835 4.8780 47.2770 ;
        RECT 4.7440 46.1835 4.7700 47.2770 ;
        RECT 4.6360 46.1835 4.6620 47.2770 ;
        RECT 4.5280 46.1835 4.5540 47.2770 ;
        RECT 4.4200 46.1835 4.4460 47.2770 ;
        RECT 4.3120 46.1835 4.3380 47.2770 ;
        RECT 4.2040 46.1835 4.2300 47.2770 ;
        RECT 4.0960 46.1835 4.1220 47.2770 ;
        RECT 3.9880 46.1835 4.0140 47.2770 ;
        RECT 3.8800 46.1835 3.9060 47.2770 ;
        RECT 3.7720 46.1835 3.7980 47.2770 ;
        RECT 3.6640 46.1835 3.6900 47.2770 ;
        RECT 3.5560 46.1835 3.5820 47.2770 ;
        RECT 3.4480 46.1835 3.4740 47.2770 ;
        RECT 3.3400 46.1835 3.3660 47.2770 ;
        RECT 3.2320 46.1835 3.2580 47.2770 ;
        RECT 3.1240 46.1835 3.1500 47.2770 ;
        RECT 3.0160 46.1835 3.0420 47.2770 ;
        RECT 2.9080 46.1835 2.9340 47.2770 ;
        RECT 2.8000 46.1835 2.8260 47.2770 ;
        RECT 2.6920 46.1835 2.7180 47.2770 ;
        RECT 2.5840 46.1835 2.6100 47.2770 ;
        RECT 2.4760 46.1835 2.5020 47.2770 ;
        RECT 2.3680 46.1835 2.3940 47.2770 ;
        RECT 2.2600 46.1835 2.2860 47.2770 ;
        RECT 2.1520 46.1835 2.1780 47.2770 ;
        RECT 2.0440 46.1835 2.0700 47.2770 ;
        RECT 1.9360 46.1835 1.9620 47.2770 ;
        RECT 1.8280 46.1835 1.8540 47.2770 ;
        RECT 1.7200 46.1835 1.7460 47.2770 ;
        RECT 1.6120 46.1835 1.6380 47.2770 ;
        RECT 1.5040 46.1835 1.5300 47.2770 ;
        RECT 1.3960 46.1835 1.4220 47.2770 ;
        RECT 1.2880 46.1835 1.3140 47.2770 ;
        RECT 1.1800 46.1835 1.2060 47.2770 ;
        RECT 1.0720 46.1835 1.0980 47.2770 ;
        RECT 0.9640 46.1835 0.9900 47.2770 ;
        RECT 0.8560 46.1835 0.8820 47.2770 ;
        RECT 0.7480 46.1835 0.7740 47.2770 ;
        RECT 0.6400 46.1835 0.6660 47.2770 ;
        RECT 0.5320 46.1835 0.5580 47.2770 ;
        RECT 0.4240 46.1835 0.4500 47.2770 ;
        RECT 0.3160 46.1835 0.3420 47.2770 ;
        RECT 0.2080 46.1835 0.2340 47.2770 ;
        RECT 0.0050 46.1835 0.0900 47.2770 ;
        RECT 8.6410 47.2635 8.7690 48.3570 ;
        RECT 8.6270 47.9290 8.7690 48.2515 ;
        RECT 8.4790 47.6560 8.5410 48.3570 ;
        RECT 8.4650 47.9655 8.5410 48.1190 ;
        RECT 8.4790 47.2635 8.5050 48.3570 ;
        RECT 8.4790 47.3845 8.5190 47.6240 ;
        RECT 8.4790 47.2635 8.5410 47.3525 ;
        RECT 8.1820 47.7140 8.3880 48.3570 ;
        RECT 8.3620 47.2635 8.3880 48.3570 ;
        RECT 8.1820 47.9910 8.4020 48.2490 ;
        RECT 8.1820 47.2635 8.2800 48.3570 ;
        RECT 7.7650 47.2635 7.8480 48.3570 ;
        RECT 7.7650 47.3520 7.8620 48.2875 ;
        RECT 16.4440 47.2635 16.5290 48.3570 ;
        RECT 16.3000 47.2635 16.3260 48.3570 ;
        RECT 16.1920 47.2635 16.2180 48.3570 ;
        RECT 16.0840 47.2635 16.1100 48.3570 ;
        RECT 15.9760 47.2635 16.0020 48.3570 ;
        RECT 15.8680 47.2635 15.8940 48.3570 ;
        RECT 15.7600 47.2635 15.7860 48.3570 ;
        RECT 15.6520 47.2635 15.6780 48.3570 ;
        RECT 15.5440 47.2635 15.5700 48.3570 ;
        RECT 15.4360 47.2635 15.4620 48.3570 ;
        RECT 15.3280 47.2635 15.3540 48.3570 ;
        RECT 15.2200 47.2635 15.2460 48.3570 ;
        RECT 15.1120 47.2635 15.1380 48.3570 ;
        RECT 15.0040 47.2635 15.0300 48.3570 ;
        RECT 14.8960 47.2635 14.9220 48.3570 ;
        RECT 14.7880 47.2635 14.8140 48.3570 ;
        RECT 14.6800 47.2635 14.7060 48.3570 ;
        RECT 14.5720 47.2635 14.5980 48.3570 ;
        RECT 14.4640 47.2635 14.4900 48.3570 ;
        RECT 14.3560 47.2635 14.3820 48.3570 ;
        RECT 14.2480 47.2635 14.2740 48.3570 ;
        RECT 14.1400 47.2635 14.1660 48.3570 ;
        RECT 14.0320 47.2635 14.0580 48.3570 ;
        RECT 13.9240 47.2635 13.9500 48.3570 ;
        RECT 13.8160 47.2635 13.8420 48.3570 ;
        RECT 13.7080 47.2635 13.7340 48.3570 ;
        RECT 13.6000 47.2635 13.6260 48.3570 ;
        RECT 13.4920 47.2635 13.5180 48.3570 ;
        RECT 13.3840 47.2635 13.4100 48.3570 ;
        RECT 13.2760 47.2635 13.3020 48.3570 ;
        RECT 13.1680 47.2635 13.1940 48.3570 ;
        RECT 13.0600 47.2635 13.0860 48.3570 ;
        RECT 12.9520 47.2635 12.9780 48.3570 ;
        RECT 12.8440 47.2635 12.8700 48.3570 ;
        RECT 12.7360 47.2635 12.7620 48.3570 ;
        RECT 12.6280 47.2635 12.6540 48.3570 ;
        RECT 12.5200 47.2635 12.5460 48.3570 ;
        RECT 12.4120 47.2635 12.4380 48.3570 ;
        RECT 12.3040 47.2635 12.3300 48.3570 ;
        RECT 12.1960 47.2635 12.2220 48.3570 ;
        RECT 12.0880 47.2635 12.1140 48.3570 ;
        RECT 11.9800 47.2635 12.0060 48.3570 ;
        RECT 11.8720 47.2635 11.8980 48.3570 ;
        RECT 11.7640 47.2635 11.7900 48.3570 ;
        RECT 11.6560 47.2635 11.6820 48.3570 ;
        RECT 11.5480 47.2635 11.5740 48.3570 ;
        RECT 11.4400 47.2635 11.4660 48.3570 ;
        RECT 11.3320 47.2635 11.3580 48.3570 ;
        RECT 11.2240 47.2635 11.2500 48.3570 ;
        RECT 11.1160 47.2635 11.1420 48.3570 ;
        RECT 11.0080 47.2635 11.0340 48.3570 ;
        RECT 10.9000 47.2635 10.9260 48.3570 ;
        RECT 10.7920 47.2635 10.8180 48.3570 ;
        RECT 10.6840 47.2635 10.7100 48.3570 ;
        RECT 10.5760 47.2635 10.6020 48.3570 ;
        RECT 10.4680 47.2635 10.4940 48.3570 ;
        RECT 10.3600 47.2635 10.3860 48.3570 ;
        RECT 10.2520 47.2635 10.2780 48.3570 ;
        RECT 10.1440 47.2635 10.1700 48.3570 ;
        RECT 10.0360 47.2635 10.0620 48.3570 ;
        RECT 9.9280 47.2635 9.9540 48.3570 ;
        RECT 9.8200 47.2635 9.8460 48.3570 ;
        RECT 9.7120 47.2635 9.7380 48.3570 ;
        RECT 9.6040 47.2635 9.6300 48.3570 ;
        RECT 9.4960 47.2635 9.5220 48.3570 ;
        RECT 9.3880 47.2635 9.4140 48.3570 ;
        RECT 9.1750 47.2635 9.2520 48.3570 ;
        RECT 7.2820 47.2635 7.3590 48.3570 ;
        RECT 7.1200 47.2635 7.1460 48.3570 ;
        RECT 7.0120 47.2635 7.0380 48.3570 ;
        RECT 6.9040 47.2635 6.9300 48.3570 ;
        RECT 6.7960 47.2635 6.8220 48.3570 ;
        RECT 6.6880 47.2635 6.7140 48.3570 ;
        RECT 6.5800 47.2635 6.6060 48.3570 ;
        RECT 6.4720 47.2635 6.4980 48.3570 ;
        RECT 6.3640 47.2635 6.3900 48.3570 ;
        RECT 6.2560 47.2635 6.2820 48.3570 ;
        RECT 6.1480 47.2635 6.1740 48.3570 ;
        RECT 6.0400 47.2635 6.0660 48.3570 ;
        RECT 5.9320 47.2635 5.9580 48.3570 ;
        RECT 5.8240 47.2635 5.8500 48.3570 ;
        RECT 5.7160 47.2635 5.7420 48.3570 ;
        RECT 5.6080 47.2635 5.6340 48.3570 ;
        RECT 5.5000 47.2635 5.5260 48.3570 ;
        RECT 5.3920 47.2635 5.4180 48.3570 ;
        RECT 5.2840 47.2635 5.3100 48.3570 ;
        RECT 5.1760 47.2635 5.2020 48.3570 ;
        RECT 5.0680 47.2635 5.0940 48.3570 ;
        RECT 4.9600 47.2635 4.9860 48.3570 ;
        RECT 4.8520 47.2635 4.8780 48.3570 ;
        RECT 4.7440 47.2635 4.7700 48.3570 ;
        RECT 4.6360 47.2635 4.6620 48.3570 ;
        RECT 4.5280 47.2635 4.5540 48.3570 ;
        RECT 4.4200 47.2635 4.4460 48.3570 ;
        RECT 4.3120 47.2635 4.3380 48.3570 ;
        RECT 4.2040 47.2635 4.2300 48.3570 ;
        RECT 4.0960 47.2635 4.1220 48.3570 ;
        RECT 3.9880 47.2635 4.0140 48.3570 ;
        RECT 3.8800 47.2635 3.9060 48.3570 ;
        RECT 3.7720 47.2635 3.7980 48.3570 ;
        RECT 3.6640 47.2635 3.6900 48.3570 ;
        RECT 3.5560 47.2635 3.5820 48.3570 ;
        RECT 3.4480 47.2635 3.4740 48.3570 ;
        RECT 3.3400 47.2635 3.3660 48.3570 ;
        RECT 3.2320 47.2635 3.2580 48.3570 ;
        RECT 3.1240 47.2635 3.1500 48.3570 ;
        RECT 3.0160 47.2635 3.0420 48.3570 ;
        RECT 2.9080 47.2635 2.9340 48.3570 ;
        RECT 2.8000 47.2635 2.8260 48.3570 ;
        RECT 2.6920 47.2635 2.7180 48.3570 ;
        RECT 2.5840 47.2635 2.6100 48.3570 ;
        RECT 2.4760 47.2635 2.5020 48.3570 ;
        RECT 2.3680 47.2635 2.3940 48.3570 ;
        RECT 2.2600 47.2635 2.2860 48.3570 ;
        RECT 2.1520 47.2635 2.1780 48.3570 ;
        RECT 2.0440 47.2635 2.0700 48.3570 ;
        RECT 1.9360 47.2635 1.9620 48.3570 ;
        RECT 1.8280 47.2635 1.8540 48.3570 ;
        RECT 1.7200 47.2635 1.7460 48.3570 ;
        RECT 1.6120 47.2635 1.6380 48.3570 ;
        RECT 1.5040 47.2635 1.5300 48.3570 ;
        RECT 1.3960 47.2635 1.4220 48.3570 ;
        RECT 1.2880 47.2635 1.3140 48.3570 ;
        RECT 1.1800 47.2635 1.2060 48.3570 ;
        RECT 1.0720 47.2635 1.0980 48.3570 ;
        RECT 0.9640 47.2635 0.9900 48.3570 ;
        RECT 0.8560 47.2635 0.8820 48.3570 ;
        RECT 0.7480 47.2635 0.7740 48.3570 ;
        RECT 0.6400 47.2635 0.6660 48.3570 ;
        RECT 0.5320 47.2635 0.5580 48.3570 ;
        RECT 0.4240 47.2635 0.4500 48.3570 ;
        RECT 0.3160 47.2635 0.3420 48.3570 ;
        RECT 0.2080 47.2635 0.2340 48.3570 ;
        RECT 0.0050 47.2635 0.0900 48.3570 ;
        RECT 8.6410 48.3435 8.7690 49.4370 ;
        RECT 8.6270 49.0090 8.7690 49.3315 ;
        RECT 8.4790 48.7360 8.5410 49.4370 ;
        RECT 8.4650 49.0455 8.5410 49.1990 ;
        RECT 8.4790 48.3435 8.5050 49.4370 ;
        RECT 8.4790 48.4645 8.5190 48.7040 ;
        RECT 8.4790 48.3435 8.5410 48.4325 ;
        RECT 8.1820 48.7940 8.3880 49.4370 ;
        RECT 8.3620 48.3435 8.3880 49.4370 ;
        RECT 8.1820 49.0710 8.4020 49.3290 ;
        RECT 8.1820 48.3435 8.2800 49.4370 ;
        RECT 7.7650 48.3435 7.8480 49.4370 ;
        RECT 7.7650 48.4320 7.8620 49.3675 ;
        RECT 16.4440 48.3435 16.5290 49.4370 ;
        RECT 16.3000 48.3435 16.3260 49.4370 ;
        RECT 16.1920 48.3435 16.2180 49.4370 ;
        RECT 16.0840 48.3435 16.1100 49.4370 ;
        RECT 15.9760 48.3435 16.0020 49.4370 ;
        RECT 15.8680 48.3435 15.8940 49.4370 ;
        RECT 15.7600 48.3435 15.7860 49.4370 ;
        RECT 15.6520 48.3435 15.6780 49.4370 ;
        RECT 15.5440 48.3435 15.5700 49.4370 ;
        RECT 15.4360 48.3435 15.4620 49.4370 ;
        RECT 15.3280 48.3435 15.3540 49.4370 ;
        RECT 15.2200 48.3435 15.2460 49.4370 ;
        RECT 15.1120 48.3435 15.1380 49.4370 ;
        RECT 15.0040 48.3435 15.0300 49.4370 ;
        RECT 14.8960 48.3435 14.9220 49.4370 ;
        RECT 14.7880 48.3435 14.8140 49.4370 ;
        RECT 14.6800 48.3435 14.7060 49.4370 ;
        RECT 14.5720 48.3435 14.5980 49.4370 ;
        RECT 14.4640 48.3435 14.4900 49.4370 ;
        RECT 14.3560 48.3435 14.3820 49.4370 ;
        RECT 14.2480 48.3435 14.2740 49.4370 ;
        RECT 14.1400 48.3435 14.1660 49.4370 ;
        RECT 14.0320 48.3435 14.0580 49.4370 ;
        RECT 13.9240 48.3435 13.9500 49.4370 ;
        RECT 13.8160 48.3435 13.8420 49.4370 ;
        RECT 13.7080 48.3435 13.7340 49.4370 ;
        RECT 13.6000 48.3435 13.6260 49.4370 ;
        RECT 13.4920 48.3435 13.5180 49.4370 ;
        RECT 13.3840 48.3435 13.4100 49.4370 ;
        RECT 13.2760 48.3435 13.3020 49.4370 ;
        RECT 13.1680 48.3435 13.1940 49.4370 ;
        RECT 13.0600 48.3435 13.0860 49.4370 ;
        RECT 12.9520 48.3435 12.9780 49.4370 ;
        RECT 12.8440 48.3435 12.8700 49.4370 ;
        RECT 12.7360 48.3435 12.7620 49.4370 ;
        RECT 12.6280 48.3435 12.6540 49.4370 ;
        RECT 12.5200 48.3435 12.5460 49.4370 ;
        RECT 12.4120 48.3435 12.4380 49.4370 ;
        RECT 12.3040 48.3435 12.3300 49.4370 ;
        RECT 12.1960 48.3435 12.2220 49.4370 ;
        RECT 12.0880 48.3435 12.1140 49.4370 ;
        RECT 11.9800 48.3435 12.0060 49.4370 ;
        RECT 11.8720 48.3435 11.8980 49.4370 ;
        RECT 11.7640 48.3435 11.7900 49.4370 ;
        RECT 11.6560 48.3435 11.6820 49.4370 ;
        RECT 11.5480 48.3435 11.5740 49.4370 ;
        RECT 11.4400 48.3435 11.4660 49.4370 ;
        RECT 11.3320 48.3435 11.3580 49.4370 ;
        RECT 11.2240 48.3435 11.2500 49.4370 ;
        RECT 11.1160 48.3435 11.1420 49.4370 ;
        RECT 11.0080 48.3435 11.0340 49.4370 ;
        RECT 10.9000 48.3435 10.9260 49.4370 ;
        RECT 10.7920 48.3435 10.8180 49.4370 ;
        RECT 10.6840 48.3435 10.7100 49.4370 ;
        RECT 10.5760 48.3435 10.6020 49.4370 ;
        RECT 10.4680 48.3435 10.4940 49.4370 ;
        RECT 10.3600 48.3435 10.3860 49.4370 ;
        RECT 10.2520 48.3435 10.2780 49.4370 ;
        RECT 10.1440 48.3435 10.1700 49.4370 ;
        RECT 10.0360 48.3435 10.0620 49.4370 ;
        RECT 9.9280 48.3435 9.9540 49.4370 ;
        RECT 9.8200 48.3435 9.8460 49.4370 ;
        RECT 9.7120 48.3435 9.7380 49.4370 ;
        RECT 9.6040 48.3435 9.6300 49.4370 ;
        RECT 9.4960 48.3435 9.5220 49.4370 ;
        RECT 9.3880 48.3435 9.4140 49.4370 ;
        RECT 9.1750 48.3435 9.2520 49.4370 ;
        RECT 7.2820 48.3435 7.3590 49.4370 ;
        RECT 7.1200 48.3435 7.1460 49.4370 ;
        RECT 7.0120 48.3435 7.0380 49.4370 ;
        RECT 6.9040 48.3435 6.9300 49.4370 ;
        RECT 6.7960 48.3435 6.8220 49.4370 ;
        RECT 6.6880 48.3435 6.7140 49.4370 ;
        RECT 6.5800 48.3435 6.6060 49.4370 ;
        RECT 6.4720 48.3435 6.4980 49.4370 ;
        RECT 6.3640 48.3435 6.3900 49.4370 ;
        RECT 6.2560 48.3435 6.2820 49.4370 ;
        RECT 6.1480 48.3435 6.1740 49.4370 ;
        RECT 6.0400 48.3435 6.0660 49.4370 ;
        RECT 5.9320 48.3435 5.9580 49.4370 ;
        RECT 5.8240 48.3435 5.8500 49.4370 ;
        RECT 5.7160 48.3435 5.7420 49.4370 ;
        RECT 5.6080 48.3435 5.6340 49.4370 ;
        RECT 5.5000 48.3435 5.5260 49.4370 ;
        RECT 5.3920 48.3435 5.4180 49.4370 ;
        RECT 5.2840 48.3435 5.3100 49.4370 ;
        RECT 5.1760 48.3435 5.2020 49.4370 ;
        RECT 5.0680 48.3435 5.0940 49.4370 ;
        RECT 4.9600 48.3435 4.9860 49.4370 ;
        RECT 4.8520 48.3435 4.8780 49.4370 ;
        RECT 4.7440 48.3435 4.7700 49.4370 ;
        RECT 4.6360 48.3435 4.6620 49.4370 ;
        RECT 4.5280 48.3435 4.5540 49.4370 ;
        RECT 4.4200 48.3435 4.4460 49.4370 ;
        RECT 4.3120 48.3435 4.3380 49.4370 ;
        RECT 4.2040 48.3435 4.2300 49.4370 ;
        RECT 4.0960 48.3435 4.1220 49.4370 ;
        RECT 3.9880 48.3435 4.0140 49.4370 ;
        RECT 3.8800 48.3435 3.9060 49.4370 ;
        RECT 3.7720 48.3435 3.7980 49.4370 ;
        RECT 3.6640 48.3435 3.6900 49.4370 ;
        RECT 3.5560 48.3435 3.5820 49.4370 ;
        RECT 3.4480 48.3435 3.4740 49.4370 ;
        RECT 3.3400 48.3435 3.3660 49.4370 ;
        RECT 3.2320 48.3435 3.2580 49.4370 ;
        RECT 3.1240 48.3435 3.1500 49.4370 ;
        RECT 3.0160 48.3435 3.0420 49.4370 ;
        RECT 2.9080 48.3435 2.9340 49.4370 ;
        RECT 2.8000 48.3435 2.8260 49.4370 ;
        RECT 2.6920 48.3435 2.7180 49.4370 ;
        RECT 2.5840 48.3435 2.6100 49.4370 ;
        RECT 2.4760 48.3435 2.5020 49.4370 ;
        RECT 2.3680 48.3435 2.3940 49.4370 ;
        RECT 2.2600 48.3435 2.2860 49.4370 ;
        RECT 2.1520 48.3435 2.1780 49.4370 ;
        RECT 2.0440 48.3435 2.0700 49.4370 ;
        RECT 1.9360 48.3435 1.9620 49.4370 ;
        RECT 1.8280 48.3435 1.8540 49.4370 ;
        RECT 1.7200 48.3435 1.7460 49.4370 ;
        RECT 1.6120 48.3435 1.6380 49.4370 ;
        RECT 1.5040 48.3435 1.5300 49.4370 ;
        RECT 1.3960 48.3435 1.4220 49.4370 ;
        RECT 1.2880 48.3435 1.3140 49.4370 ;
        RECT 1.1800 48.3435 1.2060 49.4370 ;
        RECT 1.0720 48.3435 1.0980 49.4370 ;
        RECT 0.9640 48.3435 0.9900 49.4370 ;
        RECT 0.8560 48.3435 0.8820 49.4370 ;
        RECT 0.7480 48.3435 0.7740 49.4370 ;
        RECT 0.6400 48.3435 0.6660 49.4370 ;
        RECT 0.5320 48.3435 0.5580 49.4370 ;
        RECT 0.4240 48.3435 0.4500 49.4370 ;
        RECT 0.3160 48.3435 0.3420 49.4370 ;
        RECT 0.2080 48.3435 0.2340 49.4370 ;
        RECT 0.0050 48.3435 0.0900 49.4370 ;
        RECT 8.6410 49.4235 8.7690 50.5170 ;
        RECT 8.6270 50.0890 8.7690 50.4115 ;
        RECT 8.4790 49.8160 8.5410 50.5170 ;
        RECT 8.4650 50.1255 8.5410 50.2790 ;
        RECT 8.4790 49.4235 8.5050 50.5170 ;
        RECT 8.4790 49.5445 8.5190 49.7840 ;
        RECT 8.4790 49.4235 8.5410 49.5125 ;
        RECT 8.1820 49.8740 8.3880 50.5170 ;
        RECT 8.3620 49.4235 8.3880 50.5170 ;
        RECT 8.1820 50.1510 8.4020 50.4090 ;
        RECT 8.1820 49.4235 8.2800 50.5170 ;
        RECT 7.7650 49.4235 7.8480 50.5170 ;
        RECT 7.7650 49.5120 7.8620 50.4475 ;
        RECT 16.4440 49.4235 16.5290 50.5170 ;
        RECT 16.3000 49.4235 16.3260 50.5170 ;
        RECT 16.1920 49.4235 16.2180 50.5170 ;
        RECT 16.0840 49.4235 16.1100 50.5170 ;
        RECT 15.9760 49.4235 16.0020 50.5170 ;
        RECT 15.8680 49.4235 15.8940 50.5170 ;
        RECT 15.7600 49.4235 15.7860 50.5170 ;
        RECT 15.6520 49.4235 15.6780 50.5170 ;
        RECT 15.5440 49.4235 15.5700 50.5170 ;
        RECT 15.4360 49.4235 15.4620 50.5170 ;
        RECT 15.3280 49.4235 15.3540 50.5170 ;
        RECT 15.2200 49.4235 15.2460 50.5170 ;
        RECT 15.1120 49.4235 15.1380 50.5170 ;
        RECT 15.0040 49.4235 15.0300 50.5170 ;
        RECT 14.8960 49.4235 14.9220 50.5170 ;
        RECT 14.7880 49.4235 14.8140 50.5170 ;
        RECT 14.6800 49.4235 14.7060 50.5170 ;
        RECT 14.5720 49.4235 14.5980 50.5170 ;
        RECT 14.4640 49.4235 14.4900 50.5170 ;
        RECT 14.3560 49.4235 14.3820 50.5170 ;
        RECT 14.2480 49.4235 14.2740 50.5170 ;
        RECT 14.1400 49.4235 14.1660 50.5170 ;
        RECT 14.0320 49.4235 14.0580 50.5170 ;
        RECT 13.9240 49.4235 13.9500 50.5170 ;
        RECT 13.8160 49.4235 13.8420 50.5170 ;
        RECT 13.7080 49.4235 13.7340 50.5170 ;
        RECT 13.6000 49.4235 13.6260 50.5170 ;
        RECT 13.4920 49.4235 13.5180 50.5170 ;
        RECT 13.3840 49.4235 13.4100 50.5170 ;
        RECT 13.2760 49.4235 13.3020 50.5170 ;
        RECT 13.1680 49.4235 13.1940 50.5170 ;
        RECT 13.0600 49.4235 13.0860 50.5170 ;
        RECT 12.9520 49.4235 12.9780 50.5170 ;
        RECT 12.8440 49.4235 12.8700 50.5170 ;
        RECT 12.7360 49.4235 12.7620 50.5170 ;
        RECT 12.6280 49.4235 12.6540 50.5170 ;
        RECT 12.5200 49.4235 12.5460 50.5170 ;
        RECT 12.4120 49.4235 12.4380 50.5170 ;
        RECT 12.3040 49.4235 12.3300 50.5170 ;
        RECT 12.1960 49.4235 12.2220 50.5170 ;
        RECT 12.0880 49.4235 12.1140 50.5170 ;
        RECT 11.9800 49.4235 12.0060 50.5170 ;
        RECT 11.8720 49.4235 11.8980 50.5170 ;
        RECT 11.7640 49.4235 11.7900 50.5170 ;
        RECT 11.6560 49.4235 11.6820 50.5170 ;
        RECT 11.5480 49.4235 11.5740 50.5170 ;
        RECT 11.4400 49.4235 11.4660 50.5170 ;
        RECT 11.3320 49.4235 11.3580 50.5170 ;
        RECT 11.2240 49.4235 11.2500 50.5170 ;
        RECT 11.1160 49.4235 11.1420 50.5170 ;
        RECT 11.0080 49.4235 11.0340 50.5170 ;
        RECT 10.9000 49.4235 10.9260 50.5170 ;
        RECT 10.7920 49.4235 10.8180 50.5170 ;
        RECT 10.6840 49.4235 10.7100 50.5170 ;
        RECT 10.5760 49.4235 10.6020 50.5170 ;
        RECT 10.4680 49.4235 10.4940 50.5170 ;
        RECT 10.3600 49.4235 10.3860 50.5170 ;
        RECT 10.2520 49.4235 10.2780 50.5170 ;
        RECT 10.1440 49.4235 10.1700 50.5170 ;
        RECT 10.0360 49.4235 10.0620 50.5170 ;
        RECT 9.9280 49.4235 9.9540 50.5170 ;
        RECT 9.8200 49.4235 9.8460 50.5170 ;
        RECT 9.7120 49.4235 9.7380 50.5170 ;
        RECT 9.6040 49.4235 9.6300 50.5170 ;
        RECT 9.4960 49.4235 9.5220 50.5170 ;
        RECT 9.3880 49.4235 9.4140 50.5170 ;
        RECT 9.1750 49.4235 9.2520 50.5170 ;
        RECT 7.2820 49.4235 7.3590 50.5170 ;
        RECT 7.1200 49.4235 7.1460 50.5170 ;
        RECT 7.0120 49.4235 7.0380 50.5170 ;
        RECT 6.9040 49.4235 6.9300 50.5170 ;
        RECT 6.7960 49.4235 6.8220 50.5170 ;
        RECT 6.6880 49.4235 6.7140 50.5170 ;
        RECT 6.5800 49.4235 6.6060 50.5170 ;
        RECT 6.4720 49.4235 6.4980 50.5170 ;
        RECT 6.3640 49.4235 6.3900 50.5170 ;
        RECT 6.2560 49.4235 6.2820 50.5170 ;
        RECT 6.1480 49.4235 6.1740 50.5170 ;
        RECT 6.0400 49.4235 6.0660 50.5170 ;
        RECT 5.9320 49.4235 5.9580 50.5170 ;
        RECT 5.8240 49.4235 5.8500 50.5170 ;
        RECT 5.7160 49.4235 5.7420 50.5170 ;
        RECT 5.6080 49.4235 5.6340 50.5170 ;
        RECT 5.5000 49.4235 5.5260 50.5170 ;
        RECT 5.3920 49.4235 5.4180 50.5170 ;
        RECT 5.2840 49.4235 5.3100 50.5170 ;
        RECT 5.1760 49.4235 5.2020 50.5170 ;
        RECT 5.0680 49.4235 5.0940 50.5170 ;
        RECT 4.9600 49.4235 4.9860 50.5170 ;
        RECT 4.8520 49.4235 4.8780 50.5170 ;
        RECT 4.7440 49.4235 4.7700 50.5170 ;
        RECT 4.6360 49.4235 4.6620 50.5170 ;
        RECT 4.5280 49.4235 4.5540 50.5170 ;
        RECT 4.4200 49.4235 4.4460 50.5170 ;
        RECT 4.3120 49.4235 4.3380 50.5170 ;
        RECT 4.2040 49.4235 4.2300 50.5170 ;
        RECT 4.0960 49.4235 4.1220 50.5170 ;
        RECT 3.9880 49.4235 4.0140 50.5170 ;
        RECT 3.8800 49.4235 3.9060 50.5170 ;
        RECT 3.7720 49.4235 3.7980 50.5170 ;
        RECT 3.6640 49.4235 3.6900 50.5170 ;
        RECT 3.5560 49.4235 3.5820 50.5170 ;
        RECT 3.4480 49.4235 3.4740 50.5170 ;
        RECT 3.3400 49.4235 3.3660 50.5170 ;
        RECT 3.2320 49.4235 3.2580 50.5170 ;
        RECT 3.1240 49.4235 3.1500 50.5170 ;
        RECT 3.0160 49.4235 3.0420 50.5170 ;
        RECT 2.9080 49.4235 2.9340 50.5170 ;
        RECT 2.8000 49.4235 2.8260 50.5170 ;
        RECT 2.6920 49.4235 2.7180 50.5170 ;
        RECT 2.5840 49.4235 2.6100 50.5170 ;
        RECT 2.4760 49.4235 2.5020 50.5170 ;
        RECT 2.3680 49.4235 2.3940 50.5170 ;
        RECT 2.2600 49.4235 2.2860 50.5170 ;
        RECT 2.1520 49.4235 2.1780 50.5170 ;
        RECT 2.0440 49.4235 2.0700 50.5170 ;
        RECT 1.9360 49.4235 1.9620 50.5170 ;
        RECT 1.8280 49.4235 1.8540 50.5170 ;
        RECT 1.7200 49.4235 1.7460 50.5170 ;
        RECT 1.6120 49.4235 1.6380 50.5170 ;
        RECT 1.5040 49.4235 1.5300 50.5170 ;
        RECT 1.3960 49.4235 1.4220 50.5170 ;
        RECT 1.2880 49.4235 1.3140 50.5170 ;
        RECT 1.1800 49.4235 1.2060 50.5170 ;
        RECT 1.0720 49.4235 1.0980 50.5170 ;
        RECT 0.9640 49.4235 0.9900 50.5170 ;
        RECT 0.8560 49.4235 0.8820 50.5170 ;
        RECT 0.7480 49.4235 0.7740 50.5170 ;
        RECT 0.6400 49.4235 0.6660 50.5170 ;
        RECT 0.5320 49.4235 0.5580 50.5170 ;
        RECT 0.4240 49.4235 0.4500 50.5170 ;
        RECT 0.3160 49.4235 0.3420 50.5170 ;
        RECT 0.2080 49.4235 0.2340 50.5170 ;
        RECT 0.0050 49.4235 0.0900 50.5170 ;
        RECT 8.6410 50.5035 8.7690 51.5970 ;
        RECT 8.6270 51.1690 8.7690 51.4915 ;
        RECT 8.4790 50.8960 8.5410 51.5970 ;
        RECT 8.4650 51.2055 8.5410 51.3590 ;
        RECT 8.4790 50.5035 8.5050 51.5970 ;
        RECT 8.4790 50.6245 8.5190 50.8640 ;
        RECT 8.4790 50.5035 8.5410 50.5925 ;
        RECT 8.1820 50.9540 8.3880 51.5970 ;
        RECT 8.3620 50.5035 8.3880 51.5970 ;
        RECT 8.1820 51.2310 8.4020 51.4890 ;
        RECT 8.1820 50.5035 8.2800 51.5970 ;
        RECT 7.7650 50.5035 7.8480 51.5970 ;
        RECT 7.7650 50.5920 7.8620 51.5275 ;
        RECT 16.4440 50.5035 16.5290 51.5970 ;
        RECT 16.3000 50.5035 16.3260 51.5970 ;
        RECT 16.1920 50.5035 16.2180 51.5970 ;
        RECT 16.0840 50.5035 16.1100 51.5970 ;
        RECT 15.9760 50.5035 16.0020 51.5970 ;
        RECT 15.8680 50.5035 15.8940 51.5970 ;
        RECT 15.7600 50.5035 15.7860 51.5970 ;
        RECT 15.6520 50.5035 15.6780 51.5970 ;
        RECT 15.5440 50.5035 15.5700 51.5970 ;
        RECT 15.4360 50.5035 15.4620 51.5970 ;
        RECT 15.3280 50.5035 15.3540 51.5970 ;
        RECT 15.2200 50.5035 15.2460 51.5970 ;
        RECT 15.1120 50.5035 15.1380 51.5970 ;
        RECT 15.0040 50.5035 15.0300 51.5970 ;
        RECT 14.8960 50.5035 14.9220 51.5970 ;
        RECT 14.7880 50.5035 14.8140 51.5970 ;
        RECT 14.6800 50.5035 14.7060 51.5970 ;
        RECT 14.5720 50.5035 14.5980 51.5970 ;
        RECT 14.4640 50.5035 14.4900 51.5970 ;
        RECT 14.3560 50.5035 14.3820 51.5970 ;
        RECT 14.2480 50.5035 14.2740 51.5970 ;
        RECT 14.1400 50.5035 14.1660 51.5970 ;
        RECT 14.0320 50.5035 14.0580 51.5970 ;
        RECT 13.9240 50.5035 13.9500 51.5970 ;
        RECT 13.8160 50.5035 13.8420 51.5970 ;
        RECT 13.7080 50.5035 13.7340 51.5970 ;
        RECT 13.6000 50.5035 13.6260 51.5970 ;
        RECT 13.4920 50.5035 13.5180 51.5970 ;
        RECT 13.3840 50.5035 13.4100 51.5970 ;
        RECT 13.2760 50.5035 13.3020 51.5970 ;
        RECT 13.1680 50.5035 13.1940 51.5970 ;
        RECT 13.0600 50.5035 13.0860 51.5970 ;
        RECT 12.9520 50.5035 12.9780 51.5970 ;
        RECT 12.8440 50.5035 12.8700 51.5970 ;
        RECT 12.7360 50.5035 12.7620 51.5970 ;
        RECT 12.6280 50.5035 12.6540 51.5970 ;
        RECT 12.5200 50.5035 12.5460 51.5970 ;
        RECT 12.4120 50.5035 12.4380 51.5970 ;
        RECT 12.3040 50.5035 12.3300 51.5970 ;
        RECT 12.1960 50.5035 12.2220 51.5970 ;
        RECT 12.0880 50.5035 12.1140 51.5970 ;
        RECT 11.9800 50.5035 12.0060 51.5970 ;
        RECT 11.8720 50.5035 11.8980 51.5970 ;
        RECT 11.7640 50.5035 11.7900 51.5970 ;
        RECT 11.6560 50.5035 11.6820 51.5970 ;
        RECT 11.5480 50.5035 11.5740 51.5970 ;
        RECT 11.4400 50.5035 11.4660 51.5970 ;
        RECT 11.3320 50.5035 11.3580 51.5970 ;
        RECT 11.2240 50.5035 11.2500 51.5970 ;
        RECT 11.1160 50.5035 11.1420 51.5970 ;
        RECT 11.0080 50.5035 11.0340 51.5970 ;
        RECT 10.9000 50.5035 10.9260 51.5970 ;
        RECT 10.7920 50.5035 10.8180 51.5970 ;
        RECT 10.6840 50.5035 10.7100 51.5970 ;
        RECT 10.5760 50.5035 10.6020 51.5970 ;
        RECT 10.4680 50.5035 10.4940 51.5970 ;
        RECT 10.3600 50.5035 10.3860 51.5970 ;
        RECT 10.2520 50.5035 10.2780 51.5970 ;
        RECT 10.1440 50.5035 10.1700 51.5970 ;
        RECT 10.0360 50.5035 10.0620 51.5970 ;
        RECT 9.9280 50.5035 9.9540 51.5970 ;
        RECT 9.8200 50.5035 9.8460 51.5970 ;
        RECT 9.7120 50.5035 9.7380 51.5970 ;
        RECT 9.6040 50.5035 9.6300 51.5970 ;
        RECT 9.4960 50.5035 9.5220 51.5970 ;
        RECT 9.3880 50.5035 9.4140 51.5970 ;
        RECT 9.1750 50.5035 9.2520 51.5970 ;
        RECT 7.2820 50.5035 7.3590 51.5970 ;
        RECT 7.1200 50.5035 7.1460 51.5970 ;
        RECT 7.0120 50.5035 7.0380 51.5970 ;
        RECT 6.9040 50.5035 6.9300 51.5970 ;
        RECT 6.7960 50.5035 6.8220 51.5970 ;
        RECT 6.6880 50.5035 6.7140 51.5970 ;
        RECT 6.5800 50.5035 6.6060 51.5970 ;
        RECT 6.4720 50.5035 6.4980 51.5970 ;
        RECT 6.3640 50.5035 6.3900 51.5970 ;
        RECT 6.2560 50.5035 6.2820 51.5970 ;
        RECT 6.1480 50.5035 6.1740 51.5970 ;
        RECT 6.0400 50.5035 6.0660 51.5970 ;
        RECT 5.9320 50.5035 5.9580 51.5970 ;
        RECT 5.8240 50.5035 5.8500 51.5970 ;
        RECT 5.7160 50.5035 5.7420 51.5970 ;
        RECT 5.6080 50.5035 5.6340 51.5970 ;
        RECT 5.5000 50.5035 5.5260 51.5970 ;
        RECT 5.3920 50.5035 5.4180 51.5970 ;
        RECT 5.2840 50.5035 5.3100 51.5970 ;
        RECT 5.1760 50.5035 5.2020 51.5970 ;
        RECT 5.0680 50.5035 5.0940 51.5970 ;
        RECT 4.9600 50.5035 4.9860 51.5970 ;
        RECT 4.8520 50.5035 4.8780 51.5970 ;
        RECT 4.7440 50.5035 4.7700 51.5970 ;
        RECT 4.6360 50.5035 4.6620 51.5970 ;
        RECT 4.5280 50.5035 4.5540 51.5970 ;
        RECT 4.4200 50.5035 4.4460 51.5970 ;
        RECT 4.3120 50.5035 4.3380 51.5970 ;
        RECT 4.2040 50.5035 4.2300 51.5970 ;
        RECT 4.0960 50.5035 4.1220 51.5970 ;
        RECT 3.9880 50.5035 4.0140 51.5970 ;
        RECT 3.8800 50.5035 3.9060 51.5970 ;
        RECT 3.7720 50.5035 3.7980 51.5970 ;
        RECT 3.6640 50.5035 3.6900 51.5970 ;
        RECT 3.5560 50.5035 3.5820 51.5970 ;
        RECT 3.4480 50.5035 3.4740 51.5970 ;
        RECT 3.3400 50.5035 3.3660 51.5970 ;
        RECT 3.2320 50.5035 3.2580 51.5970 ;
        RECT 3.1240 50.5035 3.1500 51.5970 ;
        RECT 3.0160 50.5035 3.0420 51.5970 ;
        RECT 2.9080 50.5035 2.9340 51.5970 ;
        RECT 2.8000 50.5035 2.8260 51.5970 ;
        RECT 2.6920 50.5035 2.7180 51.5970 ;
        RECT 2.5840 50.5035 2.6100 51.5970 ;
        RECT 2.4760 50.5035 2.5020 51.5970 ;
        RECT 2.3680 50.5035 2.3940 51.5970 ;
        RECT 2.2600 50.5035 2.2860 51.5970 ;
        RECT 2.1520 50.5035 2.1780 51.5970 ;
        RECT 2.0440 50.5035 2.0700 51.5970 ;
        RECT 1.9360 50.5035 1.9620 51.5970 ;
        RECT 1.8280 50.5035 1.8540 51.5970 ;
        RECT 1.7200 50.5035 1.7460 51.5970 ;
        RECT 1.6120 50.5035 1.6380 51.5970 ;
        RECT 1.5040 50.5035 1.5300 51.5970 ;
        RECT 1.3960 50.5035 1.4220 51.5970 ;
        RECT 1.2880 50.5035 1.3140 51.5970 ;
        RECT 1.1800 50.5035 1.2060 51.5970 ;
        RECT 1.0720 50.5035 1.0980 51.5970 ;
        RECT 0.9640 50.5035 0.9900 51.5970 ;
        RECT 0.8560 50.5035 0.8820 51.5970 ;
        RECT 0.7480 50.5035 0.7740 51.5970 ;
        RECT 0.6400 50.5035 0.6660 51.5970 ;
        RECT 0.5320 50.5035 0.5580 51.5970 ;
        RECT 0.4240 50.5035 0.4500 51.5970 ;
        RECT 0.3160 50.5035 0.3420 51.5970 ;
        RECT 0.2080 50.5035 0.2340 51.5970 ;
        RECT 0.0050 50.5035 0.0900 51.5970 ;
        RECT 8.6410 51.5835 8.7690 52.6770 ;
        RECT 8.6270 52.2490 8.7690 52.5715 ;
        RECT 8.4790 51.9760 8.5410 52.6770 ;
        RECT 8.4650 52.2855 8.5410 52.4390 ;
        RECT 8.4790 51.5835 8.5050 52.6770 ;
        RECT 8.4790 51.7045 8.5190 51.9440 ;
        RECT 8.4790 51.5835 8.5410 51.6725 ;
        RECT 8.1820 52.0340 8.3880 52.6770 ;
        RECT 8.3620 51.5835 8.3880 52.6770 ;
        RECT 8.1820 52.3110 8.4020 52.5690 ;
        RECT 8.1820 51.5835 8.2800 52.6770 ;
        RECT 7.7650 51.5835 7.8480 52.6770 ;
        RECT 7.7650 51.6720 7.8620 52.6075 ;
        RECT 16.4440 51.5835 16.5290 52.6770 ;
        RECT 16.3000 51.5835 16.3260 52.6770 ;
        RECT 16.1920 51.5835 16.2180 52.6770 ;
        RECT 16.0840 51.5835 16.1100 52.6770 ;
        RECT 15.9760 51.5835 16.0020 52.6770 ;
        RECT 15.8680 51.5835 15.8940 52.6770 ;
        RECT 15.7600 51.5835 15.7860 52.6770 ;
        RECT 15.6520 51.5835 15.6780 52.6770 ;
        RECT 15.5440 51.5835 15.5700 52.6770 ;
        RECT 15.4360 51.5835 15.4620 52.6770 ;
        RECT 15.3280 51.5835 15.3540 52.6770 ;
        RECT 15.2200 51.5835 15.2460 52.6770 ;
        RECT 15.1120 51.5835 15.1380 52.6770 ;
        RECT 15.0040 51.5835 15.0300 52.6770 ;
        RECT 14.8960 51.5835 14.9220 52.6770 ;
        RECT 14.7880 51.5835 14.8140 52.6770 ;
        RECT 14.6800 51.5835 14.7060 52.6770 ;
        RECT 14.5720 51.5835 14.5980 52.6770 ;
        RECT 14.4640 51.5835 14.4900 52.6770 ;
        RECT 14.3560 51.5835 14.3820 52.6770 ;
        RECT 14.2480 51.5835 14.2740 52.6770 ;
        RECT 14.1400 51.5835 14.1660 52.6770 ;
        RECT 14.0320 51.5835 14.0580 52.6770 ;
        RECT 13.9240 51.5835 13.9500 52.6770 ;
        RECT 13.8160 51.5835 13.8420 52.6770 ;
        RECT 13.7080 51.5835 13.7340 52.6770 ;
        RECT 13.6000 51.5835 13.6260 52.6770 ;
        RECT 13.4920 51.5835 13.5180 52.6770 ;
        RECT 13.3840 51.5835 13.4100 52.6770 ;
        RECT 13.2760 51.5835 13.3020 52.6770 ;
        RECT 13.1680 51.5835 13.1940 52.6770 ;
        RECT 13.0600 51.5835 13.0860 52.6770 ;
        RECT 12.9520 51.5835 12.9780 52.6770 ;
        RECT 12.8440 51.5835 12.8700 52.6770 ;
        RECT 12.7360 51.5835 12.7620 52.6770 ;
        RECT 12.6280 51.5835 12.6540 52.6770 ;
        RECT 12.5200 51.5835 12.5460 52.6770 ;
        RECT 12.4120 51.5835 12.4380 52.6770 ;
        RECT 12.3040 51.5835 12.3300 52.6770 ;
        RECT 12.1960 51.5835 12.2220 52.6770 ;
        RECT 12.0880 51.5835 12.1140 52.6770 ;
        RECT 11.9800 51.5835 12.0060 52.6770 ;
        RECT 11.8720 51.5835 11.8980 52.6770 ;
        RECT 11.7640 51.5835 11.7900 52.6770 ;
        RECT 11.6560 51.5835 11.6820 52.6770 ;
        RECT 11.5480 51.5835 11.5740 52.6770 ;
        RECT 11.4400 51.5835 11.4660 52.6770 ;
        RECT 11.3320 51.5835 11.3580 52.6770 ;
        RECT 11.2240 51.5835 11.2500 52.6770 ;
        RECT 11.1160 51.5835 11.1420 52.6770 ;
        RECT 11.0080 51.5835 11.0340 52.6770 ;
        RECT 10.9000 51.5835 10.9260 52.6770 ;
        RECT 10.7920 51.5835 10.8180 52.6770 ;
        RECT 10.6840 51.5835 10.7100 52.6770 ;
        RECT 10.5760 51.5835 10.6020 52.6770 ;
        RECT 10.4680 51.5835 10.4940 52.6770 ;
        RECT 10.3600 51.5835 10.3860 52.6770 ;
        RECT 10.2520 51.5835 10.2780 52.6770 ;
        RECT 10.1440 51.5835 10.1700 52.6770 ;
        RECT 10.0360 51.5835 10.0620 52.6770 ;
        RECT 9.9280 51.5835 9.9540 52.6770 ;
        RECT 9.8200 51.5835 9.8460 52.6770 ;
        RECT 9.7120 51.5835 9.7380 52.6770 ;
        RECT 9.6040 51.5835 9.6300 52.6770 ;
        RECT 9.4960 51.5835 9.5220 52.6770 ;
        RECT 9.3880 51.5835 9.4140 52.6770 ;
        RECT 9.1750 51.5835 9.2520 52.6770 ;
        RECT 7.2820 51.5835 7.3590 52.6770 ;
        RECT 7.1200 51.5835 7.1460 52.6770 ;
        RECT 7.0120 51.5835 7.0380 52.6770 ;
        RECT 6.9040 51.5835 6.9300 52.6770 ;
        RECT 6.7960 51.5835 6.8220 52.6770 ;
        RECT 6.6880 51.5835 6.7140 52.6770 ;
        RECT 6.5800 51.5835 6.6060 52.6770 ;
        RECT 6.4720 51.5835 6.4980 52.6770 ;
        RECT 6.3640 51.5835 6.3900 52.6770 ;
        RECT 6.2560 51.5835 6.2820 52.6770 ;
        RECT 6.1480 51.5835 6.1740 52.6770 ;
        RECT 6.0400 51.5835 6.0660 52.6770 ;
        RECT 5.9320 51.5835 5.9580 52.6770 ;
        RECT 5.8240 51.5835 5.8500 52.6770 ;
        RECT 5.7160 51.5835 5.7420 52.6770 ;
        RECT 5.6080 51.5835 5.6340 52.6770 ;
        RECT 5.5000 51.5835 5.5260 52.6770 ;
        RECT 5.3920 51.5835 5.4180 52.6770 ;
        RECT 5.2840 51.5835 5.3100 52.6770 ;
        RECT 5.1760 51.5835 5.2020 52.6770 ;
        RECT 5.0680 51.5835 5.0940 52.6770 ;
        RECT 4.9600 51.5835 4.9860 52.6770 ;
        RECT 4.8520 51.5835 4.8780 52.6770 ;
        RECT 4.7440 51.5835 4.7700 52.6770 ;
        RECT 4.6360 51.5835 4.6620 52.6770 ;
        RECT 4.5280 51.5835 4.5540 52.6770 ;
        RECT 4.4200 51.5835 4.4460 52.6770 ;
        RECT 4.3120 51.5835 4.3380 52.6770 ;
        RECT 4.2040 51.5835 4.2300 52.6770 ;
        RECT 4.0960 51.5835 4.1220 52.6770 ;
        RECT 3.9880 51.5835 4.0140 52.6770 ;
        RECT 3.8800 51.5835 3.9060 52.6770 ;
        RECT 3.7720 51.5835 3.7980 52.6770 ;
        RECT 3.6640 51.5835 3.6900 52.6770 ;
        RECT 3.5560 51.5835 3.5820 52.6770 ;
        RECT 3.4480 51.5835 3.4740 52.6770 ;
        RECT 3.3400 51.5835 3.3660 52.6770 ;
        RECT 3.2320 51.5835 3.2580 52.6770 ;
        RECT 3.1240 51.5835 3.1500 52.6770 ;
        RECT 3.0160 51.5835 3.0420 52.6770 ;
        RECT 2.9080 51.5835 2.9340 52.6770 ;
        RECT 2.8000 51.5835 2.8260 52.6770 ;
        RECT 2.6920 51.5835 2.7180 52.6770 ;
        RECT 2.5840 51.5835 2.6100 52.6770 ;
        RECT 2.4760 51.5835 2.5020 52.6770 ;
        RECT 2.3680 51.5835 2.3940 52.6770 ;
        RECT 2.2600 51.5835 2.2860 52.6770 ;
        RECT 2.1520 51.5835 2.1780 52.6770 ;
        RECT 2.0440 51.5835 2.0700 52.6770 ;
        RECT 1.9360 51.5835 1.9620 52.6770 ;
        RECT 1.8280 51.5835 1.8540 52.6770 ;
        RECT 1.7200 51.5835 1.7460 52.6770 ;
        RECT 1.6120 51.5835 1.6380 52.6770 ;
        RECT 1.5040 51.5835 1.5300 52.6770 ;
        RECT 1.3960 51.5835 1.4220 52.6770 ;
        RECT 1.2880 51.5835 1.3140 52.6770 ;
        RECT 1.1800 51.5835 1.2060 52.6770 ;
        RECT 1.0720 51.5835 1.0980 52.6770 ;
        RECT 0.9640 51.5835 0.9900 52.6770 ;
        RECT 0.8560 51.5835 0.8820 52.6770 ;
        RECT 0.7480 51.5835 0.7740 52.6770 ;
        RECT 0.6400 51.5835 0.6660 52.6770 ;
        RECT 0.5320 51.5835 0.5580 52.6770 ;
        RECT 0.4240 51.5835 0.4500 52.6770 ;
        RECT 0.3160 51.5835 0.3420 52.6770 ;
        RECT 0.2080 51.5835 0.2340 52.6770 ;
        RECT 0.0050 51.5835 0.0900 52.6770 ;
        RECT 8.6410 52.6635 8.7690 53.7570 ;
        RECT 8.6270 53.3290 8.7690 53.6515 ;
        RECT 8.4790 53.0560 8.5410 53.7570 ;
        RECT 8.4650 53.3655 8.5410 53.5190 ;
        RECT 8.4790 52.6635 8.5050 53.7570 ;
        RECT 8.4790 52.7845 8.5190 53.0240 ;
        RECT 8.4790 52.6635 8.5410 52.7525 ;
        RECT 8.1820 53.1140 8.3880 53.7570 ;
        RECT 8.3620 52.6635 8.3880 53.7570 ;
        RECT 8.1820 53.3910 8.4020 53.6490 ;
        RECT 8.1820 52.6635 8.2800 53.7570 ;
        RECT 7.7650 52.6635 7.8480 53.7570 ;
        RECT 7.7650 52.7520 7.8620 53.6875 ;
        RECT 16.4440 52.6635 16.5290 53.7570 ;
        RECT 16.3000 52.6635 16.3260 53.7570 ;
        RECT 16.1920 52.6635 16.2180 53.7570 ;
        RECT 16.0840 52.6635 16.1100 53.7570 ;
        RECT 15.9760 52.6635 16.0020 53.7570 ;
        RECT 15.8680 52.6635 15.8940 53.7570 ;
        RECT 15.7600 52.6635 15.7860 53.7570 ;
        RECT 15.6520 52.6635 15.6780 53.7570 ;
        RECT 15.5440 52.6635 15.5700 53.7570 ;
        RECT 15.4360 52.6635 15.4620 53.7570 ;
        RECT 15.3280 52.6635 15.3540 53.7570 ;
        RECT 15.2200 52.6635 15.2460 53.7570 ;
        RECT 15.1120 52.6635 15.1380 53.7570 ;
        RECT 15.0040 52.6635 15.0300 53.7570 ;
        RECT 14.8960 52.6635 14.9220 53.7570 ;
        RECT 14.7880 52.6635 14.8140 53.7570 ;
        RECT 14.6800 52.6635 14.7060 53.7570 ;
        RECT 14.5720 52.6635 14.5980 53.7570 ;
        RECT 14.4640 52.6635 14.4900 53.7570 ;
        RECT 14.3560 52.6635 14.3820 53.7570 ;
        RECT 14.2480 52.6635 14.2740 53.7570 ;
        RECT 14.1400 52.6635 14.1660 53.7570 ;
        RECT 14.0320 52.6635 14.0580 53.7570 ;
        RECT 13.9240 52.6635 13.9500 53.7570 ;
        RECT 13.8160 52.6635 13.8420 53.7570 ;
        RECT 13.7080 52.6635 13.7340 53.7570 ;
        RECT 13.6000 52.6635 13.6260 53.7570 ;
        RECT 13.4920 52.6635 13.5180 53.7570 ;
        RECT 13.3840 52.6635 13.4100 53.7570 ;
        RECT 13.2760 52.6635 13.3020 53.7570 ;
        RECT 13.1680 52.6635 13.1940 53.7570 ;
        RECT 13.0600 52.6635 13.0860 53.7570 ;
        RECT 12.9520 52.6635 12.9780 53.7570 ;
        RECT 12.8440 52.6635 12.8700 53.7570 ;
        RECT 12.7360 52.6635 12.7620 53.7570 ;
        RECT 12.6280 52.6635 12.6540 53.7570 ;
        RECT 12.5200 52.6635 12.5460 53.7570 ;
        RECT 12.4120 52.6635 12.4380 53.7570 ;
        RECT 12.3040 52.6635 12.3300 53.7570 ;
        RECT 12.1960 52.6635 12.2220 53.7570 ;
        RECT 12.0880 52.6635 12.1140 53.7570 ;
        RECT 11.9800 52.6635 12.0060 53.7570 ;
        RECT 11.8720 52.6635 11.8980 53.7570 ;
        RECT 11.7640 52.6635 11.7900 53.7570 ;
        RECT 11.6560 52.6635 11.6820 53.7570 ;
        RECT 11.5480 52.6635 11.5740 53.7570 ;
        RECT 11.4400 52.6635 11.4660 53.7570 ;
        RECT 11.3320 52.6635 11.3580 53.7570 ;
        RECT 11.2240 52.6635 11.2500 53.7570 ;
        RECT 11.1160 52.6635 11.1420 53.7570 ;
        RECT 11.0080 52.6635 11.0340 53.7570 ;
        RECT 10.9000 52.6635 10.9260 53.7570 ;
        RECT 10.7920 52.6635 10.8180 53.7570 ;
        RECT 10.6840 52.6635 10.7100 53.7570 ;
        RECT 10.5760 52.6635 10.6020 53.7570 ;
        RECT 10.4680 52.6635 10.4940 53.7570 ;
        RECT 10.3600 52.6635 10.3860 53.7570 ;
        RECT 10.2520 52.6635 10.2780 53.7570 ;
        RECT 10.1440 52.6635 10.1700 53.7570 ;
        RECT 10.0360 52.6635 10.0620 53.7570 ;
        RECT 9.9280 52.6635 9.9540 53.7570 ;
        RECT 9.8200 52.6635 9.8460 53.7570 ;
        RECT 9.7120 52.6635 9.7380 53.7570 ;
        RECT 9.6040 52.6635 9.6300 53.7570 ;
        RECT 9.4960 52.6635 9.5220 53.7570 ;
        RECT 9.3880 52.6635 9.4140 53.7570 ;
        RECT 9.1750 52.6635 9.2520 53.7570 ;
        RECT 7.2820 52.6635 7.3590 53.7570 ;
        RECT 7.1200 52.6635 7.1460 53.7570 ;
        RECT 7.0120 52.6635 7.0380 53.7570 ;
        RECT 6.9040 52.6635 6.9300 53.7570 ;
        RECT 6.7960 52.6635 6.8220 53.7570 ;
        RECT 6.6880 52.6635 6.7140 53.7570 ;
        RECT 6.5800 52.6635 6.6060 53.7570 ;
        RECT 6.4720 52.6635 6.4980 53.7570 ;
        RECT 6.3640 52.6635 6.3900 53.7570 ;
        RECT 6.2560 52.6635 6.2820 53.7570 ;
        RECT 6.1480 52.6635 6.1740 53.7570 ;
        RECT 6.0400 52.6635 6.0660 53.7570 ;
        RECT 5.9320 52.6635 5.9580 53.7570 ;
        RECT 5.8240 52.6635 5.8500 53.7570 ;
        RECT 5.7160 52.6635 5.7420 53.7570 ;
        RECT 5.6080 52.6635 5.6340 53.7570 ;
        RECT 5.5000 52.6635 5.5260 53.7570 ;
        RECT 5.3920 52.6635 5.4180 53.7570 ;
        RECT 5.2840 52.6635 5.3100 53.7570 ;
        RECT 5.1760 52.6635 5.2020 53.7570 ;
        RECT 5.0680 52.6635 5.0940 53.7570 ;
        RECT 4.9600 52.6635 4.9860 53.7570 ;
        RECT 4.8520 52.6635 4.8780 53.7570 ;
        RECT 4.7440 52.6635 4.7700 53.7570 ;
        RECT 4.6360 52.6635 4.6620 53.7570 ;
        RECT 4.5280 52.6635 4.5540 53.7570 ;
        RECT 4.4200 52.6635 4.4460 53.7570 ;
        RECT 4.3120 52.6635 4.3380 53.7570 ;
        RECT 4.2040 52.6635 4.2300 53.7570 ;
        RECT 4.0960 52.6635 4.1220 53.7570 ;
        RECT 3.9880 52.6635 4.0140 53.7570 ;
        RECT 3.8800 52.6635 3.9060 53.7570 ;
        RECT 3.7720 52.6635 3.7980 53.7570 ;
        RECT 3.6640 52.6635 3.6900 53.7570 ;
        RECT 3.5560 52.6635 3.5820 53.7570 ;
        RECT 3.4480 52.6635 3.4740 53.7570 ;
        RECT 3.3400 52.6635 3.3660 53.7570 ;
        RECT 3.2320 52.6635 3.2580 53.7570 ;
        RECT 3.1240 52.6635 3.1500 53.7570 ;
        RECT 3.0160 52.6635 3.0420 53.7570 ;
        RECT 2.9080 52.6635 2.9340 53.7570 ;
        RECT 2.8000 52.6635 2.8260 53.7570 ;
        RECT 2.6920 52.6635 2.7180 53.7570 ;
        RECT 2.5840 52.6635 2.6100 53.7570 ;
        RECT 2.4760 52.6635 2.5020 53.7570 ;
        RECT 2.3680 52.6635 2.3940 53.7570 ;
        RECT 2.2600 52.6635 2.2860 53.7570 ;
        RECT 2.1520 52.6635 2.1780 53.7570 ;
        RECT 2.0440 52.6635 2.0700 53.7570 ;
        RECT 1.9360 52.6635 1.9620 53.7570 ;
        RECT 1.8280 52.6635 1.8540 53.7570 ;
        RECT 1.7200 52.6635 1.7460 53.7570 ;
        RECT 1.6120 52.6635 1.6380 53.7570 ;
        RECT 1.5040 52.6635 1.5300 53.7570 ;
        RECT 1.3960 52.6635 1.4220 53.7570 ;
        RECT 1.2880 52.6635 1.3140 53.7570 ;
        RECT 1.1800 52.6635 1.2060 53.7570 ;
        RECT 1.0720 52.6635 1.0980 53.7570 ;
        RECT 0.9640 52.6635 0.9900 53.7570 ;
        RECT 0.8560 52.6635 0.8820 53.7570 ;
        RECT 0.7480 52.6635 0.7740 53.7570 ;
        RECT 0.6400 52.6635 0.6660 53.7570 ;
        RECT 0.5320 52.6635 0.5580 53.7570 ;
        RECT 0.4240 52.6635 0.4500 53.7570 ;
        RECT 0.3160 52.6635 0.3420 53.7570 ;
        RECT 0.2080 52.6635 0.2340 53.7570 ;
        RECT 0.0050 52.6635 0.0900 53.7570 ;
        RECT 8.6410 53.7435 8.7690 54.8370 ;
        RECT 8.6270 54.4090 8.7690 54.7315 ;
        RECT 8.4790 54.1360 8.5410 54.8370 ;
        RECT 8.4650 54.4455 8.5410 54.5990 ;
        RECT 8.4790 53.7435 8.5050 54.8370 ;
        RECT 8.4790 53.8645 8.5190 54.1040 ;
        RECT 8.4790 53.7435 8.5410 53.8325 ;
        RECT 8.1820 54.1940 8.3880 54.8370 ;
        RECT 8.3620 53.7435 8.3880 54.8370 ;
        RECT 8.1820 54.4710 8.4020 54.7290 ;
        RECT 8.1820 53.7435 8.2800 54.8370 ;
        RECT 7.7650 53.7435 7.8480 54.8370 ;
        RECT 7.7650 53.8320 7.8620 54.7675 ;
        RECT 16.4440 53.7435 16.5290 54.8370 ;
        RECT 16.3000 53.7435 16.3260 54.8370 ;
        RECT 16.1920 53.7435 16.2180 54.8370 ;
        RECT 16.0840 53.7435 16.1100 54.8370 ;
        RECT 15.9760 53.7435 16.0020 54.8370 ;
        RECT 15.8680 53.7435 15.8940 54.8370 ;
        RECT 15.7600 53.7435 15.7860 54.8370 ;
        RECT 15.6520 53.7435 15.6780 54.8370 ;
        RECT 15.5440 53.7435 15.5700 54.8370 ;
        RECT 15.4360 53.7435 15.4620 54.8370 ;
        RECT 15.3280 53.7435 15.3540 54.8370 ;
        RECT 15.2200 53.7435 15.2460 54.8370 ;
        RECT 15.1120 53.7435 15.1380 54.8370 ;
        RECT 15.0040 53.7435 15.0300 54.8370 ;
        RECT 14.8960 53.7435 14.9220 54.8370 ;
        RECT 14.7880 53.7435 14.8140 54.8370 ;
        RECT 14.6800 53.7435 14.7060 54.8370 ;
        RECT 14.5720 53.7435 14.5980 54.8370 ;
        RECT 14.4640 53.7435 14.4900 54.8370 ;
        RECT 14.3560 53.7435 14.3820 54.8370 ;
        RECT 14.2480 53.7435 14.2740 54.8370 ;
        RECT 14.1400 53.7435 14.1660 54.8370 ;
        RECT 14.0320 53.7435 14.0580 54.8370 ;
        RECT 13.9240 53.7435 13.9500 54.8370 ;
        RECT 13.8160 53.7435 13.8420 54.8370 ;
        RECT 13.7080 53.7435 13.7340 54.8370 ;
        RECT 13.6000 53.7435 13.6260 54.8370 ;
        RECT 13.4920 53.7435 13.5180 54.8370 ;
        RECT 13.3840 53.7435 13.4100 54.8370 ;
        RECT 13.2760 53.7435 13.3020 54.8370 ;
        RECT 13.1680 53.7435 13.1940 54.8370 ;
        RECT 13.0600 53.7435 13.0860 54.8370 ;
        RECT 12.9520 53.7435 12.9780 54.8370 ;
        RECT 12.8440 53.7435 12.8700 54.8370 ;
        RECT 12.7360 53.7435 12.7620 54.8370 ;
        RECT 12.6280 53.7435 12.6540 54.8370 ;
        RECT 12.5200 53.7435 12.5460 54.8370 ;
        RECT 12.4120 53.7435 12.4380 54.8370 ;
        RECT 12.3040 53.7435 12.3300 54.8370 ;
        RECT 12.1960 53.7435 12.2220 54.8370 ;
        RECT 12.0880 53.7435 12.1140 54.8370 ;
        RECT 11.9800 53.7435 12.0060 54.8370 ;
        RECT 11.8720 53.7435 11.8980 54.8370 ;
        RECT 11.7640 53.7435 11.7900 54.8370 ;
        RECT 11.6560 53.7435 11.6820 54.8370 ;
        RECT 11.5480 53.7435 11.5740 54.8370 ;
        RECT 11.4400 53.7435 11.4660 54.8370 ;
        RECT 11.3320 53.7435 11.3580 54.8370 ;
        RECT 11.2240 53.7435 11.2500 54.8370 ;
        RECT 11.1160 53.7435 11.1420 54.8370 ;
        RECT 11.0080 53.7435 11.0340 54.8370 ;
        RECT 10.9000 53.7435 10.9260 54.8370 ;
        RECT 10.7920 53.7435 10.8180 54.8370 ;
        RECT 10.6840 53.7435 10.7100 54.8370 ;
        RECT 10.5760 53.7435 10.6020 54.8370 ;
        RECT 10.4680 53.7435 10.4940 54.8370 ;
        RECT 10.3600 53.7435 10.3860 54.8370 ;
        RECT 10.2520 53.7435 10.2780 54.8370 ;
        RECT 10.1440 53.7435 10.1700 54.8370 ;
        RECT 10.0360 53.7435 10.0620 54.8370 ;
        RECT 9.9280 53.7435 9.9540 54.8370 ;
        RECT 9.8200 53.7435 9.8460 54.8370 ;
        RECT 9.7120 53.7435 9.7380 54.8370 ;
        RECT 9.6040 53.7435 9.6300 54.8370 ;
        RECT 9.4960 53.7435 9.5220 54.8370 ;
        RECT 9.3880 53.7435 9.4140 54.8370 ;
        RECT 9.1750 53.7435 9.2520 54.8370 ;
        RECT 7.2820 53.7435 7.3590 54.8370 ;
        RECT 7.1200 53.7435 7.1460 54.8370 ;
        RECT 7.0120 53.7435 7.0380 54.8370 ;
        RECT 6.9040 53.7435 6.9300 54.8370 ;
        RECT 6.7960 53.7435 6.8220 54.8370 ;
        RECT 6.6880 53.7435 6.7140 54.8370 ;
        RECT 6.5800 53.7435 6.6060 54.8370 ;
        RECT 6.4720 53.7435 6.4980 54.8370 ;
        RECT 6.3640 53.7435 6.3900 54.8370 ;
        RECT 6.2560 53.7435 6.2820 54.8370 ;
        RECT 6.1480 53.7435 6.1740 54.8370 ;
        RECT 6.0400 53.7435 6.0660 54.8370 ;
        RECT 5.9320 53.7435 5.9580 54.8370 ;
        RECT 5.8240 53.7435 5.8500 54.8370 ;
        RECT 5.7160 53.7435 5.7420 54.8370 ;
        RECT 5.6080 53.7435 5.6340 54.8370 ;
        RECT 5.5000 53.7435 5.5260 54.8370 ;
        RECT 5.3920 53.7435 5.4180 54.8370 ;
        RECT 5.2840 53.7435 5.3100 54.8370 ;
        RECT 5.1760 53.7435 5.2020 54.8370 ;
        RECT 5.0680 53.7435 5.0940 54.8370 ;
        RECT 4.9600 53.7435 4.9860 54.8370 ;
        RECT 4.8520 53.7435 4.8780 54.8370 ;
        RECT 4.7440 53.7435 4.7700 54.8370 ;
        RECT 4.6360 53.7435 4.6620 54.8370 ;
        RECT 4.5280 53.7435 4.5540 54.8370 ;
        RECT 4.4200 53.7435 4.4460 54.8370 ;
        RECT 4.3120 53.7435 4.3380 54.8370 ;
        RECT 4.2040 53.7435 4.2300 54.8370 ;
        RECT 4.0960 53.7435 4.1220 54.8370 ;
        RECT 3.9880 53.7435 4.0140 54.8370 ;
        RECT 3.8800 53.7435 3.9060 54.8370 ;
        RECT 3.7720 53.7435 3.7980 54.8370 ;
        RECT 3.6640 53.7435 3.6900 54.8370 ;
        RECT 3.5560 53.7435 3.5820 54.8370 ;
        RECT 3.4480 53.7435 3.4740 54.8370 ;
        RECT 3.3400 53.7435 3.3660 54.8370 ;
        RECT 3.2320 53.7435 3.2580 54.8370 ;
        RECT 3.1240 53.7435 3.1500 54.8370 ;
        RECT 3.0160 53.7435 3.0420 54.8370 ;
        RECT 2.9080 53.7435 2.9340 54.8370 ;
        RECT 2.8000 53.7435 2.8260 54.8370 ;
        RECT 2.6920 53.7435 2.7180 54.8370 ;
        RECT 2.5840 53.7435 2.6100 54.8370 ;
        RECT 2.4760 53.7435 2.5020 54.8370 ;
        RECT 2.3680 53.7435 2.3940 54.8370 ;
        RECT 2.2600 53.7435 2.2860 54.8370 ;
        RECT 2.1520 53.7435 2.1780 54.8370 ;
        RECT 2.0440 53.7435 2.0700 54.8370 ;
        RECT 1.9360 53.7435 1.9620 54.8370 ;
        RECT 1.8280 53.7435 1.8540 54.8370 ;
        RECT 1.7200 53.7435 1.7460 54.8370 ;
        RECT 1.6120 53.7435 1.6380 54.8370 ;
        RECT 1.5040 53.7435 1.5300 54.8370 ;
        RECT 1.3960 53.7435 1.4220 54.8370 ;
        RECT 1.2880 53.7435 1.3140 54.8370 ;
        RECT 1.1800 53.7435 1.2060 54.8370 ;
        RECT 1.0720 53.7435 1.0980 54.8370 ;
        RECT 0.9640 53.7435 0.9900 54.8370 ;
        RECT 0.8560 53.7435 0.8820 54.8370 ;
        RECT 0.7480 53.7435 0.7740 54.8370 ;
        RECT 0.6400 53.7435 0.6660 54.8370 ;
        RECT 0.5320 53.7435 0.5580 54.8370 ;
        RECT 0.4240 53.7435 0.4500 54.8370 ;
        RECT 0.3160 53.7435 0.3420 54.8370 ;
        RECT 0.2080 53.7435 0.2340 54.8370 ;
        RECT 0.0050 53.7435 0.0900 54.8370 ;
        RECT 8.6410 54.8235 8.7690 55.9170 ;
        RECT 8.6270 55.4890 8.7690 55.8115 ;
        RECT 8.4790 55.2160 8.5410 55.9170 ;
        RECT 8.4650 55.5255 8.5410 55.6790 ;
        RECT 8.4790 54.8235 8.5050 55.9170 ;
        RECT 8.4790 54.9445 8.5190 55.1840 ;
        RECT 8.4790 54.8235 8.5410 54.9125 ;
        RECT 8.1820 55.2740 8.3880 55.9170 ;
        RECT 8.3620 54.8235 8.3880 55.9170 ;
        RECT 8.1820 55.5510 8.4020 55.8090 ;
        RECT 8.1820 54.8235 8.2800 55.9170 ;
        RECT 7.7650 54.8235 7.8480 55.9170 ;
        RECT 7.7650 54.9120 7.8620 55.8475 ;
        RECT 16.4440 54.8235 16.5290 55.9170 ;
        RECT 16.3000 54.8235 16.3260 55.9170 ;
        RECT 16.1920 54.8235 16.2180 55.9170 ;
        RECT 16.0840 54.8235 16.1100 55.9170 ;
        RECT 15.9760 54.8235 16.0020 55.9170 ;
        RECT 15.8680 54.8235 15.8940 55.9170 ;
        RECT 15.7600 54.8235 15.7860 55.9170 ;
        RECT 15.6520 54.8235 15.6780 55.9170 ;
        RECT 15.5440 54.8235 15.5700 55.9170 ;
        RECT 15.4360 54.8235 15.4620 55.9170 ;
        RECT 15.3280 54.8235 15.3540 55.9170 ;
        RECT 15.2200 54.8235 15.2460 55.9170 ;
        RECT 15.1120 54.8235 15.1380 55.9170 ;
        RECT 15.0040 54.8235 15.0300 55.9170 ;
        RECT 14.8960 54.8235 14.9220 55.9170 ;
        RECT 14.7880 54.8235 14.8140 55.9170 ;
        RECT 14.6800 54.8235 14.7060 55.9170 ;
        RECT 14.5720 54.8235 14.5980 55.9170 ;
        RECT 14.4640 54.8235 14.4900 55.9170 ;
        RECT 14.3560 54.8235 14.3820 55.9170 ;
        RECT 14.2480 54.8235 14.2740 55.9170 ;
        RECT 14.1400 54.8235 14.1660 55.9170 ;
        RECT 14.0320 54.8235 14.0580 55.9170 ;
        RECT 13.9240 54.8235 13.9500 55.9170 ;
        RECT 13.8160 54.8235 13.8420 55.9170 ;
        RECT 13.7080 54.8235 13.7340 55.9170 ;
        RECT 13.6000 54.8235 13.6260 55.9170 ;
        RECT 13.4920 54.8235 13.5180 55.9170 ;
        RECT 13.3840 54.8235 13.4100 55.9170 ;
        RECT 13.2760 54.8235 13.3020 55.9170 ;
        RECT 13.1680 54.8235 13.1940 55.9170 ;
        RECT 13.0600 54.8235 13.0860 55.9170 ;
        RECT 12.9520 54.8235 12.9780 55.9170 ;
        RECT 12.8440 54.8235 12.8700 55.9170 ;
        RECT 12.7360 54.8235 12.7620 55.9170 ;
        RECT 12.6280 54.8235 12.6540 55.9170 ;
        RECT 12.5200 54.8235 12.5460 55.9170 ;
        RECT 12.4120 54.8235 12.4380 55.9170 ;
        RECT 12.3040 54.8235 12.3300 55.9170 ;
        RECT 12.1960 54.8235 12.2220 55.9170 ;
        RECT 12.0880 54.8235 12.1140 55.9170 ;
        RECT 11.9800 54.8235 12.0060 55.9170 ;
        RECT 11.8720 54.8235 11.8980 55.9170 ;
        RECT 11.7640 54.8235 11.7900 55.9170 ;
        RECT 11.6560 54.8235 11.6820 55.9170 ;
        RECT 11.5480 54.8235 11.5740 55.9170 ;
        RECT 11.4400 54.8235 11.4660 55.9170 ;
        RECT 11.3320 54.8235 11.3580 55.9170 ;
        RECT 11.2240 54.8235 11.2500 55.9170 ;
        RECT 11.1160 54.8235 11.1420 55.9170 ;
        RECT 11.0080 54.8235 11.0340 55.9170 ;
        RECT 10.9000 54.8235 10.9260 55.9170 ;
        RECT 10.7920 54.8235 10.8180 55.9170 ;
        RECT 10.6840 54.8235 10.7100 55.9170 ;
        RECT 10.5760 54.8235 10.6020 55.9170 ;
        RECT 10.4680 54.8235 10.4940 55.9170 ;
        RECT 10.3600 54.8235 10.3860 55.9170 ;
        RECT 10.2520 54.8235 10.2780 55.9170 ;
        RECT 10.1440 54.8235 10.1700 55.9170 ;
        RECT 10.0360 54.8235 10.0620 55.9170 ;
        RECT 9.9280 54.8235 9.9540 55.9170 ;
        RECT 9.8200 54.8235 9.8460 55.9170 ;
        RECT 9.7120 54.8235 9.7380 55.9170 ;
        RECT 9.6040 54.8235 9.6300 55.9170 ;
        RECT 9.4960 54.8235 9.5220 55.9170 ;
        RECT 9.3880 54.8235 9.4140 55.9170 ;
        RECT 9.1750 54.8235 9.2520 55.9170 ;
        RECT 7.2820 54.8235 7.3590 55.9170 ;
        RECT 7.1200 54.8235 7.1460 55.9170 ;
        RECT 7.0120 54.8235 7.0380 55.9170 ;
        RECT 6.9040 54.8235 6.9300 55.9170 ;
        RECT 6.7960 54.8235 6.8220 55.9170 ;
        RECT 6.6880 54.8235 6.7140 55.9170 ;
        RECT 6.5800 54.8235 6.6060 55.9170 ;
        RECT 6.4720 54.8235 6.4980 55.9170 ;
        RECT 6.3640 54.8235 6.3900 55.9170 ;
        RECT 6.2560 54.8235 6.2820 55.9170 ;
        RECT 6.1480 54.8235 6.1740 55.9170 ;
        RECT 6.0400 54.8235 6.0660 55.9170 ;
        RECT 5.9320 54.8235 5.9580 55.9170 ;
        RECT 5.8240 54.8235 5.8500 55.9170 ;
        RECT 5.7160 54.8235 5.7420 55.9170 ;
        RECT 5.6080 54.8235 5.6340 55.9170 ;
        RECT 5.5000 54.8235 5.5260 55.9170 ;
        RECT 5.3920 54.8235 5.4180 55.9170 ;
        RECT 5.2840 54.8235 5.3100 55.9170 ;
        RECT 5.1760 54.8235 5.2020 55.9170 ;
        RECT 5.0680 54.8235 5.0940 55.9170 ;
        RECT 4.9600 54.8235 4.9860 55.9170 ;
        RECT 4.8520 54.8235 4.8780 55.9170 ;
        RECT 4.7440 54.8235 4.7700 55.9170 ;
        RECT 4.6360 54.8235 4.6620 55.9170 ;
        RECT 4.5280 54.8235 4.5540 55.9170 ;
        RECT 4.4200 54.8235 4.4460 55.9170 ;
        RECT 4.3120 54.8235 4.3380 55.9170 ;
        RECT 4.2040 54.8235 4.2300 55.9170 ;
        RECT 4.0960 54.8235 4.1220 55.9170 ;
        RECT 3.9880 54.8235 4.0140 55.9170 ;
        RECT 3.8800 54.8235 3.9060 55.9170 ;
        RECT 3.7720 54.8235 3.7980 55.9170 ;
        RECT 3.6640 54.8235 3.6900 55.9170 ;
        RECT 3.5560 54.8235 3.5820 55.9170 ;
        RECT 3.4480 54.8235 3.4740 55.9170 ;
        RECT 3.3400 54.8235 3.3660 55.9170 ;
        RECT 3.2320 54.8235 3.2580 55.9170 ;
        RECT 3.1240 54.8235 3.1500 55.9170 ;
        RECT 3.0160 54.8235 3.0420 55.9170 ;
        RECT 2.9080 54.8235 2.9340 55.9170 ;
        RECT 2.8000 54.8235 2.8260 55.9170 ;
        RECT 2.6920 54.8235 2.7180 55.9170 ;
        RECT 2.5840 54.8235 2.6100 55.9170 ;
        RECT 2.4760 54.8235 2.5020 55.9170 ;
        RECT 2.3680 54.8235 2.3940 55.9170 ;
        RECT 2.2600 54.8235 2.2860 55.9170 ;
        RECT 2.1520 54.8235 2.1780 55.9170 ;
        RECT 2.0440 54.8235 2.0700 55.9170 ;
        RECT 1.9360 54.8235 1.9620 55.9170 ;
        RECT 1.8280 54.8235 1.8540 55.9170 ;
        RECT 1.7200 54.8235 1.7460 55.9170 ;
        RECT 1.6120 54.8235 1.6380 55.9170 ;
        RECT 1.5040 54.8235 1.5300 55.9170 ;
        RECT 1.3960 54.8235 1.4220 55.9170 ;
        RECT 1.2880 54.8235 1.3140 55.9170 ;
        RECT 1.1800 54.8235 1.2060 55.9170 ;
        RECT 1.0720 54.8235 1.0980 55.9170 ;
        RECT 0.9640 54.8235 0.9900 55.9170 ;
        RECT 0.8560 54.8235 0.8820 55.9170 ;
        RECT 0.7480 54.8235 0.7740 55.9170 ;
        RECT 0.6400 54.8235 0.6660 55.9170 ;
        RECT 0.5320 54.8235 0.5580 55.9170 ;
        RECT 0.4240 54.8235 0.4500 55.9170 ;
        RECT 0.3160 54.8235 0.3420 55.9170 ;
        RECT 0.2080 54.8235 0.2340 55.9170 ;
        RECT 0.0050 54.8235 0.0900 55.9170 ;
        RECT 8.6410 55.9035 8.7690 56.9970 ;
        RECT 8.6270 56.5690 8.7690 56.8915 ;
        RECT 8.4790 56.2960 8.5410 56.9970 ;
        RECT 8.4650 56.6055 8.5410 56.7590 ;
        RECT 8.4790 55.9035 8.5050 56.9970 ;
        RECT 8.4790 56.0245 8.5190 56.2640 ;
        RECT 8.4790 55.9035 8.5410 55.9925 ;
        RECT 8.1820 56.3540 8.3880 56.9970 ;
        RECT 8.3620 55.9035 8.3880 56.9970 ;
        RECT 8.1820 56.6310 8.4020 56.8890 ;
        RECT 8.1820 55.9035 8.2800 56.9970 ;
        RECT 7.7650 55.9035 7.8480 56.9970 ;
        RECT 7.7650 55.9920 7.8620 56.9275 ;
        RECT 16.4440 55.9035 16.5290 56.9970 ;
        RECT 16.3000 55.9035 16.3260 56.9970 ;
        RECT 16.1920 55.9035 16.2180 56.9970 ;
        RECT 16.0840 55.9035 16.1100 56.9970 ;
        RECT 15.9760 55.9035 16.0020 56.9970 ;
        RECT 15.8680 55.9035 15.8940 56.9970 ;
        RECT 15.7600 55.9035 15.7860 56.9970 ;
        RECT 15.6520 55.9035 15.6780 56.9970 ;
        RECT 15.5440 55.9035 15.5700 56.9970 ;
        RECT 15.4360 55.9035 15.4620 56.9970 ;
        RECT 15.3280 55.9035 15.3540 56.9970 ;
        RECT 15.2200 55.9035 15.2460 56.9970 ;
        RECT 15.1120 55.9035 15.1380 56.9970 ;
        RECT 15.0040 55.9035 15.0300 56.9970 ;
        RECT 14.8960 55.9035 14.9220 56.9970 ;
        RECT 14.7880 55.9035 14.8140 56.9970 ;
        RECT 14.6800 55.9035 14.7060 56.9970 ;
        RECT 14.5720 55.9035 14.5980 56.9970 ;
        RECT 14.4640 55.9035 14.4900 56.9970 ;
        RECT 14.3560 55.9035 14.3820 56.9970 ;
        RECT 14.2480 55.9035 14.2740 56.9970 ;
        RECT 14.1400 55.9035 14.1660 56.9970 ;
        RECT 14.0320 55.9035 14.0580 56.9970 ;
        RECT 13.9240 55.9035 13.9500 56.9970 ;
        RECT 13.8160 55.9035 13.8420 56.9970 ;
        RECT 13.7080 55.9035 13.7340 56.9970 ;
        RECT 13.6000 55.9035 13.6260 56.9970 ;
        RECT 13.4920 55.9035 13.5180 56.9970 ;
        RECT 13.3840 55.9035 13.4100 56.9970 ;
        RECT 13.2760 55.9035 13.3020 56.9970 ;
        RECT 13.1680 55.9035 13.1940 56.9970 ;
        RECT 13.0600 55.9035 13.0860 56.9970 ;
        RECT 12.9520 55.9035 12.9780 56.9970 ;
        RECT 12.8440 55.9035 12.8700 56.9970 ;
        RECT 12.7360 55.9035 12.7620 56.9970 ;
        RECT 12.6280 55.9035 12.6540 56.9970 ;
        RECT 12.5200 55.9035 12.5460 56.9970 ;
        RECT 12.4120 55.9035 12.4380 56.9970 ;
        RECT 12.3040 55.9035 12.3300 56.9970 ;
        RECT 12.1960 55.9035 12.2220 56.9970 ;
        RECT 12.0880 55.9035 12.1140 56.9970 ;
        RECT 11.9800 55.9035 12.0060 56.9970 ;
        RECT 11.8720 55.9035 11.8980 56.9970 ;
        RECT 11.7640 55.9035 11.7900 56.9970 ;
        RECT 11.6560 55.9035 11.6820 56.9970 ;
        RECT 11.5480 55.9035 11.5740 56.9970 ;
        RECT 11.4400 55.9035 11.4660 56.9970 ;
        RECT 11.3320 55.9035 11.3580 56.9970 ;
        RECT 11.2240 55.9035 11.2500 56.9970 ;
        RECT 11.1160 55.9035 11.1420 56.9970 ;
        RECT 11.0080 55.9035 11.0340 56.9970 ;
        RECT 10.9000 55.9035 10.9260 56.9970 ;
        RECT 10.7920 55.9035 10.8180 56.9970 ;
        RECT 10.6840 55.9035 10.7100 56.9970 ;
        RECT 10.5760 55.9035 10.6020 56.9970 ;
        RECT 10.4680 55.9035 10.4940 56.9970 ;
        RECT 10.3600 55.9035 10.3860 56.9970 ;
        RECT 10.2520 55.9035 10.2780 56.9970 ;
        RECT 10.1440 55.9035 10.1700 56.9970 ;
        RECT 10.0360 55.9035 10.0620 56.9970 ;
        RECT 9.9280 55.9035 9.9540 56.9970 ;
        RECT 9.8200 55.9035 9.8460 56.9970 ;
        RECT 9.7120 55.9035 9.7380 56.9970 ;
        RECT 9.6040 55.9035 9.6300 56.9970 ;
        RECT 9.4960 55.9035 9.5220 56.9970 ;
        RECT 9.3880 55.9035 9.4140 56.9970 ;
        RECT 9.1750 55.9035 9.2520 56.9970 ;
        RECT 7.2820 55.9035 7.3590 56.9970 ;
        RECT 7.1200 55.9035 7.1460 56.9970 ;
        RECT 7.0120 55.9035 7.0380 56.9970 ;
        RECT 6.9040 55.9035 6.9300 56.9970 ;
        RECT 6.7960 55.9035 6.8220 56.9970 ;
        RECT 6.6880 55.9035 6.7140 56.9970 ;
        RECT 6.5800 55.9035 6.6060 56.9970 ;
        RECT 6.4720 55.9035 6.4980 56.9970 ;
        RECT 6.3640 55.9035 6.3900 56.9970 ;
        RECT 6.2560 55.9035 6.2820 56.9970 ;
        RECT 6.1480 55.9035 6.1740 56.9970 ;
        RECT 6.0400 55.9035 6.0660 56.9970 ;
        RECT 5.9320 55.9035 5.9580 56.9970 ;
        RECT 5.8240 55.9035 5.8500 56.9970 ;
        RECT 5.7160 55.9035 5.7420 56.9970 ;
        RECT 5.6080 55.9035 5.6340 56.9970 ;
        RECT 5.5000 55.9035 5.5260 56.9970 ;
        RECT 5.3920 55.9035 5.4180 56.9970 ;
        RECT 5.2840 55.9035 5.3100 56.9970 ;
        RECT 5.1760 55.9035 5.2020 56.9970 ;
        RECT 5.0680 55.9035 5.0940 56.9970 ;
        RECT 4.9600 55.9035 4.9860 56.9970 ;
        RECT 4.8520 55.9035 4.8780 56.9970 ;
        RECT 4.7440 55.9035 4.7700 56.9970 ;
        RECT 4.6360 55.9035 4.6620 56.9970 ;
        RECT 4.5280 55.9035 4.5540 56.9970 ;
        RECT 4.4200 55.9035 4.4460 56.9970 ;
        RECT 4.3120 55.9035 4.3380 56.9970 ;
        RECT 4.2040 55.9035 4.2300 56.9970 ;
        RECT 4.0960 55.9035 4.1220 56.9970 ;
        RECT 3.9880 55.9035 4.0140 56.9970 ;
        RECT 3.8800 55.9035 3.9060 56.9970 ;
        RECT 3.7720 55.9035 3.7980 56.9970 ;
        RECT 3.6640 55.9035 3.6900 56.9970 ;
        RECT 3.5560 55.9035 3.5820 56.9970 ;
        RECT 3.4480 55.9035 3.4740 56.9970 ;
        RECT 3.3400 55.9035 3.3660 56.9970 ;
        RECT 3.2320 55.9035 3.2580 56.9970 ;
        RECT 3.1240 55.9035 3.1500 56.9970 ;
        RECT 3.0160 55.9035 3.0420 56.9970 ;
        RECT 2.9080 55.9035 2.9340 56.9970 ;
        RECT 2.8000 55.9035 2.8260 56.9970 ;
        RECT 2.6920 55.9035 2.7180 56.9970 ;
        RECT 2.5840 55.9035 2.6100 56.9970 ;
        RECT 2.4760 55.9035 2.5020 56.9970 ;
        RECT 2.3680 55.9035 2.3940 56.9970 ;
        RECT 2.2600 55.9035 2.2860 56.9970 ;
        RECT 2.1520 55.9035 2.1780 56.9970 ;
        RECT 2.0440 55.9035 2.0700 56.9970 ;
        RECT 1.9360 55.9035 1.9620 56.9970 ;
        RECT 1.8280 55.9035 1.8540 56.9970 ;
        RECT 1.7200 55.9035 1.7460 56.9970 ;
        RECT 1.6120 55.9035 1.6380 56.9970 ;
        RECT 1.5040 55.9035 1.5300 56.9970 ;
        RECT 1.3960 55.9035 1.4220 56.9970 ;
        RECT 1.2880 55.9035 1.3140 56.9970 ;
        RECT 1.1800 55.9035 1.2060 56.9970 ;
        RECT 1.0720 55.9035 1.0980 56.9970 ;
        RECT 0.9640 55.9035 0.9900 56.9970 ;
        RECT 0.8560 55.9035 0.8820 56.9970 ;
        RECT 0.7480 55.9035 0.7740 56.9970 ;
        RECT 0.6400 55.9035 0.6660 56.9970 ;
        RECT 0.5320 55.9035 0.5580 56.9970 ;
        RECT 0.4240 55.9035 0.4500 56.9970 ;
        RECT 0.3160 55.9035 0.3420 56.9970 ;
        RECT 0.2080 55.9035 0.2340 56.9970 ;
        RECT 0.0050 55.9035 0.0900 56.9970 ;
        RECT 8.6410 56.9835 8.7690 58.0770 ;
        RECT 8.6270 57.6490 8.7690 57.9715 ;
        RECT 8.4790 57.3760 8.5410 58.0770 ;
        RECT 8.4650 57.6855 8.5410 57.8390 ;
        RECT 8.4790 56.9835 8.5050 58.0770 ;
        RECT 8.4790 57.1045 8.5190 57.3440 ;
        RECT 8.4790 56.9835 8.5410 57.0725 ;
        RECT 8.1820 57.4340 8.3880 58.0770 ;
        RECT 8.3620 56.9835 8.3880 58.0770 ;
        RECT 8.1820 57.7110 8.4020 57.9690 ;
        RECT 8.1820 56.9835 8.2800 58.0770 ;
        RECT 7.7650 56.9835 7.8480 58.0770 ;
        RECT 7.7650 57.0720 7.8620 58.0075 ;
        RECT 16.4440 56.9835 16.5290 58.0770 ;
        RECT 16.3000 56.9835 16.3260 58.0770 ;
        RECT 16.1920 56.9835 16.2180 58.0770 ;
        RECT 16.0840 56.9835 16.1100 58.0770 ;
        RECT 15.9760 56.9835 16.0020 58.0770 ;
        RECT 15.8680 56.9835 15.8940 58.0770 ;
        RECT 15.7600 56.9835 15.7860 58.0770 ;
        RECT 15.6520 56.9835 15.6780 58.0770 ;
        RECT 15.5440 56.9835 15.5700 58.0770 ;
        RECT 15.4360 56.9835 15.4620 58.0770 ;
        RECT 15.3280 56.9835 15.3540 58.0770 ;
        RECT 15.2200 56.9835 15.2460 58.0770 ;
        RECT 15.1120 56.9835 15.1380 58.0770 ;
        RECT 15.0040 56.9835 15.0300 58.0770 ;
        RECT 14.8960 56.9835 14.9220 58.0770 ;
        RECT 14.7880 56.9835 14.8140 58.0770 ;
        RECT 14.6800 56.9835 14.7060 58.0770 ;
        RECT 14.5720 56.9835 14.5980 58.0770 ;
        RECT 14.4640 56.9835 14.4900 58.0770 ;
        RECT 14.3560 56.9835 14.3820 58.0770 ;
        RECT 14.2480 56.9835 14.2740 58.0770 ;
        RECT 14.1400 56.9835 14.1660 58.0770 ;
        RECT 14.0320 56.9835 14.0580 58.0770 ;
        RECT 13.9240 56.9835 13.9500 58.0770 ;
        RECT 13.8160 56.9835 13.8420 58.0770 ;
        RECT 13.7080 56.9835 13.7340 58.0770 ;
        RECT 13.6000 56.9835 13.6260 58.0770 ;
        RECT 13.4920 56.9835 13.5180 58.0770 ;
        RECT 13.3840 56.9835 13.4100 58.0770 ;
        RECT 13.2760 56.9835 13.3020 58.0770 ;
        RECT 13.1680 56.9835 13.1940 58.0770 ;
        RECT 13.0600 56.9835 13.0860 58.0770 ;
        RECT 12.9520 56.9835 12.9780 58.0770 ;
        RECT 12.8440 56.9835 12.8700 58.0770 ;
        RECT 12.7360 56.9835 12.7620 58.0770 ;
        RECT 12.6280 56.9835 12.6540 58.0770 ;
        RECT 12.5200 56.9835 12.5460 58.0770 ;
        RECT 12.4120 56.9835 12.4380 58.0770 ;
        RECT 12.3040 56.9835 12.3300 58.0770 ;
        RECT 12.1960 56.9835 12.2220 58.0770 ;
        RECT 12.0880 56.9835 12.1140 58.0770 ;
        RECT 11.9800 56.9835 12.0060 58.0770 ;
        RECT 11.8720 56.9835 11.8980 58.0770 ;
        RECT 11.7640 56.9835 11.7900 58.0770 ;
        RECT 11.6560 56.9835 11.6820 58.0770 ;
        RECT 11.5480 56.9835 11.5740 58.0770 ;
        RECT 11.4400 56.9835 11.4660 58.0770 ;
        RECT 11.3320 56.9835 11.3580 58.0770 ;
        RECT 11.2240 56.9835 11.2500 58.0770 ;
        RECT 11.1160 56.9835 11.1420 58.0770 ;
        RECT 11.0080 56.9835 11.0340 58.0770 ;
        RECT 10.9000 56.9835 10.9260 58.0770 ;
        RECT 10.7920 56.9835 10.8180 58.0770 ;
        RECT 10.6840 56.9835 10.7100 58.0770 ;
        RECT 10.5760 56.9835 10.6020 58.0770 ;
        RECT 10.4680 56.9835 10.4940 58.0770 ;
        RECT 10.3600 56.9835 10.3860 58.0770 ;
        RECT 10.2520 56.9835 10.2780 58.0770 ;
        RECT 10.1440 56.9835 10.1700 58.0770 ;
        RECT 10.0360 56.9835 10.0620 58.0770 ;
        RECT 9.9280 56.9835 9.9540 58.0770 ;
        RECT 9.8200 56.9835 9.8460 58.0770 ;
        RECT 9.7120 56.9835 9.7380 58.0770 ;
        RECT 9.6040 56.9835 9.6300 58.0770 ;
        RECT 9.4960 56.9835 9.5220 58.0770 ;
        RECT 9.3880 56.9835 9.4140 58.0770 ;
        RECT 9.1750 56.9835 9.2520 58.0770 ;
        RECT 7.2820 56.9835 7.3590 58.0770 ;
        RECT 7.1200 56.9835 7.1460 58.0770 ;
        RECT 7.0120 56.9835 7.0380 58.0770 ;
        RECT 6.9040 56.9835 6.9300 58.0770 ;
        RECT 6.7960 56.9835 6.8220 58.0770 ;
        RECT 6.6880 56.9835 6.7140 58.0770 ;
        RECT 6.5800 56.9835 6.6060 58.0770 ;
        RECT 6.4720 56.9835 6.4980 58.0770 ;
        RECT 6.3640 56.9835 6.3900 58.0770 ;
        RECT 6.2560 56.9835 6.2820 58.0770 ;
        RECT 6.1480 56.9835 6.1740 58.0770 ;
        RECT 6.0400 56.9835 6.0660 58.0770 ;
        RECT 5.9320 56.9835 5.9580 58.0770 ;
        RECT 5.8240 56.9835 5.8500 58.0770 ;
        RECT 5.7160 56.9835 5.7420 58.0770 ;
        RECT 5.6080 56.9835 5.6340 58.0770 ;
        RECT 5.5000 56.9835 5.5260 58.0770 ;
        RECT 5.3920 56.9835 5.4180 58.0770 ;
        RECT 5.2840 56.9835 5.3100 58.0770 ;
        RECT 5.1760 56.9835 5.2020 58.0770 ;
        RECT 5.0680 56.9835 5.0940 58.0770 ;
        RECT 4.9600 56.9835 4.9860 58.0770 ;
        RECT 4.8520 56.9835 4.8780 58.0770 ;
        RECT 4.7440 56.9835 4.7700 58.0770 ;
        RECT 4.6360 56.9835 4.6620 58.0770 ;
        RECT 4.5280 56.9835 4.5540 58.0770 ;
        RECT 4.4200 56.9835 4.4460 58.0770 ;
        RECT 4.3120 56.9835 4.3380 58.0770 ;
        RECT 4.2040 56.9835 4.2300 58.0770 ;
        RECT 4.0960 56.9835 4.1220 58.0770 ;
        RECT 3.9880 56.9835 4.0140 58.0770 ;
        RECT 3.8800 56.9835 3.9060 58.0770 ;
        RECT 3.7720 56.9835 3.7980 58.0770 ;
        RECT 3.6640 56.9835 3.6900 58.0770 ;
        RECT 3.5560 56.9835 3.5820 58.0770 ;
        RECT 3.4480 56.9835 3.4740 58.0770 ;
        RECT 3.3400 56.9835 3.3660 58.0770 ;
        RECT 3.2320 56.9835 3.2580 58.0770 ;
        RECT 3.1240 56.9835 3.1500 58.0770 ;
        RECT 3.0160 56.9835 3.0420 58.0770 ;
        RECT 2.9080 56.9835 2.9340 58.0770 ;
        RECT 2.8000 56.9835 2.8260 58.0770 ;
        RECT 2.6920 56.9835 2.7180 58.0770 ;
        RECT 2.5840 56.9835 2.6100 58.0770 ;
        RECT 2.4760 56.9835 2.5020 58.0770 ;
        RECT 2.3680 56.9835 2.3940 58.0770 ;
        RECT 2.2600 56.9835 2.2860 58.0770 ;
        RECT 2.1520 56.9835 2.1780 58.0770 ;
        RECT 2.0440 56.9835 2.0700 58.0770 ;
        RECT 1.9360 56.9835 1.9620 58.0770 ;
        RECT 1.8280 56.9835 1.8540 58.0770 ;
        RECT 1.7200 56.9835 1.7460 58.0770 ;
        RECT 1.6120 56.9835 1.6380 58.0770 ;
        RECT 1.5040 56.9835 1.5300 58.0770 ;
        RECT 1.3960 56.9835 1.4220 58.0770 ;
        RECT 1.2880 56.9835 1.3140 58.0770 ;
        RECT 1.1800 56.9835 1.2060 58.0770 ;
        RECT 1.0720 56.9835 1.0980 58.0770 ;
        RECT 0.9640 56.9835 0.9900 58.0770 ;
        RECT 0.8560 56.9835 0.8820 58.0770 ;
        RECT 0.7480 56.9835 0.7740 58.0770 ;
        RECT 0.6400 56.9835 0.6660 58.0770 ;
        RECT 0.5320 56.9835 0.5580 58.0770 ;
        RECT 0.4240 56.9835 0.4500 58.0770 ;
        RECT 0.3160 56.9835 0.3420 58.0770 ;
        RECT 0.2080 56.9835 0.2340 58.0770 ;
        RECT 0.0050 56.9835 0.0900 58.0770 ;
        RECT 8.6410 58.0635 8.7690 59.1570 ;
        RECT 8.6270 58.7290 8.7690 59.0515 ;
        RECT 8.4790 58.4560 8.5410 59.1570 ;
        RECT 8.4650 58.7655 8.5410 58.9190 ;
        RECT 8.4790 58.0635 8.5050 59.1570 ;
        RECT 8.4790 58.1845 8.5190 58.4240 ;
        RECT 8.4790 58.0635 8.5410 58.1525 ;
        RECT 8.1820 58.5140 8.3880 59.1570 ;
        RECT 8.3620 58.0635 8.3880 59.1570 ;
        RECT 8.1820 58.7910 8.4020 59.0490 ;
        RECT 8.1820 58.0635 8.2800 59.1570 ;
        RECT 7.7650 58.0635 7.8480 59.1570 ;
        RECT 7.7650 58.1520 7.8620 59.0875 ;
        RECT 16.4440 58.0635 16.5290 59.1570 ;
        RECT 16.3000 58.0635 16.3260 59.1570 ;
        RECT 16.1920 58.0635 16.2180 59.1570 ;
        RECT 16.0840 58.0635 16.1100 59.1570 ;
        RECT 15.9760 58.0635 16.0020 59.1570 ;
        RECT 15.8680 58.0635 15.8940 59.1570 ;
        RECT 15.7600 58.0635 15.7860 59.1570 ;
        RECT 15.6520 58.0635 15.6780 59.1570 ;
        RECT 15.5440 58.0635 15.5700 59.1570 ;
        RECT 15.4360 58.0635 15.4620 59.1570 ;
        RECT 15.3280 58.0635 15.3540 59.1570 ;
        RECT 15.2200 58.0635 15.2460 59.1570 ;
        RECT 15.1120 58.0635 15.1380 59.1570 ;
        RECT 15.0040 58.0635 15.0300 59.1570 ;
        RECT 14.8960 58.0635 14.9220 59.1570 ;
        RECT 14.7880 58.0635 14.8140 59.1570 ;
        RECT 14.6800 58.0635 14.7060 59.1570 ;
        RECT 14.5720 58.0635 14.5980 59.1570 ;
        RECT 14.4640 58.0635 14.4900 59.1570 ;
        RECT 14.3560 58.0635 14.3820 59.1570 ;
        RECT 14.2480 58.0635 14.2740 59.1570 ;
        RECT 14.1400 58.0635 14.1660 59.1570 ;
        RECT 14.0320 58.0635 14.0580 59.1570 ;
        RECT 13.9240 58.0635 13.9500 59.1570 ;
        RECT 13.8160 58.0635 13.8420 59.1570 ;
        RECT 13.7080 58.0635 13.7340 59.1570 ;
        RECT 13.6000 58.0635 13.6260 59.1570 ;
        RECT 13.4920 58.0635 13.5180 59.1570 ;
        RECT 13.3840 58.0635 13.4100 59.1570 ;
        RECT 13.2760 58.0635 13.3020 59.1570 ;
        RECT 13.1680 58.0635 13.1940 59.1570 ;
        RECT 13.0600 58.0635 13.0860 59.1570 ;
        RECT 12.9520 58.0635 12.9780 59.1570 ;
        RECT 12.8440 58.0635 12.8700 59.1570 ;
        RECT 12.7360 58.0635 12.7620 59.1570 ;
        RECT 12.6280 58.0635 12.6540 59.1570 ;
        RECT 12.5200 58.0635 12.5460 59.1570 ;
        RECT 12.4120 58.0635 12.4380 59.1570 ;
        RECT 12.3040 58.0635 12.3300 59.1570 ;
        RECT 12.1960 58.0635 12.2220 59.1570 ;
        RECT 12.0880 58.0635 12.1140 59.1570 ;
        RECT 11.9800 58.0635 12.0060 59.1570 ;
        RECT 11.8720 58.0635 11.8980 59.1570 ;
        RECT 11.7640 58.0635 11.7900 59.1570 ;
        RECT 11.6560 58.0635 11.6820 59.1570 ;
        RECT 11.5480 58.0635 11.5740 59.1570 ;
        RECT 11.4400 58.0635 11.4660 59.1570 ;
        RECT 11.3320 58.0635 11.3580 59.1570 ;
        RECT 11.2240 58.0635 11.2500 59.1570 ;
        RECT 11.1160 58.0635 11.1420 59.1570 ;
        RECT 11.0080 58.0635 11.0340 59.1570 ;
        RECT 10.9000 58.0635 10.9260 59.1570 ;
        RECT 10.7920 58.0635 10.8180 59.1570 ;
        RECT 10.6840 58.0635 10.7100 59.1570 ;
        RECT 10.5760 58.0635 10.6020 59.1570 ;
        RECT 10.4680 58.0635 10.4940 59.1570 ;
        RECT 10.3600 58.0635 10.3860 59.1570 ;
        RECT 10.2520 58.0635 10.2780 59.1570 ;
        RECT 10.1440 58.0635 10.1700 59.1570 ;
        RECT 10.0360 58.0635 10.0620 59.1570 ;
        RECT 9.9280 58.0635 9.9540 59.1570 ;
        RECT 9.8200 58.0635 9.8460 59.1570 ;
        RECT 9.7120 58.0635 9.7380 59.1570 ;
        RECT 9.6040 58.0635 9.6300 59.1570 ;
        RECT 9.4960 58.0635 9.5220 59.1570 ;
        RECT 9.3880 58.0635 9.4140 59.1570 ;
        RECT 9.1750 58.0635 9.2520 59.1570 ;
        RECT 7.2820 58.0635 7.3590 59.1570 ;
        RECT 7.1200 58.0635 7.1460 59.1570 ;
        RECT 7.0120 58.0635 7.0380 59.1570 ;
        RECT 6.9040 58.0635 6.9300 59.1570 ;
        RECT 6.7960 58.0635 6.8220 59.1570 ;
        RECT 6.6880 58.0635 6.7140 59.1570 ;
        RECT 6.5800 58.0635 6.6060 59.1570 ;
        RECT 6.4720 58.0635 6.4980 59.1570 ;
        RECT 6.3640 58.0635 6.3900 59.1570 ;
        RECT 6.2560 58.0635 6.2820 59.1570 ;
        RECT 6.1480 58.0635 6.1740 59.1570 ;
        RECT 6.0400 58.0635 6.0660 59.1570 ;
        RECT 5.9320 58.0635 5.9580 59.1570 ;
        RECT 5.8240 58.0635 5.8500 59.1570 ;
        RECT 5.7160 58.0635 5.7420 59.1570 ;
        RECT 5.6080 58.0635 5.6340 59.1570 ;
        RECT 5.5000 58.0635 5.5260 59.1570 ;
        RECT 5.3920 58.0635 5.4180 59.1570 ;
        RECT 5.2840 58.0635 5.3100 59.1570 ;
        RECT 5.1760 58.0635 5.2020 59.1570 ;
        RECT 5.0680 58.0635 5.0940 59.1570 ;
        RECT 4.9600 58.0635 4.9860 59.1570 ;
        RECT 4.8520 58.0635 4.8780 59.1570 ;
        RECT 4.7440 58.0635 4.7700 59.1570 ;
        RECT 4.6360 58.0635 4.6620 59.1570 ;
        RECT 4.5280 58.0635 4.5540 59.1570 ;
        RECT 4.4200 58.0635 4.4460 59.1570 ;
        RECT 4.3120 58.0635 4.3380 59.1570 ;
        RECT 4.2040 58.0635 4.2300 59.1570 ;
        RECT 4.0960 58.0635 4.1220 59.1570 ;
        RECT 3.9880 58.0635 4.0140 59.1570 ;
        RECT 3.8800 58.0635 3.9060 59.1570 ;
        RECT 3.7720 58.0635 3.7980 59.1570 ;
        RECT 3.6640 58.0635 3.6900 59.1570 ;
        RECT 3.5560 58.0635 3.5820 59.1570 ;
        RECT 3.4480 58.0635 3.4740 59.1570 ;
        RECT 3.3400 58.0635 3.3660 59.1570 ;
        RECT 3.2320 58.0635 3.2580 59.1570 ;
        RECT 3.1240 58.0635 3.1500 59.1570 ;
        RECT 3.0160 58.0635 3.0420 59.1570 ;
        RECT 2.9080 58.0635 2.9340 59.1570 ;
        RECT 2.8000 58.0635 2.8260 59.1570 ;
        RECT 2.6920 58.0635 2.7180 59.1570 ;
        RECT 2.5840 58.0635 2.6100 59.1570 ;
        RECT 2.4760 58.0635 2.5020 59.1570 ;
        RECT 2.3680 58.0635 2.3940 59.1570 ;
        RECT 2.2600 58.0635 2.2860 59.1570 ;
        RECT 2.1520 58.0635 2.1780 59.1570 ;
        RECT 2.0440 58.0635 2.0700 59.1570 ;
        RECT 1.9360 58.0635 1.9620 59.1570 ;
        RECT 1.8280 58.0635 1.8540 59.1570 ;
        RECT 1.7200 58.0635 1.7460 59.1570 ;
        RECT 1.6120 58.0635 1.6380 59.1570 ;
        RECT 1.5040 58.0635 1.5300 59.1570 ;
        RECT 1.3960 58.0635 1.4220 59.1570 ;
        RECT 1.2880 58.0635 1.3140 59.1570 ;
        RECT 1.1800 58.0635 1.2060 59.1570 ;
        RECT 1.0720 58.0635 1.0980 59.1570 ;
        RECT 0.9640 58.0635 0.9900 59.1570 ;
        RECT 0.8560 58.0635 0.8820 59.1570 ;
        RECT 0.7480 58.0635 0.7740 59.1570 ;
        RECT 0.6400 58.0635 0.6660 59.1570 ;
        RECT 0.5320 58.0635 0.5580 59.1570 ;
        RECT 0.4240 58.0635 0.4500 59.1570 ;
        RECT 0.3160 58.0635 0.3420 59.1570 ;
        RECT 0.2080 58.0635 0.2340 59.1570 ;
        RECT 0.0050 58.0635 0.0900 59.1570 ;
        RECT 8.6410 59.1435 8.7690 60.2370 ;
        RECT 8.6270 59.8090 8.7690 60.1315 ;
        RECT 8.4790 59.5360 8.5410 60.2370 ;
        RECT 8.4650 59.8455 8.5410 59.9990 ;
        RECT 8.4790 59.1435 8.5050 60.2370 ;
        RECT 8.4790 59.2645 8.5190 59.5040 ;
        RECT 8.4790 59.1435 8.5410 59.2325 ;
        RECT 8.1820 59.5940 8.3880 60.2370 ;
        RECT 8.3620 59.1435 8.3880 60.2370 ;
        RECT 8.1820 59.8710 8.4020 60.1290 ;
        RECT 8.1820 59.1435 8.2800 60.2370 ;
        RECT 7.7650 59.1435 7.8480 60.2370 ;
        RECT 7.7650 59.2320 7.8620 60.1675 ;
        RECT 16.4440 59.1435 16.5290 60.2370 ;
        RECT 16.3000 59.1435 16.3260 60.2370 ;
        RECT 16.1920 59.1435 16.2180 60.2370 ;
        RECT 16.0840 59.1435 16.1100 60.2370 ;
        RECT 15.9760 59.1435 16.0020 60.2370 ;
        RECT 15.8680 59.1435 15.8940 60.2370 ;
        RECT 15.7600 59.1435 15.7860 60.2370 ;
        RECT 15.6520 59.1435 15.6780 60.2370 ;
        RECT 15.5440 59.1435 15.5700 60.2370 ;
        RECT 15.4360 59.1435 15.4620 60.2370 ;
        RECT 15.3280 59.1435 15.3540 60.2370 ;
        RECT 15.2200 59.1435 15.2460 60.2370 ;
        RECT 15.1120 59.1435 15.1380 60.2370 ;
        RECT 15.0040 59.1435 15.0300 60.2370 ;
        RECT 14.8960 59.1435 14.9220 60.2370 ;
        RECT 14.7880 59.1435 14.8140 60.2370 ;
        RECT 14.6800 59.1435 14.7060 60.2370 ;
        RECT 14.5720 59.1435 14.5980 60.2370 ;
        RECT 14.4640 59.1435 14.4900 60.2370 ;
        RECT 14.3560 59.1435 14.3820 60.2370 ;
        RECT 14.2480 59.1435 14.2740 60.2370 ;
        RECT 14.1400 59.1435 14.1660 60.2370 ;
        RECT 14.0320 59.1435 14.0580 60.2370 ;
        RECT 13.9240 59.1435 13.9500 60.2370 ;
        RECT 13.8160 59.1435 13.8420 60.2370 ;
        RECT 13.7080 59.1435 13.7340 60.2370 ;
        RECT 13.6000 59.1435 13.6260 60.2370 ;
        RECT 13.4920 59.1435 13.5180 60.2370 ;
        RECT 13.3840 59.1435 13.4100 60.2370 ;
        RECT 13.2760 59.1435 13.3020 60.2370 ;
        RECT 13.1680 59.1435 13.1940 60.2370 ;
        RECT 13.0600 59.1435 13.0860 60.2370 ;
        RECT 12.9520 59.1435 12.9780 60.2370 ;
        RECT 12.8440 59.1435 12.8700 60.2370 ;
        RECT 12.7360 59.1435 12.7620 60.2370 ;
        RECT 12.6280 59.1435 12.6540 60.2370 ;
        RECT 12.5200 59.1435 12.5460 60.2370 ;
        RECT 12.4120 59.1435 12.4380 60.2370 ;
        RECT 12.3040 59.1435 12.3300 60.2370 ;
        RECT 12.1960 59.1435 12.2220 60.2370 ;
        RECT 12.0880 59.1435 12.1140 60.2370 ;
        RECT 11.9800 59.1435 12.0060 60.2370 ;
        RECT 11.8720 59.1435 11.8980 60.2370 ;
        RECT 11.7640 59.1435 11.7900 60.2370 ;
        RECT 11.6560 59.1435 11.6820 60.2370 ;
        RECT 11.5480 59.1435 11.5740 60.2370 ;
        RECT 11.4400 59.1435 11.4660 60.2370 ;
        RECT 11.3320 59.1435 11.3580 60.2370 ;
        RECT 11.2240 59.1435 11.2500 60.2370 ;
        RECT 11.1160 59.1435 11.1420 60.2370 ;
        RECT 11.0080 59.1435 11.0340 60.2370 ;
        RECT 10.9000 59.1435 10.9260 60.2370 ;
        RECT 10.7920 59.1435 10.8180 60.2370 ;
        RECT 10.6840 59.1435 10.7100 60.2370 ;
        RECT 10.5760 59.1435 10.6020 60.2370 ;
        RECT 10.4680 59.1435 10.4940 60.2370 ;
        RECT 10.3600 59.1435 10.3860 60.2370 ;
        RECT 10.2520 59.1435 10.2780 60.2370 ;
        RECT 10.1440 59.1435 10.1700 60.2370 ;
        RECT 10.0360 59.1435 10.0620 60.2370 ;
        RECT 9.9280 59.1435 9.9540 60.2370 ;
        RECT 9.8200 59.1435 9.8460 60.2370 ;
        RECT 9.7120 59.1435 9.7380 60.2370 ;
        RECT 9.6040 59.1435 9.6300 60.2370 ;
        RECT 9.4960 59.1435 9.5220 60.2370 ;
        RECT 9.3880 59.1435 9.4140 60.2370 ;
        RECT 9.1750 59.1435 9.2520 60.2370 ;
        RECT 7.2820 59.1435 7.3590 60.2370 ;
        RECT 7.1200 59.1435 7.1460 60.2370 ;
        RECT 7.0120 59.1435 7.0380 60.2370 ;
        RECT 6.9040 59.1435 6.9300 60.2370 ;
        RECT 6.7960 59.1435 6.8220 60.2370 ;
        RECT 6.6880 59.1435 6.7140 60.2370 ;
        RECT 6.5800 59.1435 6.6060 60.2370 ;
        RECT 6.4720 59.1435 6.4980 60.2370 ;
        RECT 6.3640 59.1435 6.3900 60.2370 ;
        RECT 6.2560 59.1435 6.2820 60.2370 ;
        RECT 6.1480 59.1435 6.1740 60.2370 ;
        RECT 6.0400 59.1435 6.0660 60.2370 ;
        RECT 5.9320 59.1435 5.9580 60.2370 ;
        RECT 5.8240 59.1435 5.8500 60.2370 ;
        RECT 5.7160 59.1435 5.7420 60.2370 ;
        RECT 5.6080 59.1435 5.6340 60.2370 ;
        RECT 5.5000 59.1435 5.5260 60.2370 ;
        RECT 5.3920 59.1435 5.4180 60.2370 ;
        RECT 5.2840 59.1435 5.3100 60.2370 ;
        RECT 5.1760 59.1435 5.2020 60.2370 ;
        RECT 5.0680 59.1435 5.0940 60.2370 ;
        RECT 4.9600 59.1435 4.9860 60.2370 ;
        RECT 4.8520 59.1435 4.8780 60.2370 ;
        RECT 4.7440 59.1435 4.7700 60.2370 ;
        RECT 4.6360 59.1435 4.6620 60.2370 ;
        RECT 4.5280 59.1435 4.5540 60.2370 ;
        RECT 4.4200 59.1435 4.4460 60.2370 ;
        RECT 4.3120 59.1435 4.3380 60.2370 ;
        RECT 4.2040 59.1435 4.2300 60.2370 ;
        RECT 4.0960 59.1435 4.1220 60.2370 ;
        RECT 3.9880 59.1435 4.0140 60.2370 ;
        RECT 3.8800 59.1435 3.9060 60.2370 ;
        RECT 3.7720 59.1435 3.7980 60.2370 ;
        RECT 3.6640 59.1435 3.6900 60.2370 ;
        RECT 3.5560 59.1435 3.5820 60.2370 ;
        RECT 3.4480 59.1435 3.4740 60.2370 ;
        RECT 3.3400 59.1435 3.3660 60.2370 ;
        RECT 3.2320 59.1435 3.2580 60.2370 ;
        RECT 3.1240 59.1435 3.1500 60.2370 ;
        RECT 3.0160 59.1435 3.0420 60.2370 ;
        RECT 2.9080 59.1435 2.9340 60.2370 ;
        RECT 2.8000 59.1435 2.8260 60.2370 ;
        RECT 2.6920 59.1435 2.7180 60.2370 ;
        RECT 2.5840 59.1435 2.6100 60.2370 ;
        RECT 2.4760 59.1435 2.5020 60.2370 ;
        RECT 2.3680 59.1435 2.3940 60.2370 ;
        RECT 2.2600 59.1435 2.2860 60.2370 ;
        RECT 2.1520 59.1435 2.1780 60.2370 ;
        RECT 2.0440 59.1435 2.0700 60.2370 ;
        RECT 1.9360 59.1435 1.9620 60.2370 ;
        RECT 1.8280 59.1435 1.8540 60.2370 ;
        RECT 1.7200 59.1435 1.7460 60.2370 ;
        RECT 1.6120 59.1435 1.6380 60.2370 ;
        RECT 1.5040 59.1435 1.5300 60.2370 ;
        RECT 1.3960 59.1435 1.4220 60.2370 ;
        RECT 1.2880 59.1435 1.3140 60.2370 ;
        RECT 1.1800 59.1435 1.2060 60.2370 ;
        RECT 1.0720 59.1435 1.0980 60.2370 ;
        RECT 0.9640 59.1435 0.9900 60.2370 ;
        RECT 0.8560 59.1435 0.8820 60.2370 ;
        RECT 0.7480 59.1435 0.7740 60.2370 ;
        RECT 0.6400 59.1435 0.6660 60.2370 ;
        RECT 0.5320 59.1435 0.5580 60.2370 ;
        RECT 0.4240 59.1435 0.4500 60.2370 ;
        RECT 0.3160 59.1435 0.3420 60.2370 ;
        RECT 0.2080 59.1435 0.2340 60.2370 ;
        RECT 0.0050 59.1435 0.0900 60.2370 ;
  LAYER V3 SPACING 0.018  ;
      RECT 0.0050 1.2200 16.5290 1.3500 ;
      RECT 16.4120 0.2565 16.5290 1.3500 ;
      RECT 9.3020 1.1240 16.3940 1.3500 ;
      RECT 7.9700 1.1240 9.2840 1.3500 ;
      RECT 7.2500 0.2565 7.8800 1.3500 ;
      RECT 0.1400 1.1240 7.2320 1.3500 ;
      RECT 0.0050 0.2565 0.1220 1.3500 ;
      RECT 16.3760 0.2565 16.5290 1.1720 ;
      RECT 9.3560 0.2565 16.3580 1.3500 ;
      RECT 8.6090 0.2565 9.3380 1.1720 ;
      RECT 8.4470 0.4520 8.5730 1.3500 ;
      RECT 7.1960 0.3560 8.4200 1.1720 ;
      RECT 0.1760 0.2565 7.1780 1.3500 ;
      RECT 0.0050 0.2565 0.1580 1.1720 ;
      RECT 8.5550 0.2565 16.5290 1.0760 ;
      RECT 0.0050 0.3560 8.5370 1.0760 ;
      RECT 8.3300 0.2565 16.5290 0.4280 ;
      RECT 0.0050 0.2565 8.3120 1.0760 ;
      RECT 0.0050 0.2565 16.5290 0.3320 ;
      RECT 0.0050 2.3000 16.5290 2.4300 ;
      RECT 16.4120 1.3365 16.5290 2.4300 ;
      RECT 9.3020 2.2040 16.3940 2.4300 ;
      RECT 7.9700 2.2040 9.2840 2.4300 ;
      RECT 7.2500 1.3365 7.8800 2.4300 ;
      RECT 0.1400 2.2040 7.2320 2.4300 ;
      RECT 0.0050 1.3365 0.1220 2.4300 ;
      RECT 16.3760 1.3365 16.5290 2.2520 ;
      RECT 9.3560 1.3365 16.3580 2.4300 ;
      RECT 8.6090 1.3365 9.3380 2.2520 ;
      RECT 8.4470 1.5320 8.5730 2.4300 ;
      RECT 7.1960 1.4360 8.4200 2.2520 ;
      RECT 0.1760 1.3365 7.1780 2.4300 ;
      RECT 0.0050 1.3365 0.1580 2.2520 ;
      RECT 8.5550 1.3365 16.5290 2.1560 ;
      RECT 0.0050 1.4360 8.5370 2.1560 ;
      RECT 8.3300 1.3365 16.5290 1.5080 ;
      RECT 0.0050 1.3365 8.3120 2.1560 ;
      RECT 0.0050 1.3365 16.5290 1.4120 ;
      RECT 0.0050 3.3800 16.5290 3.5100 ;
      RECT 16.4120 2.4165 16.5290 3.5100 ;
      RECT 9.3020 3.2840 16.3940 3.5100 ;
      RECT 7.9700 3.2840 9.2840 3.5100 ;
      RECT 7.2500 2.4165 7.8800 3.5100 ;
      RECT 0.1400 3.2840 7.2320 3.5100 ;
      RECT 0.0050 2.4165 0.1220 3.5100 ;
      RECT 16.3760 2.4165 16.5290 3.3320 ;
      RECT 9.3560 2.4165 16.3580 3.5100 ;
      RECT 8.6090 2.4165 9.3380 3.3320 ;
      RECT 8.4470 2.6120 8.5730 3.5100 ;
      RECT 7.1960 2.5160 8.4200 3.3320 ;
      RECT 0.1760 2.4165 7.1780 3.5100 ;
      RECT 0.0050 2.4165 0.1580 3.3320 ;
      RECT 8.5550 2.4165 16.5290 3.2360 ;
      RECT 0.0050 2.5160 8.5370 3.2360 ;
      RECT 8.3300 2.4165 16.5290 2.5880 ;
      RECT 0.0050 2.4165 8.3120 3.2360 ;
      RECT 0.0050 2.4165 16.5290 2.4920 ;
      RECT 0.0050 4.4600 16.5290 4.5900 ;
      RECT 16.4120 3.4965 16.5290 4.5900 ;
      RECT 9.3020 4.3640 16.3940 4.5900 ;
      RECT 7.9700 4.3640 9.2840 4.5900 ;
      RECT 7.2500 3.4965 7.8800 4.5900 ;
      RECT 0.1400 4.3640 7.2320 4.5900 ;
      RECT 0.0050 3.4965 0.1220 4.5900 ;
      RECT 16.3760 3.4965 16.5290 4.4120 ;
      RECT 9.3560 3.4965 16.3580 4.5900 ;
      RECT 8.6090 3.4965 9.3380 4.4120 ;
      RECT 8.4470 3.6920 8.5730 4.5900 ;
      RECT 7.1960 3.5960 8.4200 4.4120 ;
      RECT 0.1760 3.4965 7.1780 4.5900 ;
      RECT 0.0050 3.4965 0.1580 4.4120 ;
      RECT 8.5550 3.4965 16.5290 4.3160 ;
      RECT 0.0050 3.5960 8.5370 4.3160 ;
      RECT 8.3300 3.4965 16.5290 3.6680 ;
      RECT 0.0050 3.4965 8.3120 4.3160 ;
      RECT 0.0050 3.4965 16.5290 3.5720 ;
      RECT 0.0050 5.5400 16.5290 5.6700 ;
      RECT 16.4120 4.5765 16.5290 5.6700 ;
      RECT 9.3020 5.4440 16.3940 5.6700 ;
      RECT 7.9700 5.4440 9.2840 5.6700 ;
      RECT 7.2500 4.5765 7.8800 5.6700 ;
      RECT 0.1400 5.4440 7.2320 5.6700 ;
      RECT 0.0050 4.5765 0.1220 5.6700 ;
      RECT 16.3760 4.5765 16.5290 5.4920 ;
      RECT 9.3560 4.5765 16.3580 5.6700 ;
      RECT 8.6090 4.5765 9.3380 5.4920 ;
      RECT 8.4470 4.7720 8.5730 5.6700 ;
      RECT 7.1960 4.6760 8.4200 5.4920 ;
      RECT 0.1760 4.5765 7.1780 5.6700 ;
      RECT 0.0050 4.5765 0.1580 5.4920 ;
      RECT 8.5550 4.5765 16.5290 5.3960 ;
      RECT 0.0050 4.6760 8.5370 5.3960 ;
      RECT 8.3300 4.5765 16.5290 4.7480 ;
      RECT 0.0050 4.5765 8.3120 5.3960 ;
      RECT 0.0050 4.5765 16.5290 4.6520 ;
      RECT 0.0050 6.6200 16.5290 6.7500 ;
      RECT 16.4120 5.6565 16.5290 6.7500 ;
      RECT 9.3020 6.5240 16.3940 6.7500 ;
      RECT 7.9700 6.5240 9.2840 6.7500 ;
      RECT 7.2500 5.6565 7.8800 6.7500 ;
      RECT 0.1400 6.5240 7.2320 6.7500 ;
      RECT 0.0050 5.6565 0.1220 6.7500 ;
      RECT 16.3760 5.6565 16.5290 6.5720 ;
      RECT 9.3560 5.6565 16.3580 6.7500 ;
      RECT 8.6090 5.6565 9.3380 6.5720 ;
      RECT 8.4470 5.8520 8.5730 6.7500 ;
      RECT 7.1960 5.7560 8.4200 6.5720 ;
      RECT 0.1760 5.6565 7.1780 6.7500 ;
      RECT 0.0050 5.6565 0.1580 6.5720 ;
      RECT 8.5550 5.6565 16.5290 6.4760 ;
      RECT 0.0050 5.7560 8.5370 6.4760 ;
      RECT 8.3300 5.6565 16.5290 5.8280 ;
      RECT 0.0050 5.6565 8.3120 6.4760 ;
      RECT 0.0050 5.6565 16.5290 5.7320 ;
      RECT 0.0050 7.7000 16.5290 7.8300 ;
      RECT 16.4120 6.7365 16.5290 7.8300 ;
      RECT 9.3020 7.6040 16.3940 7.8300 ;
      RECT 7.9700 7.6040 9.2840 7.8300 ;
      RECT 7.2500 6.7365 7.8800 7.8300 ;
      RECT 0.1400 7.6040 7.2320 7.8300 ;
      RECT 0.0050 6.7365 0.1220 7.8300 ;
      RECT 16.3760 6.7365 16.5290 7.6520 ;
      RECT 9.3560 6.7365 16.3580 7.8300 ;
      RECT 8.6090 6.7365 9.3380 7.6520 ;
      RECT 8.4470 6.9320 8.5730 7.8300 ;
      RECT 7.1960 6.8360 8.4200 7.6520 ;
      RECT 0.1760 6.7365 7.1780 7.8300 ;
      RECT 0.0050 6.7365 0.1580 7.6520 ;
      RECT 8.5550 6.7365 16.5290 7.5560 ;
      RECT 0.0050 6.8360 8.5370 7.5560 ;
      RECT 8.3300 6.7365 16.5290 6.9080 ;
      RECT 0.0050 6.7365 8.3120 7.5560 ;
      RECT 0.0050 6.7365 16.5290 6.8120 ;
      RECT 0.0050 8.7800 16.5290 8.9100 ;
      RECT 16.4120 7.8165 16.5290 8.9100 ;
      RECT 9.3020 8.6840 16.3940 8.9100 ;
      RECT 7.9700 8.6840 9.2840 8.9100 ;
      RECT 7.2500 7.8165 7.8800 8.9100 ;
      RECT 0.1400 8.6840 7.2320 8.9100 ;
      RECT 0.0050 7.8165 0.1220 8.9100 ;
      RECT 16.3760 7.8165 16.5290 8.7320 ;
      RECT 9.3560 7.8165 16.3580 8.9100 ;
      RECT 8.6090 7.8165 9.3380 8.7320 ;
      RECT 8.4470 8.0120 8.5730 8.9100 ;
      RECT 7.1960 7.9160 8.4200 8.7320 ;
      RECT 0.1760 7.8165 7.1780 8.9100 ;
      RECT 0.0050 7.8165 0.1580 8.7320 ;
      RECT 8.5550 7.8165 16.5290 8.6360 ;
      RECT 0.0050 7.9160 8.5370 8.6360 ;
      RECT 8.3300 7.8165 16.5290 7.9880 ;
      RECT 0.0050 7.8165 8.3120 8.6360 ;
      RECT 0.0050 7.8165 16.5290 7.8920 ;
      RECT 0.0050 9.8600 16.5290 9.9900 ;
      RECT 16.4120 8.8965 16.5290 9.9900 ;
      RECT 9.3020 9.7640 16.3940 9.9900 ;
      RECT 7.9700 9.7640 9.2840 9.9900 ;
      RECT 7.2500 8.8965 7.8800 9.9900 ;
      RECT 0.1400 9.7640 7.2320 9.9900 ;
      RECT 0.0050 8.8965 0.1220 9.9900 ;
      RECT 16.3760 8.8965 16.5290 9.8120 ;
      RECT 9.3560 8.8965 16.3580 9.9900 ;
      RECT 8.6090 8.8965 9.3380 9.8120 ;
      RECT 8.4470 9.0920 8.5730 9.9900 ;
      RECT 7.1960 8.9960 8.4200 9.8120 ;
      RECT 0.1760 8.8965 7.1780 9.9900 ;
      RECT 0.0050 8.8965 0.1580 9.8120 ;
      RECT 8.5550 8.8965 16.5290 9.7160 ;
      RECT 0.0050 8.9960 8.5370 9.7160 ;
      RECT 8.3300 8.8965 16.5290 9.0680 ;
      RECT 0.0050 8.8965 8.3120 9.7160 ;
      RECT 0.0050 8.8965 16.5290 8.9720 ;
      RECT 0.0050 10.9400 16.5290 11.0700 ;
      RECT 16.4120 9.9765 16.5290 11.0700 ;
      RECT 9.3020 10.8440 16.3940 11.0700 ;
      RECT 7.9700 10.8440 9.2840 11.0700 ;
      RECT 7.2500 9.9765 7.8800 11.0700 ;
      RECT 0.1400 10.8440 7.2320 11.0700 ;
      RECT 0.0050 9.9765 0.1220 11.0700 ;
      RECT 16.3760 9.9765 16.5290 10.8920 ;
      RECT 9.3560 9.9765 16.3580 11.0700 ;
      RECT 8.6090 9.9765 9.3380 10.8920 ;
      RECT 8.4470 10.1720 8.5730 11.0700 ;
      RECT 7.1960 10.0760 8.4200 10.8920 ;
      RECT 0.1760 9.9765 7.1780 11.0700 ;
      RECT 0.0050 9.9765 0.1580 10.8920 ;
      RECT 8.5550 9.9765 16.5290 10.7960 ;
      RECT 0.0050 10.0760 8.5370 10.7960 ;
      RECT 8.3300 9.9765 16.5290 10.1480 ;
      RECT 0.0050 9.9765 8.3120 10.7960 ;
      RECT 0.0050 9.9765 16.5290 10.0520 ;
      RECT 0.0050 12.0200 16.5290 12.1500 ;
      RECT 16.4120 11.0565 16.5290 12.1500 ;
      RECT 9.3020 11.9240 16.3940 12.1500 ;
      RECT 7.9700 11.9240 9.2840 12.1500 ;
      RECT 7.2500 11.0565 7.8800 12.1500 ;
      RECT 0.1400 11.9240 7.2320 12.1500 ;
      RECT 0.0050 11.0565 0.1220 12.1500 ;
      RECT 16.3760 11.0565 16.5290 11.9720 ;
      RECT 9.3560 11.0565 16.3580 12.1500 ;
      RECT 8.6090 11.0565 9.3380 11.9720 ;
      RECT 8.4470 11.2520 8.5730 12.1500 ;
      RECT 7.1960 11.1560 8.4200 11.9720 ;
      RECT 0.1760 11.0565 7.1780 12.1500 ;
      RECT 0.0050 11.0565 0.1580 11.9720 ;
      RECT 8.5550 11.0565 16.5290 11.8760 ;
      RECT 0.0050 11.1560 8.5370 11.8760 ;
      RECT 8.3300 11.0565 16.5290 11.2280 ;
      RECT 0.0050 11.0565 8.3120 11.8760 ;
      RECT 0.0050 11.0565 16.5290 11.1320 ;
      RECT 0.0050 13.1000 16.5290 13.2300 ;
      RECT 16.4120 12.1365 16.5290 13.2300 ;
      RECT 9.3020 13.0040 16.3940 13.2300 ;
      RECT 7.9700 13.0040 9.2840 13.2300 ;
      RECT 7.2500 12.1365 7.8800 13.2300 ;
      RECT 0.1400 13.0040 7.2320 13.2300 ;
      RECT 0.0050 12.1365 0.1220 13.2300 ;
      RECT 16.3760 12.1365 16.5290 13.0520 ;
      RECT 9.3560 12.1365 16.3580 13.2300 ;
      RECT 8.6090 12.1365 9.3380 13.0520 ;
      RECT 8.4470 12.3320 8.5730 13.2300 ;
      RECT 7.1960 12.2360 8.4200 13.0520 ;
      RECT 0.1760 12.1365 7.1780 13.2300 ;
      RECT 0.0050 12.1365 0.1580 13.0520 ;
      RECT 8.5550 12.1365 16.5290 12.9560 ;
      RECT 0.0050 12.2360 8.5370 12.9560 ;
      RECT 8.3300 12.1365 16.5290 12.3080 ;
      RECT 0.0050 12.1365 8.3120 12.9560 ;
      RECT 0.0050 12.1365 16.5290 12.2120 ;
      RECT 0.0050 14.1800 16.5290 14.3100 ;
      RECT 16.4120 13.2165 16.5290 14.3100 ;
      RECT 9.3020 14.0840 16.3940 14.3100 ;
      RECT 7.9700 14.0840 9.2840 14.3100 ;
      RECT 7.2500 13.2165 7.8800 14.3100 ;
      RECT 0.1400 14.0840 7.2320 14.3100 ;
      RECT 0.0050 13.2165 0.1220 14.3100 ;
      RECT 16.3760 13.2165 16.5290 14.1320 ;
      RECT 9.3560 13.2165 16.3580 14.3100 ;
      RECT 8.6090 13.2165 9.3380 14.1320 ;
      RECT 8.4470 13.4120 8.5730 14.3100 ;
      RECT 7.1960 13.3160 8.4200 14.1320 ;
      RECT 0.1760 13.2165 7.1780 14.3100 ;
      RECT 0.0050 13.2165 0.1580 14.1320 ;
      RECT 8.5550 13.2165 16.5290 14.0360 ;
      RECT 0.0050 13.3160 8.5370 14.0360 ;
      RECT 8.3300 13.2165 16.5290 13.3880 ;
      RECT 0.0050 13.2165 8.3120 14.0360 ;
      RECT 0.0050 13.2165 16.5290 13.2920 ;
      RECT 0.0050 15.2600 16.5290 15.3900 ;
      RECT 16.4120 14.2965 16.5290 15.3900 ;
      RECT 9.3020 15.1640 16.3940 15.3900 ;
      RECT 7.9700 15.1640 9.2840 15.3900 ;
      RECT 7.2500 14.2965 7.8800 15.3900 ;
      RECT 0.1400 15.1640 7.2320 15.3900 ;
      RECT 0.0050 14.2965 0.1220 15.3900 ;
      RECT 16.3760 14.2965 16.5290 15.2120 ;
      RECT 9.3560 14.2965 16.3580 15.3900 ;
      RECT 8.6090 14.2965 9.3380 15.2120 ;
      RECT 8.4470 14.4920 8.5730 15.3900 ;
      RECT 7.1960 14.3960 8.4200 15.2120 ;
      RECT 0.1760 14.2965 7.1780 15.3900 ;
      RECT 0.0050 14.2965 0.1580 15.2120 ;
      RECT 8.5550 14.2965 16.5290 15.1160 ;
      RECT 0.0050 14.3960 8.5370 15.1160 ;
      RECT 8.3300 14.2965 16.5290 14.4680 ;
      RECT 0.0050 14.2965 8.3120 15.1160 ;
      RECT 0.0050 14.2965 16.5290 14.3720 ;
      RECT 0.0050 16.3400 16.5290 16.4700 ;
      RECT 16.4120 15.3765 16.5290 16.4700 ;
      RECT 9.3020 16.2440 16.3940 16.4700 ;
      RECT 7.9700 16.2440 9.2840 16.4700 ;
      RECT 7.2500 15.3765 7.8800 16.4700 ;
      RECT 0.1400 16.2440 7.2320 16.4700 ;
      RECT 0.0050 15.3765 0.1220 16.4700 ;
      RECT 16.3760 15.3765 16.5290 16.2920 ;
      RECT 9.3560 15.3765 16.3580 16.4700 ;
      RECT 8.6090 15.3765 9.3380 16.2920 ;
      RECT 8.4470 15.5720 8.5730 16.4700 ;
      RECT 7.1960 15.4760 8.4200 16.2920 ;
      RECT 0.1760 15.3765 7.1780 16.4700 ;
      RECT 0.0050 15.3765 0.1580 16.2920 ;
      RECT 8.5550 15.3765 16.5290 16.1960 ;
      RECT 0.0050 15.4760 8.5370 16.1960 ;
      RECT 8.3300 15.3765 16.5290 15.5480 ;
      RECT 0.0050 15.3765 8.3120 16.1960 ;
      RECT 0.0050 15.3765 16.5290 15.4520 ;
      RECT 0.0050 17.4200 16.5290 17.5500 ;
      RECT 16.4120 16.4565 16.5290 17.5500 ;
      RECT 9.3020 17.3240 16.3940 17.5500 ;
      RECT 7.9700 17.3240 9.2840 17.5500 ;
      RECT 7.2500 16.4565 7.8800 17.5500 ;
      RECT 0.1400 17.3240 7.2320 17.5500 ;
      RECT 0.0050 16.4565 0.1220 17.5500 ;
      RECT 16.3760 16.4565 16.5290 17.3720 ;
      RECT 9.3560 16.4565 16.3580 17.5500 ;
      RECT 8.6090 16.4565 9.3380 17.3720 ;
      RECT 8.4470 16.6520 8.5730 17.5500 ;
      RECT 7.1960 16.5560 8.4200 17.3720 ;
      RECT 0.1760 16.4565 7.1780 17.5500 ;
      RECT 0.0050 16.4565 0.1580 17.3720 ;
      RECT 8.5550 16.4565 16.5290 17.2760 ;
      RECT 0.0050 16.5560 8.5370 17.2760 ;
      RECT 8.3300 16.4565 16.5290 16.6280 ;
      RECT 0.0050 16.4565 8.3120 17.2760 ;
      RECT 0.0050 16.4565 16.5290 16.5320 ;
      RECT 0.0050 18.5000 16.5290 18.6300 ;
      RECT 16.4120 17.5365 16.5290 18.6300 ;
      RECT 9.3020 18.4040 16.3940 18.6300 ;
      RECT 7.9700 18.4040 9.2840 18.6300 ;
      RECT 7.2500 17.5365 7.8800 18.6300 ;
      RECT 0.1400 18.4040 7.2320 18.6300 ;
      RECT 0.0050 17.5365 0.1220 18.6300 ;
      RECT 16.3760 17.5365 16.5290 18.4520 ;
      RECT 9.3560 17.5365 16.3580 18.6300 ;
      RECT 8.6090 17.5365 9.3380 18.4520 ;
      RECT 8.4470 17.7320 8.5730 18.6300 ;
      RECT 7.1960 17.6360 8.4200 18.4520 ;
      RECT 0.1760 17.5365 7.1780 18.6300 ;
      RECT 0.0050 17.5365 0.1580 18.4520 ;
      RECT 8.5550 17.5365 16.5290 18.3560 ;
      RECT 0.0050 17.6360 8.5370 18.3560 ;
      RECT 8.3300 17.5365 16.5290 17.7080 ;
      RECT 0.0050 17.5365 8.3120 18.3560 ;
      RECT 0.0050 17.5365 16.5290 17.6120 ;
      RECT 0.0050 19.5800 16.5290 19.7100 ;
      RECT 16.4120 18.6165 16.5290 19.7100 ;
      RECT 9.3020 19.4840 16.3940 19.7100 ;
      RECT 7.9700 19.4840 9.2840 19.7100 ;
      RECT 7.2500 18.6165 7.8800 19.7100 ;
      RECT 0.1400 19.4840 7.2320 19.7100 ;
      RECT 0.0050 18.6165 0.1220 19.7100 ;
      RECT 16.3760 18.6165 16.5290 19.5320 ;
      RECT 9.3560 18.6165 16.3580 19.7100 ;
      RECT 8.6090 18.6165 9.3380 19.5320 ;
      RECT 8.4470 18.8120 8.5730 19.7100 ;
      RECT 7.1960 18.7160 8.4200 19.5320 ;
      RECT 0.1760 18.6165 7.1780 19.7100 ;
      RECT 0.0050 18.6165 0.1580 19.5320 ;
      RECT 8.5550 18.6165 16.5290 19.4360 ;
      RECT 0.0050 18.7160 8.5370 19.4360 ;
      RECT 8.3300 18.6165 16.5290 18.7880 ;
      RECT 0.0050 18.6165 8.3120 19.4360 ;
      RECT 0.0050 18.6165 16.5290 18.6920 ;
      RECT 0.0050 20.6600 16.5290 20.7900 ;
      RECT 16.4120 19.6965 16.5290 20.7900 ;
      RECT 9.3020 20.5640 16.3940 20.7900 ;
      RECT 7.9700 20.5640 9.2840 20.7900 ;
      RECT 7.2500 19.6965 7.8800 20.7900 ;
      RECT 0.1400 20.5640 7.2320 20.7900 ;
      RECT 0.0050 19.6965 0.1220 20.7900 ;
      RECT 16.3760 19.6965 16.5290 20.6120 ;
      RECT 9.3560 19.6965 16.3580 20.7900 ;
      RECT 8.6090 19.6965 9.3380 20.6120 ;
      RECT 8.4470 19.8920 8.5730 20.7900 ;
      RECT 7.1960 19.7960 8.4200 20.6120 ;
      RECT 0.1760 19.6965 7.1780 20.7900 ;
      RECT 0.0050 19.6965 0.1580 20.6120 ;
      RECT 8.5550 19.6965 16.5290 20.5160 ;
      RECT 0.0050 19.7960 8.5370 20.5160 ;
      RECT 8.3300 19.6965 16.5290 19.8680 ;
      RECT 0.0050 19.6965 8.3120 20.5160 ;
      RECT 0.0050 19.6965 16.5290 19.7720 ;
      RECT 0.0050 21.7400 16.5290 21.8700 ;
      RECT 16.4120 20.7765 16.5290 21.8700 ;
      RECT 9.3020 21.6440 16.3940 21.8700 ;
      RECT 7.9700 21.6440 9.2840 21.8700 ;
      RECT 7.2500 20.7765 7.8800 21.8700 ;
      RECT 0.1400 21.6440 7.2320 21.8700 ;
      RECT 0.0050 20.7765 0.1220 21.8700 ;
      RECT 16.3760 20.7765 16.5290 21.6920 ;
      RECT 9.3560 20.7765 16.3580 21.8700 ;
      RECT 8.6090 20.7765 9.3380 21.6920 ;
      RECT 8.4470 20.9720 8.5730 21.8700 ;
      RECT 7.1960 20.8760 8.4200 21.6920 ;
      RECT 0.1760 20.7765 7.1780 21.8700 ;
      RECT 0.0050 20.7765 0.1580 21.6920 ;
      RECT 8.5550 20.7765 16.5290 21.5960 ;
      RECT 0.0050 20.8760 8.5370 21.5960 ;
      RECT 8.3300 20.7765 16.5290 20.9480 ;
      RECT 0.0050 20.7765 8.3120 21.5960 ;
      RECT 0.0050 20.7765 16.5290 20.8520 ;
      RECT 0.0050 22.8200 16.5290 22.9500 ;
      RECT 16.4120 21.8565 16.5290 22.9500 ;
      RECT 9.3020 22.7240 16.3940 22.9500 ;
      RECT 7.9700 22.7240 9.2840 22.9500 ;
      RECT 7.2500 21.8565 7.8800 22.9500 ;
      RECT 0.1400 22.7240 7.2320 22.9500 ;
      RECT 0.0050 21.8565 0.1220 22.9500 ;
      RECT 16.3760 21.8565 16.5290 22.7720 ;
      RECT 9.3560 21.8565 16.3580 22.9500 ;
      RECT 8.6090 21.8565 9.3380 22.7720 ;
      RECT 8.4470 22.0520 8.5730 22.9500 ;
      RECT 7.1960 21.9560 8.4200 22.7720 ;
      RECT 0.1760 21.8565 7.1780 22.9500 ;
      RECT 0.0050 21.8565 0.1580 22.7720 ;
      RECT 8.5550 21.8565 16.5290 22.6760 ;
      RECT 0.0050 21.9560 8.5370 22.6760 ;
      RECT 8.3300 21.8565 16.5290 22.0280 ;
      RECT 0.0050 21.8565 8.3120 22.6760 ;
      RECT 0.0050 21.8565 16.5290 21.9320 ;
      RECT 0.0050 23.9000 16.5290 24.0300 ;
      RECT 16.4120 22.9365 16.5290 24.0300 ;
      RECT 9.3020 23.8040 16.3940 24.0300 ;
      RECT 7.9700 23.8040 9.2840 24.0300 ;
      RECT 7.2500 22.9365 7.8800 24.0300 ;
      RECT 0.1400 23.8040 7.2320 24.0300 ;
      RECT 0.0050 22.9365 0.1220 24.0300 ;
      RECT 16.3760 22.9365 16.5290 23.8520 ;
      RECT 9.3560 22.9365 16.3580 24.0300 ;
      RECT 8.6090 22.9365 9.3380 23.8520 ;
      RECT 8.4470 23.1320 8.5730 24.0300 ;
      RECT 7.1960 23.0360 8.4200 23.8520 ;
      RECT 0.1760 22.9365 7.1780 24.0300 ;
      RECT 0.0050 22.9365 0.1580 23.8520 ;
      RECT 8.5550 22.9365 16.5290 23.7560 ;
      RECT 0.0050 23.0360 8.5370 23.7560 ;
      RECT 8.3300 22.9365 16.5290 23.1080 ;
      RECT 0.0050 22.9365 8.3120 23.7560 ;
      RECT 0.0050 22.9365 16.5290 23.0120 ;
      RECT 0.0050 24.9800 16.5290 25.1100 ;
      RECT 16.4120 24.0165 16.5290 25.1100 ;
      RECT 9.3020 24.8840 16.3940 25.1100 ;
      RECT 7.9700 24.8840 9.2840 25.1100 ;
      RECT 7.2500 24.0165 7.8800 25.1100 ;
      RECT 0.1400 24.8840 7.2320 25.1100 ;
      RECT 0.0050 24.0165 0.1220 25.1100 ;
      RECT 16.3760 24.0165 16.5290 24.9320 ;
      RECT 9.3560 24.0165 16.3580 25.1100 ;
      RECT 8.6090 24.0165 9.3380 24.9320 ;
      RECT 8.4470 24.2120 8.5730 25.1100 ;
      RECT 7.1960 24.1160 8.4200 24.9320 ;
      RECT 0.1760 24.0165 7.1780 25.1100 ;
      RECT 0.0050 24.0165 0.1580 24.9320 ;
      RECT 8.5550 24.0165 16.5290 24.8360 ;
      RECT 0.0050 24.1160 8.5370 24.8360 ;
      RECT 8.3300 24.0165 16.5290 24.1880 ;
      RECT 0.0050 24.0165 8.3120 24.8360 ;
      RECT 0.0050 24.0165 16.5290 24.0920 ;
      RECT 0.0050 26.0600 16.5290 26.1900 ;
      RECT 16.4120 25.0965 16.5290 26.1900 ;
      RECT 9.3020 25.9640 16.3940 26.1900 ;
      RECT 7.9700 25.9640 9.2840 26.1900 ;
      RECT 7.2500 25.0965 7.8800 26.1900 ;
      RECT 0.1400 25.9640 7.2320 26.1900 ;
      RECT 0.0050 25.0965 0.1220 26.1900 ;
      RECT 16.3760 25.0965 16.5290 26.0120 ;
      RECT 9.3560 25.0965 16.3580 26.1900 ;
      RECT 8.6090 25.0965 9.3380 26.0120 ;
      RECT 8.4470 25.2920 8.5730 26.1900 ;
      RECT 7.1960 25.1960 8.4200 26.0120 ;
      RECT 0.1760 25.0965 7.1780 26.1900 ;
      RECT 0.0050 25.0965 0.1580 26.0120 ;
      RECT 8.5550 25.0965 16.5290 25.9160 ;
      RECT 0.0050 25.1960 8.5370 25.9160 ;
      RECT 8.3300 25.0965 16.5290 25.2680 ;
      RECT 0.0050 25.0965 8.3120 25.9160 ;
      RECT 0.0050 25.0965 16.5290 25.1720 ;
      RECT 0.0000 33.4770 16.5240 34.8105 ;
      RECT 10.8090 26.1570 16.5240 34.8105 ;
      RECT 8.6090 30.0210 16.5240 34.8105 ;
      RECT 9.5130 27.4290 16.5240 34.8105 ;
      RECT 8.5570 26.1570 8.5910 34.8105 ;
      RECT 8.5050 26.1570 8.5390 34.8105 ;
      RECT 8.4530 26.1570 8.4870 34.8105 ;
      RECT 8.4010 26.1570 8.4350 34.8105 ;
      RECT 0.0000 33.0450 8.3830 34.8105 ;
      RECT 8.1410 30.3090 16.5240 33.2610 ;
      RECT 8.0890 26.1570 8.1230 34.8105 ;
      RECT 8.0370 26.1570 8.0710 34.8105 ;
      RECT 7.9850 26.1570 8.0190 34.8105 ;
      RECT 7.9330 26.1570 7.9670 34.8105 ;
      RECT 0.0000 27.7170 7.9150 34.8105 ;
      RECT 0.0000 29.8770 8.3830 32.8290 ;
      RECT 8.1410 27.1410 9.2790 30.0930 ;
      RECT 9.3150 27.6210 16.5240 34.8105 ;
      RECT 0.0000 29.8770 9.2970 30.0930 ;
      RECT 8.1410 27.6210 16.5240 29.9970 ;
      RECT 7.4610 26.7090 8.2350 29.6610 ;
      RECT 7.2450 26.8530 7.9150 34.8105 ;
      RECT 0.0000 27.4290 7.2270 34.8105 ;
      RECT 6.8130 26.1570 7.2630 27.6930 ;
      RECT 0.0000 27.5250 9.4950 27.6930 ;
      RECT 9.2970 27.4290 16.5240 27.5970 ;
      RECT 10.5930 26.1570 10.7910 34.8105 ;
      RECT 6.8130 27.2370 10.5750 27.5010 ;
      RECT 5.9490 26.8530 6.7950 34.8105 ;
      RECT 0.0000 26.1570 5.9310 34.8105 ;
      RECT 10.3770 26.1570 16.5240 27.4050 ;
      RECT 10.1610 26.8530 16.5240 27.4050 ;
      RECT 0.0000 27.1415 10.1430 27.4050 ;
      RECT 9.9450 26.1570 10.3590 27.2130 ;
      RECT 9.3510 26.8530 16.5240 27.2130 ;
      RECT 8.6090 26.8530 9.3330 27.5010 ;
      RECT 8.1410 26.8050 8.3830 34.8105 ;
      RECT 8.2530 26.1570 8.6310 26.9250 ;
      RECT 8.6490 26.8050 9.9270 26.9255 ;
      RECT 6.5970 26.8050 7.4430 27.4050 ;
      RECT 6.1650 26.8050 6.5790 34.8105 ;
      RECT 0.0000 26.1570 6.1470 27.4050 ;
      RECT 9.7290 26.1570 16.5240 26.8290 ;
      RECT 8.2530 26.2370 9.7110 26.8290 ;
      RECT 7.2810 26.7090 8.2350 26.8290 ;
      RECT 6.3810 26.1570 7.2630 26.8290 ;
      RECT 0.0000 26.1570 6.3630 26.8290 ;
      RECT 9.2970 26.1570 16.5240 26.7810 ;
      RECT 8.1410 26.2370 16.5240 26.7810 ;
      RECT 0.0000 26.1570 7.9150 26.7810 ;
      RECT 0.0000 26.1570 9.2790 26.4930 ;
      RECT 0.0000 26.1570 16.5240 26.2130 ;
        RECT 0.0050 35.2670 16.5290 35.3970 ;
        RECT 16.4120 34.3035 16.5290 35.3970 ;
        RECT 9.3020 35.1710 16.3940 35.3970 ;
        RECT 7.9700 35.1710 9.2840 35.3970 ;
        RECT 7.2500 34.3035 7.8800 35.3970 ;
        RECT 0.1400 35.1710 7.2320 35.3970 ;
        RECT 0.0050 34.3035 0.1220 35.3970 ;
        RECT 16.3760 34.3035 16.5290 35.2190 ;
        RECT 9.3560 34.3035 16.3580 35.3970 ;
        RECT 8.6090 34.3035 9.3380 35.2190 ;
        RECT 8.4470 34.4990 8.5730 35.3970 ;
        RECT 7.1960 34.4030 8.4200 35.2190 ;
        RECT 0.1760 34.3035 7.1780 35.3970 ;
        RECT 0.0050 34.3035 0.1580 35.2190 ;
        RECT 8.5550 34.3035 16.5290 35.1230 ;
        RECT 0.0050 34.4030 8.5370 35.1230 ;
        RECT 8.3300 34.3035 16.5290 34.4750 ;
        RECT 0.0050 34.3035 8.3120 35.1230 ;
        RECT 0.0050 34.3035 16.5290 34.3790 ;
        RECT 0.0050 36.3470 16.5290 36.4770 ;
        RECT 16.4120 35.3835 16.5290 36.4770 ;
        RECT 9.3020 36.2510 16.3940 36.4770 ;
        RECT 7.9700 36.2510 9.2840 36.4770 ;
        RECT 7.2500 35.3835 7.8800 36.4770 ;
        RECT 0.1400 36.2510 7.2320 36.4770 ;
        RECT 0.0050 35.3835 0.1220 36.4770 ;
        RECT 16.3760 35.3835 16.5290 36.2990 ;
        RECT 9.3560 35.3835 16.3580 36.4770 ;
        RECT 8.6090 35.3835 9.3380 36.2990 ;
        RECT 8.4470 35.5790 8.5730 36.4770 ;
        RECT 7.1960 35.4830 8.4200 36.2990 ;
        RECT 0.1760 35.3835 7.1780 36.4770 ;
        RECT 0.0050 35.3835 0.1580 36.2990 ;
        RECT 8.5550 35.3835 16.5290 36.2030 ;
        RECT 0.0050 35.4830 8.5370 36.2030 ;
        RECT 8.3300 35.3835 16.5290 35.5550 ;
        RECT 0.0050 35.3835 8.3120 36.2030 ;
        RECT 0.0050 35.3835 16.5290 35.4590 ;
        RECT 0.0050 37.4270 16.5290 37.5570 ;
        RECT 16.4120 36.4635 16.5290 37.5570 ;
        RECT 9.3020 37.3310 16.3940 37.5570 ;
        RECT 7.9700 37.3310 9.2840 37.5570 ;
        RECT 7.2500 36.4635 7.8800 37.5570 ;
        RECT 0.1400 37.3310 7.2320 37.5570 ;
        RECT 0.0050 36.4635 0.1220 37.5570 ;
        RECT 16.3760 36.4635 16.5290 37.3790 ;
        RECT 9.3560 36.4635 16.3580 37.5570 ;
        RECT 8.6090 36.4635 9.3380 37.3790 ;
        RECT 8.4470 36.6590 8.5730 37.5570 ;
        RECT 7.1960 36.5630 8.4200 37.3790 ;
        RECT 0.1760 36.4635 7.1780 37.5570 ;
        RECT 0.0050 36.4635 0.1580 37.3790 ;
        RECT 8.5550 36.4635 16.5290 37.2830 ;
        RECT 0.0050 36.5630 8.5370 37.2830 ;
        RECT 8.3300 36.4635 16.5290 36.6350 ;
        RECT 0.0050 36.4635 8.3120 37.2830 ;
        RECT 0.0050 36.4635 16.5290 36.5390 ;
        RECT 0.0050 38.5070 16.5290 38.6370 ;
        RECT 16.4120 37.5435 16.5290 38.6370 ;
        RECT 9.3020 38.4110 16.3940 38.6370 ;
        RECT 7.9700 38.4110 9.2840 38.6370 ;
        RECT 7.2500 37.5435 7.8800 38.6370 ;
        RECT 0.1400 38.4110 7.2320 38.6370 ;
        RECT 0.0050 37.5435 0.1220 38.6370 ;
        RECT 16.3760 37.5435 16.5290 38.4590 ;
        RECT 9.3560 37.5435 16.3580 38.6370 ;
        RECT 8.6090 37.5435 9.3380 38.4590 ;
        RECT 8.4470 37.7390 8.5730 38.6370 ;
        RECT 7.1960 37.6430 8.4200 38.4590 ;
        RECT 0.1760 37.5435 7.1780 38.6370 ;
        RECT 0.0050 37.5435 0.1580 38.4590 ;
        RECT 8.5550 37.5435 16.5290 38.3630 ;
        RECT 0.0050 37.6430 8.5370 38.3630 ;
        RECT 8.3300 37.5435 16.5290 37.7150 ;
        RECT 0.0050 37.5435 8.3120 38.3630 ;
        RECT 0.0050 37.5435 16.5290 37.6190 ;
        RECT 0.0050 39.5870 16.5290 39.7170 ;
        RECT 16.4120 38.6235 16.5290 39.7170 ;
        RECT 9.3020 39.4910 16.3940 39.7170 ;
        RECT 7.9700 39.4910 9.2840 39.7170 ;
        RECT 7.2500 38.6235 7.8800 39.7170 ;
        RECT 0.1400 39.4910 7.2320 39.7170 ;
        RECT 0.0050 38.6235 0.1220 39.7170 ;
        RECT 16.3760 38.6235 16.5290 39.5390 ;
        RECT 9.3560 38.6235 16.3580 39.7170 ;
        RECT 8.6090 38.6235 9.3380 39.5390 ;
        RECT 8.4470 38.8190 8.5730 39.7170 ;
        RECT 7.1960 38.7230 8.4200 39.5390 ;
        RECT 0.1760 38.6235 7.1780 39.7170 ;
        RECT 0.0050 38.6235 0.1580 39.5390 ;
        RECT 8.5550 38.6235 16.5290 39.4430 ;
        RECT 0.0050 38.7230 8.5370 39.4430 ;
        RECT 8.3300 38.6235 16.5290 38.7950 ;
        RECT 0.0050 38.6235 8.3120 39.4430 ;
        RECT 0.0050 38.6235 16.5290 38.6990 ;
        RECT 0.0050 40.6670 16.5290 40.7970 ;
        RECT 16.4120 39.7035 16.5290 40.7970 ;
        RECT 9.3020 40.5710 16.3940 40.7970 ;
        RECT 7.9700 40.5710 9.2840 40.7970 ;
        RECT 7.2500 39.7035 7.8800 40.7970 ;
        RECT 0.1400 40.5710 7.2320 40.7970 ;
        RECT 0.0050 39.7035 0.1220 40.7970 ;
        RECT 16.3760 39.7035 16.5290 40.6190 ;
        RECT 9.3560 39.7035 16.3580 40.7970 ;
        RECT 8.6090 39.7035 9.3380 40.6190 ;
        RECT 8.4470 39.8990 8.5730 40.7970 ;
        RECT 7.1960 39.8030 8.4200 40.6190 ;
        RECT 0.1760 39.7035 7.1780 40.7970 ;
        RECT 0.0050 39.7035 0.1580 40.6190 ;
        RECT 8.5550 39.7035 16.5290 40.5230 ;
        RECT 0.0050 39.8030 8.5370 40.5230 ;
        RECT 8.3300 39.7035 16.5290 39.8750 ;
        RECT 0.0050 39.7035 8.3120 40.5230 ;
        RECT 0.0050 39.7035 16.5290 39.7790 ;
        RECT 0.0050 41.7470 16.5290 41.8770 ;
        RECT 16.4120 40.7835 16.5290 41.8770 ;
        RECT 9.3020 41.6510 16.3940 41.8770 ;
        RECT 7.9700 41.6510 9.2840 41.8770 ;
        RECT 7.2500 40.7835 7.8800 41.8770 ;
        RECT 0.1400 41.6510 7.2320 41.8770 ;
        RECT 0.0050 40.7835 0.1220 41.8770 ;
        RECT 16.3760 40.7835 16.5290 41.6990 ;
        RECT 9.3560 40.7835 16.3580 41.8770 ;
        RECT 8.6090 40.7835 9.3380 41.6990 ;
        RECT 8.4470 40.9790 8.5730 41.8770 ;
        RECT 7.1960 40.8830 8.4200 41.6990 ;
        RECT 0.1760 40.7835 7.1780 41.8770 ;
        RECT 0.0050 40.7835 0.1580 41.6990 ;
        RECT 8.5550 40.7835 16.5290 41.6030 ;
        RECT 0.0050 40.8830 8.5370 41.6030 ;
        RECT 8.3300 40.7835 16.5290 40.9550 ;
        RECT 0.0050 40.7835 8.3120 41.6030 ;
        RECT 0.0050 40.7835 16.5290 40.8590 ;
        RECT 0.0050 42.8270 16.5290 42.9570 ;
        RECT 16.4120 41.8635 16.5290 42.9570 ;
        RECT 9.3020 42.7310 16.3940 42.9570 ;
        RECT 7.9700 42.7310 9.2840 42.9570 ;
        RECT 7.2500 41.8635 7.8800 42.9570 ;
        RECT 0.1400 42.7310 7.2320 42.9570 ;
        RECT 0.0050 41.8635 0.1220 42.9570 ;
        RECT 16.3760 41.8635 16.5290 42.7790 ;
        RECT 9.3560 41.8635 16.3580 42.9570 ;
        RECT 8.6090 41.8635 9.3380 42.7790 ;
        RECT 8.4470 42.0590 8.5730 42.9570 ;
        RECT 7.1960 41.9630 8.4200 42.7790 ;
        RECT 0.1760 41.8635 7.1780 42.9570 ;
        RECT 0.0050 41.8635 0.1580 42.7790 ;
        RECT 8.5550 41.8635 16.5290 42.6830 ;
        RECT 0.0050 41.9630 8.5370 42.6830 ;
        RECT 8.3300 41.8635 16.5290 42.0350 ;
        RECT 0.0050 41.8635 8.3120 42.6830 ;
        RECT 0.0050 41.8635 16.5290 41.9390 ;
        RECT 0.0050 43.9070 16.5290 44.0370 ;
        RECT 16.4120 42.9435 16.5290 44.0370 ;
        RECT 9.3020 43.8110 16.3940 44.0370 ;
        RECT 7.9700 43.8110 9.2840 44.0370 ;
        RECT 7.2500 42.9435 7.8800 44.0370 ;
        RECT 0.1400 43.8110 7.2320 44.0370 ;
        RECT 0.0050 42.9435 0.1220 44.0370 ;
        RECT 16.3760 42.9435 16.5290 43.8590 ;
        RECT 9.3560 42.9435 16.3580 44.0370 ;
        RECT 8.6090 42.9435 9.3380 43.8590 ;
        RECT 8.4470 43.1390 8.5730 44.0370 ;
        RECT 7.1960 43.0430 8.4200 43.8590 ;
        RECT 0.1760 42.9435 7.1780 44.0370 ;
        RECT 0.0050 42.9435 0.1580 43.8590 ;
        RECT 8.5550 42.9435 16.5290 43.7630 ;
        RECT 0.0050 43.0430 8.5370 43.7630 ;
        RECT 8.3300 42.9435 16.5290 43.1150 ;
        RECT 0.0050 42.9435 8.3120 43.7630 ;
        RECT 0.0050 42.9435 16.5290 43.0190 ;
        RECT 0.0050 44.9870 16.5290 45.1170 ;
        RECT 16.4120 44.0235 16.5290 45.1170 ;
        RECT 9.3020 44.8910 16.3940 45.1170 ;
        RECT 7.9700 44.8910 9.2840 45.1170 ;
        RECT 7.2500 44.0235 7.8800 45.1170 ;
        RECT 0.1400 44.8910 7.2320 45.1170 ;
        RECT 0.0050 44.0235 0.1220 45.1170 ;
        RECT 16.3760 44.0235 16.5290 44.9390 ;
        RECT 9.3560 44.0235 16.3580 45.1170 ;
        RECT 8.6090 44.0235 9.3380 44.9390 ;
        RECT 8.4470 44.2190 8.5730 45.1170 ;
        RECT 7.1960 44.1230 8.4200 44.9390 ;
        RECT 0.1760 44.0235 7.1780 45.1170 ;
        RECT 0.0050 44.0235 0.1580 44.9390 ;
        RECT 8.5550 44.0235 16.5290 44.8430 ;
        RECT 0.0050 44.1230 8.5370 44.8430 ;
        RECT 8.3300 44.0235 16.5290 44.1950 ;
        RECT 0.0050 44.0235 8.3120 44.8430 ;
        RECT 0.0050 44.0235 16.5290 44.0990 ;
        RECT 0.0050 46.0670 16.5290 46.1970 ;
        RECT 16.4120 45.1035 16.5290 46.1970 ;
        RECT 9.3020 45.9710 16.3940 46.1970 ;
        RECT 7.9700 45.9710 9.2840 46.1970 ;
        RECT 7.2500 45.1035 7.8800 46.1970 ;
        RECT 0.1400 45.9710 7.2320 46.1970 ;
        RECT 0.0050 45.1035 0.1220 46.1970 ;
        RECT 16.3760 45.1035 16.5290 46.0190 ;
        RECT 9.3560 45.1035 16.3580 46.1970 ;
        RECT 8.6090 45.1035 9.3380 46.0190 ;
        RECT 8.4470 45.2990 8.5730 46.1970 ;
        RECT 7.1960 45.2030 8.4200 46.0190 ;
        RECT 0.1760 45.1035 7.1780 46.1970 ;
        RECT 0.0050 45.1035 0.1580 46.0190 ;
        RECT 8.5550 45.1035 16.5290 45.9230 ;
        RECT 0.0050 45.2030 8.5370 45.9230 ;
        RECT 8.3300 45.1035 16.5290 45.2750 ;
        RECT 0.0050 45.1035 8.3120 45.9230 ;
        RECT 0.0050 45.1035 16.5290 45.1790 ;
        RECT 0.0050 47.1470 16.5290 47.2770 ;
        RECT 16.4120 46.1835 16.5290 47.2770 ;
        RECT 9.3020 47.0510 16.3940 47.2770 ;
        RECT 7.9700 47.0510 9.2840 47.2770 ;
        RECT 7.2500 46.1835 7.8800 47.2770 ;
        RECT 0.1400 47.0510 7.2320 47.2770 ;
        RECT 0.0050 46.1835 0.1220 47.2770 ;
        RECT 16.3760 46.1835 16.5290 47.0990 ;
        RECT 9.3560 46.1835 16.3580 47.2770 ;
        RECT 8.6090 46.1835 9.3380 47.0990 ;
        RECT 8.4470 46.3790 8.5730 47.2770 ;
        RECT 7.1960 46.2830 8.4200 47.0990 ;
        RECT 0.1760 46.1835 7.1780 47.2770 ;
        RECT 0.0050 46.1835 0.1580 47.0990 ;
        RECT 8.5550 46.1835 16.5290 47.0030 ;
        RECT 0.0050 46.2830 8.5370 47.0030 ;
        RECT 8.3300 46.1835 16.5290 46.3550 ;
        RECT 0.0050 46.1835 8.3120 47.0030 ;
        RECT 0.0050 46.1835 16.5290 46.2590 ;
        RECT 0.0050 48.2270 16.5290 48.3570 ;
        RECT 16.4120 47.2635 16.5290 48.3570 ;
        RECT 9.3020 48.1310 16.3940 48.3570 ;
        RECT 7.9700 48.1310 9.2840 48.3570 ;
        RECT 7.2500 47.2635 7.8800 48.3570 ;
        RECT 0.1400 48.1310 7.2320 48.3570 ;
        RECT 0.0050 47.2635 0.1220 48.3570 ;
        RECT 16.3760 47.2635 16.5290 48.1790 ;
        RECT 9.3560 47.2635 16.3580 48.3570 ;
        RECT 8.6090 47.2635 9.3380 48.1790 ;
        RECT 8.4470 47.4590 8.5730 48.3570 ;
        RECT 7.1960 47.3630 8.4200 48.1790 ;
        RECT 0.1760 47.2635 7.1780 48.3570 ;
        RECT 0.0050 47.2635 0.1580 48.1790 ;
        RECT 8.5550 47.2635 16.5290 48.0830 ;
        RECT 0.0050 47.3630 8.5370 48.0830 ;
        RECT 8.3300 47.2635 16.5290 47.4350 ;
        RECT 0.0050 47.2635 8.3120 48.0830 ;
        RECT 0.0050 47.2635 16.5290 47.3390 ;
        RECT 0.0050 49.3070 16.5290 49.4370 ;
        RECT 16.4120 48.3435 16.5290 49.4370 ;
        RECT 9.3020 49.2110 16.3940 49.4370 ;
        RECT 7.9700 49.2110 9.2840 49.4370 ;
        RECT 7.2500 48.3435 7.8800 49.4370 ;
        RECT 0.1400 49.2110 7.2320 49.4370 ;
        RECT 0.0050 48.3435 0.1220 49.4370 ;
        RECT 16.3760 48.3435 16.5290 49.2590 ;
        RECT 9.3560 48.3435 16.3580 49.4370 ;
        RECT 8.6090 48.3435 9.3380 49.2590 ;
        RECT 8.4470 48.5390 8.5730 49.4370 ;
        RECT 7.1960 48.4430 8.4200 49.2590 ;
        RECT 0.1760 48.3435 7.1780 49.4370 ;
        RECT 0.0050 48.3435 0.1580 49.2590 ;
        RECT 8.5550 48.3435 16.5290 49.1630 ;
        RECT 0.0050 48.4430 8.5370 49.1630 ;
        RECT 8.3300 48.3435 16.5290 48.5150 ;
        RECT 0.0050 48.3435 8.3120 49.1630 ;
        RECT 0.0050 48.3435 16.5290 48.4190 ;
        RECT 0.0050 50.3870 16.5290 50.5170 ;
        RECT 16.4120 49.4235 16.5290 50.5170 ;
        RECT 9.3020 50.2910 16.3940 50.5170 ;
        RECT 7.9700 50.2910 9.2840 50.5170 ;
        RECT 7.2500 49.4235 7.8800 50.5170 ;
        RECT 0.1400 50.2910 7.2320 50.5170 ;
        RECT 0.0050 49.4235 0.1220 50.5170 ;
        RECT 16.3760 49.4235 16.5290 50.3390 ;
        RECT 9.3560 49.4235 16.3580 50.5170 ;
        RECT 8.6090 49.4235 9.3380 50.3390 ;
        RECT 8.4470 49.6190 8.5730 50.5170 ;
        RECT 7.1960 49.5230 8.4200 50.3390 ;
        RECT 0.1760 49.4235 7.1780 50.5170 ;
        RECT 0.0050 49.4235 0.1580 50.3390 ;
        RECT 8.5550 49.4235 16.5290 50.2430 ;
        RECT 0.0050 49.5230 8.5370 50.2430 ;
        RECT 8.3300 49.4235 16.5290 49.5950 ;
        RECT 0.0050 49.4235 8.3120 50.2430 ;
        RECT 0.0050 49.4235 16.5290 49.4990 ;
        RECT 0.0050 51.4670 16.5290 51.5970 ;
        RECT 16.4120 50.5035 16.5290 51.5970 ;
        RECT 9.3020 51.3710 16.3940 51.5970 ;
        RECT 7.9700 51.3710 9.2840 51.5970 ;
        RECT 7.2500 50.5035 7.8800 51.5970 ;
        RECT 0.1400 51.3710 7.2320 51.5970 ;
        RECT 0.0050 50.5035 0.1220 51.5970 ;
        RECT 16.3760 50.5035 16.5290 51.4190 ;
        RECT 9.3560 50.5035 16.3580 51.5970 ;
        RECT 8.6090 50.5035 9.3380 51.4190 ;
        RECT 8.4470 50.6990 8.5730 51.5970 ;
        RECT 7.1960 50.6030 8.4200 51.4190 ;
        RECT 0.1760 50.5035 7.1780 51.5970 ;
        RECT 0.0050 50.5035 0.1580 51.4190 ;
        RECT 8.5550 50.5035 16.5290 51.3230 ;
        RECT 0.0050 50.6030 8.5370 51.3230 ;
        RECT 8.3300 50.5035 16.5290 50.6750 ;
        RECT 0.0050 50.5035 8.3120 51.3230 ;
        RECT 0.0050 50.5035 16.5290 50.5790 ;
        RECT 0.0050 52.5470 16.5290 52.6770 ;
        RECT 16.4120 51.5835 16.5290 52.6770 ;
        RECT 9.3020 52.4510 16.3940 52.6770 ;
        RECT 7.9700 52.4510 9.2840 52.6770 ;
        RECT 7.2500 51.5835 7.8800 52.6770 ;
        RECT 0.1400 52.4510 7.2320 52.6770 ;
        RECT 0.0050 51.5835 0.1220 52.6770 ;
        RECT 16.3760 51.5835 16.5290 52.4990 ;
        RECT 9.3560 51.5835 16.3580 52.6770 ;
        RECT 8.6090 51.5835 9.3380 52.4990 ;
        RECT 8.4470 51.7790 8.5730 52.6770 ;
        RECT 7.1960 51.6830 8.4200 52.4990 ;
        RECT 0.1760 51.5835 7.1780 52.6770 ;
        RECT 0.0050 51.5835 0.1580 52.4990 ;
        RECT 8.5550 51.5835 16.5290 52.4030 ;
        RECT 0.0050 51.6830 8.5370 52.4030 ;
        RECT 8.3300 51.5835 16.5290 51.7550 ;
        RECT 0.0050 51.5835 8.3120 52.4030 ;
        RECT 0.0050 51.5835 16.5290 51.6590 ;
        RECT 0.0050 53.6270 16.5290 53.7570 ;
        RECT 16.4120 52.6635 16.5290 53.7570 ;
        RECT 9.3020 53.5310 16.3940 53.7570 ;
        RECT 7.9700 53.5310 9.2840 53.7570 ;
        RECT 7.2500 52.6635 7.8800 53.7570 ;
        RECT 0.1400 53.5310 7.2320 53.7570 ;
        RECT 0.0050 52.6635 0.1220 53.7570 ;
        RECT 16.3760 52.6635 16.5290 53.5790 ;
        RECT 9.3560 52.6635 16.3580 53.7570 ;
        RECT 8.6090 52.6635 9.3380 53.5790 ;
        RECT 8.4470 52.8590 8.5730 53.7570 ;
        RECT 7.1960 52.7630 8.4200 53.5790 ;
        RECT 0.1760 52.6635 7.1780 53.7570 ;
        RECT 0.0050 52.6635 0.1580 53.5790 ;
        RECT 8.5550 52.6635 16.5290 53.4830 ;
        RECT 0.0050 52.7630 8.5370 53.4830 ;
        RECT 8.3300 52.6635 16.5290 52.8350 ;
        RECT 0.0050 52.6635 8.3120 53.4830 ;
        RECT 0.0050 52.6635 16.5290 52.7390 ;
        RECT 0.0050 54.7070 16.5290 54.8370 ;
        RECT 16.4120 53.7435 16.5290 54.8370 ;
        RECT 9.3020 54.6110 16.3940 54.8370 ;
        RECT 7.9700 54.6110 9.2840 54.8370 ;
        RECT 7.2500 53.7435 7.8800 54.8370 ;
        RECT 0.1400 54.6110 7.2320 54.8370 ;
        RECT 0.0050 53.7435 0.1220 54.8370 ;
        RECT 16.3760 53.7435 16.5290 54.6590 ;
        RECT 9.3560 53.7435 16.3580 54.8370 ;
        RECT 8.6090 53.7435 9.3380 54.6590 ;
        RECT 8.4470 53.9390 8.5730 54.8370 ;
        RECT 7.1960 53.8430 8.4200 54.6590 ;
        RECT 0.1760 53.7435 7.1780 54.8370 ;
        RECT 0.0050 53.7435 0.1580 54.6590 ;
        RECT 8.5550 53.7435 16.5290 54.5630 ;
        RECT 0.0050 53.8430 8.5370 54.5630 ;
        RECT 8.3300 53.7435 16.5290 53.9150 ;
        RECT 0.0050 53.7435 8.3120 54.5630 ;
        RECT 0.0050 53.7435 16.5290 53.8190 ;
        RECT 0.0050 55.7870 16.5290 55.9170 ;
        RECT 16.4120 54.8235 16.5290 55.9170 ;
        RECT 9.3020 55.6910 16.3940 55.9170 ;
        RECT 7.9700 55.6910 9.2840 55.9170 ;
        RECT 7.2500 54.8235 7.8800 55.9170 ;
        RECT 0.1400 55.6910 7.2320 55.9170 ;
        RECT 0.0050 54.8235 0.1220 55.9170 ;
        RECT 16.3760 54.8235 16.5290 55.7390 ;
        RECT 9.3560 54.8235 16.3580 55.9170 ;
        RECT 8.6090 54.8235 9.3380 55.7390 ;
        RECT 8.4470 55.0190 8.5730 55.9170 ;
        RECT 7.1960 54.9230 8.4200 55.7390 ;
        RECT 0.1760 54.8235 7.1780 55.9170 ;
        RECT 0.0050 54.8235 0.1580 55.7390 ;
        RECT 8.5550 54.8235 16.5290 55.6430 ;
        RECT 0.0050 54.9230 8.5370 55.6430 ;
        RECT 8.3300 54.8235 16.5290 54.9950 ;
        RECT 0.0050 54.8235 8.3120 55.6430 ;
        RECT 0.0050 54.8235 16.5290 54.8990 ;
        RECT 0.0050 56.8670 16.5290 56.9970 ;
        RECT 16.4120 55.9035 16.5290 56.9970 ;
        RECT 9.3020 56.7710 16.3940 56.9970 ;
        RECT 7.9700 56.7710 9.2840 56.9970 ;
        RECT 7.2500 55.9035 7.8800 56.9970 ;
        RECT 0.1400 56.7710 7.2320 56.9970 ;
        RECT 0.0050 55.9035 0.1220 56.9970 ;
        RECT 16.3760 55.9035 16.5290 56.8190 ;
        RECT 9.3560 55.9035 16.3580 56.9970 ;
        RECT 8.6090 55.9035 9.3380 56.8190 ;
        RECT 8.4470 56.0990 8.5730 56.9970 ;
        RECT 7.1960 56.0030 8.4200 56.8190 ;
        RECT 0.1760 55.9035 7.1780 56.9970 ;
        RECT 0.0050 55.9035 0.1580 56.8190 ;
        RECT 8.5550 55.9035 16.5290 56.7230 ;
        RECT 0.0050 56.0030 8.5370 56.7230 ;
        RECT 8.3300 55.9035 16.5290 56.0750 ;
        RECT 0.0050 55.9035 8.3120 56.7230 ;
        RECT 0.0050 55.9035 16.5290 55.9790 ;
        RECT 0.0050 57.9470 16.5290 58.0770 ;
        RECT 16.4120 56.9835 16.5290 58.0770 ;
        RECT 9.3020 57.8510 16.3940 58.0770 ;
        RECT 7.9700 57.8510 9.2840 58.0770 ;
        RECT 7.2500 56.9835 7.8800 58.0770 ;
        RECT 0.1400 57.8510 7.2320 58.0770 ;
        RECT 0.0050 56.9835 0.1220 58.0770 ;
        RECT 16.3760 56.9835 16.5290 57.8990 ;
        RECT 9.3560 56.9835 16.3580 58.0770 ;
        RECT 8.6090 56.9835 9.3380 57.8990 ;
        RECT 8.4470 57.1790 8.5730 58.0770 ;
        RECT 7.1960 57.0830 8.4200 57.8990 ;
        RECT 0.1760 56.9835 7.1780 58.0770 ;
        RECT 0.0050 56.9835 0.1580 57.8990 ;
        RECT 8.5550 56.9835 16.5290 57.8030 ;
        RECT 0.0050 57.0830 8.5370 57.8030 ;
        RECT 8.3300 56.9835 16.5290 57.1550 ;
        RECT 0.0050 56.9835 8.3120 57.8030 ;
        RECT 0.0050 56.9835 16.5290 57.0590 ;
        RECT 0.0050 59.0270 16.5290 59.1570 ;
        RECT 16.4120 58.0635 16.5290 59.1570 ;
        RECT 9.3020 58.9310 16.3940 59.1570 ;
        RECT 7.9700 58.9310 9.2840 59.1570 ;
        RECT 7.2500 58.0635 7.8800 59.1570 ;
        RECT 0.1400 58.9310 7.2320 59.1570 ;
        RECT 0.0050 58.0635 0.1220 59.1570 ;
        RECT 16.3760 58.0635 16.5290 58.9790 ;
        RECT 9.3560 58.0635 16.3580 59.1570 ;
        RECT 8.6090 58.0635 9.3380 58.9790 ;
        RECT 8.4470 58.2590 8.5730 59.1570 ;
        RECT 7.1960 58.1630 8.4200 58.9790 ;
        RECT 0.1760 58.0635 7.1780 59.1570 ;
        RECT 0.0050 58.0635 0.1580 58.9790 ;
        RECT 8.5550 58.0635 16.5290 58.8830 ;
        RECT 0.0050 58.1630 8.5370 58.8830 ;
        RECT 8.3300 58.0635 16.5290 58.2350 ;
        RECT 0.0050 58.0635 8.3120 58.8830 ;
        RECT 0.0050 58.0635 16.5290 58.1390 ;
        RECT 0.0050 60.1070 16.5290 60.2370 ;
        RECT 16.4120 59.1435 16.5290 60.2370 ;
        RECT 9.3020 60.0110 16.3940 60.2370 ;
        RECT 7.9700 60.0110 9.2840 60.2370 ;
        RECT 7.2500 59.1435 7.8800 60.2370 ;
        RECT 0.1400 60.0110 7.2320 60.2370 ;
        RECT 0.0050 59.1435 0.1220 60.2370 ;
        RECT 16.3760 59.1435 16.5290 60.0590 ;
        RECT 9.3560 59.1435 16.3580 60.2370 ;
        RECT 8.6090 59.1435 9.3380 60.0590 ;
        RECT 8.4470 59.3390 8.5730 60.2370 ;
        RECT 7.1960 59.2430 8.4200 60.0590 ;
        RECT 0.1760 59.1435 7.1780 60.2370 ;
        RECT 0.0050 59.1435 0.1580 60.0590 ;
        RECT 8.5550 59.1435 16.5290 59.9630 ;
        RECT 0.0050 59.2430 8.5370 59.9630 ;
        RECT 8.3300 59.1435 16.5290 59.3150 ;
        RECT 0.0050 59.1435 8.3120 59.9630 ;
        RECT 0.0050 59.1435 16.5290 59.2190 ;
  LAYER M4  ;
      RECT 1.5690 27.8700 15.0095 27.8940 ;
      RECT 1.5690 28.1580 15.0095 28.1820 ;
      RECT 1.5690 28.5420 15.0095 28.5660 ;
      RECT 1.5690 28.6380 15.0095 28.6620 ;
      RECT 1.5690 28.9740 15.0095 28.9980 ;
      RECT 1.5690 29.3580 15.0095 29.3820 ;
      RECT 10.9550 26.8290 11.0390 26.8530 ;
      RECT 10.7670 27.2610 10.8970 27.2850 ;
      RECT 10.7750 27.9185 10.8920 27.9425 ;
      RECT 10.7750 28.2060 10.8920 28.2300 ;
      RECT 10.1360 27.2610 10.7070 27.2850 ;
      RECT 10.1960 28.0380 10.3040 28.0620 ;
      RECT 8.8630 28.4130 9.9560 28.4370 ;
      RECT 9.5510 27.9810 9.6350 28.0050 ;
      RECT 8.7670 29.1810 9.6350 29.2050 ;
      RECT 9.5510 29.2770 9.6350 29.3010 ;
      RECT 9.3730 27.5010 9.4570 27.5250 ;
      RECT 9.3350 28.8450 9.4190 28.8690 ;
      RECT 9.3350 29.5650 9.4190 29.5890 ;
      RECT 9.1570 27.4050 9.2410 27.4290 ;
      RECT 8.9430 26.1170 9.2060 26.1410 ;
      RECT 8.9430 34.7410 9.2060 34.7650 ;
      RECT 8.9590 28.8930 9.2030 28.9170 ;
      RECT 9.1190 29.0370 9.2030 29.0610 ;
      RECT 7.6630 29.2770 9.2030 29.3010 ;
      RECT 9.1190 29.5650 9.2030 29.5890 ;
      RECT 8.8850 34.6450 9.1480 34.6690 ;
      RECT 8.8840 26.0210 9.1470 26.0450 ;
      RECT 8.8460 25.9250 9.1090 25.9490 ;
      RECT 8.8460 34.4530 9.1090 34.4770 ;
      RECT 9.0110 29.9970 9.0950 30.0210 ;
      RECT 8.2390 30.3810 9.0950 30.4050 ;
      RECT 8.6230 32.6370 9.0950 32.6610 ;
      RECT 9.0110 32.7330 9.0950 32.7570 ;
      RECT 8.7980 25.8290 9.0610 25.8530 ;
      RECT 8.7980 34.3570 9.0610 34.3810 ;
      RECT 8.5750 31.7250 9.0200 31.7490 ;
      RECT 8.7540 25.7330 9.0170 25.7570 ;
      RECT 8.7540 34.6930 9.0170 34.7170 ;
      RECT 8.7050 26.0690 8.9680 26.0930 ;
      RECT 8.7050 34.5970 8.9680 34.6210 ;
      RECT 8.8360 29.0370 8.9570 29.0610 ;
      RECT 8.8150 31.1490 8.9480 31.1730 ;
      RECT 8.6580 25.9730 8.9210 25.9970 ;
      RECT 8.6580 34.5010 8.9210 34.5250 ;
      RECT 8.6230 25.6850 8.8860 25.7090 ;
      RECT 8.6230 34.4050 8.8860 34.4290 ;
      RECT 7.8070 32.7330 8.8760 32.7570 ;
      RECT 8.7920 33.8850 8.8760 33.9090 ;
      RECT 8.5670 25.5410 8.8300 25.5650 ;
      RECT 8.5670 34.3090 8.8300 34.3330 ;
      RECT 8.7190 29.9970 8.8040 30.0210 ;
      RECT 7.6150 30.5730 8.7320 30.5970 ;
      RECT 8.2600 28.4130 8.7170 28.4370 ;
      RECT 8.0870 26.2610 8.3540 26.2850 ;
      RECT 8.0870 34.1650 8.3540 34.1890 ;
      RECT 8.2240 29.9490 8.3330 29.9730 ;
      RECT 8.0640 26.1650 8.3060 26.1890 ;
      RECT 8.0640 34.7890 8.3060 34.8130 ;
      RECT 8.0080 25.6850 8.2500 25.7090 ;
      RECT 8.0370 34.8850 8.2500 34.9090 ;
      RECT 8.1530 29.5650 8.2370 29.5890 ;
      RECT 7.9540 25.7810 8.2020 25.8050 ;
      RECT 7.9540 34.7410 8.2020 34.7650 ;
      RECT 7.7200 32.1570 8.1410 32.1810 ;
      RECT 7.6880 26.1170 7.9550 26.1410 ;
      RECT 7.6880 34.8850 7.9550 34.9090 ;
      RECT 7.8280 30.7170 7.9490 30.7410 ;
      RECT 7.8200 33.8850 7.9040 33.9090 ;
      RECT 7.6540 26.0210 7.9010 26.0450 ;
      RECT 7.5870 34.4530 7.9010 34.4770 ;
      RECT 7.6280 25.9250 7.8580 25.9490 ;
      RECT 7.6160 34.7890 7.8580 34.8130 ;
      RECT 7.5750 25.8290 7.8050 25.8530 ;
      RECT 7.7210 32.3010 7.8050 32.3250 ;
      RECT 7.5250 34.3570 7.8050 34.3810 ;
      RECT 7.5300 25.7330 7.7600 25.7570 ;
      RECT 7.5300 34.6930 7.7600 34.7170 ;
      RECT 6.5680 29.5650 7.7570 29.5890 ;
      RECT 7.4920 25.9730 7.7220 25.9970 ;
      RECT 7.4920 34.5970 7.7220 34.6210 ;
      RECT 7.4740 25.8770 7.6670 25.9010 ;
      RECT 7.4740 34.5010 7.6670 34.5250 ;
      RECT 7.4250 25.7810 7.6180 25.8050 ;
      RECT 7.4250 34.4050 7.6180 34.4290 ;
      RECT 7.4290 30.4770 7.6130 30.5010 ;
      RECT 7.3730 25.6850 7.5660 25.7090 ;
      RECT 7.3730 34.3090 7.5660 34.3330 ;
      RECT 6.8890 27.7890 7.5650 27.8130 ;
      RECT 7.4290 30.5730 7.5130 30.5970 ;
      RECT 7.1600 26.2130 7.4230 26.2370 ;
      RECT 7.1925 29.9970 7.3260 30.0210 ;
      RECT 6.8510 27.9810 6.9350 28.0050 ;
  LAYER V4  ;
      RECT 11.0040 26.8290 11.0280 26.8530 ;
      RECT 11.0040 27.8700 11.0280 27.8940 ;
      RECT 10.8360 27.2610 10.8600 27.2850 ;
      RECT 10.8360 27.9185 10.8600 27.9425 ;
      RECT 10.8360 28.2060 10.8600 28.2300 ;
      RECT 10.2120 27.2610 10.2360 27.2850 ;
      RECT 10.2120 28.0380 10.2360 28.0620 ;
      RECT 9.6000 27.9810 9.6240 28.0050 ;
      RECT 9.6000 28.1580 9.6240 28.1820 ;
      RECT 9.6000 29.1810 9.6240 29.2050 ;
      RECT 9.6000 29.2770 9.6240 29.3010 ;
      RECT 9.3840 27.5010 9.4080 27.5250 ;
      RECT 9.3840 28.5420 9.4080 28.5660 ;
      RECT 9.3840 28.8450 9.4080 28.8690 ;
      RECT 9.3840 28.9740 9.4080 28.9980 ;
      RECT 9.3840 29.3580 9.4080 29.3820 ;
      RECT 9.3840 29.5650 9.4080 29.5890 ;
      RECT 9.1680 27.4050 9.1920 27.4290 ;
      RECT 9.1680 28.6380 9.1920 28.6620 ;
      RECT 9.1680 28.8930 9.1920 28.9170 ;
      RECT 9.1680 29.0370 9.1920 29.0610 ;
      RECT 9.1680 29.2770 9.1920 29.3010 ;
      RECT 9.1680 29.5650 9.1920 29.5890 ;
      RECT 9.0600 29.9970 9.0840 30.0210 ;
      RECT 9.0600 30.3810 9.0840 30.4050 ;
      RECT 9.0600 32.6370 9.0840 32.6610 ;
      RECT 9.0600 32.7330 9.0840 32.7570 ;
      RECT 8.9700 26.1170 8.9940 26.1410 ;
      RECT 8.9700 28.8930 8.9940 28.9170 ;
      RECT 8.9700 34.7410 8.9940 34.7650 ;
      RECT 8.9220 26.0210 8.9460 26.0450 ;
      RECT 8.9220 29.0370 8.9460 29.0610 ;
      RECT 8.9220 34.6450 8.9460 34.6690 ;
      RECT 8.8740 25.9250 8.8980 25.9490 ;
      RECT 8.8740 28.4130 8.8980 28.4370 ;
      RECT 8.8740 34.4530 8.8980 34.4770 ;
      RECT 8.8260 25.8290 8.8500 25.8530 ;
      RECT 8.8260 31.1490 8.8500 31.1730 ;
      RECT 8.8260 33.8850 8.8500 33.9090 ;
      RECT 8.8260 34.3570 8.8500 34.3810 ;
      RECT 8.7780 25.7330 8.8020 25.7570 ;
      RECT 8.7780 29.1810 8.8020 29.2050 ;
      RECT 8.7780 34.6930 8.8020 34.7170 ;
      RECT 8.7300 26.0690 8.7540 26.0930 ;
      RECT 8.7300 29.9970 8.7540 30.0210 ;
      RECT 8.7300 34.5970 8.7540 34.6210 ;
      RECT 8.6820 25.9730 8.7060 25.9970 ;
      RECT 8.6820 28.4130 8.7060 28.4370 ;
      RECT 8.6820 34.5010 8.7060 34.5250 ;
      RECT 8.6340 25.6850 8.6580 25.7090 ;
      RECT 8.6340 32.6370 8.6580 32.6610 ;
      RECT 8.6340 34.4050 8.6580 34.4290 ;
      RECT 8.5860 25.5410 8.6100 25.5650 ;
      RECT 8.5860 31.7250 8.6100 31.7490 ;
      RECT 8.5860 34.3090 8.6100 34.3330 ;
      RECT 8.2980 26.2610 8.3220 26.2850 ;
      RECT 8.2980 29.9490 8.3220 29.9730 ;
      RECT 8.2980 34.1650 8.3220 34.1890 ;
      RECT 8.2500 26.1650 8.2740 26.1890 ;
      RECT 8.2500 30.3810 8.2740 30.4050 ;
      RECT 8.2500 34.7890 8.2740 34.8130 ;
      RECT 8.2020 25.6850 8.2260 25.7090 ;
      RECT 8.2020 29.5650 8.2260 29.5890 ;
      RECT 8.2020 34.8850 8.2260 34.9090 ;
      RECT 8.1060 25.7810 8.1300 25.8050 ;
      RECT 8.1060 32.1570 8.1300 32.1810 ;
      RECT 8.1060 34.7410 8.1300 34.7650 ;
      RECT 7.9140 26.1170 7.9380 26.1410 ;
      RECT 7.9140 30.7170 7.9380 30.7410 ;
      RECT 7.9140 34.8850 7.9380 34.9090 ;
      RECT 7.8660 26.0210 7.8900 26.0450 ;
      RECT 7.8660 33.8850 7.8900 33.9090 ;
      RECT 7.8660 34.4530 7.8900 34.4770 ;
      RECT 7.8180 25.9250 7.8420 25.9490 ;
      RECT 7.8180 32.7330 7.8420 32.7570 ;
      RECT 7.8180 34.7890 7.8420 34.8130 ;
      RECT 7.7700 25.8290 7.7940 25.8530 ;
      RECT 7.7700 32.3010 7.7940 32.3250 ;
      RECT 7.7700 34.3570 7.7940 34.3810 ;
      RECT 7.7220 25.7330 7.7460 25.7570 ;
      RECT 7.7220 29.5650 7.7460 29.5890 ;
      RECT 7.7220 34.6930 7.7460 34.7170 ;
      RECT 7.6740 25.9730 7.6980 25.9970 ;
      RECT 7.6740 29.2770 7.6980 29.3010 ;
      RECT 7.6740 34.5970 7.6980 34.6210 ;
      RECT 7.6260 25.8770 7.6500 25.9010 ;
      RECT 7.6260 30.5730 7.6500 30.5970 ;
      RECT 7.6260 34.5010 7.6500 34.5250 ;
      RECT 7.5780 25.7810 7.6020 25.8050 ;
      RECT 7.5780 30.4770 7.6020 30.5010 ;
      RECT 7.5780 34.4050 7.6020 34.4290 ;
      RECT 7.5300 25.6850 7.5540 25.7090 ;
      RECT 7.5300 27.7890 7.5540 27.8130 ;
      RECT 7.5300 34.3090 7.5540 34.3330 ;
      RECT 7.4400 30.4770 7.4640 30.5010 ;
      RECT 7.4400 30.5730 7.4640 30.5970 ;
      RECT 7.2720 26.2130 7.2960 26.2370 ;
      RECT 7.2720 29.9970 7.2960 30.0210 ;
      RECT 6.9000 27.7890 6.9240 27.8130 ;
      RECT 6.9000 27.9810 6.9240 28.0050 ;
  LAYER M5  ;
      RECT 11.0040 26.8180 11.0280 27.9050 ;
      RECT 10.8360 27.2330 10.8600 28.2935 ;
      RECT 10.2120 27.2415 10.2360 28.0740 ;
      RECT 9.6000 27.9700 9.6240 28.1930 ;
      RECT 9.6000 29.1700 9.6240 29.3120 ;
      RECT 9.3840 27.4900 9.4080 28.5770 ;
      RECT 9.3840 28.8340 9.4080 29.0090 ;
      RECT 9.3840 29.3470 9.4080 29.6000 ;
      RECT 9.1680 27.3940 9.1920 28.6730 ;
      RECT 9.1680 28.8820 9.1920 29.0720 ;
      RECT 9.1680 29.2660 9.1920 29.6000 ;
      RECT 9.0600 29.9860 9.0840 30.4160 ;
      RECT 9.0600 32.6260 9.0840 32.7680 ;
      RECT 8.9700 26.4540 8.9940 34.0370 ;
      RECT 8.9220 26.4540 8.9460 34.0370 ;
      RECT 8.8740 26.4540 8.8980 34.0370 ;
      RECT 8.8260 26.4540 8.8500 34.0370 ;
      RECT 8.7780 26.4540 8.8020 34.0370 ;
      RECT 8.7300 26.4540 8.7540 34.0370 ;
      RECT 8.6820 26.4540 8.7060 34.0370 ;
      RECT 8.6340 26.4540 8.6580 34.0370 ;
      RECT 8.5860 26.4540 8.6100 34.0370 ;
      RECT 8.2980 26.4540 8.3220 34.0370 ;
      RECT 8.2500 26.4540 8.2740 34.0370 ;
      RECT 8.2020 26.4540 8.2260 34.0370 ;
      RECT 8.1060 26.4540 8.1300 34.0370 ;
      RECT 7.9140 26.4540 7.9380 34.0370 ;
      RECT 7.8660 26.4540 7.8900 34.0370 ;
      RECT 7.8180 26.4540 7.8420 34.0370 ;
      RECT 7.7700 26.4540 7.7940 34.0370 ;
      RECT 7.7220 26.4540 7.7460 34.0370 ;
      RECT 7.6740 26.4540 7.6980 34.0370 ;
      RECT 7.6260 25.6120 7.6500 34.6670 ;
      RECT 7.5780 25.5750 7.6020 34.6210 ;
      RECT 7.5300 25.5210 7.5540 34.5670 ;
      RECT 7.4400 30.4660 7.4640 30.6080 ;
      RECT 7.2720 26.1950 7.2960 30.0390 ;
      RECT 6.9000 27.7780 6.9240 28.0160 ;
  LAYER M2  ;
    RECT 0.108 0.036 15.8920 60.4440 ;
  LAYER M1  ;
    RECT 0.108 0.036 15.8920 60.4440 ;
  END
END srambank_128x4x48_6t122 
