VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


PROPERTYDEFINITIONS 
  MACRO CatenaDesignType STRING ; 
END PROPERTYDEFINITIONS 


MACRO srambank_256x4x18_6t122 
  CLASS BLOCK ; 
  ORIGIN 0 0 ; 
  FOREIGN srambank_256x4x18_6t122 0 0 ; 
  SIZE 121.392 BY 112.32 ; 
  SYMMETRY X Y ; 
  SITE coreSite ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.416 4.688 121.032 4.88 ; 
        RECT 0.416 9.008 121.032 9.2 ; 
        RECT 0.416 13.328 121.032 13.52 ; 
        RECT 0.416 17.648 121.032 17.84 ; 
        RECT 0.416 21.968 121.032 22.16 ; 
        RECT 0.416 26.288 121.032 26.48 ; 
        RECT 0.416 30.608 121.032 30.8 ; 
        RECT 0.416 34.928 121.032 35.12 ; 
        RECT 0.416 39.248 121.032 39.44 ; 
        RECT 0.416 76.076 121.032 76.268 ; 
        RECT 0.416 80.396 121.032 80.588 ; 
        RECT 0.416 84.716 121.032 84.908 ; 
        RECT 0.416 89.036 121.032 89.228 ; 
        RECT 0.416 93.356 121.032 93.548 ; 
        RECT 0.416 97.676 121.032 97.868 ; 
        RECT 0.416 101.996 121.032 102.188 ; 
        RECT 0.416 106.316 121.032 106.508 ; 
        RECT 0.416 110.636 121.032 110.828 ; 
      LAYER M3 ; 
        RECT 120.872 0.866 120.944 5.506 ; 
        RECT 64.784 0.868 64.856 5.504 ; 
        RECT 59.168 1.012 59.528 5.474 ; 
        RECT 56.576 0.868 56.648 5.504 ; 
        RECT 0.488 0.866 0.56 5.506 ; 
        RECT 120.872 5.186 120.944 9.826 ; 
        RECT 64.784 5.188 64.856 9.824 ; 
        RECT 59.168 5.332 59.528 9.794 ; 
        RECT 56.576 5.188 56.648 9.824 ; 
        RECT 0.488 5.186 0.56 9.826 ; 
        RECT 120.872 9.506 120.944 14.146 ; 
        RECT 64.784 9.508 64.856 14.144 ; 
        RECT 59.168 9.652 59.528 14.114 ; 
        RECT 56.576 9.508 56.648 14.144 ; 
        RECT 0.488 9.506 0.56 14.146 ; 
        RECT 120.872 13.826 120.944 18.466 ; 
        RECT 64.784 13.828 64.856 18.464 ; 
        RECT 59.168 13.972 59.528 18.434 ; 
        RECT 56.576 13.828 56.648 18.464 ; 
        RECT 0.488 13.826 0.56 18.466 ; 
        RECT 120.872 18.146 120.944 22.786 ; 
        RECT 64.784 18.148 64.856 22.784 ; 
        RECT 59.168 18.292 59.528 22.754 ; 
        RECT 56.576 18.148 56.648 22.784 ; 
        RECT 0.488 18.146 0.56 22.786 ; 
        RECT 120.872 22.466 120.944 27.106 ; 
        RECT 64.784 22.468 64.856 27.104 ; 
        RECT 59.168 22.612 59.528 27.074 ; 
        RECT 56.576 22.468 56.648 27.104 ; 
        RECT 0.488 22.466 0.56 27.106 ; 
        RECT 120.872 26.786 120.944 31.426 ; 
        RECT 64.784 26.788 64.856 31.424 ; 
        RECT 59.168 26.932 59.528 31.394 ; 
        RECT 56.576 26.788 56.648 31.424 ; 
        RECT 0.488 26.786 0.56 31.426 ; 
        RECT 120.872 31.106 120.944 35.746 ; 
        RECT 64.784 31.108 64.856 35.744 ; 
        RECT 59.168 31.252 59.528 35.714 ; 
        RECT 56.576 31.108 56.648 35.744 ; 
        RECT 0.488 31.106 0.56 35.746 ; 
        RECT 120.872 35.426 120.944 40.066 ; 
        RECT 64.784 35.428 64.856 40.064 ; 
        RECT 59.168 35.572 59.528 40.034 ; 
        RECT 56.576 35.428 56.648 40.064 ; 
        RECT 0.488 35.426 0.56 40.066 ; 
        RECT 56.196 55.22 56.268 79.474 ; 
        RECT 120.872 72.254 120.944 76.894 ; 
        RECT 64.784 72.256 64.856 76.892 ; 
        RECT 59.168 72.4 59.528 76.862 ; 
        RECT 56.576 72.256 56.648 76.892 ; 
        RECT 0.488 72.254 0.56 76.894 ; 
        RECT 120.872 76.574 120.944 81.214 ; 
        RECT 64.784 76.576 64.856 81.212 ; 
        RECT 59.168 76.72 59.528 81.182 ; 
        RECT 56.576 76.576 56.648 81.212 ; 
        RECT 0.488 76.574 0.56 81.214 ; 
        RECT 120.872 80.894 120.944 85.534 ; 
        RECT 64.784 80.896 64.856 85.532 ; 
        RECT 59.168 81.04 59.528 85.502 ; 
        RECT 56.576 80.896 56.648 85.532 ; 
        RECT 0.488 80.894 0.56 85.534 ; 
        RECT 120.872 85.214 120.944 89.854 ; 
        RECT 64.784 85.216 64.856 89.852 ; 
        RECT 59.168 85.36 59.528 89.822 ; 
        RECT 56.576 85.216 56.648 89.852 ; 
        RECT 0.488 85.214 0.56 89.854 ; 
        RECT 120.872 89.534 120.944 94.174 ; 
        RECT 64.784 89.536 64.856 94.172 ; 
        RECT 59.168 89.68 59.528 94.142 ; 
        RECT 56.576 89.536 56.648 94.172 ; 
        RECT 0.488 89.534 0.56 94.174 ; 
        RECT 120.872 93.854 120.944 98.494 ; 
        RECT 64.784 93.856 64.856 98.492 ; 
        RECT 59.168 94 59.528 98.462 ; 
        RECT 56.576 93.856 56.648 98.492 ; 
        RECT 0.488 93.854 0.56 98.494 ; 
        RECT 120.872 98.174 120.944 102.814 ; 
        RECT 64.784 98.176 64.856 102.812 ; 
        RECT 59.168 98.32 59.528 102.782 ; 
        RECT 56.576 98.176 56.648 102.812 ; 
        RECT 0.488 98.174 0.56 102.814 ; 
        RECT 120.872 102.494 120.944 107.134 ; 
        RECT 64.784 102.496 64.856 107.132 ; 
        RECT 59.168 102.64 59.528 107.102 ; 
        RECT 56.576 102.496 56.648 107.132 ; 
        RECT 0.488 102.494 0.56 107.134 ; 
        RECT 120.872 106.814 120.944 111.454 ; 
        RECT 64.784 106.816 64.856 111.452 ; 
        RECT 59.168 106.96 59.528 111.422 ; 
        RECT 56.576 106.816 56.648 111.452 ; 
        RECT 0.488 106.814 0.56 111.454 ; 
      LAYER V3 ; 
        RECT 0.488 4.688 0.56 4.88 ; 
        RECT 56.576 4.688 56.648 4.88 ; 
        RECT 59.168 4.688 59.528 4.88 ; 
        RECT 64.784 4.688 64.856 4.88 ; 
        RECT 120.872 4.688 120.944 4.88 ; 
        RECT 0.488 9.008 0.56 9.2 ; 
        RECT 56.576 9.008 56.648 9.2 ; 
        RECT 59.168 9.008 59.528 9.2 ; 
        RECT 64.784 9.008 64.856 9.2 ; 
        RECT 120.872 9.008 120.944 9.2 ; 
        RECT 0.488 13.328 0.56 13.52 ; 
        RECT 56.576 13.328 56.648 13.52 ; 
        RECT 59.168 13.328 59.528 13.52 ; 
        RECT 64.784 13.328 64.856 13.52 ; 
        RECT 120.872 13.328 120.944 13.52 ; 
        RECT 0.488 17.648 0.56 17.84 ; 
        RECT 56.576 17.648 56.648 17.84 ; 
        RECT 59.168 17.648 59.528 17.84 ; 
        RECT 64.784 17.648 64.856 17.84 ; 
        RECT 120.872 17.648 120.944 17.84 ; 
        RECT 0.488 21.968 0.56 22.16 ; 
        RECT 56.576 21.968 56.648 22.16 ; 
        RECT 59.168 21.968 59.528 22.16 ; 
        RECT 64.784 21.968 64.856 22.16 ; 
        RECT 120.872 21.968 120.944 22.16 ; 
        RECT 0.488 26.288 0.56 26.48 ; 
        RECT 56.576 26.288 56.648 26.48 ; 
        RECT 59.168 26.288 59.528 26.48 ; 
        RECT 64.784 26.288 64.856 26.48 ; 
        RECT 120.872 26.288 120.944 26.48 ; 
        RECT 0.488 30.608 0.56 30.8 ; 
        RECT 56.576 30.608 56.648 30.8 ; 
        RECT 59.168 30.608 59.528 30.8 ; 
        RECT 64.784 30.608 64.856 30.8 ; 
        RECT 120.872 30.608 120.944 30.8 ; 
        RECT 0.488 34.928 0.56 35.12 ; 
        RECT 56.576 34.928 56.648 35.12 ; 
        RECT 59.168 34.928 59.528 35.12 ; 
        RECT 64.784 34.928 64.856 35.12 ; 
        RECT 120.872 34.928 120.944 35.12 ; 
        RECT 0.488 39.248 0.56 39.44 ; 
        RECT 56.576 39.248 56.648 39.44 ; 
        RECT 59.168 39.248 59.528 39.44 ; 
        RECT 64.784 39.248 64.856 39.44 ; 
        RECT 120.872 39.248 120.944 39.44 ; 
        RECT 0.488 76.076 0.56 76.268 ; 
        RECT 56.576 76.076 56.648 76.268 ; 
        RECT 59.168 76.076 59.528 76.268 ; 
        RECT 64.784 76.076 64.856 76.268 ; 
        RECT 120.872 76.076 120.944 76.268 ; 
        RECT 0.488 80.396 0.56 80.588 ; 
        RECT 56.576 80.396 56.648 80.588 ; 
        RECT 59.168 80.396 59.528 80.588 ; 
        RECT 64.784 80.396 64.856 80.588 ; 
        RECT 120.872 80.396 120.944 80.588 ; 
        RECT 0.488 84.716 0.56 84.908 ; 
        RECT 56.576 84.716 56.648 84.908 ; 
        RECT 59.168 84.716 59.528 84.908 ; 
        RECT 64.784 84.716 64.856 84.908 ; 
        RECT 120.872 84.716 120.944 84.908 ; 
        RECT 0.488 89.036 0.56 89.228 ; 
        RECT 56.576 89.036 56.648 89.228 ; 
        RECT 59.168 89.036 59.528 89.228 ; 
        RECT 64.784 89.036 64.856 89.228 ; 
        RECT 120.872 89.036 120.944 89.228 ; 
        RECT 0.488 93.356 0.56 93.548 ; 
        RECT 56.576 93.356 56.648 93.548 ; 
        RECT 59.168 93.356 59.528 93.548 ; 
        RECT 64.784 93.356 64.856 93.548 ; 
        RECT 120.872 93.356 120.944 93.548 ; 
        RECT 0.488 97.676 0.56 97.868 ; 
        RECT 56.576 97.676 56.648 97.868 ; 
        RECT 59.168 97.676 59.528 97.868 ; 
        RECT 64.784 97.676 64.856 97.868 ; 
        RECT 120.872 97.676 120.944 97.868 ; 
        RECT 0.488 101.996 0.56 102.188 ; 
        RECT 56.576 101.996 56.648 102.188 ; 
        RECT 59.168 101.996 59.528 102.188 ; 
        RECT 64.784 101.996 64.856 102.188 ; 
        RECT 120.872 101.996 120.944 102.188 ; 
        RECT 0.488 106.316 0.56 106.508 ; 
        RECT 56.576 106.316 56.648 106.508 ; 
        RECT 59.168 106.316 59.528 106.508 ; 
        RECT 64.784 106.316 64.856 106.508 ; 
        RECT 120.872 106.316 120.944 106.508 ; 
        RECT 0.488 110.636 0.56 110.828 ; 
        RECT 56.576 110.636 56.648 110.828 ; 
        RECT 59.168 110.636 59.528 110.828 ; 
        RECT 64.784 110.636 64.856 110.828 ; 
        RECT 120.872 110.636 120.944 110.828 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE POWER ; 
    PORT 
      LAYER M4 ; 
        RECT 0.416 4.304 121.032 4.496 ; 
        RECT 0.416 8.624 121.032 8.816 ; 
        RECT 0.416 12.944 121.032 13.136 ; 
        RECT 0.416 17.264 121.032 17.456 ; 
        RECT 0.416 21.584 121.032 21.776 ; 
        RECT 0.416 25.904 121.032 26.096 ; 
        RECT 0.416 30.224 121.032 30.416 ; 
        RECT 0.416 34.544 121.032 34.736 ; 
        RECT 0.416 38.864 121.032 39.056 ; 
        RECT 41.904 43.126 79.488 43.99 ; 
        RECT 57.24 55.798 64.152 56.662 ; 
        RECT 57.24 68.47 64.152 69.334 ; 
        RECT 0.416 75.692 121.032 75.884 ; 
        RECT 0.416 80.012 121.032 80.204 ; 
        RECT 0.416 84.332 121.032 84.524 ; 
        RECT 0.416 88.652 121.032 88.844 ; 
        RECT 0.416 92.972 121.032 93.164 ; 
        RECT 0.416 97.292 121.032 97.484 ; 
        RECT 0.416 101.612 121.032 101.804 ; 
        RECT 0.416 105.932 121.032 106.124 ; 
        RECT 0.416 110.252 121.032 110.444 ; 
      LAYER M3 ; 
        RECT 120.728 0.866 120.8 5.506 ; 
        RECT 65 0.866 65.072 5.506 ; 
        RECT 61.94 1.012 62.084 5.47 ; 
        RECT 61.04 1.012 61.148 5.47 ; 
        RECT 56.36 0.866 56.432 5.506 ; 
        RECT 0.632 0.866 0.704 5.506 ; 
        RECT 120.728 5.186 120.8 9.826 ; 
        RECT 65 5.186 65.072 9.826 ; 
        RECT 61.94 5.332 62.084 9.79 ; 
        RECT 61.04 5.332 61.148 9.79 ; 
        RECT 56.36 5.186 56.432 9.826 ; 
        RECT 0.632 5.186 0.704 9.826 ; 
        RECT 120.728 9.506 120.8 14.146 ; 
        RECT 65 9.506 65.072 14.146 ; 
        RECT 61.94 9.652 62.084 14.11 ; 
        RECT 61.04 9.652 61.148 14.11 ; 
        RECT 56.36 9.506 56.432 14.146 ; 
        RECT 0.632 9.506 0.704 14.146 ; 
        RECT 120.728 13.826 120.8 18.466 ; 
        RECT 65 13.826 65.072 18.466 ; 
        RECT 61.94 13.972 62.084 18.43 ; 
        RECT 61.04 13.972 61.148 18.43 ; 
        RECT 56.36 13.826 56.432 18.466 ; 
        RECT 0.632 13.826 0.704 18.466 ; 
        RECT 120.728 18.146 120.8 22.786 ; 
        RECT 65 18.146 65.072 22.786 ; 
        RECT 61.94 18.292 62.084 22.75 ; 
        RECT 61.04 18.292 61.148 22.75 ; 
        RECT 56.36 18.146 56.432 22.786 ; 
        RECT 0.632 18.146 0.704 22.786 ; 
        RECT 120.728 22.466 120.8 27.106 ; 
        RECT 65 22.466 65.072 27.106 ; 
        RECT 61.94 22.612 62.084 27.07 ; 
        RECT 61.04 22.612 61.148 27.07 ; 
        RECT 56.36 22.466 56.432 27.106 ; 
        RECT 0.632 22.466 0.704 27.106 ; 
        RECT 120.728 26.786 120.8 31.426 ; 
        RECT 65 26.786 65.072 31.426 ; 
        RECT 61.94 26.932 62.084 31.39 ; 
        RECT 61.04 26.932 61.148 31.39 ; 
        RECT 56.36 26.786 56.432 31.426 ; 
        RECT 0.632 26.786 0.704 31.426 ; 
        RECT 120.728 31.106 120.8 35.746 ; 
        RECT 65 31.106 65.072 35.746 ; 
        RECT 61.94 31.252 62.084 35.71 ; 
        RECT 61.04 31.252 61.148 35.71 ; 
        RECT 56.36 31.106 56.432 35.746 ; 
        RECT 0.632 31.106 0.704 35.746 ; 
        RECT 120.728 35.426 120.8 40.066 ; 
        RECT 65 35.426 65.072 40.066 ; 
        RECT 61.94 35.572 62.084 40.03 ; 
        RECT 61.04 35.572 61.148 40.03 ; 
        RECT 56.36 35.426 56.432 40.066 ; 
        RECT 0.632 35.426 0.704 40.066 ; 
        RECT 64.98 39.948 65.052 72.776 ; 
        RECT 61.164 40.842 62.1 71.574 ; 
        RECT 56.34 39.948 56.412 79.474 ; 
        RECT 120.728 72.254 120.8 76.894 ; 
        RECT 65 72.254 65.072 76.894 ; 
        RECT 61.94 72.4 62.084 76.858 ; 
        RECT 61.04 72.4 61.148 76.858 ; 
        RECT 56.36 72.254 56.432 76.894 ; 
        RECT 0.632 72.254 0.704 76.894 ; 
        RECT 120.728 76.574 120.8 81.214 ; 
        RECT 65 76.574 65.072 81.214 ; 
        RECT 61.94 76.72 62.084 81.178 ; 
        RECT 61.04 76.72 61.148 81.178 ; 
        RECT 56.36 76.574 56.432 81.214 ; 
        RECT 0.632 76.574 0.704 81.214 ; 
        RECT 120.728 80.894 120.8 85.534 ; 
        RECT 65 80.894 65.072 85.534 ; 
        RECT 61.94 81.04 62.084 85.498 ; 
        RECT 61.04 81.04 61.148 85.498 ; 
        RECT 56.36 80.894 56.432 85.534 ; 
        RECT 0.632 80.894 0.704 85.534 ; 
        RECT 120.728 85.214 120.8 89.854 ; 
        RECT 65 85.214 65.072 89.854 ; 
        RECT 61.94 85.36 62.084 89.818 ; 
        RECT 61.04 85.36 61.148 89.818 ; 
        RECT 56.36 85.214 56.432 89.854 ; 
        RECT 0.632 85.214 0.704 89.854 ; 
        RECT 120.728 89.534 120.8 94.174 ; 
        RECT 65 89.534 65.072 94.174 ; 
        RECT 61.94 89.68 62.084 94.138 ; 
        RECT 61.04 89.68 61.148 94.138 ; 
        RECT 56.36 89.534 56.432 94.174 ; 
        RECT 0.632 89.534 0.704 94.174 ; 
        RECT 120.728 93.854 120.8 98.494 ; 
        RECT 65 93.854 65.072 98.494 ; 
        RECT 61.94 94 62.084 98.458 ; 
        RECT 61.04 94 61.148 98.458 ; 
        RECT 56.36 93.854 56.432 98.494 ; 
        RECT 0.632 93.854 0.704 98.494 ; 
        RECT 120.728 98.174 120.8 102.814 ; 
        RECT 65 98.174 65.072 102.814 ; 
        RECT 61.94 98.32 62.084 102.778 ; 
        RECT 61.04 98.32 61.148 102.778 ; 
        RECT 56.36 98.174 56.432 102.814 ; 
        RECT 0.632 98.174 0.704 102.814 ; 
        RECT 120.728 102.494 120.8 107.134 ; 
        RECT 65 102.494 65.072 107.134 ; 
        RECT 61.94 102.64 62.084 107.098 ; 
        RECT 61.04 102.64 61.148 107.098 ; 
        RECT 56.36 102.494 56.432 107.134 ; 
        RECT 0.632 102.494 0.704 107.134 ; 
        RECT 120.728 106.814 120.8 111.454 ; 
        RECT 65 106.814 65.072 111.454 ; 
        RECT 61.94 106.96 62.084 111.418 ; 
        RECT 61.04 106.96 61.148 111.418 ; 
        RECT 56.36 106.814 56.432 111.454 ; 
        RECT 0.632 106.814 0.704 111.454 ; 
      LAYER V3 ; 
        RECT 0.632 4.304 0.704 4.496 ; 
        RECT 56.36 4.304 56.432 4.496 ; 
        RECT 61.04 4.304 61.148 4.496 ; 
        RECT 61.94 4.304 62.084 4.496 ; 
        RECT 65 4.304 65.072 4.496 ; 
        RECT 120.728 4.304 120.8 4.496 ; 
        RECT 0.632 8.624 0.704 8.816 ; 
        RECT 56.36 8.624 56.432 8.816 ; 
        RECT 61.04 8.624 61.148 8.816 ; 
        RECT 61.94 8.624 62.084 8.816 ; 
        RECT 65 8.624 65.072 8.816 ; 
        RECT 120.728 8.624 120.8 8.816 ; 
        RECT 0.632 12.944 0.704 13.136 ; 
        RECT 56.36 12.944 56.432 13.136 ; 
        RECT 61.04 12.944 61.148 13.136 ; 
        RECT 61.94 12.944 62.084 13.136 ; 
        RECT 65 12.944 65.072 13.136 ; 
        RECT 120.728 12.944 120.8 13.136 ; 
        RECT 0.632 17.264 0.704 17.456 ; 
        RECT 56.36 17.264 56.432 17.456 ; 
        RECT 61.04 17.264 61.148 17.456 ; 
        RECT 61.94 17.264 62.084 17.456 ; 
        RECT 65 17.264 65.072 17.456 ; 
        RECT 120.728 17.264 120.8 17.456 ; 
        RECT 0.632 21.584 0.704 21.776 ; 
        RECT 56.36 21.584 56.432 21.776 ; 
        RECT 61.04 21.584 61.148 21.776 ; 
        RECT 61.94 21.584 62.084 21.776 ; 
        RECT 65 21.584 65.072 21.776 ; 
        RECT 120.728 21.584 120.8 21.776 ; 
        RECT 0.632 25.904 0.704 26.096 ; 
        RECT 56.36 25.904 56.432 26.096 ; 
        RECT 61.04 25.904 61.148 26.096 ; 
        RECT 61.94 25.904 62.084 26.096 ; 
        RECT 65 25.904 65.072 26.096 ; 
        RECT 120.728 25.904 120.8 26.096 ; 
        RECT 0.632 30.224 0.704 30.416 ; 
        RECT 56.36 30.224 56.432 30.416 ; 
        RECT 61.04 30.224 61.148 30.416 ; 
        RECT 61.94 30.224 62.084 30.416 ; 
        RECT 65 30.224 65.072 30.416 ; 
        RECT 120.728 30.224 120.8 30.416 ; 
        RECT 0.632 34.544 0.704 34.736 ; 
        RECT 56.36 34.544 56.432 34.736 ; 
        RECT 61.04 34.544 61.148 34.736 ; 
        RECT 61.94 34.544 62.084 34.736 ; 
        RECT 65 34.544 65.072 34.736 ; 
        RECT 120.728 34.544 120.8 34.736 ; 
        RECT 0.632 38.864 0.704 39.056 ; 
        RECT 56.36 38.864 56.432 39.056 ; 
        RECT 61.04 38.864 61.148 39.056 ; 
        RECT 61.94 38.864 62.084 39.056 ; 
        RECT 65 38.864 65.072 39.056 ; 
        RECT 120.728 38.864 120.8 39.056 ; 
        RECT 56.34 43.126 56.412 43.99 ; 
        RECT 61.18 68.47 61.252 69.334 ; 
        RECT 61.18 55.798 61.252 56.662 ; 
        RECT 61.18 43.126 61.252 43.99 ; 
        RECT 61.388 68.47 61.46 69.334 ; 
        RECT 61.388 55.798 61.46 56.662 ; 
        RECT 61.388 43.126 61.46 43.99 ; 
        RECT 61.596 68.47 61.668 69.334 ; 
        RECT 61.596 55.798 61.668 56.662 ; 
        RECT 61.596 43.126 61.668 43.99 ; 
        RECT 61.804 68.47 61.876 69.334 ; 
        RECT 61.804 55.798 61.876 56.662 ; 
        RECT 61.804 43.126 61.876 43.99 ; 
        RECT 62.012 68.47 62.084 69.334 ; 
        RECT 62.012 55.798 62.084 56.662 ; 
        RECT 62.012 43.126 62.084 43.99 ; 
        RECT 64.98 43.126 65.052 43.99 ; 
        RECT 0.632 75.692 0.704 75.884 ; 
        RECT 56.36 75.692 56.432 75.884 ; 
        RECT 61.04 75.692 61.148 75.884 ; 
        RECT 61.94 75.692 62.084 75.884 ; 
        RECT 65 75.692 65.072 75.884 ; 
        RECT 120.728 75.692 120.8 75.884 ; 
        RECT 0.632 80.012 0.704 80.204 ; 
        RECT 56.36 80.012 56.432 80.204 ; 
        RECT 61.04 80.012 61.148 80.204 ; 
        RECT 61.94 80.012 62.084 80.204 ; 
        RECT 65 80.012 65.072 80.204 ; 
        RECT 120.728 80.012 120.8 80.204 ; 
        RECT 0.632 84.332 0.704 84.524 ; 
        RECT 56.36 84.332 56.432 84.524 ; 
        RECT 61.04 84.332 61.148 84.524 ; 
        RECT 61.94 84.332 62.084 84.524 ; 
        RECT 65 84.332 65.072 84.524 ; 
        RECT 120.728 84.332 120.8 84.524 ; 
        RECT 0.632 88.652 0.704 88.844 ; 
        RECT 56.36 88.652 56.432 88.844 ; 
        RECT 61.04 88.652 61.148 88.844 ; 
        RECT 61.94 88.652 62.084 88.844 ; 
        RECT 65 88.652 65.072 88.844 ; 
        RECT 120.728 88.652 120.8 88.844 ; 
        RECT 0.632 92.972 0.704 93.164 ; 
        RECT 56.36 92.972 56.432 93.164 ; 
        RECT 61.04 92.972 61.148 93.164 ; 
        RECT 61.94 92.972 62.084 93.164 ; 
        RECT 65 92.972 65.072 93.164 ; 
        RECT 120.728 92.972 120.8 93.164 ; 
        RECT 0.632 97.292 0.704 97.484 ; 
        RECT 56.36 97.292 56.432 97.484 ; 
        RECT 61.04 97.292 61.148 97.484 ; 
        RECT 61.94 97.292 62.084 97.484 ; 
        RECT 65 97.292 65.072 97.484 ; 
        RECT 120.728 97.292 120.8 97.484 ; 
        RECT 0.632 101.612 0.704 101.804 ; 
        RECT 56.36 101.612 56.432 101.804 ; 
        RECT 61.04 101.612 61.148 101.804 ; 
        RECT 61.94 101.612 62.084 101.804 ; 
        RECT 65 101.612 65.072 101.804 ; 
        RECT 120.728 101.612 120.8 101.804 ; 
        RECT 0.632 105.932 0.704 106.124 ; 
        RECT 56.36 105.932 56.432 106.124 ; 
        RECT 61.04 105.932 61.148 106.124 ; 
        RECT 61.94 105.932 62.084 106.124 ; 
        RECT 65 105.932 65.072 106.124 ; 
        RECT 120.728 105.932 120.8 106.124 ; 
        RECT 0.632 110.252 0.704 110.444 ; 
        RECT 56.36 110.252 56.432 110.444 ; 
        RECT 61.04 110.252 61.148 110.444 ; 
        RECT 61.94 110.252 62.084 110.444 ; 
        RECT 65 110.252 65.072 110.444 ; 
        RECT 120.728 110.252 120.8 110.444 ; 
    END 
  END VSS 
  PIN ADDRESS[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 70.812 45.014 70.884 45.162 ; 
      LAYER M4 ; 
        RECT 70.604 45.046 70.94 45.142 ; 
      LAYER M5 ; 
        RECT 70.8 41.242 70.896 54.202 ; 
      LAYER V3 ; 
        RECT 70.812 45.046 70.884 45.142 ; 
      LAYER V4 ; 
        RECT 70.8 45.046 70.896 45.142 ; 
    END 
  END ADDRESS[0] 
  PIN ADDRESS[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 69.948 45.026 70.02 45.174 ; 
      LAYER M4 ; 
        RECT 69.74 45.046 70.076 45.142 ; 
      LAYER M5 ; 
        RECT 69.936 41.242 70.032 54.202 ; 
      LAYER V3 ; 
        RECT 69.948 45.046 70.02 45.142 ; 
      LAYER V4 ; 
        RECT 69.936 45.046 70.032 45.142 ; 
    END 
  END ADDRESS[1] 
  PIN ADDRESS[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 69.084 42.71 69.156 42.858 ; 
      LAYER M4 ; 
        RECT 68.876 42.742 69.212 42.838 ; 
      LAYER M5 ; 
        RECT 69.072 41.242 69.168 54.202 ; 
      LAYER V3 ; 
        RECT 69.084 42.742 69.156 42.838 ; 
      LAYER V4 ; 
        RECT 69.072 42.742 69.168 42.838 ; 
    END 
  END ADDRESS[2] 
  PIN ADDRESS[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 68.22 43.67 68.292 44.394 ; 
      LAYER M4 ; 
        RECT 68.012 44.278 68.348 44.374 ; 
      LAYER M5 ; 
        RECT 68.208 41.242 68.304 54.202 ; 
      LAYER V3 ; 
        RECT 68.22 44.278 68.292 44.374 ; 
      LAYER V4 ; 
        RECT 68.208 44.278 68.304 44.374 ; 
    END 
  END ADDRESS[3] 
  PIN ADDRESS[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 67.356 42.722 67.428 42.99 ; 
      LAYER M4 ; 
        RECT 67.148 42.742 67.484 42.838 ; 
      LAYER M5 ; 
        RECT 67.344 41.242 67.44 54.202 ; 
      LAYER V3 ; 
        RECT 67.356 42.742 67.428 42.838 ; 
      LAYER V4 ; 
        RECT 67.344 42.742 67.44 42.838 ; 
    END 
  END ADDRESS[4] 
  PIN ADDRESS[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 66.492 41.654 66.564 42.666 ; 
      LAYER M4 ; 
        RECT 66.284 42.55 66.62 42.646 ; 
      LAYER M5 ; 
        RECT 66.48 41.242 66.576 54.202 ; 
      LAYER V3 ; 
        RECT 66.492 42.55 66.564 42.646 ; 
      LAYER V4 ; 
        RECT 66.48 42.55 66.576 42.646 ; 
    END 
  END ADDRESS[5] 
  PIN ADDRESS[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 65.628 45.794 65.7 45.942 ; 
      LAYER M4 ; 
        RECT 65.42 45.814 65.756 45.91 ; 
      LAYER M5 ; 
        RECT 65.616 41.242 65.712 54.202 ; 
      LAYER V3 ; 
        RECT 65.628 45.814 65.7 45.91 ; 
      LAYER V4 ; 
        RECT 65.616 45.814 65.712 45.91 ; 
    END 
  END ADDRESS[6] 
  PIN ADDRESS[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 64.764 45.182 64.836 45.546 ; 
      LAYER M4 ; 
        RECT 64.556 45.43 64.892 45.526 ; 
      LAYER M5 ; 
        RECT 64.752 41.242 64.848 54.202 ; 
      LAYER V3 ; 
        RECT 64.764 45.43 64.836 45.526 ; 
      LAYER V4 ; 
        RECT 64.752 45.43 64.848 45.526 ; 
    END 
  END ADDRESS[7] 
  PIN ADDRESS[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 63.324 43.814 63.396 44.394 ; 
      LAYER M4 ; 
        RECT 63.28 44.278 64.028 44.374 ; 
      LAYER M5 ; 
        RECT 63.888 40.206 63.984 54.202 ; 
      LAYER V3 ; 
        RECT 63.324 44.278 63.396 44.374 ; 
      LAYER V4 ; 
        RECT 63.888 44.278 63.984 44.374 ; 
    END 
  END ADDRESS[8] 
  PIN ADDRESS[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 62.172 42.722 62.244 42.99 ; 
      LAYER M4 ; 
        RECT 61.036 42.742 62.288 42.838 ; 
      LAYER M5 ; 
        RECT 61.08 41.242 61.176 54.202 ; 
      LAYER V3 ; 
        RECT 62.172 42.742 62.244 42.838 ; 
      LAYER V4 ; 
        RECT 61.08 42.742 61.176 42.838 ; 
    END 
  END ADDRESS[9] 
  PIN banksel 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.588 41.654 60.66 42.666 ; 
      LAYER M4 ; 
        RECT 59.74 42.55 60.704 42.646 ; 
      LAYER M5 ; 
        RECT 59.784 41.242 59.88 54.202 ; 
      LAYER V3 ; 
        RECT 60.588 42.55 60.66 42.646 ; 
      LAYER V4 ; 
        RECT 59.784 42.55 59.88 42.646 ; 
    END 
  END banksel 
  PIN clk 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 56.556 46.178 56.628 46.374 ; 
      LAYER M4 ; 
        RECT 56.348 46.198 56.684 46.294 ; 
      LAYER M5 ; 
        RECT 56.544 41.242 56.64 54.202 ; 
      LAYER V3 ; 
        RECT 56.556 46.198 56.628 46.294 ; 
      LAYER V4 ; 
        RECT 56.544 46.198 56.64 46.294 ; 
    END 
  END clk 
  PIN write 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 57.42 42.722 57.492 42.99 ; 
      LAYER M4 ; 
        RECT 57.212 42.742 57.548 42.838 ; 
      LAYER M5 ; 
        RECT 57.408 41.242 57.504 54.202 ; 
      LAYER V3 ; 
        RECT 57.42 42.742 57.492 42.838 ; 
      LAYER V4 ; 
        RECT 57.408 42.742 57.504 42.838 ; 
    END 
  END write 
  PIN read 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 56.7 41.654 56.772 42.666 ; 
      LAYER M4 ; 
        RECT 55.636 42.55 56.816 42.646 ; 
      LAYER M5 ; 
        RECT 55.68 41.242 55.776 54.202 ; 
      LAYER V3 ; 
        RECT 56.7 42.55 56.772 42.646 ; 
      LAYER V4 ; 
        RECT 55.68 42.55 55.776 42.646 ; 
    END 
  END read 
  PIN sdel[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 54.828 45.014 54.9 45.162 ; 
      LAYER M4 ; 
        RECT 54.62 45.046 54.956 45.142 ; 
      LAYER M5 ; 
        RECT 54.816 41.242 54.912 54.202 ; 
      LAYER V3 ; 
        RECT 54.828 45.046 54.9 45.142 ; 
      LAYER V4 ; 
        RECT 54.816 45.046 54.912 45.142 ; 
    END 
  END sdel[0] 
  PIN sdel[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 53.964 42.722 54.036 43.638 ; 
      LAYER M4 ; 
        RECT 53.756 42.742 54.092 42.838 ; 
      LAYER M5 ; 
        RECT 53.952 41.242 54.048 54.202 ; 
      LAYER V3 ; 
        RECT 53.964 42.742 54.036 42.838 ; 
      LAYER V4 ; 
        RECT 53.952 42.742 54.048 42.838 ; 
    END 
  END sdel[1] 
  PIN sdel[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 53.1 41.654 53.172 42.666 ; 
      LAYER M4 ; 
        RECT 52.892 42.55 53.228 42.646 ; 
      LAYER M5 ; 
        RECT 53.088 41.242 53.184 54.202 ; 
      LAYER V3 ; 
        RECT 53.1 42.55 53.172 42.646 ; 
      LAYER V4 ; 
        RECT 53.088 42.55 53.184 42.646 ; 
    END 
  END sdel[2] 
  PIN sdel[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 52.236 42.71 52.308 42.858 ; 
      LAYER M4 ; 
        RECT 52.028 42.742 52.364 42.838 ; 
      LAYER M5 ; 
        RECT 52.224 41.242 52.32 54.202 ; 
      LAYER V3 ; 
        RECT 52.236 42.742 52.308 42.838 ; 
      LAYER V4 ; 
        RECT 52.224 42.742 52.32 42.838 ; 
    END 
  END sdel[3] 
  PIN sdel[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 51.372 45.014 51.444 45.162 ; 
      LAYER M4 ; 
        RECT 51.164 45.046 51.5 45.142 ; 
      LAYER M5 ; 
        RECT 51.36 41.242 51.456 54.202 ; 
      LAYER V3 ; 
        RECT 51.372 45.046 51.444 45.142 ; 
      LAYER V4 ; 
        RECT 51.36 45.046 51.456 45.142 ; 
    END 
  END sdel[4] 
  PIN dataout[14] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 94.498 61.868 95.456 ; 
      LAYER M4 ; 
        RECT 59.444 94.7 62.036 94.796 ; 
      LAYER V3 ; 
        RECT 61.796 94.7 61.868 94.796 ; 
    END 
  END dataout[14] 
  PIN dataout[13] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 90.178 61.868 91.136 ; 
      LAYER M4 ; 
        RECT 59.444 90.38 62.036 90.476 ; 
      LAYER V3 ; 
        RECT 61.796 90.38 61.868 90.476 ; 
    END 
  END dataout[13] 
  PIN dataout[12] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 85.858 61.868 86.816 ; 
      LAYER M4 ; 
        RECT 59.444 86.06 62.036 86.156 ; 
      LAYER V3 ; 
        RECT 61.796 86.06 61.868 86.156 ; 
    END 
  END dataout[12] 
  PIN dataout[11] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 81.538 61.868 82.496 ; 
      LAYER M4 ; 
        RECT 59.444 81.74 62.036 81.836 ; 
      LAYER V3 ; 
        RECT 61.796 81.74 61.868 81.836 ; 
    END 
  END dataout[11] 
  PIN dataout[10] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 77.218 61.868 78.176 ; 
      LAYER M4 ; 
        RECT 59.444 77.42 62.036 77.516 ; 
      LAYER V3 ; 
        RECT 61.796 77.42 61.868 77.516 ; 
    END 
  END dataout[10] 
  PIN dataout[0] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 1.51 61.868 2.468 ; 
      LAYER M4 ; 
        RECT 59.444 1.712 62.036 1.808 ; 
      LAYER V3 ; 
        RECT 61.796 1.712 61.868 1.808 ; 
    END 
  END dataout[0] 
  PIN dataout[15] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 98.818 61.868 99.776 ; 
      LAYER M4 ; 
        RECT 59.444 99.02 62.036 99.116 ; 
      LAYER V3 ; 
        RECT 61.796 99.02 61.868 99.116 ; 
    END 
  END dataout[15] 
  PIN dataout[16] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 103.138 61.868 104.096 ; 
      LAYER M4 ; 
        RECT 59.444 103.34 62.036 103.436 ; 
      LAYER V3 ; 
        RECT 61.796 103.34 61.868 103.436 ; 
    END 
  END dataout[16] 
  PIN dataout[17] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 107.458 61.868 108.416 ; 
      LAYER M4 ; 
        RECT 59.444 107.66 62.036 107.756 ; 
      LAYER V3 ; 
        RECT 61.796 107.66 61.868 107.756 ; 
    END 
  END dataout[17] 
  PIN dataout[18] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[18] 
  PIN dataout[19] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[19] 
  PIN dataout[1] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 5.83 61.868 6.788 ; 
      LAYER M4 ; 
        RECT 59.444 6.032 62.036 6.128 ; 
      LAYER V3 ; 
        RECT 61.796 6.032 61.868 6.128 ; 
    END 
  END dataout[1] 
  PIN dataout[20] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[20] 
  PIN dataout[21] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[21] 
  PIN dataout[22] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[22] 
  PIN dataout[23] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[23] 
  PIN dataout[24] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[24] 
  PIN dataout[25] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[25] 
  PIN dataout[26] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[26] 
  PIN dataout[27] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[27] 
  PIN dataout[28] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[28] 
  PIN dataout[29] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[29] 
  PIN dataout[2] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 10.15 61.868 11.108 ; 
      LAYER M4 ; 
        RECT 59.444 10.352 62.036 10.448 ; 
      LAYER V3 ; 
        RECT 61.796 10.352 61.868 10.448 ; 
    END 
  END dataout[2] 
  PIN dataout[30] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[30] 
  PIN dataout[31] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[31] 
  PIN dataout[32] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[32] 
  PIN dataout[33] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[33] 
  PIN dataout[34] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[34] 
  PIN dataout[35] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[35] 
  PIN dataout[36] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[36] 
  PIN dataout[37] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[37] 
  PIN dataout[38] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[38] 
  PIN dataout[39] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[39] 
  PIN dataout[3] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 14.47 61.868 15.428 ; 
      LAYER M4 ; 
        RECT 59.444 14.672 62.036 14.768 ; 
      LAYER V3 ; 
        RECT 61.796 14.672 61.868 14.768 ; 
    END 
  END dataout[3] 
  PIN dataout[40] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[40] 
  PIN dataout[41] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[41] 
  PIN dataout[42] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[42] 
  PIN dataout[43] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[43] 
  PIN dataout[44] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[44] 
  PIN dataout[45] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[45] 
  PIN dataout[46] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[46] 
  PIN dataout[47] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[47] 
  PIN dataout[48] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[48] 
  PIN dataout[49] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[49] 
  PIN dataout[4] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 18.79 61.868 19.748 ; 
      LAYER M4 ; 
        RECT 59.444 18.992 62.036 19.088 ; 
      LAYER V3 ; 
        RECT 61.796 18.992 61.868 19.088 ; 
    END 
  END dataout[4] 
  PIN dataout[50] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[50] 
  PIN dataout[51] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[51] 
  PIN dataout[52] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[52] 
  PIN dataout[53] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[53] 
  PIN dataout[54] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[54] 
  PIN dataout[55] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[55] 
  PIN dataout[56] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[56] 
  PIN dataout[57] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[57] 
  PIN dataout[58] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[58] 
  PIN dataout[59] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[59] 
  PIN dataout[5] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 23.11 61.868 24.068 ; 
      LAYER M4 ; 
        RECT 59.444 23.312 62.036 23.408 ; 
      LAYER V3 ; 
        RECT 61.796 23.312 61.868 23.408 ; 
    END 
  END dataout[5] 
  PIN dataout[60] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[60] 
  PIN dataout[61] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[61] 
  PIN dataout[62] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[62] 
  PIN dataout[63] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END dataout[63] 
  PIN dataout[6] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 27.43 61.868 28.388 ; 
      LAYER M4 ; 
        RECT 59.444 27.632 62.036 27.728 ; 
      LAYER V3 ; 
        RECT 61.796 27.632 61.868 27.728 ; 
    END 
  END dataout[6] 
  PIN dataout[7] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 31.75 61.868 32.708 ; 
      LAYER M4 ; 
        RECT 59.444 31.952 62.036 32.048 ; 
      LAYER V3 ; 
        RECT 61.796 31.952 61.868 32.048 ; 
    END 
  END dataout[7] 
  PIN dataout[8] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 36.07 61.868 37.028 ; 
      LAYER M4 ; 
        RECT 59.444 36.272 62.036 36.368 ; 
      LAYER V3 ; 
        RECT 61.796 36.272 61.868 36.368 ; 
    END 
  END dataout[8] 
  PIN dataout[9] 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 61.796 72.898 61.868 73.856 ; 
      LAYER M4 ; 
        RECT 59.444 73.1 62.036 73.196 ; 
      LAYER V3 ; 
        RECT 61.796 73.1 61.868 73.196 ; 
    END 
  END dataout[9] 
  PIN wd[0] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 1.08 60.968 2.7 ; 
      LAYER M4 ; 
        RECT 59.444 1.328 61.988 1.424 ; 
      LAYER V3 ; 
        RECT 60.896 1.328 60.968 1.424 ; 
    END 
  END wd[0] 
  PIN wd[10] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 76.788 60.968 78.408 ; 
      LAYER M4 ; 
        RECT 59.444 77.036 61.988 77.132 ; 
      LAYER V3 ; 
        RECT 60.896 77.036 60.968 77.132 ; 
    END 
  END wd[10] 
  PIN wd[11] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 81.108 60.968 82.728 ; 
      LAYER M4 ; 
        RECT 59.444 81.356 61.988 81.452 ; 
      LAYER V3 ; 
        RECT 60.896 81.356 60.968 81.452 ; 
    END 
  END wd[11] 
  PIN wd[12] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 85.428 60.968 87.048 ; 
      LAYER M4 ; 
        RECT 59.444 85.676 61.988 85.772 ; 
      LAYER V3 ; 
        RECT 60.896 85.676 60.968 85.772 ; 
    END 
  END wd[12] 
  PIN wd[13] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 89.748 60.968 91.368 ; 
      LAYER M4 ; 
        RECT 59.444 89.996 61.988 90.092 ; 
      LAYER V3 ; 
        RECT 60.896 89.996 60.968 90.092 ; 
    END 
  END wd[13] 
  PIN wd[14] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 94.068 60.968 95.688 ; 
      LAYER M4 ; 
        RECT 59.444 94.316 61.988 94.412 ; 
      LAYER V3 ; 
        RECT 60.896 94.316 60.968 94.412 ; 
    END 
  END wd[14] 
  PIN wd[15] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 98.388 60.968 100.008 ; 
      LAYER M4 ; 
        RECT 59.444 98.636 61.988 98.732 ; 
      LAYER V3 ; 
        RECT 60.896 98.636 60.968 98.732 ; 
    END 
  END wd[15] 
  PIN wd[16] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 102.708 60.968 104.328 ; 
      LAYER M4 ; 
        RECT 59.444 102.956 61.988 103.052 ; 
      LAYER V3 ; 
        RECT 60.896 102.956 60.968 103.052 ; 
    END 
  END wd[16] 
  PIN wd[17] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 107.028 60.968 108.648 ; 
      LAYER M4 ; 
        RECT 59.444 107.276 61.988 107.372 ; 
      LAYER V3 ; 
        RECT 60.896 107.276 60.968 107.372 ; 
    END 
  END wd[17] 
  PIN wd[18] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[18] 
  PIN wd[19] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[19] 
  PIN wd[1] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 5.4 60.968 7.02 ; 
      LAYER M4 ; 
        RECT 59.444 5.648 61.988 5.744 ; 
      LAYER V3 ; 
        RECT 60.896 5.648 60.968 5.744 ; 
    END 
  END wd[1] 
  PIN wd[20] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[20] 
  PIN wd[21] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[21] 
  PIN wd[22] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[22] 
  PIN wd[23] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[23] 
  PIN wd[24] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[24] 
  PIN wd[25] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[25] 
  PIN wd[26] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[26] 
  PIN wd[27] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[27] 
  PIN wd[28] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[28] 
  PIN wd[29] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[29] 
  PIN wd[2] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 9.72 60.968 11.34 ; 
      LAYER M4 ; 
        RECT 59.444 9.968 61.988 10.064 ; 
      LAYER V3 ; 
        RECT 60.896 9.968 60.968 10.064 ; 
    END 
  END wd[2] 
  PIN wd[30] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[30] 
  PIN wd[31] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[31] 
  PIN wd[32] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[32] 
  PIN wd[33] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[33] 
  PIN wd[34] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[34] 
  PIN wd[35] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[35] 
  PIN wd[36] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[36] 
  PIN wd[37] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[37] 
  PIN wd[38] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[38] 
  PIN wd[39] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[39] 
  PIN wd[3] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 14.04 60.968 15.66 ; 
      LAYER M4 ; 
        RECT 59.444 14.288 61.988 14.384 ; 
      LAYER V3 ; 
        RECT 60.896 14.288 60.968 14.384 ; 
    END 
  END wd[3] 
  PIN wd[40] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[40] 
  PIN wd[41] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[41] 
  PIN wd[42] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[42] 
  PIN wd[43] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[43] 
  PIN wd[44] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[44] 
  PIN wd[45] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[45] 
  PIN wd[46] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[46] 
  PIN wd[47] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[47] 
  PIN wd[48] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[48] 
  PIN wd[49] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[49] 
  PIN wd[4] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 18.36 60.968 19.98 ; 
      LAYER M4 ; 
        RECT 59.444 18.608 61.988 18.704 ; 
      LAYER V3 ; 
        RECT 60.896 18.608 60.968 18.704 ; 
    END 
  END wd[4] 
  PIN wd[50] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[50] 
  PIN wd[51] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[51] 
  PIN wd[52] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[52] 
  PIN wd[53] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[53] 
  PIN wd[54] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[54] 
  PIN wd[55] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[55] 
  PIN wd[56] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[56] 
  PIN wd[57] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[57] 
  PIN wd[58] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[58] 
  PIN wd[59] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[59] 
  PIN wd[5] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 22.68 60.968 24.3 ; 
      LAYER M4 ; 
        RECT 59.444 22.928 61.988 23.024 ; 
      LAYER V3 ; 
        RECT 60.896 22.928 60.968 23.024 ; 
    END 
  END wd[5] 
  PIN wd[60] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[60] 
  PIN wd[61] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[61] 
  PIN wd[62] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[62] 
  PIN wd[63] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
    END 
  END wd[63] 
  PIN wd[6] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 27 60.968 28.62 ; 
      LAYER M4 ; 
        RECT 59.444 27.248 61.988 27.344 ; 
      LAYER V3 ; 
        RECT 60.896 27.248 60.968 27.344 ; 
    END 
  END wd[6] 
  PIN wd[7] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 31.32 60.968 32.94 ; 
      LAYER M4 ; 
        RECT 59.444 31.568 61.988 31.664 ; 
      LAYER V3 ; 
        RECT 60.896 31.568 60.968 31.664 ; 
    END 
  END wd[7] 
  PIN wd[8] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 35.64 60.968 37.26 ; 
      LAYER M4 ; 
        RECT 59.444 35.888 61.988 35.984 ; 
      LAYER V3 ; 
        RECT 60.896 35.888 60.968 35.984 ; 
    END 
  END wd[8] 
  PIN wd[9] 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M3 ; 
        RECT 60.896 72.468 60.968 74.088 ; 
      LAYER M4 ; 
        RECT 59.444 72.716 61.988 72.812 ; 
      LAYER V3 ; 
        RECT 60.896 72.716 60.968 72.812 ; 
    END 
  END wd[9] 
OBS 
  LAYER M1 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0 40.054 121.392 74.668 ; 
        RECT 0.02 72.414 121.412 76.788 ; 
        RECT 0.02 76.734 121.412 81.108 ; 
        RECT 0.02 81.054 121.412 85.428 ; 
        RECT 0.02 85.374 121.412 89.748 ; 
        RECT 0.02 89.694 121.412 94.068 ; 
        RECT 0.02 94.014 121.412 98.388 ; 
        RECT 0.02 98.334 121.412 102.708 ; 
        RECT 0.02 102.654 121.412 107.028 ; 
        RECT 0.02 106.974 121.412 111.348 ; 
  LAYER M2 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0 40.054 121.392 74.668 ; 
        RECT 0.02 72.414 121.412 76.788 ; 
        RECT 0.02 76.734 121.412 81.108 ; 
        RECT 0.02 81.054 121.412 85.428 ; 
        RECT 0.02 85.374 121.412 89.748 ; 
        RECT 0.02 89.694 121.412 94.068 ; 
        RECT 0.02 94.014 121.412 98.388 ; 
        RECT 0.02 98.334 121.412 102.708 ; 
        RECT 0.02 102.654 121.412 107.028 ; 
        RECT 0.02 106.974 121.412 111.348 ; 
  LAYER V1 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0 40.054 121.392 74.668 ; 
        RECT 0.02 72.414 121.412 76.788 ; 
        RECT 0.02 76.734 121.412 81.108 ; 
        RECT 0.02 81.054 121.412 85.428 ; 
        RECT 0.02 85.374 121.412 89.748 ; 
        RECT 0.02 89.694 121.412 94.068 ; 
        RECT 0.02 94.014 121.412 98.388 ; 
        RECT 0.02 98.334 121.412 102.708 ; 
        RECT 0.02 102.654 121.412 107.028 ; 
        RECT 0.02 106.974 121.412 111.348 ; 
  LAYER V2 SPACING 0.072 ; 
      RECT 0.02 1.026 121.412 5.4 ; 
      RECT 0.02 5.346 121.412 9.72 ; 
      RECT 0.02 9.666 121.412 14.04 ; 
      RECT 0.02 13.986 121.412 18.36 ; 
      RECT 0.02 18.306 121.412 22.68 ; 
      RECT 0.02 22.626 121.412 27 ; 
      RECT 0.02 26.946 121.412 31.32 ; 
      RECT 0.02 31.266 121.412 35.64 ; 
      RECT 0.02 35.586 121.412 39.96 ; 
      RECT 0 40.054 121.392 74.668 ; 
        RECT 0.02 72.414 121.412 76.788 ; 
        RECT 0.02 76.734 121.412 81.108 ; 
        RECT 0.02 81.054 121.412 85.428 ; 
        RECT 0.02 85.374 121.412 89.748 ; 
        RECT 0.02 89.694 121.412 94.068 ; 
        RECT 0.02 94.014 121.412 98.388 ; 
        RECT 0.02 98.334 121.412 102.708 ; 
        RECT 0.02 102.654 121.412 107.028 ; 
        RECT 0.02 106.974 121.412 111.348 ; 
  LAYER M3 ; 
      RECT 62.444 1.38 62.516 5.122 ; 
      RECT 62.3 1.38 62.372 5.122 ; 
      RECT 62.156 3.688 62.228 4.978 ; 
      RECT 61.688 4.476 61.76 4.914 ; 
      RECT 61.652 1.51 61.724 2.468 ; 
      RECT 61.508 3.834 61.58 4.448 ; 
      RECT 61.184 3.936 61.256 4.968 ; 
      RECT 59.024 1.38 59.096 5.122 ; 
      RECT 58.88 1.38 58.952 5.122 ; 
      RECT 58.736 2.104 58.808 4.376 ; 
      RECT 62.444 5.7 62.516 9.442 ; 
      RECT 62.3 5.7 62.372 9.442 ; 
      RECT 62.156 8.008 62.228 9.298 ; 
      RECT 61.688 8.796 61.76 9.234 ; 
      RECT 61.652 5.83 61.724 6.788 ; 
      RECT 61.508 8.154 61.58 8.768 ; 
      RECT 61.184 8.256 61.256 9.288 ; 
      RECT 59.024 5.7 59.096 9.442 ; 
      RECT 58.88 5.7 58.952 9.442 ; 
      RECT 58.736 6.424 58.808 8.696 ; 
      RECT 62.444 10.02 62.516 13.762 ; 
      RECT 62.3 10.02 62.372 13.762 ; 
      RECT 62.156 12.328 62.228 13.618 ; 
      RECT 61.688 13.116 61.76 13.554 ; 
      RECT 61.652 10.15 61.724 11.108 ; 
      RECT 61.508 12.474 61.58 13.088 ; 
      RECT 61.184 12.576 61.256 13.608 ; 
      RECT 59.024 10.02 59.096 13.762 ; 
      RECT 58.88 10.02 58.952 13.762 ; 
      RECT 58.736 10.744 58.808 13.016 ; 
      RECT 62.444 14.34 62.516 18.082 ; 
      RECT 62.3 14.34 62.372 18.082 ; 
      RECT 62.156 16.648 62.228 17.938 ; 
      RECT 61.688 17.436 61.76 17.874 ; 
      RECT 61.652 14.47 61.724 15.428 ; 
      RECT 61.508 16.794 61.58 17.408 ; 
      RECT 61.184 16.896 61.256 17.928 ; 
      RECT 59.024 14.34 59.096 18.082 ; 
      RECT 58.88 14.34 58.952 18.082 ; 
      RECT 58.736 15.064 58.808 17.336 ; 
      RECT 62.444 18.66 62.516 22.402 ; 
      RECT 62.3 18.66 62.372 22.402 ; 
      RECT 62.156 20.968 62.228 22.258 ; 
      RECT 61.688 21.756 61.76 22.194 ; 
      RECT 61.652 18.79 61.724 19.748 ; 
      RECT 61.508 21.114 61.58 21.728 ; 
      RECT 61.184 21.216 61.256 22.248 ; 
      RECT 59.024 18.66 59.096 22.402 ; 
      RECT 58.88 18.66 58.952 22.402 ; 
      RECT 58.736 19.384 58.808 21.656 ; 
      RECT 62.444 22.98 62.516 26.722 ; 
      RECT 62.3 22.98 62.372 26.722 ; 
      RECT 62.156 25.288 62.228 26.578 ; 
      RECT 61.688 26.076 61.76 26.514 ; 
      RECT 61.652 23.11 61.724 24.068 ; 
      RECT 61.508 25.434 61.58 26.048 ; 
      RECT 61.184 25.536 61.256 26.568 ; 
      RECT 59.024 22.98 59.096 26.722 ; 
      RECT 58.88 22.98 58.952 26.722 ; 
      RECT 58.736 23.704 58.808 25.976 ; 
      RECT 62.444 27.3 62.516 31.042 ; 
      RECT 62.3 27.3 62.372 31.042 ; 
      RECT 62.156 29.608 62.228 30.898 ; 
      RECT 61.688 30.396 61.76 30.834 ; 
      RECT 61.652 27.43 61.724 28.388 ; 
      RECT 61.508 29.754 61.58 30.368 ; 
      RECT 61.184 29.856 61.256 30.888 ; 
      RECT 59.024 27.3 59.096 31.042 ; 
      RECT 58.88 27.3 58.952 31.042 ; 
      RECT 58.736 28.024 58.808 30.296 ; 
      RECT 62.444 31.62 62.516 35.362 ; 
      RECT 62.3 31.62 62.372 35.362 ; 
      RECT 62.156 33.928 62.228 35.218 ; 
      RECT 61.688 34.716 61.76 35.154 ; 
      RECT 61.652 31.75 61.724 32.708 ; 
      RECT 61.508 34.074 61.58 34.688 ; 
      RECT 61.184 34.176 61.256 35.208 ; 
      RECT 59.024 31.62 59.096 35.362 ; 
      RECT 58.88 31.62 58.952 35.362 ; 
      RECT 58.736 32.344 58.808 34.616 ; 
      RECT 62.444 35.94 62.516 39.682 ; 
      RECT 62.3 35.94 62.372 39.682 ; 
      RECT 62.156 38.248 62.228 39.538 ; 
      RECT 61.688 39.036 61.76 39.474 ; 
      RECT 61.652 36.07 61.724 37.028 ; 
      RECT 61.508 38.394 61.58 39.008 ; 
      RECT 61.184 38.496 61.256 39.528 ; 
      RECT 59.024 35.94 59.096 39.682 ; 
      RECT 58.88 35.94 58.952 39.682 ; 
      RECT 58.736 36.664 58.808 38.936 ; 
      RECT 120.852 39.294 120.924 72.776 ; 
      RECT 120.708 39.294 120.78 72.776 ; 
      RECT 120.276 39.294 120.348 54.258 ; 
      RECT 119.844 39.294 119.916 54.258 ; 
      RECT 119.412 39.294 119.484 54.258 ; 
      RECT 118.98 39.294 119.052 54.258 ; 
      RECT 118.548 39.294 118.62 54.258 ; 
      RECT 118.116 39.294 118.188 54.258 ; 
      RECT 117.684 39.294 117.756 54.258 ; 
      RECT 117.252 39.294 117.324 54.258 ; 
      RECT 116.82 39.294 116.892 54.258 ; 
      RECT 116.388 39.294 116.46 54.258 ; 
      RECT 115.956 39.294 116.028 54.258 ; 
      RECT 115.524 39.294 115.596 54.258 ; 
      RECT 115.092 39.294 115.164 54.258 ; 
      RECT 114.66 39.294 114.732 54.258 ; 
      RECT 114.228 39.294 114.3 54.258 ; 
      RECT 113.796 39.294 113.868 54.258 ; 
      RECT 113.364 39.294 113.436 54.258 ; 
      RECT 112.932 39.294 113.004 54.258 ; 
      RECT 112.5 39.294 112.572 54.258 ; 
      RECT 112.068 39.294 112.14 54.258 ; 
      RECT 111.636 39.294 111.708 54.258 ; 
      RECT 111.204 39.294 111.276 54.258 ; 
      RECT 110.772 39.294 110.844 54.258 ; 
      RECT 110.34 39.294 110.412 54.258 ; 
      RECT 109.908 39.294 109.98 54.258 ; 
      RECT 109.476 39.294 109.548 54.258 ; 
      RECT 109.044 39.294 109.116 54.258 ; 
      RECT 108.612 39.294 108.684 54.258 ; 
      RECT 108.18 39.294 108.252 54.258 ; 
      RECT 107.748 39.294 107.82 54.258 ; 
      RECT 107.316 39.294 107.388 54.258 ; 
      RECT 106.884 39.294 106.956 54.258 ; 
      RECT 106.452 39.294 106.524 54.258 ; 
      RECT 106.02 39.294 106.092 54.258 ; 
      RECT 105.588 39.294 105.66 54.258 ; 
      RECT 105.156 39.294 105.228 54.258 ; 
      RECT 104.724 39.294 104.796 54.258 ; 
      RECT 104.292 39.294 104.364 54.258 ; 
      RECT 103.86 39.294 103.932 54.258 ; 
      RECT 103.428 39.294 103.5 54.258 ; 
      RECT 102.996 39.294 103.068 54.258 ; 
      RECT 102.564 39.294 102.636 54.258 ; 
      RECT 102.132 39.294 102.204 54.258 ; 
      RECT 101.7 39.294 101.772 54.258 ; 
      RECT 101.268 39.294 101.34 54.258 ; 
      RECT 100.836 39.294 100.908 54.258 ; 
      RECT 100.404 39.294 100.476 54.258 ; 
      RECT 99.972 39.294 100.044 54.258 ; 
      RECT 99.54 39.294 99.612 54.258 ; 
      RECT 99.108 39.294 99.18 54.258 ; 
      RECT 98.676 39.294 98.748 54.258 ; 
      RECT 98.244 39.294 98.316 54.258 ; 
      RECT 97.812 39.294 97.884 54.258 ; 
      RECT 97.38 39.294 97.452 54.258 ; 
      RECT 96.948 39.294 97.02 54.258 ; 
      RECT 96.516 39.294 96.588 54.258 ; 
      RECT 96.084 39.294 96.156 54.258 ; 
      RECT 95.652 39.294 95.724 54.258 ; 
      RECT 95.22 39.294 95.292 54.258 ; 
      RECT 94.788 39.294 94.86 54.258 ; 
      RECT 94.356 39.294 94.428 54.258 ; 
      RECT 93.924 39.294 93.996 54.258 ; 
      RECT 93.492 39.294 93.564 54.258 ; 
      RECT 93.06 39.294 93.132 54.258 ; 
      RECT 92.628 39.294 92.7 54.258 ; 
      RECT 92.196 39.294 92.268 54.258 ; 
      RECT 91.764 39.294 91.836 54.258 ; 
      RECT 91.332 39.294 91.404 54.258 ; 
      RECT 90.9 39.294 90.972 54.258 ; 
      RECT 90.468 39.294 90.54 54.258 ; 
      RECT 90.036 39.294 90.108 54.258 ; 
      RECT 89.604 39.294 89.676 54.258 ; 
      RECT 89.172 39.294 89.244 54.258 ; 
      RECT 88.74 39.294 88.812 54.258 ; 
      RECT 88.308 39.294 88.38 54.258 ; 
      RECT 87.876 39.294 87.948 54.258 ; 
      RECT 87.444 39.294 87.516 54.258 ; 
      RECT 87.012 39.294 87.084 54.258 ; 
      RECT 86.58 39.294 86.652 54.258 ; 
      RECT 86.148 39.294 86.22 54.258 ; 
      RECT 85.716 39.294 85.788 54.258 ; 
      RECT 85.284 39.294 85.356 54.258 ; 
      RECT 84.852 39.294 84.924 54.258 ; 
      RECT 84.42 39.294 84.492 54.258 ; 
      RECT 83.988 39.294 84.06 54.258 ; 
      RECT 83.556 39.294 83.628 54.258 ; 
      RECT 83.124 39.294 83.196 54.258 ; 
      RECT 82.692 39.294 82.764 54.258 ; 
      RECT 82.26 39.294 82.332 54.258 ; 
      RECT 81.828 39.294 81.9 54.258 ; 
      RECT 81.396 39.294 81.468 54.258 ; 
      RECT 80.964 39.294 81.036 54.258 ; 
      RECT 80.532 39.294 80.604 54.258 ; 
      RECT 80.1 39.294 80.172 54.258 ; 
      RECT 79.668 39.294 79.74 54.258 ; 
      RECT 79.236 39.948 79.308 41.348 ; 
      RECT 78.804 39.294 78.876 54.258 ; 
      RECT 78.372 39.294 78.444 54.258 ; 
      RECT 77.94 39.294 78.012 54.258 ; 
      RECT 77.508 39.294 77.58 54.258 ; 
      RECT 77.076 39.294 77.148 54.258 ; 
      RECT 76.644 39.294 76.716 54.258 ; 
      RECT 76.212 39.294 76.284 54.258 ; 
      RECT 75.78 39.294 75.852 54.258 ; 
      RECT 75.348 39.294 75.42 54.258 ; 
      RECT 74.916 39.294 74.988 54.258 ; 
      RECT 74.484 39.294 74.556 54.258 ; 
      RECT 74.052 39.294 74.124 54.258 ; 
      RECT 73.62 39.294 73.692 54.258 ; 
      RECT 73.188 39.294 73.26 54.258 ; 
      RECT 72.756 39.294 72.828 54.258 ; 
      RECT 72.324 39.294 72.396 54.258 ; 
      RECT 71.892 39.294 71.964 54.258 ; 
      RECT 71.46 39.294 71.532 54.258 ; 
      RECT 71.028 39.294 71.1 54.258 ; 
      RECT 70.596 39.294 70.668 54.258 ; 
      RECT 70.164 39.294 70.236 54.258 ; 
      RECT 69.732 39.294 69.804 54.258 ; 
      RECT 69.3 39.294 69.372 54.258 ; 
      RECT 68.868 39.294 68.94 54.258 ; 
      RECT 68.436 39.294 68.508 54.258 ; 
      RECT 68.004 39.294 68.076 54.258 ; 
      RECT 67.572 39.294 67.644 54.258 ; 
      RECT 67.14 39.294 67.212 54.258 ; 
      RECT 66.708 39.294 66.78 54.258 ; 
      RECT 66.276 39.294 66.348 54.258 ; 
      RECT 65.844 39.294 65.916 54.258 ; 
      RECT 65.7 55.102 65.772 57.9208 ; 
      RECT 65.7 60.874 65.772 65.518 ; 
      RECT 65.628 42.59 65.7 45.294 ; 
      RECT 65.628 48.278 65.7 49.47 ; 
      RECT 65.628 52.742 65.7 53.79 ; 
      RECT 65.556 55.356 65.628 58.116 ; 
      RECT 65.556 58.32 65.628 62.262 ; 
      RECT 65.556 62.426 65.628 64.894 ; 
      RECT 65.412 39.294 65.484 72.776 ; 
      RECT 65.268 56.446 65.34 56.778 ; 
      RECT 65.196 43.022 65.268 45.546 ; 
      RECT 65.196 47.198 65.268 47.958 ; 
      RECT 65.196 50.726 65.268 50.922 ; 
      RECT 65.196 53.654 65.268 53.802 ; 
      RECT 65.124 55.226 65.196 69.598 ; 
      RECT 64.764 40.08 64.836 40.632 ; 
      RECT 64.764 41.51 64.836 44.718 ; 
      RECT 64.764 46.91 64.836 49.182 ; 
      RECT 64.764 55.226 64.836 69.598 ; 
      RECT 64.62 47.198 64.692 48.678 ; 
      RECT 64.476 44.606 64.548 45.15 ; 
      RECT 64.476 48.566 64.548 49.47 ; 
      RECT 64.476 53.534 64.548 53.79 ; 
      RECT 64.332 45.014 64.404 45.162 ; 
      RECT 64.332 51.518 64.404 51.69 ; 
      RECT 64.332 53.654 64.404 53.802 ; 
      RECT 64.188 46.262 64.26 48.246 ; 
      RECT 64.188 48.422 64.26 49.182 ; 
      RECT 64.188 52.262 64.26 53.502 ; 
      RECT 64.044 45.83 64.116 50.818 ; 
      RECT 60.156 40.054 60.228 40.67 ; 
      RECT 60.012 40.054 60.084 40.254 ; 
      RECT 59.724 40.054 59.796 40.34 ; 
      RECT 57.132 44.606 57.204 46.23 ; 
      RECT 56.988 49.046 57.06 49.194 ; 
      RECT 56.844 44.75 56.916 47.166 ; 
      RECT 56.7 44.102 56.772 44.358 ; 
      RECT 56.556 40.266 56.628 40.47 ; 
      RECT 56.556 52.742 56.628 53.502 ; 
      RECT 56.556 55.226 56.628 69.598 ; 
      RECT 56.124 41.942 56.196 42.702 ; 
      RECT 56.124 45.038 56.196 54.078 ; 
      RECT 56.052 56.446 56.124 56.778 ; 
      RECT 55.908 39.948 55.98 72.776 ; 
      RECT 55.764 55.356 55.836 58.116 ; 
      RECT 55.764 58.32 55.836 62.262 ; 
      RECT 55.764 62.426 55.836 64.894 ; 
      RECT 55.692 41.942 55.764 43.926 ; 
      RECT 55.692 47.054 55.764 49.326 ; 
      RECT 55.692 50.582 55.764 53.502 ; 
      RECT 55.62 55.102 55.692 57.9208 ; 
      RECT 55.62 60.874 55.692 65.518 ; 
      RECT 55.476 39.948 55.548 41.348 ; 
      RECT 55.476 54.124 55.548 72.776 ; 
      RECT 55.044 39.948 55.116 41.348 ; 
      RECT 54.612 39.948 54.684 41.348 ; 
      RECT 54.18 39.948 54.252 41.348 ; 
      RECT 53.748 39.948 53.82 41.348 ; 
      RECT 53.316 39.948 53.388 41.348 ; 
      RECT 52.884 39.948 52.956 41.348 ; 
      RECT 52.452 39.948 52.524 41.348 ; 
      RECT 52.02 39.948 52.092 41.348 ; 
      RECT 51.588 39.948 51.66 41.348 ; 
      RECT 51.156 39.948 51.228 41.348 ; 
      RECT 50.724 39.948 50.796 41.348 ; 
      RECT 50.292 39.948 50.364 41.348 ; 
      RECT 49.86 39.948 49.932 41.348 ; 
      RECT 49.428 39.948 49.5 41.348 ; 
      RECT 48.996 39.948 49.068 41.348 ; 
      RECT 48.564 39.948 48.636 41.348 ; 
      RECT 48.132 39.948 48.204 41.348 ; 
      RECT 47.7 39.948 47.772 41.348 ; 
      RECT 47.268 39.948 47.34 41.348 ; 
      RECT 46.836 39.948 46.908 41.348 ; 
      RECT 46.404 39.948 46.476 41.348 ; 
      RECT 45.972 39.948 46.044 41.348 ; 
      RECT 45.54 39.948 45.612 41.348 ; 
      RECT 45.108 39.948 45.18 41.348 ; 
      RECT 44.676 39.948 44.748 41.348 ; 
      RECT 44.244 39.948 44.316 41.348 ; 
      RECT 43.812 39.948 43.884 41.348 ; 
      RECT 43.38 39.948 43.452 41.348 ; 
      RECT 42.948 39.948 43.02 41.348 ; 
      RECT 42.516 39.948 42.588 41.348 ; 
      RECT 42.084 39.948 42.156 41.348 ; 
      RECT 41.652 39.948 41.724 41.348 ; 
      RECT 41.22 39.948 41.292 41.348 ; 
      RECT 40.788 39.948 40.86 41.348 ; 
      RECT 40.356 39.948 40.428 41.348 ; 
      RECT 39.924 39.948 39.996 41.348 ; 
      RECT 39.492 39.948 39.564 41.348 ; 
      RECT 39.06 39.948 39.132 41.348 ; 
      RECT 38.628 39.948 38.7 41.348 ; 
      RECT 38.196 39.948 38.268 41.348 ; 
      RECT 37.764 39.948 37.836 41.348 ; 
      RECT 37.332 39.948 37.404 41.348 ; 
      RECT 36.9 39.948 36.972 41.348 ; 
      RECT 36.468 39.948 36.54 41.348 ; 
      RECT 36.036 39.948 36.108 41.348 ; 
      RECT 35.604 39.948 35.676 41.348 ; 
      RECT 35.172 39.948 35.244 41.348 ; 
      RECT 34.74 39.948 34.812 41.348 ; 
      RECT 34.308 39.948 34.38 41.348 ; 
      RECT 33.876 39.948 33.948 41.348 ; 
      RECT 33.444 39.948 33.516 41.348 ; 
      RECT 33.012 39.948 33.084 41.348 ; 
      RECT 32.58 39.948 32.652 41.348 ; 
      RECT 32.148 39.948 32.22 41.348 ; 
      RECT 31.716 39.948 31.788 41.348 ; 
      RECT 31.284 39.948 31.356 41.348 ; 
      RECT 30.852 39.948 30.924 41.348 ; 
      RECT 30.42 39.948 30.492 41.348 ; 
      RECT 29.988 39.948 30.06 41.348 ; 
      RECT 29.556 39.948 29.628 41.348 ; 
      RECT 29.124 39.948 29.196 41.348 ; 
      RECT 28.692 39.948 28.764 41.348 ; 
      RECT 28.26 39.948 28.332 41.348 ; 
      RECT 27.828 39.948 27.9 41.348 ; 
      RECT 27.396 39.948 27.468 41.348 ; 
      RECT 26.964 39.948 27.036 41.348 ; 
      RECT 26.532 39.948 26.604 41.348 ; 
      RECT 26.1 39.948 26.172 41.348 ; 
      RECT 25.668 39.948 25.74 41.348 ; 
      RECT 25.236 39.948 25.308 41.348 ; 
      RECT 24.804 39.948 24.876 41.348 ; 
      RECT 24.372 39.948 24.444 41.348 ; 
      RECT 23.94 39.948 24.012 41.348 ; 
      RECT 23.508 39.948 23.58 41.348 ; 
      RECT 23.076 39.948 23.148 41.348 ; 
      RECT 22.644 39.948 22.716 41.348 ; 
      RECT 22.212 39.948 22.284 41.348 ; 
      RECT 21.78 39.948 21.852 41.348 ; 
      RECT 21.348 39.948 21.42 41.348 ; 
      RECT 20.916 39.948 20.988 41.348 ; 
      RECT 20.484 39.948 20.556 41.348 ; 
      RECT 20.052 39.948 20.124 41.348 ; 
      RECT 19.62 39.948 19.692 41.348 ; 
      RECT 19.188 39.948 19.26 41.348 ; 
      RECT 18.756 39.948 18.828 41.348 ; 
      RECT 18.324 39.948 18.396 41.348 ; 
      RECT 17.892 39.948 17.964 41.348 ; 
      RECT 17.46 39.948 17.532 41.348 ; 
      RECT 17.028 39.948 17.1 41.348 ; 
      RECT 16.596 39.948 16.668 41.348 ; 
      RECT 16.164 39.948 16.236 41.348 ; 
      RECT 15.732 39.948 15.804 41.348 ; 
      RECT 15.3 39.948 15.372 41.348 ; 
      RECT 14.868 39.948 14.94 41.348 ; 
      RECT 14.436 39.948 14.508 41.348 ; 
      RECT 14.004 39.948 14.076 41.348 ; 
      RECT 13.572 39.948 13.644 41.348 ; 
      RECT 13.14 39.948 13.212 41.348 ; 
      RECT 12.708 39.948 12.78 41.348 ; 
      RECT 12.276 39.948 12.348 41.348 ; 
      RECT 11.844 39.948 11.916 41.348 ; 
      RECT 11.412 39.948 11.484 41.348 ; 
      RECT 10.98 39.948 11.052 41.348 ; 
      RECT 10.548 39.948 10.62 41.348 ; 
      RECT 10.116 39.948 10.188 41.348 ; 
      RECT 9.684 39.948 9.756 41.348 ; 
      RECT 9.252 39.948 9.324 41.348 ; 
      RECT 8.82 39.948 8.892 41.348 ; 
      RECT 8.388 39.948 8.46 41.348 ; 
      RECT 7.956 39.948 8.028 41.348 ; 
      RECT 7.524 39.948 7.596 41.348 ; 
      RECT 7.092 39.948 7.164 41.348 ; 
      RECT 6.66 39.948 6.732 41.348 ; 
      RECT 6.228 39.948 6.3 41.348 ; 
      RECT 5.796 39.948 5.868 41.348 ; 
      RECT 5.364 39.948 5.436 41.348 ; 
      RECT 4.932 39.948 5.004 41.348 ; 
      RECT 4.5 39.948 4.572 41.348 ; 
      RECT 4.068 39.948 4.14 41.348 ; 
      RECT 3.636 39.948 3.708 41.348 ; 
      RECT 3.204 39.948 3.276 41.348 ; 
      RECT 2.772 39.948 2.844 41.348 ; 
      RECT 2.34 39.948 2.412 41.348 ; 
      RECT 1.908 39.948 1.98 41.348 ; 
      RECT 1.476 39.948 1.548 41.348 ; 
      RECT 1.044 39.948 1.116 41.348 ; 
      RECT 0.612 39.948 0.684 72.776 ; 
      RECT 0.468 39.948 0.54 72.776 ; 
        RECT 62.444 72.768 62.516 76.51 ; 
        RECT 62.3 72.768 62.372 76.51 ; 
        RECT 62.156 75.076 62.228 76.366 ; 
        RECT 61.688 75.864 61.76 76.302 ; 
        RECT 61.652 72.898 61.724 73.856 ; 
        RECT 61.508 75.222 61.58 75.836 ; 
        RECT 61.184 75.324 61.256 76.356 ; 
        RECT 59.024 72.768 59.096 76.51 ; 
        RECT 58.88 72.768 58.952 76.51 ; 
        RECT 58.736 73.492 58.808 75.764 ; 
        RECT 62.444 77.088 62.516 80.83 ; 
        RECT 62.3 77.088 62.372 80.83 ; 
        RECT 62.156 79.396 62.228 80.686 ; 
        RECT 61.688 80.184 61.76 80.622 ; 
        RECT 61.652 77.218 61.724 78.176 ; 
        RECT 61.508 79.542 61.58 80.156 ; 
        RECT 61.184 79.644 61.256 80.676 ; 
        RECT 59.024 77.088 59.096 80.83 ; 
        RECT 58.88 77.088 58.952 80.83 ; 
        RECT 58.736 77.812 58.808 80.084 ; 
        RECT 62.444 81.408 62.516 85.15 ; 
        RECT 62.3 81.408 62.372 85.15 ; 
        RECT 62.156 83.716 62.228 85.006 ; 
        RECT 61.688 84.504 61.76 84.942 ; 
        RECT 61.652 81.538 61.724 82.496 ; 
        RECT 61.508 83.862 61.58 84.476 ; 
        RECT 61.184 83.964 61.256 84.996 ; 
        RECT 59.024 81.408 59.096 85.15 ; 
        RECT 58.88 81.408 58.952 85.15 ; 
        RECT 58.736 82.132 58.808 84.404 ; 
        RECT 62.444 85.728 62.516 89.47 ; 
        RECT 62.3 85.728 62.372 89.47 ; 
        RECT 62.156 88.036 62.228 89.326 ; 
        RECT 61.688 88.824 61.76 89.262 ; 
        RECT 61.652 85.858 61.724 86.816 ; 
        RECT 61.508 88.182 61.58 88.796 ; 
        RECT 61.184 88.284 61.256 89.316 ; 
        RECT 59.024 85.728 59.096 89.47 ; 
        RECT 58.88 85.728 58.952 89.47 ; 
        RECT 58.736 86.452 58.808 88.724 ; 
        RECT 62.444 90.048 62.516 93.79 ; 
        RECT 62.3 90.048 62.372 93.79 ; 
        RECT 62.156 92.356 62.228 93.646 ; 
        RECT 61.688 93.144 61.76 93.582 ; 
        RECT 61.652 90.178 61.724 91.136 ; 
        RECT 61.508 92.502 61.58 93.116 ; 
        RECT 61.184 92.604 61.256 93.636 ; 
        RECT 59.024 90.048 59.096 93.79 ; 
        RECT 58.88 90.048 58.952 93.79 ; 
        RECT 58.736 90.772 58.808 93.044 ; 
        RECT 62.444 94.368 62.516 98.11 ; 
        RECT 62.3 94.368 62.372 98.11 ; 
        RECT 62.156 96.676 62.228 97.966 ; 
        RECT 61.688 97.464 61.76 97.902 ; 
        RECT 61.652 94.498 61.724 95.456 ; 
        RECT 61.508 96.822 61.58 97.436 ; 
        RECT 61.184 96.924 61.256 97.956 ; 
        RECT 59.024 94.368 59.096 98.11 ; 
        RECT 58.88 94.368 58.952 98.11 ; 
        RECT 58.736 95.092 58.808 97.364 ; 
        RECT 62.444 98.688 62.516 102.43 ; 
        RECT 62.3 98.688 62.372 102.43 ; 
        RECT 62.156 100.996 62.228 102.286 ; 
        RECT 61.688 101.784 61.76 102.222 ; 
        RECT 61.652 98.818 61.724 99.776 ; 
        RECT 61.508 101.142 61.58 101.756 ; 
        RECT 61.184 101.244 61.256 102.276 ; 
        RECT 59.024 98.688 59.096 102.43 ; 
        RECT 58.88 98.688 58.952 102.43 ; 
        RECT 58.736 99.412 58.808 101.684 ; 
        RECT 62.444 103.008 62.516 106.75 ; 
        RECT 62.3 103.008 62.372 106.75 ; 
        RECT 62.156 105.316 62.228 106.606 ; 
        RECT 61.688 106.104 61.76 106.542 ; 
        RECT 61.652 103.138 61.724 104.096 ; 
        RECT 61.508 105.462 61.58 106.076 ; 
        RECT 61.184 105.564 61.256 106.596 ; 
        RECT 59.024 103.008 59.096 106.75 ; 
        RECT 58.88 103.008 58.952 106.75 ; 
        RECT 58.736 103.732 58.808 106.004 ; 
        RECT 62.444 107.328 62.516 111.07 ; 
        RECT 62.3 107.328 62.372 111.07 ; 
        RECT 62.156 109.636 62.228 110.926 ; 
        RECT 61.688 110.424 61.76 110.862 ; 
        RECT 61.652 107.458 61.724 108.416 ; 
        RECT 61.508 109.782 61.58 110.396 ; 
        RECT 61.184 109.884 61.256 110.916 ; 
        RECT 59.024 107.328 59.096 111.07 ; 
        RECT 58.88 107.328 58.952 111.07 ; 
        RECT 58.736 108.052 58.808 110.324 ; 
  LAYER M3 SPACING 0.072 ; 
      RECT 62.212 1.026 62.724 5.4 ; 
      RECT 62.156 3.688 62.724 4.978 ; 
      RECT 61.276 2.596 61.812 5.4 ; 
      RECT 61.184 3.936 61.812 4.968 ; 
      RECT 61.276 1.026 61.668 5.4 ; 
      RECT 61.276 1.51 61.724 2.468 ; 
      RECT 61.276 1.026 61.812 1.382 ; 
      RECT 60.376 2.828 60.912 5.4 ; 
      RECT 60.376 1.026 60.768 5.4 ; 
      RECT 58.708 1.026 59.04 5.4 ; 
      RECT 58.708 1.38 59.096 5.122 ; 
      RECT 121.072 1.026 121.412 5.4 ; 
      RECT 120.496 1.026 120.6 5.4 ; 
      RECT 120.064 1.026 120.168 5.4 ; 
      RECT 119.632 1.026 119.736 5.4 ; 
      RECT 119.2 1.026 119.304 5.4 ; 
      RECT 118.768 1.026 118.872 5.4 ; 
      RECT 118.336 1.026 118.44 5.4 ; 
      RECT 117.904 1.026 118.008 5.4 ; 
      RECT 117.472 1.026 117.576 5.4 ; 
      RECT 117.04 1.026 117.144 5.4 ; 
      RECT 116.608 1.026 116.712 5.4 ; 
      RECT 116.176 1.026 116.28 5.4 ; 
      RECT 115.744 1.026 115.848 5.4 ; 
      RECT 115.312 1.026 115.416 5.4 ; 
      RECT 114.88 1.026 114.984 5.4 ; 
      RECT 114.448 1.026 114.552 5.4 ; 
      RECT 114.016 1.026 114.12 5.4 ; 
      RECT 113.584 1.026 113.688 5.4 ; 
      RECT 113.152 1.026 113.256 5.4 ; 
      RECT 112.72 1.026 112.824 5.4 ; 
      RECT 112.288 1.026 112.392 5.4 ; 
      RECT 111.856 1.026 111.96 5.4 ; 
      RECT 111.424 1.026 111.528 5.4 ; 
      RECT 110.992 1.026 111.096 5.4 ; 
      RECT 110.56 1.026 110.664 5.4 ; 
      RECT 110.128 1.026 110.232 5.4 ; 
      RECT 109.696 1.026 109.8 5.4 ; 
      RECT 109.264 1.026 109.368 5.4 ; 
      RECT 108.832 1.026 108.936 5.4 ; 
      RECT 108.4 1.026 108.504 5.4 ; 
      RECT 107.968 1.026 108.072 5.4 ; 
      RECT 107.536 1.026 107.64 5.4 ; 
      RECT 107.104 1.026 107.208 5.4 ; 
      RECT 106.672 1.026 106.776 5.4 ; 
      RECT 106.24 1.026 106.344 5.4 ; 
      RECT 105.808 1.026 105.912 5.4 ; 
      RECT 105.376 1.026 105.48 5.4 ; 
      RECT 104.944 1.026 105.048 5.4 ; 
      RECT 104.512 1.026 104.616 5.4 ; 
      RECT 104.08 1.026 104.184 5.4 ; 
      RECT 103.648 1.026 103.752 5.4 ; 
      RECT 103.216 1.026 103.32 5.4 ; 
      RECT 102.784 1.026 102.888 5.4 ; 
      RECT 102.352 1.026 102.456 5.4 ; 
      RECT 101.92 1.026 102.024 5.4 ; 
      RECT 101.488 1.026 101.592 5.4 ; 
      RECT 101.056 1.026 101.16 5.4 ; 
      RECT 100.624 1.026 100.728 5.4 ; 
      RECT 100.192 1.026 100.296 5.4 ; 
      RECT 99.76 1.026 99.864 5.4 ; 
      RECT 99.328 1.026 99.432 5.4 ; 
      RECT 98.896 1.026 99 5.4 ; 
      RECT 98.464 1.026 98.568 5.4 ; 
      RECT 98.032 1.026 98.136 5.4 ; 
      RECT 97.6 1.026 97.704 5.4 ; 
      RECT 97.168 1.026 97.272 5.4 ; 
      RECT 96.736 1.026 96.84 5.4 ; 
      RECT 96.304 1.026 96.408 5.4 ; 
      RECT 95.872 1.026 95.976 5.4 ; 
      RECT 95.44 1.026 95.544 5.4 ; 
      RECT 95.008 1.026 95.112 5.4 ; 
      RECT 94.576 1.026 94.68 5.4 ; 
      RECT 94.144 1.026 94.248 5.4 ; 
      RECT 93.712 1.026 93.816 5.4 ; 
      RECT 93.28 1.026 93.384 5.4 ; 
      RECT 92.848 1.026 92.952 5.4 ; 
      RECT 92.416 1.026 92.52 5.4 ; 
      RECT 91.984 1.026 92.088 5.4 ; 
      RECT 91.552 1.026 91.656 5.4 ; 
      RECT 91.12 1.026 91.224 5.4 ; 
      RECT 90.688 1.026 90.792 5.4 ; 
      RECT 90.256 1.026 90.36 5.4 ; 
      RECT 89.824 1.026 89.928 5.4 ; 
      RECT 89.392 1.026 89.496 5.4 ; 
      RECT 88.96 1.026 89.064 5.4 ; 
      RECT 88.528 1.026 88.632 5.4 ; 
      RECT 88.096 1.026 88.2 5.4 ; 
      RECT 87.664 1.026 87.768 5.4 ; 
      RECT 87.232 1.026 87.336 5.4 ; 
      RECT 86.8 1.026 86.904 5.4 ; 
      RECT 86.368 1.026 86.472 5.4 ; 
      RECT 85.936 1.026 86.04 5.4 ; 
      RECT 85.504 1.026 85.608 5.4 ; 
      RECT 85.072 1.026 85.176 5.4 ; 
      RECT 84.64 1.026 84.744 5.4 ; 
      RECT 84.208 1.026 84.312 5.4 ; 
      RECT 83.776 1.026 83.88 5.4 ; 
      RECT 83.344 1.026 83.448 5.4 ; 
      RECT 82.912 1.026 83.016 5.4 ; 
      RECT 82.48 1.026 82.584 5.4 ; 
      RECT 82.048 1.026 82.152 5.4 ; 
      RECT 81.616 1.026 81.72 5.4 ; 
      RECT 81.184 1.026 81.288 5.4 ; 
      RECT 80.752 1.026 80.856 5.4 ; 
      RECT 80.32 1.026 80.424 5.4 ; 
      RECT 79.888 1.026 79.992 5.4 ; 
      RECT 79.456 1.026 79.56 5.4 ; 
      RECT 79.024 1.026 79.128 5.4 ; 
      RECT 78.592 1.026 78.696 5.4 ; 
      RECT 78.16 1.026 78.264 5.4 ; 
      RECT 77.728 1.026 77.832 5.4 ; 
      RECT 77.296 1.026 77.4 5.4 ; 
      RECT 76.864 1.026 76.968 5.4 ; 
      RECT 76.432 1.026 76.536 5.4 ; 
      RECT 76 1.026 76.104 5.4 ; 
      RECT 75.568 1.026 75.672 5.4 ; 
      RECT 75.136 1.026 75.24 5.4 ; 
      RECT 74.704 1.026 74.808 5.4 ; 
      RECT 74.272 1.026 74.376 5.4 ; 
      RECT 73.84 1.026 73.944 5.4 ; 
      RECT 73.408 1.026 73.512 5.4 ; 
      RECT 72.976 1.026 73.08 5.4 ; 
      RECT 72.544 1.026 72.648 5.4 ; 
      RECT 72.112 1.026 72.216 5.4 ; 
      RECT 71.68 1.026 71.784 5.4 ; 
      RECT 71.248 1.026 71.352 5.4 ; 
      RECT 70.816 1.026 70.92 5.4 ; 
      RECT 70.384 1.026 70.488 5.4 ; 
      RECT 69.952 1.026 70.056 5.4 ; 
      RECT 69.52 1.026 69.624 5.4 ; 
      RECT 69.088 1.026 69.192 5.4 ; 
      RECT 68.656 1.026 68.76 5.4 ; 
      RECT 68.224 1.026 68.328 5.4 ; 
      RECT 67.792 1.026 67.896 5.4 ; 
      RECT 67.36 1.026 67.464 5.4 ; 
      RECT 66.928 1.026 67.032 5.4 ; 
      RECT 66.496 1.026 66.6 5.4 ; 
      RECT 66.064 1.026 66.168 5.4 ; 
      RECT 65.632 1.026 65.736 5.4 ; 
      RECT 65.2 1.026 65.304 5.4 ; 
      RECT 64.348 1.026 64.656 5.4 ; 
      RECT 56.776 1.026 57.084 5.4 ; 
      RECT 56.128 1.026 56.232 5.4 ; 
      RECT 55.696 1.026 55.8 5.4 ; 
      RECT 55.264 1.026 55.368 5.4 ; 
      RECT 54.832 1.026 54.936 5.4 ; 
      RECT 54.4 1.026 54.504 5.4 ; 
      RECT 53.968 1.026 54.072 5.4 ; 
      RECT 53.536 1.026 53.64 5.4 ; 
      RECT 53.104 1.026 53.208 5.4 ; 
      RECT 52.672 1.026 52.776 5.4 ; 
      RECT 52.24 1.026 52.344 5.4 ; 
      RECT 51.808 1.026 51.912 5.4 ; 
      RECT 51.376 1.026 51.48 5.4 ; 
      RECT 50.944 1.026 51.048 5.4 ; 
      RECT 50.512 1.026 50.616 5.4 ; 
      RECT 50.08 1.026 50.184 5.4 ; 
      RECT 49.648 1.026 49.752 5.4 ; 
      RECT 49.216 1.026 49.32 5.4 ; 
      RECT 48.784 1.026 48.888 5.4 ; 
      RECT 48.352 1.026 48.456 5.4 ; 
      RECT 47.92 1.026 48.024 5.4 ; 
      RECT 47.488 1.026 47.592 5.4 ; 
      RECT 47.056 1.026 47.16 5.4 ; 
      RECT 46.624 1.026 46.728 5.4 ; 
      RECT 46.192 1.026 46.296 5.4 ; 
      RECT 45.76 1.026 45.864 5.4 ; 
      RECT 45.328 1.026 45.432 5.4 ; 
      RECT 44.896 1.026 45 5.4 ; 
      RECT 44.464 1.026 44.568 5.4 ; 
      RECT 44.032 1.026 44.136 5.4 ; 
      RECT 43.6 1.026 43.704 5.4 ; 
      RECT 43.168 1.026 43.272 5.4 ; 
      RECT 42.736 1.026 42.84 5.4 ; 
      RECT 42.304 1.026 42.408 5.4 ; 
      RECT 41.872 1.026 41.976 5.4 ; 
      RECT 41.44 1.026 41.544 5.4 ; 
      RECT 41.008 1.026 41.112 5.4 ; 
      RECT 40.576 1.026 40.68 5.4 ; 
      RECT 40.144 1.026 40.248 5.4 ; 
      RECT 39.712 1.026 39.816 5.4 ; 
      RECT 39.28 1.026 39.384 5.4 ; 
      RECT 38.848 1.026 38.952 5.4 ; 
      RECT 38.416 1.026 38.52 5.4 ; 
      RECT 37.984 1.026 38.088 5.4 ; 
      RECT 37.552 1.026 37.656 5.4 ; 
      RECT 37.12 1.026 37.224 5.4 ; 
      RECT 36.688 1.026 36.792 5.4 ; 
      RECT 36.256 1.026 36.36 5.4 ; 
      RECT 35.824 1.026 35.928 5.4 ; 
      RECT 35.392 1.026 35.496 5.4 ; 
      RECT 34.96 1.026 35.064 5.4 ; 
      RECT 34.528 1.026 34.632 5.4 ; 
      RECT 34.096 1.026 34.2 5.4 ; 
      RECT 33.664 1.026 33.768 5.4 ; 
      RECT 33.232 1.026 33.336 5.4 ; 
      RECT 32.8 1.026 32.904 5.4 ; 
      RECT 32.368 1.026 32.472 5.4 ; 
      RECT 31.936 1.026 32.04 5.4 ; 
      RECT 31.504 1.026 31.608 5.4 ; 
      RECT 31.072 1.026 31.176 5.4 ; 
      RECT 30.64 1.026 30.744 5.4 ; 
      RECT 30.208 1.026 30.312 5.4 ; 
      RECT 29.776 1.026 29.88 5.4 ; 
      RECT 29.344 1.026 29.448 5.4 ; 
      RECT 28.912 1.026 29.016 5.4 ; 
      RECT 28.48 1.026 28.584 5.4 ; 
      RECT 28.048 1.026 28.152 5.4 ; 
      RECT 27.616 1.026 27.72 5.4 ; 
      RECT 27.184 1.026 27.288 5.4 ; 
      RECT 26.752 1.026 26.856 5.4 ; 
      RECT 26.32 1.026 26.424 5.4 ; 
      RECT 25.888 1.026 25.992 5.4 ; 
      RECT 25.456 1.026 25.56 5.4 ; 
      RECT 25.024 1.026 25.128 5.4 ; 
      RECT 24.592 1.026 24.696 5.4 ; 
      RECT 24.16 1.026 24.264 5.4 ; 
      RECT 23.728 1.026 23.832 5.4 ; 
      RECT 23.296 1.026 23.4 5.4 ; 
      RECT 22.864 1.026 22.968 5.4 ; 
      RECT 22.432 1.026 22.536 5.4 ; 
      RECT 22 1.026 22.104 5.4 ; 
      RECT 21.568 1.026 21.672 5.4 ; 
      RECT 21.136 1.026 21.24 5.4 ; 
      RECT 20.704 1.026 20.808 5.4 ; 
      RECT 20.272 1.026 20.376 5.4 ; 
      RECT 19.84 1.026 19.944 5.4 ; 
      RECT 19.408 1.026 19.512 5.4 ; 
      RECT 18.976 1.026 19.08 5.4 ; 
      RECT 18.544 1.026 18.648 5.4 ; 
      RECT 18.112 1.026 18.216 5.4 ; 
      RECT 17.68 1.026 17.784 5.4 ; 
      RECT 17.248 1.026 17.352 5.4 ; 
      RECT 16.816 1.026 16.92 5.4 ; 
      RECT 16.384 1.026 16.488 5.4 ; 
      RECT 15.952 1.026 16.056 5.4 ; 
      RECT 15.52 1.026 15.624 5.4 ; 
      RECT 15.088 1.026 15.192 5.4 ; 
      RECT 14.656 1.026 14.76 5.4 ; 
      RECT 14.224 1.026 14.328 5.4 ; 
      RECT 13.792 1.026 13.896 5.4 ; 
      RECT 13.36 1.026 13.464 5.4 ; 
      RECT 12.928 1.026 13.032 5.4 ; 
      RECT 12.496 1.026 12.6 5.4 ; 
      RECT 12.064 1.026 12.168 5.4 ; 
      RECT 11.632 1.026 11.736 5.4 ; 
      RECT 11.2 1.026 11.304 5.4 ; 
      RECT 10.768 1.026 10.872 5.4 ; 
      RECT 10.336 1.026 10.44 5.4 ; 
      RECT 9.904 1.026 10.008 5.4 ; 
      RECT 9.472 1.026 9.576 5.4 ; 
      RECT 9.04 1.026 9.144 5.4 ; 
      RECT 8.608 1.026 8.712 5.4 ; 
      RECT 8.176 1.026 8.28 5.4 ; 
      RECT 7.744 1.026 7.848 5.4 ; 
      RECT 7.312 1.026 7.416 5.4 ; 
      RECT 6.88 1.026 6.984 5.4 ; 
      RECT 6.448 1.026 6.552 5.4 ; 
      RECT 6.016 1.026 6.12 5.4 ; 
      RECT 5.584 1.026 5.688 5.4 ; 
      RECT 5.152 1.026 5.256 5.4 ; 
      RECT 4.72 1.026 4.824 5.4 ; 
      RECT 4.288 1.026 4.392 5.4 ; 
      RECT 3.856 1.026 3.96 5.4 ; 
      RECT 3.424 1.026 3.528 5.4 ; 
      RECT 2.992 1.026 3.096 5.4 ; 
      RECT 2.56 1.026 2.664 5.4 ; 
      RECT 2.128 1.026 2.232 5.4 ; 
      RECT 1.696 1.026 1.8 5.4 ; 
      RECT 1.264 1.026 1.368 5.4 ; 
      RECT 0.832 1.026 0.936 5.4 ; 
      RECT 0.02 1.026 0.36 5.4 ; 
      RECT 62.212 5.346 62.724 9.72 ; 
      RECT 62.156 8.008 62.724 9.298 ; 
      RECT 61.276 6.916 61.812 9.72 ; 
      RECT 61.184 8.256 61.812 9.288 ; 
      RECT 61.276 5.346 61.668 9.72 ; 
      RECT 61.276 5.83 61.724 6.788 ; 
      RECT 61.276 5.346 61.812 5.702 ; 
      RECT 60.376 7.148 60.912 9.72 ; 
      RECT 60.376 5.346 60.768 9.72 ; 
      RECT 58.708 5.346 59.04 9.72 ; 
      RECT 58.708 5.7 59.096 9.442 ; 
      RECT 121.072 5.346 121.412 9.72 ; 
      RECT 120.496 5.346 120.6 9.72 ; 
      RECT 120.064 5.346 120.168 9.72 ; 
      RECT 119.632 5.346 119.736 9.72 ; 
      RECT 119.2 5.346 119.304 9.72 ; 
      RECT 118.768 5.346 118.872 9.72 ; 
      RECT 118.336 5.346 118.44 9.72 ; 
      RECT 117.904 5.346 118.008 9.72 ; 
      RECT 117.472 5.346 117.576 9.72 ; 
      RECT 117.04 5.346 117.144 9.72 ; 
      RECT 116.608 5.346 116.712 9.72 ; 
      RECT 116.176 5.346 116.28 9.72 ; 
      RECT 115.744 5.346 115.848 9.72 ; 
      RECT 115.312 5.346 115.416 9.72 ; 
      RECT 114.88 5.346 114.984 9.72 ; 
      RECT 114.448 5.346 114.552 9.72 ; 
      RECT 114.016 5.346 114.12 9.72 ; 
      RECT 113.584 5.346 113.688 9.72 ; 
      RECT 113.152 5.346 113.256 9.72 ; 
      RECT 112.72 5.346 112.824 9.72 ; 
      RECT 112.288 5.346 112.392 9.72 ; 
      RECT 111.856 5.346 111.96 9.72 ; 
      RECT 111.424 5.346 111.528 9.72 ; 
      RECT 110.992 5.346 111.096 9.72 ; 
      RECT 110.56 5.346 110.664 9.72 ; 
      RECT 110.128 5.346 110.232 9.72 ; 
      RECT 109.696 5.346 109.8 9.72 ; 
      RECT 109.264 5.346 109.368 9.72 ; 
      RECT 108.832 5.346 108.936 9.72 ; 
      RECT 108.4 5.346 108.504 9.72 ; 
      RECT 107.968 5.346 108.072 9.72 ; 
      RECT 107.536 5.346 107.64 9.72 ; 
      RECT 107.104 5.346 107.208 9.72 ; 
      RECT 106.672 5.346 106.776 9.72 ; 
      RECT 106.24 5.346 106.344 9.72 ; 
      RECT 105.808 5.346 105.912 9.72 ; 
      RECT 105.376 5.346 105.48 9.72 ; 
      RECT 104.944 5.346 105.048 9.72 ; 
      RECT 104.512 5.346 104.616 9.72 ; 
      RECT 104.08 5.346 104.184 9.72 ; 
      RECT 103.648 5.346 103.752 9.72 ; 
      RECT 103.216 5.346 103.32 9.72 ; 
      RECT 102.784 5.346 102.888 9.72 ; 
      RECT 102.352 5.346 102.456 9.72 ; 
      RECT 101.92 5.346 102.024 9.72 ; 
      RECT 101.488 5.346 101.592 9.72 ; 
      RECT 101.056 5.346 101.16 9.72 ; 
      RECT 100.624 5.346 100.728 9.72 ; 
      RECT 100.192 5.346 100.296 9.72 ; 
      RECT 99.76 5.346 99.864 9.72 ; 
      RECT 99.328 5.346 99.432 9.72 ; 
      RECT 98.896 5.346 99 9.72 ; 
      RECT 98.464 5.346 98.568 9.72 ; 
      RECT 98.032 5.346 98.136 9.72 ; 
      RECT 97.6 5.346 97.704 9.72 ; 
      RECT 97.168 5.346 97.272 9.72 ; 
      RECT 96.736 5.346 96.84 9.72 ; 
      RECT 96.304 5.346 96.408 9.72 ; 
      RECT 95.872 5.346 95.976 9.72 ; 
      RECT 95.44 5.346 95.544 9.72 ; 
      RECT 95.008 5.346 95.112 9.72 ; 
      RECT 94.576 5.346 94.68 9.72 ; 
      RECT 94.144 5.346 94.248 9.72 ; 
      RECT 93.712 5.346 93.816 9.72 ; 
      RECT 93.28 5.346 93.384 9.72 ; 
      RECT 92.848 5.346 92.952 9.72 ; 
      RECT 92.416 5.346 92.52 9.72 ; 
      RECT 91.984 5.346 92.088 9.72 ; 
      RECT 91.552 5.346 91.656 9.72 ; 
      RECT 91.12 5.346 91.224 9.72 ; 
      RECT 90.688 5.346 90.792 9.72 ; 
      RECT 90.256 5.346 90.36 9.72 ; 
      RECT 89.824 5.346 89.928 9.72 ; 
      RECT 89.392 5.346 89.496 9.72 ; 
      RECT 88.96 5.346 89.064 9.72 ; 
      RECT 88.528 5.346 88.632 9.72 ; 
      RECT 88.096 5.346 88.2 9.72 ; 
      RECT 87.664 5.346 87.768 9.72 ; 
      RECT 87.232 5.346 87.336 9.72 ; 
      RECT 86.8 5.346 86.904 9.72 ; 
      RECT 86.368 5.346 86.472 9.72 ; 
      RECT 85.936 5.346 86.04 9.72 ; 
      RECT 85.504 5.346 85.608 9.72 ; 
      RECT 85.072 5.346 85.176 9.72 ; 
      RECT 84.64 5.346 84.744 9.72 ; 
      RECT 84.208 5.346 84.312 9.72 ; 
      RECT 83.776 5.346 83.88 9.72 ; 
      RECT 83.344 5.346 83.448 9.72 ; 
      RECT 82.912 5.346 83.016 9.72 ; 
      RECT 82.48 5.346 82.584 9.72 ; 
      RECT 82.048 5.346 82.152 9.72 ; 
      RECT 81.616 5.346 81.72 9.72 ; 
      RECT 81.184 5.346 81.288 9.72 ; 
      RECT 80.752 5.346 80.856 9.72 ; 
      RECT 80.32 5.346 80.424 9.72 ; 
      RECT 79.888 5.346 79.992 9.72 ; 
      RECT 79.456 5.346 79.56 9.72 ; 
      RECT 79.024 5.346 79.128 9.72 ; 
      RECT 78.592 5.346 78.696 9.72 ; 
      RECT 78.16 5.346 78.264 9.72 ; 
      RECT 77.728 5.346 77.832 9.72 ; 
      RECT 77.296 5.346 77.4 9.72 ; 
      RECT 76.864 5.346 76.968 9.72 ; 
      RECT 76.432 5.346 76.536 9.72 ; 
      RECT 76 5.346 76.104 9.72 ; 
      RECT 75.568 5.346 75.672 9.72 ; 
      RECT 75.136 5.346 75.24 9.72 ; 
      RECT 74.704 5.346 74.808 9.72 ; 
      RECT 74.272 5.346 74.376 9.72 ; 
      RECT 73.84 5.346 73.944 9.72 ; 
      RECT 73.408 5.346 73.512 9.72 ; 
      RECT 72.976 5.346 73.08 9.72 ; 
      RECT 72.544 5.346 72.648 9.72 ; 
      RECT 72.112 5.346 72.216 9.72 ; 
      RECT 71.68 5.346 71.784 9.72 ; 
      RECT 71.248 5.346 71.352 9.72 ; 
      RECT 70.816 5.346 70.92 9.72 ; 
      RECT 70.384 5.346 70.488 9.72 ; 
      RECT 69.952 5.346 70.056 9.72 ; 
      RECT 69.52 5.346 69.624 9.72 ; 
      RECT 69.088 5.346 69.192 9.72 ; 
      RECT 68.656 5.346 68.76 9.72 ; 
      RECT 68.224 5.346 68.328 9.72 ; 
      RECT 67.792 5.346 67.896 9.72 ; 
      RECT 67.36 5.346 67.464 9.72 ; 
      RECT 66.928 5.346 67.032 9.72 ; 
      RECT 66.496 5.346 66.6 9.72 ; 
      RECT 66.064 5.346 66.168 9.72 ; 
      RECT 65.632 5.346 65.736 9.72 ; 
      RECT 65.2 5.346 65.304 9.72 ; 
      RECT 64.348 5.346 64.656 9.72 ; 
      RECT 56.776 5.346 57.084 9.72 ; 
      RECT 56.128 5.346 56.232 9.72 ; 
      RECT 55.696 5.346 55.8 9.72 ; 
      RECT 55.264 5.346 55.368 9.72 ; 
      RECT 54.832 5.346 54.936 9.72 ; 
      RECT 54.4 5.346 54.504 9.72 ; 
      RECT 53.968 5.346 54.072 9.72 ; 
      RECT 53.536 5.346 53.64 9.72 ; 
      RECT 53.104 5.346 53.208 9.72 ; 
      RECT 52.672 5.346 52.776 9.72 ; 
      RECT 52.24 5.346 52.344 9.72 ; 
      RECT 51.808 5.346 51.912 9.72 ; 
      RECT 51.376 5.346 51.48 9.72 ; 
      RECT 50.944 5.346 51.048 9.72 ; 
      RECT 50.512 5.346 50.616 9.72 ; 
      RECT 50.08 5.346 50.184 9.72 ; 
      RECT 49.648 5.346 49.752 9.72 ; 
      RECT 49.216 5.346 49.32 9.72 ; 
      RECT 48.784 5.346 48.888 9.72 ; 
      RECT 48.352 5.346 48.456 9.72 ; 
      RECT 47.92 5.346 48.024 9.72 ; 
      RECT 47.488 5.346 47.592 9.72 ; 
      RECT 47.056 5.346 47.16 9.72 ; 
      RECT 46.624 5.346 46.728 9.72 ; 
      RECT 46.192 5.346 46.296 9.72 ; 
      RECT 45.76 5.346 45.864 9.72 ; 
      RECT 45.328 5.346 45.432 9.72 ; 
      RECT 44.896 5.346 45 9.72 ; 
      RECT 44.464 5.346 44.568 9.72 ; 
      RECT 44.032 5.346 44.136 9.72 ; 
      RECT 43.6 5.346 43.704 9.72 ; 
      RECT 43.168 5.346 43.272 9.72 ; 
      RECT 42.736 5.346 42.84 9.72 ; 
      RECT 42.304 5.346 42.408 9.72 ; 
      RECT 41.872 5.346 41.976 9.72 ; 
      RECT 41.44 5.346 41.544 9.72 ; 
      RECT 41.008 5.346 41.112 9.72 ; 
      RECT 40.576 5.346 40.68 9.72 ; 
      RECT 40.144 5.346 40.248 9.72 ; 
      RECT 39.712 5.346 39.816 9.72 ; 
      RECT 39.28 5.346 39.384 9.72 ; 
      RECT 38.848 5.346 38.952 9.72 ; 
      RECT 38.416 5.346 38.52 9.72 ; 
      RECT 37.984 5.346 38.088 9.72 ; 
      RECT 37.552 5.346 37.656 9.72 ; 
      RECT 37.12 5.346 37.224 9.72 ; 
      RECT 36.688 5.346 36.792 9.72 ; 
      RECT 36.256 5.346 36.36 9.72 ; 
      RECT 35.824 5.346 35.928 9.72 ; 
      RECT 35.392 5.346 35.496 9.72 ; 
      RECT 34.96 5.346 35.064 9.72 ; 
      RECT 34.528 5.346 34.632 9.72 ; 
      RECT 34.096 5.346 34.2 9.72 ; 
      RECT 33.664 5.346 33.768 9.72 ; 
      RECT 33.232 5.346 33.336 9.72 ; 
      RECT 32.8 5.346 32.904 9.72 ; 
      RECT 32.368 5.346 32.472 9.72 ; 
      RECT 31.936 5.346 32.04 9.72 ; 
      RECT 31.504 5.346 31.608 9.72 ; 
      RECT 31.072 5.346 31.176 9.72 ; 
      RECT 30.64 5.346 30.744 9.72 ; 
      RECT 30.208 5.346 30.312 9.72 ; 
      RECT 29.776 5.346 29.88 9.72 ; 
      RECT 29.344 5.346 29.448 9.72 ; 
      RECT 28.912 5.346 29.016 9.72 ; 
      RECT 28.48 5.346 28.584 9.72 ; 
      RECT 28.048 5.346 28.152 9.72 ; 
      RECT 27.616 5.346 27.72 9.72 ; 
      RECT 27.184 5.346 27.288 9.72 ; 
      RECT 26.752 5.346 26.856 9.72 ; 
      RECT 26.32 5.346 26.424 9.72 ; 
      RECT 25.888 5.346 25.992 9.72 ; 
      RECT 25.456 5.346 25.56 9.72 ; 
      RECT 25.024 5.346 25.128 9.72 ; 
      RECT 24.592 5.346 24.696 9.72 ; 
      RECT 24.16 5.346 24.264 9.72 ; 
      RECT 23.728 5.346 23.832 9.72 ; 
      RECT 23.296 5.346 23.4 9.72 ; 
      RECT 22.864 5.346 22.968 9.72 ; 
      RECT 22.432 5.346 22.536 9.72 ; 
      RECT 22 5.346 22.104 9.72 ; 
      RECT 21.568 5.346 21.672 9.72 ; 
      RECT 21.136 5.346 21.24 9.72 ; 
      RECT 20.704 5.346 20.808 9.72 ; 
      RECT 20.272 5.346 20.376 9.72 ; 
      RECT 19.84 5.346 19.944 9.72 ; 
      RECT 19.408 5.346 19.512 9.72 ; 
      RECT 18.976 5.346 19.08 9.72 ; 
      RECT 18.544 5.346 18.648 9.72 ; 
      RECT 18.112 5.346 18.216 9.72 ; 
      RECT 17.68 5.346 17.784 9.72 ; 
      RECT 17.248 5.346 17.352 9.72 ; 
      RECT 16.816 5.346 16.92 9.72 ; 
      RECT 16.384 5.346 16.488 9.72 ; 
      RECT 15.952 5.346 16.056 9.72 ; 
      RECT 15.52 5.346 15.624 9.72 ; 
      RECT 15.088 5.346 15.192 9.72 ; 
      RECT 14.656 5.346 14.76 9.72 ; 
      RECT 14.224 5.346 14.328 9.72 ; 
      RECT 13.792 5.346 13.896 9.72 ; 
      RECT 13.36 5.346 13.464 9.72 ; 
      RECT 12.928 5.346 13.032 9.72 ; 
      RECT 12.496 5.346 12.6 9.72 ; 
      RECT 12.064 5.346 12.168 9.72 ; 
      RECT 11.632 5.346 11.736 9.72 ; 
      RECT 11.2 5.346 11.304 9.72 ; 
      RECT 10.768 5.346 10.872 9.72 ; 
      RECT 10.336 5.346 10.44 9.72 ; 
      RECT 9.904 5.346 10.008 9.72 ; 
      RECT 9.472 5.346 9.576 9.72 ; 
      RECT 9.04 5.346 9.144 9.72 ; 
      RECT 8.608 5.346 8.712 9.72 ; 
      RECT 8.176 5.346 8.28 9.72 ; 
      RECT 7.744 5.346 7.848 9.72 ; 
      RECT 7.312 5.346 7.416 9.72 ; 
      RECT 6.88 5.346 6.984 9.72 ; 
      RECT 6.448 5.346 6.552 9.72 ; 
      RECT 6.016 5.346 6.12 9.72 ; 
      RECT 5.584 5.346 5.688 9.72 ; 
      RECT 5.152 5.346 5.256 9.72 ; 
      RECT 4.72 5.346 4.824 9.72 ; 
      RECT 4.288 5.346 4.392 9.72 ; 
      RECT 3.856 5.346 3.96 9.72 ; 
      RECT 3.424 5.346 3.528 9.72 ; 
      RECT 2.992 5.346 3.096 9.72 ; 
      RECT 2.56 5.346 2.664 9.72 ; 
      RECT 2.128 5.346 2.232 9.72 ; 
      RECT 1.696 5.346 1.8 9.72 ; 
      RECT 1.264 5.346 1.368 9.72 ; 
      RECT 0.832 5.346 0.936 9.72 ; 
      RECT 0.02 5.346 0.36 9.72 ; 
      RECT 62.212 9.666 62.724 14.04 ; 
      RECT 62.156 12.328 62.724 13.618 ; 
      RECT 61.276 11.236 61.812 14.04 ; 
      RECT 61.184 12.576 61.812 13.608 ; 
      RECT 61.276 9.666 61.668 14.04 ; 
      RECT 61.276 10.15 61.724 11.108 ; 
      RECT 61.276 9.666 61.812 10.022 ; 
      RECT 60.376 11.468 60.912 14.04 ; 
      RECT 60.376 9.666 60.768 14.04 ; 
      RECT 58.708 9.666 59.04 14.04 ; 
      RECT 58.708 10.02 59.096 13.762 ; 
      RECT 121.072 9.666 121.412 14.04 ; 
      RECT 120.496 9.666 120.6 14.04 ; 
      RECT 120.064 9.666 120.168 14.04 ; 
      RECT 119.632 9.666 119.736 14.04 ; 
      RECT 119.2 9.666 119.304 14.04 ; 
      RECT 118.768 9.666 118.872 14.04 ; 
      RECT 118.336 9.666 118.44 14.04 ; 
      RECT 117.904 9.666 118.008 14.04 ; 
      RECT 117.472 9.666 117.576 14.04 ; 
      RECT 117.04 9.666 117.144 14.04 ; 
      RECT 116.608 9.666 116.712 14.04 ; 
      RECT 116.176 9.666 116.28 14.04 ; 
      RECT 115.744 9.666 115.848 14.04 ; 
      RECT 115.312 9.666 115.416 14.04 ; 
      RECT 114.88 9.666 114.984 14.04 ; 
      RECT 114.448 9.666 114.552 14.04 ; 
      RECT 114.016 9.666 114.12 14.04 ; 
      RECT 113.584 9.666 113.688 14.04 ; 
      RECT 113.152 9.666 113.256 14.04 ; 
      RECT 112.72 9.666 112.824 14.04 ; 
      RECT 112.288 9.666 112.392 14.04 ; 
      RECT 111.856 9.666 111.96 14.04 ; 
      RECT 111.424 9.666 111.528 14.04 ; 
      RECT 110.992 9.666 111.096 14.04 ; 
      RECT 110.56 9.666 110.664 14.04 ; 
      RECT 110.128 9.666 110.232 14.04 ; 
      RECT 109.696 9.666 109.8 14.04 ; 
      RECT 109.264 9.666 109.368 14.04 ; 
      RECT 108.832 9.666 108.936 14.04 ; 
      RECT 108.4 9.666 108.504 14.04 ; 
      RECT 107.968 9.666 108.072 14.04 ; 
      RECT 107.536 9.666 107.64 14.04 ; 
      RECT 107.104 9.666 107.208 14.04 ; 
      RECT 106.672 9.666 106.776 14.04 ; 
      RECT 106.24 9.666 106.344 14.04 ; 
      RECT 105.808 9.666 105.912 14.04 ; 
      RECT 105.376 9.666 105.48 14.04 ; 
      RECT 104.944 9.666 105.048 14.04 ; 
      RECT 104.512 9.666 104.616 14.04 ; 
      RECT 104.08 9.666 104.184 14.04 ; 
      RECT 103.648 9.666 103.752 14.04 ; 
      RECT 103.216 9.666 103.32 14.04 ; 
      RECT 102.784 9.666 102.888 14.04 ; 
      RECT 102.352 9.666 102.456 14.04 ; 
      RECT 101.92 9.666 102.024 14.04 ; 
      RECT 101.488 9.666 101.592 14.04 ; 
      RECT 101.056 9.666 101.16 14.04 ; 
      RECT 100.624 9.666 100.728 14.04 ; 
      RECT 100.192 9.666 100.296 14.04 ; 
      RECT 99.76 9.666 99.864 14.04 ; 
      RECT 99.328 9.666 99.432 14.04 ; 
      RECT 98.896 9.666 99 14.04 ; 
      RECT 98.464 9.666 98.568 14.04 ; 
      RECT 98.032 9.666 98.136 14.04 ; 
      RECT 97.6 9.666 97.704 14.04 ; 
      RECT 97.168 9.666 97.272 14.04 ; 
      RECT 96.736 9.666 96.84 14.04 ; 
      RECT 96.304 9.666 96.408 14.04 ; 
      RECT 95.872 9.666 95.976 14.04 ; 
      RECT 95.44 9.666 95.544 14.04 ; 
      RECT 95.008 9.666 95.112 14.04 ; 
      RECT 94.576 9.666 94.68 14.04 ; 
      RECT 94.144 9.666 94.248 14.04 ; 
      RECT 93.712 9.666 93.816 14.04 ; 
      RECT 93.28 9.666 93.384 14.04 ; 
      RECT 92.848 9.666 92.952 14.04 ; 
      RECT 92.416 9.666 92.52 14.04 ; 
      RECT 91.984 9.666 92.088 14.04 ; 
      RECT 91.552 9.666 91.656 14.04 ; 
      RECT 91.12 9.666 91.224 14.04 ; 
      RECT 90.688 9.666 90.792 14.04 ; 
      RECT 90.256 9.666 90.36 14.04 ; 
      RECT 89.824 9.666 89.928 14.04 ; 
      RECT 89.392 9.666 89.496 14.04 ; 
      RECT 88.96 9.666 89.064 14.04 ; 
      RECT 88.528 9.666 88.632 14.04 ; 
      RECT 88.096 9.666 88.2 14.04 ; 
      RECT 87.664 9.666 87.768 14.04 ; 
      RECT 87.232 9.666 87.336 14.04 ; 
      RECT 86.8 9.666 86.904 14.04 ; 
      RECT 86.368 9.666 86.472 14.04 ; 
      RECT 85.936 9.666 86.04 14.04 ; 
      RECT 85.504 9.666 85.608 14.04 ; 
      RECT 85.072 9.666 85.176 14.04 ; 
      RECT 84.64 9.666 84.744 14.04 ; 
      RECT 84.208 9.666 84.312 14.04 ; 
      RECT 83.776 9.666 83.88 14.04 ; 
      RECT 83.344 9.666 83.448 14.04 ; 
      RECT 82.912 9.666 83.016 14.04 ; 
      RECT 82.48 9.666 82.584 14.04 ; 
      RECT 82.048 9.666 82.152 14.04 ; 
      RECT 81.616 9.666 81.72 14.04 ; 
      RECT 81.184 9.666 81.288 14.04 ; 
      RECT 80.752 9.666 80.856 14.04 ; 
      RECT 80.32 9.666 80.424 14.04 ; 
      RECT 79.888 9.666 79.992 14.04 ; 
      RECT 79.456 9.666 79.56 14.04 ; 
      RECT 79.024 9.666 79.128 14.04 ; 
      RECT 78.592 9.666 78.696 14.04 ; 
      RECT 78.16 9.666 78.264 14.04 ; 
      RECT 77.728 9.666 77.832 14.04 ; 
      RECT 77.296 9.666 77.4 14.04 ; 
      RECT 76.864 9.666 76.968 14.04 ; 
      RECT 76.432 9.666 76.536 14.04 ; 
      RECT 76 9.666 76.104 14.04 ; 
      RECT 75.568 9.666 75.672 14.04 ; 
      RECT 75.136 9.666 75.24 14.04 ; 
      RECT 74.704 9.666 74.808 14.04 ; 
      RECT 74.272 9.666 74.376 14.04 ; 
      RECT 73.84 9.666 73.944 14.04 ; 
      RECT 73.408 9.666 73.512 14.04 ; 
      RECT 72.976 9.666 73.08 14.04 ; 
      RECT 72.544 9.666 72.648 14.04 ; 
      RECT 72.112 9.666 72.216 14.04 ; 
      RECT 71.68 9.666 71.784 14.04 ; 
      RECT 71.248 9.666 71.352 14.04 ; 
      RECT 70.816 9.666 70.92 14.04 ; 
      RECT 70.384 9.666 70.488 14.04 ; 
      RECT 69.952 9.666 70.056 14.04 ; 
      RECT 69.52 9.666 69.624 14.04 ; 
      RECT 69.088 9.666 69.192 14.04 ; 
      RECT 68.656 9.666 68.76 14.04 ; 
      RECT 68.224 9.666 68.328 14.04 ; 
      RECT 67.792 9.666 67.896 14.04 ; 
      RECT 67.36 9.666 67.464 14.04 ; 
      RECT 66.928 9.666 67.032 14.04 ; 
      RECT 66.496 9.666 66.6 14.04 ; 
      RECT 66.064 9.666 66.168 14.04 ; 
      RECT 65.632 9.666 65.736 14.04 ; 
      RECT 65.2 9.666 65.304 14.04 ; 
      RECT 64.348 9.666 64.656 14.04 ; 
      RECT 56.776 9.666 57.084 14.04 ; 
      RECT 56.128 9.666 56.232 14.04 ; 
      RECT 55.696 9.666 55.8 14.04 ; 
      RECT 55.264 9.666 55.368 14.04 ; 
      RECT 54.832 9.666 54.936 14.04 ; 
      RECT 54.4 9.666 54.504 14.04 ; 
      RECT 53.968 9.666 54.072 14.04 ; 
      RECT 53.536 9.666 53.64 14.04 ; 
      RECT 53.104 9.666 53.208 14.04 ; 
      RECT 52.672 9.666 52.776 14.04 ; 
      RECT 52.24 9.666 52.344 14.04 ; 
      RECT 51.808 9.666 51.912 14.04 ; 
      RECT 51.376 9.666 51.48 14.04 ; 
      RECT 50.944 9.666 51.048 14.04 ; 
      RECT 50.512 9.666 50.616 14.04 ; 
      RECT 50.08 9.666 50.184 14.04 ; 
      RECT 49.648 9.666 49.752 14.04 ; 
      RECT 49.216 9.666 49.32 14.04 ; 
      RECT 48.784 9.666 48.888 14.04 ; 
      RECT 48.352 9.666 48.456 14.04 ; 
      RECT 47.92 9.666 48.024 14.04 ; 
      RECT 47.488 9.666 47.592 14.04 ; 
      RECT 47.056 9.666 47.16 14.04 ; 
      RECT 46.624 9.666 46.728 14.04 ; 
      RECT 46.192 9.666 46.296 14.04 ; 
      RECT 45.76 9.666 45.864 14.04 ; 
      RECT 45.328 9.666 45.432 14.04 ; 
      RECT 44.896 9.666 45 14.04 ; 
      RECT 44.464 9.666 44.568 14.04 ; 
      RECT 44.032 9.666 44.136 14.04 ; 
      RECT 43.6 9.666 43.704 14.04 ; 
      RECT 43.168 9.666 43.272 14.04 ; 
      RECT 42.736 9.666 42.84 14.04 ; 
      RECT 42.304 9.666 42.408 14.04 ; 
      RECT 41.872 9.666 41.976 14.04 ; 
      RECT 41.44 9.666 41.544 14.04 ; 
      RECT 41.008 9.666 41.112 14.04 ; 
      RECT 40.576 9.666 40.68 14.04 ; 
      RECT 40.144 9.666 40.248 14.04 ; 
      RECT 39.712 9.666 39.816 14.04 ; 
      RECT 39.28 9.666 39.384 14.04 ; 
      RECT 38.848 9.666 38.952 14.04 ; 
      RECT 38.416 9.666 38.52 14.04 ; 
      RECT 37.984 9.666 38.088 14.04 ; 
      RECT 37.552 9.666 37.656 14.04 ; 
      RECT 37.12 9.666 37.224 14.04 ; 
      RECT 36.688 9.666 36.792 14.04 ; 
      RECT 36.256 9.666 36.36 14.04 ; 
      RECT 35.824 9.666 35.928 14.04 ; 
      RECT 35.392 9.666 35.496 14.04 ; 
      RECT 34.96 9.666 35.064 14.04 ; 
      RECT 34.528 9.666 34.632 14.04 ; 
      RECT 34.096 9.666 34.2 14.04 ; 
      RECT 33.664 9.666 33.768 14.04 ; 
      RECT 33.232 9.666 33.336 14.04 ; 
      RECT 32.8 9.666 32.904 14.04 ; 
      RECT 32.368 9.666 32.472 14.04 ; 
      RECT 31.936 9.666 32.04 14.04 ; 
      RECT 31.504 9.666 31.608 14.04 ; 
      RECT 31.072 9.666 31.176 14.04 ; 
      RECT 30.64 9.666 30.744 14.04 ; 
      RECT 30.208 9.666 30.312 14.04 ; 
      RECT 29.776 9.666 29.88 14.04 ; 
      RECT 29.344 9.666 29.448 14.04 ; 
      RECT 28.912 9.666 29.016 14.04 ; 
      RECT 28.48 9.666 28.584 14.04 ; 
      RECT 28.048 9.666 28.152 14.04 ; 
      RECT 27.616 9.666 27.72 14.04 ; 
      RECT 27.184 9.666 27.288 14.04 ; 
      RECT 26.752 9.666 26.856 14.04 ; 
      RECT 26.32 9.666 26.424 14.04 ; 
      RECT 25.888 9.666 25.992 14.04 ; 
      RECT 25.456 9.666 25.56 14.04 ; 
      RECT 25.024 9.666 25.128 14.04 ; 
      RECT 24.592 9.666 24.696 14.04 ; 
      RECT 24.16 9.666 24.264 14.04 ; 
      RECT 23.728 9.666 23.832 14.04 ; 
      RECT 23.296 9.666 23.4 14.04 ; 
      RECT 22.864 9.666 22.968 14.04 ; 
      RECT 22.432 9.666 22.536 14.04 ; 
      RECT 22 9.666 22.104 14.04 ; 
      RECT 21.568 9.666 21.672 14.04 ; 
      RECT 21.136 9.666 21.24 14.04 ; 
      RECT 20.704 9.666 20.808 14.04 ; 
      RECT 20.272 9.666 20.376 14.04 ; 
      RECT 19.84 9.666 19.944 14.04 ; 
      RECT 19.408 9.666 19.512 14.04 ; 
      RECT 18.976 9.666 19.08 14.04 ; 
      RECT 18.544 9.666 18.648 14.04 ; 
      RECT 18.112 9.666 18.216 14.04 ; 
      RECT 17.68 9.666 17.784 14.04 ; 
      RECT 17.248 9.666 17.352 14.04 ; 
      RECT 16.816 9.666 16.92 14.04 ; 
      RECT 16.384 9.666 16.488 14.04 ; 
      RECT 15.952 9.666 16.056 14.04 ; 
      RECT 15.52 9.666 15.624 14.04 ; 
      RECT 15.088 9.666 15.192 14.04 ; 
      RECT 14.656 9.666 14.76 14.04 ; 
      RECT 14.224 9.666 14.328 14.04 ; 
      RECT 13.792 9.666 13.896 14.04 ; 
      RECT 13.36 9.666 13.464 14.04 ; 
      RECT 12.928 9.666 13.032 14.04 ; 
      RECT 12.496 9.666 12.6 14.04 ; 
      RECT 12.064 9.666 12.168 14.04 ; 
      RECT 11.632 9.666 11.736 14.04 ; 
      RECT 11.2 9.666 11.304 14.04 ; 
      RECT 10.768 9.666 10.872 14.04 ; 
      RECT 10.336 9.666 10.44 14.04 ; 
      RECT 9.904 9.666 10.008 14.04 ; 
      RECT 9.472 9.666 9.576 14.04 ; 
      RECT 9.04 9.666 9.144 14.04 ; 
      RECT 8.608 9.666 8.712 14.04 ; 
      RECT 8.176 9.666 8.28 14.04 ; 
      RECT 7.744 9.666 7.848 14.04 ; 
      RECT 7.312 9.666 7.416 14.04 ; 
      RECT 6.88 9.666 6.984 14.04 ; 
      RECT 6.448 9.666 6.552 14.04 ; 
      RECT 6.016 9.666 6.12 14.04 ; 
      RECT 5.584 9.666 5.688 14.04 ; 
      RECT 5.152 9.666 5.256 14.04 ; 
      RECT 4.72 9.666 4.824 14.04 ; 
      RECT 4.288 9.666 4.392 14.04 ; 
      RECT 3.856 9.666 3.96 14.04 ; 
      RECT 3.424 9.666 3.528 14.04 ; 
      RECT 2.992 9.666 3.096 14.04 ; 
      RECT 2.56 9.666 2.664 14.04 ; 
      RECT 2.128 9.666 2.232 14.04 ; 
      RECT 1.696 9.666 1.8 14.04 ; 
      RECT 1.264 9.666 1.368 14.04 ; 
      RECT 0.832 9.666 0.936 14.04 ; 
      RECT 0.02 9.666 0.36 14.04 ; 
      RECT 62.212 13.986 62.724 18.36 ; 
      RECT 62.156 16.648 62.724 17.938 ; 
      RECT 61.276 15.556 61.812 18.36 ; 
      RECT 61.184 16.896 61.812 17.928 ; 
      RECT 61.276 13.986 61.668 18.36 ; 
      RECT 61.276 14.47 61.724 15.428 ; 
      RECT 61.276 13.986 61.812 14.342 ; 
      RECT 60.376 15.788 60.912 18.36 ; 
      RECT 60.376 13.986 60.768 18.36 ; 
      RECT 58.708 13.986 59.04 18.36 ; 
      RECT 58.708 14.34 59.096 18.082 ; 
      RECT 121.072 13.986 121.412 18.36 ; 
      RECT 120.496 13.986 120.6 18.36 ; 
      RECT 120.064 13.986 120.168 18.36 ; 
      RECT 119.632 13.986 119.736 18.36 ; 
      RECT 119.2 13.986 119.304 18.36 ; 
      RECT 118.768 13.986 118.872 18.36 ; 
      RECT 118.336 13.986 118.44 18.36 ; 
      RECT 117.904 13.986 118.008 18.36 ; 
      RECT 117.472 13.986 117.576 18.36 ; 
      RECT 117.04 13.986 117.144 18.36 ; 
      RECT 116.608 13.986 116.712 18.36 ; 
      RECT 116.176 13.986 116.28 18.36 ; 
      RECT 115.744 13.986 115.848 18.36 ; 
      RECT 115.312 13.986 115.416 18.36 ; 
      RECT 114.88 13.986 114.984 18.36 ; 
      RECT 114.448 13.986 114.552 18.36 ; 
      RECT 114.016 13.986 114.12 18.36 ; 
      RECT 113.584 13.986 113.688 18.36 ; 
      RECT 113.152 13.986 113.256 18.36 ; 
      RECT 112.72 13.986 112.824 18.36 ; 
      RECT 112.288 13.986 112.392 18.36 ; 
      RECT 111.856 13.986 111.96 18.36 ; 
      RECT 111.424 13.986 111.528 18.36 ; 
      RECT 110.992 13.986 111.096 18.36 ; 
      RECT 110.56 13.986 110.664 18.36 ; 
      RECT 110.128 13.986 110.232 18.36 ; 
      RECT 109.696 13.986 109.8 18.36 ; 
      RECT 109.264 13.986 109.368 18.36 ; 
      RECT 108.832 13.986 108.936 18.36 ; 
      RECT 108.4 13.986 108.504 18.36 ; 
      RECT 107.968 13.986 108.072 18.36 ; 
      RECT 107.536 13.986 107.64 18.36 ; 
      RECT 107.104 13.986 107.208 18.36 ; 
      RECT 106.672 13.986 106.776 18.36 ; 
      RECT 106.24 13.986 106.344 18.36 ; 
      RECT 105.808 13.986 105.912 18.36 ; 
      RECT 105.376 13.986 105.48 18.36 ; 
      RECT 104.944 13.986 105.048 18.36 ; 
      RECT 104.512 13.986 104.616 18.36 ; 
      RECT 104.08 13.986 104.184 18.36 ; 
      RECT 103.648 13.986 103.752 18.36 ; 
      RECT 103.216 13.986 103.32 18.36 ; 
      RECT 102.784 13.986 102.888 18.36 ; 
      RECT 102.352 13.986 102.456 18.36 ; 
      RECT 101.92 13.986 102.024 18.36 ; 
      RECT 101.488 13.986 101.592 18.36 ; 
      RECT 101.056 13.986 101.16 18.36 ; 
      RECT 100.624 13.986 100.728 18.36 ; 
      RECT 100.192 13.986 100.296 18.36 ; 
      RECT 99.76 13.986 99.864 18.36 ; 
      RECT 99.328 13.986 99.432 18.36 ; 
      RECT 98.896 13.986 99 18.36 ; 
      RECT 98.464 13.986 98.568 18.36 ; 
      RECT 98.032 13.986 98.136 18.36 ; 
      RECT 97.6 13.986 97.704 18.36 ; 
      RECT 97.168 13.986 97.272 18.36 ; 
      RECT 96.736 13.986 96.84 18.36 ; 
      RECT 96.304 13.986 96.408 18.36 ; 
      RECT 95.872 13.986 95.976 18.36 ; 
      RECT 95.44 13.986 95.544 18.36 ; 
      RECT 95.008 13.986 95.112 18.36 ; 
      RECT 94.576 13.986 94.68 18.36 ; 
      RECT 94.144 13.986 94.248 18.36 ; 
      RECT 93.712 13.986 93.816 18.36 ; 
      RECT 93.28 13.986 93.384 18.36 ; 
      RECT 92.848 13.986 92.952 18.36 ; 
      RECT 92.416 13.986 92.52 18.36 ; 
      RECT 91.984 13.986 92.088 18.36 ; 
      RECT 91.552 13.986 91.656 18.36 ; 
      RECT 91.12 13.986 91.224 18.36 ; 
      RECT 90.688 13.986 90.792 18.36 ; 
      RECT 90.256 13.986 90.36 18.36 ; 
      RECT 89.824 13.986 89.928 18.36 ; 
      RECT 89.392 13.986 89.496 18.36 ; 
      RECT 88.96 13.986 89.064 18.36 ; 
      RECT 88.528 13.986 88.632 18.36 ; 
      RECT 88.096 13.986 88.2 18.36 ; 
      RECT 87.664 13.986 87.768 18.36 ; 
      RECT 87.232 13.986 87.336 18.36 ; 
      RECT 86.8 13.986 86.904 18.36 ; 
      RECT 86.368 13.986 86.472 18.36 ; 
      RECT 85.936 13.986 86.04 18.36 ; 
      RECT 85.504 13.986 85.608 18.36 ; 
      RECT 85.072 13.986 85.176 18.36 ; 
      RECT 84.64 13.986 84.744 18.36 ; 
      RECT 84.208 13.986 84.312 18.36 ; 
      RECT 83.776 13.986 83.88 18.36 ; 
      RECT 83.344 13.986 83.448 18.36 ; 
      RECT 82.912 13.986 83.016 18.36 ; 
      RECT 82.48 13.986 82.584 18.36 ; 
      RECT 82.048 13.986 82.152 18.36 ; 
      RECT 81.616 13.986 81.72 18.36 ; 
      RECT 81.184 13.986 81.288 18.36 ; 
      RECT 80.752 13.986 80.856 18.36 ; 
      RECT 80.32 13.986 80.424 18.36 ; 
      RECT 79.888 13.986 79.992 18.36 ; 
      RECT 79.456 13.986 79.56 18.36 ; 
      RECT 79.024 13.986 79.128 18.36 ; 
      RECT 78.592 13.986 78.696 18.36 ; 
      RECT 78.16 13.986 78.264 18.36 ; 
      RECT 77.728 13.986 77.832 18.36 ; 
      RECT 77.296 13.986 77.4 18.36 ; 
      RECT 76.864 13.986 76.968 18.36 ; 
      RECT 76.432 13.986 76.536 18.36 ; 
      RECT 76 13.986 76.104 18.36 ; 
      RECT 75.568 13.986 75.672 18.36 ; 
      RECT 75.136 13.986 75.24 18.36 ; 
      RECT 74.704 13.986 74.808 18.36 ; 
      RECT 74.272 13.986 74.376 18.36 ; 
      RECT 73.84 13.986 73.944 18.36 ; 
      RECT 73.408 13.986 73.512 18.36 ; 
      RECT 72.976 13.986 73.08 18.36 ; 
      RECT 72.544 13.986 72.648 18.36 ; 
      RECT 72.112 13.986 72.216 18.36 ; 
      RECT 71.68 13.986 71.784 18.36 ; 
      RECT 71.248 13.986 71.352 18.36 ; 
      RECT 70.816 13.986 70.92 18.36 ; 
      RECT 70.384 13.986 70.488 18.36 ; 
      RECT 69.952 13.986 70.056 18.36 ; 
      RECT 69.52 13.986 69.624 18.36 ; 
      RECT 69.088 13.986 69.192 18.36 ; 
      RECT 68.656 13.986 68.76 18.36 ; 
      RECT 68.224 13.986 68.328 18.36 ; 
      RECT 67.792 13.986 67.896 18.36 ; 
      RECT 67.36 13.986 67.464 18.36 ; 
      RECT 66.928 13.986 67.032 18.36 ; 
      RECT 66.496 13.986 66.6 18.36 ; 
      RECT 66.064 13.986 66.168 18.36 ; 
      RECT 65.632 13.986 65.736 18.36 ; 
      RECT 65.2 13.986 65.304 18.36 ; 
      RECT 64.348 13.986 64.656 18.36 ; 
      RECT 56.776 13.986 57.084 18.36 ; 
      RECT 56.128 13.986 56.232 18.36 ; 
      RECT 55.696 13.986 55.8 18.36 ; 
      RECT 55.264 13.986 55.368 18.36 ; 
      RECT 54.832 13.986 54.936 18.36 ; 
      RECT 54.4 13.986 54.504 18.36 ; 
      RECT 53.968 13.986 54.072 18.36 ; 
      RECT 53.536 13.986 53.64 18.36 ; 
      RECT 53.104 13.986 53.208 18.36 ; 
      RECT 52.672 13.986 52.776 18.36 ; 
      RECT 52.24 13.986 52.344 18.36 ; 
      RECT 51.808 13.986 51.912 18.36 ; 
      RECT 51.376 13.986 51.48 18.36 ; 
      RECT 50.944 13.986 51.048 18.36 ; 
      RECT 50.512 13.986 50.616 18.36 ; 
      RECT 50.08 13.986 50.184 18.36 ; 
      RECT 49.648 13.986 49.752 18.36 ; 
      RECT 49.216 13.986 49.32 18.36 ; 
      RECT 48.784 13.986 48.888 18.36 ; 
      RECT 48.352 13.986 48.456 18.36 ; 
      RECT 47.92 13.986 48.024 18.36 ; 
      RECT 47.488 13.986 47.592 18.36 ; 
      RECT 47.056 13.986 47.16 18.36 ; 
      RECT 46.624 13.986 46.728 18.36 ; 
      RECT 46.192 13.986 46.296 18.36 ; 
      RECT 45.76 13.986 45.864 18.36 ; 
      RECT 45.328 13.986 45.432 18.36 ; 
      RECT 44.896 13.986 45 18.36 ; 
      RECT 44.464 13.986 44.568 18.36 ; 
      RECT 44.032 13.986 44.136 18.36 ; 
      RECT 43.6 13.986 43.704 18.36 ; 
      RECT 43.168 13.986 43.272 18.36 ; 
      RECT 42.736 13.986 42.84 18.36 ; 
      RECT 42.304 13.986 42.408 18.36 ; 
      RECT 41.872 13.986 41.976 18.36 ; 
      RECT 41.44 13.986 41.544 18.36 ; 
      RECT 41.008 13.986 41.112 18.36 ; 
      RECT 40.576 13.986 40.68 18.36 ; 
      RECT 40.144 13.986 40.248 18.36 ; 
      RECT 39.712 13.986 39.816 18.36 ; 
      RECT 39.28 13.986 39.384 18.36 ; 
      RECT 38.848 13.986 38.952 18.36 ; 
      RECT 38.416 13.986 38.52 18.36 ; 
      RECT 37.984 13.986 38.088 18.36 ; 
      RECT 37.552 13.986 37.656 18.36 ; 
      RECT 37.12 13.986 37.224 18.36 ; 
      RECT 36.688 13.986 36.792 18.36 ; 
      RECT 36.256 13.986 36.36 18.36 ; 
      RECT 35.824 13.986 35.928 18.36 ; 
      RECT 35.392 13.986 35.496 18.36 ; 
      RECT 34.96 13.986 35.064 18.36 ; 
      RECT 34.528 13.986 34.632 18.36 ; 
      RECT 34.096 13.986 34.2 18.36 ; 
      RECT 33.664 13.986 33.768 18.36 ; 
      RECT 33.232 13.986 33.336 18.36 ; 
      RECT 32.8 13.986 32.904 18.36 ; 
      RECT 32.368 13.986 32.472 18.36 ; 
      RECT 31.936 13.986 32.04 18.36 ; 
      RECT 31.504 13.986 31.608 18.36 ; 
      RECT 31.072 13.986 31.176 18.36 ; 
      RECT 30.64 13.986 30.744 18.36 ; 
      RECT 30.208 13.986 30.312 18.36 ; 
      RECT 29.776 13.986 29.88 18.36 ; 
      RECT 29.344 13.986 29.448 18.36 ; 
      RECT 28.912 13.986 29.016 18.36 ; 
      RECT 28.48 13.986 28.584 18.36 ; 
      RECT 28.048 13.986 28.152 18.36 ; 
      RECT 27.616 13.986 27.72 18.36 ; 
      RECT 27.184 13.986 27.288 18.36 ; 
      RECT 26.752 13.986 26.856 18.36 ; 
      RECT 26.32 13.986 26.424 18.36 ; 
      RECT 25.888 13.986 25.992 18.36 ; 
      RECT 25.456 13.986 25.56 18.36 ; 
      RECT 25.024 13.986 25.128 18.36 ; 
      RECT 24.592 13.986 24.696 18.36 ; 
      RECT 24.16 13.986 24.264 18.36 ; 
      RECT 23.728 13.986 23.832 18.36 ; 
      RECT 23.296 13.986 23.4 18.36 ; 
      RECT 22.864 13.986 22.968 18.36 ; 
      RECT 22.432 13.986 22.536 18.36 ; 
      RECT 22 13.986 22.104 18.36 ; 
      RECT 21.568 13.986 21.672 18.36 ; 
      RECT 21.136 13.986 21.24 18.36 ; 
      RECT 20.704 13.986 20.808 18.36 ; 
      RECT 20.272 13.986 20.376 18.36 ; 
      RECT 19.84 13.986 19.944 18.36 ; 
      RECT 19.408 13.986 19.512 18.36 ; 
      RECT 18.976 13.986 19.08 18.36 ; 
      RECT 18.544 13.986 18.648 18.36 ; 
      RECT 18.112 13.986 18.216 18.36 ; 
      RECT 17.68 13.986 17.784 18.36 ; 
      RECT 17.248 13.986 17.352 18.36 ; 
      RECT 16.816 13.986 16.92 18.36 ; 
      RECT 16.384 13.986 16.488 18.36 ; 
      RECT 15.952 13.986 16.056 18.36 ; 
      RECT 15.52 13.986 15.624 18.36 ; 
      RECT 15.088 13.986 15.192 18.36 ; 
      RECT 14.656 13.986 14.76 18.36 ; 
      RECT 14.224 13.986 14.328 18.36 ; 
      RECT 13.792 13.986 13.896 18.36 ; 
      RECT 13.36 13.986 13.464 18.36 ; 
      RECT 12.928 13.986 13.032 18.36 ; 
      RECT 12.496 13.986 12.6 18.36 ; 
      RECT 12.064 13.986 12.168 18.36 ; 
      RECT 11.632 13.986 11.736 18.36 ; 
      RECT 11.2 13.986 11.304 18.36 ; 
      RECT 10.768 13.986 10.872 18.36 ; 
      RECT 10.336 13.986 10.44 18.36 ; 
      RECT 9.904 13.986 10.008 18.36 ; 
      RECT 9.472 13.986 9.576 18.36 ; 
      RECT 9.04 13.986 9.144 18.36 ; 
      RECT 8.608 13.986 8.712 18.36 ; 
      RECT 8.176 13.986 8.28 18.36 ; 
      RECT 7.744 13.986 7.848 18.36 ; 
      RECT 7.312 13.986 7.416 18.36 ; 
      RECT 6.88 13.986 6.984 18.36 ; 
      RECT 6.448 13.986 6.552 18.36 ; 
      RECT 6.016 13.986 6.12 18.36 ; 
      RECT 5.584 13.986 5.688 18.36 ; 
      RECT 5.152 13.986 5.256 18.36 ; 
      RECT 4.72 13.986 4.824 18.36 ; 
      RECT 4.288 13.986 4.392 18.36 ; 
      RECT 3.856 13.986 3.96 18.36 ; 
      RECT 3.424 13.986 3.528 18.36 ; 
      RECT 2.992 13.986 3.096 18.36 ; 
      RECT 2.56 13.986 2.664 18.36 ; 
      RECT 2.128 13.986 2.232 18.36 ; 
      RECT 1.696 13.986 1.8 18.36 ; 
      RECT 1.264 13.986 1.368 18.36 ; 
      RECT 0.832 13.986 0.936 18.36 ; 
      RECT 0.02 13.986 0.36 18.36 ; 
      RECT 62.212 18.306 62.724 22.68 ; 
      RECT 62.156 20.968 62.724 22.258 ; 
      RECT 61.276 19.876 61.812 22.68 ; 
      RECT 61.184 21.216 61.812 22.248 ; 
      RECT 61.276 18.306 61.668 22.68 ; 
      RECT 61.276 18.79 61.724 19.748 ; 
      RECT 61.276 18.306 61.812 18.662 ; 
      RECT 60.376 20.108 60.912 22.68 ; 
      RECT 60.376 18.306 60.768 22.68 ; 
      RECT 58.708 18.306 59.04 22.68 ; 
      RECT 58.708 18.66 59.096 22.402 ; 
      RECT 121.072 18.306 121.412 22.68 ; 
      RECT 120.496 18.306 120.6 22.68 ; 
      RECT 120.064 18.306 120.168 22.68 ; 
      RECT 119.632 18.306 119.736 22.68 ; 
      RECT 119.2 18.306 119.304 22.68 ; 
      RECT 118.768 18.306 118.872 22.68 ; 
      RECT 118.336 18.306 118.44 22.68 ; 
      RECT 117.904 18.306 118.008 22.68 ; 
      RECT 117.472 18.306 117.576 22.68 ; 
      RECT 117.04 18.306 117.144 22.68 ; 
      RECT 116.608 18.306 116.712 22.68 ; 
      RECT 116.176 18.306 116.28 22.68 ; 
      RECT 115.744 18.306 115.848 22.68 ; 
      RECT 115.312 18.306 115.416 22.68 ; 
      RECT 114.88 18.306 114.984 22.68 ; 
      RECT 114.448 18.306 114.552 22.68 ; 
      RECT 114.016 18.306 114.12 22.68 ; 
      RECT 113.584 18.306 113.688 22.68 ; 
      RECT 113.152 18.306 113.256 22.68 ; 
      RECT 112.72 18.306 112.824 22.68 ; 
      RECT 112.288 18.306 112.392 22.68 ; 
      RECT 111.856 18.306 111.96 22.68 ; 
      RECT 111.424 18.306 111.528 22.68 ; 
      RECT 110.992 18.306 111.096 22.68 ; 
      RECT 110.56 18.306 110.664 22.68 ; 
      RECT 110.128 18.306 110.232 22.68 ; 
      RECT 109.696 18.306 109.8 22.68 ; 
      RECT 109.264 18.306 109.368 22.68 ; 
      RECT 108.832 18.306 108.936 22.68 ; 
      RECT 108.4 18.306 108.504 22.68 ; 
      RECT 107.968 18.306 108.072 22.68 ; 
      RECT 107.536 18.306 107.64 22.68 ; 
      RECT 107.104 18.306 107.208 22.68 ; 
      RECT 106.672 18.306 106.776 22.68 ; 
      RECT 106.24 18.306 106.344 22.68 ; 
      RECT 105.808 18.306 105.912 22.68 ; 
      RECT 105.376 18.306 105.48 22.68 ; 
      RECT 104.944 18.306 105.048 22.68 ; 
      RECT 104.512 18.306 104.616 22.68 ; 
      RECT 104.08 18.306 104.184 22.68 ; 
      RECT 103.648 18.306 103.752 22.68 ; 
      RECT 103.216 18.306 103.32 22.68 ; 
      RECT 102.784 18.306 102.888 22.68 ; 
      RECT 102.352 18.306 102.456 22.68 ; 
      RECT 101.92 18.306 102.024 22.68 ; 
      RECT 101.488 18.306 101.592 22.68 ; 
      RECT 101.056 18.306 101.16 22.68 ; 
      RECT 100.624 18.306 100.728 22.68 ; 
      RECT 100.192 18.306 100.296 22.68 ; 
      RECT 99.76 18.306 99.864 22.68 ; 
      RECT 99.328 18.306 99.432 22.68 ; 
      RECT 98.896 18.306 99 22.68 ; 
      RECT 98.464 18.306 98.568 22.68 ; 
      RECT 98.032 18.306 98.136 22.68 ; 
      RECT 97.6 18.306 97.704 22.68 ; 
      RECT 97.168 18.306 97.272 22.68 ; 
      RECT 96.736 18.306 96.84 22.68 ; 
      RECT 96.304 18.306 96.408 22.68 ; 
      RECT 95.872 18.306 95.976 22.68 ; 
      RECT 95.44 18.306 95.544 22.68 ; 
      RECT 95.008 18.306 95.112 22.68 ; 
      RECT 94.576 18.306 94.68 22.68 ; 
      RECT 94.144 18.306 94.248 22.68 ; 
      RECT 93.712 18.306 93.816 22.68 ; 
      RECT 93.28 18.306 93.384 22.68 ; 
      RECT 92.848 18.306 92.952 22.68 ; 
      RECT 92.416 18.306 92.52 22.68 ; 
      RECT 91.984 18.306 92.088 22.68 ; 
      RECT 91.552 18.306 91.656 22.68 ; 
      RECT 91.12 18.306 91.224 22.68 ; 
      RECT 90.688 18.306 90.792 22.68 ; 
      RECT 90.256 18.306 90.36 22.68 ; 
      RECT 89.824 18.306 89.928 22.68 ; 
      RECT 89.392 18.306 89.496 22.68 ; 
      RECT 88.96 18.306 89.064 22.68 ; 
      RECT 88.528 18.306 88.632 22.68 ; 
      RECT 88.096 18.306 88.2 22.68 ; 
      RECT 87.664 18.306 87.768 22.68 ; 
      RECT 87.232 18.306 87.336 22.68 ; 
      RECT 86.8 18.306 86.904 22.68 ; 
      RECT 86.368 18.306 86.472 22.68 ; 
      RECT 85.936 18.306 86.04 22.68 ; 
      RECT 85.504 18.306 85.608 22.68 ; 
      RECT 85.072 18.306 85.176 22.68 ; 
      RECT 84.64 18.306 84.744 22.68 ; 
      RECT 84.208 18.306 84.312 22.68 ; 
      RECT 83.776 18.306 83.88 22.68 ; 
      RECT 83.344 18.306 83.448 22.68 ; 
      RECT 82.912 18.306 83.016 22.68 ; 
      RECT 82.48 18.306 82.584 22.68 ; 
      RECT 82.048 18.306 82.152 22.68 ; 
      RECT 81.616 18.306 81.72 22.68 ; 
      RECT 81.184 18.306 81.288 22.68 ; 
      RECT 80.752 18.306 80.856 22.68 ; 
      RECT 80.32 18.306 80.424 22.68 ; 
      RECT 79.888 18.306 79.992 22.68 ; 
      RECT 79.456 18.306 79.56 22.68 ; 
      RECT 79.024 18.306 79.128 22.68 ; 
      RECT 78.592 18.306 78.696 22.68 ; 
      RECT 78.16 18.306 78.264 22.68 ; 
      RECT 77.728 18.306 77.832 22.68 ; 
      RECT 77.296 18.306 77.4 22.68 ; 
      RECT 76.864 18.306 76.968 22.68 ; 
      RECT 76.432 18.306 76.536 22.68 ; 
      RECT 76 18.306 76.104 22.68 ; 
      RECT 75.568 18.306 75.672 22.68 ; 
      RECT 75.136 18.306 75.24 22.68 ; 
      RECT 74.704 18.306 74.808 22.68 ; 
      RECT 74.272 18.306 74.376 22.68 ; 
      RECT 73.84 18.306 73.944 22.68 ; 
      RECT 73.408 18.306 73.512 22.68 ; 
      RECT 72.976 18.306 73.08 22.68 ; 
      RECT 72.544 18.306 72.648 22.68 ; 
      RECT 72.112 18.306 72.216 22.68 ; 
      RECT 71.68 18.306 71.784 22.68 ; 
      RECT 71.248 18.306 71.352 22.68 ; 
      RECT 70.816 18.306 70.92 22.68 ; 
      RECT 70.384 18.306 70.488 22.68 ; 
      RECT 69.952 18.306 70.056 22.68 ; 
      RECT 69.52 18.306 69.624 22.68 ; 
      RECT 69.088 18.306 69.192 22.68 ; 
      RECT 68.656 18.306 68.76 22.68 ; 
      RECT 68.224 18.306 68.328 22.68 ; 
      RECT 67.792 18.306 67.896 22.68 ; 
      RECT 67.36 18.306 67.464 22.68 ; 
      RECT 66.928 18.306 67.032 22.68 ; 
      RECT 66.496 18.306 66.6 22.68 ; 
      RECT 66.064 18.306 66.168 22.68 ; 
      RECT 65.632 18.306 65.736 22.68 ; 
      RECT 65.2 18.306 65.304 22.68 ; 
      RECT 64.348 18.306 64.656 22.68 ; 
      RECT 56.776 18.306 57.084 22.68 ; 
      RECT 56.128 18.306 56.232 22.68 ; 
      RECT 55.696 18.306 55.8 22.68 ; 
      RECT 55.264 18.306 55.368 22.68 ; 
      RECT 54.832 18.306 54.936 22.68 ; 
      RECT 54.4 18.306 54.504 22.68 ; 
      RECT 53.968 18.306 54.072 22.68 ; 
      RECT 53.536 18.306 53.64 22.68 ; 
      RECT 53.104 18.306 53.208 22.68 ; 
      RECT 52.672 18.306 52.776 22.68 ; 
      RECT 52.24 18.306 52.344 22.68 ; 
      RECT 51.808 18.306 51.912 22.68 ; 
      RECT 51.376 18.306 51.48 22.68 ; 
      RECT 50.944 18.306 51.048 22.68 ; 
      RECT 50.512 18.306 50.616 22.68 ; 
      RECT 50.08 18.306 50.184 22.68 ; 
      RECT 49.648 18.306 49.752 22.68 ; 
      RECT 49.216 18.306 49.32 22.68 ; 
      RECT 48.784 18.306 48.888 22.68 ; 
      RECT 48.352 18.306 48.456 22.68 ; 
      RECT 47.92 18.306 48.024 22.68 ; 
      RECT 47.488 18.306 47.592 22.68 ; 
      RECT 47.056 18.306 47.16 22.68 ; 
      RECT 46.624 18.306 46.728 22.68 ; 
      RECT 46.192 18.306 46.296 22.68 ; 
      RECT 45.76 18.306 45.864 22.68 ; 
      RECT 45.328 18.306 45.432 22.68 ; 
      RECT 44.896 18.306 45 22.68 ; 
      RECT 44.464 18.306 44.568 22.68 ; 
      RECT 44.032 18.306 44.136 22.68 ; 
      RECT 43.6 18.306 43.704 22.68 ; 
      RECT 43.168 18.306 43.272 22.68 ; 
      RECT 42.736 18.306 42.84 22.68 ; 
      RECT 42.304 18.306 42.408 22.68 ; 
      RECT 41.872 18.306 41.976 22.68 ; 
      RECT 41.44 18.306 41.544 22.68 ; 
      RECT 41.008 18.306 41.112 22.68 ; 
      RECT 40.576 18.306 40.68 22.68 ; 
      RECT 40.144 18.306 40.248 22.68 ; 
      RECT 39.712 18.306 39.816 22.68 ; 
      RECT 39.28 18.306 39.384 22.68 ; 
      RECT 38.848 18.306 38.952 22.68 ; 
      RECT 38.416 18.306 38.52 22.68 ; 
      RECT 37.984 18.306 38.088 22.68 ; 
      RECT 37.552 18.306 37.656 22.68 ; 
      RECT 37.12 18.306 37.224 22.68 ; 
      RECT 36.688 18.306 36.792 22.68 ; 
      RECT 36.256 18.306 36.36 22.68 ; 
      RECT 35.824 18.306 35.928 22.68 ; 
      RECT 35.392 18.306 35.496 22.68 ; 
      RECT 34.96 18.306 35.064 22.68 ; 
      RECT 34.528 18.306 34.632 22.68 ; 
      RECT 34.096 18.306 34.2 22.68 ; 
      RECT 33.664 18.306 33.768 22.68 ; 
      RECT 33.232 18.306 33.336 22.68 ; 
      RECT 32.8 18.306 32.904 22.68 ; 
      RECT 32.368 18.306 32.472 22.68 ; 
      RECT 31.936 18.306 32.04 22.68 ; 
      RECT 31.504 18.306 31.608 22.68 ; 
      RECT 31.072 18.306 31.176 22.68 ; 
      RECT 30.64 18.306 30.744 22.68 ; 
      RECT 30.208 18.306 30.312 22.68 ; 
      RECT 29.776 18.306 29.88 22.68 ; 
      RECT 29.344 18.306 29.448 22.68 ; 
      RECT 28.912 18.306 29.016 22.68 ; 
      RECT 28.48 18.306 28.584 22.68 ; 
      RECT 28.048 18.306 28.152 22.68 ; 
      RECT 27.616 18.306 27.72 22.68 ; 
      RECT 27.184 18.306 27.288 22.68 ; 
      RECT 26.752 18.306 26.856 22.68 ; 
      RECT 26.32 18.306 26.424 22.68 ; 
      RECT 25.888 18.306 25.992 22.68 ; 
      RECT 25.456 18.306 25.56 22.68 ; 
      RECT 25.024 18.306 25.128 22.68 ; 
      RECT 24.592 18.306 24.696 22.68 ; 
      RECT 24.16 18.306 24.264 22.68 ; 
      RECT 23.728 18.306 23.832 22.68 ; 
      RECT 23.296 18.306 23.4 22.68 ; 
      RECT 22.864 18.306 22.968 22.68 ; 
      RECT 22.432 18.306 22.536 22.68 ; 
      RECT 22 18.306 22.104 22.68 ; 
      RECT 21.568 18.306 21.672 22.68 ; 
      RECT 21.136 18.306 21.24 22.68 ; 
      RECT 20.704 18.306 20.808 22.68 ; 
      RECT 20.272 18.306 20.376 22.68 ; 
      RECT 19.84 18.306 19.944 22.68 ; 
      RECT 19.408 18.306 19.512 22.68 ; 
      RECT 18.976 18.306 19.08 22.68 ; 
      RECT 18.544 18.306 18.648 22.68 ; 
      RECT 18.112 18.306 18.216 22.68 ; 
      RECT 17.68 18.306 17.784 22.68 ; 
      RECT 17.248 18.306 17.352 22.68 ; 
      RECT 16.816 18.306 16.92 22.68 ; 
      RECT 16.384 18.306 16.488 22.68 ; 
      RECT 15.952 18.306 16.056 22.68 ; 
      RECT 15.52 18.306 15.624 22.68 ; 
      RECT 15.088 18.306 15.192 22.68 ; 
      RECT 14.656 18.306 14.76 22.68 ; 
      RECT 14.224 18.306 14.328 22.68 ; 
      RECT 13.792 18.306 13.896 22.68 ; 
      RECT 13.36 18.306 13.464 22.68 ; 
      RECT 12.928 18.306 13.032 22.68 ; 
      RECT 12.496 18.306 12.6 22.68 ; 
      RECT 12.064 18.306 12.168 22.68 ; 
      RECT 11.632 18.306 11.736 22.68 ; 
      RECT 11.2 18.306 11.304 22.68 ; 
      RECT 10.768 18.306 10.872 22.68 ; 
      RECT 10.336 18.306 10.44 22.68 ; 
      RECT 9.904 18.306 10.008 22.68 ; 
      RECT 9.472 18.306 9.576 22.68 ; 
      RECT 9.04 18.306 9.144 22.68 ; 
      RECT 8.608 18.306 8.712 22.68 ; 
      RECT 8.176 18.306 8.28 22.68 ; 
      RECT 7.744 18.306 7.848 22.68 ; 
      RECT 7.312 18.306 7.416 22.68 ; 
      RECT 6.88 18.306 6.984 22.68 ; 
      RECT 6.448 18.306 6.552 22.68 ; 
      RECT 6.016 18.306 6.12 22.68 ; 
      RECT 5.584 18.306 5.688 22.68 ; 
      RECT 5.152 18.306 5.256 22.68 ; 
      RECT 4.72 18.306 4.824 22.68 ; 
      RECT 4.288 18.306 4.392 22.68 ; 
      RECT 3.856 18.306 3.96 22.68 ; 
      RECT 3.424 18.306 3.528 22.68 ; 
      RECT 2.992 18.306 3.096 22.68 ; 
      RECT 2.56 18.306 2.664 22.68 ; 
      RECT 2.128 18.306 2.232 22.68 ; 
      RECT 1.696 18.306 1.8 22.68 ; 
      RECT 1.264 18.306 1.368 22.68 ; 
      RECT 0.832 18.306 0.936 22.68 ; 
      RECT 0.02 18.306 0.36 22.68 ; 
      RECT 62.212 22.626 62.724 27 ; 
      RECT 62.156 25.288 62.724 26.578 ; 
      RECT 61.276 24.196 61.812 27 ; 
      RECT 61.184 25.536 61.812 26.568 ; 
      RECT 61.276 22.626 61.668 27 ; 
      RECT 61.276 23.11 61.724 24.068 ; 
      RECT 61.276 22.626 61.812 22.982 ; 
      RECT 60.376 24.428 60.912 27 ; 
      RECT 60.376 22.626 60.768 27 ; 
      RECT 58.708 22.626 59.04 27 ; 
      RECT 58.708 22.98 59.096 26.722 ; 
      RECT 121.072 22.626 121.412 27 ; 
      RECT 120.496 22.626 120.6 27 ; 
      RECT 120.064 22.626 120.168 27 ; 
      RECT 119.632 22.626 119.736 27 ; 
      RECT 119.2 22.626 119.304 27 ; 
      RECT 118.768 22.626 118.872 27 ; 
      RECT 118.336 22.626 118.44 27 ; 
      RECT 117.904 22.626 118.008 27 ; 
      RECT 117.472 22.626 117.576 27 ; 
      RECT 117.04 22.626 117.144 27 ; 
      RECT 116.608 22.626 116.712 27 ; 
      RECT 116.176 22.626 116.28 27 ; 
      RECT 115.744 22.626 115.848 27 ; 
      RECT 115.312 22.626 115.416 27 ; 
      RECT 114.88 22.626 114.984 27 ; 
      RECT 114.448 22.626 114.552 27 ; 
      RECT 114.016 22.626 114.12 27 ; 
      RECT 113.584 22.626 113.688 27 ; 
      RECT 113.152 22.626 113.256 27 ; 
      RECT 112.72 22.626 112.824 27 ; 
      RECT 112.288 22.626 112.392 27 ; 
      RECT 111.856 22.626 111.96 27 ; 
      RECT 111.424 22.626 111.528 27 ; 
      RECT 110.992 22.626 111.096 27 ; 
      RECT 110.56 22.626 110.664 27 ; 
      RECT 110.128 22.626 110.232 27 ; 
      RECT 109.696 22.626 109.8 27 ; 
      RECT 109.264 22.626 109.368 27 ; 
      RECT 108.832 22.626 108.936 27 ; 
      RECT 108.4 22.626 108.504 27 ; 
      RECT 107.968 22.626 108.072 27 ; 
      RECT 107.536 22.626 107.64 27 ; 
      RECT 107.104 22.626 107.208 27 ; 
      RECT 106.672 22.626 106.776 27 ; 
      RECT 106.24 22.626 106.344 27 ; 
      RECT 105.808 22.626 105.912 27 ; 
      RECT 105.376 22.626 105.48 27 ; 
      RECT 104.944 22.626 105.048 27 ; 
      RECT 104.512 22.626 104.616 27 ; 
      RECT 104.08 22.626 104.184 27 ; 
      RECT 103.648 22.626 103.752 27 ; 
      RECT 103.216 22.626 103.32 27 ; 
      RECT 102.784 22.626 102.888 27 ; 
      RECT 102.352 22.626 102.456 27 ; 
      RECT 101.92 22.626 102.024 27 ; 
      RECT 101.488 22.626 101.592 27 ; 
      RECT 101.056 22.626 101.16 27 ; 
      RECT 100.624 22.626 100.728 27 ; 
      RECT 100.192 22.626 100.296 27 ; 
      RECT 99.76 22.626 99.864 27 ; 
      RECT 99.328 22.626 99.432 27 ; 
      RECT 98.896 22.626 99 27 ; 
      RECT 98.464 22.626 98.568 27 ; 
      RECT 98.032 22.626 98.136 27 ; 
      RECT 97.6 22.626 97.704 27 ; 
      RECT 97.168 22.626 97.272 27 ; 
      RECT 96.736 22.626 96.84 27 ; 
      RECT 96.304 22.626 96.408 27 ; 
      RECT 95.872 22.626 95.976 27 ; 
      RECT 95.44 22.626 95.544 27 ; 
      RECT 95.008 22.626 95.112 27 ; 
      RECT 94.576 22.626 94.68 27 ; 
      RECT 94.144 22.626 94.248 27 ; 
      RECT 93.712 22.626 93.816 27 ; 
      RECT 93.28 22.626 93.384 27 ; 
      RECT 92.848 22.626 92.952 27 ; 
      RECT 92.416 22.626 92.52 27 ; 
      RECT 91.984 22.626 92.088 27 ; 
      RECT 91.552 22.626 91.656 27 ; 
      RECT 91.12 22.626 91.224 27 ; 
      RECT 90.688 22.626 90.792 27 ; 
      RECT 90.256 22.626 90.36 27 ; 
      RECT 89.824 22.626 89.928 27 ; 
      RECT 89.392 22.626 89.496 27 ; 
      RECT 88.96 22.626 89.064 27 ; 
      RECT 88.528 22.626 88.632 27 ; 
      RECT 88.096 22.626 88.2 27 ; 
      RECT 87.664 22.626 87.768 27 ; 
      RECT 87.232 22.626 87.336 27 ; 
      RECT 86.8 22.626 86.904 27 ; 
      RECT 86.368 22.626 86.472 27 ; 
      RECT 85.936 22.626 86.04 27 ; 
      RECT 85.504 22.626 85.608 27 ; 
      RECT 85.072 22.626 85.176 27 ; 
      RECT 84.64 22.626 84.744 27 ; 
      RECT 84.208 22.626 84.312 27 ; 
      RECT 83.776 22.626 83.88 27 ; 
      RECT 83.344 22.626 83.448 27 ; 
      RECT 82.912 22.626 83.016 27 ; 
      RECT 82.48 22.626 82.584 27 ; 
      RECT 82.048 22.626 82.152 27 ; 
      RECT 81.616 22.626 81.72 27 ; 
      RECT 81.184 22.626 81.288 27 ; 
      RECT 80.752 22.626 80.856 27 ; 
      RECT 80.32 22.626 80.424 27 ; 
      RECT 79.888 22.626 79.992 27 ; 
      RECT 79.456 22.626 79.56 27 ; 
      RECT 79.024 22.626 79.128 27 ; 
      RECT 78.592 22.626 78.696 27 ; 
      RECT 78.16 22.626 78.264 27 ; 
      RECT 77.728 22.626 77.832 27 ; 
      RECT 77.296 22.626 77.4 27 ; 
      RECT 76.864 22.626 76.968 27 ; 
      RECT 76.432 22.626 76.536 27 ; 
      RECT 76 22.626 76.104 27 ; 
      RECT 75.568 22.626 75.672 27 ; 
      RECT 75.136 22.626 75.24 27 ; 
      RECT 74.704 22.626 74.808 27 ; 
      RECT 74.272 22.626 74.376 27 ; 
      RECT 73.84 22.626 73.944 27 ; 
      RECT 73.408 22.626 73.512 27 ; 
      RECT 72.976 22.626 73.08 27 ; 
      RECT 72.544 22.626 72.648 27 ; 
      RECT 72.112 22.626 72.216 27 ; 
      RECT 71.68 22.626 71.784 27 ; 
      RECT 71.248 22.626 71.352 27 ; 
      RECT 70.816 22.626 70.92 27 ; 
      RECT 70.384 22.626 70.488 27 ; 
      RECT 69.952 22.626 70.056 27 ; 
      RECT 69.52 22.626 69.624 27 ; 
      RECT 69.088 22.626 69.192 27 ; 
      RECT 68.656 22.626 68.76 27 ; 
      RECT 68.224 22.626 68.328 27 ; 
      RECT 67.792 22.626 67.896 27 ; 
      RECT 67.36 22.626 67.464 27 ; 
      RECT 66.928 22.626 67.032 27 ; 
      RECT 66.496 22.626 66.6 27 ; 
      RECT 66.064 22.626 66.168 27 ; 
      RECT 65.632 22.626 65.736 27 ; 
      RECT 65.2 22.626 65.304 27 ; 
      RECT 64.348 22.626 64.656 27 ; 
      RECT 56.776 22.626 57.084 27 ; 
      RECT 56.128 22.626 56.232 27 ; 
      RECT 55.696 22.626 55.8 27 ; 
      RECT 55.264 22.626 55.368 27 ; 
      RECT 54.832 22.626 54.936 27 ; 
      RECT 54.4 22.626 54.504 27 ; 
      RECT 53.968 22.626 54.072 27 ; 
      RECT 53.536 22.626 53.64 27 ; 
      RECT 53.104 22.626 53.208 27 ; 
      RECT 52.672 22.626 52.776 27 ; 
      RECT 52.24 22.626 52.344 27 ; 
      RECT 51.808 22.626 51.912 27 ; 
      RECT 51.376 22.626 51.48 27 ; 
      RECT 50.944 22.626 51.048 27 ; 
      RECT 50.512 22.626 50.616 27 ; 
      RECT 50.08 22.626 50.184 27 ; 
      RECT 49.648 22.626 49.752 27 ; 
      RECT 49.216 22.626 49.32 27 ; 
      RECT 48.784 22.626 48.888 27 ; 
      RECT 48.352 22.626 48.456 27 ; 
      RECT 47.92 22.626 48.024 27 ; 
      RECT 47.488 22.626 47.592 27 ; 
      RECT 47.056 22.626 47.16 27 ; 
      RECT 46.624 22.626 46.728 27 ; 
      RECT 46.192 22.626 46.296 27 ; 
      RECT 45.76 22.626 45.864 27 ; 
      RECT 45.328 22.626 45.432 27 ; 
      RECT 44.896 22.626 45 27 ; 
      RECT 44.464 22.626 44.568 27 ; 
      RECT 44.032 22.626 44.136 27 ; 
      RECT 43.6 22.626 43.704 27 ; 
      RECT 43.168 22.626 43.272 27 ; 
      RECT 42.736 22.626 42.84 27 ; 
      RECT 42.304 22.626 42.408 27 ; 
      RECT 41.872 22.626 41.976 27 ; 
      RECT 41.44 22.626 41.544 27 ; 
      RECT 41.008 22.626 41.112 27 ; 
      RECT 40.576 22.626 40.68 27 ; 
      RECT 40.144 22.626 40.248 27 ; 
      RECT 39.712 22.626 39.816 27 ; 
      RECT 39.28 22.626 39.384 27 ; 
      RECT 38.848 22.626 38.952 27 ; 
      RECT 38.416 22.626 38.52 27 ; 
      RECT 37.984 22.626 38.088 27 ; 
      RECT 37.552 22.626 37.656 27 ; 
      RECT 37.12 22.626 37.224 27 ; 
      RECT 36.688 22.626 36.792 27 ; 
      RECT 36.256 22.626 36.36 27 ; 
      RECT 35.824 22.626 35.928 27 ; 
      RECT 35.392 22.626 35.496 27 ; 
      RECT 34.96 22.626 35.064 27 ; 
      RECT 34.528 22.626 34.632 27 ; 
      RECT 34.096 22.626 34.2 27 ; 
      RECT 33.664 22.626 33.768 27 ; 
      RECT 33.232 22.626 33.336 27 ; 
      RECT 32.8 22.626 32.904 27 ; 
      RECT 32.368 22.626 32.472 27 ; 
      RECT 31.936 22.626 32.04 27 ; 
      RECT 31.504 22.626 31.608 27 ; 
      RECT 31.072 22.626 31.176 27 ; 
      RECT 30.64 22.626 30.744 27 ; 
      RECT 30.208 22.626 30.312 27 ; 
      RECT 29.776 22.626 29.88 27 ; 
      RECT 29.344 22.626 29.448 27 ; 
      RECT 28.912 22.626 29.016 27 ; 
      RECT 28.48 22.626 28.584 27 ; 
      RECT 28.048 22.626 28.152 27 ; 
      RECT 27.616 22.626 27.72 27 ; 
      RECT 27.184 22.626 27.288 27 ; 
      RECT 26.752 22.626 26.856 27 ; 
      RECT 26.32 22.626 26.424 27 ; 
      RECT 25.888 22.626 25.992 27 ; 
      RECT 25.456 22.626 25.56 27 ; 
      RECT 25.024 22.626 25.128 27 ; 
      RECT 24.592 22.626 24.696 27 ; 
      RECT 24.16 22.626 24.264 27 ; 
      RECT 23.728 22.626 23.832 27 ; 
      RECT 23.296 22.626 23.4 27 ; 
      RECT 22.864 22.626 22.968 27 ; 
      RECT 22.432 22.626 22.536 27 ; 
      RECT 22 22.626 22.104 27 ; 
      RECT 21.568 22.626 21.672 27 ; 
      RECT 21.136 22.626 21.24 27 ; 
      RECT 20.704 22.626 20.808 27 ; 
      RECT 20.272 22.626 20.376 27 ; 
      RECT 19.84 22.626 19.944 27 ; 
      RECT 19.408 22.626 19.512 27 ; 
      RECT 18.976 22.626 19.08 27 ; 
      RECT 18.544 22.626 18.648 27 ; 
      RECT 18.112 22.626 18.216 27 ; 
      RECT 17.68 22.626 17.784 27 ; 
      RECT 17.248 22.626 17.352 27 ; 
      RECT 16.816 22.626 16.92 27 ; 
      RECT 16.384 22.626 16.488 27 ; 
      RECT 15.952 22.626 16.056 27 ; 
      RECT 15.52 22.626 15.624 27 ; 
      RECT 15.088 22.626 15.192 27 ; 
      RECT 14.656 22.626 14.76 27 ; 
      RECT 14.224 22.626 14.328 27 ; 
      RECT 13.792 22.626 13.896 27 ; 
      RECT 13.36 22.626 13.464 27 ; 
      RECT 12.928 22.626 13.032 27 ; 
      RECT 12.496 22.626 12.6 27 ; 
      RECT 12.064 22.626 12.168 27 ; 
      RECT 11.632 22.626 11.736 27 ; 
      RECT 11.2 22.626 11.304 27 ; 
      RECT 10.768 22.626 10.872 27 ; 
      RECT 10.336 22.626 10.44 27 ; 
      RECT 9.904 22.626 10.008 27 ; 
      RECT 9.472 22.626 9.576 27 ; 
      RECT 9.04 22.626 9.144 27 ; 
      RECT 8.608 22.626 8.712 27 ; 
      RECT 8.176 22.626 8.28 27 ; 
      RECT 7.744 22.626 7.848 27 ; 
      RECT 7.312 22.626 7.416 27 ; 
      RECT 6.88 22.626 6.984 27 ; 
      RECT 6.448 22.626 6.552 27 ; 
      RECT 6.016 22.626 6.12 27 ; 
      RECT 5.584 22.626 5.688 27 ; 
      RECT 5.152 22.626 5.256 27 ; 
      RECT 4.72 22.626 4.824 27 ; 
      RECT 4.288 22.626 4.392 27 ; 
      RECT 3.856 22.626 3.96 27 ; 
      RECT 3.424 22.626 3.528 27 ; 
      RECT 2.992 22.626 3.096 27 ; 
      RECT 2.56 22.626 2.664 27 ; 
      RECT 2.128 22.626 2.232 27 ; 
      RECT 1.696 22.626 1.8 27 ; 
      RECT 1.264 22.626 1.368 27 ; 
      RECT 0.832 22.626 0.936 27 ; 
      RECT 0.02 22.626 0.36 27 ; 
      RECT 62.212 26.946 62.724 31.32 ; 
      RECT 62.156 29.608 62.724 30.898 ; 
      RECT 61.276 28.516 61.812 31.32 ; 
      RECT 61.184 29.856 61.812 30.888 ; 
      RECT 61.276 26.946 61.668 31.32 ; 
      RECT 61.276 27.43 61.724 28.388 ; 
      RECT 61.276 26.946 61.812 27.302 ; 
      RECT 60.376 28.748 60.912 31.32 ; 
      RECT 60.376 26.946 60.768 31.32 ; 
      RECT 58.708 26.946 59.04 31.32 ; 
      RECT 58.708 27.3 59.096 31.042 ; 
      RECT 121.072 26.946 121.412 31.32 ; 
      RECT 120.496 26.946 120.6 31.32 ; 
      RECT 120.064 26.946 120.168 31.32 ; 
      RECT 119.632 26.946 119.736 31.32 ; 
      RECT 119.2 26.946 119.304 31.32 ; 
      RECT 118.768 26.946 118.872 31.32 ; 
      RECT 118.336 26.946 118.44 31.32 ; 
      RECT 117.904 26.946 118.008 31.32 ; 
      RECT 117.472 26.946 117.576 31.32 ; 
      RECT 117.04 26.946 117.144 31.32 ; 
      RECT 116.608 26.946 116.712 31.32 ; 
      RECT 116.176 26.946 116.28 31.32 ; 
      RECT 115.744 26.946 115.848 31.32 ; 
      RECT 115.312 26.946 115.416 31.32 ; 
      RECT 114.88 26.946 114.984 31.32 ; 
      RECT 114.448 26.946 114.552 31.32 ; 
      RECT 114.016 26.946 114.12 31.32 ; 
      RECT 113.584 26.946 113.688 31.32 ; 
      RECT 113.152 26.946 113.256 31.32 ; 
      RECT 112.72 26.946 112.824 31.32 ; 
      RECT 112.288 26.946 112.392 31.32 ; 
      RECT 111.856 26.946 111.96 31.32 ; 
      RECT 111.424 26.946 111.528 31.32 ; 
      RECT 110.992 26.946 111.096 31.32 ; 
      RECT 110.56 26.946 110.664 31.32 ; 
      RECT 110.128 26.946 110.232 31.32 ; 
      RECT 109.696 26.946 109.8 31.32 ; 
      RECT 109.264 26.946 109.368 31.32 ; 
      RECT 108.832 26.946 108.936 31.32 ; 
      RECT 108.4 26.946 108.504 31.32 ; 
      RECT 107.968 26.946 108.072 31.32 ; 
      RECT 107.536 26.946 107.64 31.32 ; 
      RECT 107.104 26.946 107.208 31.32 ; 
      RECT 106.672 26.946 106.776 31.32 ; 
      RECT 106.24 26.946 106.344 31.32 ; 
      RECT 105.808 26.946 105.912 31.32 ; 
      RECT 105.376 26.946 105.48 31.32 ; 
      RECT 104.944 26.946 105.048 31.32 ; 
      RECT 104.512 26.946 104.616 31.32 ; 
      RECT 104.08 26.946 104.184 31.32 ; 
      RECT 103.648 26.946 103.752 31.32 ; 
      RECT 103.216 26.946 103.32 31.32 ; 
      RECT 102.784 26.946 102.888 31.32 ; 
      RECT 102.352 26.946 102.456 31.32 ; 
      RECT 101.92 26.946 102.024 31.32 ; 
      RECT 101.488 26.946 101.592 31.32 ; 
      RECT 101.056 26.946 101.16 31.32 ; 
      RECT 100.624 26.946 100.728 31.32 ; 
      RECT 100.192 26.946 100.296 31.32 ; 
      RECT 99.76 26.946 99.864 31.32 ; 
      RECT 99.328 26.946 99.432 31.32 ; 
      RECT 98.896 26.946 99 31.32 ; 
      RECT 98.464 26.946 98.568 31.32 ; 
      RECT 98.032 26.946 98.136 31.32 ; 
      RECT 97.6 26.946 97.704 31.32 ; 
      RECT 97.168 26.946 97.272 31.32 ; 
      RECT 96.736 26.946 96.84 31.32 ; 
      RECT 96.304 26.946 96.408 31.32 ; 
      RECT 95.872 26.946 95.976 31.32 ; 
      RECT 95.44 26.946 95.544 31.32 ; 
      RECT 95.008 26.946 95.112 31.32 ; 
      RECT 94.576 26.946 94.68 31.32 ; 
      RECT 94.144 26.946 94.248 31.32 ; 
      RECT 93.712 26.946 93.816 31.32 ; 
      RECT 93.28 26.946 93.384 31.32 ; 
      RECT 92.848 26.946 92.952 31.32 ; 
      RECT 92.416 26.946 92.52 31.32 ; 
      RECT 91.984 26.946 92.088 31.32 ; 
      RECT 91.552 26.946 91.656 31.32 ; 
      RECT 91.12 26.946 91.224 31.32 ; 
      RECT 90.688 26.946 90.792 31.32 ; 
      RECT 90.256 26.946 90.36 31.32 ; 
      RECT 89.824 26.946 89.928 31.32 ; 
      RECT 89.392 26.946 89.496 31.32 ; 
      RECT 88.96 26.946 89.064 31.32 ; 
      RECT 88.528 26.946 88.632 31.32 ; 
      RECT 88.096 26.946 88.2 31.32 ; 
      RECT 87.664 26.946 87.768 31.32 ; 
      RECT 87.232 26.946 87.336 31.32 ; 
      RECT 86.8 26.946 86.904 31.32 ; 
      RECT 86.368 26.946 86.472 31.32 ; 
      RECT 85.936 26.946 86.04 31.32 ; 
      RECT 85.504 26.946 85.608 31.32 ; 
      RECT 85.072 26.946 85.176 31.32 ; 
      RECT 84.64 26.946 84.744 31.32 ; 
      RECT 84.208 26.946 84.312 31.32 ; 
      RECT 83.776 26.946 83.88 31.32 ; 
      RECT 83.344 26.946 83.448 31.32 ; 
      RECT 82.912 26.946 83.016 31.32 ; 
      RECT 82.48 26.946 82.584 31.32 ; 
      RECT 82.048 26.946 82.152 31.32 ; 
      RECT 81.616 26.946 81.72 31.32 ; 
      RECT 81.184 26.946 81.288 31.32 ; 
      RECT 80.752 26.946 80.856 31.32 ; 
      RECT 80.32 26.946 80.424 31.32 ; 
      RECT 79.888 26.946 79.992 31.32 ; 
      RECT 79.456 26.946 79.56 31.32 ; 
      RECT 79.024 26.946 79.128 31.32 ; 
      RECT 78.592 26.946 78.696 31.32 ; 
      RECT 78.16 26.946 78.264 31.32 ; 
      RECT 77.728 26.946 77.832 31.32 ; 
      RECT 77.296 26.946 77.4 31.32 ; 
      RECT 76.864 26.946 76.968 31.32 ; 
      RECT 76.432 26.946 76.536 31.32 ; 
      RECT 76 26.946 76.104 31.32 ; 
      RECT 75.568 26.946 75.672 31.32 ; 
      RECT 75.136 26.946 75.24 31.32 ; 
      RECT 74.704 26.946 74.808 31.32 ; 
      RECT 74.272 26.946 74.376 31.32 ; 
      RECT 73.84 26.946 73.944 31.32 ; 
      RECT 73.408 26.946 73.512 31.32 ; 
      RECT 72.976 26.946 73.08 31.32 ; 
      RECT 72.544 26.946 72.648 31.32 ; 
      RECT 72.112 26.946 72.216 31.32 ; 
      RECT 71.68 26.946 71.784 31.32 ; 
      RECT 71.248 26.946 71.352 31.32 ; 
      RECT 70.816 26.946 70.92 31.32 ; 
      RECT 70.384 26.946 70.488 31.32 ; 
      RECT 69.952 26.946 70.056 31.32 ; 
      RECT 69.52 26.946 69.624 31.32 ; 
      RECT 69.088 26.946 69.192 31.32 ; 
      RECT 68.656 26.946 68.76 31.32 ; 
      RECT 68.224 26.946 68.328 31.32 ; 
      RECT 67.792 26.946 67.896 31.32 ; 
      RECT 67.36 26.946 67.464 31.32 ; 
      RECT 66.928 26.946 67.032 31.32 ; 
      RECT 66.496 26.946 66.6 31.32 ; 
      RECT 66.064 26.946 66.168 31.32 ; 
      RECT 65.632 26.946 65.736 31.32 ; 
      RECT 65.2 26.946 65.304 31.32 ; 
      RECT 64.348 26.946 64.656 31.32 ; 
      RECT 56.776 26.946 57.084 31.32 ; 
      RECT 56.128 26.946 56.232 31.32 ; 
      RECT 55.696 26.946 55.8 31.32 ; 
      RECT 55.264 26.946 55.368 31.32 ; 
      RECT 54.832 26.946 54.936 31.32 ; 
      RECT 54.4 26.946 54.504 31.32 ; 
      RECT 53.968 26.946 54.072 31.32 ; 
      RECT 53.536 26.946 53.64 31.32 ; 
      RECT 53.104 26.946 53.208 31.32 ; 
      RECT 52.672 26.946 52.776 31.32 ; 
      RECT 52.24 26.946 52.344 31.32 ; 
      RECT 51.808 26.946 51.912 31.32 ; 
      RECT 51.376 26.946 51.48 31.32 ; 
      RECT 50.944 26.946 51.048 31.32 ; 
      RECT 50.512 26.946 50.616 31.32 ; 
      RECT 50.08 26.946 50.184 31.32 ; 
      RECT 49.648 26.946 49.752 31.32 ; 
      RECT 49.216 26.946 49.32 31.32 ; 
      RECT 48.784 26.946 48.888 31.32 ; 
      RECT 48.352 26.946 48.456 31.32 ; 
      RECT 47.92 26.946 48.024 31.32 ; 
      RECT 47.488 26.946 47.592 31.32 ; 
      RECT 47.056 26.946 47.16 31.32 ; 
      RECT 46.624 26.946 46.728 31.32 ; 
      RECT 46.192 26.946 46.296 31.32 ; 
      RECT 45.76 26.946 45.864 31.32 ; 
      RECT 45.328 26.946 45.432 31.32 ; 
      RECT 44.896 26.946 45 31.32 ; 
      RECT 44.464 26.946 44.568 31.32 ; 
      RECT 44.032 26.946 44.136 31.32 ; 
      RECT 43.6 26.946 43.704 31.32 ; 
      RECT 43.168 26.946 43.272 31.32 ; 
      RECT 42.736 26.946 42.84 31.32 ; 
      RECT 42.304 26.946 42.408 31.32 ; 
      RECT 41.872 26.946 41.976 31.32 ; 
      RECT 41.44 26.946 41.544 31.32 ; 
      RECT 41.008 26.946 41.112 31.32 ; 
      RECT 40.576 26.946 40.68 31.32 ; 
      RECT 40.144 26.946 40.248 31.32 ; 
      RECT 39.712 26.946 39.816 31.32 ; 
      RECT 39.28 26.946 39.384 31.32 ; 
      RECT 38.848 26.946 38.952 31.32 ; 
      RECT 38.416 26.946 38.52 31.32 ; 
      RECT 37.984 26.946 38.088 31.32 ; 
      RECT 37.552 26.946 37.656 31.32 ; 
      RECT 37.12 26.946 37.224 31.32 ; 
      RECT 36.688 26.946 36.792 31.32 ; 
      RECT 36.256 26.946 36.36 31.32 ; 
      RECT 35.824 26.946 35.928 31.32 ; 
      RECT 35.392 26.946 35.496 31.32 ; 
      RECT 34.96 26.946 35.064 31.32 ; 
      RECT 34.528 26.946 34.632 31.32 ; 
      RECT 34.096 26.946 34.2 31.32 ; 
      RECT 33.664 26.946 33.768 31.32 ; 
      RECT 33.232 26.946 33.336 31.32 ; 
      RECT 32.8 26.946 32.904 31.32 ; 
      RECT 32.368 26.946 32.472 31.32 ; 
      RECT 31.936 26.946 32.04 31.32 ; 
      RECT 31.504 26.946 31.608 31.32 ; 
      RECT 31.072 26.946 31.176 31.32 ; 
      RECT 30.64 26.946 30.744 31.32 ; 
      RECT 30.208 26.946 30.312 31.32 ; 
      RECT 29.776 26.946 29.88 31.32 ; 
      RECT 29.344 26.946 29.448 31.32 ; 
      RECT 28.912 26.946 29.016 31.32 ; 
      RECT 28.48 26.946 28.584 31.32 ; 
      RECT 28.048 26.946 28.152 31.32 ; 
      RECT 27.616 26.946 27.72 31.32 ; 
      RECT 27.184 26.946 27.288 31.32 ; 
      RECT 26.752 26.946 26.856 31.32 ; 
      RECT 26.32 26.946 26.424 31.32 ; 
      RECT 25.888 26.946 25.992 31.32 ; 
      RECT 25.456 26.946 25.56 31.32 ; 
      RECT 25.024 26.946 25.128 31.32 ; 
      RECT 24.592 26.946 24.696 31.32 ; 
      RECT 24.16 26.946 24.264 31.32 ; 
      RECT 23.728 26.946 23.832 31.32 ; 
      RECT 23.296 26.946 23.4 31.32 ; 
      RECT 22.864 26.946 22.968 31.32 ; 
      RECT 22.432 26.946 22.536 31.32 ; 
      RECT 22 26.946 22.104 31.32 ; 
      RECT 21.568 26.946 21.672 31.32 ; 
      RECT 21.136 26.946 21.24 31.32 ; 
      RECT 20.704 26.946 20.808 31.32 ; 
      RECT 20.272 26.946 20.376 31.32 ; 
      RECT 19.84 26.946 19.944 31.32 ; 
      RECT 19.408 26.946 19.512 31.32 ; 
      RECT 18.976 26.946 19.08 31.32 ; 
      RECT 18.544 26.946 18.648 31.32 ; 
      RECT 18.112 26.946 18.216 31.32 ; 
      RECT 17.68 26.946 17.784 31.32 ; 
      RECT 17.248 26.946 17.352 31.32 ; 
      RECT 16.816 26.946 16.92 31.32 ; 
      RECT 16.384 26.946 16.488 31.32 ; 
      RECT 15.952 26.946 16.056 31.32 ; 
      RECT 15.52 26.946 15.624 31.32 ; 
      RECT 15.088 26.946 15.192 31.32 ; 
      RECT 14.656 26.946 14.76 31.32 ; 
      RECT 14.224 26.946 14.328 31.32 ; 
      RECT 13.792 26.946 13.896 31.32 ; 
      RECT 13.36 26.946 13.464 31.32 ; 
      RECT 12.928 26.946 13.032 31.32 ; 
      RECT 12.496 26.946 12.6 31.32 ; 
      RECT 12.064 26.946 12.168 31.32 ; 
      RECT 11.632 26.946 11.736 31.32 ; 
      RECT 11.2 26.946 11.304 31.32 ; 
      RECT 10.768 26.946 10.872 31.32 ; 
      RECT 10.336 26.946 10.44 31.32 ; 
      RECT 9.904 26.946 10.008 31.32 ; 
      RECT 9.472 26.946 9.576 31.32 ; 
      RECT 9.04 26.946 9.144 31.32 ; 
      RECT 8.608 26.946 8.712 31.32 ; 
      RECT 8.176 26.946 8.28 31.32 ; 
      RECT 7.744 26.946 7.848 31.32 ; 
      RECT 7.312 26.946 7.416 31.32 ; 
      RECT 6.88 26.946 6.984 31.32 ; 
      RECT 6.448 26.946 6.552 31.32 ; 
      RECT 6.016 26.946 6.12 31.32 ; 
      RECT 5.584 26.946 5.688 31.32 ; 
      RECT 5.152 26.946 5.256 31.32 ; 
      RECT 4.72 26.946 4.824 31.32 ; 
      RECT 4.288 26.946 4.392 31.32 ; 
      RECT 3.856 26.946 3.96 31.32 ; 
      RECT 3.424 26.946 3.528 31.32 ; 
      RECT 2.992 26.946 3.096 31.32 ; 
      RECT 2.56 26.946 2.664 31.32 ; 
      RECT 2.128 26.946 2.232 31.32 ; 
      RECT 1.696 26.946 1.8 31.32 ; 
      RECT 1.264 26.946 1.368 31.32 ; 
      RECT 0.832 26.946 0.936 31.32 ; 
      RECT 0.02 26.946 0.36 31.32 ; 
      RECT 62.212 31.266 62.724 35.64 ; 
      RECT 62.156 33.928 62.724 35.218 ; 
      RECT 61.276 32.836 61.812 35.64 ; 
      RECT 61.184 34.176 61.812 35.208 ; 
      RECT 61.276 31.266 61.668 35.64 ; 
      RECT 61.276 31.75 61.724 32.708 ; 
      RECT 61.276 31.266 61.812 31.622 ; 
      RECT 60.376 33.068 60.912 35.64 ; 
      RECT 60.376 31.266 60.768 35.64 ; 
      RECT 58.708 31.266 59.04 35.64 ; 
      RECT 58.708 31.62 59.096 35.362 ; 
      RECT 121.072 31.266 121.412 35.64 ; 
      RECT 120.496 31.266 120.6 35.64 ; 
      RECT 120.064 31.266 120.168 35.64 ; 
      RECT 119.632 31.266 119.736 35.64 ; 
      RECT 119.2 31.266 119.304 35.64 ; 
      RECT 118.768 31.266 118.872 35.64 ; 
      RECT 118.336 31.266 118.44 35.64 ; 
      RECT 117.904 31.266 118.008 35.64 ; 
      RECT 117.472 31.266 117.576 35.64 ; 
      RECT 117.04 31.266 117.144 35.64 ; 
      RECT 116.608 31.266 116.712 35.64 ; 
      RECT 116.176 31.266 116.28 35.64 ; 
      RECT 115.744 31.266 115.848 35.64 ; 
      RECT 115.312 31.266 115.416 35.64 ; 
      RECT 114.88 31.266 114.984 35.64 ; 
      RECT 114.448 31.266 114.552 35.64 ; 
      RECT 114.016 31.266 114.12 35.64 ; 
      RECT 113.584 31.266 113.688 35.64 ; 
      RECT 113.152 31.266 113.256 35.64 ; 
      RECT 112.72 31.266 112.824 35.64 ; 
      RECT 112.288 31.266 112.392 35.64 ; 
      RECT 111.856 31.266 111.96 35.64 ; 
      RECT 111.424 31.266 111.528 35.64 ; 
      RECT 110.992 31.266 111.096 35.64 ; 
      RECT 110.56 31.266 110.664 35.64 ; 
      RECT 110.128 31.266 110.232 35.64 ; 
      RECT 109.696 31.266 109.8 35.64 ; 
      RECT 109.264 31.266 109.368 35.64 ; 
      RECT 108.832 31.266 108.936 35.64 ; 
      RECT 108.4 31.266 108.504 35.64 ; 
      RECT 107.968 31.266 108.072 35.64 ; 
      RECT 107.536 31.266 107.64 35.64 ; 
      RECT 107.104 31.266 107.208 35.64 ; 
      RECT 106.672 31.266 106.776 35.64 ; 
      RECT 106.24 31.266 106.344 35.64 ; 
      RECT 105.808 31.266 105.912 35.64 ; 
      RECT 105.376 31.266 105.48 35.64 ; 
      RECT 104.944 31.266 105.048 35.64 ; 
      RECT 104.512 31.266 104.616 35.64 ; 
      RECT 104.08 31.266 104.184 35.64 ; 
      RECT 103.648 31.266 103.752 35.64 ; 
      RECT 103.216 31.266 103.32 35.64 ; 
      RECT 102.784 31.266 102.888 35.64 ; 
      RECT 102.352 31.266 102.456 35.64 ; 
      RECT 101.92 31.266 102.024 35.64 ; 
      RECT 101.488 31.266 101.592 35.64 ; 
      RECT 101.056 31.266 101.16 35.64 ; 
      RECT 100.624 31.266 100.728 35.64 ; 
      RECT 100.192 31.266 100.296 35.64 ; 
      RECT 99.76 31.266 99.864 35.64 ; 
      RECT 99.328 31.266 99.432 35.64 ; 
      RECT 98.896 31.266 99 35.64 ; 
      RECT 98.464 31.266 98.568 35.64 ; 
      RECT 98.032 31.266 98.136 35.64 ; 
      RECT 97.6 31.266 97.704 35.64 ; 
      RECT 97.168 31.266 97.272 35.64 ; 
      RECT 96.736 31.266 96.84 35.64 ; 
      RECT 96.304 31.266 96.408 35.64 ; 
      RECT 95.872 31.266 95.976 35.64 ; 
      RECT 95.44 31.266 95.544 35.64 ; 
      RECT 95.008 31.266 95.112 35.64 ; 
      RECT 94.576 31.266 94.68 35.64 ; 
      RECT 94.144 31.266 94.248 35.64 ; 
      RECT 93.712 31.266 93.816 35.64 ; 
      RECT 93.28 31.266 93.384 35.64 ; 
      RECT 92.848 31.266 92.952 35.64 ; 
      RECT 92.416 31.266 92.52 35.64 ; 
      RECT 91.984 31.266 92.088 35.64 ; 
      RECT 91.552 31.266 91.656 35.64 ; 
      RECT 91.12 31.266 91.224 35.64 ; 
      RECT 90.688 31.266 90.792 35.64 ; 
      RECT 90.256 31.266 90.36 35.64 ; 
      RECT 89.824 31.266 89.928 35.64 ; 
      RECT 89.392 31.266 89.496 35.64 ; 
      RECT 88.96 31.266 89.064 35.64 ; 
      RECT 88.528 31.266 88.632 35.64 ; 
      RECT 88.096 31.266 88.2 35.64 ; 
      RECT 87.664 31.266 87.768 35.64 ; 
      RECT 87.232 31.266 87.336 35.64 ; 
      RECT 86.8 31.266 86.904 35.64 ; 
      RECT 86.368 31.266 86.472 35.64 ; 
      RECT 85.936 31.266 86.04 35.64 ; 
      RECT 85.504 31.266 85.608 35.64 ; 
      RECT 85.072 31.266 85.176 35.64 ; 
      RECT 84.64 31.266 84.744 35.64 ; 
      RECT 84.208 31.266 84.312 35.64 ; 
      RECT 83.776 31.266 83.88 35.64 ; 
      RECT 83.344 31.266 83.448 35.64 ; 
      RECT 82.912 31.266 83.016 35.64 ; 
      RECT 82.48 31.266 82.584 35.64 ; 
      RECT 82.048 31.266 82.152 35.64 ; 
      RECT 81.616 31.266 81.72 35.64 ; 
      RECT 81.184 31.266 81.288 35.64 ; 
      RECT 80.752 31.266 80.856 35.64 ; 
      RECT 80.32 31.266 80.424 35.64 ; 
      RECT 79.888 31.266 79.992 35.64 ; 
      RECT 79.456 31.266 79.56 35.64 ; 
      RECT 79.024 31.266 79.128 35.64 ; 
      RECT 78.592 31.266 78.696 35.64 ; 
      RECT 78.16 31.266 78.264 35.64 ; 
      RECT 77.728 31.266 77.832 35.64 ; 
      RECT 77.296 31.266 77.4 35.64 ; 
      RECT 76.864 31.266 76.968 35.64 ; 
      RECT 76.432 31.266 76.536 35.64 ; 
      RECT 76 31.266 76.104 35.64 ; 
      RECT 75.568 31.266 75.672 35.64 ; 
      RECT 75.136 31.266 75.24 35.64 ; 
      RECT 74.704 31.266 74.808 35.64 ; 
      RECT 74.272 31.266 74.376 35.64 ; 
      RECT 73.84 31.266 73.944 35.64 ; 
      RECT 73.408 31.266 73.512 35.64 ; 
      RECT 72.976 31.266 73.08 35.64 ; 
      RECT 72.544 31.266 72.648 35.64 ; 
      RECT 72.112 31.266 72.216 35.64 ; 
      RECT 71.68 31.266 71.784 35.64 ; 
      RECT 71.248 31.266 71.352 35.64 ; 
      RECT 70.816 31.266 70.92 35.64 ; 
      RECT 70.384 31.266 70.488 35.64 ; 
      RECT 69.952 31.266 70.056 35.64 ; 
      RECT 69.52 31.266 69.624 35.64 ; 
      RECT 69.088 31.266 69.192 35.64 ; 
      RECT 68.656 31.266 68.76 35.64 ; 
      RECT 68.224 31.266 68.328 35.64 ; 
      RECT 67.792 31.266 67.896 35.64 ; 
      RECT 67.36 31.266 67.464 35.64 ; 
      RECT 66.928 31.266 67.032 35.64 ; 
      RECT 66.496 31.266 66.6 35.64 ; 
      RECT 66.064 31.266 66.168 35.64 ; 
      RECT 65.632 31.266 65.736 35.64 ; 
      RECT 65.2 31.266 65.304 35.64 ; 
      RECT 64.348 31.266 64.656 35.64 ; 
      RECT 56.776 31.266 57.084 35.64 ; 
      RECT 56.128 31.266 56.232 35.64 ; 
      RECT 55.696 31.266 55.8 35.64 ; 
      RECT 55.264 31.266 55.368 35.64 ; 
      RECT 54.832 31.266 54.936 35.64 ; 
      RECT 54.4 31.266 54.504 35.64 ; 
      RECT 53.968 31.266 54.072 35.64 ; 
      RECT 53.536 31.266 53.64 35.64 ; 
      RECT 53.104 31.266 53.208 35.64 ; 
      RECT 52.672 31.266 52.776 35.64 ; 
      RECT 52.24 31.266 52.344 35.64 ; 
      RECT 51.808 31.266 51.912 35.64 ; 
      RECT 51.376 31.266 51.48 35.64 ; 
      RECT 50.944 31.266 51.048 35.64 ; 
      RECT 50.512 31.266 50.616 35.64 ; 
      RECT 50.08 31.266 50.184 35.64 ; 
      RECT 49.648 31.266 49.752 35.64 ; 
      RECT 49.216 31.266 49.32 35.64 ; 
      RECT 48.784 31.266 48.888 35.64 ; 
      RECT 48.352 31.266 48.456 35.64 ; 
      RECT 47.92 31.266 48.024 35.64 ; 
      RECT 47.488 31.266 47.592 35.64 ; 
      RECT 47.056 31.266 47.16 35.64 ; 
      RECT 46.624 31.266 46.728 35.64 ; 
      RECT 46.192 31.266 46.296 35.64 ; 
      RECT 45.76 31.266 45.864 35.64 ; 
      RECT 45.328 31.266 45.432 35.64 ; 
      RECT 44.896 31.266 45 35.64 ; 
      RECT 44.464 31.266 44.568 35.64 ; 
      RECT 44.032 31.266 44.136 35.64 ; 
      RECT 43.6 31.266 43.704 35.64 ; 
      RECT 43.168 31.266 43.272 35.64 ; 
      RECT 42.736 31.266 42.84 35.64 ; 
      RECT 42.304 31.266 42.408 35.64 ; 
      RECT 41.872 31.266 41.976 35.64 ; 
      RECT 41.44 31.266 41.544 35.64 ; 
      RECT 41.008 31.266 41.112 35.64 ; 
      RECT 40.576 31.266 40.68 35.64 ; 
      RECT 40.144 31.266 40.248 35.64 ; 
      RECT 39.712 31.266 39.816 35.64 ; 
      RECT 39.28 31.266 39.384 35.64 ; 
      RECT 38.848 31.266 38.952 35.64 ; 
      RECT 38.416 31.266 38.52 35.64 ; 
      RECT 37.984 31.266 38.088 35.64 ; 
      RECT 37.552 31.266 37.656 35.64 ; 
      RECT 37.12 31.266 37.224 35.64 ; 
      RECT 36.688 31.266 36.792 35.64 ; 
      RECT 36.256 31.266 36.36 35.64 ; 
      RECT 35.824 31.266 35.928 35.64 ; 
      RECT 35.392 31.266 35.496 35.64 ; 
      RECT 34.96 31.266 35.064 35.64 ; 
      RECT 34.528 31.266 34.632 35.64 ; 
      RECT 34.096 31.266 34.2 35.64 ; 
      RECT 33.664 31.266 33.768 35.64 ; 
      RECT 33.232 31.266 33.336 35.64 ; 
      RECT 32.8 31.266 32.904 35.64 ; 
      RECT 32.368 31.266 32.472 35.64 ; 
      RECT 31.936 31.266 32.04 35.64 ; 
      RECT 31.504 31.266 31.608 35.64 ; 
      RECT 31.072 31.266 31.176 35.64 ; 
      RECT 30.64 31.266 30.744 35.64 ; 
      RECT 30.208 31.266 30.312 35.64 ; 
      RECT 29.776 31.266 29.88 35.64 ; 
      RECT 29.344 31.266 29.448 35.64 ; 
      RECT 28.912 31.266 29.016 35.64 ; 
      RECT 28.48 31.266 28.584 35.64 ; 
      RECT 28.048 31.266 28.152 35.64 ; 
      RECT 27.616 31.266 27.72 35.64 ; 
      RECT 27.184 31.266 27.288 35.64 ; 
      RECT 26.752 31.266 26.856 35.64 ; 
      RECT 26.32 31.266 26.424 35.64 ; 
      RECT 25.888 31.266 25.992 35.64 ; 
      RECT 25.456 31.266 25.56 35.64 ; 
      RECT 25.024 31.266 25.128 35.64 ; 
      RECT 24.592 31.266 24.696 35.64 ; 
      RECT 24.16 31.266 24.264 35.64 ; 
      RECT 23.728 31.266 23.832 35.64 ; 
      RECT 23.296 31.266 23.4 35.64 ; 
      RECT 22.864 31.266 22.968 35.64 ; 
      RECT 22.432 31.266 22.536 35.64 ; 
      RECT 22 31.266 22.104 35.64 ; 
      RECT 21.568 31.266 21.672 35.64 ; 
      RECT 21.136 31.266 21.24 35.64 ; 
      RECT 20.704 31.266 20.808 35.64 ; 
      RECT 20.272 31.266 20.376 35.64 ; 
      RECT 19.84 31.266 19.944 35.64 ; 
      RECT 19.408 31.266 19.512 35.64 ; 
      RECT 18.976 31.266 19.08 35.64 ; 
      RECT 18.544 31.266 18.648 35.64 ; 
      RECT 18.112 31.266 18.216 35.64 ; 
      RECT 17.68 31.266 17.784 35.64 ; 
      RECT 17.248 31.266 17.352 35.64 ; 
      RECT 16.816 31.266 16.92 35.64 ; 
      RECT 16.384 31.266 16.488 35.64 ; 
      RECT 15.952 31.266 16.056 35.64 ; 
      RECT 15.52 31.266 15.624 35.64 ; 
      RECT 15.088 31.266 15.192 35.64 ; 
      RECT 14.656 31.266 14.76 35.64 ; 
      RECT 14.224 31.266 14.328 35.64 ; 
      RECT 13.792 31.266 13.896 35.64 ; 
      RECT 13.36 31.266 13.464 35.64 ; 
      RECT 12.928 31.266 13.032 35.64 ; 
      RECT 12.496 31.266 12.6 35.64 ; 
      RECT 12.064 31.266 12.168 35.64 ; 
      RECT 11.632 31.266 11.736 35.64 ; 
      RECT 11.2 31.266 11.304 35.64 ; 
      RECT 10.768 31.266 10.872 35.64 ; 
      RECT 10.336 31.266 10.44 35.64 ; 
      RECT 9.904 31.266 10.008 35.64 ; 
      RECT 9.472 31.266 9.576 35.64 ; 
      RECT 9.04 31.266 9.144 35.64 ; 
      RECT 8.608 31.266 8.712 35.64 ; 
      RECT 8.176 31.266 8.28 35.64 ; 
      RECT 7.744 31.266 7.848 35.64 ; 
      RECT 7.312 31.266 7.416 35.64 ; 
      RECT 6.88 31.266 6.984 35.64 ; 
      RECT 6.448 31.266 6.552 35.64 ; 
      RECT 6.016 31.266 6.12 35.64 ; 
      RECT 5.584 31.266 5.688 35.64 ; 
      RECT 5.152 31.266 5.256 35.64 ; 
      RECT 4.72 31.266 4.824 35.64 ; 
      RECT 4.288 31.266 4.392 35.64 ; 
      RECT 3.856 31.266 3.96 35.64 ; 
      RECT 3.424 31.266 3.528 35.64 ; 
      RECT 2.992 31.266 3.096 35.64 ; 
      RECT 2.56 31.266 2.664 35.64 ; 
      RECT 2.128 31.266 2.232 35.64 ; 
      RECT 1.696 31.266 1.8 35.64 ; 
      RECT 1.264 31.266 1.368 35.64 ; 
      RECT 0.832 31.266 0.936 35.64 ; 
      RECT 0.02 31.266 0.36 35.64 ; 
      RECT 62.212 35.586 62.724 39.96 ; 
      RECT 62.156 38.248 62.724 39.538 ; 
      RECT 61.276 37.156 61.812 39.96 ; 
      RECT 61.184 38.496 61.812 39.528 ; 
      RECT 61.276 35.586 61.668 39.96 ; 
      RECT 61.276 36.07 61.724 37.028 ; 
      RECT 61.276 35.586 61.812 35.942 ; 
      RECT 60.376 37.388 60.912 39.96 ; 
      RECT 60.376 35.586 60.768 39.96 ; 
      RECT 58.708 35.586 59.04 39.96 ; 
      RECT 58.708 35.94 59.096 39.682 ; 
      RECT 121.072 35.586 121.412 39.96 ; 
      RECT 120.496 35.586 120.6 39.96 ; 
      RECT 120.064 35.586 120.168 39.96 ; 
      RECT 119.632 35.586 119.736 39.96 ; 
      RECT 119.2 35.586 119.304 39.96 ; 
      RECT 118.768 35.586 118.872 39.96 ; 
      RECT 118.336 35.586 118.44 39.96 ; 
      RECT 117.904 35.586 118.008 39.96 ; 
      RECT 117.472 35.586 117.576 39.96 ; 
      RECT 117.04 35.586 117.144 39.96 ; 
      RECT 116.608 35.586 116.712 39.96 ; 
      RECT 116.176 35.586 116.28 39.96 ; 
      RECT 115.744 35.586 115.848 39.96 ; 
      RECT 115.312 35.586 115.416 39.96 ; 
      RECT 114.88 35.586 114.984 39.96 ; 
      RECT 114.448 35.586 114.552 39.96 ; 
      RECT 114.016 35.586 114.12 39.96 ; 
      RECT 113.584 35.586 113.688 39.96 ; 
      RECT 113.152 35.586 113.256 39.96 ; 
      RECT 112.72 35.586 112.824 39.96 ; 
      RECT 112.288 35.586 112.392 39.96 ; 
      RECT 111.856 35.586 111.96 39.96 ; 
      RECT 111.424 35.586 111.528 39.96 ; 
      RECT 110.992 35.586 111.096 39.96 ; 
      RECT 110.56 35.586 110.664 39.96 ; 
      RECT 110.128 35.586 110.232 39.96 ; 
      RECT 109.696 35.586 109.8 39.96 ; 
      RECT 109.264 35.586 109.368 39.96 ; 
      RECT 108.832 35.586 108.936 39.96 ; 
      RECT 108.4 35.586 108.504 39.96 ; 
      RECT 107.968 35.586 108.072 39.96 ; 
      RECT 107.536 35.586 107.64 39.96 ; 
      RECT 107.104 35.586 107.208 39.96 ; 
      RECT 106.672 35.586 106.776 39.96 ; 
      RECT 106.24 35.586 106.344 39.96 ; 
      RECT 105.808 35.586 105.912 39.96 ; 
      RECT 105.376 35.586 105.48 39.96 ; 
      RECT 104.944 35.586 105.048 39.96 ; 
      RECT 104.512 35.586 104.616 39.96 ; 
      RECT 104.08 35.586 104.184 39.96 ; 
      RECT 103.648 35.586 103.752 39.96 ; 
      RECT 103.216 35.586 103.32 39.96 ; 
      RECT 102.784 35.586 102.888 39.96 ; 
      RECT 102.352 35.586 102.456 39.96 ; 
      RECT 101.92 35.586 102.024 39.96 ; 
      RECT 101.488 35.586 101.592 39.96 ; 
      RECT 101.056 35.586 101.16 39.96 ; 
      RECT 100.624 35.586 100.728 39.96 ; 
      RECT 100.192 35.586 100.296 39.96 ; 
      RECT 99.76 35.586 99.864 39.96 ; 
      RECT 99.328 35.586 99.432 39.96 ; 
      RECT 98.896 35.586 99 39.96 ; 
      RECT 98.464 35.586 98.568 39.96 ; 
      RECT 98.032 35.586 98.136 39.96 ; 
      RECT 97.6 35.586 97.704 39.96 ; 
      RECT 97.168 35.586 97.272 39.96 ; 
      RECT 96.736 35.586 96.84 39.96 ; 
      RECT 96.304 35.586 96.408 39.96 ; 
      RECT 95.872 35.586 95.976 39.96 ; 
      RECT 95.44 35.586 95.544 39.96 ; 
      RECT 95.008 35.586 95.112 39.96 ; 
      RECT 94.576 35.586 94.68 39.96 ; 
      RECT 94.144 35.586 94.248 39.96 ; 
      RECT 93.712 35.586 93.816 39.96 ; 
      RECT 93.28 35.586 93.384 39.96 ; 
      RECT 92.848 35.586 92.952 39.96 ; 
      RECT 92.416 35.586 92.52 39.96 ; 
      RECT 91.984 35.586 92.088 39.96 ; 
      RECT 91.552 35.586 91.656 39.96 ; 
      RECT 91.12 35.586 91.224 39.96 ; 
      RECT 90.688 35.586 90.792 39.96 ; 
      RECT 90.256 35.586 90.36 39.96 ; 
      RECT 89.824 35.586 89.928 39.96 ; 
      RECT 89.392 35.586 89.496 39.96 ; 
      RECT 88.96 35.586 89.064 39.96 ; 
      RECT 88.528 35.586 88.632 39.96 ; 
      RECT 88.096 35.586 88.2 39.96 ; 
      RECT 87.664 35.586 87.768 39.96 ; 
      RECT 87.232 35.586 87.336 39.96 ; 
      RECT 86.8 35.586 86.904 39.96 ; 
      RECT 86.368 35.586 86.472 39.96 ; 
      RECT 85.936 35.586 86.04 39.96 ; 
      RECT 85.504 35.586 85.608 39.96 ; 
      RECT 85.072 35.586 85.176 39.96 ; 
      RECT 84.64 35.586 84.744 39.96 ; 
      RECT 84.208 35.586 84.312 39.96 ; 
      RECT 83.776 35.586 83.88 39.96 ; 
      RECT 83.344 35.586 83.448 39.96 ; 
      RECT 82.912 35.586 83.016 39.96 ; 
      RECT 82.48 35.586 82.584 39.96 ; 
      RECT 82.048 35.586 82.152 39.96 ; 
      RECT 81.616 35.586 81.72 39.96 ; 
      RECT 81.184 35.586 81.288 39.96 ; 
      RECT 80.752 35.586 80.856 39.96 ; 
      RECT 80.32 35.586 80.424 39.96 ; 
      RECT 79.888 35.586 79.992 39.96 ; 
      RECT 79.456 35.586 79.56 39.96 ; 
      RECT 79.024 35.586 79.128 39.96 ; 
      RECT 78.592 35.586 78.696 39.96 ; 
      RECT 78.16 35.586 78.264 39.96 ; 
      RECT 77.728 35.586 77.832 39.96 ; 
      RECT 77.296 35.586 77.4 39.96 ; 
      RECT 76.864 35.586 76.968 39.96 ; 
      RECT 76.432 35.586 76.536 39.96 ; 
      RECT 76 35.586 76.104 39.96 ; 
      RECT 75.568 35.586 75.672 39.96 ; 
      RECT 75.136 35.586 75.24 39.96 ; 
      RECT 74.704 35.586 74.808 39.96 ; 
      RECT 74.272 35.586 74.376 39.96 ; 
      RECT 73.84 35.586 73.944 39.96 ; 
      RECT 73.408 35.586 73.512 39.96 ; 
      RECT 72.976 35.586 73.08 39.96 ; 
      RECT 72.544 35.586 72.648 39.96 ; 
      RECT 72.112 35.586 72.216 39.96 ; 
      RECT 71.68 35.586 71.784 39.96 ; 
      RECT 71.248 35.586 71.352 39.96 ; 
      RECT 70.816 35.586 70.92 39.96 ; 
      RECT 70.384 35.586 70.488 39.96 ; 
      RECT 69.952 35.586 70.056 39.96 ; 
      RECT 69.52 35.586 69.624 39.96 ; 
      RECT 69.088 35.586 69.192 39.96 ; 
      RECT 68.656 35.586 68.76 39.96 ; 
      RECT 68.224 35.586 68.328 39.96 ; 
      RECT 67.792 35.586 67.896 39.96 ; 
      RECT 67.36 35.586 67.464 39.96 ; 
      RECT 66.928 35.586 67.032 39.96 ; 
      RECT 66.496 35.586 66.6 39.96 ; 
      RECT 66.064 35.586 66.168 39.96 ; 
      RECT 65.632 35.586 65.736 39.96 ; 
      RECT 65.2 35.586 65.304 39.96 ; 
      RECT 64.348 35.586 64.656 39.96 ; 
      RECT 56.776 35.586 57.084 39.96 ; 
      RECT 56.128 35.586 56.232 39.96 ; 
      RECT 55.696 35.586 55.8 39.96 ; 
      RECT 55.264 35.586 55.368 39.96 ; 
      RECT 54.832 35.586 54.936 39.96 ; 
      RECT 54.4 35.586 54.504 39.96 ; 
      RECT 53.968 35.586 54.072 39.96 ; 
      RECT 53.536 35.586 53.64 39.96 ; 
      RECT 53.104 35.586 53.208 39.96 ; 
      RECT 52.672 35.586 52.776 39.96 ; 
      RECT 52.24 35.586 52.344 39.96 ; 
      RECT 51.808 35.586 51.912 39.96 ; 
      RECT 51.376 35.586 51.48 39.96 ; 
      RECT 50.944 35.586 51.048 39.96 ; 
      RECT 50.512 35.586 50.616 39.96 ; 
      RECT 50.08 35.586 50.184 39.96 ; 
      RECT 49.648 35.586 49.752 39.96 ; 
      RECT 49.216 35.586 49.32 39.96 ; 
      RECT 48.784 35.586 48.888 39.96 ; 
      RECT 48.352 35.586 48.456 39.96 ; 
      RECT 47.92 35.586 48.024 39.96 ; 
      RECT 47.488 35.586 47.592 39.96 ; 
      RECT 47.056 35.586 47.16 39.96 ; 
      RECT 46.624 35.586 46.728 39.96 ; 
      RECT 46.192 35.586 46.296 39.96 ; 
      RECT 45.76 35.586 45.864 39.96 ; 
      RECT 45.328 35.586 45.432 39.96 ; 
      RECT 44.896 35.586 45 39.96 ; 
      RECT 44.464 35.586 44.568 39.96 ; 
      RECT 44.032 35.586 44.136 39.96 ; 
      RECT 43.6 35.586 43.704 39.96 ; 
      RECT 43.168 35.586 43.272 39.96 ; 
      RECT 42.736 35.586 42.84 39.96 ; 
      RECT 42.304 35.586 42.408 39.96 ; 
      RECT 41.872 35.586 41.976 39.96 ; 
      RECT 41.44 35.586 41.544 39.96 ; 
      RECT 41.008 35.586 41.112 39.96 ; 
      RECT 40.576 35.586 40.68 39.96 ; 
      RECT 40.144 35.586 40.248 39.96 ; 
      RECT 39.712 35.586 39.816 39.96 ; 
      RECT 39.28 35.586 39.384 39.96 ; 
      RECT 38.848 35.586 38.952 39.96 ; 
      RECT 38.416 35.586 38.52 39.96 ; 
      RECT 37.984 35.586 38.088 39.96 ; 
      RECT 37.552 35.586 37.656 39.96 ; 
      RECT 37.12 35.586 37.224 39.96 ; 
      RECT 36.688 35.586 36.792 39.96 ; 
      RECT 36.256 35.586 36.36 39.96 ; 
      RECT 35.824 35.586 35.928 39.96 ; 
      RECT 35.392 35.586 35.496 39.96 ; 
      RECT 34.96 35.586 35.064 39.96 ; 
      RECT 34.528 35.586 34.632 39.96 ; 
      RECT 34.096 35.586 34.2 39.96 ; 
      RECT 33.664 35.586 33.768 39.96 ; 
      RECT 33.232 35.586 33.336 39.96 ; 
      RECT 32.8 35.586 32.904 39.96 ; 
      RECT 32.368 35.586 32.472 39.96 ; 
      RECT 31.936 35.586 32.04 39.96 ; 
      RECT 31.504 35.586 31.608 39.96 ; 
      RECT 31.072 35.586 31.176 39.96 ; 
      RECT 30.64 35.586 30.744 39.96 ; 
      RECT 30.208 35.586 30.312 39.96 ; 
      RECT 29.776 35.586 29.88 39.96 ; 
      RECT 29.344 35.586 29.448 39.96 ; 
      RECT 28.912 35.586 29.016 39.96 ; 
      RECT 28.48 35.586 28.584 39.96 ; 
      RECT 28.048 35.586 28.152 39.96 ; 
      RECT 27.616 35.586 27.72 39.96 ; 
      RECT 27.184 35.586 27.288 39.96 ; 
      RECT 26.752 35.586 26.856 39.96 ; 
      RECT 26.32 35.586 26.424 39.96 ; 
      RECT 25.888 35.586 25.992 39.96 ; 
      RECT 25.456 35.586 25.56 39.96 ; 
      RECT 25.024 35.586 25.128 39.96 ; 
      RECT 24.592 35.586 24.696 39.96 ; 
      RECT 24.16 35.586 24.264 39.96 ; 
      RECT 23.728 35.586 23.832 39.96 ; 
      RECT 23.296 35.586 23.4 39.96 ; 
      RECT 22.864 35.586 22.968 39.96 ; 
      RECT 22.432 35.586 22.536 39.96 ; 
      RECT 22 35.586 22.104 39.96 ; 
      RECT 21.568 35.586 21.672 39.96 ; 
      RECT 21.136 35.586 21.24 39.96 ; 
      RECT 20.704 35.586 20.808 39.96 ; 
      RECT 20.272 35.586 20.376 39.96 ; 
      RECT 19.84 35.586 19.944 39.96 ; 
      RECT 19.408 35.586 19.512 39.96 ; 
      RECT 18.976 35.586 19.08 39.96 ; 
      RECT 18.544 35.586 18.648 39.96 ; 
      RECT 18.112 35.586 18.216 39.96 ; 
      RECT 17.68 35.586 17.784 39.96 ; 
      RECT 17.248 35.586 17.352 39.96 ; 
      RECT 16.816 35.586 16.92 39.96 ; 
      RECT 16.384 35.586 16.488 39.96 ; 
      RECT 15.952 35.586 16.056 39.96 ; 
      RECT 15.52 35.586 15.624 39.96 ; 
      RECT 15.088 35.586 15.192 39.96 ; 
      RECT 14.656 35.586 14.76 39.96 ; 
      RECT 14.224 35.586 14.328 39.96 ; 
      RECT 13.792 35.586 13.896 39.96 ; 
      RECT 13.36 35.586 13.464 39.96 ; 
      RECT 12.928 35.586 13.032 39.96 ; 
      RECT 12.496 35.586 12.6 39.96 ; 
      RECT 12.064 35.586 12.168 39.96 ; 
      RECT 11.632 35.586 11.736 39.96 ; 
      RECT 11.2 35.586 11.304 39.96 ; 
      RECT 10.768 35.586 10.872 39.96 ; 
      RECT 10.336 35.586 10.44 39.96 ; 
      RECT 9.904 35.586 10.008 39.96 ; 
      RECT 9.472 35.586 9.576 39.96 ; 
      RECT 9.04 35.586 9.144 39.96 ; 
      RECT 8.608 35.586 8.712 39.96 ; 
      RECT 8.176 35.586 8.28 39.96 ; 
      RECT 7.744 35.586 7.848 39.96 ; 
      RECT 7.312 35.586 7.416 39.96 ; 
      RECT 6.88 35.586 6.984 39.96 ; 
      RECT 6.448 35.586 6.552 39.96 ; 
      RECT 6.016 35.586 6.12 39.96 ; 
      RECT 5.584 35.586 5.688 39.96 ; 
      RECT 5.152 35.586 5.256 39.96 ; 
      RECT 4.72 35.586 4.824 39.96 ; 
      RECT 4.288 35.586 4.392 39.96 ; 
      RECT 3.856 35.586 3.96 39.96 ; 
      RECT 3.424 35.586 3.528 39.96 ; 
      RECT 2.992 35.586 3.096 39.96 ; 
      RECT 2.56 35.586 2.664 39.96 ; 
      RECT 2.128 35.586 2.232 39.96 ; 
      RECT 1.696 35.586 1.8 39.96 ; 
      RECT 1.264 35.586 1.368 39.96 ; 
      RECT 0.832 35.586 0.936 39.96 ; 
      RECT 0.02 35.586 0.36 39.96 ; 
      RECT 56.54 72.904 121.392 74.668 ; 
      RECT 71.012 40.054 121.392 74.668 ; 
      RECT 65.18 46.07 121.392 74.668 ; 
      RECT 70.148 45.29 121.392 74.668 ; 
      RECT 56.54 71.702 64.852 74.668 ; 
      RECT 62.228 45.674 64.852 74.668 ; 
      RECT 56.54 46.502 61.036 74.668 ; 
      RECT 60.788 40.054 61.036 74.668 ; 
      RECT 62.172 66.638 64.852 71.07 ; 
      RECT 65.124 55.226 121.392 69.598 ; 
      RECT 56.54 67.574 61.092 68.622 ; 
      RECT 62.172 56.486 64.852 65.814 ; 
      RECT 56.54 57.998 61.092 63.222 ; 
      RECT 56.54 47.342 61.092 57.822 ; 
      RECT 62.172 45.182 64.636 52.326 ; 
      RECT 56.756 46.262 61.092 47.022 ; 
      RECT 56.756 43.118 61.036 74.668 ; 
      RECT 57.62 42.794 61.036 74.668 ; 
      RECT 56.756 45.182 61.092 46.086 ; 
      RECT 65.828 45.302 121.392 74.668 ; 
      RECT 65.18 40.054 65.5 74.668 ; 
      RECT 56.54 42.794 57.292 46.05 ; 
      RECT 65.18 40.054 66.364 45.666 ; 
      RECT 65.18 44.522 69.82 45.666 ; 
      RECT 70.148 40.054 70.684 74.668 ; 
      RECT 62.228 44.522 64.636 74.668 ; 
      RECT 63.524 40.054 64.852 45.054 ; 
      RECT 65.18 44.522 70.684 44.898 ; 
      RECT 69.284 40.054 121.392 44.886 ; 
      RECT 56.54 44.606 61.092 44.862 ; 
      RECT 68.42 42.986 121.392 44.886 ; 
      RECT 65.18 43.118 68.092 45.666 ; 
      RECT 62.228 43.118 63.196 74.668 ; 
      RECT 57.62 43.022 61.092 44.07 ; 
      RECT 62.372 40.054 64.852 43.686 ; 
      RECT 67.556 40.054 68.956 43.542 ; 
      RECT 65.18 42.794 67.228 45.666 ; 
      RECT 66.692 40.054 67.228 74.668 ; 
      RECT 57.62 40.054 60.46 74.668 ; 
      RECT 56.9 40.054 57.292 74.668 ; 
      RECT 66.692 40.054 68.956 42.594 ; 
      RECT 62.228 40.054 64.852 42.594 ; 
      RECT 56.9 40.054 60.46 42.594 ; 
      RECT 66.692 40.054 121.392 42.582 ; 
      RECT 62.172 41.942 64.852 42.558 ; 
      RECT 65.18 40.054 121.392 41.526 ; 
      RECT 56.54 40.054 61.036 41.526 ; 
      RECT 56.54 40.054 64.852 40.714 ; 
      RECT 71.028 39.294 71.1 74.668 ; 
      RECT 70.596 39.294 70.668 74.668 ; 
      RECT 70.164 39.294 70.236 74.668 ; 
      RECT 69.732 39.294 69.804 74.668 ; 
      RECT 69.3 39.294 69.372 74.668 ; 
      RECT 68.868 39.294 68.94 74.668 ; 
      RECT 68.436 39.294 68.508 74.668 ; 
      RECT 68.004 39.294 68.076 74.668 ; 
      RECT 67.572 39.294 67.644 74.668 ; 
      RECT 67.14 39.294 67.212 74.668 ; 
      RECT 66.708 39.294 66.78 74.668 ; 
      RECT 66.276 39.294 66.348 74.668 ; 
      RECT 65.844 39.294 65.916 74.668 ; 
      RECT 65.412 39.294 65.484 74.668 ; 
      RECT 0 45.29 56.068 74.668 ; 
      RECT 0 56.446 56.124 56.778 ; 
      RECT 55.028 40.054 56.212 55.092 ; 
      RECT 51.572 43.766 54.7 74.668 ; 
      RECT 0 40.054 51.244 74.668 ; 
      RECT 54.164 40.054 56.212 44.886 ; 
      RECT 0 42.986 53.836 44.886 ; 
      RECT 53.3 40.054 53.836 74.668 ; 
      RECT 52.436 42.794 53.836 74.668 ; 
      RECT 0 40.054 52.108 44.886 ; 
      RECT 52.436 40.054 52.972 74.668 ; 
      RECT 53.3 40.054 56.212 42.594 ; 
      RECT 0 40.054 52.972 42.582 ; 
      RECT 0 40.054 56.212 41.526 ; 
      RECT 53.316 39.948 53.388 74.668 ; 
      RECT 52.884 39.948 52.956 74.668 ; 
        RECT 62.212 72.414 62.724 76.788 ; 
        RECT 62.156 75.076 62.724 76.366 ; 
        RECT 61.276 73.984 61.812 76.788 ; 
        RECT 61.184 75.324 61.812 76.356 ; 
        RECT 61.276 72.414 61.668 76.788 ; 
        RECT 61.276 72.898 61.724 73.856 ; 
        RECT 61.276 72.414 61.812 72.77 ; 
        RECT 60.376 74.216 60.912 76.788 ; 
        RECT 60.376 72.414 60.768 76.788 ; 
        RECT 58.708 72.414 59.04 76.788 ; 
        RECT 58.708 72.768 59.096 76.51 ; 
        RECT 121.072 72.414 121.412 76.788 ; 
        RECT 120.496 72.414 120.6 76.788 ; 
        RECT 120.064 72.414 120.168 76.788 ; 
        RECT 119.632 72.414 119.736 76.788 ; 
        RECT 119.2 72.414 119.304 76.788 ; 
        RECT 118.768 72.414 118.872 76.788 ; 
        RECT 118.336 72.414 118.44 76.788 ; 
        RECT 117.904 72.414 118.008 76.788 ; 
        RECT 117.472 72.414 117.576 76.788 ; 
        RECT 117.04 72.414 117.144 76.788 ; 
        RECT 116.608 72.414 116.712 76.788 ; 
        RECT 116.176 72.414 116.28 76.788 ; 
        RECT 115.744 72.414 115.848 76.788 ; 
        RECT 115.312 72.414 115.416 76.788 ; 
        RECT 114.88 72.414 114.984 76.788 ; 
        RECT 114.448 72.414 114.552 76.788 ; 
        RECT 114.016 72.414 114.12 76.788 ; 
        RECT 113.584 72.414 113.688 76.788 ; 
        RECT 113.152 72.414 113.256 76.788 ; 
        RECT 112.72 72.414 112.824 76.788 ; 
        RECT 112.288 72.414 112.392 76.788 ; 
        RECT 111.856 72.414 111.96 76.788 ; 
        RECT 111.424 72.414 111.528 76.788 ; 
        RECT 110.992 72.414 111.096 76.788 ; 
        RECT 110.56 72.414 110.664 76.788 ; 
        RECT 110.128 72.414 110.232 76.788 ; 
        RECT 109.696 72.414 109.8 76.788 ; 
        RECT 109.264 72.414 109.368 76.788 ; 
        RECT 108.832 72.414 108.936 76.788 ; 
        RECT 108.4 72.414 108.504 76.788 ; 
        RECT 107.968 72.414 108.072 76.788 ; 
        RECT 107.536 72.414 107.64 76.788 ; 
        RECT 107.104 72.414 107.208 76.788 ; 
        RECT 106.672 72.414 106.776 76.788 ; 
        RECT 106.24 72.414 106.344 76.788 ; 
        RECT 105.808 72.414 105.912 76.788 ; 
        RECT 105.376 72.414 105.48 76.788 ; 
        RECT 104.944 72.414 105.048 76.788 ; 
        RECT 104.512 72.414 104.616 76.788 ; 
        RECT 104.08 72.414 104.184 76.788 ; 
        RECT 103.648 72.414 103.752 76.788 ; 
        RECT 103.216 72.414 103.32 76.788 ; 
        RECT 102.784 72.414 102.888 76.788 ; 
        RECT 102.352 72.414 102.456 76.788 ; 
        RECT 101.92 72.414 102.024 76.788 ; 
        RECT 101.488 72.414 101.592 76.788 ; 
        RECT 101.056 72.414 101.16 76.788 ; 
        RECT 100.624 72.414 100.728 76.788 ; 
        RECT 100.192 72.414 100.296 76.788 ; 
        RECT 99.76 72.414 99.864 76.788 ; 
        RECT 99.328 72.414 99.432 76.788 ; 
        RECT 98.896 72.414 99 76.788 ; 
        RECT 98.464 72.414 98.568 76.788 ; 
        RECT 98.032 72.414 98.136 76.788 ; 
        RECT 97.6 72.414 97.704 76.788 ; 
        RECT 97.168 72.414 97.272 76.788 ; 
        RECT 96.736 72.414 96.84 76.788 ; 
        RECT 96.304 72.414 96.408 76.788 ; 
        RECT 95.872 72.414 95.976 76.788 ; 
        RECT 95.44 72.414 95.544 76.788 ; 
        RECT 95.008 72.414 95.112 76.788 ; 
        RECT 94.576 72.414 94.68 76.788 ; 
        RECT 94.144 72.414 94.248 76.788 ; 
        RECT 93.712 72.414 93.816 76.788 ; 
        RECT 93.28 72.414 93.384 76.788 ; 
        RECT 92.848 72.414 92.952 76.788 ; 
        RECT 92.416 72.414 92.52 76.788 ; 
        RECT 91.984 72.414 92.088 76.788 ; 
        RECT 91.552 72.414 91.656 76.788 ; 
        RECT 91.12 72.414 91.224 76.788 ; 
        RECT 90.688 72.414 90.792 76.788 ; 
        RECT 90.256 72.414 90.36 76.788 ; 
        RECT 89.824 72.414 89.928 76.788 ; 
        RECT 89.392 72.414 89.496 76.788 ; 
        RECT 88.96 72.414 89.064 76.788 ; 
        RECT 88.528 72.414 88.632 76.788 ; 
        RECT 88.096 72.414 88.2 76.788 ; 
        RECT 87.664 72.414 87.768 76.788 ; 
        RECT 87.232 72.414 87.336 76.788 ; 
        RECT 86.8 72.414 86.904 76.788 ; 
        RECT 86.368 72.414 86.472 76.788 ; 
        RECT 85.936 72.414 86.04 76.788 ; 
        RECT 85.504 72.414 85.608 76.788 ; 
        RECT 85.072 72.414 85.176 76.788 ; 
        RECT 84.64 72.414 84.744 76.788 ; 
        RECT 84.208 72.414 84.312 76.788 ; 
        RECT 83.776 72.414 83.88 76.788 ; 
        RECT 83.344 72.414 83.448 76.788 ; 
        RECT 82.912 72.414 83.016 76.788 ; 
        RECT 82.48 72.414 82.584 76.788 ; 
        RECT 82.048 72.414 82.152 76.788 ; 
        RECT 81.616 72.414 81.72 76.788 ; 
        RECT 81.184 72.414 81.288 76.788 ; 
        RECT 80.752 72.414 80.856 76.788 ; 
        RECT 80.32 72.414 80.424 76.788 ; 
        RECT 79.888 72.414 79.992 76.788 ; 
        RECT 79.456 72.414 79.56 76.788 ; 
        RECT 79.024 72.414 79.128 76.788 ; 
        RECT 78.592 72.414 78.696 76.788 ; 
        RECT 78.16 72.414 78.264 76.788 ; 
        RECT 77.728 72.414 77.832 76.788 ; 
        RECT 77.296 72.414 77.4 76.788 ; 
        RECT 76.864 72.414 76.968 76.788 ; 
        RECT 76.432 72.414 76.536 76.788 ; 
        RECT 76 72.414 76.104 76.788 ; 
        RECT 75.568 72.414 75.672 76.788 ; 
        RECT 75.136 72.414 75.24 76.788 ; 
        RECT 74.704 72.414 74.808 76.788 ; 
        RECT 74.272 72.414 74.376 76.788 ; 
        RECT 73.84 72.414 73.944 76.788 ; 
        RECT 73.408 72.414 73.512 76.788 ; 
        RECT 72.976 72.414 73.08 76.788 ; 
        RECT 72.544 72.414 72.648 76.788 ; 
        RECT 72.112 72.414 72.216 76.788 ; 
        RECT 71.68 72.414 71.784 76.788 ; 
        RECT 71.248 72.414 71.352 76.788 ; 
        RECT 70.816 72.414 70.92 76.788 ; 
        RECT 70.384 72.414 70.488 76.788 ; 
        RECT 69.952 72.414 70.056 76.788 ; 
        RECT 69.52 72.414 69.624 76.788 ; 
        RECT 69.088 72.414 69.192 76.788 ; 
        RECT 68.656 72.414 68.76 76.788 ; 
        RECT 68.224 72.414 68.328 76.788 ; 
        RECT 67.792 72.414 67.896 76.788 ; 
        RECT 67.36 72.414 67.464 76.788 ; 
        RECT 66.928 72.414 67.032 76.788 ; 
        RECT 66.496 72.414 66.6 76.788 ; 
        RECT 66.064 72.414 66.168 76.788 ; 
        RECT 65.632 72.414 65.736 76.788 ; 
        RECT 65.2 72.414 65.304 76.788 ; 
        RECT 64.348 72.414 64.656 76.788 ; 
        RECT 56.776 72.414 57.084 76.788 ; 
        RECT 56.128 72.414 56.232 76.788 ; 
        RECT 55.696 72.414 55.8 76.788 ; 
        RECT 55.264 72.414 55.368 76.788 ; 
        RECT 54.832 72.414 54.936 76.788 ; 
        RECT 54.4 72.414 54.504 76.788 ; 
        RECT 53.968 72.414 54.072 76.788 ; 
        RECT 53.536 72.414 53.64 76.788 ; 
        RECT 53.104 72.414 53.208 76.788 ; 
        RECT 52.672 72.414 52.776 76.788 ; 
        RECT 52.24 72.414 52.344 76.788 ; 
        RECT 51.808 72.414 51.912 76.788 ; 
        RECT 51.376 72.414 51.48 76.788 ; 
        RECT 50.944 72.414 51.048 76.788 ; 
        RECT 50.512 72.414 50.616 76.788 ; 
        RECT 50.08 72.414 50.184 76.788 ; 
        RECT 49.648 72.414 49.752 76.788 ; 
        RECT 49.216 72.414 49.32 76.788 ; 
        RECT 48.784 72.414 48.888 76.788 ; 
        RECT 48.352 72.414 48.456 76.788 ; 
        RECT 47.92 72.414 48.024 76.788 ; 
        RECT 47.488 72.414 47.592 76.788 ; 
        RECT 47.056 72.414 47.16 76.788 ; 
        RECT 46.624 72.414 46.728 76.788 ; 
        RECT 46.192 72.414 46.296 76.788 ; 
        RECT 45.76 72.414 45.864 76.788 ; 
        RECT 45.328 72.414 45.432 76.788 ; 
        RECT 44.896 72.414 45 76.788 ; 
        RECT 44.464 72.414 44.568 76.788 ; 
        RECT 44.032 72.414 44.136 76.788 ; 
        RECT 43.6 72.414 43.704 76.788 ; 
        RECT 43.168 72.414 43.272 76.788 ; 
        RECT 42.736 72.414 42.84 76.788 ; 
        RECT 42.304 72.414 42.408 76.788 ; 
        RECT 41.872 72.414 41.976 76.788 ; 
        RECT 41.44 72.414 41.544 76.788 ; 
        RECT 41.008 72.414 41.112 76.788 ; 
        RECT 40.576 72.414 40.68 76.788 ; 
        RECT 40.144 72.414 40.248 76.788 ; 
        RECT 39.712 72.414 39.816 76.788 ; 
        RECT 39.28 72.414 39.384 76.788 ; 
        RECT 38.848 72.414 38.952 76.788 ; 
        RECT 38.416 72.414 38.52 76.788 ; 
        RECT 37.984 72.414 38.088 76.788 ; 
        RECT 37.552 72.414 37.656 76.788 ; 
        RECT 37.12 72.414 37.224 76.788 ; 
        RECT 36.688 72.414 36.792 76.788 ; 
        RECT 36.256 72.414 36.36 76.788 ; 
        RECT 35.824 72.414 35.928 76.788 ; 
        RECT 35.392 72.414 35.496 76.788 ; 
        RECT 34.96 72.414 35.064 76.788 ; 
        RECT 34.528 72.414 34.632 76.788 ; 
        RECT 34.096 72.414 34.2 76.788 ; 
        RECT 33.664 72.414 33.768 76.788 ; 
        RECT 33.232 72.414 33.336 76.788 ; 
        RECT 32.8 72.414 32.904 76.788 ; 
        RECT 32.368 72.414 32.472 76.788 ; 
        RECT 31.936 72.414 32.04 76.788 ; 
        RECT 31.504 72.414 31.608 76.788 ; 
        RECT 31.072 72.414 31.176 76.788 ; 
        RECT 30.64 72.414 30.744 76.788 ; 
        RECT 30.208 72.414 30.312 76.788 ; 
        RECT 29.776 72.414 29.88 76.788 ; 
        RECT 29.344 72.414 29.448 76.788 ; 
        RECT 28.912 72.414 29.016 76.788 ; 
        RECT 28.48 72.414 28.584 76.788 ; 
        RECT 28.048 72.414 28.152 76.788 ; 
        RECT 27.616 72.414 27.72 76.788 ; 
        RECT 27.184 72.414 27.288 76.788 ; 
        RECT 26.752 72.414 26.856 76.788 ; 
        RECT 26.32 72.414 26.424 76.788 ; 
        RECT 25.888 72.414 25.992 76.788 ; 
        RECT 25.456 72.414 25.56 76.788 ; 
        RECT 25.024 72.414 25.128 76.788 ; 
        RECT 24.592 72.414 24.696 76.788 ; 
        RECT 24.16 72.414 24.264 76.788 ; 
        RECT 23.728 72.414 23.832 76.788 ; 
        RECT 23.296 72.414 23.4 76.788 ; 
        RECT 22.864 72.414 22.968 76.788 ; 
        RECT 22.432 72.414 22.536 76.788 ; 
        RECT 22 72.414 22.104 76.788 ; 
        RECT 21.568 72.414 21.672 76.788 ; 
        RECT 21.136 72.414 21.24 76.788 ; 
        RECT 20.704 72.414 20.808 76.788 ; 
        RECT 20.272 72.414 20.376 76.788 ; 
        RECT 19.84 72.414 19.944 76.788 ; 
        RECT 19.408 72.414 19.512 76.788 ; 
        RECT 18.976 72.414 19.08 76.788 ; 
        RECT 18.544 72.414 18.648 76.788 ; 
        RECT 18.112 72.414 18.216 76.788 ; 
        RECT 17.68 72.414 17.784 76.788 ; 
        RECT 17.248 72.414 17.352 76.788 ; 
        RECT 16.816 72.414 16.92 76.788 ; 
        RECT 16.384 72.414 16.488 76.788 ; 
        RECT 15.952 72.414 16.056 76.788 ; 
        RECT 15.52 72.414 15.624 76.788 ; 
        RECT 15.088 72.414 15.192 76.788 ; 
        RECT 14.656 72.414 14.76 76.788 ; 
        RECT 14.224 72.414 14.328 76.788 ; 
        RECT 13.792 72.414 13.896 76.788 ; 
        RECT 13.36 72.414 13.464 76.788 ; 
        RECT 12.928 72.414 13.032 76.788 ; 
        RECT 12.496 72.414 12.6 76.788 ; 
        RECT 12.064 72.414 12.168 76.788 ; 
        RECT 11.632 72.414 11.736 76.788 ; 
        RECT 11.2 72.414 11.304 76.788 ; 
        RECT 10.768 72.414 10.872 76.788 ; 
        RECT 10.336 72.414 10.44 76.788 ; 
        RECT 9.904 72.414 10.008 76.788 ; 
        RECT 9.472 72.414 9.576 76.788 ; 
        RECT 9.04 72.414 9.144 76.788 ; 
        RECT 8.608 72.414 8.712 76.788 ; 
        RECT 8.176 72.414 8.28 76.788 ; 
        RECT 7.744 72.414 7.848 76.788 ; 
        RECT 7.312 72.414 7.416 76.788 ; 
        RECT 6.88 72.414 6.984 76.788 ; 
        RECT 6.448 72.414 6.552 76.788 ; 
        RECT 6.016 72.414 6.12 76.788 ; 
        RECT 5.584 72.414 5.688 76.788 ; 
        RECT 5.152 72.414 5.256 76.788 ; 
        RECT 4.72 72.414 4.824 76.788 ; 
        RECT 4.288 72.414 4.392 76.788 ; 
        RECT 3.856 72.414 3.96 76.788 ; 
        RECT 3.424 72.414 3.528 76.788 ; 
        RECT 2.992 72.414 3.096 76.788 ; 
        RECT 2.56 72.414 2.664 76.788 ; 
        RECT 2.128 72.414 2.232 76.788 ; 
        RECT 1.696 72.414 1.8 76.788 ; 
        RECT 1.264 72.414 1.368 76.788 ; 
        RECT 0.832 72.414 0.936 76.788 ; 
        RECT 0.02 72.414 0.36 76.788 ; 
        RECT 62.212 76.734 62.724 81.108 ; 
        RECT 62.156 79.396 62.724 80.686 ; 
        RECT 61.276 78.304 61.812 81.108 ; 
        RECT 61.184 79.644 61.812 80.676 ; 
        RECT 61.276 76.734 61.668 81.108 ; 
        RECT 61.276 77.218 61.724 78.176 ; 
        RECT 61.276 76.734 61.812 77.09 ; 
        RECT 60.376 78.536 60.912 81.108 ; 
        RECT 60.376 76.734 60.768 81.108 ; 
        RECT 58.708 76.734 59.04 81.108 ; 
        RECT 58.708 77.088 59.096 80.83 ; 
        RECT 121.072 76.734 121.412 81.108 ; 
        RECT 120.496 76.734 120.6 81.108 ; 
        RECT 120.064 76.734 120.168 81.108 ; 
        RECT 119.632 76.734 119.736 81.108 ; 
        RECT 119.2 76.734 119.304 81.108 ; 
        RECT 118.768 76.734 118.872 81.108 ; 
        RECT 118.336 76.734 118.44 81.108 ; 
        RECT 117.904 76.734 118.008 81.108 ; 
        RECT 117.472 76.734 117.576 81.108 ; 
        RECT 117.04 76.734 117.144 81.108 ; 
        RECT 116.608 76.734 116.712 81.108 ; 
        RECT 116.176 76.734 116.28 81.108 ; 
        RECT 115.744 76.734 115.848 81.108 ; 
        RECT 115.312 76.734 115.416 81.108 ; 
        RECT 114.88 76.734 114.984 81.108 ; 
        RECT 114.448 76.734 114.552 81.108 ; 
        RECT 114.016 76.734 114.12 81.108 ; 
        RECT 113.584 76.734 113.688 81.108 ; 
        RECT 113.152 76.734 113.256 81.108 ; 
        RECT 112.72 76.734 112.824 81.108 ; 
        RECT 112.288 76.734 112.392 81.108 ; 
        RECT 111.856 76.734 111.96 81.108 ; 
        RECT 111.424 76.734 111.528 81.108 ; 
        RECT 110.992 76.734 111.096 81.108 ; 
        RECT 110.56 76.734 110.664 81.108 ; 
        RECT 110.128 76.734 110.232 81.108 ; 
        RECT 109.696 76.734 109.8 81.108 ; 
        RECT 109.264 76.734 109.368 81.108 ; 
        RECT 108.832 76.734 108.936 81.108 ; 
        RECT 108.4 76.734 108.504 81.108 ; 
        RECT 107.968 76.734 108.072 81.108 ; 
        RECT 107.536 76.734 107.64 81.108 ; 
        RECT 107.104 76.734 107.208 81.108 ; 
        RECT 106.672 76.734 106.776 81.108 ; 
        RECT 106.24 76.734 106.344 81.108 ; 
        RECT 105.808 76.734 105.912 81.108 ; 
        RECT 105.376 76.734 105.48 81.108 ; 
        RECT 104.944 76.734 105.048 81.108 ; 
        RECT 104.512 76.734 104.616 81.108 ; 
        RECT 104.08 76.734 104.184 81.108 ; 
        RECT 103.648 76.734 103.752 81.108 ; 
        RECT 103.216 76.734 103.32 81.108 ; 
        RECT 102.784 76.734 102.888 81.108 ; 
        RECT 102.352 76.734 102.456 81.108 ; 
        RECT 101.92 76.734 102.024 81.108 ; 
        RECT 101.488 76.734 101.592 81.108 ; 
        RECT 101.056 76.734 101.16 81.108 ; 
        RECT 100.624 76.734 100.728 81.108 ; 
        RECT 100.192 76.734 100.296 81.108 ; 
        RECT 99.76 76.734 99.864 81.108 ; 
        RECT 99.328 76.734 99.432 81.108 ; 
        RECT 98.896 76.734 99 81.108 ; 
        RECT 98.464 76.734 98.568 81.108 ; 
        RECT 98.032 76.734 98.136 81.108 ; 
        RECT 97.6 76.734 97.704 81.108 ; 
        RECT 97.168 76.734 97.272 81.108 ; 
        RECT 96.736 76.734 96.84 81.108 ; 
        RECT 96.304 76.734 96.408 81.108 ; 
        RECT 95.872 76.734 95.976 81.108 ; 
        RECT 95.44 76.734 95.544 81.108 ; 
        RECT 95.008 76.734 95.112 81.108 ; 
        RECT 94.576 76.734 94.68 81.108 ; 
        RECT 94.144 76.734 94.248 81.108 ; 
        RECT 93.712 76.734 93.816 81.108 ; 
        RECT 93.28 76.734 93.384 81.108 ; 
        RECT 92.848 76.734 92.952 81.108 ; 
        RECT 92.416 76.734 92.52 81.108 ; 
        RECT 91.984 76.734 92.088 81.108 ; 
        RECT 91.552 76.734 91.656 81.108 ; 
        RECT 91.12 76.734 91.224 81.108 ; 
        RECT 90.688 76.734 90.792 81.108 ; 
        RECT 90.256 76.734 90.36 81.108 ; 
        RECT 89.824 76.734 89.928 81.108 ; 
        RECT 89.392 76.734 89.496 81.108 ; 
        RECT 88.96 76.734 89.064 81.108 ; 
        RECT 88.528 76.734 88.632 81.108 ; 
        RECT 88.096 76.734 88.2 81.108 ; 
        RECT 87.664 76.734 87.768 81.108 ; 
        RECT 87.232 76.734 87.336 81.108 ; 
        RECT 86.8 76.734 86.904 81.108 ; 
        RECT 86.368 76.734 86.472 81.108 ; 
        RECT 85.936 76.734 86.04 81.108 ; 
        RECT 85.504 76.734 85.608 81.108 ; 
        RECT 85.072 76.734 85.176 81.108 ; 
        RECT 84.64 76.734 84.744 81.108 ; 
        RECT 84.208 76.734 84.312 81.108 ; 
        RECT 83.776 76.734 83.88 81.108 ; 
        RECT 83.344 76.734 83.448 81.108 ; 
        RECT 82.912 76.734 83.016 81.108 ; 
        RECT 82.48 76.734 82.584 81.108 ; 
        RECT 82.048 76.734 82.152 81.108 ; 
        RECT 81.616 76.734 81.72 81.108 ; 
        RECT 81.184 76.734 81.288 81.108 ; 
        RECT 80.752 76.734 80.856 81.108 ; 
        RECT 80.32 76.734 80.424 81.108 ; 
        RECT 79.888 76.734 79.992 81.108 ; 
        RECT 79.456 76.734 79.56 81.108 ; 
        RECT 79.024 76.734 79.128 81.108 ; 
        RECT 78.592 76.734 78.696 81.108 ; 
        RECT 78.16 76.734 78.264 81.108 ; 
        RECT 77.728 76.734 77.832 81.108 ; 
        RECT 77.296 76.734 77.4 81.108 ; 
        RECT 76.864 76.734 76.968 81.108 ; 
        RECT 76.432 76.734 76.536 81.108 ; 
        RECT 76 76.734 76.104 81.108 ; 
        RECT 75.568 76.734 75.672 81.108 ; 
        RECT 75.136 76.734 75.24 81.108 ; 
        RECT 74.704 76.734 74.808 81.108 ; 
        RECT 74.272 76.734 74.376 81.108 ; 
        RECT 73.84 76.734 73.944 81.108 ; 
        RECT 73.408 76.734 73.512 81.108 ; 
        RECT 72.976 76.734 73.08 81.108 ; 
        RECT 72.544 76.734 72.648 81.108 ; 
        RECT 72.112 76.734 72.216 81.108 ; 
        RECT 71.68 76.734 71.784 81.108 ; 
        RECT 71.248 76.734 71.352 81.108 ; 
        RECT 70.816 76.734 70.92 81.108 ; 
        RECT 70.384 76.734 70.488 81.108 ; 
        RECT 69.952 76.734 70.056 81.108 ; 
        RECT 69.52 76.734 69.624 81.108 ; 
        RECT 69.088 76.734 69.192 81.108 ; 
        RECT 68.656 76.734 68.76 81.108 ; 
        RECT 68.224 76.734 68.328 81.108 ; 
        RECT 67.792 76.734 67.896 81.108 ; 
        RECT 67.36 76.734 67.464 81.108 ; 
        RECT 66.928 76.734 67.032 81.108 ; 
        RECT 66.496 76.734 66.6 81.108 ; 
        RECT 66.064 76.734 66.168 81.108 ; 
        RECT 65.632 76.734 65.736 81.108 ; 
        RECT 65.2 76.734 65.304 81.108 ; 
        RECT 64.348 76.734 64.656 81.108 ; 
        RECT 56.776 76.734 57.084 81.108 ; 
        RECT 56.128 76.734 56.232 81.108 ; 
        RECT 55.696 76.734 55.8 81.108 ; 
        RECT 55.264 76.734 55.368 81.108 ; 
        RECT 54.832 76.734 54.936 81.108 ; 
        RECT 54.4 76.734 54.504 81.108 ; 
        RECT 53.968 76.734 54.072 81.108 ; 
        RECT 53.536 76.734 53.64 81.108 ; 
        RECT 53.104 76.734 53.208 81.108 ; 
        RECT 52.672 76.734 52.776 81.108 ; 
        RECT 52.24 76.734 52.344 81.108 ; 
        RECT 51.808 76.734 51.912 81.108 ; 
        RECT 51.376 76.734 51.48 81.108 ; 
        RECT 50.944 76.734 51.048 81.108 ; 
        RECT 50.512 76.734 50.616 81.108 ; 
        RECT 50.08 76.734 50.184 81.108 ; 
        RECT 49.648 76.734 49.752 81.108 ; 
        RECT 49.216 76.734 49.32 81.108 ; 
        RECT 48.784 76.734 48.888 81.108 ; 
        RECT 48.352 76.734 48.456 81.108 ; 
        RECT 47.92 76.734 48.024 81.108 ; 
        RECT 47.488 76.734 47.592 81.108 ; 
        RECT 47.056 76.734 47.16 81.108 ; 
        RECT 46.624 76.734 46.728 81.108 ; 
        RECT 46.192 76.734 46.296 81.108 ; 
        RECT 45.76 76.734 45.864 81.108 ; 
        RECT 45.328 76.734 45.432 81.108 ; 
        RECT 44.896 76.734 45 81.108 ; 
        RECT 44.464 76.734 44.568 81.108 ; 
        RECT 44.032 76.734 44.136 81.108 ; 
        RECT 43.6 76.734 43.704 81.108 ; 
        RECT 43.168 76.734 43.272 81.108 ; 
        RECT 42.736 76.734 42.84 81.108 ; 
        RECT 42.304 76.734 42.408 81.108 ; 
        RECT 41.872 76.734 41.976 81.108 ; 
        RECT 41.44 76.734 41.544 81.108 ; 
        RECT 41.008 76.734 41.112 81.108 ; 
        RECT 40.576 76.734 40.68 81.108 ; 
        RECT 40.144 76.734 40.248 81.108 ; 
        RECT 39.712 76.734 39.816 81.108 ; 
        RECT 39.28 76.734 39.384 81.108 ; 
        RECT 38.848 76.734 38.952 81.108 ; 
        RECT 38.416 76.734 38.52 81.108 ; 
        RECT 37.984 76.734 38.088 81.108 ; 
        RECT 37.552 76.734 37.656 81.108 ; 
        RECT 37.12 76.734 37.224 81.108 ; 
        RECT 36.688 76.734 36.792 81.108 ; 
        RECT 36.256 76.734 36.36 81.108 ; 
        RECT 35.824 76.734 35.928 81.108 ; 
        RECT 35.392 76.734 35.496 81.108 ; 
        RECT 34.96 76.734 35.064 81.108 ; 
        RECT 34.528 76.734 34.632 81.108 ; 
        RECT 34.096 76.734 34.2 81.108 ; 
        RECT 33.664 76.734 33.768 81.108 ; 
        RECT 33.232 76.734 33.336 81.108 ; 
        RECT 32.8 76.734 32.904 81.108 ; 
        RECT 32.368 76.734 32.472 81.108 ; 
        RECT 31.936 76.734 32.04 81.108 ; 
        RECT 31.504 76.734 31.608 81.108 ; 
        RECT 31.072 76.734 31.176 81.108 ; 
        RECT 30.64 76.734 30.744 81.108 ; 
        RECT 30.208 76.734 30.312 81.108 ; 
        RECT 29.776 76.734 29.88 81.108 ; 
        RECT 29.344 76.734 29.448 81.108 ; 
        RECT 28.912 76.734 29.016 81.108 ; 
        RECT 28.48 76.734 28.584 81.108 ; 
        RECT 28.048 76.734 28.152 81.108 ; 
        RECT 27.616 76.734 27.72 81.108 ; 
        RECT 27.184 76.734 27.288 81.108 ; 
        RECT 26.752 76.734 26.856 81.108 ; 
        RECT 26.32 76.734 26.424 81.108 ; 
        RECT 25.888 76.734 25.992 81.108 ; 
        RECT 25.456 76.734 25.56 81.108 ; 
        RECT 25.024 76.734 25.128 81.108 ; 
        RECT 24.592 76.734 24.696 81.108 ; 
        RECT 24.16 76.734 24.264 81.108 ; 
        RECT 23.728 76.734 23.832 81.108 ; 
        RECT 23.296 76.734 23.4 81.108 ; 
        RECT 22.864 76.734 22.968 81.108 ; 
        RECT 22.432 76.734 22.536 81.108 ; 
        RECT 22 76.734 22.104 81.108 ; 
        RECT 21.568 76.734 21.672 81.108 ; 
        RECT 21.136 76.734 21.24 81.108 ; 
        RECT 20.704 76.734 20.808 81.108 ; 
        RECT 20.272 76.734 20.376 81.108 ; 
        RECT 19.84 76.734 19.944 81.108 ; 
        RECT 19.408 76.734 19.512 81.108 ; 
        RECT 18.976 76.734 19.08 81.108 ; 
        RECT 18.544 76.734 18.648 81.108 ; 
        RECT 18.112 76.734 18.216 81.108 ; 
        RECT 17.68 76.734 17.784 81.108 ; 
        RECT 17.248 76.734 17.352 81.108 ; 
        RECT 16.816 76.734 16.92 81.108 ; 
        RECT 16.384 76.734 16.488 81.108 ; 
        RECT 15.952 76.734 16.056 81.108 ; 
        RECT 15.52 76.734 15.624 81.108 ; 
        RECT 15.088 76.734 15.192 81.108 ; 
        RECT 14.656 76.734 14.76 81.108 ; 
        RECT 14.224 76.734 14.328 81.108 ; 
        RECT 13.792 76.734 13.896 81.108 ; 
        RECT 13.36 76.734 13.464 81.108 ; 
        RECT 12.928 76.734 13.032 81.108 ; 
        RECT 12.496 76.734 12.6 81.108 ; 
        RECT 12.064 76.734 12.168 81.108 ; 
        RECT 11.632 76.734 11.736 81.108 ; 
        RECT 11.2 76.734 11.304 81.108 ; 
        RECT 10.768 76.734 10.872 81.108 ; 
        RECT 10.336 76.734 10.44 81.108 ; 
        RECT 9.904 76.734 10.008 81.108 ; 
        RECT 9.472 76.734 9.576 81.108 ; 
        RECT 9.04 76.734 9.144 81.108 ; 
        RECT 8.608 76.734 8.712 81.108 ; 
        RECT 8.176 76.734 8.28 81.108 ; 
        RECT 7.744 76.734 7.848 81.108 ; 
        RECT 7.312 76.734 7.416 81.108 ; 
        RECT 6.88 76.734 6.984 81.108 ; 
        RECT 6.448 76.734 6.552 81.108 ; 
        RECT 6.016 76.734 6.12 81.108 ; 
        RECT 5.584 76.734 5.688 81.108 ; 
        RECT 5.152 76.734 5.256 81.108 ; 
        RECT 4.72 76.734 4.824 81.108 ; 
        RECT 4.288 76.734 4.392 81.108 ; 
        RECT 3.856 76.734 3.96 81.108 ; 
        RECT 3.424 76.734 3.528 81.108 ; 
        RECT 2.992 76.734 3.096 81.108 ; 
        RECT 2.56 76.734 2.664 81.108 ; 
        RECT 2.128 76.734 2.232 81.108 ; 
        RECT 1.696 76.734 1.8 81.108 ; 
        RECT 1.264 76.734 1.368 81.108 ; 
        RECT 0.832 76.734 0.936 81.108 ; 
        RECT 0.02 76.734 0.36 81.108 ; 
        RECT 62.212 81.054 62.724 85.428 ; 
        RECT 62.156 83.716 62.724 85.006 ; 
        RECT 61.276 82.624 61.812 85.428 ; 
        RECT 61.184 83.964 61.812 84.996 ; 
        RECT 61.276 81.054 61.668 85.428 ; 
        RECT 61.276 81.538 61.724 82.496 ; 
        RECT 61.276 81.054 61.812 81.41 ; 
        RECT 60.376 82.856 60.912 85.428 ; 
        RECT 60.376 81.054 60.768 85.428 ; 
        RECT 58.708 81.054 59.04 85.428 ; 
        RECT 58.708 81.408 59.096 85.15 ; 
        RECT 121.072 81.054 121.412 85.428 ; 
        RECT 120.496 81.054 120.6 85.428 ; 
        RECT 120.064 81.054 120.168 85.428 ; 
        RECT 119.632 81.054 119.736 85.428 ; 
        RECT 119.2 81.054 119.304 85.428 ; 
        RECT 118.768 81.054 118.872 85.428 ; 
        RECT 118.336 81.054 118.44 85.428 ; 
        RECT 117.904 81.054 118.008 85.428 ; 
        RECT 117.472 81.054 117.576 85.428 ; 
        RECT 117.04 81.054 117.144 85.428 ; 
        RECT 116.608 81.054 116.712 85.428 ; 
        RECT 116.176 81.054 116.28 85.428 ; 
        RECT 115.744 81.054 115.848 85.428 ; 
        RECT 115.312 81.054 115.416 85.428 ; 
        RECT 114.88 81.054 114.984 85.428 ; 
        RECT 114.448 81.054 114.552 85.428 ; 
        RECT 114.016 81.054 114.12 85.428 ; 
        RECT 113.584 81.054 113.688 85.428 ; 
        RECT 113.152 81.054 113.256 85.428 ; 
        RECT 112.72 81.054 112.824 85.428 ; 
        RECT 112.288 81.054 112.392 85.428 ; 
        RECT 111.856 81.054 111.96 85.428 ; 
        RECT 111.424 81.054 111.528 85.428 ; 
        RECT 110.992 81.054 111.096 85.428 ; 
        RECT 110.56 81.054 110.664 85.428 ; 
        RECT 110.128 81.054 110.232 85.428 ; 
        RECT 109.696 81.054 109.8 85.428 ; 
        RECT 109.264 81.054 109.368 85.428 ; 
        RECT 108.832 81.054 108.936 85.428 ; 
        RECT 108.4 81.054 108.504 85.428 ; 
        RECT 107.968 81.054 108.072 85.428 ; 
        RECT 107.536 81.054 107.64 85.428 ; 
        RECT 107.104 81.054 107.208 85.428 ; 
        RECT 106.672 81.054 106.776 85.428 ; 
        RECT 106.24 81.054 106.344 85.428 ; 
        RECT 105.808 81.054 105.912 85.428 ; 
        RECT 105.376 81.054 105.48 85.428 ; 
        RECT 104.944 81.054 105.048 85.428 ; 
        RECT 104.512 81.054 104.616 85.428 ; 
        RECT 104.08 81.054 104.184 85.428 ; 
        RECT 103.648 81.054 103.752 85.428 ; 
        RECT 103.216 81.054 103.32 85.428 ; 
        RECT 102.784 81.054 102.888 85.428 ; 
        RECT 102.352 81.054 102.456 85.428 ; 
        RECT 101.92 81.054 102.024 85.428 ; 
        RECT 101.488 81.054 101.592 85.428 ; 
        RECT 101.056 81.054 101.16 85.428 ; 
        RECT 100.624 81.054 100.728 85.428 ; 
        RECT 100.192 81.054 100.296 85.428 ; 
        RECT 99.76 81.054 99.864 85.428 ; 
        RECT 99.328 81.054 99.432 85.428 ; 
        RECT 98.896 81.054 99 85.428 ; 
        RECT 98.464 81.054 98.568 85.428 ; 
        RECT 98.032 81.054 98.136 85.428 ; 
        RECT 97.6 81.054 97.704 85.428 ; 
        RECT 97.168 81.054 97.272 85.428 ; 
        RECT 96.736 81.054 96.84 85.428 ; 
        RECT 96.304 81.054 96.408 85.428 ; 
        RECT 95.872 81.054 95.976 85.428 ; 
        RECT 95.44 81.054 95.544 85.428 ; 
        RECT 95.008 81.054 95.112 85.428 ; 
        RECT 94.576 81.054 94.68 85.428 ; 
        RECT 94.144 81.054 94.248 85.428 ; 
        RECT 93.712 81.054 93.816 85.428 ; 
        RECT 93.28 81.054 93.384 85.428 ; 
        RECT 92.848 81.054 92.952 85.428 ; 
        RECT 92.416 81.054 92.52 85.428 ; 
        RECT 91.984 81.054 92.088 85.428 ; 
        RECT 91.552 81.054 91.656 85.428 ; 
        RECT 91.12 81.054 91.224 85.428 ; 
        RECT 90.688 81.054 90.792 85.428 ; 
        RECT 90.256 81.054 90.36 85.428 ; 
        RECT 89.824 81.054 89.928 85.428 ; 
        RECT 89.392 81.054 89.496 85.428 ; 
        RECT 88.96 81.054 89.064 85.428 ; 
        RECT 88.528 81.054 88.632 85.428 ; 
        RECT 88.096 81.054 88.2 85.428 ; 
        RECT 87.664 81.054 87.768 85.428 ; 
        RECT 87.232 81.054 87.336 85.428 ; 
        RECT 86.8 81.054 86.904 85.428 ; 
        RECT 86.368 81.054 86.472 85.428 ; 
        RECT 85.936 81.054 86.04 85.428 ; 
        RECT 85.504 81.054 85.608 85.428 ; 
        RECT 85.072 81.054 85.176 85.428 ; 
        RECT 84.64 81.054 84.744 85.428 ; 
        RECT 84.208 81.054 84.312 85.428 ; 
        RECT 83.776 81.054 83.88 85.428 ; 
        RECT 83.344 81.054 83.448 85.428 ; 
        RECT 82.912 81.054 83.016 85.428 ; 
        RECT 82.48 81.054 82.584 85.428 ; 
        RECT 82.048 81.054 82.152 85.428 ; 
        RECT 81.616 81.054 81.72 85.428 ; 
        RECT 81.184 81.054 81.288 85.428 ; 
        RECT 80.752 81.054 80.856 85.428 ; 
        RECT 80.32 81.054 80.424 85.428 ; 
        RECT 79.888 81.054 79.992 85.428 ; 
        RECT 79.456 81.054 79.56 85.428 ; 
        RECT 79.024 81.054 79.128 85.428 ; 
        RECT 78.592 81.054 78.696 85.428 ; 
        RECT 78.16 81.054 78.264 85.428 ; 
        RECT 77.728 81.054 77.832 85.428 ; 
        RECT 77.296 81.054 77.4 85.428 ; 
        RECT 76.864 81.054 76.968 85.428 ; 
        RECT 76.432 81.054 76.536 85.428 ; 
        RECT 76 81.054 76.104 85.428 ; 
        RECT 75.568 81.054 75.672 85.428 ; 
        RECT 75.136 81.054 75.24 85.428 ; 
        RECT 74.704 81.054 74.808 85.428 ; 
        RECT 74.272 81.054 74.376 85.428 ; 
        RECT 73.84 81.054 73.944 85.428 ; 
        RECT 73.408 81.054 73.512 85.428 ; 
        RECT 72.976 81.054 73.08 85.428 ; 
        RECT 72.544 81.054 72.648 85.428 ; 
        RECT 72.112 81.054 72.216 85.428 ; 
        RECT 71.68 81.054 71.784 85.428 ; 
        RECT 71.248 81.054 71.352 85.428 ; 
        RECT 70.816 81.054 70.92 85.428 ; 
        RECT 70.384 81.054 70.488 85.428 ; 
        RECT 69.952 81.054 70.056 85.428 ; 
        RECT 69.52 81.054 69.624 85.428 ; 
        RECT 69.088 81.054 69.192 85.428 ; 
        RECT 68.656 81.054 68.76 85.428 ; 
        RECT 68.224 81.054 68.328 85.428 ; 
        RECT 67.792 81.054 67.896 85.428 ; 
        RECT 67.36 81.054 67.464 85.428 ; 
        RECT 66.928 81.054 67.032 85.428 ; 
        RECT 66.496 81.054 66.6 85.428 ; 
        RECT 66.064 81.054 66.168 85.428 ; 
        RECT 65.632 81.054 65.736 85.428 ; 
        RECT 65.2 81.054 65.304 85.428 ; 
        RECT 64.348 81.054 64.656 85.428 ; 
        RECT 56.776 81.054 57.084 85.428 ; 
        RECT 56.128 81.054 56.232 85.428 ; 
        RECT 55.696 81.054 55.8 85.428 ; 
        RECT 55.264 81.054 55.368 85.428 ; 
        RECT 54.832 81.054 54.936 85.428 ; 
        RECT 54.4 81.054 54.504 85.428 ; 
        RECT 53.968 81.054 54.072 85.428 ; 
        RECT 53.536 81.054 53.64 85.428 ; 
        RECT 53.104 81.054 53.208 85.428 ; 
        RECT 52.672 81.054 52.776 85.428 ; 
        RECT 52.24 81.054 52.344 85.428 ; 
        RECT 51.808 81.054 51.912 85.428 ; 
        RECT 51.376 81.054 51.48 85.428 ; 
        RECT 50.944 81.054 51.048 85.428 ; 
        RECT 50.512 81.054 50.616 85.428 ; 
        RECT 50.08 81.054 50.184 85.428 ; 
        RECT 49.648 81.054 49.752 85.428 ; 
        RECT 49.216 81.054 49.32 85.428 ; 
        RECT 48.784 81.054 48.888 85.428 ; 
        RECT 48.352 81.054 48.456 85.428 ; 
        RECT 47.92 81.054 48.024 85.428 ; 
        RECT 47.488 81.054 47.592 85.428 ; 
        RECT 47.056 81.054 47.16 85.428 ; 
        RECT 46.624 81.054 46.728 85.428 ; 
        RECT 46.192 81.054 46.296 85.428 ; 
        RECT 45.76 81.054 45.864 85.428 ; 
        RECT 45.328 81.054 45.432 85.428 ; 
        RECT 44.896 81.054 45 85.428 ; 
        RECT 44.464 81.054 44.568 85.428 ; 
        RECT 44.032 81.054 44.136 85.428 ; 
        RECT 43.6 81.054 43.704 85.428 ; 
        RECT 43.168 81.054 43.272 85.428 ; 
        RECT 42.736 81.054 42.84 85.428 ; 
        RECT 42.304 81.054 42.408 85.428 ; 
        RECT 41.872 81.054 41.976 85.428 ; 
        RECT 41.44 81.054 41.544 85.428 ; 
        RECT 41.008 81.054 41.112 85.428 ; 
        RECT 40.576 81.054 40.68 85.428 ; 
        RECT 40.144 81.054 40.248 85.428 ; 
        RECT 39.712 81.054 39.816 85.428 ; 
        RECT 39.28 81.054 39.384 85.428 ; 
        RECT 38.848 81.054 38.952 85.428 ; 
        RECT 38.416 81.054 38.52 85.428 ; 
        RECT 37.984 81.054 38.088 85.428 ; 
        RECT 37.552 81.054 37.656 85.428 ; 
        RECT 37.12 81.054 37.224 85.428 ; 
        RECT 36.688 81.054 36.792 85.428 ; 
        RECT 36.256 81.054 36.36 85.428 ; 
        RECT 35.824 81.054 35.928 85.428 ; 
        RECT 35.392 81.054 35.496 85.428 ; 
        RECT 34.96 81.054 35.064 85.428 ; 
        RECT 34.528 81.054 34.632 85.428 ; 
        RECT 34.096 81.054 34.2 85.428 ; 
        RECT 33.664 81.054 33.768 85.428 ; 
        RECT 33.232 81.054 33.336 85.428 ; 
        RECT 32.8 81.054 32.904 85.428 ; 
        RECT 32.368 81.054 32.472 85.428 ; 
        RECT 31.936 81.054 32.04 85.428 ; 
        RECT 31.504 81.054 31.608 85.428 ; 
        RECT 31.072 81.054 31.176 85.428 ; 
        RECT 30.64 81.054 30.744 85.428 ; 
        RECT 30.208 81.054 30.312 85.428 ; 
        RECT 29.776 81.054 29.88 85.428 ; 
        RECT 29.344 81.054 29.448 85.428 ; 
        RECT 28.912 81.054 29.016 85.428 ; 
        RECT 28.48 81.054 28.584 85.428 ; 
        RECT 28.048 81.054 28.152 85.428 ; 
        RECT 27.616 81.054 27.72 85.428 ; 
        RECT 27.184 81.054 27.288 85.428 ; 
        RECT 26.752 81.054 26.856 85.428 ; 
        RECT 26.32 81.054 26.424 85.428 ; 
        RECT 25.888 81.054 25.992 85.428 ; 
        RECT 25.456 81.054 25.56 85.428 ; 
        RECT 25.024 81.054 25.128 85.428 ; 
        RECT 24.592 81.054 24.696 85.428 ; 
        RECT 24.16 81.054 24.264 85.428 ; 
        RECT 23.728 81.054 23.832 85.428 ; 
        RECT 23.296 81.054 23.4 85.428 ; 
        RECT 22.864 81.054 22.968 85.428 ; 
        RECT 22.432 81.054 22.536 85.428 ; 
        RECT 22 81.054 22.104 85.428 ; 
        RECT 21.568 81.054 21.672 85.428 ; 
        RECT 21.136 81.054 21.24 85.428 ; 
        RECT 20.704 81.054 20.808 85.428 ; 
        RECT 20.272 81.054 20.376 85.428 ; 
        RECT 19.84 81.054 19.944 85.428 ; 
        RECT 19.408 81.054 19.512 85.428 ; 
        RECT 18.976 81.054 19.08 85.428 ; 
        RECT 18.544 81.054 18.648 85.428 ; 
        RECT 18.112 81.054 18.216 85.428 ; 
        RECT 17.68 81.054 17.784 85.428 ; 
        RECT 17.248 81.054 17.352 85.428 ; 
        RECT 16.816 81.054 16.92 85.428 ; 
        RECT 16.384 81.054 16.488 85.428 ; 
        RECT 15.952 81.054 16.056 85.428 ; 
        RECT 15.52 81.054 15.624 85.428 ; 
        RECT 15.088 81.054 15.192 85.428 ; 
        RECT 14.656 81.054 14.76 85.428 ; 
        RECT 14.224 81.054 14.328 85.428 ; 
        RECT 13.792 81.054 13.896 85.428 ; 
        RECT 13.36 81.054 13.464 85.428 ; 
        RECT 12.928 81.054 13.032 85.428 ; 
        RECT 12.496 81.054 12.6 85.428 ; 
        RECT 12.064 81.054 12.168 85.428 ; 
        RECT 11.632 81.054 11.736 85.428 ; 
        RECT 11.2 81.054 11.304 85.428 ; 
        RECT 10.768 81.054 10.872 85.428 ; 
        RECT 10.336 81.054 10.44 85.428 ; 
        RECT 9.904 81.054 10.008 85.428 ; 
        RECT 9.472 81.054 9.576 85.428 ; 
        RECT 9.04 81.054 9.144 85.428 ; 
        RECT 8.608 81.054 8.712 85.428 ; 
        RECT 8.176 81.054 8.28 85.428 ; 
        RECT 7.744 81.054 7.848 85.428 ; 
        RECT 7.312 81.054 7.416 85.428 ; 
        RECT 6.88 81.054 6.984 85.428 ; 
        RECT 6.448 81.054 6.552 85.428 ; 
        RECT 6.016 81.054 6.12 85.428 ; 
        RECT 5.584 81.054 5.688 85.428 ; 
        RECT 5.152 81.054 5.256 85.428 ; 
        RECT 4.72 81.054 4.824 85.428 ; 
        RECT 4.288 81.054 4.392 85.428 ; 
        RECT 3.856 81.054 3.96 85.428 ; 
        RECT 3.424 81.054 3.528 85.428 ; 
        RECT 2.992 81.054 3.096 85.428 ; 
        RECT 2.56 81.054 2.664 85.428 ; 
        RECT 2.128 81.054 2.232 85.428 ; 
        RECT 1.696 81.054 1.8 85.428 ; 
        RECT 1.264 81.054 1.368 85.428 ; 
        RECT 0.832 81.054 0.936 85.428 ; 
        RECT 0.02 81.054 0.36 85.428 ; 
        RECT 62.212 85.374 62.724 89.748 ; 
        RECT 62.156 88.036 62.724 89.326 ; 
        RECT 61.276 86.944 61.812 89.748 ; 
        RECT 61.184 88.284 61.812 89.316 ; 
        RECT 61.276 85.374 61.668 89.748 ; 
        RECT 61.276 85.858 61.724 86.816 ; 
        RECT 61.276 85.374 61.812 85.73 ; 
        RECT 60.376 87.176 60.912 89.748 ; 
        RECT 60.376 85.374 60.768 89.748 ; 
        RECT 58.708 85.374 59.04 89.748 ; 
        RECT 58.708 85.728 59.096 89.47 ; 
        RECT 121.072 85.374 121.412 89.748 ; 
        RECT 120.496 85.374 120.6 89.748 ; 
        RECT 120.064 85.374 120.168 89.748 ; 
        RECT 119.632 85.374 119.736 89.748 ; 
        RECT 119.2 85.374 119.304 89.748 ; 
        RECT 118.768 85.374 118.872 89.748 ; 
        RECT 118.336 85.374 118.44 89.748 ; 
        RECT 117.904 85.374 118.008 89.748 ; 
        RECT 117.472 85.374 117.576 89.748 ; 
        RECT 117.04 85.374 117.144 89.748 ; 
        RECT 116.608 85.374 116.712 89.748 ; 
        RECT 116.176 85.374 116.28 89.748 ; 
        RECT 115.744 85.374 115.848 89.748 ; 
        RECT 115.312 85.374 115.416 89.748 ; 
        RECT 114.88 85.374 114.984 89.748 ; 
        RECT 114.448 85.374 114.552 89.748 ; 
        RECT 114.016 85.374 114.12 89.748 ; 
        RECT 113.584 85.374 113.688 89.748 ; 
        RECT 113.152 85.374 113.256 89.748 ; 
        RECT 112.72 85.374 112.824 89.748 ; 
        RECT 112.288 85.374 112.392 89.748 ; 
        RECT 111.856 85.374 111.96 89.748 ; 
        RECT 111.424 85.374 111.528 89.748 ; 
        RECT 110.992 85.374 111.096 89.748 ; 
        RECT 110.56 85.374 110.664 89.748 ; 
        RECT 110.128 85.374 110.232 89.748 ; 
        RECT 109.696 85.374 109.8 89.748 ; 
        RECT 109.264 85.374 109.368 89.748 ; 
        RECT 108.832 85.374 108.936 89.748 ; 
        RECT 108.4 85.374 108.504 89.748 ; 
        RECT 107.968 85.374 108.072 89.748 ; 
        RECT 107.536 85.374 107.64 89.748 ; 
        RECT 107.104 85.374 107.208 89.748 ; 
        RECT 106.672 85.374 106.776 89.748 ; 
        RECT 106.24 85.374 106.344 89.748 ; 
        RECT 105.808 85.374 105.912 89.748 ; 
        RECT 105.376 85.374 105.48 89.748 ; 
        RECT 104.944 85.374 105.048 89.748 ; 
        RECT 104.512 85.374 104.616 89.748 ; 
        RECT 104.08 85.374 104.184 89.748 ; 
        RECT 103.648 85.374 103.752 89.748 ; 
        RECT 103.216 85.374 103.32 89.748 ; 
        RECT 102.784 85.374 102.888 89.748 ; 
        RECT 102.352 85.374 102.456 89.748 ; 
        RECT 101.92 85.374 102.024 89.748 ; 
        RECT 101.488 85.374 101.592 89.748 ; 
        RECT 101.056 85.374 101.16 89.748 ; 
        RECT 100.624 85.374 100.728 89.748 ; 
        RECT 100.192 85.374 100.296 89.748 ; 
        RECT 99.76 85.374 99.864 89.748 ; 
        RECT 99.328 85.374 99.432 89.748 ; 
        RECT 98.896 85.374 99 89.748 ; 
        RECT 98.464 85.374 98.568 89.748 ; 
        RECT 98.032 85.374 98.136 89.748 ; 
        RECT 97.6 85.374 97.704 89.748 ; 
        RECT 97.168 85.374 97.272 89.748 ; 
        RECT 96.736 85.374 96.84 89.748 ; 
        RECT 96.304 85.374 96.408 89.748 ; 
        RECT 95.872 85.374 95.976 89.748 ; 
        RECT 95.44 85.374 95.544 89.748 ; 
        RECT 95.008 85.374 95.112 89.748 ; 
        RECT 94.576 85.374 94.68 89.748 ; 
        RECT 94.144 85.374 94.248 89.748 ; 
        RECT 93.712 85.374 93.816 89.748 ; 
        RECT 93.28 85.374 93.384 89.748 ; 
        RECT 92.848 85.374 92.952 89.748 ; 
        RECT 92.416 85.374 92.52 89.748 ; 
        RECT 91.984 85.374 92.088 89.748 ; 
        RECT 91.552 85.374 91.656 89.748 ; 
        RECT 91.12 85.374 91.224 89.748 ; 
        RECT 90.688 85.374 90.792 89.748 ; 
        RECT 90.256 85.374 90.36 89.748 ; 
        RECT 89.824 85.374 89.928 89.748 ; 
        RECT 89.392 85.374 89.496 89.748 ; 
        RECT 88.96 85.374 89.064 89.748 ; 
        RECT 88.528 85.374 88.632 89.748 ; 
        RECT 88.096 85.374 88.2 89.748 ; 
        RECT 87.664 85.374 87.768 89.748 ; 
        RECT 87.232 85.374 87.336 89.748 ; 
        RECT 86.8 85.374 86.904 89.748 ; 
        RECT 86.368 85.374 86.472 89.748 ; 
        RECT 85.936 85.374 86.04 89.748 ; 
        RECT 85.504 85.374 85.608 89.748 ; 
        RECT 85.072 85.374 85.176 89.748 ; 
        RECT 84.64 85.374 84.744 89.748 ; 
        RECT 84.208 85.374 84.312 89.748 ; 
        RECT 83.776 85.374 83.88 89.748 ; 
        RECT 83.344 85.374 83.448 89.748 ; 
        RECT 82.912 85.374 83.016 89.748 ; 
        RECT 82.48 85.374 82.584 89.748 ; 
        RECT 82.048 85.374 82.152 89.748 ; 
        RECT 81.616 85.374 81.72 89.748 ; 
        RECT 81.184 85.374 81.288 89.748 ; 
        RECT 80.752 85.374 80.856 89.748 ; 
        RECT 80.32 85.374 80.424 89.748 ; 
        RECT 79.888 85.374 79.992 89.748 ; 
        RECT 79.456 85.374 79.56 89.748 ; 
        RECT 79.024 85.374 79.128 89.748 ; 
        RECT 78.592 85.374 78.696 89.748 ; 
        RECT 78.16 85.374 78.264 89.748 ; 
        RECT 77.728 85.374 77.832 89.748 ; 
        RECT 77.296 85.374 77.4 89.748 ; 
        RECT 76.864 85.374 76.968 89.748 ; 
        RECT 76.432 85.374 76.536 89.748 ; 
        RECT 76 85.374 76.104 89.748 ; 
        RECT 75.568 85.374 75.672 89.748 ; 
        RECT 75.136 85.374 75.24 89.748 ; 
        RECT 74.704 85.374 74.808 89.748 ; 
        RECT 74.272 85.374 74.376 89.748 ; 
        RECT 73.84 85.374 73.944 89.748 ; 
        RECT 73.408 85.374 73.512 89.748 ; 
        RECT 72.976 85.374 73.08 89.748 ; 
        RECT 72.544 85.374 72.648 89.748 ; 
        RECT 72.112 85.374 72.216 89.748 ; 
        RECT 71.68 85.374 71.784 89.748 ; 
        RECT 71.248 85.374 71.352 89.748 ; 
        RECT 70.816 85.374 70.92 89.748 ; 
        RECT 70.384 85.374 70.488 89.748 ; 
        RECT 69.952 85.374 70.056 89.748 ; 
        RECT 69.52 85.374 69.624 89.748 ; 
        RECT 69.088 85.374 69.192 89.748 ; 
        RECT 68.656 85.374 68.76 89.748 ; 
        RECT 68.224 85.374 68.328 89.748 ; 
        RECT 67.792 85.374 67.896 89.748 ; 
        RECT 67.36 85.374 67.464 89.748 ; 
        RECT 66.928 85.374 67.032 89.748 ; 
        RECT 66.496 85.374 66.6 89.748 ; 
        RECT 66.064 85.374 66.168 89.748 ; 
        RECT 65.632 85.374 65.736 89.748 ; 
        RECT 65.2 85.374 65.304 89.748 ; 
        RECT 64.348 85.374 64.656 89.748 ; 
        RECT 56.776 85.374 57.084 89.748 ; 
        RECT 56.128 85.374 56.232 89.748 ; 
        RECT 55.696 85.374 55.8 89.748 ; 
        RECT 55.264 85.374 55.368 89.748 ; 
        RECT 54.832 85.374 54.936 89.748 ; 
        RECT 54.4 85.374 54.504 89.748 ; 
        RECT 53.968 85.374 54.072 89.748 ; 
        RECT 53.536 85.374 53.64 89.748 ; 
        RECT 53.104 85.374 53.208 89.748 ; 
        RECT 52.672 85.374 52.776 89.748 ; 
        RECT 52.24 85.374 52.344 89.748 ; 
        RECT 51.808 85.374 51.912 89.748 ; 
        RECT 51.376 85.374 51.48 89.748 ; 
        RECT 50.944 85.374 51.048 89.748 ; 
        RECT 50.512 85.374 50.616 89.748 ; 
        RECT 50.08 85.374 50.184 89.748 ; 
        RECT 49.648 85.374 49.752 89.748 ; 
        RECT 49.216 85.374 49.32 89.748 ; 
        RECT 48.784 85.374 48.888 89.748 ; 
        RECT 48.352 85.374 48.456 89.748 ; 
        RECT 47.92 85.374 48.024 89.748 ; 
        RECT 47.488 85.374 47.592 89.748 ; 
        RECT 47.056 85.374 47.16 89.748 ; 
        RECT 46.624 85.374 46.728 89.748 ; 
        RECT 46.192 85.374 46.296 89.748 ; 
        RECT 45.76 85.374 45.864 89.748 ; 
        RECT 45.328 85.374 45.432 89.748 ; 
        RECT 44.896 85.374 45 89.748 ; 
        RECT 44.464 85.374 44.568 89.748 ; 
        RECT 44.032 85.374 44.136 89.748 ; 
        RECT 43.6 85.374 43.704 89.748 ; 
        RECT 43.168 85.374 43.272 89.748 ; 
        RECT 42.736 85.374 42.84 89.748 ; 
        RECT 42.304 85.374 42.408 89.748 ; 
        RECT 41.872 85.374 41.976 89.748 ; 
        RECT 41.44 85.374 41.544 89.748 ; 
        RECT 41.008 85.374 41.112 89.748 ; 
        RECT 40.576 85.374 40.68 89.748 ; 
        RECT 40.144 85.374 40.248 89.748 ; 
        RECT 39.712 85.374 39.816 89.748 ; 
        RECT 39.28 85.374 39.384 89.748 ; 
        RECT 38.848 85.374 38.952 89.748 ; 
        RECT 38.416 85.374 38.52 89.748 ; 
        RECT 37.984 85.374 38.088 89.748 ; 
        RECT 37.552 85.374 37.656 89.748 ; 
        RECT 37.12 85.374 37.224 89.748 ; 
        RECT 36.688 85.374 36.792 89.748 ; 
        RECT 36.256 85.374 36.36 89.748 ; 
        RECT 35.824 85.374 35.928 89.748 ; 
        RECT 35.392 85.374 35.496 89.748 ; 
        RECT 34.96 85.374 35.064 89.748 ; 
        RECT 34.528 85.374 34.632 89.748 ; 
        RECT 34.096 85.374 34.2 89.748 ; 
        RECT 33.664 85.374 33.768 89.748 ; 
        RECT 33.232 85.374 33.336 89.748 ; 
        RECT 32.8 85.374 32.904 89.748 ; 
        RECT 32.368 85.374 32.472 89.748 ; 
        RECT 31.936 85.374 32.04 89.748 ; 
        RECT 31.504 85.374 31.608 89.748 ; 
        RECT 31.072 85.374 31.176 89.748 ; 
        RECT 30.64 85.374 30.744 89.748 ; 
        RECT 30.208 85.374 30.312 89.748 ; 
        RECT 29.776 85.374 29.88 89.748 ; 
        RECT 29.344 85.374 29.448 89.748 ; 
        RECT 28.912 85.374 29.016 89.748 ; 
        RECT 28.48 85.374 28.584 89.748 ; 
        RECT 28.048 85.374 28.152 89.748 ; 
        RECT 27.616 85.374 27.72 89.748 ; 
        RECT 27.184 85.374 27.288 89.748 ; 
        RECT 26.752 85.374 26.856 89.748 ; 
        RECT 26.32 85.374 26.424 89.748 ; 
        RECT 25.888 85.374 25.992 89.748 ; 
        RECT 25.456 85.374 25.56 89.748 ; 
        RECT 25.024 85.374 25.128 89.748 ; 
        RECT 24.592 85.374 24.696 89.748 ; 
        RECT 24.16 85.374 24.264 89.748 ; 
        RECT 23.728 85.374 23.832 89.748 ; 
        RECT 23.296 85.374 23.4 89.748 ; 
        RECT 22.864 85.374 22.968 89.748 ; 
        RECT 22.432 85.374 22.536 89.748 ; 
        RECT 22 85.374 22.104 89.748 ; 
        RECT 21.568 85.374 21.672 89.748 ; 
        RECT 21.136 85.374 21.24 89.748 ; 
        RECT 20.704 85.374 20.808 89.748 ; 
        RECT 20.272 85.374 20.376 89.748 ; 
        RECT 19.84 85.374 19.944 89.748 ; 
        RECT 19.408 85.374 19.512 89.748 ; 
        RECT 18.976 85.374 19.08 89.748 ; 
        RECT 18.544 85.374 18.648 89.748 ; 
        RECT 18.112 85.374 18.216 89.748 ; 
        RECT 17.68 85.374 17.784 89.748 ; 
        RECT 17.248 85.374 17.352 89.748 ; 
        RECT 16.816 85.374 16.92 89.748 ; 
        RECT 16.384 85.374 16.488 89.748 ; 
        RECT 15.952 85.374 16.056 89.748 ; 
        RECT 15.52 85.374 15.624 89.748 ; 
        RECT 15.088 85.374 15.192 89.748 ; 
        RECT 14.656 85.374 14.76 89.748 ; 
        RECT 14.224 85.374 14.328 89.748 ; 
        RECT 13.792 85.374 13.896 89.748 ; 
        RECT 13.36 85.374 13.464 89.748 ; 
        RECT 12.928 85.374 13.032 89.748 ; 
        RECT 12.496 85.374 12.6 89.748 ; 
        RECT 12.064 85.374 12.168 89.748 ; 
        RECT 11.632 85.374 11.736 89.748 ; 
        RECT 11.2 85.374 11.304 89.748 ; 
        RECT 10.768 85.374 10.872 89.748 ; 
        RECT 10.336 85.374 10.44 89.748 ; 
        RECT 9.904 85.374 10.008 89.748 ; 
        RECT 9.472 85.374 9.576 89.748 ; 
        RECT 9.04 85.374 9.144 89.748 ; 
        RECT 8.608 85.374 8.712 89.748 ; 
        RECT 8.176 85.374 8.28 89.748 ; 
        RECT 7.744 85.374 7.848 89.748 ; 
        RECT 7.312 85.374 7.416 89.748 ; 
        RECT 6.88 85.374 6.984 89.748 ; 
        RECT 6.448 85.374 6.552 89.748 ; 
        RECT 6.016 85.374 6.12 89.748 ; 
        RECT 5.584 85.374 5.688 89.748 ; 
        RECT 5.152 85.374 5.256 89.748 ; 
        RECT 4.72 85.374 4.824 89.748 ; 
        RECT 4.288 85.374 4.392 89.748 ; 
        RECT 3.856 85.374 3.96 89.748 ; 
        RECT 3.424 85.374 3.528 89.748 ; 
        RECT 2.992 85.374 3.096 89.748 ; 
        RECT 2.56 85.374 2.664 89.748 ; 
        RECT 2.128 85.374 2.232 89.748 ; 
        RECT 1.696 85.374 1.8 89.748 ; 
        RECT 1.264 85.374 1.368 89.748 ; 
        RECT 0.832 85.374 0.936 89.748 ; 
        RECT 0.02 85.374 0.36 89.748 ; 
        RECT 62.212 89.694 62.724 94.068 ; 
        RECT 62.156 92.356 62.724 93.646 ; 
        RECT 61.276 91.264 61.812 94.068 ; 
        RECT 61.184 92.604 61.812 93.636 ; 
        RECT 61.276 89.694 61.668 94.068 ; 
        RECT 61.276 90.178 61.724 91.136 ; 
        RECT 61.276 89.694 61.812 90.05 ; 
        RECT 60.376 91.496 60.912 94.068 ; 
        RECT 60.376 89.694 60.768 94.068 ; 
        RECT 58.708 89.694 59.04 94.068 ; 
        RECT 58.708 90.048 59.096 93.79 ; 
        RECT 121.072 89.694 121.412 94.068 ; 
        RECT 120.496 89.694 120.6 94.068 ; 
        RECT 120.064 89.694 120.168 94.068 ; 
        RECT 119.632 89.694 119.736 94.068 ; 
        RECT 119.2 89.694 119.304 94.068 ; 
        RECT 118.768 89.694 118.872 94.068 ; 
        RECT 118.336 89.694 118.44 94.068 ; 
        RECT 117.904 89.694 118.008 94.068 ; 
        RECT 117.472 89.694 117.576 94.068 ; 
        RECT 117.04 89.694 117.144 94.068 ; 
        RECT 116.608 89.694 116.712 94.068 ; 
        RECT 116.176 89.694 116.28 94.068 ; 
        RECT 115.744 89.694 115.848 94.068 ; 
        RECT 115.312 89.694 115.416 94.068 ; 
        RECT 114.88 89.694 114.984 94.068 ; 
        RECT 114.448 89.694 114.552 94.068 ; 
        RECT 114.016 89.694 114.12 94.068 ; 
        RECT 113.584 89.694 113.688 94.068 ; 
        RECT 113.152 89.694 113.256 94.068 ; 
        RECT 112.72 89.694 112.824 94.068 ; 
        RECT 112.288 89.694 112.392 94.068 ; 
        RECT 111.856 89.694 111.96 94.068 ; 
        RECT 111.424 89.694 111.528 94.068 ; 
        RECT 110.992 89.694 111.096 94.068 ; 
        RECT 110.56 89.694 110.664 94.068 ; 
        RECT 110.128 89.694 110.232 94.068 ; 
        RECT 109.696 89.694 109.8 94.068 ; 
        RECT 109.264 89.694 109.368 94.068 ; 
        RECT 108.832 89.694 108.936 94.068 ; 
        RECT 108.4 89.694 108.504 94.068 ; 
        RECT 107.968 89.694 108.072 94.068 ; 
        RECT 107.536 89.694 107.64 94.068 ; 
        RECT 107.104 89.694 107.208 94.068 ; 
        RECT 106.672 89.694 106.776 94.068 ; 
        RECT 106.24 89.694 106.344 94.068 ; 
        RECT 105.808 89.694 105.912 94.068 ; 
        RECT 105.376 89.694 105.48 94.068 ; 
        RECT 104.944 89.694 105.048 94.068 ; 
        RECT 104.512 89.694 104.616 94.068 ; 
        RECT 104.08 89.694 104.184 94.068 ; 
        RECT 103.648 89.694 103.752 94.068 ; 
        RECT 103.216 89.694 103.32 94.068 ; 
        RECT 102.784 89.694 102.888 94.068 ; 
        RECT 102.352 89.694 102.456 94.068 ; 
        RECT 101.92 89.694 102.024 94.068 ; 
        RECT 101.488 89.694 101.592 94.068 ; 
        RECT 101.056 89.694 101.16 94.068 ; 
        RECT 100.624 89.694 100.728 94.068 ; 
        RECT 100.192 89.694 100.296 94.068 ; 
        RECT 99.76 89.694 99.864 94.068 ; 
        RECT 99.328 89.694 99.432 94.068 ; 
        RECT 98.896 89.694 99 94.068 ; 
        RECT 98.464 89.694 98.568 94.068 ; 
        RECT 98.032 89.694 98.136 94.068 ; 
        RECT 97.6 89.694 97.704 94.068 ; 
        RECT 97.168 89.694 97.272 94.068 ; 
        RECT 96.736 89.694 96.84 94.068 ; 
        RECT 96.304 89.694 96.408 94.068 ; 
        RECT 95.872 89.694 95.976 94.068 ; 
        RECT 95.44 89.694 95.544 94.068 ; 
        RECT 95.008 89.694 95.112 94.068 ; 
        RECT 94.576 89.694 94.68 94.068 ; 
        RECT 94.144 89.694 94.248 94.068 ; 
        RECT 93.712 89.694 93.816 94.068 ; 
        RECT 93.28 89.694 93.384 94.068 ; 
        RECT 92.848 89.694 92.952 94.068 ; 
        RECT 92.416 89.694 92.52 94.068 ; 
        RECT 91.984 89.694 92.088 94.068 ; 
        RECT 91.552 89.694 91.656 94.068 ; 
        RECT 91.12 89.694 91.224 94.068 ; 
        RECT 90.688 89.694 90.792 94.068 ; 
        RECT 90.256 89.694 90.36 94.068 ; 
        RECT 89.824 89.694 89.928 94.068 ; 
        RECT 89.392 89.694 89.496 94.068 ; 
        RECT 88.96 89.694 89.064 94.068 ; 
        RECT 88.528 89.694 88.632 94.068 ; 
        RECT 88.096 89.694 88.2 94.068 ; 
        RECT 87.664 89.694 87.768 94.068 ; 
        RECT 87.232 89.694 87.336 94.068 ; 
        RECT 86.8 89.694 86.904 94.068 ; 
        RECT 86.368 89.694 86.472 94.068 ; 
        RECT 85.936 89.694 86.04 94.068 ; 
        RECT 85.504 89.694 85.608 94.068 ; 
        RECT 85.072 89.694 85.176 94.068 ; 
        RECT 84.64 89.694 84.744 94.068 ; 
        RECT 84.208 89.694 84.312 94.068 ; 
        RECT 83.776 89.694 83.88 94.068 ; 
        RECT 83.344 89.694 83.448 94.068 ; 
        RECT 82.912 89.694 83.016 94.068 ; 
        RECT 82.48 89.694 82.584 94.068 ; 
        RECT 82.048 89.694 82.152 94.068 ; 
        RECT 81.616 89.694 81.72 94.068 ; 
        RECT 81.184 89.694 81.288 94.068 ; 
        RECT 80.752 89.694 80.856 94.068 ; 
        RECT 80.32 89.694 80.424 94.068 ; 
        RECT 79.888 89.694 79.992 94.068 ; 
        RECT 79.456 89.694 79.56 94.068 ; 
        RECT 79.024 89.694 79.128 94.068 ; 
        RECT 78.592 89.694 78.696 94.068 ; 
        RECT 78.16 89.694 78.264 94.068 ; 
        RECT 77.728 89.694 77.832 94.068 ; 
        RECT 77.296 89.694 77.4 94.068 ; 
        RECT 76.864 89.694 76.968 94.068 ; 
        RECT 76.432 89.694 76.536 94.068 ; 
        RECT 76 89.694 76.104 94.068 ; 
        RECT 75.568 89.694 75.672 94.068 ; 
        RECT 75.136 89.694 75.24 94.068 ; 
        RECT 74.704 89.694 74.808 94.068 ; 
        RECT 74.272 89.694 74.376 94.068 ; 
        RECT 73.84 89.694 73.944 94.068 ; 
        RECT 73.408 89.694 73.512 94.068 ; 
        RECT 72.976 89.694 73.08 94.068 ; 
        RECT 72.544 89.694 72.648 94.068 ; 
        RECT 72.112 89.694 72.216 94.068 ; 
        RECT 71.68 89.694 71.784 94.068 ; 
        RECT 71.248 89.694 71.352 94.068 ; 
        RECT 70.816 89.694 70.92 94.068 ; 
        RECT 70.384 89.694 70.488 94.068 ; 
        RECT 69.952 89.694 70.056 94.068 ; 
        RECT 69.52 89.694 69.624 94.068 ; 
        RECT 69.088 89.694 69.192 94.068 ; 
        RECT 68.656 89.694 68.76 94.068 ; 
        RECT 68.224 89.694 68.328 94.068 ; 
        RECT 67.792 89.694 67.896 94.068 ; 
        RECT 67.36 89.694 67.464 94.068 ; 
        RECT 66.928 89.694 67.032 94.068 ; 
        RECT 66.496 89.694 66.6 94.068 ; 
        RECT 66.064 89.694 66.168 94.068 ; 
        RECT 65.632 89.694 65.736 94.068 ; 
        RECT 65.2 89.694 65.304 94.068 ; 
        RECT 64.348 89.694 64.656 94.068 ; 
        RECT 56.776 89.694 57.084 94.068 ; 
        RECT 56.128 89.694 56.232 94.068 ; 
        RECT 55.696 89.694 55.8 94.068 ; 
        RECT 55.264 89.694 55.368 94.068 ; 
        RECT 54.832 89.694 54.936 94.068 ; 
        RECT 54.4 89.694 54.504 94.068 ; 
        RECT 53.968 89.694 54.072 94.068 ; 
        RECT 53.536 89.694 53.64 94.068 ; 
        RECT 53.104 89.694 53.208 94.068 ; 
        RECT 52.672 89.694 52.776 94.068 ; 
        RECT 52.24 89.694 52.344 94.068 ; 
        RECT 51.808 89.694 51.912 94.068 ; 
        RECT 51.376 89.694 51.48 94.068 ; 
        RECT 50.944 89.694 51.048 94.068 ; 
        RECT 50.512 89.694 50.616 94.068 ; 
        RECT 50.08 89.694 50.184 94.068 ; 
        RECT 49.648 89.694 49.752 94.068 ; 
        RECT 49.216 89.694 49.32 94.068 ; 
        RECT 48.784 89.694 48.888 94.068 ; 
        RECT 48.352 89.694 48.456 94.068 ; 
        RECT 47.92 89.694 48.024 94.068 ; 
        RECT 47.488 89.694 47.592 94.068 ; 
        RECT 47.056 89.694 47.16 94.068 ; 
        RECT 46.624 89.694 46.728 94.068 ; 
        RECT 46.192 89.694 46.296 94.068 ; 
        RECT 45.76 89.694 45.864 94.068 ; 
        RECT 45.328 89.694 45.432 94.068 ; 
        RECT 44.896 89.694 45 94.068 ; 
        RECT 44.464 89.694 44.568 94.068 ; 
        RECT 44.032 89.694 44.136 94.068 ; 
        RECT 43.6 89.694 43.704 94.068 ; 
        RECT 43.168 89.694 43.272 94.068 ; 
        RECT 42.736 89.694 42.84 94.068 ; 
        RECT 42.304 89.694 42.408 94.068 ; 
        RECT 41.872 89.694 41.976 94.068 ; 
        RECT 41.44 89.694 41.544 94.068 ; 
        RECT 41.008 89.694 41.112 94.068 ; 
        RECT 40.576 89.694 40.68 94.068 ; 
        RECT 40.144 89.694 40.248 94.068 ; 
        RECT 39.712 89.694 39.816 94.068 ; 
        RECT 39.28 89.694 39.384 94.068 ; 
        RECT 38.848 89.694 38.952 94.068 ; 
        RECT 38.416 89.694 38.52 94.068 ; 
        RECT 37.984 89.694 38.088 94.068 ; 
        RECT 37.552 89.694 37.656 94.068 ; 
        RECT 37.12 89.694 37.224 94.068 ; 
        RECT 36.688 89.694 36.792 94.068 ; 
        RECT 36.256 89.694 36.36 94.068 ; 
        RECT 35.824 89.694 35.928 94.068 ; 
        RECT 35.392 89.694 35.496 94.068 ; 
        RECT 34.96 89.694 35.064 94.068 ; 
        RECT 34.528 89.694 34.632 94.068 ; 
        RECT 34.096 89.694 34.2 94.068 ; 
        RECT 33.664 89.694 33.768 94.068 ; 
        RECT 33.232 89.694 33.336 94.068 ; 
        RECT 32.8 89.694 32.904 94.068 ; 
        RECT 32.368 89.694 32.472 94.068 ; 
        RECT 31.936 89.694 32.04 94.068 ; 
        RECT 31.504 89.694 31.608 94.068 ; 
        RECT 31.072 89.694 31.176 94.068 ; 
        RECT 30.64 89.694 30.744 94.068 ; 
        RECT 30.208 89.694 30.312 94.068 ; 
        RECT 29.776 89.694 29.88 94.068 ; 
        RECT 29.344 89.694 29.448 94.068 ; 
        RECT 28.912 89.694 29.016 94.068 ; 
        RECT 28.48 89.694 28.584 94.068 ; 
        RECT 28.048 89.694 28.152 94.068 ; 
        RECT 27.616 89.694 27.72 94.068 ; 
        RECT 27.184 89.694 27.288 94.068 ; 
        RECT 26.752 89.694 26.856 94.068 ; 
        RECT 26.32 89.694 26.424 94.068 ; 
        RECT 25.888 89.694 25.992 94.068 ; 
        RECT 25.456 89.694 25.56 94.068 ; 
        RECT 25.024 89.694 25.128 94.068 ; 
        RECT 24.592 89.694 24.696 94.068 ; 
        RECT 24.16 89.694 24.264 94.068 ; 
        RECT 23.728 89.694 23.832 94.068 ; 
        RECT 23.296 89.694 23.4 94.068 ; 
        RECT 22.864 89.694 22.968 94.068 ; 
        RECT 22.432 89.694 22.536 94.068 ; 
        RECT 22 89.694 22.104 94.068 ; 
        RECT 21.568 89.694 21.672 94.068 ; 
        RECT 21.136 89.694 21.24 94.068 ; 
        RECT 20.704 89.694 20.808 94.068 ; 
        RECT 20.272 89.694 20.376 94.068 ; 
        RECT 19.84 89.694 19.944 94.068 ; 
        RECT 19.408 89.694 19.512 94.068 ; 
        RECT 18.976 89.694 19.08 94.068 ; 
        RECT 18.544 89.694 18.648 94.068 ; 
        RECT 18.112 89.694 18.216 94.068 ; 
        RECT 17.68 89.694 17.784 94.068 ; 
        RECT 17.248 89.694 17.352 94.068 ; 
        RECT 16.816 89.694 16.92 94.068 ; 
        RECT 16.384 89.694 16.488 94.068 ; 
        RECT 15.952 89.694 16.056 94.068 ; 
        RECT 15.52 89.694 15.624 94.068 ; 
        RECT 15.088 89.694 15.192 94.068 ; 
        RECT 14.656 89.694 14.76 94.068 ; 
        RECT 14.224 89.694 14.328 94.068 ; 
        RECT 13.792 89.694 13.896 94.068 ; 
        RECT 13.36 89.694 13.464 94.068 ; 
        RECT 12.928 89.694 13.032 94.068 ; 
        RECT 12.496 89.694 12.6 94.068 ; 
        RECT 12.064 89.694 12.168 94.068 ; 
        RECT 11.632 89.694 11.736 94.068 ; 
        RECT 11.2 89.694 11.304 94.068 ; 
        RECT 10.768 89.694 10.872 94.068 ; 
        RECT 10.336 89.694 10.44 94.068 ; 
        RECT 9.904 89.694 10.008 94.068 ; 
        RECT 9.472 89.694 9.576 94.068 ; 
        RECT 9.04 89.694 9.144 94.068 ; 
        RECT 8.608 89.694 8.712 94.068 ; 
        RECT 8.176 89.694 8.28 94.068 ; 
        RECT 7.744 89.694 7.848 94.068 ; 
        RECT 7.312 89.694 7.416 94.068 ; 
        RECT 6.88 89.694 6.984 94.068 ; 
        RECT 6.448 89.694 6.552 94.068 ; 
        RECT 6.016 89.694 6.12 94.068 ; 
        RECT 5.584 89.694 5.688 94.068 ; 
        RECT 5.152 89.694 5.256 94.068 ; 
        RECT 4.72 89.694 4.824 94.068 ; 
        RECT 4.288 89.694 4.392 94.068 ; 
        RECT 3.856 89.694 3.96 94.068 ; 
        RECT 3.424 89.694 3.528 94.068 ; 
        RECT 2.992 89.694 3.096 94.068 ; 
        RECT 2.56 89.694 2.664 94.068 ; 
        RECT 2.128 89.694 2.232 94.068 ; 
        RECT 1.696 89.694 1.8 94.068 ; 
        RECT 1.264 89.694 1.368 94.068 ; 
        RECT 0.832 89.694 0.936 94.068 ; 
        RECT 0.02 89.694 0.36 94.068 ; 
        RECT 62.212 94.014 62.724 98.388 ; 
        RECT 62.156 96.676 62.724 97.966 ; 
        RECT 61.276 95.584 61.812 98.388 ; 
        RECT 61.184 96.924 61.812 97.956 ; 
        RECT 61.276 94.014 61.668 98.388 ; 
        RECT 61.276 94.498 61.724 95.456 ; 
        RECT 61.276 94.014 61.812 94.37 ; 
        RECT 60.376 95.816 60.912 98.388 ; 
        RECT 60.376 94.014 60.768 98.388 ; 
        RECT 58.708 94.014 59.04 98.388 ; 
        RECT 58.708 94.368 59.096 98.11 ; 
        RECT 121.072 94.014 121.412 98.388 ; 
        RECT 120.496 94.014 120.6 98.388 ; 
        RECT 120.064 94.014 120.168 98.388 ; 
        RECT 119.632 94.014 119.736 98.388 ; 
        RECT 119.2 94.014 119.304 98.388 ; 
        RECT 118.768 94.014 118.872 98.388 ; 
        RECT 118.336 94.014 118.44 98.388 ; 
        RECT 117.904 94.014 118.008 98.388 ; 
        RECT 117.472 94.014 117.576 98.388 ; 
        RECT 117.04 94.014 117.144 98.388 ; 
        RECT 116.608 94.014 116.712 98.388 ; 
        RECT 116.176 94.014 116.28 98.388 ; 
        RECT 115.744 94.014 115.848 98.388 ; 
        RECT 115.312 94.014 115.416 98.388 ; 
        RECT 114.88 94.014 114.984 98.388 ; 
        RECT 114.448 94.014 114.552 98.388 ; 
        RECT 114.016 94.014 114.12 98.388 ; 
        RECT 113.584 94.014 113.688 98.388 ; 
        RECT 113.152 94.014 113.256 98.388 ; 
        RECT 112.72 94.014 112.824 98.388 ; 
        RECT 112.288 94.014 112.392 98.388 ; 
        RECT 111.856 94.014 111.96 98.388 ; 
        RECT 111.424 94.014 111.528 98.388 ; 
        RECT 110.992 94.014 111.096 98.388 ; 
        RECT 110.56 94.014 110.664 98.388 ; 
        RECT 110.128 94.014 110.232 98.388 ; 
        RECT 109.696 94.014 109.8 98.388 ; 
        RECT 109.264 94.014 109.368 98.388 ; 
        RECT 108.832 94.014 108.936 98.388 ; 
        RECT 108.4 94.014 108.504 98.388 ; 
        RECT 107.968 94.014 108.072 98.388 ; 
        RECT 107.536 94.014 107.64 98.388 ; 
        RECT 107.104 94.014 107.208 98.388 ; 
        RECT 106.672 94.014 106.776 98.388 ; 
        RECT 106.24 94.014 106.344 98.388 ; 
        RECT 105.808 94.014 105.912 98.388 ; 
        RECT 105.376 94.014 105.48 98.388 ; 
        RECT 104.944 94.014 105.048 98.388 ; 
        RECT 104.512 94.014 104.616 98.388 ; 
        RECT 104.08 94.014 104.184 98.388 ; 
        RECT 103.648 94.014 103.752 98.388 ; 
        RECT 103.216 94.014 103.32 98.388 ; 
        RECT 102.784 94.014 102.888 98.388 ; 
        RECT 102.352 94.014 102.456 98.388 ; 
        RECT 101.92 94.014 102.024 98.388 ; 
        RECT 101.488 94.014 101.592 98.388 ; 
        RECT 101.056 94.014 101.16 98.388 ; 
        RECT 100.624 94.014 100.728 98.388 ; 
        RECT 100.192 94.014 100.296 98.388 ; 
        RECT 99.76 94.014 99.864 98.388 ; 
        RECT 99.328 94.014 99.432 98.388 ; 
        RECT 98.896 94.014 99 98.388 ; 
        RECT 98.464 94.014 98.568 98.388 ; 
        RECT 98.032 94.014 98.136 98.388 ; 
        RECT 97.6 94.014 97.704 98.388 ; 
        RECT 97.168 94.014 97.272 98.388 ; 
        RECT 96.736 94.014 96.84 98.388 ; 
        RECT 96.304 94.014 96.408 98.388 ; 
        RECT 95.872 94.014 95.976 98.388 ; 
        RECT 95.44 94.014 95.544 98.388 ; 
        RECT 95.008 94.014 95.112 98.388 ; 
        RECT 94.576 94.014 94.68 98.388 ; 
        RECT 94.144 94.014 94.248 98.388 ; 
        RECT 93.712 94.014 93.816 98.388 ; 
        RECT 93.28 94.014 93.384 98.388 ; 
        RECT 92.848 94.014 92.952 98.388 ; 
        RECT 92.416 94.014 92.52 98.388 ; 
        RECT 91.984 94.014 92.088 98.388 ; 
        RECT 91.552 94.014 91.656 98.388 ; 
        RECT 91.12 94.014 91.224 98.388 ; 
        RECT 90.688 94.014 90.792 98.388 ; 
        RECT 90.256 94.014 90.36 98.388 ; 
        RECT 89.824 94.014 89.928 98.388 ; 
        RECT 89.392 94.014 89.496 98.388 ; 
        RECT 88.96 94.014 89.064 98.388 ; 
        RECT 88.528 94.014 88.632 98.388 ; 
        RECT 88.096 94.014 88.2 98.388 ; 
        RECT 87.664 94.014 87.768 98.388 ; 
        RECT 87.232 94.014 87.336 98.388 ; 
        RECT 86.8 94.014 86.904 98.388 ; 
        RECT 86.368 94.014 86.472 98.388 ; 
        RECT 85.936 94.014 86.04 98.388 ; 
        RECT 85.504 94.014 85.608 98.388 ; 
        RECT 85.072 94.014 85.176 98.388 ; 
        RECT 84.64 94.014 84.744 98.388 ; 
        RECT 84.208 94.014 84.312 98.388 ; 
        RECT 83.776 94.014 83.88 98.388 ; 
        RECT 83.344 94.014 83.448 98.388 ; 
        RECT 82.912 94.014 83.016 98.388 ; 
        RECT 82.48 94.014 82.584 98.388 ; 
        RECT 82.048 94.014 82.152 98.388 ; 
        RECT 81.616 94.014 81.72 98.388 ; 
        RECT 81.184 94.014 81.288 98.388 ; 
        RECT 80.752 94.014 80.856 98.388 ; 
        RECT 80.32 94.014 80.424 98.388 ; 
        RECT 79.888 94.014 79.992 98.388 ; 
        RECT 79.456 94.014 79.56 98.388 ; 
        RECT 79.024 94.014 79.128 98.388 ; 
        RECT 78.592 94.014 78.696 98.388 ; 
        RECT 78.16 94.014 78.264 98.388 ; 
        RECT 77.728 94.014 77.832 98.388 ; 
        RECT 77.296 94.014 77.4 98.388 ; 
        RECT 76.864 94.014 76.968 98.388 ; 
        RECT 76.432 94.014 76.536 98.388 ; 
        RECT 76 94.014 76.104 98.388 ; 
        RECT 75.568 94.014 75.672 98.388 ; 
        RECT 75.136 94.014 75.24 98.388 ; 
        RECT 74.704 94.014 74.808 98.388 ; 
        RECT 74.272 94.014 74.376 98.388 ; 
        RECT 73.84 94.014 73.944 98.388 ; 
        RECT 73.408 94.014 73.512 98.388 ; 
        RECT 72.976 94.014 73.08 98.388 ; 
        RECT 72.544 94.014 72.648 98.388 ; 
        RECT 72.112 94.014 72.216 98.388 ; 
        RECT 71.68 94.014 71.784 98.388 ; 
        RECT 71.248 94.014 71.352 98.388 ; 
        RECT 70.816 94.014 70.92 98.388 ; 
        RECT 70.384 94.014 70.488 98.388 ; 
        RECT 69.952 94.014 70.056 98.388 ; 
        RECT 69.52 94.014 69.624 98.388 ; 
        RECT 69.088 94.014 69.192 98.388 ; 
        RECT 68.656 94.014 68.76 98.388 ; 
        RECT 68.224 94.014 68.328 98.388 ; 
        RECT 67.792 94.014 67.896 98.388 ; 
        RECT 67.36 94.014 67.464 98.388 ; 
        RECT 66.928 94.014 67.032 98.388 ; 
        RECT 66.496 94.014 66.6 98.388 ; 
        RECT 66.064 94.014 66.168 98.388 ; 
        RECT 65.632 94.014 65.736 98.388 ; 
        RECT 65.2 94.014 65.304 98.388 ; 
        RECT 64.348 94.014 64.656 98.388 ; 
        RECT 56.776 94.014 57.084 98.388 ; 
        RECT 56.128 94.014 56.232 98.388 ; 
        RECT 55.696 94.014 55.8 98.388 ; 
        RECT 55.264 94.014 55.368 98.388 ; 
        RECT 54.832 94.014 54.936 98.388 ; 
        RECT 54.4 94.014 54.504 98.388 ; 
        RECT 53.968 94.014 54.072 98.388 ; 
        RECT 53.536 94.014 53.64 98.388 ; 
        RECT 53.104 94.014 53.208 98.388 ; 
        RECT 52.672 94.014 52.776 98.388 ; 
        RECT 52.24 94.014 52.344 98.388 ; 
        RECT 51.808 94.014 51.912 98.388 ; 
        RECT 51.376 94.014 51.48 98.388 ; 
        RECT 50.944 94.014 51.048 98.388 ; 
        RECT 50.512 94.014 50.616 98.388 ; 
        RECT 50.08 94.014 50.184 98.388 ; 
        RECT 49.648 94.014 49.752 98.388 ; 
        RECT 49.216 94.014 49.32 98.388 ; 
        RECT 48.784 94.014 48.888 98.388 ; 
        RECT 48.352 94.014 48.456 98.388 ; 
        RECT 47.92 94.014 48.024 98.388 ; 
        RECT 47.488 94.014 47.592 98.388 ; 
        RECT 47.056 94.014 47.16 98.388 ; 
        RECT 46.624 94.014 46.728 98.388 ; 
        RECT 46.192 94.014 46.296 98.388 ; 
        RECT 45.76 94.014 45.864 98.388 ; 
        RECT 45.328 94.014 45.432 98.388 ; 
        RECT 44.896 94.014 45 98.388 ; 
        RECT 44.464 94.014 44.568 98.388 ; 
        RECT 44.032 94.014 44.136 98.388 ; 
        RECT 43.6 94.014 43.704 98.388 ; 
        RECT 43.168 94.014 43.272 98.388 ; 
        RECT 42.736 94.014 42.84 98.388 ; 
        RECT 42.304 94.014 42.408 98.388 ; 
        RECT 41.872 94.014 41.976 98.388 ; 
        RECT 41.44 94.014 41.544 98.388 ; 
        RECT 41.008 94.014 41.112 98.388 ; 
        RECT 40.576 94.014 40.68 98.388 ; 
        RECT 40.144 94.014 40.248 98.388 ; 
        RECT 39.712 94.014 39.816 98.388 ; 
        RECT 39.28 94.014 39.384 98.388 ; 
        RECT 38.848 94.014 38.952 98.388 ; 
        RECT 38.416 94.014 38.52 98.388 ; 
        RECT 37.984 94.014 38.088 98.388 ; 
        RECT 37.552 94.014 37.656 98.388 ; 
        RECT 37.12 94.014 37.224 98.388 ; 
        RECT 36.688 94.014 36.792 98.388 ; 
        RECT 36.256 94.014 36.36 98.388 ; 
        RECT 35.824 94.014 35.928 98.388 ; 
        RECT 35.392 94.014 35.496 98.388 ; 
        RECT 34.96 94.014 35.064 98.388 ; 
        RECT 34.528 94.014 34.632 98.388 ; 
        RECT 34.096 94.014 34.2 98.388 ; 
        RECT 33.664 94.014 33.768 98.388 ; 
        RECT 33.232 94.014 33.336 98.388 ; 
        RECT 32.8 94.014 32.904 98.388 ; 
        RECT 32.368 94.014 32.472 98.388 ; 
        RECT 31.936 94.014 32.04 98.388 ; 
        RECT 31.504 94.014 31.608 98.388 ; 
        RECT 31.072 94.014 31.176 98.388 ; 
        RECT 30.64 94.014 30.744 98.388 ; 
        RECT 30.208 94.014 30.312 98.388 ; 
        RECT 29.776 94.014 29.88 98.388 ; 
        RECT 29.344 94.014 29.448 98.388 ; 
        RECT 28.912 94.014 29.016 98.388 ; 
        RECT 28.48 94.014 28.584 98.388 ; 
        RECT 28.048 94.014 28.152 98.388 ; 
        RECT 27.616 94.014 27.72 98.388 ; 
        RECT 27.184 94.014 27.288 98.388 ; 
        RECT 26.752 94.014 26.856 98.388 ; 
        RECT 26.32 94.014 26.424 98.388 ; 
        RECT 25.888 94.014 25.992 98.388 ; 
        RECT 25.456 94.014 25.56 98.388 ; 
        RECT 25.024 94.014 25.128 98.388 ; 
        RECT 24.592 94.014 24.696 98.388 ; 
        RECT 24.16 94.014 24.264 98.388 ; 
        RECT 23.728 94.014 23.832 98.388 ; 
        RECT 23.296 94.014 23.4 98.388 ; 
        RECT 22.864 94.014 22.968 98.388 ; 
        RECT 22.432 94.014 22.536 98.388 ; 
        RECT 22 94.014 22.104 98.388 ; 
        RECT 21.568 94.014 21.672 98.388 ; 
        RECT 21.136 94.014 21.24 98.388 ; 
        RECT 20.704 94.014 20.808 98.388 ; 
        RECT 20.272 94.014 20.376 98.388 ; 
        RECT 19.84 94.014 19.944 98.388 ; 
        RECT 19.408 94.014 19.512 98.388 ; 
        RECT 18.976 94.014 19.08 98.388 ; 
        RECT 18.544 94.014 18.648 98.388 ; 
        RECT 18.112 94.014 18.216 98.388 ; 
        RECT 17.68 94.014 17.784 98.388 ; 
        RECT 17.248 94.014 17.352 98.388 ; 
        RECT 16.816 94.014 16.92 98.388 ; 
        RECT 16.384 94.014 16.488 98.388 ; 
        RECT 15.952 94.014 16.056 98.388 ; 
        RECT 15.52 94.014 15.624 98.388 ; 
        RECT 15.088 94.014 15.192 98.388 ; 
        RECT 14.656 94.014 14.76 98.388 ; 
        RECT 14.224 94.014 14.328 98.388 ; 
        RECT 13.792 94.014 13.896 98.388 ; 
        RECT 13.36 94.014 13.464 98.388 ; 
        RECT 12.928 94.014 13.032 98.388 ; 
        RECT 12.496 94.014 12.6 98.388 ; 
        RECT 12.064 94.014 12.168 98.388 ; 
        RECT 11.632 94.014 11.736 98.388 ; 
        RECT 11.2 94.014 11.304 98.388 ; 
        RECT 10.768 94.014 10.872 98.388 ; 
        RECT 10.336 94.014 10.44 98.388 ; 
        RECT 9.904 94.014 10.008 98.388 ; 
        RECT 9.472 94.014 9.576 98.388 ; 
        RECT 9.04 94.014 9.144 98.388 ; 
        RECT 8.608 94.014 8.712 98.388 ; 
        RECT 8.176 94.014 8.28 98.388 ; 
        RECT 7.744 94.014 7.848 98.388 ; 
        RECT 7.312 94.014 7.416 98.388 ; 
        RECT 6.88 94.014 6.984 98.388 ; 
        RECT 6.448 94.014 6.552 98.388 ; 
        RECT 6.016 94.014 6.12 98.388 ; 
        RECT 5.584 94.014 5.688 98.388 ; 
        RECT 5.152 94.014 5.256 98.388 ; 
        RECT 4.72 94.014 4.824 98.388 ; 
        RECT 4.288 94.014 4.392 98.388 ; 
        RECT 3.856 94.014 3.96 98.388 ; 
        RECT 3.424 94.014 3.528 98.388 ; 
        RECT 2.992 94.014 3.096 98.388 ; 
        RECT 2.56 94.014 2.664 98.388 ; 
        RECT 2.128 94.014 2.232 98.388 ; 
        RECT 1.696 94.014 1.8 98.388 ; 
        RECT 1.264 94.014 1.368 98.388 ; 
        RECT 0.832 94.014 0.936 98.388 ; 
        RECT 0.02 94.014 0.36 98.388 ; 
        RECT 62.212 98.334 62.724 102.708 ; 
        RECT 62.156 100.996 62.724 102.286 ; 
        RECT 61.276 99.904 61.812 102.708 ; 
        RECT 61.184 101.244 61.812 102.276 ; 
        RECT 61.276 98.334 61.668 102.708 ; 
        RECT 61.276 98.818 61.724 99.776 ; 
        RECT 61.276 98.334 61.812 98.69 ; 
        RECT 60.376 100.136 60.912 102.708 ; 
        RECT 60.376 98.334 60.768 102.708 ; 
        RECT 58.708 98.334 59.04 102.708 ; 
        RECT 58.708 98.688 59.096 102.43 ; 
        RECT 121.072 98.334 121.412 102.708 ; 
        RECT 120.496 98.334 120.6 102.708 ; 
        RECT 120.064 98.334 120.168 102.708 ; 
        RECT 119.632 98.334 119.736 102.708 ; 
        RECT 119.2 98.334 119.304 102.708 ; 
        RECT 118.768 98.334 118.872 102.708 ; 
        RECT 118.336 98.334 118.44 102.708 ; 
        RECT 117.904 98.334 118.008 102.708 ; 
        RECT 117.472 98.334 117.576 102.708 ; 
        RECT 117.04 98.334 117.144 102.708 ; 
        RECT 116.608 98.334 116.712 102.708 ; 
        RECT 116.176 98.334 116.28 102.708 ; 
        RECT 115.744 98.334 115.848 102.708 ; 
        RECT 115.312 98.334 115.416 102.708 ; 
        RECT 114.88 98.334 114.984 102.708 ; 
        RECT 114.448 98.334 114.552 102.708 ; 
        RECT 114.016 98.334 114.12 102.708 ; 
        RECT 113.584 98.334 113.688 102.708 ; 
        RECT 113.152 98.334 113.256 102.708 ; 
        RECT 112.72 98.334 112.824 102.708 ; 
        RECT 112.288 98.334 112.392 102.708 ; 
        RECT 111.856 98.334 111.96 102.708 ; 
        RECT 111.424 98.334 111.528 102.708 ; 
        RECT 110.992 98.334 111.096 102.708 ; 
        RECT 110.56 98.334 110.664 102.708 ; 
        RECT 110.128 98.334 110.232 102.708 ; 
        RECT 109.696 98.334 109.8 102.708 ; 
        RECT 109.264 98.334 109.368 102.708 ; 
        RECT 108.832 98.334 108.936 102.708 ; 
        RECT 108.4 98.334 108.504 102.708 ; 
        RECT 107.968 98.334 108.072 102.708 ; 
        RECT 107.536 98.334 107.64 102.708 ; 
        RECT 107.104 98.334 107.208 102.708 ; 
        RECT 106.672 98.334 106.776 102.708 ; 
        RECT 106.24 98.334 106.344 102.708 ; 
        RECT 105.808 98.334 105.912 102.708 ; 
        RECT 105.376 98.334 105.48 102.708 ; 
        RECT 104.944 98.334 105.048 102.708 ; 
        RECT 104.512 98.334 104.616 102.708 ; 
        RECT 104.08 98.334 104.184 102.708 ; 
        RECT 103.648 98.334 103.752 102.708 ; 
        RECT 103.216 98.334 103.32 102.708 ; 
        RECT 102.784 98.334 102.888 102.708 ; 
        RECT 102.352 98.334 102.456 102.708 ; 
        RECT 101.92 98.334 102.024 102.708 ; 
        RECT 101.488 98.334 101.592 102.708 ; 
        RECT 101.056 98.334 101.16 102.708 ; 
        RECT 100.624 98.334 100.728 102.708 ; 
        RECT 100.192 98.334 100.296 102.708 ; 
        RECT 99.76 98.334 99.864 102.708 ; 
        RECT 99.328 98.334 99.432 102.708 ; 
        RECT 98.896 98.334 99 102.708 ; 
        RECT 98.464 98.334 98.568 102.708 ; 
        RECT 98.032 98.334 98.136 102.708 ; 
        RECT 97.6 98.334 97.704 102.708 ; 
        RECT 97.168 98.334 97.272 102.708 ; 
        RECT 96.736 98.334 96.84 102.708 ; 
        RECT 96.304 98.334 96.408 102.708 ; 
        RECT 95.872 98.334 95.976 102.708 ; 
        RECT 95.44 98.334 95.544 102.708 ; 
        RECT 95.008 98.334 95.112 102.708 ; 
        RECT 94.576 98.334 94.68 102.708 ; 
        RECT 94.144 98.334 94.248 102.708 ; 
        RECT 93.712 98.334 93.816 102.708 ; 
        RECT 93.28 98.334 93.384 102.708 ; 
        RECT 92.848 98.334 92.952 102.708 ; 
        RECT 92.416 98.334 92.52 102.708 ; 
        RECT 91.984 98.334 92.088 102.708 ; 
        RECT 91.552 98.334 91.656 102.708 ; 
        RECT 91.12 98.334 91.224 102.708 ; 
        RECT 90.688 98.334 90.792 102.708 ; 
        RECT 90.256 98.334 90.36 102.708 ; 
        RECT 89.824 98.334 89.928 102.708 ; 
        RECT 89.392 98.334 89.496 102.708 ; 
        RECT 88.96 98.334 89.064 102.708 ; 
        RECT 88.528 98.334 88.632 102.708 ; 
        RECT 88.096 98.334 88.2 102.708 ; 
        RECT 87.664 98.334 87.768 102.708 ; 
        RECT 87.232 98.334 87.336 102.708 ; 
        RECT 86.8 98.334 86.904 102.708 ; 
        RECT 86.368 98.334 86.472 102.708 ; 
        RECT 85.936 98.334 86.04 102.708 ; 
        RECT 85.504 98.334 85.608 102.708 ; 
        RECT 85.072 98.334 85.176 102.708 ; 
        RECT 84.64 98.334 84.744 102.708 ; 
        RECT 84.208 98.334 84.312 102.708 ; 
        RECT 83.776 98.334 83.88 102.708 ; 
        RECT 83.344 98.334 83.448 102.708 ; 
        RECT 82.912 98.334 83.016 102.708 ; 
        RECT 82.48 98.334 82.584 102.708 ; 
        RECT 82.048 98.334 82.152 102.708 ; 
        RECT 81.616 98.334 81.72 102.708 ; 
        RECT 81.184 98.334 81.288 102.708 ; 
        RECT 80.752 98.334 80.856 102.708 ; 
        RECT 80.32 98.334 80.424 102.708 ; 
        RECT 79.888 98.334 79.992 102.708 ; 
        RECT 79.456 98.334 79.56 102.708 ; 
        RECT 79.024 98.334 79.128 102.708 ; 
        RECT 78.592 98.334 78.696 102.708 ; 
        RECT 78.16 98.334 78.264 102.708 ; 
        RECT 77.728 98.334 77.832 102.708 ; 
        RECT 77.296 98.334 77.4 102.708 ; 
        RECT 76.864 98.334 76.968 102.708 ; 
        RECT 76.432 98.334 76.536 102.708 ; 
        RECT 76 98.334 76.104 102.708 ; 
        RECT 75.568 98.334 75.672 102.708 ; 
        RECT 75.136 98.334 75.24 102.708 ; 
        RECT 74.704 98.334 74.808 102.708 ; 
        RECT 74.272 98.334 74.376 102.708 ; 
        RECT 73.84 98.334 73.944 102.708 ; 
        RECT 73.408 98.334 73.512 102.708 ; 
        RECT 72.976 98.334 73.08 102.708 ; 
        RECT 72.544 98.334 72.648 102.708 ; 
        RECT 72.112 98.334 72.216 102.708 ; 
        RECT 71.68 98.334 71.784 102.708 ; 
        RECT 71.248 98.334 71.352 102.708 ; 
        RECT 70.816 98.334 70.92 102.708 ; 
        RECT 70.384 98.334 70.488 102.708 ; 
        RECT 69.952 98.334 70.056 102.708 ; 
        RECT 69.52 98.334 69.624 102.708 ; 
        RECT 69.088 98.334 69.192 102.708 ; 
        RECT 68.656 98.334 68.76 102.708 ; 
        RECT 68.224 98.334 68.328 102.708 ; 
        RECT 67.792 98.334 67.896 102.708 ; 
        RECT 67.36 98.334 67.464 102.708 ; 
        RECT 66.928 98.334 67.032 102.708 ; 
        RECT 66.496 98.334 66.6 102.708 ; 
        RECT 66.064 98.334 66.168 102.708 ; 
        RECT 65.632 98.334 65.736 102.708 ; 
        RECT 65.2 98.334 65.304 102.708 ; 
        RECT 64.348 98.334 64.656 102.708 ; 
        RECT 56.776 98.334 57.084 102.708 ; 
        RECT 56.128 98.334 56.232 102.708 ; 
        RECT 55.696 98.334 55.8 102.708 ; 
        RECT 55.264 98.334 55.368 102.708 ; 
        RECT 54.832 98.334 54.936 102.708 ; 
        RECT 54.4 98.334 54.504 102.708 ; 
        RECT 53.968 98.334 54.072 102.708 ; 
        RECT 53.536 98.334 53.64 102.708 ; 
        RECT 53.104 98.334 53.208 102.708 ; 
        RECT 52.672 98.334 52.776 102.708 ; 
        RECT 52.24 98.334 52.344 102.708 ; 
        RECT 51.808 98.334 51.912 102.708 ; 
        RECT 51.376 98.334 51.48 102.708 ; 
        RECT 50.944 98.334 51.048 102.708 ; 
        RECT 50.512 98.334 50.616 102.708 ; 
        RECT 50.08 98.334 50.184 102.708 ; 
        RECT 49.648 98.334 49.752 102.708 ; 
        RECT 49.216 98.334 49.32 102.708 ; 
        RECT 48.784 98.334 48.888 102.708 ; 
        RECT 48.352 98.334 48.456 102.708 ; 
        RECT 47.92 98.334 48.024 102.708 ; 
        RECT 47.488 98.334 47.592 102.708 ; 
        RECT 47.056 98.334 47.16 102.708 ; 
        RECT 46.624 98.334 46.728 102.708 ; 
        RECT 46.192 98.334 46.296 102.708 ; 
        RECT 45.76 98.334 45.864 102.708 ; 
        RECT 45.328 98.334 45.432 102.708 ; 
        RECT 44.896 98.334 45 102.708 ; 
        RECT 44.464 98.334 44.568 102.708 ; 
        RECT 44.032 98.334 44.136 102.708 ; 
        RECT 43.6 98.334 43.704 102.708 ; 
        RECT 43.168 98.334 43.272 102.708 ; 
        RECT 42.736 98.334 42.84 102.708 ; 
        RECT 42.304 98.334 42.408 102.708 ; 
        RECT 41.872 98.334 41.976 102.708 ; 
        RECT 41.44 98.334 41.544 102.708 ; 
        RECT 41.008 98.334 41.112 102.708 ; 
        RECT 40.576 98.334 40.68 102.708 ; 
        RECT 40.144 98.334 40.248 102.708 ; 
        RECT 39.712 98.334 39.816 102.708 ; 
        RECT 39.28 98.334 39.384 102.708 ; 
        RECT 38.848 98.334 38.952 102.708 ; 
        RECT 38.416 98.334 38.52 102.708 ; 
        RECT 37.984 98.334 38.088 102.708 ; 
        RECT 37.552 98.334 37.656 102.708 ; 
        RECT 37.12 98.334 37.224 102.708 ; 
        RECT 36.688 98.334 36.792 102.708 ; 
        RECT 36.256 98.334 36.36 102.708 ; 
        RECT 35.824 98.334 35.928 102.708 ; 
        RECT 35.392 98.334 35.496 102.708 ; 
        RECT 34.96 98.334 35.064 102.708 ; 
        RECT 34.528 98.334 34.632 102.708 ; 
        RECT 34.096 98.334 34.2 102.708 ; 
        RECT 33.664 98.334 33.768 102.708 ; 
        RECT 33.232 98.334 33.336 102.708 ; 
        RECT 32.8 98.334 32.904 102.708 ; 
        RECT 32.368 98.334 32.472 102.708 ; 
        RECT 31.936 98.334 32.04 102.708 ; 
        RECT 31.504 98.334 31.608 102.708 ; 
        RECT 31.072 98.334 31.176 102.708 ; 
        RECT 30.64 98.334 30.744 102.708 ; 
        RECT 30.208 98.334 30.312 102.708 ; 
        RECT 29.776 98.334 29.88 102.708 ; 
        RECT 29.344 98.334 29.448 102.708 ; 
        RECT 28.912 98.334 29.016 102.708 ; 
        RECT 28.48 98.334 28.584 102.708 ; 
        RECT 28.048 98.334 28.152 102.708 ; 
        RECT 27.616 98.334 27.72 102.708 ; 
        RECT 27.184 98.334 27.288 102.708 ; 
        RECT 26.752 98.334 26.856 102.708 ; 
        RECT 26.32 98.334 26.424 102.708 ; 
        RECT 25.888 98.334 25.992 102.708 ; 
        RECT 25.456 98.334 25.56 102.708 ; 
        RECT 25.024 98.334 25.128 102.708 ; 
        RECT 24.592 98.334 24.696 102.708 ; 
        RECT 24.16 98.334 24.264 102.708 ; 
        RECT 23.728 98.334 23.832 102.708 ; 
        RECT 23.296 98.334 23.4 102.708 ; 
        RECT 22.864 98.334 22.968 102.708 ; 
        RECT 22.432 98.334 22.536 102.708 ; 
        RECT 22 98.334 22.104 102.708 ; 
        RECT 21.568 98.334 21.672 102.708 ; 
        RECT 21.136 98.334 21.24 102.708 ; 
        RECT 20.704 98.334 20.808 102.708 ; 
        RECT 20.272 98.334 20.376 102.708 ; 
        RECT 19.84 98.334 19.944 102.708 ; 
        RECT 19.408 98.334 19.512 102.708 ; 
        RECT 18.976 98.334 19.08 102.708 ; 
        RECT 18.544 98.334 18.648 102.708 ; 
        RECT 18.112 98.334 18.216 102.708 ; 
        RECT 17.68 98.334 17.784 102.708 ; 
        RECT 17.248 98.334 17.352 102.708 ; 
        RECT 16.816 98.334 16.92 102.708 ; 
        RECT 16.384 98.334 16.488 102.708 ; 
        RECT 15.952 98.334 16.056 102.708 ; 
        RECT 15.52 98.334 15.624 102.708 ; 
        RECT 15.088 98.334 15.192 102.708 ; 
        RECT 14.656 98.334 14.76 102.708 ; 
        RECT 14.224 98.334 14.328 102.708 ; 
        RECT 13.792 98.334 13.896 102.708 ; 
        RECT 13.36 98.334 13.464 102.708 ; 
        RECT 12.928 98.334 13.032 102.708 ; 
        RECT 12.496 98.334 12.6 102.708 ; 
        RECT 12.064 98.334 12.168 102.708 ; 
        RECT 11.632 98.334 11.736 102.708 ; 
        RECT 11.2 98.334 11.304 102.708 ; 
        RECT 10.768 98.334 10.872 102.708 ; 
        RECT 10.336 98.334 10.44 102.708 ; 
        RECT 9.904 98.334 10.008 102.708 ; 
        RECT 9.472 98.334 9.576 102.708 ; 
        RECT 9.04 98.334 9.144 102.708 ; 
        RECT 8.608 98.334 8.712 102.708 ; 
        RECT 8.176 98.334 8.28 102.708 ; 
        RECT 7.744 98.334 7.848 102.708 ; 
        RECT 7.312 98.334 7.416 102.708 ; 
        RECT 6.88 98.334 6.984 102.708 ; 
        RECT 6.448 98.334 6.552 102.708 ; 
        RECT 6.016 98.334 6.12 102.708 ; 
        RECT 5.584 98.334 5.688 102.708 ; 
        RECT 5.152 98.334 5.256 102.708 ; 
        RECT 4.72 98.334 4.824 102.708 ; 
        RECT 4.288 98.334 4.392 102.708 ; 
        RECT 3.856 98.334 3.96 102.708 ; 
        RECT 3.424 98.334 3.528 102.708 ; 
        RECT 2.992 98.334 3.096 102.708 ; 
        RECT 2.56 98.334 2.664 102.708 ; 
        RECT 2.128 98.334 2.232 102.708 ; 
        RECT 1.696 98.334 1.8 102.708 ; 
        RECT 1.264 98.334 1.368 102.708 ; 
        RECT 0.832 98.334 0.936 102.708 ; 
        RECT 0.02 98.334 0.36 102.708 ; 
        RECT 62.212 102.654 62.724 107.028 ; 
        RECT 62.156 105.316 62.724 106.606 ; 
        RECT 61.276 104.224 61.812 107.028 ; 
        RECT 61.184 105.564 61.812 106.596 ; 
        RECT 61.276 102.654 61.668 107.028 ; 
        RECT 61.276 103.138 61.724 104.096 ; 
        RECT 61.276 102.654 61.812 103.01 ; 
        RECT 60.376 104.456 60.912 107.028 ; 
        RECT 60.376 102.654 60.768 107.028 ; 
        RECT 58.708 102.654 59.04 107.028 ; 
        RECT 58.708 103.008 59.096 106.75 ; 
        RECT 121.072 102.654 121.412 107.028 ; 
        RECT 120.496 102.654 120.6 107.028 ; 
        RECT 120.064 102.654 120.168 107.028 ; 
        RECT 119.632 102.654 119.736 107.028 ; 
        RECT 119.2 102.654 119.304 107.028 ; 
        RECT 118.768 102.654 118.872 107.028 ; 
        RECT 118.336 102.654 118.44 107.028 ; 
        RECT 117.904 102.654 118.008 107.028 ; 
        RECT 117.472 102.654 117.576 107.028 ; 
        RECT 117.04 102.654 117.144 107.028 ; 
        RECT 116.608 102.654 116.712 107.028 ; 
        RECT 116.176 102.654 116.28 107.028 ; 
        RECT 115.744 102.654 115.848 107.028 ; 
        RECT 115.312 102.654 115.416 107.028 ; 
        RECT 114.88 102.654 114.984 107.028 ; 
        RECT 114.448 102.654 114.552 107.028 ; 
        RECT 114.016 102.654 114.12 107.028 ; 
        RECT 113.584 102.654 113.688 107.028 ; 
        RECT 113.152 102.654 113.256 107.028 ; 
        RECT 112.72 102.654 112.824 107.028 ; 
        RECT 112.288 102.654 112.392 107.028 ; 
        RECT 111.856 102.654 111.96 107.028 ; 
        RECT 111.424 102.654 111.528 107.028 ; 
        RECT 110.992 102.654 111.096 107.028 ; 
        RECT 110.56 102.654 110.664 107.028 ; 
        RECT 110.128 102.654 110.232 107.028 ; 
        RECT 109.696 102.654 109.8 107.028 ; 
        RECT 109.264 102.654 109.368 107.028 ; 
        RECT 108.832 102.654 108.936 107.028 ; 
        RECT 108.4 102.654 108.504 107.028 ; 
        RECT 107.968 102.654 108.072 107.028 ; 
        RECT 107.536 102.654 107.64 107.028 ; 
        RECT 107.104 102.654 107.208 107.028 ; 
        RECT 106.672 102.654 106.776 107.028 ; 
        RECT 106.24 102.654 106.344 107.028 ; 
        RECT 105.808 102.654 105.912 107.028 ; 
        RECT 105.376 102.654 105.48 107.028 ; 
        RECT 104.944 102.654 105.048 107.028 ; 
        RECT 104.512 102.654 104.616 107.028 ; 
        RECT 104.08 102.654 104.184 107.028 ; 
        RECT 103.648 102.654 103.752 107.028 ; 
        RECT 103.216 102.654 103.32 107.028 ; 
        RECT 102.784 102.654 102.888 107.028 ; 
        RECT 102.352 102.654 102.456 107.028 ; 
        RECT 101.92 102.654 102.024 107.028 ; 
        RECT 101.488 102.654 101.592 107.028 ; 
        RECT 101.056 102.654 101.16 107.028 ; 
        RECT 100.624 102.654 100.728 107.028 ; 
        RECT 100.192 102.654 100.296 107.028 ; 
        RECT 99.76 102.654 99.864 107.028 ; 
        RECT 99.328 102.654 99.432 107.028 ; 
        RECT 98.896 102.654 99 107.028 ; 
        RECT 98.464 102.654 98.568 107.028 ; 
        RECT 98.032 102.654 98.136 107.028 ; 
        RECT 97.6 102.654 97.704 107.028 ; 
        RECT 97.168 102.654 97.272 107.028 ; 
        RECT 96.736 102.654 96.84 107.028 ; 
        RECT 96.304 102.654 96.408 107.028 ; 
        RECT 95.872 102.654 95.976 107.028 ; 
        RECT 95.44 102.654 95.544 107.028 ; 
        RECT 95.008 102.654 95.112 107.028 ; 
        RECT 94.576 102.654 94.68 107.028 ; 
        RECT 94.144 102.654 94.248 107.028 ; 
        RECT 93.712 102.654 93.816 107.028 ; 
        RECT 93.28 102.654 93.384 107.028 ; 
        RECT 92.848 102.654 92.952 107.028 ; 
        RECT 92.416 102.654 92.52 107.028 ; 
        RECT 91.984 102.654 92.088 107.028 ; 
        RECT 91.552 102.654 91.656 107.028 ; 
        RECT 91.12 102.654 91.224 107.028 ; 
        RECT 90.688 102.654 90.792 107.028 ; 
        RECT 90.256 102.654 90.36 107.028 ; 
        RECT 89.824 102.654 89.928 107.028 ; 
        RECT 89.392 102.654 89.496 107.028 ; 
        RECT 88.96 102.654 89.064 107.028 ; 
        RECT 88.528 102.654 88.632 107.028 ; 
        RECT 88.096 102.654 88.2 107.028 ; 
        RECT 87.664 102.654 87.768 107.028 ; 
        RECT 87.232 102.654 87.336 107.028 ; 
        RECT 86.8 102.654 86.904 107.028 ; 
        RECT 86.368 102.654 86.472 107.028 ; 
        RECT 85.936 102.654 86.04 107.028 ; 
        RECT 85.504 102.654 85.608 107.028 ; 
        RECT 85.072 102.654 85.176 107.028 ; 
        RECT 84.64 102.654 84.744 107.028 ; 
        RECT 84.208 102.654 84.312 107.028 ; 
        RECT 83.776 102.654 83.88 107.028 ; 
        RECT 83.344 102.654 83.448 107.028 ; 
        RECT 82.912 102.654 83.016 107.028 ; 
        RECT 82.48 102.654 82.584 107.028 ; 
        RECT 82.048 102.654 82.152 107.028 ; 
        RECT 81.616 102.654 81.72 107.028 ; 
        RECT 81.184 102.654 81.288 107.028 ; 
        RECT 80.752 102.654 80.856 107.028 ; 
        RECT 80.32 102.654 80.424 107.028 ; 
        RECT 79.888 102.654 79.992 107.028 ; 
        RECT 79.456 102.654 79.56 107.028 ; 
        RECT 79.024 102.654 79.128 107.028 ; 
        RECT 78.592 102.654 78.696 107.028 ; 
        RECT 78.16 102.654 78.264 107.028 ; 
        RECT 77.728 102.654 77.832 107.028 ; 
        RECT 77.296 102.654 77.4 107.028 ; 
        RECT 76.864 102.654 76.968 107.028 ; 
        RECT 76.432 102.654 76.536 107.028 ; 
        RECT 76 102.654 76.104 107.028 ; 
        RECT 75.568 102.654 75.672 107.028 ; 
        RECT 75.136 102.654 75.24 107.028 ; 
        RECT 74.704 102.654 74.808 107.028 ; 
        RECT 74.272 102.654 74.376 107.028 ; 
        RECT 73.84 102.654 73.944 107.028 ; 
        RECT 73.408 102.654 73.512 107.028 ; 
        RECT 72.976 102.654 73.08 107.028 ; 
        RECT 72.544 102.654 72.648 107.028 ; 
        RECT 72.112 102.654 72.216 107.028 ; 
        RECT 71.68 102.654 71.784 107.028 ; 
        RECT 71.248 102.654 71.352 107.028 ; 
        RECT 70.816 102.654 70.92 107.028 ; 
        RECT 70.384 102.654 70.488 107.028 ; 
        RECT 69.952 102.654 70.056 107.028 ; 
        RECT 69.52 102.654 69.624 107.028 ; 
        RECT 69.088 102.654 69.192 107.028 ; 
        RECT 68.656 102.654 68.76 107.028 ; 
        RECT 68.224 102.654 68.328 107.028 ; 
        RECT 67.792 102.654 67.896 107.028 ; 
        RECT 67.36 102.654 67.464 107.028 ; 
        RECT 66.928 102.654 67.032 107.028 ; 
        RECT 66.496 102.654 66.6 107.028 ; 
        RECT 66.064 102.654 66.168 107.028 ; 
        RECT 65.632 102.654 65.736 107.028 ; 
        RECT 65.2 102.654 65.304 107.028 ; 
        RECT 64.348 102.654 64.656 107.028 ; 
        RECT 56.776 102.654 57.084 107.028 ; 
        RECT 56.128 102.654 56.232 107.028 ; 
        RECT 55.696 102.654 55.8 107.028 ; 
        RECT 55.264 102.654 55.368 107.028 ; 
        RECT 54.832 102.654 54.936 107.028 ; 
        RECT 54.4 102.654 54.504 107.028 ; 
        RECT 53.968 102.654 54.072 107.028 ; 
        RECT 53.536 102.654 53.64 107.028 ; 
        RECT 53.104 102.654 53.208 107.028 ; 
        RECT 52.672 102.654 52.776 107.028 ; 
        RECT 52.24 102.654 52.344 107.028 ; 
        RECT 51.808 102.654 51.912 107.028 ; 
        RECT 51.376 102.654 51.48 107.028 ; 
        RECT 50.944 102.654 51.048 107.028 ; 
        RECT 50.512 102.654 50.616 107.028 ; 
        RECT 50.08 102.654 50.184 107.028 ; 
        RECT 49.648 102.654 49.752 107.028 ; 
        RECT 49.216 102.654 49.32 107.028 ; 
        RECT 48.784 102.654 48.888 107.028 ; 
        RECT 48.352 102.654 48.456 107.028 ; 
        RECT 47.92 102.654 48.024 107.028 ; 
        RECT 47.488 102.654 47.592 107.028 ; 
        RECT 47.056 102.654 47.16 107.028 ; 
        RECT 46.624 102.654 46.728 107.028 ; 
        RECT 46.192 102.654 46.296 107.028 ; 
        RECT 45.76 102.654 45.864 107.028 ; 
        RECT 45.328 102.654 45.432 107.028 ; 
        RECT 44.896 102.654 45 107.028 ; 
        RECT 44.464 102.654 44.568 107.028 ; 
        RECT 44.032 102.654 44.136 107.028 ; 
        RECT 43.6 102.654 43.704 107.028 ; 
        RECT 43.168 102.654 43.272 107.028 ; 
        RECT 42.736 102.654 42.84 107.028 ; 
        RECT 42.304 102.654 42.408 107.028 ; 
        RECT 41.872 102.654 41.976 107.028 ; 
        RECT 41.44 102.654 41.544 107.028 ; 
        RECT 41.008 102.654 41.112 107.028 ; 
        RECT 40.576 102.654 40.68 107.028 ; 
        RECT 40.144 102.654 40.248 107.028 ; 
        RECT 39.712 102.654 39.816 107.028 ; 
        RECT 39.28 102.654 39.384 107.028 ; 
        RECT 38.848 102.654 38.952 107.028 ; 
        RECT 38.416 102.654 38.52 107.028 ; 
        RECT 37.984 102.654 38.088 107.028 ; 
        RECT 37.552 102.654 37.656 107.028 ; 
        RECT 37.12 102.654 37.224 107.028 ; 
        RECT 36.688 102.654 36.792 107.028 ; 
        RECT 36.256 102.654 36.36 107.028 ; 
        RECT 35.824 102.654 35.928 107.028 ; 
        RECT 35.392 102.654 35.496 107.028 ; 
        RECT 34.96 102.654 35.064 107.028 ; 
        RECT 34.528 102.654 34.632 107.028 ; 
        RECT 34.096 102.654 34.2 107.028 ; 
        RECT 33.664 102.654 33.768 107.028 ; 
        RECT 33.232 102.654 33.336 107.028 ; 
        RECT 32.8 102.654 32.904 107.028 ; 
        RECT 32.368 102.654 32.472 107.028 ; 
        RECT 31.936 102.654 32.04 107.028 ; 
        RECT 31.504 102.654 31.608 107.028 ; 
        RECT 31.072 102.654 31.176 107.028 ; 
        RECT 30.64 102.654 30.744 107.028 ; 
        RECT 30.208 102.654 30.312 107.028 ; 
        RECT 29.776 102.654 29.88 107.028 ; 
        RECT 29.344 102.654 29.448 107.028 ; 
        RECT 28.912 102.654 29.016 107.028 ; 
        RECT 28.48 102.654 28.584 107.028 ; 
        RECT 28.048 102.654 28.152 107.028 ; 
        RECT 27.616 102.654 27.72 107.028 ; 
        RECT 27.184 102.654 27.288 107.028 ; 
        RECT 26.752 102.654 26.856 107.028 ; 
        RECT 26.32 102.654 26.424 107.028 ; 
        RECT 25.888 102.654 25.992 107.028 ; 
        RECT 25.456 102.654 25.56 107.028 ; 
        RECT 25.024 102.654 25.128 107.028 ; 
        RECT 24.592 102.654 24.696 107.028 ; 
        RECT 24.16 102.654 24.264 107.028 ; 
        RECT 23.728 102.654 23.832 107.028 ; 
        RECT 23.296 102.654 23.4 107.028 ; 
        RECT 22.864 102.654 22.968 107.028 ; 
        RECT 22.432 102.654 22.536 107.028 ; 
        RECT 22 102.654 22.104 107.028 ; 
        RECT 21.568 102.654 21.672 107.028 ; 
        RECT 21.136 102.654 21.24 107.028 ; 
        RECT 20.704 102.654 20.808 107.028 ; 
        RECT 20.272 102.654 20.376 107.028 ; 
        RECT 19.84 102.654 19.944 107.028 ; 
        RECT 19.408 102.654 19.512 107.028 ; 
        RECT 18.976 102.654 19.08 107.028 ; 
        RECT 18.544 102.654 18.648 107.028 ; 
        RECT 18.112 102.654 18.216 107.028 ; 
        RECT 17.68 102.654 17.784 107.028 ; 
        RECT 17.248 102.654 17.352 107.028 ; 
        RECT 16.816 102.654 16.92 107.028 ; 
        RECT 16.384 102.654 16.488 107.028 ; 
        RECT 15.952 102.654 16.056 107.028 ; 
        RECT 15.52 102.654 15.624 107.028 ; 
        RECT 15.088 102.654 15.192 107.028 ; 
        RECT 14.656 102.654 14.76 107.028 ; 
        RECT 14.224 102.654 14.328 107.028 ; 
        RECT 13.792 102.654 13.896 107.028 ; 
        RECT 13.36 102.654 13.464 107.028 ; 
        RECT 12.928 102.654 13.032 107.028 ; 
        RECT 12.496 102.654 12.6 107.028 ; 
        RECT 12.064 102.654 12.168 107.028 ; 
        RECT 11.632 102.654 11.736 107.028 ; 
        RECT 11.2 102.654 11.304 107.028 ; 
        RECT 10.768 102.654 10.872 107.028 ; 
        RECT 10.336 102.654 10.44 107.028 ; 
        RECT 9.904 102.654 10.008 107.028 ; 
        RECT 9.472 102.654 9.576 107.028 ; 
        RECT 9.04 102.654 9.144 107.028 ; 
        RECT 8.608 102.654 8.712 107.028 ; 
        RECT 8.176 102.654 8.28 107.028 ; 
        RECT 7.744 102.654 7.848 107.028 ; 
        RECT 7.312 102.654 7.416 107.028 ; 
        RECT 6.88 102.654 6.984 107.028 ; 
        RECT 6.448 102.654 6.552 107.028 ; 
        RECT 6.016 102.654 6.12 107.028 ; 
        RECT 5.584 102.654 5.688 107.028 ; 
        RECT 5.152 102.654 5.256 107.028 ; 
        RECT 4.72 102.654 4.824 107.028 ; 
        RECT 4.288 102.654 4.392 107.028 ; 
        RECT 3.856 102.654 3.96 107.028 ; 
        RECT 3.424 102.654 3.528 107.028 ; 
        RECT 2.992 102.654 3.096 107.028 ; 
        RECT 2.56 102.654 2.664 107.028 ; 
        RECT 2.128 102.654 2.232 107.028 ; 
        RECT 1.696 102.654 1.8 107.028 ; 
        RECT 1.264 102.654 1.368 107.028 ; 
        RECT 0.832 102.654 0.936 107.028 ; 
        RECT 0.02 102.654 0.36 107.028 ; 
        RECT 62.212 106.974 62.724 111.348 ; 
        RECT 62.156 109.636 62.724 110.926 ; 
        RECT 61.276 108.544 61.812 111.348 ; 
        RECT 61.184 109.884 61.812 110.916 ; 
        RECT 61.276 106.974 61.668 111.348 ; 
        RECT 61.276 107.458 61.724 108.416 ; 
        RECT 61.276 106.974 61.812 107.33 ; 
        RECT 60.376 108.776 60.912 111.348 ; 
        RECT 60.376 106.974 60.768 111.348 ; 
        RECT 58.708 106.974 59.04 111.348 ; 
        RECT 58.708 107.328 59.096 111.07 ; 
        RECT 121.072 106.974 121.412 111.348 ; 
        RECT 120.496 106.974 120.6 111.348 ; 
        RECT 120.064 106.974 120.168 111.348 ; 
        RECT 119.632 106.974 119.736 111.348 ; 
        RECT 119.2 106.974 119.304 111.348 ; 
        RECT 118.768 106.974 118.872 111.348 ; 
        RECT 118.336 106.974 118.44 111.348 ; 
        RECT 117.904 106.974 118.008 111.348 ; 
        RECT 117.472 106.974 117.576 111.348 ; 
        RECT 117.04 106.974 117.144 111.348 ; 
        RECT 116.608 106.974 116.712 111.348 ; 
        RECT 116.176 106.974 116.28 111.348 ; 
        RECT 115.744 106.974 115.848 111.348 ; 
        RECT 115.312 106.974 115.416 111.348 ; 
        RECT 114.88 106.974 114.984 111.348 ; 
        RECT 114.448 106.974 114.552 111.348 ; 
        RECT 114.016 106.974 114.12 111.348 ; 
        RECT 113.584 106.974 113.688 111.348 ; 
        RECT 113.152 106.974 113.256 111.348 ; 
        RECT 112.72 106.974 112.824 111.348 ; 
        RECT 112.288 106.974 112.392 111.348 ; 
        RECT 111.856 106.974 111.96 111.348 ; 
        RECT 111.424 106.974 111.528 111.348 ; 
        RECT 110.992 106.974 111.096 111.348 ; 
        RECT 110.56 106.974 110.664 111.348 ; 
        RECT 110.128 106.974 110.232 111.348 ; 
        RECT 109.696 106.974 109.8 111.348 ; 
        RECT 109.264 106.974 109.368 111.348 ; 
        RECT 108.832 106.974 108.936 111.348 ; 
        RECT 108.4 106.974 108.504 111.348 ; 
        RECT 107.968 106.974 108.072 111.348 ; 
        RECT 107.536 106.974 107.64 111.348 ; 
        RECT 107.104 106.974 107.208 111.348 ; 
        RECT 106.672 106.974 106.776 111.348 ; 
        RECT 106.24 106.974 106.344 111.348 ; 
        RECT 105.808 106.974 105.912 111.348 ; 
        RECT 105.376 106.974 105.48 111.348 ; 
        RECT 104.944 106.974 105.048 111.348 ; 
        RECT 104.512 106.974 104.616 111.348 ; 
        RECT 104.08 106.974 104.184 111.348 ; 
        RECT 103.648 106.974 103.752 111.348 ; 
        RECT 103.216 106.974 103.32 111.348 ; 
        RECT 102.784 106.974 102.888 111.348 ; 
        RECT 102.352 106.974 102.456 111.348 ; 
        RECT 101.92 106.974 102.024 111.348 ; 
        RECT 101.488 106.974 101.592 111.348 ; 
        RECT 101.056 106.974 101.16 111.348 ; 
        RECT 100.624 106.974 100.728 111.348 ; 
        RECT 100.192 106.974 100.296 111.348 ; 
        RECT 99.76 106.974 99.864 111.348 ; 
        RECT 99.328 106.974 99.432 111.348 ; 
        RECT 98.896 106.974 99 111.348 ; 
        RECT 98.464 106.974 98.568 111.348 ; 
        RECT 98.032 106.974 98.136 111.348 ; 
        RECT 97.6 106.974 97.704 111.348 ; 
        RECT 97.168 106.974 97.272 111.348 ; 
        RECT 96.736 106.974 96.84 111.348 ; 
        RECT 96.304 106.974 96.408 111.348 ; 
        RECT 95.872 106.974 95.976 111.348 ; 
        RECT 95.44 106.974 95.544 111.348 ; 
        RECT 95.008 106.974 95.112 111.348 ; 
        RECT 94.576 106.974 94.68 111.348 ; 
        RECT 94.144 106.974 94.248 111.348 ; 
        RECT 93.712 106.974 93.816 111.348 ; 
        RECT 93.28 106.974 93.384 111.348 ; 
        RECT 92.848 106.974 92.952 111.348 ; 
        RECT 92.416 106.974 92.52 111.348 ; 
        RECT 91.984 106.974 92.088 111.348 ; 
        RECT 91.552 106.974 91.656 111.348 ; 
        RECT 91.12 106.974 91.224 111.348 ; 
        RECT 90.688 106.974 90.792 111.348 ; 
        RECT 90.256 106.974 90.36 111.348 ; 
        RECT 89.824 106.974 89.928 111.348 ; 
        RECT 89.392 106.974 89.496 111.348 ; 
        RECT 88.96 106.974 89.064 111.348 ; 
        RECT 88.528 106.974 88.632 111.348 ; 
        RECT 88.096 106.974 88.2 111.348 ; 
        RECT 87.664 106.974 87.768 111.348 ; 
        RECT 87.232 106.974 87.336 111.348 ; 
        RECT 86.8 106.974 86.904 111.348 ; 
        RECT 86.368 106.974 86.472 111.348 ; 
        RECT 85.936 106.974 86.04 111.348 ; 
        RECT 85.504 106.974 85.608 111.348 ; 
        RECT 85.072 106.974 85.176 111.348 ; 
        RECT 84.64 106.974 84.744 111.348 ; 
        RECT 84.208 106.974 84.312 111.348 ; 
        RECT 83.776 106.974 83.88 111.348 ; 
        RECT 83.344 106.974 83.448 111.348 ; 
        RECT 82.912 106.974 83.016 111.348 ; 
        RECT 82.48 106.974 82.584 111.348 ; 
        RECT 82.048 106.974 82.152 111.348 ; 
        RECT 81.616 106.974 81.72 111.348 ; 
        RECT 81.184 106.974 81.288 111.348 ; 
        RECT 80.752 106.974 80.856 111.348 ; 
        RECT 80.32 106.974 80.424 111.348 ; 
        RECT 79.888 106.974 79.992 111.348 ; 
        RECT 79.456 106.974 79.56 111.348 ; 
        RECT 79.024 106.974 79.128 111.348 ; 
        RECT 78.592 106.974 78.696 111.348 ; 
        RECT 78.16 106.974 78.264 111.348 ; 
        RECT 77.728 106.974 77.832 111.348 ; 
        RECT 77.296 106.974 77.4 111.348 ; 
        RECT 76.864 106.974 76.968 111.348 ; 
        RECT 76.432 106.974 76.536 111.348 ; 
        RECT 76 106.974 76.104 111.348 ; 
        RECT 75.568 106.974 75.672 111.348 ; 
        RECT 75.136 106.974 75.24 111.348 ; 
        RECT 74.704 106.974 74.808 111.348 ; 
        RECT 74.272 106.974 74.376 111.348 ; 
        RECT 73.84 106.974 73.944 111.348 ; 
        RECT 73.408 106.974 73.512 111.348 ; 
        RECT 72.976 106.974 73.08 111.348 ; 
        RECT 72.544 106.974 72.648 111.348 ; 
        RECT 72.112 106.974 72.216 111.348 ; 
        RECT 71.68 106.974 71.784 111.348 ; 
        RECT 71.248 106.974 71.352 111.348 ; 
        RECT 70.816 106.974 70.92 111.348 ; 
        RECT 70.384 106.974 70.488 111.348 ; 
        RECT 69.952 106.974 70.056 111.348 ; 
        RECT 69.52 106.974 69.624 111.348 ; 
        RECT 69.088 106.974 69.192 111.348 ; 
        RECT 68.656 106.974 68.76 111.348 ; 
        RECT 68.224 106.974 68.328 111.348 ; 
        RECT 67.792 106.974 67.896 111.348 ; 
        RECT 67.36 106.974 67.464 111.348 ; 
        RECT 66.928 106.974 67.032 111.348 ; 
        RECT 66.496 106.974 66.6 111.348 ; 
        RECT 66.064 106.974 66.168 111.348 ; 
        RECT 65.632 106.974 65.736 111.348 ; 
        RECT 65.2 106.974 65.304 111.348 ; 
        RECT 64.348 106.974 64.656 111.348 ; 
        RECT 56.776 106.974 57.084 111.348 ; 
        RECT 56.128 106.974 56.232 111.348 ; 
        RECT 55.696 106.974 55.8 111.348 ; 
        RECT 55.264 106.974 55.368 111.348 ; 
        RECT 54.832 106.974 54.936 111.348 ; 
        RECT 54.4 106.974 54.504 111.348 ; 
        RECT 53.968 106.974 54.072 111.348 ; 
        RECT 53.536 106.974 53.64 111.348 ; 
        RECT 53.104 106.974 53.208 111.348 ; 
        RECT 52.672 106.974 52.776 111.348 ; 
        RECT 52.24 106.974 52.344 111.348 ; 
        RECT 51.808 106.974 51.912 111.348 ; 
        RECT 51.376 106.974 51.48 111.348 ; 
        RECT 50.944 106.974 51.048 111.348 ; 
        RECT 50.512 106.974 50.616 111.348 ; 
        RECT 50.08 106.974 50.184 111.348 ; 
        RECT 49.648 106.974 49.752 111.348 ; 
        RECT 49.216 106.974 49.32 111.348 ; 
        RECT 48.784 106.974 48.888 111.348 ; 
        RECT 48.352 106.974 48.456 111.348 ; 
        RECT 47.92 106.974 48.024 111.348 ; 
        RECT 47.488 106.974 47.592 111.348 ; 
        RECT 47.056 106.974 47.16 111.348 ; 
        RECT 46.624 106.974 46.728 111.348 ; 
        RECT 46.192 106.974 46.296 111.348 ; 
        RECT 45.76 106.974 45.864 111.348 ; 
        RECT 45.328 106.974 45.432 111.348 ; 
        RECT 44.896 106.974 45 111.348 ; 
        RECT 44.464 106.974 44.568 111.348 ; 
        RECT 44.032 106.974 44.136 111.348 ; 
        RECT 43.6 106.974 43.704 111.348 ; 
        RECT 43.168 106.974 43.272 111.348 ; 
        RECT 42.736 106.974 42.84 111.348 ; 
        RECT 42.304 106.974 42.408 111.348 ; 
        RECT 41.872 106.974 41.976 111.348 ; 
        RECT 41.44 106.974 41.544 111.348 ; 
        RECT 41.008 106.974 41.112 111.348 ; 
        RECT 40.576 106.974 40.68 111.348 ; 
        RECT 40.144 106.974 40.248 111.348 ; 
        RECT 39.712 106.974 39.816 111.348 ; 
        RECT 39.28 106.974 39.384 111.348 ; 
        RECT 38.848 106.974 38.952 111.348 ; 
        RECT 38.416 106.974 38.52 111.348 ; 
        RECT 37.984 106.974 38.088 111.348 ; 
        RECT 37.552 106.974 37.656 111.348 ; 
        RECT 37.12 106.974 37.224 111.348 ; 
        RECT 36.688 106.974 36.792 111.348 ; 
        RECT 36.256 106.974 36.36 111.348 ; 
        RECT 35.824 106.974 35.928 111.348 ; 
        RECT 35.392 106.974 35.496 111.348 ; 
        RECT 34.96 106.974 35.064 111.348 ; 
        RECT 34.528 106.974 34.632 111.348 ; 
        RECT 34.096 106.974 34.2 111.348 ; 
        RECT 33.664 106.974 33.768 111.348 ; 
        RECT 33.232 106.974 33.336 111.348 ; 
        RECT 32.8 106.974 32.904 111.348 ; 
        RECT 32.368 106.974 32.472 111.348 ; 
        RECT 31.936 106.974 32.04 111.348 ; 
        RECT 31.504 106.974 31.608 111.348 ; 
        RECT 31.072 106.974 31.176 111.348 ; 
        RECT 30.64 106.974 30.744 111.348 ; 
        RECT 30.208 106.974 30.312 111.348 ; 
        RECT 29.776 106.974 29.88 111.348 ; 
        RECT 29.344 106.974 29.448 111.348 ; 
        RECT 28.912 106.974 29.016 111.348 ; 
        RECT 28.48 106.974 28.584 111.348 ; 
        RECT 28.048 106.974 28.152 111.348 ; 
        RECT 27.616 106.974 27.72 111.348 ; 
        RECT 27.184 106.974 27.288 111.348 ; 
        RECT 26.752 106.974 26.856 111.348 ; 
        RECT 26.32 106.974 26.424 111.348 ; 
        RECT 25.888 106.974 25.992 111.348 ; 
        RECT 25.456 106.974 25.56 111.348 ; 
        RECT 25.024 106.974 25.128 111.348 ; 
        RECT 24.592 106.974 24.696 111.348 ; 
        RECT 24.16 106.974 24.264 111.348 ; 
        RECT 23.728 106.974 23.832 111.348 ; 
        RECT 23.296 106.974 23.4 111.348 ; 
        RECT 22.864 106.974 22.968 111.348 ; 
        RECT 22.432 106.974 22.536 111.348 ; 
        RECT 22 106.974 22.104 111.348 ; 
        RECT 21.568 106.974 21.672 111.348 ; 
        RECT 21.136 106.974 21.24 111.348 ; 
        RECT 20.704 106.974 20.808 111.348 ; 
        RECT 20.272 106.974 20.376 111.348 ; 
        RECT 19.84 106.974 19.944 111.348 ; 
        RECT 19.408 106.974 19.512 111.348 ; 
        RECT 18.976 106.974 19.08 111.348 ; 
        RECT 18.544 106.974 18.648 111.348 ; 
        RECT 18.112 106.974 18.216 111.348 ; 
        RECT 17.68 106.974 17.784 111.348 ; 
        RECT 17.248 106.974 17.352 111.348 ; 
        RECT 16.816 106.974 16.92 111.348 ; 
        RECT 16.384 106.974 16.488 111.348 ; 
        RECT 15.952 106.974 16.056 111.348 ; 
        RECT 15.52 106.974 15.624 111.348 ; 
        RECT 15.088 106.974 15.192 111.348 ; 
        RECT 14.656 106.974 14.76 111.348 ; 
        RECT 14.224 106.974 14.328 111.348 ; 
        RECT 13.792 106.974 13.896 111.348 ; 
        RECT 13.36 106.974 13.464 111.348 ; 
        RECT 12.928 106.974 13.032 111.348 ; 
        RECT 12.496 106.974 12.6 111.348 ; 
        RECT 12.064 106.974 12.168 111.348 ; 
        RECT 11.632 106.974 11.736 111.348 ; 
        RECT 11.2 106.974 11.304 111.348 ; 
        RECT 10.768 106.974 10.872 111.348 ; 
        RECT 10.336 106.974 10.44 111.348 ; 
        RECT 9.904 106.974 10.008 111.348 ; 
        RECT 9.472 106.974 9.576 111.348 ; 
        RECT 9.04 106.974 9.144 111.348 ; 
        RECT 8.608 106.974 8.712 111.348 ; 
        RECT 8.176 106.974 8.28 111.348 ; 
        RECT 7.744 106.974 7.848 111.348 ; 
        RECT 7.312 106.974 7.416 111.348 ; 
        RECT 6.88 106.974 6.984 111.348 ; 
        RECT 6.448 106.974 6.552 111.348 ; 
        RECT 6.016 106.974 6.12 111.348 ; 
        RECT 5.584 106.974 5.688 111.348 ; 
        RECT 5.152 106.974 5.256 111.348 ; 
        RECT 4.72 106.974 4.824 111.348 ; 
        RECT 4.288 106.974 4.392 111.348 ; 
        RECT 3.856 106.974 3.96 111.348 ; 
        RECT 3.424 106.974 3.528 111.348 ; 
        RECT 2.992 106.974 3.096 111.348 ; 
        RECT 2.56 106.974 2.664 111.348 ; 
        RECT 2.128 106.974 2.232 111.348 ; 
        RECT 1.696 106.974 1.8 111.348 ; 
        RECT 1.264 106.974 1.368 111.348 ; 
        RECT 0.832 106.974 0.936 111.348 ; 
        RECT 0.02 106.974 0.36 111.348 ; 
  LAYER V3 SPACING 0.072 ; 
      RECT 0.02 4.88 121.412 5.4 ; 
      RECT 120.944 1.026 121.412 5.4 ; 
      RECT 64.856 4.496 120.872 5.4 ; 
      RECT 59.528 4.496 64.784 5.4 ; 
      RECT 56.648 1.026 59.168 5.4 ; 
      RECT 0.56 4.496 56.576 5.4 ; 
      RECT 0.02 1.026 0.488 5.4 ; 
      RECT 120.8 1.026 121.412 4.688 ; 
      RECT 65.072 1.026 120.728 5.4 ; 
      RECT 62.084 1.026 65 4.688 ; 
      RECT 61.148 1.808 61.94 5.4 ; 
      RECT 56.432 1.424 61.04 4.688 ; 
      RECT 0.704 1.026 56.36 5.4 ; 
      RECT 0.02 1.026 0.632 4.688 ; 
      RECT 61.868 1.026 121.412 4.304 ; 
      RECT 0.02 1.424 61.796 4.304 ; 
      RECT 60.968 1.026 121.412 1.712 ; 
      RECT 0.02 1.026 60.896 4.304 ; 
      RECT 0.02 1.026 121.412 1.328 ; 
      RECT 0.02 9.2 121.412 9.72 ; 
      RECT 120.944 5.346 121.412 9.72 ; 
      RECT 64.856 8.816 120.872 9.72 ; 
      RECT 59.528 8.816 64.784 9.72 ; 
      RECT 56.648 5.346 59.168 9.72 ; 
      RECT 0.56 8.816 56.576 9.72 ; 
      RECT 0.02 5.346 0.488 9.72 ; 
      RECT 120.8 5.346 121.412 9.008 ; 
      RECT 65.072 5.346 120.728 9.72 ; 
      RECT 62.084 5.346 65 9.008 ; 
      RECT 61.148 6.128 61.94 9.72 ; 
      RECT 56.432 5.744 61.04 9.008 ; 
      RECT 0.704 5.346 56.36 9.72 ; 
      RECT 0.02 5.346 0.632 9.008 ; 
      RECT 61.868 5.346 121.412 8.624 ; 
      RECT 0.02 5.744 61.796 8.624 ; 
      RECT 60.968 5.346 121.412 6.032 ; 
      RECT 0.02 5.346 60.896 8.624 ; 
      RECT 0.02 5.346 121.412 5.648 ; 
      RECT 0.02 13.52 121.412 14.04 ; 
      RECT 120.944 9.666 121.412 14.04 ; 
      RECT 64.856 13.136 120.872 14.04 ; 
      RECT 59.528 13.136 64.784 14.04 ; 
      RECT 56.648 9.666 59.168 14.04 ; 
      RECT 0.56 13.136 56.576 14.04 ; 
      RECT 0.02 9.666 0.488 14.04 ; 
      RECT 120.8 9.666 121.412 13.328 ; 
      RECT 65.072 9.666 120.728 14.04 ; 
      RECT 62.084 9.666 65 13.328 ; 
      RECT 61.148 10.448 61.94 14.04 ; 
      RECT 56.432 10.064 61.04 13.328 ; 
      RECT 0.704 9.666 56.36 14.04 ; 
      RECT 0.02 9.666 0.632 13.328 ; 
      RECT 61.868 9.666 121.412 12.944 ; 
      RECT 0.02 10.064 61.796 12.944 ; 
      RECT 60.968 9.666 121.412 10.352 ; 
      RECT 0.02 9.666 60.896 12.944 ; 
      RECT 0.02 9.666 121.412 9.968 ; 
      RECT 0.02 17.84 121.412 18.36 ; 
      RECT 120.944 13.986 121.412 18.36 ; 
      RECT 64.856 17.456 120.872 18.36 ; 
      RECT 59.528 17.456 64.784 18.36 ; 
      RECT 56.648 13.986 59.168 18.36 ; 
      RECT 0.56 17.456 56.576 18.36 ; 
      RECT 0.02 13.986 0.488 18.36 ; 
      RECT 120.8 13.986 121.412 17.648 ; 
      RECT 65.072 13.986 120.728 18.36 ; 
      RECT 62.084 13.986 65 17.648 ; 
      RECT 61.148 14.768 61.94 18.36 ; 
      RECT 56.432 14.384 61.04 17.648 ; 
      RECT 0.704 13.986 56.36 18.36 ; 
      RECT 0.02 13.986 0.632 17.648 ; 
      RECT 61.868 13.986 121.412 17.264 ; 
      RECT 0.02 14.384 61.796 17.264 ; 
      RECT 60.968 13.986 121.412 14.672 ; 
      RECT 0.02 13.986 60.896 17.264 ; 
      RECT 0.02 13.986 121.412 14.288 ; 
      RECT 0.02 22.16 121.412 22.68 ; 
      RECT 120.944 18.306 121.412 22.68 ; 
      RECT 64.856 21.776 120.872 22.68 ; 
      RECT 59.528 21.776 64.784 22.68 ; 
      RECT 56.648 18.306 59.168 22.68 ; 
      RECT 0.56 21.776 56.576 22.68 ; 
      RECT 0.02 18.306 0.488 22.68 ; 
      RECT 120.8 18.306 121.412 21.968 ; 
      RECT 65.072 18.306 120.728 22.68 ; 
      RECT 62.084 18.306 65 21.968 ; 
      RECT 61.148 19.088 61.94 22.68 ; 
      RECT 56.432 18.704 61.04 21.968 ; 
      RECT 0.704 18.306 56.36 22.68 ; 
      RECT 0.02 18.306 0.632 21.968 ; 
      RECT 61.868 18.306 121.412 21.584 ; 
      RECT 0.02 18.704 61.796 21.584 ; 
      RECT 60.968 18.306 121.412 18.992 ; 
      RECT 0.02 18.306 60.896 21.584 ; 
      RECT 0.02 18.306 121.412 18.608 ; 
      RECT 0.02 26.48 121.412 27 ; 
      RECT 120.944 22.626 121.412 27 ; 
      RECT 64.856 26.096 120.872 27 ; 
      RECT 59.528 26.096 64.784 27 ; 
      RECT 56.648 22.626 59.168 27 ; 
      RECT 0.56 26.096 56.576 27 ; 
      RECT 0.02 22.626 0.488 27 ; 
      RECT 120.8 22.626 121.412 26.288 ; 
      RECT 65.072 22.626 120.728 27 ; 
      RECT 62.084 22.626 65 26.288 ; 
      RECT 61.148 23.408 61.94 27 ; 
      RECT 56.432 23.024 61.04 26.288 ; 
      RECT 0.704 22.626 56.36 27 ; 
      RECT 0.02 22.626 0.632 26.288 ; 
      RECT 61.868 22.626 121.412 25.904 ; 
      RECT 0.02 23.024 61.796 25.904 ; 
      RECT 60.968 22.626 121.412 23.312 ; 
      RECT 0.02 22.626 60.896 25.904 ; 
      RECT 0.02 22.626 121.412 22.928 ; 
      RECT 0.02 30.8 121.412 31.32 ; 
      RECT 120.944 26.946 121.412 31.32 ; 
      RECT 64.856 30.416 120.872 31.32 ; 
      RECT 59.528 30.416 64.784 31.32 ; 
      RECT 56.648 26.946 59.168 31.32 ; 
      RECT 0.56 30.416 56.576 31.32 ; 
      RECT 0.02 26.946 0.488 31.32 ; 
      RECT 120.8 26.946 121.412 30.608 ; 
      RECT 65.072 26.946 120.728 31.32 ; 
      RECT 62.084 26.946 65 30.608 ; 
      RECT 61.148 27.728 61.94 31.32 ; 
      RECT 56.432 27.344 61.04 30.608 ; 
      RECT 0.704 26.946 56.36 31.32 ; 
      RECT 0.02 26.946 0.632 30.608 ; 
      RECT 61.868 26.946 121.412 30.224 ; 
      RECT 0.02 27.344 61.796 30.224 ; 
      RECT 60.968 26.946 121.412 27.632 ; 
      RECT 0.02 26.946 60.896 30.224 ; 
      RECT 0.02 26.946 121.412 27.248 ; 
      RECT 0.02 35.12 121.412 35.64 ; 
      RECT 120.944 31.266 121.412 35.64 ; 
      RECT 64.856 34.736 120.872 35.64 ; 
      RECT 59.528 34.736 64.784 35.64 ; 
      RECT 56.648 31.266 59.168 35.64 ; 
      RECT 0.56 34.736 56.576 35.64 ; 
      RECT 0.02 31.266 0.488 35.64 ; 
      RECT 120.8 31.266 121.412 34.928 ; 
      RECT 65.072 31.266 120.728 35.64 ; 
      RECT 62.084 31.266 65 34.928 ; 
      RECT 61.148 32.048 61.94 35.64 ; 
      RECT 56.432 31.664 61.04 34.928 ; 
      RECT 0.704 31.266 56.36 35.64 ; 
      RECT 0.02 31.266 0.632 34.928 ; 
      RECT 61.868 31.266 121.412 34.544 ; 
      RECT 0.02 31.664 61.796 34.544 ; 
      RECT 60.968 31.266 121.412 31.952 ; 
      RECT 0.02 31.266 60.896 34.544 ; 
      RECT 0.02 31.266 121.412 31.568 ; 
      RECT 0.02 39.44 121.412 39.96 ; 
      RECT 120.944 35.586 121.412 39.96 ; 
      RECT 64.856 39.056 120.872 39.96 ; 
      RECT 59.528 39.056 64.784 39.96 ; 
      RECT 56.648 35.586 59.168 39.96 ; 
      RECT 0.56 39.056 56.576 39.96 ; 
      RECT 0.02 35.586 0.488 39.96 ; 
      RECT 120.8 35.586 121.412 39.248 ; 
      RECT 65.072 35.586 120.728 39.96 ; 
      RECT 62.084 35.586 65 39.248 ; 
      RECT 61.148 36.368 61.94 39.96 ; 
      RECT 56.432 35.984 61.04 39.248 ; 
      RECT 0.704 35.586 56.36 39.96 ; 
      RECT 0.02 35.586 0.632 39.248 ; 
      RECT 61.868 35.586 121.412 38.864 ; 
      RECT 0.02 35.984 61.796 38.864 ; 
      RECT 60.968 35.586 121.412 36.272 ; 
      RECT 0.02 35.586 60.896 38.864 ; 
      RECT 0.02 35.586 121.412 35.888 ; 
      RECT 0 69.334 121.392 74.668 ; 
      RECT 70.884 40.054 121.392 74.668 ; 
      RECT 62.084 45.91 121.392 74.668 ; 
      RECT 65.7 45.142 121.392 74.668 ; 
      RECT 61.876 40.054 62.012 74.668 ; 
      RECT 61.668 40.054 61.804 74.668 ; 
      RECT 61.46 40.054 61.596 74.668 ; 
      RECT 61.252 40.054 61.388 74.668 ; 
      RECT 0 46.294 61.18 74.668 ; 
      RECT 0 56.662 121.392 68.47 ; 
      RECT 56.628 43.99 63.324 55.798 ; 
      RECT 0 45.142 56.556 74.668 ; 
      RECT 0 45.526 65.628 46.198 ; 
      RECT 64.836 45.142 121.392 45.814 ; 
      RECT 0 45.142 64.764 46.198 ; 
      RECT 70.02 40.054 70.812 74.668 ; 
      RECT 54.9 44.374 69.948 45.43 ; 
      RECT 51.444 42.838 54.828 74.668 ; 
      RECT 0 40.054 51.372 74.668 ; 
      RECT 69.156 40.054 121.392 45.046 ; 
      RECT 68.292 42.838 121.392 45.046 ; 
      RECT 63.396 43.99 68.22 45.43 ; 
      RECT 0 43.99 63.324 45.046 ; 
      RECT 67.428 40.054 69.084 44.278 ; 
      RECT 65.052 42.838 121.392 44.278 ; 
      RECT 62.084 42.838 64.98 44.278 ; 
      RECT 56.412 42.838 61.18 46.198 ; 
      RECT 0 42.838 56.34 45.046 ; 
      RECT 62.244 42.646 67.356 43.126 ; 
      RECT 57.492 42.646 62.172 43.126 ; 
      RECT 54.036 42.646 57.42 43.126 ; 
      RECT 52.308 42.646 53.964 74.668 ; 
      RECT 0 40.054 52.236 45.046 ; 
      RECT 66.564 40.054 121.392 42.742 ; 
      RECT 60.66 40.054 66.492 42.742 ; 
      RECT 56.772 40.054 60.588 42.742 ; 
      RECT 53.172 40.054 56.7 42.742 ; 
      RECT 0 40.054 53.1 42.742 ; 
      RECT 0 40.054 121.392 42.55 ; 
        RECT 0.02 76.268 121.412 76.788 ; 
        RECT 120.944 72.414 121.412 76.788 ; 
        RECT 64.856 75.884 120.872 76.788 ; 
        RECT 59.528 75.884 64.784 76.788 ; 
        RECT 56.648 72.414 59.168 76.788 ; 
        RECT 0.56 75.884 56.576 76.788 ; 
        RECT 0.02 72.414 0.488 76.788 ; 
        RECT 120.8 72.414 121.412 76.076 ; 
        RECT 65.072 72.414 120.728 76.788 ; 
        RECT 62.084 72.414 65 76.076 ; 
        RECT 61.148 73.196 61.94 76.788 ; 
        RECT 56.432 72.812 61.04 76.076 ; 
        RECT 0.704 72.414 56.36 76.788 ; 
        RECT 0.02 72.414 0.632 76.076 ; 
        RECT 61.868 72.414 121.412 75.692 ; 
        RECT 0.02 72.812 61.796 75.692 ; 
        RECT 60.968 72.414 121.412 73.1 ; 
        RECT 0.02 72.414 60.896 75.692 ; 
        RECT 0.02 72.414 121.412 72.716 ; 
        RECT 0.02 80.588 121.412 81.108 ; 
        RECT 120.944 76.734 121.412 81.108 ; 
        RECT 64.856 80.204 120.872 81.108 ; 
        RECT 59.528 80.204 64.784 81.108 ; 
        RECT 56.648 76.734 59.168 81.108 ; 
        RECT 0.56 80.204 56.576 81.108 ; 
        RECT 0.02 76.734 0.488 81.108 ; 
        RECT 120.8 76.734 121.412 80.396 ; 
        RECT 65.072 76.734 120.728 81.108 ; 
        RECT 62.084 76.734 65 80.396 ; 
        RECT 61.148 77.516 61.94 81.108 ; 
        RECT 56.432 77.132 61.04 80.396 ; 
        RECT 0.704 76.734 56.36 81.108 ; 
        RECT 0.02 76.734 0.632 80.396 ; 
        RECT 61.868 76.734 121.412 80.012 ; 
        RECT 0.02 77.132 61.796 80.012 ; 
        RECT 60.968 76.734 121.412 77.42 ; 
        RECT 0.02 76.734 60.896 80.012 ; 
        RECT 0.02 76.734 121.412 77.036 ; 
        RECT 0.02 84.908 121.412 85.428 ; 
        RECT 120.944 81.054 121.412 85.428 ; 
        RECT 64.856 84.524 120.872 85.428 ; 
        RECT 59.528 84.524 64.784 85.428 ; 
        RECT 56.648 81.054 59.168 85.428 ; 
        RECT 0.56 84.524 56.576 85.428 ; 
        RECT 0.02 81.054 0.488 85.428 ; 
        RECT 120.8 81.054 121.412 84.716 ; 
        RECT 65.072 81.054 120.728 85.428 ; 
        RECT 62.084 81.054 65 84.716 ; 
        RECT 61.148 81.836 61.94 85.428 ; 
        RECT 56.432 81.452 61.04 84.716 ; 
        RECT 0.704 81.054 56.36 85.428 ; 
        RECT 0.02 81.054 0.632 84.716 ; 
        RECT 61.868 81.054 121.412 84.332 ; 
        RECT 0.02 81.452 61.796 84.332 ; 
        RECT 60.968 81.054 121.412 81.74 ; 
        RECT 0.02 81.054 60.896 84.332 ; 
        RECT 0.02 81.054 121.412 81.356 ; 
        RECT 0.02 89.228 121.412 89.748 ; 
        RECT 120.944 85.374 121.412 89.748 ; 
        RECT 64.856 88.844 120.872 89.748 ; 
        RECT 59.528 88.844 64.784 89.748 ; 
        RECT 56.648 85.374 59.168 89.748 ; 
        RECT 0.56 88.844 56.576 89.748 ; 
        RECT 0.02 85.374 0.488 89.748 ; 
        RECT 120.8 85.374 121.412 89.036 ; 
        RECT 65.072 85.374 120.728 89.748 ; 
        RECT 62.084 85.374 65 89.036 ; 
        RECT 61.148 86.156 61.94 89.748 ; 
        RECT 56.432 85.772 61.04 89.036 ; 
        RECT 0.704 85.374 56.36 89.748 ; 
        RECT 0.02 85.374 0.632 89.036 ; 
        RECT 61.868 85.374 121.412 88.652 ; 
        RECT 0.02 85.772 61.796 88.652 ; 
        RECT 60.968 85.374 121.412 86.06 ; 
        RECT 0.02 85.374 60.896 88.652 ; 
        RECT 0.02 85.374 121.412 85.676 ; 
        RECT 0.02 93.548 121.412 94.068 ; 
        RECT 120.944 89.694 121.412 94.068 ; 
        RECT 64.856 93.164 120.872 94.068 ; 
        RECT 59.528 93.164 64.784 94.068 ; 
        RECT 56.648 89.694 59.168 94.068 ; 
        RECT 0.56 93.164 56.576 94.068 ; 
        RECT 0.02 89.694 0.488 94.068 ; 
        RECT 120.8 89.694 121.412 93.356 ; 
        RECT 65.072 89.694 120.728 94.068 ; 
        RECT 62.084 89.694 65 93.356 ; 
        RECT 61.148 90.476 61.94 94.068 ; 
        RECT 56.432 90.092 61.04 93.356 ; 
        RECT 0.704 89.694 56.36 94.068 ; 
        RECT 0.02 89.694 0.632 93.356 ; 
        RECT 61.868 89.694 121.412 92.972 ; 
        RECT 0.02 90.092 61.796 92.972 ; 
        RECT 60.968 89.694 121.412 90.38 ; 
        RECT 0.02 89.694 60.896 92.972 ; 
        RECT 0.02 89.694 121.412 89.996 ; 
        RECT 0.02 97.868 121.412 98.388 ; 
        RECT 120.944 94.014 121.412 98.388 ; 
        RECT 64.856 97.484 120.872 98.388 ; 
        RECT 59.528 97.484 64.784 98.388 ; 
        RECT 56.648 94.014 59.168 98.388 ; 
        RECT 0.56 97.484 56.576 98.388 ; 
        RECT 0.02 94.014 0.488 98.388 ; 
        RECT 120.8 94.014 121.412 97.676 ; 
        RECT 65.072 94.014 120.728 98.388 ; 
        RECT 62.084 94.014 65 97.676 ; 
        RECT 61.148 94.796 61.94 98.388 ; 
        RECT 56.432 94.412 61.04 97.676 ; 
        RECT 0.704 94.014 56.36 98.388 ; 
        RECT 0.02 94.014 0.632 97.676 ; 
        RECT 61.868 94.014 121.412 97.292 ; 
        RECT 0.02 94.412 61.796 97.292 ; 
        RECT 60.968 94.014 121.412 94.7 ; 
        RECT 0.02 94.014 60.896 97.292 ; 
        RECT 0.02 94.014 121.412 94.316 ; 
        RECT 0.02 102.188 121.412 102.708 ; 
        RECT 120.944 98.334 121.412 102.708 ; 
        RECT 64.856 101.804 120.872 102.708 ; 
        RECT 59.528 101.804 64.784 102.708 ; 
        RECT 56.648 98.334 59.168 102.708 ; 
        RECT 0.56 101.804 56.576 102.708 ; 
        RECT 0.02 98.334 0.488 102.708 ; 
        RECT 120.8 98.334 121.412 101.996 ; 
        RECT 65.072 98.334 120.728 102.708 ; 
        RECT 62.084 98.334 65 101.996 ; 
        RECT 61.148 99.116 61.94 102.708 ; 
        RECT 56.432 98.732 61.04 101.996 ; 
        RECT 0.704 98.334 56.36 102.708 ; 
        RECT 0.02 98.334 0.632 101.996 ; 
        RECT 61.868 98.334 121.412 101.612 ; 
        RECT 0.02 98.732 61.796 101.612 ; 
        RECT 60.968 98.334 121.412 99.02 ; 
        RECT 0.02 98.334 60.896 101.612 ; 
        RECT 0.02 98.334 121.412 98.636 ; 
        RECT 0.02 106.508 121.412 107.028 ; 
        RECT 120.944 102.654 121.412 107.028 ; 
        RECT 64.856 106.124 120.872 107.028 ; 
        RECT 59.528 106.124 64.784 107.028 ; 
        RECT 56.648 102.654 59.168 107.028 ; 
        RECT 0.56 106.124 56.576 107.028 ; 
        RECT 0.02 102.654 0.488 107.028 ; 
        RECT 120.8 102.654 121.412 106.316 ; 
        RECT 65.072 102.654 120.728 107.028 ; 
        RECT 62.084 102.654 65 106.316 ; 
        RECT 61.148 103.436 61.94 107.028 ; 
        RECT 56.432 103.052 61.04 106.316 ; 
        RECT 0.704 102.654 56.36 107.028 ; 
        RECT 0.02 102.654 0.632 106.316 ; 
        RECT 61.868 102.654 121.412 105.932 ; 
        RECT 0.02 103.052 61.796 105.932 ; 
        RECT 60.968 102.654 121.412 103.34 ; 
        RECT 0.02 102.654 60.896 105.932 ; 
        RECT 0.02 102.654 121.412 102.956 ; 
        RECT 0.02 110.828 121.412 111.348 ; 
        RECT 120.944 106.974 121.412 111.348 ; 
        RECT 64.856 110.444 120.872 111.348 ; 
        RECT 59.528 110.444 64.784 111.348 ; 
        RECT 56.648 106.974 59.168 111.348 ; 
        RECT 0.56 110.444 56.576 111.348 ; 
        RECT 0.02 106.974 0.488 111.348 ; 
        RECT 120.8 106.974 121.412 110.636 ; 
        RECT 65.072 106.974 120.728 111.348 ; 
        RECT 62.084 106.974 65 110.636 ; 
        RECT 61.148 107.756 61.94 111.348 ; 
        RECT 56.432 107.372 61.04 110.636 ; 
        RECT 0.704 106.974 56.36 111.348 ; 
        RECT 0.02 106.974 0.632 110.636 ; 
        RECT 61.868 106.974 121.412 110.252 ; 
        RECT 0.02 107.372 61.796 110.252 ; 
        RECT 60.968 106.974 121.412 107.66 ; 
        RECT 0.02 106.974 60.896 110.252 ; 
        RECT 0.02 106.974 121.412 107.276 ; 
  LAYER M4 ; 
      RECT 6.4 46.906 115.342 47.002 ; 
      RECT 6.4 48.058 115.342 48.154 ; 
      RECT 6.4 49.594 115.342 49.69 ; 
      RECT 6.4 49.978 115.342 50.074 ; 
      RECT 6.4 51.322 115.342 51.418 ; 
      RECT 6.4 52.858 115.342 52.954 ; 
      RECT 6.4 53.242 115.342 53.338 ; 
      RECT 41.904 41.398 79.488 42.262 ; 
      RECT 71.468 42.742 71.804 42.838 ; 
      RECT 70.714 44.47 71.234 44.566 ; 
      RECT 70.748 48.25 71.216 48.346 ; 
      RECT 70.746 47.1 71.214 47.196 ; 
      RECT 68.15 44.47 70.434 44.566 ; 
      RECT 68.39 47.53 68.822 47.626 ; 
      RECT 63.1 49.078 67.472 49.174 ; 
      RECT 65.852 47.35 66.188 47.446 ; 
      RECT 62.716 52.15 66.188 52.246 ; 
      RECT 65.852 52.534 66.188 52.63 ; 
      RECT 65.14 45.43 65.476 45.526 ; 
      RECT 64.988 50.806 65.324 50.902 ; 
      RECT 64.988 53.686 65.324 53.782 ; 
      RECT 63.912 40.278 64.964 40.374 ; 
      RECT 64.436 55.414 64.884 55.51 ; 
      RECT 64.276 45.046 64.612 45.142 ; 
      RECT 63.42 39.894 64.472 39.99 ; 
      RECT 63.42 74.314 64.472 74.41 ; 
      RECT 63.484 50.998 64.46 51.094 ; 
      RECT 64.124 51.574 64.46 51.67 ; 
      RECT 58.3 52.534 64.46 52.63 ; 
      RECT 64.124 53.686 64.46 53.782 ; 
      RECT 63.188 73.93 64.24 74.026 ; 
      RECT 63.184 39.51 64.236 39.606 ; 
      RECT 57.24 54.07 64.152 54.934 ; 
      RECT 57.24 66.742 64.152 67.606 ; 
      RECT 63.032 39.126 64.084 39.222 ; 
      RECT 63.032 73.162 64.084 73.258 ; 
      RECT 63.692 55.414 64.028 55.51 ; 
      RECT 60.604 56.95 64.028 57.046 ; 
      RECT 62.14 65.974 64.028 66.07 ; 
      RECT 63.692 66.358 64.028 66.454 ; 
      RECT 62.84 38.742 63.892 38.838 ; 
      RECT 62.84 72.778 63.892 72.874 ; 
      RECT 61.948 62.326 63.728 62.422 ; 
      RECT 62.664 38.358 63.716 38.454 ; 
      RECT 62.664 74.122 63.716 74.218 ; 
      RECT 62.468 39.702 63.52 39.798 ; 
      RECT 62.468 73.738 63.52 73.834 ; 
      RECT 62.992 51.574 63.476 51.67 ; 
      RECT 62.908 60.022 63.44 60.118 ; 
      RECT 62.28 39.318 63.332 39.414 ; 
      RECT 62.28 73.354 63.332 73.45 ; 
      RECT 62.14 38.166 63.192 38.262 ; 
      RECT 62.14 72.97 63.192 73.066 ; 
      RECT 58.876 66.358 63.152 66.454 ; 
      RECT 62.816 70.966 63.152 71.062 ; 
      RECT 61.916 37.59 62.968 37.686 ; 
      RECT 61.916 72.586 62.968 72.682 ; 
      RECT 62.524 55.414 62.864 55.51 ; 
      RECT 58.108 57.718 62.576 57.814 ; 
      RECT 60.688 49.078 62.516 49.174 ; 
      RECT 59.996 40.47 61.064 40.566 ; 
      RECT 59.996 72.01 61.064 72.106 ; 
      RECT 60.544 55.222 60.98 55.318 ; 
      RECT 59.904 40.086 60.872 40.182 ; 
      RECT 59.904 74.506 60.872 74.602 ; 
      RECT 59.68 38.166 60.648 38.262 ; 
      RECT 59.796 74.89 60.648 74.986 ; 
      RECT 60.26 53.686 60.596 53.782 ; 
      RECT 59.464 38.55 60.456 38.646 ; 
      RECT 59.464 74.314 60.456 74.41 ; 
      RECT 58.528 64.054 60.212 64.15 ; 
      RECT 58.4 39.894 59.468 39.99 ; 
      RECT 58.4 74.89 59.468 74.986 ; 
      RECT 58.96 58.294 59.444 58.39 ; 
      RECT 58.928 70.966 59.264 71.062 ; 
      RECT 58.264 39.51 59.252 39.606 ; 
      RECT 57.996 73.162 59.252 73.258 ; 
      RECT 58.16 39.126 59.08 39.222 ; 
      RECT 58.112 74.506 59.08 74.602 ; 
      RECT 57.948 38.742 58.868 38.838 ; 
      RECT 58.532 64.63 58.868 64.726 ; 
      RECT 57.748 72.778 58.868 72.874 ; 
      RECT 57.768 38.358 58.688 38.454 ; 
      RECT 57.768 74.122 58.688 74.218 ; 
      RECT 53.92 53.686 58.676 53.782 ; 
      RECT 57.616 39.318 58.536 39.414 ; 
      RECT 57.616 73.738 58.536 73.834 ; 
      RECT 57.544 38.934 58.316 39.03 ; 
      RECT 57.544 73.354 58.316 73.45 ; 
      RECT 57.348 38.55 58.12 38.646 ; 
      RECT 57.348 72.97 58.12 73.066 ; 
      RECT 57.364 57.334 58.1 57.43 ; 
      RECT 57.14 38.166 57.912 38.262 ; 
      RECT 57.14 72.586 57.912 72.682 ; 
      RECT 55.204 46.582 57.908 46.678 ; 
      RECT 57.364 57.718 57.7 57.814 ; 
      RECT 56.288 40.278 57.34 40.374 ; 
      RECT 56.78 49.078 57.116 49.174 ; 
      RECT 56.504 55.414 56.952 55.51 ; 
      RECT 55.052 47.35 55.388 47.446 ; 
  LAYER V4 ; 
      RECT 71.664 42.742 71.76 42.838 ; 
      RECT 71.664 46.906 71.76 47.002 ; 
      RECT 70.992 47.1 71.088 47.196 ; 
      RECT 70.992 48.25 71.088 48.346 ; 
      RECT 70.99 44.47 71.086 44.566 ; 
      RECT 68.454 44.47 68.55 44.566 ; 
      RECT 68.454 47.53 68.55 47.626 ; 
      RECT 66.048 47.35 66.144 47.446 ; 
      RECT 66.048 48.058 66.144 48.154 ; 
      RECT 66.048 52.15 66.144 52.246 ; 
      RECT 66.048 52.534 66.144 52.63 ; 
      RECT 65.184 45.43 65.28 45.526 ; 
      RECT 65.184 49.594 65.28 49.69 ; 
      RECT 65.184 50.806 65.28 50.902 ; 
      RECT 65.184 51.322 65.28 51.418 ; 
      RECT 65.184 52.858 65.28 52.954 ; 
      RECT 65.184 53.686 65.28 53.782 ; 
      RECT 64.508 40.278 64.604 40.374 ; 
      RECT 64.512 41.398 64.604 42.262 ; 
      RECT 64.508 55.414 64.604 55.51 ; 
      RECT 64.32 45.046 64.416 45.142 ; 
      RECT 64.32 49.978 64.416 50.074 ; 
      RECT 64.32 50.998 64.416 51.094 ; 
      RECT 64.32 51.574 64.416 51.67 ; 
      RECT 64.32 52.534 64.416 52.63 ; 
      RECT 64.32 53.686 64.416 53.782 ; 
      RECT 63.888 55.414 63.984 55.51 ; 
      RECT 63.888 56.95 63.984 57.046 ; 
      RECT 63.888 65.974 63.984 66.07 ; 
      RECT 63.888 66.358 63.984 66.454 ; 
      RECT 63.528 39.894 63.624 39.99 ; 
      RECT 63.528 50.998 63.624 51.094 ; 
      RECT 63.528 74.314 63.624 74.41 ; 
      RECT 63.336 39.51 63.432 39.606 ; 
      RECT 63.336 51.574 63.432 51.67 ; 
      RECT 63.336 73.93 63.432 74.026 ; 
      RECT 63.144 39.126 63.24 39.222 ; 
      RECT 63.144 49.078 63.24 49.174 ; 
      RECT 63.144 73.162 63.24 73.258 ; 
      RECT 62.952 38.742 63.048 38.838 ; 
      RECT 62.952 60.022 63.048 60.118 ; 
      RECT 62.952 70.966 63.048 71.062 ; 
      RECT 62.952 72.778 63.048 72.874 ; 
      RECT 62.76 38.358 62.856 38.454 ; 
      RECT 62.76 52.15 62.856 52.246 ; 
      RECT 62.76 74.122 62.856 74.218 ; 
      RECT 62.568 39.702 62.664 39.798 ; 
      RECT 62.568 55.414 62.664 55.51 ; 
      RECT 62.568 73.738 62.664 73.834 ; 
      RECT 62.376 39.318 62.472 39.414 ; 
      RECT 62.376 49.078 62.472 49.174 ; 
      RECT 62.376 73.354 62.472 73.45 ; 
      RECT 62.184 38.166 62.28 38.262 ; 
      RECT 62.184 65.974 62.28 66.07 ; 
      RECT 62.184 72.97 62.28 73.066 ; 
      RECT 61.992 37.59 62.088 37.686 ; 
      RECT 61.992 62.326 62.088 62.422 ; 
      RECT 61.992 72.586 62.088 72.682 ; 
      RECT 60.84 40.47 60.936 40.566 ; 
      RECT 60.84 55.222 60.936 55.318 ; 
      RECT 60.84 72.01 60.936 72.106 ; 
      RECT 60.648 40.086 60.744 40.182 ; 
      RECT 60.648 56.95 60.744 57.046 ; 
      RECT 60.648 74.506 60.744 74.602 ; 
      RECT 60.456 38.166 60.552 38.262 ; 
      RECT 60.456 53.686 60.552 53.782 ; 
      RECT 60.456 74.89 60.552 74.986 ; 
      RECT 60.072 38.55 60.168 38.646 ; 
      RECT 60.072 64.054 60.168 64.15 ; 
      RECT 60.072 74.314 60.168 74.41 ; 
      RECT 59.304 39.894 59.4 39.99 ; 
      RECT 59.304 58.294 59.4 58.39 ; 
      RECT 59.304 74.89 59.4 74.986 ; 
      RECT 59.112 39.51 59.208 39.606 ; 
      RECT 59.112 70.966 59.208 71.062 ; 
      RECT 59.112 73.162 59.208 73.258 ; 
      RECT 58.92 39.126 59.016 39.222 ; 
      RECT 58.92 66.358 59.016 66.454 ; 
      RECT 58.92 74.506 59.016 74.602 ; 
      RECT 58.728 38.742 58.824 38.838 ; 
      RECT 58.728 64.63 58.824 64.726 ; 
      RECT 58.728 72.778 58.824 72.874 ; 
      RECT 58.536 38.358 58.632 38.454 ; 
      RECT 58.536 53.686 58.632 53.782 ; 
      RECT 58.536 74.122 58.632 74.218 ; 
      RECT 58.344 39.318 58.44 39.414 ; 
      RECT 58.344 52.534 58.44 52.63 ; 
      RECT 58.344 73.738 58.44 73.834 ; 
      RECT 58.152 38.934 58.248 39.03 ; 
      RECT 58.152 57.718 58.248 57.814 ; 
      RECT 58.152 73.354 58.248 73.45 ; 
      RECT 57.96 38.55 58.056 38.646 ; 
      RECT 57.96 57.334 58.056 57.43 ; 
      RECT 57.96 72.97 58.056 73.066 ; 
      RECT 57.768 38.166 57.864 38.262 ; 
      RECT 57.768 46.582 57.864 46.678 ; 
      RECT 57.768 72.586 57.864 72.682 ; 
      RECT 57.408 57.334 57.504 57.43 ; 
      RECT 57.408 57.718 57.504 57.814 ; 
      RECT 56.976 49.078 57.072 49.174 ; 
      RECT 56.976 53.242 57.072 53.338 ; 
      RECT 56.736 40.278 56.832 40.374 ; 
      RECT 56.74 41.398 56.832 42.262 ; 
      RECT 56.736 55.414 56.832 55.51 ; 
      RECT 55.248 46.582 55.344 46.678 ; 
      RECT 55.248 47.35 55.344 47.446 ; 
  LAYER M5 ; 
      RECT 71.664 42.698 71.76 47.046 ; 
      RECT 70.99 44.288 71.086 48.53 ; 
      RECT 68.454 44.304 68.55 47.788 ; 
      RECT 66.048 47.306 66.144 48.198 ; 
      RECT 66.048 52.106 66.144 52.674 ; 
      RECT 65.184 45.386 65.28 49.734 ; 
      RECT 65.184 50.762 65.28 51.462 ; 
      RECT 65.184 52.814 65.28 53.826 ; 
      RECT 64.508 40.206 64.604 55.582 ; 
      RECT 64.32 45.002 64.416 50.118 ; 
      RECT 64.32 50.954 64.416 51.714 ; 
      RECT 64.32 52.49 64.416 53.826 ; 
      RECT 63.888 55.37 63.984 57.09 ; 
      RECT 63.888 65.93 63.984 66.498 ; 
      RECT 63.528 37.284 63.624 75.29 ; 
      RECT 63.336 37.284 63.432 75.286 ; 
      RECT 63.144 37.284 63.24 75.286 ; 
      RECT 62.952 37.284 63.048 75.17 ; 
      RECT 62.76 37.284 62.856 75.158 ; 
      RECT 62.568 37.284 62.664 75.166 ; 
      RECT 62.376 37.284 62.472 75.138 ; 
      RECT 62.184 37.284 62.28 75.202 ; 
      RECT 61.992 37.284 62.088 75.198 ; 
      RECT 60.84 38.106 60.936 75.422 ; 
      RECT 60.648 38.11 60.744 75.426 ; 
      RECT 60.456 38.106 60.552 75.422 ; 
      RECT 60.072 38.17 60.168 75.426 ; 
      RECT 59.304 38.166 59.4 75.238 ; 
      RECT 59.112 38.166 59.208 75.238 ; 
      RECT 58.92 38.166 59.016 75.238 ; 
      RECT 58.728 38.166 58.824 75.238 ; 
      RECT 58.536 38.166 58.632 75.238 ; 
      RECT 58.344 38.05 58.44 75.238 ; 
      RECT 58.152 37.874 58.248 74.094 ; 
      RECT 57.96 37.726 58.056 73.91 ; 
      RECT 57.768 37.51 57.864 73.694 ; 
      RECT 57.408 57.29 57.504 57.858 ; 
      RECT 56.976 49.034 57.072 53.382 ; 
      RECT 56.736 40.206 56.832 55.582 ; 
      RECT 55.248 46.538 55.344 47.49 ; 
  LAYER M2 ; 
    RECT 0.432 0.144 120.96 112.176 ; 
  LAYER M1 ; 
    RECT 0.432 0.144 120.96 112.176 ; 
  END 
END srambank_256x4x18_6t122 
