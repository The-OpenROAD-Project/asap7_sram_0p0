VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO srambank_256x4x20_6t122
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN srambank_256x4x20_6t122 0 0 ;
  SIZE 30.348 BY 30.240000000000002 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1040 1.1720 30.2580 1.2200 ;
        RECT 0.1040 2.2520 30.2580 2.3000 ;
        RECT 0.1040 3.3320 30.2580 3.3800 ;
        RECT 0.1040 4.4120 30.2580 4.4600 ;
        RECT 0.1040 5.4920 30.2580 5.5400 ;
        RECT 0.1040 6.5720 30.2580 6.6200 ;
        RECT 0.1040 7.6520 30.2580 7.7000 ;
        RECT 0.1040 8.7320 30.2580 8.7800 ;
        RECT 0.1040 9.8120 30.2580 9.8600 ;
        RECT 0.1040 10.8920 30.2580 10.9400 ;
        RECT 0.1040 20.0990 30.2580 20.1470 ;
        RECT 0.1040 21.1790 30.2580 21.2270 ;
        RECT 0.1040 22.2590 30.2580 22.3070 ;
        RECT 0.1040 23.3390 30.2580 23.3870 ;
        RECT 0.1040 24.4190 30.2580 24.4670 ;
        RECT 0.1040 25.4990 30.2580 25.5470 ;
        RECT 0.1040 26.5790 30.2580 26.6270 ;
        RECT 0.1040 27.6590 30.2580 27.7070 ;
        RECT 0.1040 28.7390 30.2580 28.7870 ;
        RECT 0.1040 29.8190 30.2580 29.8670 ;
      LAYER M3  ;
        RECT 30.2180 0.2165 30.2360 1.3765 ;
        RECT 16.1960 0.2170 16.2140 1.3760 ;
        RECT 14.7920 0.2530 14.8820 1.3685 ;
        RECT 14.1440 0.2170 14.1620 1.3760 ;
        RECT 0.1220 0.2165 0.1400 1.3765 ;
        RECT 30.2180 1.2965 30.2360 2.4565 ;
        RECT 16.1960 1.2970 16.2140 2.4560 ;
        RECT 14.7920 1.3330 14.8820 2.4485 ;
        RECT 14.1440 1.2970 14.1620 2.4560 ;
        RECT 0.1220 1.2965 0.1400 2.4565 ;
        RECT 30.2180 2.3765 30.2360 3.5365 ;
        RECT 16.1960 2.3770 16.2140 3.5360 ;
        RECT 14.7920 2.4130 14.8820 3.5285 ;
        RECT 14.1440 2.3770 14.1620 3.5360 ;
        RECT 0.1220 2.3765 0.1400 3.5365 ;
        RECT 30.2180 3.4565 30.2360 4.6165 ;
        RECT 16.1960 3.4570 16.2140 4.6160 ;
        RECT 14.7920 3.4930 14.8820 4.6085 ;
        RECT 14.1440 3.4570 14.1620 4.6160 ;
        RECT 0.1220 3.4565 0.1400 4.6165 ;
        RECT 30.2180 4.5365 30.2360 5.6965 ;
        RECT 16.1960 4.5370 16.2140 5.6960 ;
        RECT 14.7920 4.5730 14.8820 5.6885 ;
        RECT 14.1440 4.5370 14.1620 5.6960 ;
        RECT 0.1220 4.5365 0.1400 5.6965 ;
        RECT 30.2180 5.6165 30.2360 6.7765 ;
        RECT 16.1960 5.6170 16.2140 6.7760 ;
        RECT 14.7920 5.6530 14.8820 6.7685 ;
        RECT 14.1440 5.6170 14.1620 6.7760 ;
        RECT 0.1220 5.6165 0.1400 6.7765 ;
        RECT 30.2180 6.6965 30.2360 7.8565 ;
        RECT 16.1960 6.6970 16.2140 7.8560 ;
        RECT 14.7920 6.7330 14.8820 7.8485 ;
        RECT 14.1440 6.6970 14.1620 7.8560 ;
        RECT 0.1220 6.6965 0.1400 7.8565 ;
        RECT 30.2180 7.7765 30.2360 8.9365 ;
        RECT 16.1960 7.7770 16.2140 8.9360 ;
        RECT 14.7920 7.8130 14.8820 8.9285 ;
        RECT 14.1440 7.7770 14.1620 8.9360 ;
        RECT 0.1220 7.7765 0.1400 8.9365 ;
        RECT 30.2180 8.8565 30.2360 10.0165 ;
        RECT 16.1960 8.8570 16.2140 10.0160 ;
        RECT 14.7920 8.8930 14.8820 10.0085 ;
        RECT 14.1440 8.8570 14.1620 10.0160 ;
        RECT 0.1220 8.8565 0.1400 10.0165 ;
        RECT 30.2180 9.9365 30.2360 11.0965 ;
        RECT 16.1960 9.9370 16.2140 11.0960 ;
        RECT 14.7920 9.9730 14.8820 11.0885 ;
        RECT 14.1440 9.9370 14.1620 11.0960 ;
        RECT 0.1220 9.9365 0.1400 11.0965 ;
        RECT 14.0490 14.8850 14.0670 20.9485 ;
        RECT 30.2180 19.1435 30.2360 20.3035 ;
        RECT 16.1960 19.1440 16.2140 20.3030 ;
        RECT 14.7920 19.1800 14.8820 20.2955 ;
        RECT 14.1440 19.1440 14.1620 20.3030 ;
        RECT 0.1220 19.1435 0.1400 20.3035 ;
        RECT 30.2180 20.2235 30.2360 21.3835 ;
        RECT 16.1960 20.2240 16.2140 21.3830 ;
        RECT 14.7920 20.2600 14.8820 21.3755 ;
        RECT 14.1440 20.2240 14.1620 21.3830 ;
        RECT 0.1220 20.2235 0.1400 21.3835 ;
        RECT 30.2180 21.3035 30.2360 22.4635 ;
        RECT 16.1960 21.3040 16.2140 22.4630 ;
        RECT 14.7920 21.3400 14.8820 22.4555 ;
        RECT 14.1440 21.3040 14.1620 22.4630 ;
        RECT 0.1220 21.3035 0.1400 22.4635 ;
        RECT 30.2180 22.3835 30.2360 23.5435 ;
        RECT 16.1960 22.3840 16.2140 23.5430 ;
        RECT 14.7920 22.4200 14.8820 23.5355 ;
        RECT 14.1440 22.3840 14.1620 23.5430 ;
        RECT 0.1220 22.3835 0.1400 23.5435 ;
        RECT 30.2180 23.4635 30.2360 24.6235 ;
        RECT 16.1960 23.4640 16.2140 24.6230 ;
        RECT 14.7920 23.5000 14.8820 24.6155 ;
        RECT 14.1440 23.4640 14.1620 24.6230 ;
        RECT 0.1220 23.4635 0.1400 24.6235 ;
        RECT 30.2180 24.5435 30.2360 25.7035 ;
        RECT 16.1960 24.5440 16.2140 25.7030 ;
        RECT 14.7920 24.5800 14.8820 25.6955 ;
        RECT 14.1440 24.5440 14.1620 25.7030 ;
        RECT 0.1220 24.5435 0.1400 25.7035 ;
        RECT 30.2180 25.6235 30.2360 26.7835 ;
        RECT 16.1960 25.6240 16.2140 26.7830 ;
        RECT 14.7920 25.6600 14.8820 26.7755 ;
        RECT 14.1440 25.6240 14.1620 26.7830 ;
        RECT 0.1220 25.6235 0.1400 26.7835 ;
        RECT 30.2180 26.7035 30.2360 27.8635 ;
        RECT 16.1960 26.7040 16.2140 27.8630 ;
        RECT 14.7920 26.7400 14.8820 27.8555 ;
        RECT 14.1440 26.7040 14.1620 27.8630 ;
        RECT 0.1220 26.7035 0.1400 27.8635 ;
        RECT 30.2180 27.7835 30.2360 28.9435 ;
        RECT 16.1960 27.7840 16.2140 28.9430 ;
        RECT 14.7920 27.8200 14.8820 28.9355 ;
        RECT 14.1440 27.7840 14.1620 28.9430 ;
        RECT 0.1220 27.7835 0.1400 28.9435 ;
        RECT 30.2180 28.8635 30.2360 30.0235 ;
        RECT 16.1960 28.8640 16.2140 30.0230 ;
        RECT 14.7920 28.9000 14.8820 30.0155 ;
        RECT 14.1440 28.8640 14.1620 30.0230 ;
        RECT 0.1220 28.8635 0.1400 30.0235 ;
      LAYER V3  ;
        RECT 0.1220 1.1720 0.1400 1.2200 ;
        RECT 14.1440 1.1720 14.1620 1.2200 ;
        RECT 14.7920 1.1720 14.8820 1.2200 ;
        RECT 16.1960 1.1720 16.2140 1.2200 ;
        RECT 30.2180 1.1720 30.2360 1.2200 ;
        RECT 0.1220 2.2520 0.1400 2.3000 ;
        RECT 14.1440 2.2520 14.1620 2.3000 ;
        RECT 14.7920 2.2520 14.8820 2.3000 ;
        RECT 16.1960 2.2520 16.2140 2.3000 ;
        RECT 30.2180 2.2520 30.2360 2.3000 ;
        RECT 0.1220 3.3320 0.1400 3.3800 ;
        RECT 14.1440 3.3320 14.1620 3.3800 ;
        RECT 14.7920 3.3320 14.8820 3.3800 ;
        RECT 16.1960 3.3320 16.2140 3.3800 ;
        RECT 30.2180 3.3320 30.2360 3.3800 ;
        RECT 0.1220 4.4120 0.1400 4.4600 ;
        RECT 14.1440 4.4120 14.1620 4.4600 ;
        RECT 14.7920 4.4120 14.8820 4.4600 ;
        RECT 16.1960 4.4120 16.2140 4.4600 ;
        RECT 30.2180 4.4120 30.2360 4.4600 ;
        RECT 0.1220 5.4920 0.1400 5.5400 ;
        RECT 14.1440 5.4920 14.1620 5.5400 ;
        RECT 14.7920 5.4920 14.8820 5.5400 ;
        RECT 16.1960 5.4920 16.2140 5.5400 ;
        RECT 30.2180 5.4920 30.2360 5.5400 ;
        RECT 0.1220 6.5720 0.1400 6.6200 ;
        RECT 14.1440 6.5720 14.1620 6.6200 ;
        RECT 14.7920 6.5720 14.8820 6.6200 ;
        RECT 16.1960 6.5720 16.2140 6.6200 ;
        RECT 30.2180 6.5720 30.2360 6.6200 ;
        RECT 0.1220 7.6520 0.1400 7.7000 ;
        RECT 14.1440 7.6520 14.1620 7.7000 ;
        RECT 14.7920 7.6520 14.8820 7.7000 ;
        RECT 16.1960 7.6520 16.2140 7.7000 ;
        RECT 30.2180 7.6520 30.2360 7.7000 ;
        RECT 0.1220 8.7320 0.1400 8.7800 ;
        RECT 14.1440 8.7320 14.1620 8.7800 ;
        RECT 14.7920 8.7320 14.8820 8.7800 ;
        RECT 16.1960 8.7320 16.2140 8.7800 ;
        RECT 30.2180 8.7320 30.2360 8.7800 ;
        RECT 0.1220 9.8120 0.1400 9.8600 ;
        RECT 14.1440 9.8120 14.1620 9.8600 ;
        RECT 14.7920 9.8120 14.8820 9.8600 ;
        RECT 16.1960 9.8120 16.2140 9.8600 ;
        RECT 30.2180 9.8120 30.2360 9.8600 ;
        RECT 0.1220 10.8920 0.1400 10.9400 ;
        RECT 14.1440 10.8920 14.1620 10.9400 ;
        RECT 14.7920 10.8920 14.8820 10.9400 ;
        RECT 16.1960 10.8920 16.2140 10.9400 ;
        RECT 30.2180 10.8920 30.2360 10.9400 ;
        RECT 0.1220 20.0990 0.1400 20.1470 ;
        RECT 14.1440 20.0990 14.1620 20.1470 ;
        RECT 14.7920 20.0990 14.8820 20.1470 ;
        RECT 16.1960 20.0990 16.2140 20.1470 ;
        RECT 30.2180 20.0990 30.2360 20.1470 ;
        RECT 0.1220 21.1790 0.1400 21.2270 ;
        RECT 14.1440 21.1790 14.1620 21.2270 ;
        RECT 14.7920 21.1790 14.8820 21.2270 ;
        RECT 16.1960 21.1790 16.2140 21.2270 ;
        RECT 30.2180 21.1790 30.2360 21.2270 ;
        RECT 0.1220 22.2590 0.1400 22.3070 ;
        RECT 14.1440 22.2590 14.1620 22.3070 ;
        RECT 14.7920 22.2590 14.8820 22.3070 ;
        RECT 16.1960 22.2590 16.2140 22.3070 ;
        RECT 30.2180 22.2590 30.2360 22.3070 ;
        RECT 0.1220 23.3390 0.1400 23.3870 ;
        RECT 14.1440 23.3390 14.1620 23.3870 ;
        RECT 14.7920 23.3390 14.8820 23.3870 ;
        RECT 16.1960 23.3390 16.2140 23.3870 ;
        RECT 30.2180 23.3390 30.2360 23.3870 ;
        RECT 0.1220 24.4190 0.1400 24.4670 ;
        RECT 14.1440 24.4190 14.1620 24.4670 ;
        RECT 14.7920 24.4190 14.8820 24.4670 ;
        RECT 16.1960 24.4190 16.2140 24.4670 ;
        RECT 30.2180 24.4190 30.2360 24.4670 ;
        RECT 0.1220 25.4990 0.1400 25.5470 ;
        RECT 14.1440 25.4990 14.1620 25.5470 ;
        RECT 14.7920 25.4990 14.8820 25.5470 ;
        RECT 16.1960 25.4990 16.2140 25.5470 ;
        RECT 30.2180 25.4990 30.2360 25.5470 ;
        RECT 0.1220 26.5790 0.1400 26.6270 ;
        RECT 14.1440 26.5790 14.1620 26.6270 ;
        RECT 14.7920 26.5790 14.8820 26.6270 ;
        RECT 16.1960 26.5790 16.2140 26.6270 ;
        RECT 30.2180 26.5790 30.2360 26.6270 ;
        RECT 0.1220 27.6590 0.1400 27.7070 ;
        RECT 14.1440 27.6590 14.1620 27.7070 ;
        RECT 14.7920 27.6590 14.8820 27.7070 ;
        RECT 16.1960 27.6590 16.2140 27.7070 ;
        RECT 30.2180 27.6590 30.2360 27.7070 ;
        RECT 0.1220 28.7390 0.1400 28.7870 ;
        RECT 14.1440 28.7390 14.1620 28.7870 ;
        RECT 14.7920 28.7390 14.8820 28.7870 ;
        RECT 16.1960 28.7390 16.2140 28.7870 ;
        RECT 30.2180 28.7390 30.2360 28.7870 ;
        RECT 0.1220 29.8190 0.1400 29.8670 ;
        RECT 14.1440 29.8190 14.1620 29.8670 ;
        RECT 14.7920 29.8190 14.8820 29.8670 ;
        RECT 16.1960 29.8190 16.2140 29.8670 ;
        RECT 30.2180 29.8190 30.2360 29.8670 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4  ;
        RECT 0.1040 1.0760 30.2580 1.1240 ;
        RECT 0.1040 2.1560 30.2580 2.2040 ;
        RECT 0.1040 3.2360 30.2580 3.2840 ;
        RECT 0.1040 4.3160 30.2580 4.3640 ;
        RECT 0.1040 5.3960 30.2580 5.4440 ;
        RECT 0.1040 6.4760 30.2580 6.5240 ;
        RECT 0.1040 7.5560 30.2580 7.6040 ;
        RECT 0.1040 8.6360 30.2580 8.6840 ;
        RECT 0.1040 9.7160 30.2580 9.7640 ;
        RECT 0.1040 10.7960 30.2580 10.8440 ;
        RECT 10.4760 11.8615 19.8720 12.0775 ;
        RECT 14.3100 15.0295 16.0380 15.2455 ;
        RECT 14.3100 18.1975 16.0380 18.4135 ;
        RECT 0.1040 20.0030 30.2580 20.0510 ;
        RECT 0.1040 21.0830 30.2580 21.1310 ;
        RECT 0.1040 22.1630 30.2580 22.2110 ;
        RECT 0.1040 23.2430 30.2580 23.2910 ;
        RECT 0.1040 24.3230 30.2580 24.3710 ;
        RECT 0.1040 25.4030 30.2580 25.4510 ;
        RECT 0.1040 26.4830 30.2580 26.5310 ;
        RECT 0.1040 27.5630 30.2580 27.6110 ;
        RECT 0.1040 28.6430 30.2580 28.6910 ;
        RECT 0.1040 29.7230 30.2580 29.7710 ;
      LAYER M3  ;
        RECT 30.1820 0.2165 30.2000 1.3765 ;
        RECT 16.2500 0.2165 16.2680 1.3765 ;
        RECT 15.4850 0.2530 15.5210 1.3675 ;
        RECT 15.2600 0.2530 15.2870 1.3675 ;
        RECT 14.0900 0.2165 14.1080 1.3765 ;
        RECT 0.1580 0.2165 0.1760 1.3765 ;
        RECT 30.1820 1.2965 30.2000 2.4565 ;
        RECT 16.2500 1.2965 16.2680 2.4565 ;
        RECT 15.4850 1.3330 15.5210 2.4475 ;
        RECT 15.2600 1.3330 15.2870 2.4475 ;
        RECT 14.0900 1.2965 14.1080 2.4565 ;
        RECT 0.1580 1.2965 0.1760 2.4565 ;
        RECT 30.1820 2.3765 30.2000 3.5365 ;
        RECT 16.2500 2.3765 16.2680 3.5365 ;
        RECT 15.4850 2.4130 15.5210 3.5275 ;
        RECT 15.2600 2.4130 15.2870 3.5275 ;
        RECT 14.0900 2.3765 14.1080 3.5365 ;
        RECT 0.1580 2.3765 0.1760 3.5365 ;
        RECT 30.1820 3.4565 30.2000 4.6165 ;
        RECT 16.2500 3.4565 16.2680 4.6165 ;
        RECT 15.4850 3.4930 15.5210 4.6075 ;
        RECT 15.2600 3.4930 15.2870 4.6075 ;
        RECT 14.0900 3.4565 14.1080 4.6165 ;
        RECT 0.1580 3.4565 0.1760 4.6165 ;
        RECT 30.1820 4.5365 30.2000 5.6965 ;
        RECT 16.2500 4.5365 16.2680 5.6965 ;
        RECT 15.4850 4.5730 15.5210 5.6875 ;
        RECT 15.2600 4.5730 15.2870 5.6875 ;
        RECT 14.0900 4.5365 14.1080 5.6965 ;
        RECT 0.1580 4.5365 0.1760 5.6965 ;
        RECT 30.1820 5.6165 30.2000 6.7765 ;
        RECT 16.2500 5.6165 16.2680 6.7765 ;
        RECT 15.4850 5.6530 15.5210 6.7675 ;
        RECT 15.2600 5.6530 15.2870 6.7675 ;
        RECT 14.0900 5.6165 14.1080 6.7765 ;
        RECT 0.1580 5.6165 0.1760 6.7765 ;
        RECT 30.1820 6.6965 30.2000 7.8565 ;
        RECT 16.2500 6.6965 16.2680 7.8565 ;
        RECT 15.4850 6.7330 15.5210 7.8475 ;
        RECT 15.2600 6.7330 15.2870 7.8475 ;
        RECT 14.0900 6.6965 14.1080 7.8565 ;
        RECT 0.1580 6.6965 0.1760 7.8565 ;
        RECT 30.1820 7.7765 30.2000 8.9365 ;
        RECT 16.2500 7.7765 16.2680 8.9365 ;
        RECT 15.4850 7.8130 15.5210 8.9275 ;
        RECT 15.2600 7.8130 15.2870 8.9275 ;
        RECT 14.0900 7.7765 14.1080 8.9365 ;
        RECT 0.1580 7.7765 0.1760 8.9365 ;
        RECT 30.1820 8.8565 30.2000 10.0165 ;
        RECT 16.2500 8.8565 16.2680 10.0165 ;
        RECT 15.4850 8.8930 15.5210 10.0075 ;
        RECT 15.2600 8.8930 15.2870 10.0075 ;
        RECT 14.0900 8.8565 14.1080 10.0165 ;
        RECT 0.1580 8.8565 0.1760 10.0165 ;
        RECT 30.1820 9.9365 30.2000 11.0965 ;
        RECT 16.2500 9.9365 16.2680 11.0965 ;
        RECT 15.4850 9.9730 15.5210 11.0875 ;
        RECT 15.2600 9.9730 15.2870 11.0875 ;
        RECT 14.0900 9.9365 14.1080 11.0965 ;
        RECT 0.1580 9.9365 0.1760 11.0965 ;
        RECT 16.2450 11.0670 16.2630 19.2740 ;
        RECT 15.2910 11.2905 15.5250 18.9735 ;
        RECT 14.0850 11.0670 14.1030 20.9485 ;
        RECT 30.1820 19.1435 30.2000 20.3035 ;
        RECT 16.2500 19.1435 16.2680 20.3035 ;
        RECT 15.4850 19.1800 15.5210 20.2945 ;
        RECT 15.2600 19.1800 15.2870 20.2945 ;
        RECT 14.0900 19.1435 14.1080 20.3035 ;
        RECT 0.1580 19.1435 0.1760 20.3035 ;
        RECT 30.1820 20.2235 30.2000 21.3835 ;
        RECT 16.2500 20.2235 16.2680 21.3835 ;
        RECT 15.4850 20.2600 15.5210 21.3745 ;
        RECT 15.2600 20.2600 15.2870 21.3745 ;
        RECT 14.0900 20.2235 14.1080 21.3835 ;
        RECT 0.1580 20.2235 0.1760 21.3835 ;
        RECT 30.1820 21.3035 30.2000 22.4635 ;
        RECT 16.2500 21.3035 16.2680 22.4635 ;
        RECT 15.4850 21.3400 15.5210 22.4545 ;
        RECT 15.2600 21.3400 15.2870 22.4545 ;
        RECT 14.0900 21.3035 14.1080 22.4635 ;
        RECT 0.1580 21.3035 0.1760 22.4635 ;
        RECT 30.1820 22.3835 30.2000 23.5435 ;
        RECT 16.2500 22.3835 16.2680 23.5435 ;
        RECT 15.4850 22.4200 15.5210 23.5345 ;
        RECT 15.2600 22.4200 15.2870 23.5345 ;
        RECT 14.0900 22.3835 14.1080 23.5435 ;
        RECT 0.1580 22.3835 0.1760 23.5435 ;
        RECT 30.1820 23.4635 30.2000 24.6235 ;
        RECT 16.2500 23.4635 16.2680 24.6235 ;
        RECT 15.4850 23.5000 15.5210 24.6145 ;
        RECT 15.2600 23.5000 15.2870 24.6145 ;
        RECT 14.0900 23.4635 14.1080 24.6235 ;
        RECT 0.1580 23.4635 0.1760 24.6235 ;
        RECT 30.1820 24.5435 30.2000 25.7035 ;
        RECT 16.2500 24.5435 16.2680 25.7035 ;
        RECT 15.4850 24.5800 15.5210 25.6945 ;
        RECT 15.2600 24.5800 15.2870 25.6945 ;
        RECT 14.0900 24.5435 14.1080 25.7035 ;
        RECT 0.1580 24.5435 0.1760 25.7035 ;
        RECT 30.1820 25.6235 30.2000 26.7835 ;
        RECT 16.2500 25.6235 16.2680 26.7835 ;
        RECT 15.4850 25.6600 15.5210 26.7745 ;
        RECT 15.2600 25.6600 15.2870 26.7745 ;
        RECT 14.0900 25.6235 14.1080 26.7835 ;
        RECT 0.1580 25.6235 0.1760 26.7835 ;
        RECT 30.1820 26.7035 30.2000 27.8635 ;
        RECT 16.2500 26.7035 16.2680 27.8635 ;
        RECT 15.4850 26.7400 15.5210 27.8545 ;
        RECT 15.2600 26.7400 15.2870 27.8545 ;
        RECT 14.0900 26.7035 14.1080 27.8635 ;
        RECT 0.1580 26.7035 0.1760 27.8635 ;
        RECT 30.1820 27.7835 30.2000 28.9435 ;
        RECT 16.2500 27.7835 16.2680 28.9435 ;
        RECT 15.4850 27.8200 15.5210 28.9345 ;
        RECT 15.2600 27.8200 15.2870 28.9345 ;
        RECT 14.0900 27.7835 14.1080 28.9435 ;
        RECT 0.1580 27.7835 0.1760 28.9435 ;
        RECT 30.1820 28.8635 30.2000 30.0235 ;
        RECT 16.2500 28.8635 16.2680 30.0235 ;
        RECT 15.4850 28.9000 15.5210 30.0145 ;
        RECT 15.2600 28.9000 15.2870 30.0145 ;
        RECT 14.0900 28.8635 14.1080 30.0235 ;
        RECT 0.1580 28.8635 0.1760 30.0235 ;
      LAYER V3  ;
        RECT 0.1580 1.0760 0.1760 1.1240 ;
        RECT 14.0900 1.0760 14.1080 1.1240 ;
        RECT 15.2600 1.0760 15.2870 1.1240 ;
        RECT 15.4850 1.0760 15.5210 1.1240 ;
        RECT 16.2500 1.0760 16.2680 1.1240 ;
        RECT 30.1820 1.0760 30.2000 1.1240 ;
        RECT 0.1580 2.1560 0.1760 2.2040 ;
        RECT 14.0900 2.1560 14.1080 2.2040 ;
        RECT 15.2600 2.1560 15.2870 2.2040 ;
        RECT 15.4850 2.1560 15.5210 2.2040 ;
        RECT 16.2500 2.1560 16.2680 2.2040 ;
        RECT 30.1820 2.1560 30.2000 2.2040 ;
        RECT 0.1580 3.2360 0.1760 3.2840 ;
        RECT 14.0900 3.2360 14.1080 3.2840 ;
        RECT 15.2600 3.2360 15.2870 3.2840 ;
        RECT 15.4850 3.2360 15.5210 3.2840 ;
        RECT 16.2500 3.2360 16.2680 3.2840 ;
        RECT 30.1820 3.2360 30.2000 3.2840 ;
        RECT 0.1580 4.3160 0.1760 4.3640 ;
        RECT 14.0900 4.3160 14.1080 4.3640 ;
        RECT 15.2600 4.3160 15.2870 4.3640 ;
        RECT 15.4850 4.3160 15.5210 4.3640 ;
        RECT 16.2500 4.3160 16.2680 4.3640 ;
        RECT 30.1820 4.3160 30.2000 4.3640 ;
        RECT 0.1580 5.3960 0.1760 5.4440 ;
        RECT 14.0900 5.3960 14.1080 5.4440 ;
        RECT 15.2600 5.3960 15.2870 5.4440 ;
        RECT 15.4850 5.3960 15.5210 5.4440 ;
        RECT 16.2500 5.3960 16.2680 5.4440 ;
        RECT 30.1820 5.3960 30.2000 5.4440 ;
        RECT 0.1580 6.4760 0.1760 6.5240 ;
        RECT 14.0900 6.4760 14.1080 6.5240 ;
        RECT 15.2600 6.4760 15.2870 6.5240 ;
        RECT 15.4850 6.4760 15.5210 6.5240 ;
        RECT 16.2500 6.4760 16.2680 6.5240 ;
        RECT 30.1820 6.4760 30.2000 6.5240 ;
        RECT 0.1580 7.5560 0.1760 7.6040 ;
        RECT 14.0900 7.5560 14.1080 7.6040 ;
        RECT 15.2600 7.5560 15.2870 7.6040 ;
        RECT 15.4850 7.5560 15.5210 7.6040 ;
        RECT 16.2500 7.5560 16.2680 7.6040 ;
        RECT 30.1820 7.5560 30.2000 7.6040 ;
        RECT 0.1580 8.6360 0.1760 8.6840 ;
        RECT 14.0900 8.6360 14.1080 8.6840 ;
        RECT 15.2600 8.6360 15.2870 8.6840 ;
        RECT 15.4850 8.6360 15.5210 8.6840 ;
        RECT 16.2500 8.6360 16.2680 8.6840 ;
        RECT 30.1820 8.6360 30.2000 8.6840 ;
        RECT 0.1580 9.7160 0.1760 9.7640 ;
        RECT 14.0900 9.7160 14.1080 9.7640 ;
        RECT 15.2600 9.7160 15.2870 9.7640 ;
        RECT 15.4850 9.7160 15.5210 9.7640 ;
        RECT 16.2500 9.7160 16.2680 9.7640 ;
        RECT 30.1820 9.7160 30.2000 9.7640 ;
        RECT 0.1580 10.7960 0.1760 10.8440 ;
        RECT 14.0900 10.7960 14.1080 10.8440 ;
        RECT 15.2600 10.7960 15.2870 10.8440 ;
        RECT 15.4850 10.7960 15.5210 10.8440 ;
        RECT 16.2500 10.7960 16.2680 10.8440 ;
        RECT 30.1820 10.7960 30.2000 10.8440 ;
        RECT 14.0850 11.8615 14.1030 12.0775 ;
        RECT 15.2950 18.1975 15.3130 18.4135 ;
        RECT 15.2950 15.0295 15.3130 15.2455 ;
        RECT 15.2950 11.8615 15.3130 12.0775 ;
        RECT 15.3470 18.1975 15.3650 18.4135 ;
        RECT 15.3470 15.0295 15.3650 15.2455 ;
        RECT 15.3470 11.8615 15.3650 12.0775 ;
        RECT 15.3990 18.1975 15.4170 18.4135 ;
        RECT 15.3990 15.0295 15.4170 15.2455 ;
        RECT 15.3990 11.8615 15.4170 12.0775 ;
        RECT 15.4510 18.1975 15.4690 18.4135 ;
        RECT 15.4510 15.0295 15.4690 15.2455 ;
        RECT 15.4510 11.8615 15.4690 12.0775 ;
        RECT 15.5030 18.1975 15.5210 18.4135 ;
        RECT 15.5030 15.0295 15.5210 15.2455 ;
        RECT 15.5030 11.8615 15.5210 12.0775 ;
        RECT 16.2450 11.8615 16.2630 12.0775 ;
        RECT 0.1580 20.0030 0.1760 20.0510 ;
        RECT 14.0900 20.0030 14.1080 20.0510 ;
        RECT 15.2600 20.0030 15.2870 20.0510 ;
        RECT 15.4850 20.0030 15.5210 20.0510 ;
        RECT 16.2500 20.0030 16.2680 20.0510 ;
        RECT 30.1820 20.0030 30.2000 20.0510 ;
        RECT 0.1580 21.0830 0.1760 21.1310 ;
        RECT 14.0900 21.0830 14.1080 21.1310 ;
        RECT 15.2600 21.0830 15.2870 21.1310 ;
        RECT 15.4850 21.0830 15.5210 21.1310 ;
        RECT 16.2500 21.0830 16.2680 21.1310 ;
        RECT 30.1820 21.0830 30.2000 21.1310 ;
        RECT 0.1580 22.1630 0.1760 22.2110 ;
        RECT 14.0900 22.1630 14.1080 22.2110 ;
        RECT 15.2600 22.1630 15.2870 22.2110 ;
        RECT 15.4850 22.1630 15.5210 22.2110 ;
        RECT 16.2500 22.1630 16.2680 22.2110 ;
        RECT 30.1820 22.1630 30.2000 22.2110 ;
        RECT 0.1580 23.2430 0.1760 23.2910 ;
        RECT 14.0900 23.2430 14.1080 23.2910 ;
        RECT 15.2600 23.2430 15.2870 23.2910 ;
        RECT 15.4850 23.2430 15.5210 23.2910 ;
        RECT 16.2500 23.2430 16.2680 23.2910 ;
        RECT 30.1820 23.2430 30.2000 23.2910 ;
        RECT 0.1580 24.3230 0.1760 24.3710 ;
        RECT 14.0900 24.3230 14.1080 24.3710 ;
        RECT 15.2600 24.3230 15.2870 24.3710 ;
        RECT 15.4850 24.3230 15.5210 24.3710 ;
        RECT 16.2500 24.3230 16.2680 24.3710 ;
        RECT 30.1820 24.3230 30.2000 24.3710 ;
        RECT 0.1580 25.4030 0.1760 25.4510 ;
        RECT 14.0900 25.4030 14.1080 25.4510 ;
        RECT 15.2600 25.4030 15.2870 25.4510 ;
        RECT 15.4850 25.4030 15.5210 25.4510 ;
        RECT 16.2500 25.4030 16.2680 25.4510 ;
        RECT 30.1820 25.4030 30.2000 25.4510 ;
        RECT 0.1580 26.4830 0.1760 26.5310 ;
        RECT 14.0900 26.4830 14.1080 26.5310 ;
        RECT 15.2600 26.4830 15.2870 26.5310 ;
        RECT 15.4850 26.4830 15.5210 26.5310 ;
        RECT 16.2500 26.4830 16.2680 26.5310 ;
        RECT 30.1820 26.4830 30.2000 26.5310 ;
        RECT 0.1580 27.5630 0.1760 27.6110 ;
        RECT 14.0900 27.5630 14.1080 27.6110 ;
        RECT 15.2600 27.5630 15.2870 27.6110 ;
        RECT 15.4850 27.5630 15.5210 27.6110 ;
        RECT 16.2500 27.5630 16.2680 27.6110 ;
        RECT 30.1820 27.5630 30.2000 27.6110 ;
        RECT 0.1580 28.6430 0.1760 28.6910 ;
        RECT 14.0900 28.6430 14.1080 28.6910 ;
        RECT 15.2600 28.6430 15.2870 28.6910 ;
        RECT 15.4850 28.6430 15.5210 28.6910 ;
        RECT 16.2500 28.6430 16.2680 28.6910 ;
        RECT 30.1820 28.6430 30.2000 28.6910 ;
        RECT 0.1580 29.7230 0.1760 29.7710 ;
        RECT 14.0900 29.7230 14.1080 29.7710 ;
        RECT 15.2600 29.7230 15.2870 29.7710 ;
        RECT 15.4850 29.7230 15.5210 29.7710 ;
        RECT 16.2500 29.7230 16.2680 29.7710 ;
        RECT 30.1820 29.7230 30.2000 29.7710 ;
    END
  END VSS
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.7030 12.3335 17.7210 12.3705 ;
      LAYER M4  ;
        RECT 17.6510 12.3415 17.7350 12.3655 ;
      LAYER M5  ;
        RECT 17.7000 11.3905 17.7240 14.6305 ;
      LAYER V3  ;
        RECT 17.7030 12.3415 17.7210 12.3655 ;
      LAYER V4  ;
        RECT 17.7000 12.3415 17.7240 12.3655 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.4870 12.3365 17.5050 12.3735 ;
      LAYER M4  ;
        RECT 17.4350 12.3415 17.5190 12.3655 ;
      LAYER M5  ;
        RECT 17.4840 11.3905 17.5080 14.6305 ;
      LAYER V3  ;
        RECT 17.4870 12.3415 17.5050 12.3655 ;
      LAYER V4  ;
        RECT 17.4840 12.3415 17.5080 12.3655 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.2710 11.7575 17.2890 11.7945 ;
      LAYER M4  ;
        RECT 17.2190 11.7655 17.3030 11.7895 ;
      LAYER M5  ;
        RECT 17.2680 11.3905 17.2920 14.6305 ;
      LAYER V3  ;
        RECT 17.2710 11.7655 17.2890 11.7895 ;
      LAYER V4  ;
        RECT 17.2680 11.7655 17.2920 11.7895 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 17.0550 11.9975 17.0730 12.1785 ;
      LAYER M4  ;
        RECT 17.0030 12.1495 17.0870 12.1735 ;
      LAYER M5  ;
        RECT 17.0520 11.3905 17.0760 14.6305 ;
      LAYER V3  ;
        RECT 17.0550 12.1495 17.0730 12.1735 ;
      LAYER V4  ;
        RECT 17.0520 12.1495 17.0760 12.1735 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.8390 11.7605 16.8570 11.8275 ;
      LAYER M4  ;
        RECT 16.7870 11.7655 16.8710 11.7895 ;
      LAYER M5  ;
        RECT 16.8360 11.3905 16.8600 14.6305 ;
      LAYER V3  ;
        RECT 16.8390 11.7655 16.8570 11.7895 ;
      LAYER V4  ;
        RECT 16.8360 11.7655 16.8600 11.7895 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.6230 11.4935 16.6410 11.7465 ;
      LAYER M4  ;
        RECT 16.5710 11.7175 16.6550 11.7415 ;
      LAYER M5  ;
        RECT 16.6200 11.3905 16.6440 14.6305 ;
      LAYER V3  ;
        RECT 16.6230 11.7175 16.6410 11.7415 ;
      LAYER V4  ;
        RECT 16.6200 11.7175 16.6440 11.7415 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.4070 12.5285 16.4250 12.5655 ;
      LAYER M4  ;
        RECT 16.3550 12.5335 16.4390 12.5575 ;
      LAYER M5  ;
        RECT 16.4040 11.3905 16.4280 14.6305 ;
      LAYER V3  ;
        RECT 16.4070 12.5335 16.4250 12.5575 ;
      LAYER V4  ;
        RECT 16.4040 12.5335 16.4280 12.5575 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 16.1910 12.3755 16.2090 12.4665 ;
      LAYER M4  ;
        RECT 16.1390 12.4375 16.2230 12.4615 ;
      LAYER M5  ;
        RECT 16.1880 11.3905 16.2120 14.6305 ;
      LAYER V3  ;
        RECT 16.1910 12.4375 16.2090 12.4615 ;
      LAYER V4  ;
        RECT 16.1880 12.4375 16.2120 12.4615 ;
    END
  END ADDRESS[7]
  PIN ADDRESS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.8310 12.0335 15.8490 12.1785 ;
      LAYER M4  ;
        RECT 15.8200 12.1495 16.0070 12.1735 ;
      LAYER M5  ;
        RECT 15.9720 11.1315 15.9960 14.6305 ;
      LAYER V3  ;
        RECT 15.8310 12.1495 15.8490 12.1735 ;
      LAYER V4  ;
        RECT 15.9720 12.1495 15.9960 12.1735 ;
    END
  END ADDRESS[8]
  PIN ADDRESS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.5430 11.7605 15.5610 11.8275 ;
      LAYER M4  ;
        RECT 15.2590 11.7655 15.5720 11.7895 ;
      LAYER M5  ;
        RECT 15.2700 11.3905 15.2940 14.6305 ;
      LAYER V3  ;
        RECT 15.5430 11.7655 15.5610 11.7895 ;
      LAYER V4  ;
        RECT 15.2700 11.7655 15.2940 11.7895 ;
    END
  END ADDRESS[9]
  PIN banksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.1470 11.4935 15.1650 11.7465 ;
      LAYER M4  ;
        RECT 14.9350 11.7175 15.1760 11.7415 ;
      LAYER M5  ;
        RECT 14.9460 11.3905 14.9700 14.6305 ;
      LAYER V3  ;
        RECT 15.1470 11.7175 15.1650 11.7415 ;
      LAYER V4  ;
        RECT 14.9460 11.7175 14.9700 11.7415 ;
    END
  END banksel
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.1390 12.6245 14.1570 12.6735 ;
      LAYER M4  ;
        RECT 14.0870 12.6295 14.1710 12.6535 ;
      LAYER M5  ;
        RECT 14.1360 11.3905 14.1600 14.6305 ;
      LAYER V3  ;
        RECT 14.1390 12.6295 14.1570 12.6535 ;
      LAYER V4  ;
        RECT 14.1360 12.6295 14.1600 12.6535 ;
    END
  END clk
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.3550 11.7605 14.3730 11.8275 ;
      LAYER M4  ;
        RECT 14.3030 11.7655 14.3870 11.7895 ;
      LAYER M5  ;
        RECT 14.3520 11.3905 14.3760 14.6305 ;
      LAYER V3  ;
        RECT 14.3550 11.7655 14.3730 11.7895 ;
      LAYER V4  ;
        RECT 14.3520 11.7655 14.3760 11.7895 ;
    END
  END write
  PIN read
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 14.1750 11.4935 14.1930 11.7465 ;
      LAYER M4  ;
        RECT 13.9090 11.7175 14.2040 11.7415 ;
      LAYER M5  ;
        RECT 13.9200 11.3905 13.9440 14.6305 ;
      LAYER V3  ;
        RECT 14.1750 11.7175 14.1930 11.7415 ;
      LAYER V4  ;
        RECT 13.9200 11.7175 13.9440 11.7415 ;
    END
  END read
  PIN sdel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.7070 12.3335 13.7250 12.3705 ;
      LAYER M4  ;
        RECT 13.6550 12.3415 13.7390 12.3655 ;
      LAYER M5  ;
        RECT 13.7040 11.3905 13.7280 14.6305 ;
      LAYER V3  ;
        RECT 13.7070 12.3415 13.7250 12.3655 ;
      LAYER V4  ;
        RECT 13.7040 12.3415 13.7280 12.3655 ;
    END
  END sdel[0]
  PIN sdel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.4910 11.7605 13.5090 11.9895 ;
      LAYER M4  ;
        RECT 13.4390 11.7655 13.5230 11.7895 ;
      LAYER M5  ;
        RECT 13.4880 11.3905 13.5120 14.6305 ;
      LAYER V3  ;
        RECT 13.4910 11.7655 13.5090 11.7895 ;
      LAYER V4  ;
        RECT 13.4880 11.7655 13.5120 11.7895 ;
    END
  END sdel[1]
  PIN sdel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.2750 11.4935 13.2930 11.7465 ;
      LAYER M4  ;
        RECT 13.2230 11.7175 13.3070 11.7415 ;
      LAYER M5  ;
        RECT 13.2720 11.3905 13.2960 14.6305 ;
      LAYER V3  ;
        RECT 13.2750 11.7175 13.2930 11.7415 ;
      LAYER V4  ;
        RECT 13.2720 11.7175 13.2960 11.7415 ;
    END
  END sdel[2]
  PIN sdel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 13.0590 11.7575 13.0770 11.7945 ;
      LAYER M4  ;
        RECT 13.0070 11.7655 13.0910 11.7895 ;
      LAYER M5  ;
        RECT 13.0560 11.3905 13.0800 14.6305 ;
      LAYER V3  ;
        RECT 13.0590 11.7655 13.0770 11.7895 ;
      LAYER V4  ;
        RECT 13.0560 11.7655 13.0800 11.7895 ;
    END
  END sdel[3]
  PIN sdel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 12.8430 12.3335 12.8610 12.3705 ;
      LAYER M4  ;
        RECT 12.7910 12.3415 12.8750 12.3655 ;
      LAYER M5  ;
        RECT 12.8400 11.3905 12.8640 14.6305 ;
      LAYER V3  ;
        RECT 12.8430 12.3415 12.8610 12.3655 ;
      LAYER V4  ;
        RECT 12.8400 12.3415 12.8640 12.3655 ;
    END
  END sdel[4]
  PIN dataout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 23.6245 15.4670 23.8640 ;
      LAYER M4  ;
        RECT 14.8610 23.6750 15.5090 23.6990 ;
      LAYER V3  ;
        RECT 15.4490 23.6750 15.4670 23.6990 ;
    END
  END dataout[14]
  PIN dataout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 22.5445 15.4670 22.7840 ;
      LAYER M4  ;
        RECT 14.8610 22.5950 15.5090 22.6190 ;
      LAYER V3  ;
        RECT 15.4490 22.5950 15.4670 22.6190 ;
    END
  END dataout[13]
  PIN dataout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 21.4645 15.4670 21.7040 ;
      LAYER M4  ;
        RECT 14.8610 21.5150 15.5090 21.5390 ;
      LAYER V3  ;
        RECT 15.4490 21.5150 15.4670 21.5390 ;
    END
  END dataout[12]
  PIN dataout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 20.3845 15.4670 20.6240 ;
      LAYER M4  ;
        RECT 14.8610 20.4350 15.5090 20.4590 ;
      LAYER V3  ;
        RECT 15.4490 20.4350 15.4670 20.4590 ;
    END
  END dataout[11]
  PIN dataout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 19.3045 15.4670 19.5440 ;
      LAYER M4  ;
        RECT 14.8610 19.3550 15.5090 19.3790 ;
      LAYER V3  ;
        RECT 15.4490 19.3550 15.4670 19.3790 ;
    END
  END dataout[10]
  PIN dataout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 0.3775 15.4670 0.6170 ;
      LAYER M4  ;
        RECT 14.8610 0.4280 15.5090 0.4520 ;
      LAYER V3  ;
        RECT 15.4490 0.4280 15.4670 0.4520 ;
    END
  END dataout[0]
  PIN dataout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 24.7045 15.4670 24.9440 ;
      LAYER M4  ;
        RECT 14.8610 24.7550 15.5090 24.7790 ;
      LAYER V3  ;
        RECT 15.4490 24.7550 15.4670 24.7790 ;
    END
  END dataout[15]
  PIN dataout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 25.7845 15.4670 26.0240 ;
      LAYER M4  ;
        RECT 14.8610 25.8350 15.5090 25.8590 ;
      LAYER V3  ;
        RECT 15.4490 25.8350 15.4670 25.8590 ;
    END
  END dataout[16]
  PIN dataout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 26.8645 15.4670 27.1040 ;
      LAYER M4  ;
        RECT 14.8610 26.9150 15.5090 26.9390 ;
      LAYER V3  ;
        RECT 15.4490 26.9150 15.4670 26.9390 ;
    END
  END dataout[17]
  PIN dataout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 27.9445 15.4670 28.1840 ;
      LAYER M4  ;
        RECT 14.8610 27.9950 15.5090 28.0190 ;
      LAYER V3  ;
        RECT 15.4490 27.9950 15.4670 28.0190 ;
    END
  END dataout[18]
  PIN dataout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 29.0245 15.4670 29.2640 ;
      LAYER M4  ;
        RECT 14.8610 29.0750 15.5090 29.0990 ;
      LAYER V3  ;
        RECT 15.4490 29.0750 15.4670 29.0990 ;
    END
  END dataout[19]
  PIN dataout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 1.4575 15.4670 1.6970 ;
      LAYER M4  ;
        RECT 14.8610 1.5080 15.5090 1.5320 ;
      LAYER V3  ;
        RECT 15.4490 1.5080 15.4670 1.5320 ;
    END
  END dataout[1]
  PIN dataout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[20]
  PIN dataout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[21]
  PIN dataout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[22]
  PIN dataout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[23]
  PIN dataout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[24]
  PIN dataout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[25]
  PIN dataout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[26]
  PIN dataout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[27]
  PIN dataout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[28]
  PIN dataout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[29]
  PIN dataout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 2.5375 15.4670 2.7770 ;
      LAYER M4  ;
        RECT 14.8610 2.5880 15.5090 2.6120 ;
      LAYER V3  ;
        RECT 15.4490 2.5880 15.4670 2.6120 ;
    END
  END dataout[2]
  PIN dataout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[30]
  PIN dataout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[31]
  PIN dataout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[32]
  PIN dataout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[33]
  PIN dataout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[34]
  PIN dataout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[35]
  PIN dataout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[36]
  PIN dataout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[37]
  PIN dataout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[38]
  PIN dataout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[39]
  PIN dataout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 3.6175 15.4670 3.8570 ;
      LAYER M4  ;
        RECT 14.8610 3.6680 15.5090 3.6920 ;
      LAYER V3  ;
        RECT 15.4490 3.6680 15.4670 3.6920 ;
    END
  END dataout[3]
  PIN dataout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[40]
  PIN dataout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[41]
  PIN dataout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[42]
  PIN dataout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[43]
  PIN dataout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[44]
  PIN dataout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[45]
  PIN dataout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[46]
  PIN dataout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[47]
  PIN dataout[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[48]
  PIN dataout[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[49]
  PIN dataout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 4.6975 15.4670 4.9370 ;
      LAYER M4  ;
        RECT 14.8610 4.7480 15.5090 4.7720 ;
      LAYER V3  ;
        RECT 15.4490 4.7480 15.4670 4.7720 ;
    END
  END dataout[4]
  PIN dataout[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[50]
  PIN dataout[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[51]
  PIN dataout[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[52]
  PIN dataout[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[53]
  PIN dataout[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[54]
  PIN dataout[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[55]
  PIN dataout[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[56]
  PIN dataout[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[57]
  PIN dataout[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[58]
  PIN dataout[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[59]
  PIN dataout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 5.7775 15.4670 6.0170 ;
      LAYER M4  ;
        RECT 14.8610 5.8280 15.5090 5.8520 ;
      LAYER V3  ;
        RECT 15.4490 5.8280 15.4670 5.8520 ;
    END
  END dataout[5]
  PIN dataout[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[60]
  PIN dataout[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[61]
  PIN dataout[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[62]
  PIN dataout[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END dataout[63]
  PIN dataout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 6.8575 15.4670 7.0970 ;
      LAYER M4  ;
        RECT 14.8610 6.9080 15.5090 6.9320 ;
      LAYER V3  ;
        RECT 15.4490 6.9080 15.4670 6.9320 ;
    END
  END dataout[6]
  PIN dataout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 7.9375 15.4670 8.1770 ;
      LAYER M4  ;
        RECT 14.8610 7.9880 15.5090 8.0120 ;
      LAYER V3  ;
        RECT 15.4490 7.9880 15.4670 8.0120 ;
    END
  END dataout[7]
  PIN dataout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 9.0175 15.4670 9.2570 ;
      LAYER M4  ;
        RECT 14.8610 9.0680 15.5090 9.0920 ;
      LAYER V3  ;
        RECT 15.4490 9.0680 15.4670 9.0920 ;
    END
  END dataout[8]
  PIN dataout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.4490 10.0975 15.4670 10.3370 ;
      LAYER M4  ;
        RECT 14.8610 10.1480 15.5090 10.1720 ;
      LAYER V3  ;
        RECT 15.4490 10.1480 15.4670 10.1720 ;
    END
  END dataout[9]
  PIN wd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 0.2700 15.2420 0.6750 ;
      LAYER M4  ;
        RECT 14.8610 0.3320 15.4970 0.3560 ;
      LAYER V3  ;
        RECT 15.2240 0.3320 15.2420 0.3560 ;
    END
  END wd[0]
  PIN wd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 19.1970 15.2420 19.6020 ;
      LAYER M4  ;
        RECT 14.8610 19.2590 15.4970 19.2830 ;
      LAYER V3  ;
        RECT 15.2240 19.2590 15.2420 19.2830 ;
    END
  END wd[10]
  PIN wd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 20.2770 15.2420 20.6820 ;
      LAYER M4  ;
        RECT 14.8610 20.3390 15.4970 20.3630 ;
      LAYER V3  ;
        RECT 15.2240 20.3390 15.2420 20.3630 ;
    END
  END wd[11]
  PIN wd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 21.3570 15.2420 21.7620 ;
      LAYER M4  ;
        RECT 14.8610 21.4190 15.4970 21.4430 ;
      LAYER V3  ;
        RECT 15.2240 21.4190 15.2420 21.4430 ;
    END
  END wd[12]
  PIN wd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 22.4370 15.2420 22.8420 ;
      LAYER M4  ;
        RECT 14.8610 22.4990 15.4970 22.5230 ;
      LAYER V3  ;
        RECT 15.2240 22.4990 15.2420 22.5230 ;
    END
  END wd[13]
  PIN wd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 23.5170 15.2420 23.9220 ;
      LAYER M4  ;
        RECT 14.8610 23.5790 15.4970 23.6030 ;
      LAYER V3  ;
        RECT 15.2240 23.5790 15.2420 23.6030 ;
    END
  END wd[14]
  PIN wd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 24.5970 15.2420 25.0020 ;
      LAYER M4  ;
        RECT 14.8610 24.6590 15.4970 24.6830 ;
      LAYER V3  ;
        RECT 15.2240 24.6590 15.2420 24.6830 ;
    END
  END wd[15]
  PIN wd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 25.6770 15.2420 26.0820 ;
      LAYER M4  ;
        RECT 14.8610 25.7390 15.4970 25.7630 ;
      LAYER V3  ;
        RECT 15.2240 25.7390 15.2420 25.7630 ;
    END
  END wd[16]
  PIN wd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 26.7570 15.2420 27.1620 ;
      LAYER M4  ;
        RECT 14.8610 26.8190 15.4970 26.8430 ;
      LAYER V3  ;
        RECT 15.2240 26.8190 15.2420 26.8430 ;
    END
  END wd[17]
  PIN wd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 27.8370 15.2420 28.2420 ;
      LAYER M4  ;
        RECT 14.8610 27.8990 15.4970 27.9230 ;
      LAYER V3  ;
        RECT 15.2240 27.8990 15.2420 27.9230 ;
    END
  END wd[18]
  PIN wd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 28.9170 15.2420 29.3220 ;
      LAYER M4  ;
        RECT 14.8610 28.9790 15.4970 29.0030 ;
      LAYER V3  ;
        RECT 15.2240 28.9790 15.2420 29.0030 ;
    END
  END wd[19]
  PIN wd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 1.3500 15.2420 1.7550 ;
      LAYER M4  ;
        RECT 14.8610 1.4120 15.4970 1.4360 ;
      LAYER V3  ;
        RECT 15.2240 1.4120 15.2420 1.4360 ;
    END
  END wd[1]
  PIN wd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[20]
  PIN wd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[21]
  PIN wd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[22]
  PIN wd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[23]
  PIN wd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[24]
  PIN wd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[25]
  PIN wd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[26]
  PIN wd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[27]
  PIN wd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[28]
  PIN wd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[29]
  PIN wd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 2.4300 15.2420 2.8350 ;
      LAYER M4  ;
        RECT 14.8610 2.4920 15.4970 2.5160 ;
      LAYER V3  ;
        RECT 15.2240 2.4920 15.2420 2.5160 ;
    END
  END wd[2]
  PIN wd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[30]
  PIN wd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[31]
  PIN wd[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[32]
  PIN wd[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[33]
  PIN wd[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[34]
  PIN wd[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[35]
  PIN wd[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[36]
  PIN wd[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[37]
  PIN wd[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[38]
  PIN wd[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[39]
  PIN wd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 3.5100 15.2420 3.9150 ;
      LAYER M4  ;
        RECT 14.8610 3.5720 15.4970 3.5960 ;
      LAYER V3  ;
        RECT 15.2240 3.5720 15.2420 3.5960 ;
    END
  END wd[3]
  PIN wd[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[40]
  PIN wd[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[41]
  PIN wd[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[42]
  PIN wd[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[43]
  PIN wd[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[44]
  PIN wd[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[45]
  PIN wd[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[46]
  PIN wd[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[47]
  PIN wd[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[48]
  PIN wd[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[49]
  PIN wd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 4.5900 15.2420 4.9950 ;
      LAYER M4  ;
        RECT 14.8610 4.6520 15.4970 4.6760 ;
      LAYER V3  ;
        RECT 15.2240 4.6520 15.2420 4.6760 ;
    END
  END wd[4]
  PIN wd[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[50]
  PIN wd[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[51]
  PIN wd[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[52]
  PIN wd[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[53]
  PIN wd[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[54]
  PIN wd[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[55]
  PIN wd[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[56]
  PIN wd[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[57]
  PIN wd[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[58]
  PIN wd[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[59]
  PIN wd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 5.6700 15.2420 6.0750 ;
      LAYER M4  ;
        RECT 14.8610 5.7320 15.4970 5.7560 ;
      LAYER V3  ;
        RECT 15.2240 5.7320 15.2420 5.7560 ;
    END
  END wd[5]
  PIN wd[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[60]
  PIN wd[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[61]
  PIN wd[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[62]
  PIN wd[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
    END
  END wd[63]
  PIN wd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 6.7500 15.2420 7.1550 ;
      LAYER M4  ;
        RECT 14.8610 6.8120 15.4970 6.8360 ;
      LAYER V3  ;
        RECT 15.2240 6.8120 15.2420 6.8360 ;
    END
  END wd[6]
  PIN wd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 7.8300 15.2420 8.2350 ;
      LAYER M4  ;
        RECT 14.8610 7.8920 15.4970 7.9160 ;
      LAYER V3  ;
        RECT 15.2240 7.8920 15.2420 7.9160 ;
    END
  END wd[7]
  PIN wd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 8.9100 15.2420 9.3150 ;
      LAYER M4  ;
        RECT 14.8610 8.9720 15.4970 8.9960 ;
      LAYER V3  ;
        RECT 15.2240 8.9720 15.2420 8.9960 ;
    END
  END wd[8]
  PIN wd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3  ;
        RECT 15.2240 9.9900 15.2420 10.3950 ;
      LAYER M4  ;
        RECT 14.8610 10.0520 15.4970 10.0760 ;
      LAYER V3  ;
        RECT 15.2240 10.0520 15.2420 10.0760 ;
    END
  END wd[9]
OBS
  LAYER M1 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0000 11.0935 30.3480 19.7470 ;
        RECT 0.0050 19.1835 30.3530 20.2770 ;
        RECT 0.0050 20.2635 30.3530 21.3570 ;
        RECT 0.0050 21.3435 30.3530 22.4370 ;
        RECT 0.0050 22.4235 30.3530 23.5170 ;
        RECT 0.0050 23.5035 30.3530 24.5970 ;
        RECT 0.0050 24.5835 30.3530 25.6770 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
  LAYER M2 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0000 11.0935 30.3480 19.7470 ;
        RECT 0.0050 19.1835 30.3530 20.2770 ;
        RECT 0.0050 20.2635 30.3530 21.3570 ;
        RECT 0.0050 21.3435 30.3530 22.4370 ;
        RECT 0.0050 22.4235 30.3530 23.5170 ;
        RECT 0.0050 23.5035 30.3530 24.5970 ;
        RECT 0.0050 24.5835 30.3530 25.6770 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
  LAYER V1 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0000 11.0935 30.3480 19.7470 ;
        RECT 0.0050 19.1835 30.3530 20.2770 ;
        RECT 0.0050 20.2635 30.3530 21.3570 ;
        RECT 0.0050 21.3435 30.3530 22.4370 ;
        RECT 0.0050 22.4235 30.3530 23.5170 ;
        RECT 0.0050 23.5035 30.3530 24.5970 ;
        RECT 0.0050 24.5835 30.3530 25.6770 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
  LAYER V2 SPACING 0.018  ;
      RECT 0.0050 0.2565 30.3530 1.3500 ;
      RECT 0.0050 1.3365 30.3530 2.4300 ;
      RECT 0.0050 2.4165 30.3530 3.5100 ;
      RECT 0.0050 3.4965 30.3530 4.5900 ;
      RECT 0.0050 4.5765 30.3530 5.6700 ;
      RECT 0.0050 5.6565 30.3530 6.7500 ;
      RECT 0.0050 6.7365 30.3530 7.8300 ;
      RECT 0.0050 7.8165 30.3530 8.9100 ;
      RECT 0.0050 8.8965 30.3530 9.9900 ;
      RECT 0.0050 9.9765 30.3530 11.0700 ;
      RECT 0.0000 11.0935 30.3480 19.7470 ;
        RECT 0.0050 19.1835 30.3530 20.2770 ;
        RECT 0.0050 20.2635 30.3530 21.3570 ;
        RECT 0.0050 21.3435 30.3530 22.4370 ;
        RECT 0.0050 22.4235 30.3530 23.5170 ;
        RECT 0.0050 23.5035 30.3530 24.5970 ;
        RECT 0.0050 24.5835 30.3530 25.6770 ;
        RECT 0.0050 25.6635 30.3530 26.7570 ;
        RECT 0.0050 26.7435 30.3530 27.8370 ;
        RECT 0.0050 27.8235 30.3530 28.9170 ;
        RECT 0.0050 28.9035 30.3530 29.9970 ;
  LAYER M3  ;
      RECT 15.6110 0.3450 15.6290 1.2805 ;
      RECT 15.5750 0.3450 15.5930 1.2805 ;
      RECT 15.5390 0.9220 15.5570 1.2445 ;
      RECT 15.4220 1.1190 15.4400 1.2285 ;
      RECT 15.4130 0.3775 15.4310 0.6170 ;
      RECT 15.3770 0.9585 15.3950 1.1120 ;
      RECT 15.2960 0.9840 15.3140 1.2420 ;
      RECT 14.7560 0.3450 14.7740 1.2805 ;
      RECT 14.7200 0.3450 14.7380 1.2805 ;
      RECT 14.6840 0.5260 14.7020 1.0940 ;
      RECT 15.6110 1.4250 15.6290 2.3605 ;
      RECT 15.5750 1.4250 15.5930 2.3605 ;
      RECT 15.5390 2.0020 15.5570 2.3245 ;
      RECT 15.4220 2.1990 15.4400 2.3085 ;
      RECT 15.4130 1.4575 15.4310 1.6970 ;
      RECT 15.3770 2.0385 15.3950 2.1920 ;
      RECT 15.2960 2.0640 15.3140 2.3220 ;
      RECT 14.7560 1.4250 14.7740 2.3605 ;
      RECT 14.7200 1.4250 14.7380 2.3605 ;
      RECT 14.6840 1.6060 14.7020 2.1740 ;
      RECT 15.6110 2.5050 15.6290 3.4405 ;
      RECT 15.5750 2.5050 15.5930 3.4405 ;
      RECT 15.5390 3.0820 15.5570 3.4045 ;
      RECT 15.4220 3.2790 15.4400 3.3885 ;
      RECT 15.4130 2.5375 15.4310 2.7770 ;
      RECT 15.3770 3.1185 15.3950 3.2720 ;
      RECT 15.2960 3.1440 15.3140 3.4020 ;
      RECT 14.7560 2.5050 14.7740 3.4405 ;
      RECT 14.7200 2.5050 14.7380 3.4405 ;
      RECT 14.6840 2.6860 14.7020 3.2540 ;
      RECT 15.6110 3.5850 15.6290 4.5205 ;
      RECT 15.5750 3.5850 15.5930 4.5205 ;
      RECT 15.5390 4.1620 15.5570 4.4845 ;
      RECT 15.4220 4.3590 15.4400 4.4685 ;
      RECT 15.4130 3.6175 15.4310 3.8570 ;
      RECT 15.3770 4.1985 15.3950 4.3520 ;
      RECT 15.2960 4.2240 15.3140 4.4820 ;
      RECT 14.7560 3.5850 14.7740 4.5205 ;
      RECT 14.7200 3.5850 14.7380 4.5205 ;
      RECT 14.6840 3.7660 14.7020 4.3340 ;
      RECT 15.6110 4.6650 15.6290 5.6005 ;
      RECT 15.5750 4.6650 15.5930 5.6005 ;
      RECT 15.5390 5.2420 15.5570 5.5645 ;
      RECT 15.4220 5.4390 15.4400 5.5485 ;
      RECT 15.4130 4.6975 15.4310 4.9370 ;
      RECT 15.3770 5.2785 15.3950 5.4320 ;
      RECT 15.2960 5.3040 15.3140 5.5620 ;
      RECT 14.7560 4.6650 14.7740 5.6005 ;
      RECT 14.7200 4.6650 14.7380 5.6005 ;
      RECT 14.6840 4.8460 14.7020 5.4140 ;
      RECT 15.6110 5.7450 15.6290 6.6805 ;
      RECT 15.5750 5.7450 15.5930 6.6805 ;
      RECT 15.5390 6.3220 15.5570 6.6445 ;
      RECT 15.4220 6.5190 15.4400 6.6285 ;
      RECT 15.4130 5.7775 15.4310 6.0170 ;
      RECT 15.3770 6.3585 15.3950 6.5120 ;
      RECT 15.2960 6.3840 15.3140 6.6420 ;
      RECT 14.7560 5.7450 14.7740 6.6805 ;
      RECT 14.7200 5.7450 14.7380 6.6805 ;
      RECT 14.6840 5.9260 14.7020 6.4940 ;
      RECT 15.6110 6.8250 15.6290 7.7605 ;
      RECT 15.5750 6.8250 15.5930 7.7605 ;
      RECT 15.5390 7.4020 15.5570 7.7245 ;
      RECT 15.4220 7.5990 15.4400 7.7085 ;
      RECT 15.4130 6.8575 15.4310 7.0970 ;
      RECT 15.3770 7.4385 15.3950 7.5920 ;
      RECT 15.2960 7.4640 15.3140 7.7220 ;
      RECT 14.7560 6.8250 14.7740 7.7605 ;
      RECT 14.7200 6.8250 14.7380 7.7605 ;
      RECT 14.6840 7.0060 14.7020 7.5740 ;
      RECT 15.6110 7.9050 15.6290 8.8405 ;
      RECT 15.5750 7.9050 15.5930 8.8405 ;
      RECT 15.5390 8.4820 15.5570 8.8045 ;
      RECT 15.4220 8.6790 15.4400 8.7885 ;
      RECT 15.4130 7.9375 15.4310 8.1770 ;
      RECT 15.3770 8.5185 15.3950 8.6720 ;
      RECT 15.2960 8.5440 15.3140 8.8020 ;
      RECT 14.7560 7.9050 14.7740 8.8405 ;
      RECT 14.7200 7.9050 14.7380 8.8405 ;
      RECT 14.6840 8.0860 14.7020 8.6540 ;
      RECT 15.6110 8.9850 15.6290 9.9205 ;
      RECT 15.5750 8.9850 15.5930 9.9205 ;
      RECT 15.5390 9.5620 15.5570 9.8845 ;
      RECT 15.4220 9.7590 15.4400 9.8685 ;
      RECT 15.4130 9.0175 15.4310 9.2570 ;
      RECT 15.3770 9.5985 15.3950 9.7520 ;
      RECT 15.2960 9.6240 15.3140 9.8820 ;
      RECT 14.7560 8.9850 14.7740 9.9205 ;
      RECT 14.7200 8.9850 14.7380 9.9205 ;
      RECT 14.6840 9.1660 14.7020 9.7340 ;
      RECT 15.6110 10.0650 15.6290 11.0005 ;
      RECT 15.5750 10.0650 15.5930 11.0005 ;
      RECT 15.5390 10.6420 15.5570 10.9645 ;
      RECT 15.4220 10.8390 15.4400 10.9485 ;
      RECT 15.4130 10.0975 15.4310 10.3370 ;
      RECT 15.3770 10.6785 15.3950 10.8320 ;
      RECT 15.2960 10.7040 15.3140 10.9620 ;
      RECT 14.7560 10.0650 14.7740 11.0005 ;
      RECT 14.7200 10.0650 14.7380 11.0005 ;
      RECT 14.6840 10.2460 14.7020 10.8140 ;
      RECT 30.2130 10.9035 30.2310 19.2740 ;
      RECT 30.1770 10.9035 30.1950 19.2740 ;
      RECT 30.0690 10.9035 30.0870 14.6445 ;
      RECT 29.9610 10.9035 29.9790 14.6445 ;
      RECT 29.8530 10.9035 29.8710 14.6445 ;
      RECT 29.7450 10.9035 29.7630 14.6445 ;
      RECT 29.6370 10.9035 29.6550 14.6445 ;
      RECT 29.5290 10.9035 29.5470 14.6445 ;
      RECT 29.4210 10.9035 29.4390 14.6445 ;
      RECT 29.3130 10.9035 29.3310 14.6445 ;
      RECT 29.2050 10.9035 29.2230 14.6445 ;
      RECT 29.0970 10.9035 29.1150 14.6445 ;
      RECT 28.9890 10.9035 29.0070 14.6445 ;
      RECT 28.8810 10.9035 28.8990 14.6445 ;
      RECT 28.7730 10.9035 28.7910 14.6445 ;
      RECT 28.6650 10.9035 28.6830 14.6445 ;
      RECT 28.5570 10.9035 28.5750 14.6445 ;
      RECT 28.4490 10.9035 28.4670 14.6445 ;
      RECT 28.3410 10.9035 28.3590 14.6445 ;
      RECT 28.2330 10.9035 28.2510 14.6445 ;
      RECT 28.1250 10.9035 28.1430 14.6445 ;
      RECT 28.0170 10.9035 28.0350 14.6445 ;
      RECT 27.9090 10.9035 27.9270 14.6445 ;
      RECT 27.8010 10.9035 27.8190 14.6445 ;
      RECT 27.6930 10.9035 27.7110 14.6445 ;
      RECT 27.5850 10.9035 27.6030 14.6445 ;
      RECT 27.4770 10.9035 27.4950 14.6445 ;
      RECT 27.3690 10.9035 27.3870 14.6445 ;
      RECT 27.2610 10.9035 27.2790 14.6445 ;
      RECT 27.1530 10.9035 27.1710 14.6445 ;
      RECT 27.0450 10.9035 27.0630 14.6445 ;
      RECT 26.9370 10.9035 26.9550 14.6445 ;
      RECT 26.8290 10.9035 26.8470 14.6445 ;
      RECT 26.7210 10.9035 26.7390 14.6445 ;
      RECT 26.6130 10.9035 26.6310 14.6445 ;
      RECT 26.5050 10.9035 26.5230 14.6445 ;
      RECT 26.3970 10.9035 26.4150 14.6445 ;
      RECT 26.2890 10.9035 26.3070 14.6445 ;
      RECT 26.1810 10.9035 26.1990 14.6445 ;
      RECT 26.0730 10.9035 26.0910 14.6445 ;
      RECT 25.9650 10.9035 25.9830 14.6445 ;
      RECT 25.8570 10.9035 25.8750 14.6445 ;
      RECT 25.7490 10.9035 25.7670 14.6445 ;
      RECT 25.6410 10.9035 25.6590 14.6445 ;
      RECT 25.5330 10.9035 25.5510 14.6445 ;
      RECT 25.4250 10.9035 25.4430 14.6445 ;
      RECT 25.3170 10.9035 25.3350 14.6445 ;
      RECT 25.2090 10.9035 25.2270 14.6445 ;
      RECT 25.1010 10.9035 25.1190 14.6445 ;
      RECT 24.9930 10.9035 25.0110 14.6445 ;
      RECT 24.8850 10.9035 24.9030 14.6445 ;
      RECT 24.7770 10.9035 24.7950 14.6445 ;
      RECT 24.6690 10.9035 24.6870 14.6445 ;
      RECT 24.5610 10.9035 24.5790 14.6445 ;
      RECT 24.4530 10.9035 24.4710 14.6445 ;
      RECT 24.3450 10.9035 24.3630 14.6445 ;
      RECT 24.2370 10.9035 24.2550 14.6445 ;
      RECT 24.1290 10.9035 24.1470 14.6445 ;
      RECT 24.0210 10.9035 24.0390 14.6445 ;
      RECT 23.9130 10.9035 23.9310 14.6445 ;
      RECT 23.8050 10.9035 23.8230 14.6445 ;
      RECT 23.6970 10.9035 23.7150 14.6445 ;
      RECT 23.5890 10.9035 23.6070 14.6445 ;
      RECT 23.4810 10.9035 23.4990 14.6445 ;
      RECT 23.3730 10.9035 23.3910 14.6445 ;
      RECT 23.2650 10.9035 23.2830 14.6445 ;
      RECT 23.1570 10.9035 23.1750 14.6445 ;
      RECT 23.0490 10.9035 23.0670 14.6445 ;
      RECT 22.9410 10.9035 22.9590 14.6445 ;
      RECT 22.8330 10.9035 22.8510 14.6445 ;
      RECT 22.7250 10.9035 22.7430 14.6445 ;
      RECT 22.6170 10.9035 22.6350 14.6445 ;
      RECT 22.5090 10.9035 22.5270 14.6445 ;
      RECT 22.4010 10.9035 22.4190 14.6445 ;
      RECT 22.2930 10.9035 22.3110 14.6445 ;
      RECT 22.1850 10.9035 22.2030 14.6445 ;
      RECT 22.0770 10.9035 22.0950 14.6445 ;
      RECT 21.9690 10.9035 21.9870 14.6445 ;
      RECT 21.8610 10.9035 21.8790 14.6445 ;
      RECT 21.7530 10.9035 21.7710 14.6445 ;
      RECT 21.6450 10.9035 21.6630 14.6445 ;
      RECT 21.5370 10.9035 21.5550 14.6445 ;
      RECT 21.4290 10.9035 21.4470 14.6445 ;
      RECT 21.3210 10.9035 21.3390 14.6445 ;
      RECT 21.2130 10.9035 21.2310 14.6445 ;
      RECT 21.1050 10.9035 21.1230 14.6445 ;
      RECT 20.9970 10.9035 21.0150 14.6445 ;
      RECT 20.8890 10.9035 20.9070 14.6445 ;
      RECT 20.7810 10.9035 20.7990 14.6445 ;
      RECT 20.6730 10.9035 20.6910 14.6445 ;
      RECT 20.5650 10.9035 20.5830 14.6445 ;
      RECT 20.4570 10.9035 20.4750 14.6445 ;
      RECT 20.3490 10.9035 20.3670 14.6445 ;
      RECT 20.2410 10.9035 20.2590 14.6445 ;
      RECT 20.1330 10.9035 20.1510 14.6445 ;
      RECT 20.0250 10.9035 20.0430 14.6445 ;
      RECT 19.9170 10.9035 19.9350 14.6445 ;
      RECT 19.8090 11.0670 19.8270 11.4170 ;
      RECT 19.7010 10.9035 19.7190 14.6445 ;
      RECT 19.5930 10.9035 19.6110 14.6445 ;
      RECT 19.4850 10.9035 19.5030 14.6445 ;
      RECT 19.3770 10.9035 19.3950 14.6445 ;
      RECT 19.2690 10.9035 19.2870 14.6445 ;
      RECT 19.1610 10.9035 19.1790 14.6445 ;
      RECT 19.0530 10.9035 19.0710 14.6445 ;
      RECT 18.9450 10.9035 18.9630 14.6445 ;
      RECT 18.8370 10.9035 18.8550 14.6445 ;
      RECT 18.7290 10.9035 18.7470 14.6445 ;
      RECT 18.6210 10.9035 18.6390 14.6445 ;
      RECT 18.5130 10.9035 18.5310 14.6445 ;
      RECT 18.4050 10.9035 18.4230 14.6445 ;
      RECT 18.2970 10.9035 18.3150 14.6445 ;
      RECT 18.1890 10.9035 18.2070 14.6445 ;
      RECT 18.0810 10.9035 18.0990 14.6445 ;
      RECT 17.9730 10.9035 17.9910 14.6445 ;
      RECT 17.8650 10.9035 17.8830 14.6445 ;
      RECT 17.7570 10.9035 17.7750 14.6445 ;
      RECT 17.6490 10.9035 17.6670 14.6445 ;
      RECT 17.5410 10.9035 17.5590 14.6445 ;
      RECT 17.4330 10.9035 17.4510 14.6445 ;
      RECT 17.3250 10.9035 17.3430 14.6445 ;
      RECT 17.2170 10.9035 17.2350 14.6445 ;
      RECT 17.1090 10.9035 17.1270 14.6445 ;
      RECT 17.0010 10.9035 17.0190 14.6445 ;
      RECT 16.8930 10.9035 16.9110 14.6445 ;
      RECT 16.7850 10.9035 16.8030 14.6445 ;
      RECT 16.6770 10.9035 16.6950 14.6445 ;
      RECT 16.5690 10.9035 16.5870 14.6445 ;
      RECT 16.4610 10.9035 16.4790 14.6445 ;
      RECT 16.4250 14.8555 16.4430 15.5602 ;
      RECT 16.4250 16.2985 16.4430 17.4595 ;
      RECT 16.4070 11.7275 16.4250 12.4035 ;
      RECT 16.4070 13.1495 16.4250 13.4475 ;
      RECT 16.4070 14.2655 16.4250 14.5275 ;
      RECT 16.3890 14.9190 16.4070 15.6090 ;
      RECT 16.3890 15.6600 16.4070 16.6455 ;
      RECT 16.3890 16.6865 16.4070 17.3035 ;
      RECT 16.3530 10.9035 16.3710 19.2740 ;
      RECT 16.3170 15.1915 16.3350 15.2745 ;
      RECT 16.2990 11.8355 16.3170 12.4665 ;
      RECT 16.2990 12.8795 16.3170 13.0695 ;
      RECT 16.2990 13.7615 16.3170 13.8105 ;
      RECT 16.2990 14.4935 16.3170 14.5305 ;
      RECT 16.2810 14.8865 16.2990 18.4795 ;
      RECT 16.1910 11.1000 16.2090 11.2380 ;
      RECT 16.1910 11.4575 16.2090 12.2595 ;
      RECT 16.1910 12.8075 16.2090 13.3755 ;
      RECT 16.1910 14.8865 16.2090 18.4795 ;
      RECT 16.1550 12.8795 16.1730 13.2495 ;
      RECT 16.1190 12.2315 16.1370 12.3675 ;
      RECT 16.1190 13.2215 16.1370 13.4475 ;
      RECT 16.1190 14.4635 16.1370 14.5275 ;
      RECT 16.0830 12.3335 16.1010 12.3705 ;
      RECT 16.0830 13.9595 16.1010 14.0025 ;
      RECT 16.0830 14.4935 16.1010 14.5305 ;
      RECT 16.0470 12.6455 16.0650 13.1415 ;
      RECT 16.0470 13.1855 16.0650 13.3755 ;
      RECT 16.0470 14.1455 16.0650 14.4555 ;
      RECT 16.0110 12.5375 16.0290 13.7845 ;
      RECT 15.0390 11.0935 15.0570 11.2475 ;
      RECT 15.0030 11.0935 15.0210 11.1435 ;
      RECT 14.9310 11.0935 14.9490 11.1650 ;
      RECT 14.2830 12.2315 14.3010 12.6375 ;
      RECT 14.2470 13.3415 14.2650 13.3785 ;
      RECT 14.2110 12.2675 14.2290 12.8715 ;
      RECT 14.1750 12.1055 14.1930 12.1695 ;
      RECT 14.1390 11.1465 14.1570 11.1975 ;
      RECT 14.1390 14.2655 14.1570 14.4555 ;
      RECT 14.1390 14.8865 14.1570 18.4795 ;
      RECT 14.0310 11.5655 14.0490 11.7555 ;
      RECT 14.0310 12.3395 14.0490 14.5995 ;
      RECT 14.0130 15.1915 14.0310 15.2745 ;
      RECT 13.9770 11.0670 13.9950 19.2740 ;
      RECT 13.9410 14.9190 13.9590 15.6090 ;
      RECT 13.9410 15.6600 13.9590 16.6455 ;
      RECT 13.9410 16.6865 13.9590 17.3035 ;
      RECT 13.9230 11.5655 13.9410 12.0615 ;
      RECT 13.9230 12.8435 13.9410 13.4115 ;
      RECT 13.9230 13.7255 13.9410 14.4555 ;
      RECT 13.9050 14.8555 13.9230 15.5602 ;
      RECT 13.9050 16.2985 13.9230 17.4595 ;
      RECT 13.8690 11.0670 13.8870 11.4170 ;
      RECT 13.8690 14.6110 13.8870 19.2740 ;
      RECT 13.7610 11.0670 13.7790 11.4170 ;
      RECT 13.6530 11.0670 13.6710 11.4170 ;
      RECT 13.5450 11.0670 13.5630 11.4170 ;
      RECT 13.4370 11.0670 13.4550 11.4170 ;
      RECT 13.3290 11.0670 13.3470 11.4170 ;
      RECT 13.2210 11.0670 13.2390 11.4170 ;
      RECT 13.1130 11.0670 13.1310 11.4170 ;
      RECT 13.0050 11.0670 13.0230 11.4170 ;
      RECT 12.8970 11.0670 12.9150 11.4170 ;
      RECT 12.7890 11.0670 12.8070 11.4170 ;
      RECT 12.6810 11.0670 12.6990 11.4170 ;
      RECT 12.5730 11.0670 12.5910 11.4170 ;
      RECT 12.4650 11.0670 12.4830 11.4170 ;
      RECT 12.3570 11.0670 12.3750 11.4170 ;
      RECT 12.2490 11.0670 12.2670 11.4170 ;
      RECT 12.1410 11.0670 12.1590 11.4170 ;
      RECT 12.0330 11.0670 12.0510 11.4170 ;
      RECT 11.9250 11.0670 11.9430 11.4170 ;
      RECT 11.8170 11.0670 11.8350 11.4170 ;
      RECT 11.7090 11.0670 11.7270 11.4170 ;
      RECT 11.6010 11.0670 11.6190 11.4170 ;
      RECT 11.4930 11.0670 11.5110 11.4170 ;
      RECT 11.3850 11.0670 11.4030 11.4170 ;
      RECT 11.2770 11.0670 11.2950 11.4170 ;
      RECT 11.1690 11.0670 11.1870 11.4170 ;
      RECT 11.0610 11.0670 11.0790 11.4170 ;
      RECT 10.9530 11.0670 10.9710 11.4170 ;
      RECT 10.8450 11.0670 10.8630 11.4170 ;
      RECT 10.7370 11.0670 10.7550 11.4170 ;
      RECT 10.6290 11.0670 10.6470 11.4170 ;
      RECT 10.5210 11.0670 10.5390 11.4170 ;
      RECT 10.4130 11.0670 10.4310 11.4170 ;
      RECT 10.3050 11.0670 10.3230 11.4170 ;
      RECT 10.1970 11.0670 10.2150 11.4170 ;
      RECT 10.0890 11.0670 10.1070 11.4170 ;
      RECT 9.9810 11.0670 9.9990 11.4170 ;
      RECT 9.8730 11.0670 9.8910 11.4170 ;
      RECT 9.7650 11.0670 9.7830 11.4170 ;
      RECT 9.6570 11.0670 9.6750 11.4170 ;
      RECT 9.5490 11.0670 9.5670 11.4170 ;
      RECT 9.4410 11.0670 9.4590 11.4170 ;
      RECT 9.3330 11.0670 9.3510 11.4170 ;
      RECT 9.2250 11.0670 9.2430 11.4170 ;
      RECT 9.1170 11.0670 9.1350 11.4170 ;
      RECT 9.0090 11.0670 9.0270 11.4170 ;
      RECT 8.9010 11.0670 8.9190 11.4170 ;
      RECT 8.7930 11.0670 8.8110 11.4170 ;
      RECT 8.6850 11.0670 8.7030 11.4170 ;
      RECT 8.5770 11.0670 8.5950 11.4170 ;
      RECT 8.4690 11.0670 8.4870 11.4170 ;
      RECT 8.3610 11.0670 8.3790 11.4170 ;
      RECT 8.2530 11.0670 8.2710 11.4170 ;
      RECT 8.1450 11.0670 8.1630 11.4170 ;
      RECT 8.0370 11.0670 8.0550 11.4170 ;
      RECT 7.9290 11.0670 7.9470 11.4170 ;
      RECT 7.8210 11.0670 7.8390 11.4170 ;
      RECT 7.7130 11.0670 7.7310 11.4170 ;
      RECT 7.6050 11.0670 7.6230 11.4170 ;
      RECT 7.4970 11.0670 7.5150 11.4170 ;
      RECT 7.3890 11.0670 7.4070 11.4170 ;
      RECT 7.2810 11.0670 7.2990 11.4170 ;
      RECT 7.1730 11.0670 7.1910 11.4170 ;
      RECT 7.0650 11.0670 7.0830 11.4170 ;
      RECT 6.9570 11.0670 6.9750 11.4170 ;
      RECT 6.8490 11.0670 6.8670 11.4170 ;
      RECT 6.7410 11.0670 6.7590 11.4170 ;
      RECT 6.6330 11.0670 6.6510 11.4170 ;
      RECT 6.5250 11.0670 6.5430 11.4170 ;
      RECT 6.4170 11.0670 6.4350 11.4170 ;
      RECT 6.3090 11.0670 6.3270 11.4170 ;
      RECT 6.2010 11.0670 6.2190 11.4170 ;
      RECT 6.0930 11.0670 6.1110 11.4170 ;
      RECT 5.9850 11.0670 6.0030 11.4170 ;
      RECT 5.8770 11.0670 5.8950 11.4170 ;
      RECT 5.7690 11.0670 5.7870 11.4170 ;
      RECT 5.6610 11.0670 5.6790 11.4170 ;
      RECT 5.5530 11.0670 5.5710 11.4170 ;
      RECT 5.4450 11.0670 5.4630 11.4170 ;
      RECT 5.3370 11.0670 5.3550 11.4170 ;
      RECT 5.2290 11.0670 5.2470 11.4170 ;
      RECT 5.1210 11.0670 5.1390 11.4170 ;
      RECT 5.0130 11.0670 5.0310 11.4170 ;
      RECT 4.9050 11.0670 4.9230 11.4170 ;
      RECT 4.7970 11.0670 4.8150 11.4170 ;
      RECT 4.6890 11.0670 4.7070 11.4170 ;
      RECT 4.5810 11.0670 4.5990 11.4170 ;
      RECT 4.4730 11.0670 4.4910 11.4170 ;
      RECT 4.3650 11.0670 4.3830 11.4170 ;
      RECT 4.2570 11.0670 4.2750 11.4170 ;
      RECT 4.1490 11.0670 4.1670 11.4170 ;
      RECT 4.0410 11.0670 4.0590 11.4170 ;
      RECT 3.9330 11.0670 3.9510 11.4170 ;
      RECT 3.8250 11.0670 3.8430 11.4170 ;
      RECT 3.7170 11.0670 3.7350 11.4170 ;
      RECT 3.6090 11.0670 3.6270 11.4170 ;
      RECT 3.5010 11.0670 3.5190 11.4170 ;
      RECT 3.3930 11.0670 3.4110 11.4170 ;
      RECT 3.2850 11.0670 3.3030 11.4170 ;
      RECT 3.1770 11.0670 3.1950 11.4170 ;
      RECT 3.0690 11.0670 3.0870 11.4170 ;
      RECT 2.9610 11.0670 2.9790 11.4170 ;
      RECT 2.8530 11.0670 2.8710 11.4170 ;
      RECT 2.7450 11.0670 2.7630 11.4170 ;
      RECT 2.6370 11.0670 2.6550 11.4170 ;
      RECT 2.5290 11.0670 2.5470 11.4170 ;
      RECT 2.4210 11.0670 2.4390 11.4170 ;
      RECT 2.3130 11.0670 2.3310 11.4170 ;
      RECT 2.2050 11.0670 2.2230 11.4170 ;
      RECT 2.0970 11.0670 2.1150 11.4170 ;
      RECT 1.9890 11.0670 2.0070 11.4170 ;
      RECT 1.8810 11.0670 1.8990 11.4170 ;
      RECT 1.7730 11.0670 1.7910 11.4170 ;
      RECT 1.6650 11.0670 1.6830 11.4170 ;
      RECT 1.5570 11.0670 1.5750 11.4170 ;
      RECT 1.4490 11.0670 1.4670 11.4170 ;
      RECT 1.3410 11.0670 1.3590 11.4170 ;
      RECT 1.2330 11.0670 1.2510 11.4170 ;
      RECT 1.1250 11.0670 1.1430 11.4170 ;
      RECT 1.0170 11.0670 1.0350 11.4170 ;
      RECT 0.9090 11.0670 0.9270 11.4170 ;
      RECT 0.8010 11.0670 0.8190 11.4170 ;
      RECT 0.6930 11.0670 0.7110 11.4170 ;
      RECT 0.5850 11.0670 0.6030 11.4170 ;
      RECT 0.4770 11.0670 0.4950 11.4170 ;
      RECT 0.3690 11.0670 0.3870 11.4170 ;
      RECT 0.2610 11.0670 0.2790 11.4170 ;
      RECT 0.1530 11.0670 0.1710 19.2740 ;
      RECT 0.1170 11.0670 0.1350 19.2740 ;
        RECT 15.6110 19.2720 15.6290 20.2075 ;
        RECT 15.5750 19.2720 15.5930 20.2075 ;
        RECT 15.5390 19.8490 15.5570 20.1715 ;
        RECT 15.4220 20.0460 15.4400 20.1555 ;
        RECT 15.4130 19.3045 15.4310 19.5440 ;
        RECT 15.3770 19.8855 15.3950 20.0390 ;
        RECT 15.2960 19.9110 15.3140 20.1690 ;
        RECT 14.7560 19.2720 14.7740 20.2075 ;
        RECT 14.7200 19.2720 14.7380 20.2075 ;
        RECT 14.6840 19.4530 14.7020 20.0210 ;
        RECT 15.6110 20.3520 15.6290 21.2875 ;
        RECT 15.5750 20.3520 15.5930 21.2875 ;
        RECT 15.5390 20.9290 15.5570 21.2515 ;
        RECT 15.4220 21.1260 15.4400 21.2355 ;
        RECT 15.4130 20.3845 15.4310 20.6240 ;
        RECT 15.3770 20.9655 15.3950 21.1190 ;
        RECT 15.2960 20.9910 15.3140 21.2490 ;
        RECT 14.7560 20.3520 14.7740 21.2875 ;
        RECT 14.7200 20.3520 14.7380 21.2875 ;
        RECT 14.6840 20.5330 14.7020 21.1010 ;
        RECT 15.6110 21.4320 15.6290 22.3675 ;
        RECT 15.5750 21.4320 15.5930 22.3675 ;
        RECT 15.5390 22.0090 15.5570 22.3315 ;
        RECT 15.4220 22.2060 15.4400 22.3155 ;
        RECT 15.4130 21.4645 15.4310 21.7040 ;
        RECT 15.3770 22.0455 15.3950 22.1990 ;
        RECT 15.2960 22.0710 15.3140 22.3290 ;
        RECT 14.7560 21.4320 14.7740 22.3675 ;
        RECT 14.7200 21.4320 14.7380 22.3675 ;
        RECT 14.6840 21.6130 14.7020 22.1810 ;
        RECT 15.6110 22.5120 15.6290 23.4475 ;
        RECT 15.5750 22.5120 15.5930 23.4475 ;
        RECT 15.5390 23.0890 15.5570 23.4115 ;
        RECT 15.4220 23.2860 15.4400 23.3955 ;
        RECT 15.4130 22.5445 15.4310 22.7840 ;
        RECT 15.3770 23.1255 15.3950 23.2790 ;
        RECT 15.2960 23.1510 15.3140 23.4090 ;
        RECT 14.7560 22.5120 14.7740 23.4475 ;
        RECT 14.7200 22.5120 14.7380 23.4475 ;
        RECT 14.6840 22.6930 14.7020 23.2610 ;
        RECT 15.6110 23.5920 15.6290 24.5275 ;
        RECT 15.5750 23.5920 15.5930 24.5275 ;
        RECT 15.5390 24.1690 15.5570 24.4915 ;
        RECT 15.4220 24.3660 15.4400 24.4755 ;
        RECT 15.4130 23.6245 15.4310 23.8640 ;
        RECT 15.3770 24.2055 15.3950 24.3590 ;
        RECT 15.2960 24.2310 15.3140 24.4890 ;
        RECT 14.7560 23.5920 14.7740 24.5275 ;
        RECT 14.7200 23.5920 14.7380 24.5275 ;
        RECT 14.6840 23.7730 14.7020 24.3410 ;
        RECT 15.6110 24.6720 15.6290 25.6075 ;
        RECT 15.5750 24.6720 15.5930 25.6075 ;
        RECT 15.5390 25.2490 15.5570 25.5715 ;
        RECT 15.4220 25.4460 15.4400 25.5555 ;
        RECT 15.4130 24.7045 15.4310 24.9440 ;
        RECT 15.3770 25.2855 15.3950 25.4390 ;
        RECT 15.2960 25.3110 15.3140 25.5690 ;
        RECT 14.7560 24.6720 14.7740 25.6075 ;
        RECT 14.7200 24.6720 14.7380 25.6075 ;
        RECT 14.6840 24.8530 14.7020 25.4210 ;
        RECT 15.6110 25.7520 15.6290 26.6875 ;
        RECT 15.5750 25.7520 15.5930 26.6875 ;
        RECT 15.5390 26.3290 15.5570 26.6515 ;
        RECT 15.4220 26.5260 15.4400 26.6355 ;
        RECT 15.4130 25.7845 15.4310 26.0240 ;
        RECT 15.3770 26.3655 15.3950 26.5190 ;
        RECT 15.2960 26.3910 15.3140 26.6490 ;
        RECT 14.7560 25.7520 14.7740 26.6875 ;
        RECT 14.7200 25.7520 14.7380 26.6875 ;
        RECT 14.6840 25.9330 14.7020 26.5010 ;
        RECT 15.6110 26.8320 15.6290 27.7675 ;
        RECT 15.5750 26.8320 15.5930 27.7675 ;
        RECT 15.5390 27.4090 15.5570 27.7315 ;
        RECT 15.4220 27.6060 15.4400 27.7155 ;
        RECT 15.4130 26.8645 15.4310 27.1040 ;
        RECT 15.3770 27.4455 15.3950 27.5990 ;
        RECT 15.2960 27.4710 15.3140 27.7290 ;
        RECT 14.7560 26.8320 14.7740 27.7675 ;
        RECT 14.7200 26.8320 14.7380 27.7675 ;
        RECT 14.6840 27.0130 14.7020 27.5810 ;
        RECT 15.6110 27.9120 15.6290 28.8475 ;
        RECT 15.5750 27.9120 15.5930 28.8475 ;
        RECT 15.5390 28.4890 15.5570 28.8115 ;
        RECT 15.4220 28.6860 15.4400 28.7955 ;
        RECT 15.4130 27.9445 15.4310 28.1840 ;
        RECT 15.3770 28.5255 15.3950 28.6790 ;
        RECT 15.2960 28.5510 15.3140 28.8090 ;
        RECT 14.7560 27.9120 14.7740 28.8475 ;
        RECT 14.7200 27.9120 14.7380 28.8475 ;
        RECT 14.6840 28.0930 14.7020 28.6610 ;
        RECT 15.6110 28.9920 15.6290 29.9275 ;
        RECT 15.5750 28.9920 15.5930 29.9275 ;
        RECT 15.5390 29.5690 15.5570 29.8915 ;
        RECT 15.4220 29.7660 15.4400 29.8755 ;
        RECT 15.4130 29.0245 15.4310 29.2640 ;
        RECT 15.3770 29.6055 15.3950 29.7590 ;
        RECT 15.2960 29.6310 15.3140 29.8890 ;
        RECT 14.7560 28.9920 14.7740 29.9275 ;
        RECT 14.7200 28.9920 14.7380 29.9275 ;
        RECT 14.6840 29.1730 14.7020 29.7410 ;
  LAYER M3 SPACING 0.018  ;
      RECT 15.5530 0.2565 15.6810 1.3500 ;
      RECT 15.5390 0.9220 15.6810 1.2445 ;
      RECT 15.3190 0.6490 15.4530 1.3500 ;
      RECT 15.2960 0.9840 15.4530 1.2420 ;
      RECT 15.3190 0.2565 15.4170 1.3500 ;
      RECT 15.3190 0.3775 15.4310 0.6170 ;
      RECT 15.3190 0.2565 15.4530 0.3455 ;
      RECT 15.0940 0.7070 15.2280 1.3500 ;
      RECT 15.0940 0.2565 15.1920 1.3500 ;
      RECT 14.6770 0.2565 14.7600 1.3500 ;
      RECT 14.6770 0.3450 14.7740 1.2805 ;
      RECT 30.2680 0.2565 30.3530 1.3500 ;
      RECT 30.1240 0.2565 30.1500 1.3500 ;
      RECT 30.0160 0.2565 30.0420 1.3500 ;
      RECT 29.9080 0.2565 29.9340 1.3500 ;
      RECT 29.8000 0.2565 29.8260 1.3500 ;
      RECT 29.6920 0.2565 29.7180 1.3500 ;
      RECT 29.5840 0.2565 29.6100 1.3500 ;
      RECT 29.4760 0.2565 29.5020 1.3500 ;
      RECT 29.3680 0.2565 29.3940 1.3500 ;
      RECT 29.2600 0.2565 29.2860 1.3500 ;
      RECT 29.1520 0.2565 29.1780 1.3500 ;
      RECT 29.0440 0.2565 29.0700 1.3500 ;
      RECT 28.9360 0.2565 28.9620 1.3500 ;
      RECT 28.8280 0.2565 28.8540 1.3500 ;
      RECT 28.7200 0.2565 28.7460 1.3500 ;
      RECT 28.6120 0.2565 28.6380 1.3500 ;
      RECT 28.5040 0.2565 28.5300 1.3500 ;
      RECT 28.3960 0.2565 28.4220 1.3500 ;
      RECT 28.2880 0.2565 28.3140 1.3500 ;
      RECT 28.1800 0.2565 28.2060 1.3500 ;
      RECT 28.0720 0.2565 28.0980 1.3500 ;
      RECT 27.9640 0.2565 27.9900 1.3500 ;
      RECT 27.8560 0.2565 27.8820 1.3500 ;
      RECT 27.7480 0.2565 27.7740 1.3500 ;
      RECT 27.6400 0.2565 27.6660 1.3500 ;
      RECT 27.5320 0.2565 27.5580 1.3500 ;
      RECT 27.4240 0.2565 27.4500 1.3500 ;
      RECT 27.3160 0.2565 27.3420 1.3500 ;
      RECT 27.2080 0.2565 27.2340 1.3500 ;
      RECT 27.1000 0.2565 27.1260 1.3500 ;
      RECT 26.9920 0.2565 27.0180 1.3500 ;
      RECT 26.8840 0.2565 26.9100 1.3500 ;
      RECT 26.7760 0.2565 26.8020 1.3500 ;
      RECT 26.6680 0.2565 26.6940 1.3500 ;
      RECT 26.5600 0.2565 26.5860 1.3500 ;
      RECT 26.4520 0.2565 26.4780 1.3500 ;
      RECT 26.3440 0.2565 26.3700 1.3500 ;
      RECT 26.2360 0.2565 26.2620 1.3500 ;
      RECT 26.1280 0.2565 26.1540 1.3500 ;
      RECT 26.0200 0.2565 26.0460 1.3500 ;
      RECT 25.9120 0.2565 25.9380 1.3500 ;
      RECT 25.8040 0.2565 25.8300 1.3500 ;
      RECT 25.6960 0.2565 25.7220 1.3500 ;
      RECT 25.5880 0.2565 25.6140 1.3500 ;
      RECT 25.4800 0.2565 25.5060 1.3500 ;
      RECT 25.3720 0.2565 25.3980 1.3500 ;
      RECT 25.2640 0.2565 25.2900 1.3500 ;
      RECT 25.1560 0.2565 25.1820 1.3500 ;
      RECT 25.0480 0.2565 25.0740 1.3500 ;
      RECT 24.9400 0.2565 24.9660 1.3500 ;
      RECT 24.8320 0.2565 24.8580 1.3500 ;
      RECT 24.7240 0.2565 24.7500 1.3500 ;
      RECT 24.6160 0.2565 24.6420 1.3500 ;
      RECT 24.5080 0.2565 24.5340 1.3500 ;
      RECT 24.4000 0.2565 24.4260 1.3500 ;
      RECT 24.2920 0.2565 24.3180 1.3500 ;
      RECT 24.1840 0.2565 24.2100 1.3500 ;
      RECT 24.0760 0.2565 24.1020 1.3500 ;
      RECT 23.9680 0.2565 23.9940 1.3500 ;
      RECT 23.8600 0.2565 23.8860 1.3500 ;
      RECT 23.7520 0.2565 23.7780 1.3500 ;
      RECT 23.6440 0.2565 23.6700 1.3500 ;
      RECT 23.5360 0.2565 23.5620 1.3500 ;
      RECT 23.4280 0.2565 23.4540 1.3500 ;
      RECT 23.3200 0.2565 23.3460 1.3500 ;
      RECT 23.2120 0.2565 23.2380 1.3500 ;
      RECT 23.1040 0.2565 23.1300 1.3500 ;
      RECT 22.9960 0.2565 23.0220 1.3500 ;
      RECT 22.8880 0.2565 22.9140 1.3500 ;
      RECT 22.7800 0.2565 22.8060 1.3500 ;
      RECT 22.6720 0.2565 22.6980 1.3500 ;
      RECT 22.5640 0.2565 22.5900 1.3500 ;
      RECT 22.4560 0.2565 22.4820 1.3500 ;
      RECT 22.3480 0.2565 22.3740 1.3500 ;
      RECT 22.2400 0.2565 22.2660 1.3500 ;
      RECT 22.1320 0.2565 22.1580 1.3500 ;
      RECT 22.0240 0.2565 22.0500 1.3500 ;
      RECT 21.9160 0.2565 21.9420 1.3500 ;
      RECT 21.8080 0.2565 21.8340 1.3500 ;
      RECT 21.7000 0.2565 21.7260 1.3500 ;
      RECT 21.5920 0.2565 21.6180 1.3500 ;
      RECT 21.4840 0.2565 21.5100 1.3500 ;
      RECT 21.3760 0.2565 21.4020 1.3500 ;
      RECT 21.2680 0.2565 21.2940 1.3500 ;
      RECT 21.1600 0.2565 21.1860 1.3500 ;
      RECT 21.0520 0.2565 21.0780 1.3500 ;
      RECT 20.9440 0.2565 20.9700 1.3500 ;
      RECT 20.8360 0.2565 20.8620 1.3500 ;
      RECT 20.7280 0.2565 20.7540 1.3500 ;
      RECT 20.6200 0.2565 20.6460 1.3500 ;
      RECT 20.5120 0.2565 20.5380 1.3500 ;
      RECT 20.4040 0.2565 20.4300 1.3500 ;
      RECT 20.2960 0.2565 20.3220 1.3500 ;
      RECT 20.1880 0.2565 20.2140 1.3500 ;
      RECT 20.0800 0.2565 20.1060 1.3500 ;
      RECT 19.9720 0.2565 19.9980 1.3500 ;
      RECT 19.8640 0.2565 19.8900 1.3500 ;
      RECT 19.7560 0.2565 19.7820 1.3500 ;
      RECT 19.6480 0.2565 19.6740 1.3500 ;
      RECT 19.5400 0.2565 19.5660 1.3500 ;
      RECT 19.4320 0.2565 19.4580 1.3500 ;
      RECT 19.3240 0.2565 19.3500 1.3500 ;
      RECT 19.2160 0.2565 19.2420 1.3500 ;
      RECT 19.1080 0.2565 19.1340 1.3500 ;
      RECT 19.0000 0.2565 19.0260 1.3500 ;
      RECT 18.8920 0.2565 18.9180 1.3500 ;
      RECT 18.7840 0.2565 18.8100 1.3500 ;
      RECT 18.6760 0.2565 18.7020 1.3500 ;
      RECT 18.5680 0.2565 18.5940 1.3500 ;
      RECT 18.4600 0.2565 18.4860 1.3500 ;
      RECT 18.3520 0.2565 18.3780 1.3500 ;
      RECT 18.2440 0.2565 18.2700 1.3500 ;
      RECT 18.1360 0.2565 18.1620 1.3500 ;
      RECT 18.0280 0.2565 18.0540 1.3500 ;
      RECT 17.9200 0.2565 17.9460 1.3500 ;
      RECT 17.8120 0.2565 17.8380 1.3500 ;
      RECT 17.7040 0.2565 17.7300 1.3500 ;
      RECT 17.5960 0.2565 17.6220 1.3500 ;
      RECT 17.4880 0.2565 17.5140 1.3500 ;
      RECT 17.3800 0.2565 17.4060 1.3500 ;
      RECT 17.2720 0.2565 17.2980 1.3500 ;
      RECT 17.1640 0.2565 17.1900 1.3500 ;
      RECT 17.0560 0.2565 17.0820 1.3500 ;
      RECT 16.9480 0.2565 16.9740 1.3500 ;
      RECT 16.8400 0.2565 16.8660 1.3500 ;
      RECT 16.7320 0.2565 16.7580 1.3500 ;
      RECT 16.6240 0.2565 16.6500 1.3500 ;
      RECT 16.5160 0.2565 16.5420 1.3500 ;
      RECT 16.4080 0.2565 16.4340 1.3500 ;
      RECT 16.3000 0.2565 16.3260 1.3500 ;
      RECT 16.0870 0.2565 16.1640 1.3500 ;
      RECT 14.1940 0.2565 14.2710 1.3500 ;
      RECT 14.0320 0.2565 14.0580 1.3500 ;
      RECT 13.9240 0.2565 13.9500 1.3500 ;
      RECT 13.8160 0.2565 13.8420 1.3500 ;
      RECT 13.7080 0.2565 13.7340 1.3500 ;
      RECT 13.6000 0.2565 13.6260 1.3500 ;
      RECT 13.4920 0.2565 13.5180 1.3500 ;
      RECT 13.3840 0.2565 13.4100 1.3500 ;
      RECT 13.2760 0.2565 13.3020 1.3500 ;
      RECT 13.1680 0.2565 13.1940 1.3500 ;
      RECT 13.0600 0.2565 13.0860 1.3500 ;
      RECT 12.9520 0.2565 12.9780 1.3500 ;
      RECT 12.8440 0.2565 12.8700 1.3500 ;
      RECT 12.7360 0.2565 12.7620 1.3500 ;
      RECT 12.6280 0.2565 12.6540 1.3500 ;
      RECT 12.5200 0.2565 12.5460 1.3500 ;
      RECT 12.4120 0.2565 12.4380 1.3500 ;
      RECT 12.3040 0.2565 12.3300 1.3500 ;
      RECT 12.1960 0.2565 12.2220 1.3500 ;
      RECT 12.0880 0.2565 12.1140 1.3500 ;
      RECT 11.9800 0.2565 12.0060 1.3500 ;
      RECT 11.8720 0.2565 11.8980 1.3500 ;
      RECT 11.7640 0.2565 11.7900 1.3500 ;
      RECT 11.6560 0.2565 11.6820 1.3500 ;
      RECT 11.5480 0.2565 11.5740 1.3500 ;
      RECT 11.4400 0.2565 11.4660 1.3500 ;
      RECT 11.3320 0.2565 11.3580 1.3500 ;
      RECT 11.2240 0.2565 11.2500 1.3500 ;
      RECT 11.1160 0.2565 11.1420 1.3500 ;
      RECT 11.0080 0.2565 11.0340 1.3500 ;
      RECT 10.9000 0.2565 10.9260 1.3500 ;
      RECT 10.7920 0.2565 10.8180 1.3500 ;
      RECT 10.6840 0.2565 10.7100 1.3500 ;
      RECT 10.5760 0.2565 10.6020 1.3500 ;
      RECT 10.4680 0.2565 10.4940 1.3500 ;
      RECT 10.3600 0.2565 10.3860 1.3500 ;
      RECT 10.2520 0.2565 10.2780 1.3500 ;
      RECT 10.1440 0.2565 10.1700 1.3500 ;
      RECT 10.0360 0.2565 10.0620 1.3500 ;
      RECT 9.9280 0.2565 9.9540 1.3500 ;
      RECT 9.8200 0.2565 9.8460 1.3500 ;
      RECT 9.7120 0.2565 9.7380 1.3500 ;
      RECT 9.6040 0.2565 9.6300 1.3500 ;
      RECT 9.4960 0.2565 9.5220 1.3500 ;
      RECT 9.3880 0.2565 9.4140 1.3500 ;
      RECT 9.2800 0.2565 9.3060 1.3500 ;
      RECT 9.1720 0.2565 9.1980 1.3500 ;
      RECT 9.0640 0.2565 9.0900 1.3500 ;
      RECT 8.9560 0.2565 8.9820 1.3500 ;
      RECT 8.8480 0.2565 8.8740 1.3500 ;
      RECT 8.7400 0.2565 8.7660 1.3500 ;
      RECT 8.6320 0.2565 8.6580 1.3500 ;
      RECT 8.5240 0.2565 8.5500 1.3500 ;
      RECT 8.4160 0.2565 8.4420 1.3500 ;
      RECT 8.3080 0.2565 8.3340 1.3500 ;
      RECT 8.2000 0.2565 8.2260 1.3500 ;
      RECT 8.0920 0.2565 8.1180 1.3500 ;
      RECT 7.9840 0.2565 8.0100 1.3500 ;
      RECT 7.8760 0.2565 7.9020 1.3500 ;
      RECT 7.7680 0.2565 7.7940 1.3500 ;
      RECT 7.6600 0.2565 7.6860 1.3500 ;
      RECT 7.5520 0.2565 7.5780 1.3500 ;
      RECT 7.4440 0.2565 7.4700 1.3500 ;
      RECT 7.3360 0.2565 7.3620 1.3500 ;
      RECT 7.2280 0.2565 7.2540 1.3500 ;
      RECT 7.1200 0.2565 7.1460 1.3500 ;
      RECT 7.0120 0.2565 7.0380 1.3500 ;
      RECT 6.9040 0.2565 6.9300 1.3500 ;
      RECT 6.7960 0.2565 6.8220 1.3500 ;
      RECT 6.6880 0.2565 6.7140 1.3500 ;
      RECT 6.5800 0.2565 6.6060 1.3500 ;
      RECT 6.4720 0.2565 6.4980 1.3500 ;
      RECT 6.3640 0.2565 6.3900 1.3500 ;
      RECT 6.2560 0.2565 6.2820 1.3500 ;
      RECT 6.1480 0.2565 6.1740 1.3500 ;
      RECT 6.0400 0.2565 6.0660 1.3500 ;
      RECT 5.9320 0.2565 5.9580 1.3500 ;
      RECT 5.8240 0.2565 5.8500 1.3500 ;
      RECT 5.7160 0.2565 5.7420 1.3500 ;
      RECT 5.6080 0.2565 5.6340 1.3500 ;
      RECT 5.5000 0.2565 5.5260 1.3500 ;
      RECT 5.3920 0.2565 5.4180 1.3500 ;
      RECT 5.2840 0.2565 5.3100 1.3500 ;
      RECT 5.1760 0.2565 5.2020 1.3500 ;
      RECT 5.0680 0.2565 5.0940 1.3500 ;
      RECT 4.9600 0.2565 4.9860 1.3500 ;
      RECT 4.8520 0.2565 4.8780 1.3500 ;
      RECT 4.7440 0.2565 4.7700 1.3500 ;
      RECT 4.6360 0.2565 4.6620 1.3500 ;
      RECT 4.5280 0.2565 4.5540 1.3500 ;
      RECT 4.4200 0.2565 4.4460 1.3500 ;
      RECT 4.3120 0.2565 4.3380 1.3500 ;
      RECT 4.2040 0.2565 4.2300 1.3500 ;
      RECT 4.0960 0.2565 4.1220 1.3500 ;
      RECT 3.9880 0.2565 4.0140 1.3500 ;
      RECT 3.8800 0.2565 3.9060 1.3500 ;
      RECT 3.7720 0.2565 3.7980 1.3500 ;
      RECT 3.6640 0.2565 3.6900 1.3500 ;
      RECT 3.5560 0.2565 3.5820 1.3500 ;
      RECT 3.4480 0.2565 3.4740 1.3500 ;
      RECT 3.3400 0.2565 3.3660 1.3500 ;
      RECT 3.2320 0.2565 3.2580 1.3500 ;
      RECT 3.1240 0.2565 3.1500 1.3500 ;
      RECT 3.0160 0.2565 3.0420 1.3500 ;
      RECT 2.9080 0.2565 2.9340 1.3500 ;
      RECT 2.8000 0.2565 2.8260 1.3500 ;
      RECT 2.6920 0.2565 2.7180 1.3500 ;
      RECT 2.5840 0.2565 2.6100 1.3500 ;
      RECT 2.4760 0.2565 2.5020 1.3500 ;
      RECT 2.3680 0.2565 2.3940 1.3500 ;
      RECT 2.2600 0.2565 2.2860 1.3500 ;
      RECT 2.1520 0.2565 2.1780 1.3500 ;
      RECT 2.0440 0.2565 2.0700 1.3500 ;
      RECT 1.9360 0.2565 1.9620 1.3500 ;
      RECT 1.8280 0.2565 1.8540 1.3500 ;
      RECT 1.7200 0.2565 1.7460 1.3500 ;
      RECT 1.6120 0.2565 1.6380 1.3500 ;
      RECT 1.5040 0.2565 1.5300 1.3500 ;
      RECT 1.3960 0.2565 1.4220 1.3500 ;
      RECT 1.2880 0.2565 1.3140 1.3500 ;
      RECT 1.1800 0.2565 1.2060 1.3500 ;
      RECT 1.0720 0.2565 1.0980 1.3500 ;
      RECT 0.9640 0.2565 0.9900 1.3500 ;
      RECT 0.8560 0.2565 0.8820 1.3500 ;
      RECT 0.7480 0.2565 0.7740 1.3500 ;
      RECT 0.6400 0.2565 0.6660 1.3500 ;
      RECT 0.5320 0.2565 0.5580 1.3500 ;
      RECT 0.4240 0.2565 0.4500 1.3500 ;
      RECT 0.3160 0.2565 0.3420 1.3500 ;
      RECT 0.2080 0.2565 0.2340 1.3500 ;
      RECT 0.0050 0.2565 0.0900 1.3500 ;
      RECT 15.5530 1.3365 15.6810 2.4300 ;
      RECT 15.5390 2.0020 15.6810 2.3245 ;
      RECT 15.3190 1.7290 15.4530 2.4300 ;
      RECT 15.2960 2.0640 15.4530 2.3220 ;
      RECT 15.3190 1.3365 15.4170 2.4300 ;
      RECT 15.3190 1.4575 15.4310 1.6970 ;
      RECT 15.3190 1.3365 15.4530 1.4255 ;
      RECT 15.0940 1.7870 15.2280 2.4300 ;
      RECT 15.0940 1.3365 15.1920 2.4300 ;
      RECT 14.6770 1.3365 14.7600 2.4300 ;
      RECT 14.6770 1.4250 14.7740 2.3605 ;
      RECT 30.2680 1.3365 30.3530 2.4300 ;
      RECT 30.1240 1.3365 30.1500 2.4300 ;
      RECT 30.0160 1.3365 30.0420 2.4300 ;
      RECT 29.9080 1.3365 29.9340 2.4300 ;
      RECT 29.8000 1.3365 29.8260 2.4300 ;
      RECT 29.6920 1.3365 29.7180 2.4300 ;
      RECT 29.5840 1.3365 29.6100 2.4300 ;
      RECT 29.4760 1.3365 29.5020 2.4300 ;
      RECT 29.3680 1.3365 29.3940 2.4300 ;
      RECT 29.2600 1.3365 29.2860 2.4300 ;
      RECT 29.1520 1.3365 29.1780 2.4300 ;
      RECT 29.0440 1.3365 29.0700 2.4300 ;
      RECT 28.9360 1.3365 28.9620 2.4300 ;
      RECT 28.8280 1.3365 28.8540 2.4300 ;
      RECT 28.7200 1.3365 28.7460 2.4300 ;
      RECT 28.6120 1.3365 28.6380 2.4300 ;
      RECT 28.5040 1.3365 28.5300 2.4300 ;
      RECT 28.3960 1.3365 28.4220 2.4300 ;
      RECT 28.2880 1.3365 28.3140 2.4300 ;
      RECT 28.1800 1.3365 28.2060 2.4300 ;
      RECT 28.0720 1.3365 28.0980 2.4300 ;
      RECT 27.9640 1.3365 27.9900 2.4300 ;
      RECT 27.8560 1.3365 27.8820 2.4300 ;
      RECT 27.7480 1.3365 27.7740 2.4300 ;
      RECT 27.6400 1.3365 27.6660 2.4300 ;
      RECT 27.5320 1.3365 27.5580 2.4300 ;
      RECT 27.4240 1.3365 27.4500 2.4300 ;
      RECT 27.3160 1.3365 27.3420 2.4300 ;
      RECT 27.2080 1.3365 27.2340 2.4300 ;
      RECT 27.1000 1.3365 27.1260 2.4300 ;
      RECT 26.9920 1.3365 27.0180 2.4300 ;
      RECT 26.8840 1.3365 26.9100 2.4300 ;
      RECT 26.7760 1.3365 26.8020 2.4300 ;
      RECT 26.6680 1.3365 26.6940 2.4300 ;
      RECT 26.5600 1.3365 26.5860 2.4300 ;
      RECT 26.4520 1.3365 26.4780 2.4300 ;
      RECT 26.3440 1.3365 26.3700 2.4300 ;
      RECT 26.2360 1.3365 26.2620 2.4300 ;
      RECT 26.1280 1.3365 26.1540 2.4300 ;
      RECT 26.0200 1.3365 26.0460 2.4300 ;
      RECT 25.9120 1.3365 25.9380 2.4300 ;
      RECT 25.8040 1.3365 25.8300 2.4300 ;
      RECT 25.6960 1.3365 25.7220 2.4300 ;
      RECT 25.5880 1.3365 25.6140 2.4300 ;
      RECT 25.4800 1.3365 25.5060 2.4300 ;
      RECT 25.3720 1.3365 25.3980 2.4300 ;
      RECT 25.2640 1.3365 25.2900 2.4300 ;
      RECT 25.1560 1.3365 25.1820 2.4300 ;
      RECT 25.0480 1.3365 25.0740 2.4300 ;
      RECT 24.9400 1.3365 24.9660 2.4300 ;
      RECT 24.8320 1.3365 24.8580 2.4300 ;
      RECT 24.7240 1.3365 24.7500 2.4300 ;
      RECT 24.6160 1.3365 24.6420 2.4300 ;
      RECT 24.5080 1.3365 24.5340 2.4300 ;
      RECT 24.4000 1.3365 24.4260 2.4300 ;
      RECT 24.2920 1.3365 24.3180 2.4300 ;
      RECT 24.1840 1.3365 24.2100 2.4300 ;
      RECT 24.0760 1.3365 24.1020 2.4300 ;
      RECT 23.9680 1.3365 23.9940 2.4300 ;
      RECT 23.8600 1.3365 23.8860 2.4300 ;
      RECT 23.7520 1.3365 23.7780 2.4300 ;
      RECT 23.6440 1.3365 23.6700 2.4300 ;
      RECT 23.5360 1.3365 23.5620 2.4300 ;
      RECT 23.4280 1.3365 23.4540 2.4300 ;
      RECT 23.3200 1.3365 23.3460 2.4300 ;
      RECT 23.2120 1.3365 23.2380 2.4300 ;
      RECT 23.1040 1.3365 23.1300 2.4300 ;
      RECT 22.9960 1.3365 23.0220 2.4300 ;
      RECT 22.8880 1.3365 22.9140 2.4300 ;
      RECT 22.7800 1.3365 22.8060 2.4300 ;
      RECT 22.6720 1.3365 22.6980 2.4300 ;
      RECT 22.5640 1.3365 22.5900 2.4300 ;
      RECT 22.4560 1.3365 22.4820 2.4300 ;
      RECT 22.3480 1.3365 22.3740 2.4300 ;
      RECT 22.2400 1.3365 22.2660 2.4300 ;
      RECT 22.1320 1.3365 22.1580 2.4300 ;
      RECT 22.0240 1.3365 22.0500 2.4300 ;
      RECT 21.9160 1.3365 21.9420 2.4300 ;
      RECT 21.8080 1.3365 21.8340 2.4300 ;
      RECT 21.7000 1.3365 21.7260 2.4300 ;
      RECT 21.5920 1.3365 21.6180 2.4300 ;
      RECT 21.4840 1.3365 21.5100 2.4300 ;
      RECT 21.3760 1.3365 21.4020 2.4300 ;
      RECT 21.2680 1.3365 21.2940 2.4300 ;
      RECT 21.1600 1.3365 21.1860 2.4300 ;
      RECT 21.0520 1.3365 21.0780 2.4300 ;
      RECT 20.9440 1.3365 20.9700 2.4300 ;
      RECT 20.8360 1.3365 20.8620 2.4300 ;
      RECT 20.7280 1.3365 20.7540 2.4300 ;
      RECT 20.6200 1.3365 20.6460 2.4300 ;
      RECT 20.5120 1.3365 20.5380 2.4300 ;
      RECT 20.4040 1.3365 20.4300 2.4300 ;
      RECT 20.2960 1.3365 20.3220 2.4300 ;
      RECT 20.1880 1.3365 20.2140 2.4300 ;
      RECT 20.0800 1.3365 20.1060 2.4300 ;
      RECT 19.9720 1.3365 19.9980 2.4300 ;
      RECT 19.8640 1.3365 19.8900 2.4300 ;
      RECT 19.7560 1.3365 19.7820 2.4300 ;
      RECT 19.6480 1.3365 19.6740 2.4300 ;
      RECT 19.5400 1.3365 19.5660 2.4300 ;
      RECT 19.4320 1.3365 19.4580 2.4300 ;
      RECT 19.3240 1.3365 19.3500 2.4300 ;
      RECT 19.2160 1.3365 19.2420 2.4300 ;
      RECT 19.1080 1.3365 19.1340 2.4300 ;
      RECT 19.0000 1.3365 19.0260 2.4300 ;
      RECT 18.8920 1.3365 18.9180 2.4300 ;
      RECT 18.7840 1.3365 18.8100 2.4300 ;
      RECT 18.6760 1.3365 18.7020 2.4300 ;
      RECT 18.5680 1.3365 18.5940 2.4300 ;
      RECT 18.4600 1.3365 18.4860 2.4300 ;
      RECT 18.3520 1.3365 18.3780 2.4300 ;
      RECT 18.2440 1.3365 18.2700 2.4300 ;
      RECT 18.1360 1.3365 18.1620 2.4300 ;
      RECT 18.0280 1.3365 18.0540 2.4300 ;
      RECT 17.9200 1.3365 17.9460 2.4300 ;
      RECT 17.8120 1.3365 17.8380 2.4300 ;
      RECT 17.7040 1.3365 17.7300 2.4300 ;
      RECT 17.5960 1.3365 17.6220 2.4300 ;
      RECT 17.4880 1.3365 17.5140 2.4300 ;
      RECT 17.3800 1.3365 17.4060 2.4300 ;
      RECT 17.2720 1.3365 17.2980 2.4300 ;
      RECT 17.1640 1.3365 17.1900 2.4300 ;
      RECT 17.0560 1.3365 17.0820 2.4300 ;
      RECT 16.9480 1.3365 16.9740 2.4300 ;
      RECT 16.8400 1.3365 16.8660 2.4300 ;
      RECT 16.7320 1.3365 16.7580 2.4300 ;
      RECT 16.6240 1.3365 16.6500 2.4300 ;
      RECT 16.5160 1.3365 16.5420 2.4300 ;
      RECT 16.4080 1.3365 16.4340 2.4300 ;
      RECT 16.3000 1.3365 16.3260 2.4300 ;
      RECT 16.0870 1.3365 16.1640 2.4300 ;
      RECT 14.1940 1.3365 14.2710 2.4300 ;
      RECT 14.0320 1.3365 14.0580 2.4300 ;
      RECT 13.9240 1.3365 13.9500 2.4300 ;
      RECT 13.8160 1.3365 13.8420 2.4300 ;
      RECT 13.7080 1.3365 13.7340 2.4300 ;
      RECT 13.6000 1.3365 13.6260 2.4300 ;
      RECT 13.4920 1.3365 13.5180 2.4300 ;
      RECT 13.3840 1.3365 13.4100 2.4300 ;
      RECT 13.2760 1.3365 13.3020 2.4300 ;
      RECT 13.1680 1.3365 13.1940 2.4300 ;
      RECT 13.0600 1.3365 13.0860 2.4300 ;
      RECT 12.9520 1.3365 12.9780 2.4300 ;
      RECT 12.8440 1.3365 12.8700 2.4300 ;
      RECT 12.7360 1.3365 12.7620 2.4300 ;
      RECT 12.6280 1.3365 12.6540 2.4300 ;
      RECT 12.5200 1.3365 12.5460 2.4300 ;
      RECT 12.4120 1.3365 12.4380 2.4300 ;
      RECT 12.3040 1.3365 12.3300 2.4300 ;
      RECT 12.1960 1.3365 12.2220 2.4300 ;
      RECT 12.0880 1.3365 12.1140 2.4300 ;
      RECT 11.9800 1.3365 12.0060 2.4300 ;
      RECT 11.8720 1.3365 11.8980 2.4300 ;
      RECT 11.7640 1.3365 11.7900 2.4300 ;
      RECT 11.6560 1.3365 11.6820 2.4300 ;
      RECT 11.5480 1.3365 11.5740 2.4300 ;
      RECT 11.4400 1.3365 11.4660 2.4300 ;
      RECT 11.3320 1.3365 11.3580 2.4300 ;
      RECT 11.2240 1.3365 11.2500 2.4300 ;
      RECT 11.1160 1.3365 11.1420 2.4300 ;
      RECT 11.0080 1.3365 11.0340 2.4300 ;
      RECT 10.9000 1.3365 10.9260 2.4300 ;
      RECT 10.7920 1.3365 10.8180 2.4300 ;
      RECT 10.6840 1.3365 10.7100 2.4300 ;
      RECT 10.5760 1.3365 10.6020 2.4300 ;
      RECT 10.4680 1.3365 10.4940 2.4300 ;
      RECT 10.3600 1.3365 10.3860 2.4300 ;
      RECT 10.2520 1.3365 10.2780 2.4300 ;
      RECT 10.1440 1.3365 10.1700 2.4300 ;
      RECT 10.0360 1.3365 10.0620 2.4300 ;
      RECT 9.9280 1.3365 9.9540 2.4300 ;
      RECT 9.8200 1.3365 9.8460 2.4300 ;
      RECT 9.7120 1.3365 9.7380 2.4300 ;
      RECT 9.6040 1.3365 9.6300 2.4300 ;
      RECT 9.4960 1.3365 9.5220 2.4300 ;
      RECT 9.3880 1.3365 9.4140 2.4300 ;
      RECT 9.2800 1.3365 9.3060 2.4300 ;
      RECT 9.1720 1.3365 9.1980 2.4300 ;
      RECT 9.0640 1.3365 9.0900 2.4300 ;
      RECT 8.9560 1.3365 8.9820 2.4300 ;
      RECT 8.8480 1.3365 8.8740 2.4300 ;
      RECT 8.7400 1.3365 8.7660 2.4300 ;
      RECT 8.6320 1.3365 8.6580 2.4300 ;
      RECT 8.5240 1.3365 8.5500 2.4300 ;
      RECT 8.4160 1.3365 8.4420 2.4300 ;
      RECT 8.3080 1.3365 8.3340 2.4300 ;
      RECT 8.2000 1.3365 8.2260 2.4300 ;
      RECT 8.0920 1.3365 8.1180 2.4300 ;
      RECT 7.9840 1.3365 8.0100 2.4300 ;
      RECT 7.8760 1.3365 7.9020 2.4300 ;
      RECT 7.7680 1.3365 7.7940 2.4300 ;
      RECT 7.6600 1.3365 7.6860 2.4300 ;
      RECT 7.5520 1.3365 7.5780 2.4300 ;
      RECT 7.4440 1.3365 7.4700 2.4300 ;
      RECT 7.3360 1.3365 7.3620 2.4300 ;
      RECT 7.2280 1.3365 7.2540 2.4300 ;
      RECT 7.1200 1.3365 7.1460 2.4300 ;
      RECT 7.0120 1.3365 7.0380 2.4300 ;
      RECT 6.9040 1.3365 6.9300 2.4300 ;
      RECT 6.7960 1.3365 6.8220 2.4300 ;
      RECT 6.6880 1.3365 6.7140 2.4300 ;
      RECT 6.5800 1.3365 6.6060 2.4300 ;
      RECT 6.4720 1.3365 6.4980 2.4300 ;
      RECT 6.3640 1.3365 6.3900 2.4300 ;
      RECT 6.2560 1.3365 6.2820 2.4300 ;
      RECT 6.1480 1.3365 6.1740 2.4300 ;
      RECT 6.0400 1.3365 6.0660 2.4300 ;
      RECT 5.9320 1.3365 5.9580 2.4300 ;
      RECT 5.8240 1.3365 5.8500 2.4300 ;
      RECT 5.7160 1.3365 5.7420 2.4300 ;
      RECT 5.6080 1.3365 5.6340 2.4300 ;
      RECT 5.5000 1.3365 5.5260 2.4300 ;
      RECT 5.3920 1.3365 5.4180 2.4300 ;
      RECT 5.2840 1.3365 5.3100 2.4300 ;
      RECT 5.1760 1.3365 5.2020 2.4300 ;
      RECT 5.0680 1.3365 5.0940 2.4300 ;
      RECT 4.9600 1.3365 4.9860 2.4300 ;
      RECT 4.8520 1.3365 4.8780 2.4300 ;
      RECT 4.7440 1.3365 4.7700 2.4300 ;
      RECT 4.6360 1.3365 4.6620 2.4300 ;
      RECT 4.5280 1.3365 4.5540 2.4300 ;
      RECT 4.4200 1.3365 4.4460 2.4300 ;
      RECT 4.3120 1.3365 4.3380 2.4300 ;
      RECT 4.2040 1.3365 4.2300 2.4300 ;
      RECT 4.0960 1.3365 4.1220 2.4300 ;
      RECT 3.9880 1.3365 4.0140 2.4300 ;
      RECT 3.8800 1.3365 3.9060 2.4300 ;
      RECT 3.7720 1.3365 3.7980 2.4300 ;
      RECT 3.6640 1.3365 3.6900 2.4300 ;
      RECT 3.5560 1.3365 3.5820 2.4300 ;
      RECT 3.4480 1.3365 3.4740 2.4300 ;
      RECT 3.3400 1.3365 3.3660 2.4300 ;
      RECT 3.2320 1.3365 3.2580 2.4300 ;
      RECT 3.1240 1.3365 3.1500 2.4300 ;
      RECT 3.0160 1.3365 3.0420 2.4300 ;
      RECT 2.9080 1.3365 2.9340 2.4300 ;
      RECT 2.8000 1.3365 2.8260 2.4300 ;
      RECT 2.6920 1.3365 2.7180 2.4300 ;
      RECT 2.5840 1.3365 2.6100 2.4300 ;
      RECT 2.4760 1.3365 2.5020 2.4300 ;
      RECT 2.3680 1.3365 2.3940 2.4300 ;
      RECT 2.2600 1.3365 2.2860 2.4300 ;
      RECT 2.1520 1.3365 2.1780 2.4300 ;
      RECT 2.0440 1.3365 2.0700 2.4300 ;
      RECT 1.9360 1.3365 1.9620 2.4300 ;
      RECT 1.8280 1.3365 1.8540 2.4300 ;
      RECT 1.7200 1.3365 1.7460 2.4300 ;
      RECT 1.6120 1.3365 1.6380 2.4300 ;
      RECT 1.5040 1.3365 1.5300 2.4300 ;
      RECT 1.3960 1.3365 1.4220 2.4300 ;
      RECT 1.2880 1.3365 1.3140 2.4300 ;
      RECT 1.1800 1.3365 1.2060 2.4300 ;
      RECT 1.0720 1.3365 1.0980 2.4300 ;
      RECT 0.9640 1.3365 0.9900 2.4300 ;
      RECT 0.8560 1.3365 0.8820 2.4300 ;
      RECT 0.7480 1.3365 0.7740 2.4300 ;
      RECT 0.6400 1.3365 0.6660 2.4300 ;
      RECT 0.5320 1.3365 0.5580 2.4300 ;
      RECT 0.4240 1.3365 0.4500 2.4300 ;
      RECT 0.3160 1.3365 0.3420 2.4300 ;
      RECT 0.2080 1.3365 0.2340 2.4300 ;
      RECT 0.0050 1.3365 0.0900 2.4300 ;
      RECT 15.5530 2.4165 15.6810 3.5100 ;
      RECT 15.5390 3.0820 15.6810 3.4045 ;
      RECT 15.3190 2.8090 15.4530 3.5100 ;
      RECT 15.2960 3.1440 15.4530 3.4020 ;
      RECT 15.3190 2.4165 15.4170 3.5100 ;
      RECT 15.3190 2.5375 15.4310 2.7770 ;
      RECT 15.3190 2.4165 15.4530 2.5055 ;
      RECT 15.0940 2.8670 15.2280 3.5100 ;
      RECT 15.0940 2.4165 15.1920 3.5100 ;
      RECT 14.6770 2.4165 14.7600 3.5100 ;
      RECT 14.6770 2.5050 14.7740 3.4405 ;
      RECT 30.2680 2.4165 30.3530 3.5100 ;
      RECT 30.1240 2.4165 30.1500 3.5100 ;
      RECT 30.0160 2.4165 30.0420 3.5100 ;
      RECT 29.9080 2.4165 29.9340 3.5100 ;
      RECT 29.8000 2.4165 29.8260 3.5100 ;
      RECT 29.6920 2.4165 29.7180 3.5100 ;
      RECT 29.5840 2.4165 29.6100 3.5100 ;
      RECT 29.4760 2.4165 29.5020 3.5100 ;
      RECT 29.3680 2.4165 29.3940 3.5100 ;
      RECT 29.2600 2.4165 29.2860 3.5100 ;
      RECT 29.1520 2.4165 29.1780 3.5100 ;
      RECT 29.0440 2.4165 29.0700 3.5100 ;
      RECT 28.9360 2.4165 28.9620 3.5100 ;
      RECT 28.8280 2.4165 28.8540 3.5100 ;
      RECT 28.7200 2.4165 28.7460 3.5100 ;
      RECT 28.6120 2.4165 28.6380 3.5100 ;
      RECT 28.5040 2.4165 28.5300 3.5100 ;
      RECT 28.3960 2.4165 28.4220 3.5100 ;
      RECT 28.2880 2.4165 28.3140 3.5100 ;
      RECT 28.1800 2.4165 28.2060 3.5100 ;
      RECT 28.0720 2.4165 28.0980 3.5100 ;
      RECT 27.9640 2.4165 27.9900 3.5100 ;
      RECT 27.8560 2.4165 27.8820 3.5100 ;
      RECT 27.7480 2.4165 27.7740 3.5100 ;
      RECT 27.6400 2.4165 27.6660 3.5100 ;
      RECT 27.5320 2.4165 27.5580 3.5100 ;
      RECT 27.4240 2.4165 27.4500 3.5100 ;
      RECT 27.3160 2.4165 27.3420 3.5100 ;
      RECT 27.2080 2.4165 27.2340 3.5100 ;
      RECT 27.1000 2.4165 27.1260 3.5100 ;
      RECT 26.9920 2.4165 27.0180 3.5100 ;
      RECT 26.8840 2.4165 26.9100 3.5100 ;
      RECT 26.7760 2.4165 26.8020 3.5100 ;
      RECT 26.6680 2.4165 26.6940 3.5100 ;
      RECT 26.5600 2.4165 26.5860 3.5100 ;
      RECT 26.4520 2.4165 26.4780 3.5100 ;
      RECT 26.3440 2.4165 26.3700 3.5100 ;
      RECT 26.2360 2.4165 26.2620 3.5100 ;
      RECT 26.1280 2.4165 26.1540 3.5100 ;
      RECT 26.0200 2.4165 26.0460 3.5100 ;
      RECT 25.9120 2.4165 25.9380 3.5100 ;
      RECT 25.8040 2.4165 25.8300 3.5100 ;
      RECT 25.6960 2.4165 25.7220 3.5100 ;
      RECT 25.5880 2.4165 25.6140 3.5100 ;
      RECT 25.4800 2.4165 25.5060 3.5100 ;
      RECT 25.3720 2.4165 25.3980 3.5100 ;
      RECT 25.2640 2.4165 25.2900 3.5100 ;
      RECT 25.1560 2.4165 25.1820 3.5100 ;
      RECT 25.0480 2.4165 25.0740 3.5100 ;
      RECT 24.9400 2.4165 24.9660 3.5100 ;
      RECT 24.8320 2.4165 24.8580 3.5100 ;
      RECT 24.7240 2.4165 24.7500 3.5100 ;
      RECT 24.6160 2.4165 24.6420 3.5100 ;
      RECT 24.5080 2.4165 24.5340 3.5100 ;
      RECT 24.4000 2.4165 24.4260 3.5100 ;
      RECT 24.2920 2.4165 24.3180 3.5100 ;
      RECT 24.1840 2.4165 24.2100 3.5100 ;
      RECT 24.0760 2.4165 24.1020 3.5100 ;
      RECT 23.9680 2.4165 23.9940 3.5100 ;
      RECT 23.8600 2.4165 23.8860 3.5100 ;
      RECT 23.7520 2.4165 23.7780 3.5100 ;
      RECT 23.6440 2.4165 23.6700 3.5100 ;
      RECT 23.5360 2.4165 23.5620 3.5100 ;
      RECT 23.4280 2.4165 23.4540 3.5100 ;
      RECT 23.3200 2.4165 23.3460 3.5100 ;
      RECT 23.2120 2.4165 23.2380 3.5100 ;
      RECT 23.1040 2.4165 23.1300 3.5100 ;
      RECT 22.9960 2.4165 23.0220 3.5100 ;
      RECT 22.8880 2.4165 22.9140 3.5100 ;
      RECT 22.7800 2.4165 22.8060 3.5100 ;
      RECT 22.6720 2.4165 22.6980 3.5100 ;
      RECT 22.5640 2.4165 22.5900 3.5100 ;
      RECT 22.4560 2.4165 22.4820 3.5100 ;
      RECT 22.3480 2.4165 22.3740 3.5100 ;
      RECT 22.2400 2.4165 22.2660 3.5100 ;
      RECT 22.1320 2.4165 22.1580 3.5100 ;
      RECT 22.0240 2.4165 22.0500 3.5100 ;
      RECT 21.9160 2.4165 21.9420 3.5100 ;
      RECT 21.8080 2.4165 21.8340 3.5100 ;
      RECT 21.7000 2.4165 21.7260 3.5100 ;
      RECT 21.5920 2.4165 21.6180 3.5100 ;
      RECT 21.4840 2.4165 21.5100 3.5100 ;
      RECT 21.3760 2.4165 21.4020 3.5100 ;
      RECT 21.2680 2.4165 21.2940 3.5100 ;
      RECT 21.1600 2.4165 21.1860 3.5100 ;
      RECT 21.0520 2.4165 21.0780 3.5100 ;
      RECT 20.9440 2.4165 20.9700 3.5100 ;
      RECT 20.8360 2.4165 20.8620 3.5100 ;
      RECT 20.7280 2.4165 20.7540 3.5100 ;
      RECT 20.6200 2.4165 20.6460 3.5100 ;
      RECT 20.5120 2.4165 20.5380 3.5100 ;
      RECT 20.4040 2.4165 20.4300 3.5100 ;
      RECT 20.2960 2.4165 20.3220 3.5100 ;
      RECT 20.1880 2.4165 20.2140 3.5100 ;
      RECT 20.0800 2.4165 20.1060 3.5100 ;
      RECT 19.9720 2.4165 19.9980 3.5100 ;
      RECT 19.8640 2.4165 19.8900 3.5100 ;
      RECT 19.7560 2.4165 19.7820 3.5100 ;
      RECT 19.6480 2.4165 19.6740 3.5100 ;
      RECT 19.5400 2.4165 19.5660 3.5100 ;
      RECT 19.4320 2.4165 19.4580 3.5100 ;
      RECT 19.3240 2.4165 19.3500 3.5100 ;
      RECT 19.2160 2.4165 19.2420 3.5100 ;
      RECT 19.1080 2.4165 19.1340 3.5100 ;
      RECT 19.0000 2.4165 19.0260 3.5100 ;
      RECT 18.8920 2.4165 18.9180 3.5100 ;
      RECT 18.7840 2.4165 18.8100 3.5100 ;
      RECT 18.6760 2.4165 18.7020 3.5100 ;
      RECT 18.5680 2.4165 18.5940 3.5100 ;
      RECT 18.4600 2.4165 18.4860 3.5100 ;
      RECT 18.3520 2.4165 18.3780 3.5100 ;
      RECT 18.2440 2.4165 18.2700 3.5100 ;
      RECT 18.1360 2.4165 18.1620 3.5100 ;
      RECT 18.0280 2.4165 18.0540 3.5100 ;
      RECT 17.9200 2.4165 17.9460 3.5100 ;
      RECT 17.8120 2.4165 17.8380 3.5100 ;
      RECT 17.7040 2.4165 17.7300 3.5100 ;
      RECT 17.5960 2.4165 17.6220 3.5100 ;
      RECT 17.4880 2.4165 17.5140 3.5100 ;
      RECT 17.3800 2.4165 17.4060 3.5100 ;
      RECT 17.2720 2.4165 17.2980 3.5100 ;
      RECT 17.1640 2.4165 17.1900 3.5100 ;
      RECT 17.0560 2.4165 17.0820 3.5100 ;
      RECT 16.9480 2.4165 16.9740 3.5100 ;
      RECT 16.8400 2.4165 16.8660 3.5100 ;
      RECT 16.7320 2.4165 16.7580 3.5100 ;
      RECT 16.6240 2.4165 16.6500 3.5100 ;
      RECT 16.5160 2.4165 16.5420 3.5100 ;
      RECT 16.4080 2.4165 16.4340 3.5100 ;
      RECT 16.3000 2.4165 16.3260 3.5100 ;
      RECT 16.0870 2.4165 16.1640 3.5100 ;
      RECT 14.1940 2.4165 14.2710 3.5100 ;
      RECT 14.0320 2.4165 14.0580 3.5100 ;
      RECT 13.9240 2.4165 13.9500 3.5100 ;
      RECT 13.8160 2.4165 13.8420 3.5100 ;
      RECT 13.7080 2.4165 13.7340 3.5100 ;
      RECT 13.6000 2.4165 13.6260 3.5100 ;
      RECT 13.4920 2.4165 13.5180 3.5100 ;
      RECT 13.3840 2.4165 13.4100 3.5100 ;
      RECT 13.2760 2.4165 13.3020 3.5100 ;
      RECT 13.1680 2.4165 13.1940 3.5100 ;
      RECT 13.0600 2.4165 13.0860 3.5100 ;
      RECT 12.9520 2.4165 12.9780 3.5100 ;
      RECT 12.8440 2.4165 12.8700 3.5100 ;
      RECT 12.7360 2.4165 12.7620 3.5100 ;
      RECT 12.6280 2.4165 12.6540 3.5100 ;
      RECT 12.5200 2.4165 12.5460 3.5100 ;
      RECT 12.4120 2.4165 12.4380 3.5100 ;
      RECT 12.3040 2.4165 12.3300 3.5100 ;
      RECT 12.1960 2.4165 12.2220 3.5100 ;
      RECT 12.0880 2.4165 12.1140 3.5100 ;
      RECT 11.9800 2.4165 12.0060 3.5100 ;
      RECT 11.8720 2.4165 11.8980 3.5100 ;
      RECT 11.7640 2.4165 11.7900 3.5100 ;
      RECT 11.6560 2.4165 11.6820 3.5100 ;
      RECT 11.5480 2.4165 11.5740 3.5100 ;
      RECT 11.4400 2.4165 11.4660 3.5100 ;
      RECT 11.3320 2.4165 11.3580 3.5100 ;
      RECT 11.2240 2.4165 11.2500 3.5100 ;
      RECT 11.1160 2.4165 11.1420 3.5100 ;
      RECT 11.0080 2.4165 11.0340 3.5100 ;
      RECT 10.9000 2.4165 10.9260 3.5100 ;
      RECT 10.7920 2.4165 10.8180 3.5100 ;
      RECT 10.6840 2.4165 10.7100 3.5100 ;
      RECT 10.5760 2.4165 10.6020 3.5100 ;
      RECT 10.4680 2.4165 10.4940 3.5100 ;
      RECT 10.3600 2.4165 10.3860 3.5100 ;
      RECT 10.2520 2.4165 10.2780 3.5100 ;
      RECT 10.1440 2.4165 10.1700 3.5100 ;
      RECT 10.0360 2.4165 10.0620 3.5100 ;
      RECT 9.9280 2.4165 9.9540 3.5100 ;
      RECT 9.8200 2.4165 9.8460 3.5100 ;
      RECT 9.7120 2.4165 9.7380 3.5100 ;
      RECT 9.6040 2.4165 9.6300 3.5100 ;
      RECT 9.4960 2.4165 9.5220 3.5100 ;
      RECT 9.3880 2.4165 9.4140 3.5100 ;
      RECT 9.2800 2.4165 9.3060 3.5100 ;
      RECT 9.1720 2.4165 9.1980 3.5100 ;
      RECT 9.0640 2.4165 9.0900 3.5100 ;
      RECT 8.9560 2.4165 8.9820 3.5100 ;
      RECT 8.8480 2.4165 8.8740 3.5100 ;
      RECT 8.7400 2.4165 8.7660 3.5100 ;
      RECT 8.6320 2.4165 8.6580 3.5100 ;
      RECT 8.5240 2.4165 8.5500 3.5100 ;
      RECT 8.4160 2.4165 8.4420 3.5100 ;
      RECT 8.3080 2.4165 8.3340 3.5100 ;
      RECT 8.2000 2.4165 8.2260 3.5100 ;
      RECT 8.0920 2.4165 8.1180 3.5100 ;
      RECT 7.9840 2.4165 8.0100 3.5100 ;
      RECT 7.8760 2.4165 7.9020 3.5100 ;
      RECT 7.7680 2.4165 7.7940 3.5100 ;
      RECT 7.6600 2.4165 7.6860 3.5100 ;
      RECT 7.5520 2.4165 7.5780 3.5100 ;
      RECT 7.4440 2.4165 7.4700 3.5100 ;
      RECT 7.3360 2.4165 7.3620 3.5100 ;
      RECT 7.2280 2.4165 7.2540 3.5100 ;
      RECT 7.1200 2.4165 7.1460 3.5100 ;
      RECT 7.0120 2.4165 7.0380 3.5100 ;
      RECT 6.9040 2.4165 6.9300 3.5100 ;
      RECT 6.7960 2.4165 6.8220 3.5100 ;
      RECT 6.6880 2.4165 6.7140 3.5100 ;
      RECT 6.5800 2.4165 6.6060 3.5100 ;
      RECT 6.4720 2.4165 6.4980 3.5100 ;
      RECT 6.3640 2.4165 6.3900 3.5100 ;
      RECT 6.2560 2.4165 6.2820 3.5100 ;
      RECT 6.1480 2.4165 6.1740 3.5100 ;
      RECT 6.0400 2.4165 6.0660 3.5100 ;
      RECT 5.9320 2.4165 5.9580 3.5100 ;
      RECT 5.8240 2.4165 5.8500 3.5100 ;
      RECT 5.7160 2.4165 5.7420 3.5100 ;
      RECT 5.6080 2.4165 5.6340 3.5100 ;
      RECT 5.5000 2.4165 5.5260 3.5100 ;
      RECT 5.3920 2.4165 5.4180 3.5100 ;
      RECT 5.2840 2.4165 5.3100 3.5100 ;
      RECT 5.1760 2.4165 5.2020 3.5100 ;
      RECT 5.0680 2.4165 5.0940 3.5100 ;
      RECT 4.9600 2.4165 4.9860 3.5100 ;
      RECT 4.8520 2.4165 4.8780 3.5100 ;
      RECT 4.7440 2.4165 4.7700 3.5100 ;
      RECT 4.6360 2.4165 4.6620 3.5100 ;
      RECT 4.5280 2.4165 4.5540 3.5100 ;
      RECT 4.4200 2.4165 4.4460 3.5100 ;
      RECT 4.3120 2.4165 4.3380 3.5100 ;
      RECT 4.2040 2.4165 4.2300 3.5100 ;
      RECT 4.0960 2.4165 4.1220 3.5100 ;
      RECT 3.9880 2.4165 4.0140 3.5100 ;
      RECT 3.8800 2.4165 3.9060 3.5100 ;
      RECT 3.7720 2.4165 3.7980 3.5100 ;
      RECT 3.6640 2.4165 3.6900 3.5100 ;
      RECT 3.5560 2.4165 3.5820 3.5100 ;
      RECT 3.4480 2.4165 3.4740 3.5100 ;
      RECT 3.3400 2.4165 3.3660 3.5100 ;
      RECT 3.2320 2.4165 3.2580 3.5100 ;
      RECT 3.1240 2.4165 3.1500 3.5100 ;
      RECT 3.0160 2.4165 3.0420 3.5100 ;
      RECT 2.9080 2.4165 2.9340 3.5100 ;
      RECT 2.8000 2.4165 2.8260 3.5100 ;
      RECT 2.6920 2.4165 2.7180 3.5100 ;
      RECT 2.5840 2.4165 2.6100 3.5100 ;
      RECT 2.4760 2.4165 2.5020 3.5100 ;
      RECT 2.3680 2.4165 2.3940 3.5100 ;
      RECT 2.2600 2.4165 2.2860 3.5100 ;
      RECT 2.1520 2.4165 2.1780 3.5100 ;
      RECT 2.0440 2.4165 2.0700 3.5100 ;
      RECT 1.9360 2.4165 1.9620 3.5100 ;
      RECT 1.8280 2.4165 1.8540 3.5100 ;
      RECT 1.7200 2.4165 1.7460 3.5100 ;
      RECT 1.6120 2.4165 1.6380 3.5100 ;
      RECT 1.5040 2.4165 1.5300 3.5100 ;
      RECT 1.3960 2.4165 1.4220 3.5100 ;
      RECT 1.2880 2.4165 1.3140 3.5100 ;
      RECT 1.1800 2.4165 1.2060 3.5100 ;
      RECT 1.0720 2.4165 1.0980 3.5100 ;
      RECT 0.9640 2.4165 0.9900 3.5100 ;
      RECT 0.8560 2.4165 0.8820 3.5100 ;
      RECT 0.7480 2.4165 0.7740 3.5100 ;
      RECT 0.6400 2.4165 0.6660 3.5100 ;
      RECT 0.5320 2.4165 0.5580 3.5100 ;
      RECT 0.4240 2.4165 0.4500 3.5100 ;
      RECT 0.3160 2.4165 0.3420 3.5100 ;
      RECT 0.2080 2.4165 0.2340 3.5100 ;
      RECT 0.0050 2.4165 0.0900 3.5100 ;
      RECT 15.5530 3.4965 15.6810 4.5900 ;
      RECT 15.5390 4.1620 15.6810 4.4845 ;
      RECT 15.3190 3.8890 15.4530 4.5900 ;
      RECT 15.2960 4.2240 15.4530 4.4820 ;
      RECT 15.3190 3.4965 15.4170 4.5900 ;
      RECT 15.3190 3.6175 15.4310 3.8570 ;
      RECT 15.3190 3.4965 15.4530 3.5855 ;
      RECT 15.0940 3.9470 15.2280 4.5900 ;
      RECT 15.0940 3.4965 15.1920 4.5900 ;
      RECT 14.6770 3.4965 14.7600 4.5900 ;
      RECT 14.6770 3.5850 14.7740 4.5205 ;
      RECT 30.2680 3.4965 30.3530 4.5900 ;
      RECT 30.1240 3.4965 30.1500 4.5900 ;
      RECT 30.0160 3.4965 30.0420 4.5900 ;
      RECT 29.9080 3.4965 29.9340 4.5900 ;
      RECT 29.8000 3.4965 29.8260 4.5900 ;
      RECT 29.6920 3.4965 29.7180 4.5900 ;
      RECT 29.5840 3.4965 29.6100 4.5900 ;
      RECT 29.4760 3.4965 29.5020 4.5900 ;
      RECT 29.3680 3.4965 29.3940 4.5900 ;
      RECT 29.2600 3.4965 29.2860 4.5900 ;
      RECT 29.1520 3.4965 29.1780 4.5900 ;
      RECT 29.0440 3.4965 29.0700 4.5900 ;
      RECT 28.9360 3.4965 28.9620 4.5900 ;
      RECT 28.8280 3.4965 28.8540 4.5900 ;
      RECT 28.7200 3.4965 28.7460 4.5900 ;
      RECT 28.6120 3.4965 28.6380 4.5900 ;
      RECT 28.5040 3.4965 28.5300 4.5900 ;
      RECT 28.3960 3.4965 28.4220 4.5900 ;
      RECT 28.2880 3.4965 28.3140 4.5900 ;
      RECT 28.1800 3.4965 28.2060 4.5900 ;
      RECT 28.0720 3.4965 28.0980 4.5900 ;
      RECT 27.9640 3.4965 27.9900 4.5900 ;
      RECT 27.8560 3.4965 27.8820 4.5900 ;
      RECT 27.7480 3.4965 27.7740 4.5900 ;
      RECT 27.6400 3.4965 27.6660 4.5900 ;
      RECT 27.5320 3.4965 27.5580 4.5900 ;
      RECT 27.4240 3.4965 27.4500 4.5900 ;
      RECT 27.3160 3.4965 27.3420 4.5900 ;
      RECT 27.2080 3.4965 27.2340 4.5900 ;
      RECT 27.1000 3.4965 27.1260 4.5900 ;
      RECT 26.9920 3.4965 27.0180 4.5900 ;
      RECT 26.8840 3.4965 26.9100 4.5900 ;
      RECT 26.7760 3.4965 26.8020 4.5900 ;
      RECT 26.6680 3.4965 26.6940 4.5900 ;
      RECT 26.5600 3.4965 26.5860 4.5900 ;
      RECT 26.4520 3.4965 26.4780 4.5900 ;
      RECT 26.3440 3.4965 26.3700 4.5900 ;
      RECT 26.2360 3.4965 26.2620 4.5900 ;
      RECT 26.1280 3.4965 26.1540 4.5900 ;
      RECT 26.0200 3.4965 26.0460 4.5900 ;
      RECT 25.9120 3.4965 25.9380 4.5900 ;
      RECT 25.8040 3.4965 25.8300 4.5900 ;
      RECT 25.6960 3.4965 25.7220 4.5900 ;
      RECT 25.5880 3.4965 25.6140 4.5900 ;
      RECT 25.4800 3.4965 25.5060 4.5900 ;
      RECT 25.3720 3.4965 25.3980 4.5900 ;
      RECT 25.2640 3.4965 25.2900 4.5900 ;
      RECT 25.1560 3.4965 25.1820 4.5900 ;
      RECT 25.0480 3.4965 25.0740 4.5900 ;
      RECT 24.9400 3.4965 24.9660 4.5900 ;
      RECT 24.8320 3.4965 24.8580 4.5900 ;
      RECT 24.7240 3.4965 24.7500 4.5900 ;
      RECT 24.6160 3.4965 24.6420 4.5900 ;
      RECT 24.5080 3.4965 24.5340 4.5900 ;
      RECT 24.4000 3.4965 24.4260 4.5900 ;
      RECT 24.2920 3.4965 24.3180 4.5900 ;
      RECT 24.1840 3.4965 24.2100 4.5900 ;
      RECT 24.0760 3.4965 24.1020 4.5900 ;
      RECT 23.9680 3.4965 23.9940 4.5900 ;
      RECT 23.8600 3.4965 23.8860 4.5900 ;
      RECT 23.7520 3.4965 23.7780 4.5900 ;
      RECT 23.6440 3.4965 23.6700 4.5900 ;
      RECT 23.5360 3.4965 23.5620 4.5900 ;
      RECT 23.4280 3.4965 23.4540 4.5900 ;
      RECT 23.3200 3.4965 23.3460 4.5900 ;
      RECT 23.2120 3.4965 23.2380 4.5900 ;
      RECT 23.1040 3.4965 23.1300 4.5900 ;
      RECT 22.9960 3.4965 23.0220 4.5900 ;
      RECT 22.8880 3.4965 22.9140 4.5900 ;
      RECT 22.7800 3.4965 22.8060 4.5900 ;
      RECT 22.6720 3.4965 22.6980 4.5900 ;
      RECT 22.5640 3.4965 22.5900 4.5900 ;
      RECT 22.4560 3.4965 22.4820 4.5900 ;
      RECT 22.3480 3.4965 22.3740 4.5900 ;
      RECT 22.2400 3.4965 22.2660 4.5900 ;
      RECT 22.1320 3.4965 22.1580 4.5900 ;
      RECT 22.0240 3.4965 22.0500 4.5900 ;
      RECT 21.9160 3.4965 21.9420 4.5900 ;
      RECT 21.8080 3.4965 21.8340 4.5900 ;
      RECT 21.7000 3.4965 21.7260 4.5900 ;
      RECT 21.5920 3.4965 21.6180 4.5900 ;
      RECT 21.4840 3.4965 21.5100 4.5900 ;
      RECT 21.3760 3.4965 21.4020 4.5900 ;
      RECT 21.2680 3.4965 21.2940 4.5900 ;
      RECT 21.1600 3.4965 21.1860 4.5900 ;
      RECT 21.0520 3.4965 21.0780 4.5900 ;
      RECT 20.9440 3.4965 20.9700 4.5900 ;
      RECT 20.8360 3.4965 20.8620 4.5900 ;
      RECT 20.7280 3.4965 20.7540 4.5900 ;
      RECT 20.6200 3.4965 20.6460 4.5900 ;
      RECT 20.5120 3.4965 20.5380 4.5900 ;
      RECT 20.4040 3.4965 20.4300 4.5900 ;
      RECT 20.2960 3.4965 20.3220 4.5900 ;
      RECT 20.1880 3.4965 20.2140 4.5900 ;
      RECT 20.0800 3.4965 20.1060 4.5900 ;
      RECT 19.9720 3.4965 19.9980 4.5900 ;
      RECT 19.8640 3.4965 19.8900 4.5900 ;
      RECT 19.7560 3.4965 19.7820 4.5900 ;
      RECT 19.6480 3.4965 19.6740 4.5900 ;
      RECT 19.5400 3.4965 19.5660 4.5900 ;
      RECT 19.4320 3.4965 19.4580 4.5900 ;
      RECT 19.3240 3.4965 19.3500 4.5900 ;
      RECT 19.2160 3.4965 19.2420 4.5900 ;
      RECT 19.1080 3.4965 19.1340 4.5900 ;
      RECT 19.0000 3.4965 19.0260 4.5900 ;
      RECT 18.8920 3.4965 18.9180 4.5900 ;
      RECT 18.7840 3.4965 18.8100 4.5900 ;
      RECT 18.6760 3.4965 18.7020 4.5900 ;
      RECT 18.5680 3.4965 18.5940 4.5900 ;
      RECT 18.4600 3.4965 18.4860 4.5900 ;
      RECT 18.3520 3.4965 18.3780 4.5900 ;
      RECT 18.2440 3.4965 18.2700 4.5900 ;
      RECT 18.1360 3.4965 18.1620 4.5900 ;
      RECT 18.0280 3.4965 18.0540 4.5900 ;
      RECT 17.9200 3.4965 17.9460 4.5900 ;
      RECT 17.8120 3.4965 17.8380 4.5900 ;
      RECT 17.7040 3.4965 17.7300 4.5900 ;
      RECT 17.5960 3.4965 17.6220 4.5900 ;
      RECT 17.4880 3.4965 17.5140 4.5900 ;
      RECT 17.3800 3.4965 17.4060 4.5900 ;
      RECT 17.2720 3.4965 17.2980 4.5900 ;
      RECT 17.1640 3.4965 17.1900 4.5900 ;
      RECT 17.0560 3.4965 17.0820 4.5900 ;
      RECT 16.9480 3.4965 16.9740 4.5900 ;
      RECT 16.8400 3.4965 16.8660 4.5900 ;
      RECT 16.7320 3.4965 16.7580 4.5900 ;
      RECT 16.6240 3.4965 16.6500 4.5900 ;
      RECT 16.5160 3.4965 16.5420 4.5900 ;
      RECT 16.4080 3.4965 16.4340 4.5900 ;
      RECT 16.3000 3.4965 16.3260 4.5900 ;
      RECT 16.0870 3.4965 16.1640 4.5900 ;
      RECT 14.1940 3.4965 14.2710 4.5900 ;
      RECT 14.0320 3.4965 14.0580 4.5900 ;
      RECT 13.9240 3.4965 13.9500 4.5900 ;
      RECT 13.8160 3.4965 13.8420 4.5900 ;
      RECT 13.7080 3.4965 13.7340 4.5900 ;
      RECT 13.6000 3.4965 13.6260 4.5900 ;
      RECT 13.4920 3.4965 13.5180 4.5900 ;
      RECT 13.3840 3.4965 13.4100 4.5900 ;
      RECT 13.2760 3.4965 13.3020 4.5900 ;
      RECT 13.1680 3.4965 13.1940 4.5900 ;
      RECT 13.0600 3.4965 13.0860 4.5900 ;
      RECT 12.9520 3.4965 12.9780 4.5900 ;
      RECT 12.8440 3.4965 12.8700 4.5900 ;
      RECT 12.7360 3.4965 12.7620 4.5900 ;
      RECT 12.6280 3.4965 12.6540 4.5900 ;
      RECT 12.5200 3.4965 12.5460 4.5900 ;
      RECT 12.4120 3.4965 12.4380 4.5900 ;
      RECT 12.3040 3.4965 12.3300 4.5900 ;
      RECT 12.1960 3.4965 12.2220 4.5900 ;
      RECT 12.0880 3.4965 12.1140 4.5900 ;
      RECT 11.9800 3.4965 12.0060 4.5900 ;
      RECT 11.8720 3.4965 11.8980 4.5900 ;
      RECT 11.7640 3.4965 11.7900 4.5900 ;
      RECT 11.6560 3.4965 11.6820 4.5900 ;
      RECT 11.5480 3.4965 11.5740 4.5900 ;
      RECT 11.4400 3.4965 11.4660 4.5900 ;
      RECT 11.3320 3.4965 11.3580 4.5900 ;
      RECT 11.2240 3.4965 11.2500 4.5900 ;
      RECT 11.1160 3.4965 11.1420 4.5900 ;
      RECT 11.0080 3.4965 11.0340 4.5900 ;
      RECT 10.9000 3.4965 10.9260 4.5900 ;
      RECT 10.7920 3.4965 10.8180 4.5900 ;
      RECT 10.6840 3.4965 10.7100 4.5900 ;
      RECT 10.5760 3.4965 10.6020 4.5900 ;
      RECT 10.4680 3.4965 10.4940 4.5900 ;
      RECT 10.3600 3.4965 10.3860 4.5900 ;
      RECT 10.2520 3.4965 10.2780 4.5900 ;
      RECT 10.1440 3.4965 10.1700 4.5900 ;
      RECT 10.0360 3.4965 10.0620 4.5900 ;
      RECT 9.9280 3.4965 9.9540 4.5900 ;
      RECT 9.8200 3.4965 9.8460 4.5900 ;
      RECT 9.7120 3.4965 9.7380 4.5900 ;
      RECT 9.6040 3.4965 9.6300 4.5900 ;
      RECT 9.4960 3.4965 9.5220 4.5900 ;
      RECT 9.3880 3.4965 9.4140 4.5900 ;
      RECT 9.2800 3.4965 9.3060 4.5900 ;
      RECT 9.1720 3.4965 9.1980 4.5900 ;
      RECT 9.0640 3.4965 9.0900 4.5900 ;
      RECT 8.9560 3.4965 8.9820 4.5900 ;
      RECT 8.8480 3.4965 8.8740 4.5900 ;
      RECT 8.7400 3.4965 8.7660 4.5900 ;
      RECT 8.6320 3.4965 8.6580 4.5900 ;
      RECT 8.5240 3.4965 8.5500 4.5900 ;
      RECT 8.4160 3.4965 8.4420 4.5900 ;
      RECT 8.3080 3.4965 8.3340 4.5900 ;
      RECT 8.2000 3.4965 8.2260 4.5900 ;
      RECT 8.0920 3.4965 8.1180 4.5900 ;
      RECT 7.9840 3.4965 8.0100 4.5900 ;
      RECT 7.8760 3.4965 7.9020 4.5900 ;
      RECT 7.7680 3.4965 7.7940 4.5900 ;
      RECT 7.6600 3.4965 7.6860 4.5900 ;
      RECT 7.5520 3.4965 7.5780 4.5900 ;
      RECT 7.4440 3.4965 7.4700 4.5900 ;
      RECT 7.3360 3.4965 7.3620 4.5900 ;
      RECT 7.2280 3.4965 7.2540 4.5900 ;
      RECT 7.1200 3.4965 7.1460 4.5900 ;
      RECT 7.0120 3.4965 7.0380 4.5900 ;
      RECT 6.9040 3.4965 6.9300 4.5900 ;
      RECT 6.7960 3.4965 6.8220 4.5900 ;
      RECT 6.6880 3.4965 6.7140 4.5900 ;
      RECT 6.5800 3.4965 6.6060 4.5900 ;
      RECT 6.4720 3.4965 6.4980 4.5900 ;
      RECT 6.3640 3.4965 6.3900 4.5900 ;
      RECT 6.2560 3.4965 6.2820 4.5900 ;
      RECT 6.1480 3.4965 6.1740 4.5900 ;
      RECT 6.0400 3.4965 6.0660 4.5900 ;
      RECT 5.9320 3.4965 5.9580 4.5900 ;
      RECT 5.8240 3.4965 5.8500 4.5900 ;
      RECT 5.7160 3.4965 5.7420 4.5900 ;
      RECT 5.6080 3.4965 5.6340 4.5900 ;
      RECT 5.5000 3.4965 5.5260 4.5900 ;
      RECT 5.3920 3.4965 5.4180 4.5900 ;
      RECT 5.2840 3.4965 5.3100 4.5900 ;
      RECT 5.1760 3.4965 5.2020 4.5900 ;
      RECT 5.0680 3.4965 5.0940 4.5900 ;
      RECT 4.9600 3.4965 4.9860 4.5900 ;
      RECT 4.8520 3.4965 4.8780 4.5900 ;
      RECT 4.7440 3.4965 4.7700 4.5900 ;
      RECT 4.6360 3.4965 4.6620 4.5900 ;
      RECT 4.5280 3.4965 4.5540 4.5900 ;
      RECT 4.4200 3.4965 4.4460 4.5900 ;
      RECT 4.3120 3.4965 4.3380 4.5900 ;
      RECT 4.2040 3.4965 4.2300 4.5900 ;
      RECT 4.0960 3.4965 4.1220 4.5900 ;
      RECT 3.9880 3.4965 4.0140 4.5900 ;
      RECT 3.8800 3.4965 3.9060 4.5900 ;
      RECT 3.7720 3.4965 3.7980 4.5900 ;
      RECT 3.6640 3.4965 3.6900 4.5900 ;
      RECT 3.5560 3.4965 3.5820 4.5900 ;
      RECT 3.4480 3.4965 3.4740 4.5900 ;
      RECT 3.3400 3.4965 3.3660 4.5900 ;
      RECT 3.2320 3.4965 3.2580 4.5900 ;
      RECT 3.1240 3.4965 3.1500 4.5900 ;
      RECT 3.0160 3.4965 3.0420 4.5900 ;
      RECT 2.9080 3.4965 2.9340 4.5900 ;
      RECT 2.8000 3.4965 2.8260 4.5900 ;
      RECT 2.6920 3.4965 2.7180 4.5900 ;
      RECT 2.5840 3.4965 2.6100 4.5900 ;
      RECT 2.4760 3.4965 2.5020 4.5900 ;
      RECT 2.3680 3.4965 2.3940 4.5900 ;
      RECT 2.2600 3.4965 2.2860 4.5900 ;
      RECT 2.1520 3.4965 2.1780 4.5900 ;
      RECT 2.0440 3.4965 2.0700 4.5900 ;
      RECT 1.9360 3.4965 1.9620 4.5900 ;
      RECT 1.8280 3.4965 1.8540 4.5900 ;
      RECT 1.7200 3.4965 1.7460 4.5900 ;
      RECT 1.6120 3.4965 1.6380 4.5900 ;
      RECT 1.5040 3.4965 1.5300 4.5900 ;
      RECT 1.3960 3.4965 1.4220 4.5900 ;
      RECT 1.2880 3.4965 1.3140 4.5900 ;
      RECT 1.1800 3.4965 1.2060 4.5900 ;
      RECT 1.0720 3.4965 1.0980 4.5900 ;
      RECT 0.9640 3.4965 0.9900 4.5900 ;
      RECT 0.8560 3.4965 0.8820 4.5900 ;
      RECT 0.7480 3.4965 0.7740 4.5900 ;
      RECT 0.6400 3.4965 0.6660 4.5900 ;
      RECT 0.5320 3.4965 0.5580 4.5900 ;
      RECT 0.4240 3.4965 0.4500 4.5900 ;
      RECT 0.3160 3.4965 0.3420 4.5900 ;
      RECT 0.2080 3.4965 0.2340 4.5900 ;
      RECT 0.0050 3.4965 0.0900 4.5900 ;
      RECT 15.5530 4.5765 15.6810 5.6700 ;
      RECT 15.5390 5.2420 15.6810 5.5645 ;
      RECT 15.3190 4.9690 15.4530 5.6700 ;
      RECT 15.2960 5.3040 15.4530 5.5620 ;
      RECT 15.3190 4.5765 15.4170 5.6700 ;
      RECT 15.3190 4.6975 15.4310 4.9370 ;
      RECT 15.3190 4.5765 15.4530 4.6655 ;
      RECT 15.0940 5.0270 15.2280 5.6700 ;
      RECT 15.0940 4.5765 15.1920 5.6700 ;
      RECT 14.6770 4.5765 14.7600 5.6700 ;
      RECT 14.6770 4.6650 14.7740 5.6005 ;
      RECT 30.2680 4.5765 30.3530 5.6700 ;
      RECT 30.1240 4.5765 30.1500 5.6700 ;
      RECT 30.0160 4.5765 30.0420 5.6700 ;
      RECT 29.9080 4.5765 29.9340 5.6700 ;
      RECT 29.8000 4.5765 29.8260 5.6700 ;
      RECT 29.6920 4.5765 29.7180 5.6700 ;
      RECT 29.5840 4.5765 29.6100 5.6700 ;
      RECT 29.4760 4.5765 29.5020 5.6700 ;
      RECT 29.3680 4.5765 29.3940 5.6700 ;
      RECT 29.2600 4.5765 29.2860 5.6700 ;
      RECT 29.1520 4.5765 29.1780 5.6700 ;
      RECT 29.0440 4.5765 29.0700 5.6700 ;
      RECT 28.9360 4.5765 28.9620 5.6700 ;
      RECT 28.8280 4.5765 28.8540 5.6700 ;
      RECT 28.7200 4.5765 28.7460 5.6700 ;
      RECT 28.6120 4.5765 28.6380 5.6700 ;
      RECT 28.5040 4.5765 28.5300 5.6700 ;
      RECT 28.3960 4.5765 28.4220 5.6700 ;
      RECT 28.2880 4.5765 28.3140 5.6700 ;
      RECT 28.1800 4.5765 28.2060 5.6700 ;
      RECT 28.0720 4.5765 28.0980 5.6700 ;
      RECT 27.9640 4.5765 27.9900 5.6700 ;
      RECT 27.8560 4.5765 27.8820 5.6700 ;
      RECT 27.7480 4.5765 27.7740 5.6700 ;
      RECT 27.6400 4.5765 27.6660 5.6700 ;
      RECT 27.5320 4.5765 27.5580 5.6700 ;
      RECT 27.4240 4.5765 27.4500 5.6700 ;
      RECT 27.3160 4.5765 27.3420 5.6700 ;
      RECT 27.2080 4.5765 27.2340 5.6700 ;
      RECT 27.1000 4.5765 27.1260 5.6700 ;
      RECT 26.9920 4.5765 27.0180 5.6700 ;
      RECT 26.8840 4.5765 26.9100 5.6700 ;
      RECT 26.7760 4.5765 26.8020 5.6700 ;
      RECT 26.6680 4.5765 26.6940 5.6700 ;
      RECT 26.5600 4.5765 26.5860 5.6700 ;
      RECT 26.4520 4.5765 26.4780 5.6700 ;
      RECT 26.3440 4.5765 26.3700 5.6700 ;
      RECT 26.2360 4.5765 26.2620 5.6700 ;
      RECT 26.1280 4.5765 26.1540 5.6700 ;
      RECT 26.0200 4.5765 26.0460 5.6700 ;
      RECT 25.9120 4.5765 25.9380 5.6700 ;
      RECT 25.8040 4.5765 25.8300 5.6700 ;
      RECT 25.6960 4.5765 25.7220 5.6700 ;
      RECT 25.5880 4.5765 25.6140 5.6700 ;
      RECT 25.4800 4.5765 25.5060 5.6700 ;
      RECT 25.3720 4.5765 25.3980 5.6700 ;
      RECT 25.2640 4.5765 25.2900 5.6700 ;
      RECT 25.1560 4.5765 25.1820 5.6700 ;
      RECT 25.0480 4.5765 25.0740 5.6700 ;
      RECT 24.9400 4.5765 24.9660 5.6700 ;
      RECT 24.8320 4.5765 24.8580 5.6700 ;
      RECT 24.7240 4.5765 24.7500 5.6700 ;
      RECT 24.6160 4.5765 24.6420 5.6700 ;
      RECT 24.5080 4.5765 24.5340 5.6700 ;
      RECT 24.4000 4.5765 24.4260 5.6700 ;
      RECT 24.2920 4.5765 24.3180 5.6700 ;
      RECT 24.1840 4.5765 24.2100 5.6700 ;
      RECT 24.0760 4.5765 24.1020 5.6700 ;
      RECT 23.9680 4.5765 23.9940 5.6700 ;
      RECT 23.8600 4.5765 23.8860 5.6700 ;
      RECT 23.7520 4.5765 23.7780 5.6700 ;
      RECT 23.6440 4.5765 23.6700 5.6700 ;
      RECT 23.5360 4.5765 23.5620 5.6700 ;
      RECT 23.4280 4.5765 23.4540 5.6700 ;
      RECT 23.3200 4.5765 23.3460 5.6700 ;
      RECT 23.2120 4.5765 23.2380 5.6700 ;
      RECT 23.1040 4.5765 23.1300 5.6700 ;
      RECT 22.9960 4.5765 23.0220 5.6700 ;
      RECT 22.8880 4.5765 22.9140 5.6700 ;
      RECT 22.7800 4.5765 22.8060 5.6700 ;
      RECT 22.6720 4.5765 22.6980 5.6700 ;
      RECT 22.5640 4.5765 22.5900 5.6700 ;
      RECT 22.4560 4.5765 22.4820 5.6700 ;
      RECT 22.3480 4.5765 22.3740 5.6700 ;
      RECT 22.2400 4.5765 22.2660 5.6700 ;
      RECT 22.1320 4.5765 22.1580 5.6700 ;
      RECT 22.0240 4.5765 22.0500 5.6700 ;
      RECT 21.9160 4.5765 21.9420 5.6700 ;
      RECT 21.8080 4.5765 21.8340 5.6700 ;
      RECT 21.7000 4.5765 21.7260 5.6700 ;
      RECT 21.5920 4.5765 21.6180 5.6700 ;
      RECT 21.4840 4.5765 21.5100 5.6700 ;
      RECT 21.3760 4.5765 21.4020 5.6700 ;
      RECT 21.2680 4.5765 21.2940 5.6700 ;
      RECT 21.1600 4.5765 21.1860 5.6700 ;
      RECT 21.0520 4.5765 21.0780 5.6700 ;
      RECT 20.9440 4.5765 20.9700 5.6700 ;
      RECT 20.8360 4.5765 20.8620 5.6700 ;
      RECT 20.7280 4.5765 20.7540 5.6700 ;
      RECT 20.6200 4.5765 20.6460 5.6700 ;
      RECT 20.5120 4.5765 20.5380 5.6700 ;
      RECT 20.4040 4.5765 20.4300 5.6700 ;
      RECT 20.2960 4.5765 20.3220 5.6700 ;
      RECT 20.1880 4.5765 20.2140 5.6700 ;
      RECT 20.0800 4.5765 20.1060 5.6700 ;
      RECT 19.9720 4.5765 19.9980 5.6700 ;
      RECT 19.8640 4.5765 19.8900 5.6700 ;
      RECT 19.7560 4.5765 19.7820 5.6700 ;
      RECT 19.6480 4.5765 19.6740 5.6700 ;
      RECT 19.5400 4.5765 19.5660 5.6700 ;
      RECT 19.4320 4.5765 19.4580 5.6700 ;
      RECT 19.3240 4.5765 19.3500 5.6700 ;
      RECT 19.2160 4.5765 19.2420 5.6700 ;
      RECT 19.1080 4.5765 19.1340 5.6700 ;
      RECT 19.0000 4.5765 19.0260 5.6700 ;
      RECT 18.8920 4.5765 18.9180 5.6700 ;
      RECT 18.7840 4.5765 18.8100 5.6700 ;
      RECT 18.6760 4.5765 18.7020 5.6700 ;
      RECT 18.5680 4.5765 18.5940 5.6700 ;
      RECT 18.4600 4.5765 18.4860 5.6700 ;
      RECT 18.3520 4.5765 18.3780 5.6700 ;
      RECT 18.2440 4.5765 18.2700 5.6700 ;
      RECT 18.1360 4.5765 18.1620 5.6700 ;
      RECT 18.0280 4.5765 18.0540 5.6700 ;
      RECT 17.9200 4.5765 17.9460 5.6700 ;
      RECT 17.8120 4.5765 17.8380 5.6700 ;
      RECT 17.7040 4.5765 17.7300 5.6700 ;
      RECT 17.5960 4.5765 17.6220 5.6700 ;
      RECT 17.4880 4.5765 17.5140 5.6700 ;
      RECT 17.3800 4.5765 17.4060 5.6700 ;
      RECT 17.2720 4.5765 17.2980 5.6700 ;
      RECT 17.1640 4.5765 17.1900 5.6700 ;
      RECT 17.0560 4.5765 17.0820 5.6700 ;
      RECT 16.9480 4.5765 16.9740 5.6700 ;
      RECT 16.8400 4.5765 16.8660 5.6700 ;
      RECT 16.7320 4.5765 16.7580 5.6700 ;
      RECT 16.6240 4.5765 16.6500 5.6700 ;
      RECT 16.5160 4.5765 16.5420 5.6700 ;
      RECT 16.4080 4.5765 16.4340 5.6700 ;
      RECT 16.3000 4.5765 16.3260 5.6700 ;
      RECT 16.0870 4.5765 16.1640 5.6700 ;
      RECT 14.1940 4.5765 14.2710 5.6700 ;
      RECT 14.0320 4.5765 14.0580 5.6700 ;
      RECT 13.9240 4.5765 13.9500 5.6700 ;
      RECT 13.8160 4.5765 13.8420 5.6700 ;
      RECT 13.7080 4.5765 13.7340 5.6700 ;
      RECT 13.6000 4.5765 13.6260 5.6700 ;
      RECT 13.4920 4.5765 13.5180 5.6700 ;
      RECT 13.3840 4.5765 13.4100 5.6700 ;
      RECT 13.2760 4.5765 13.3020 5.6700 ;
      RECT 13.1680 4.5765 13.1940 5.6700 ;
      RECT 13.0600 4.5765 13.0860 5.6700 ;
      RECT 12.9520 4.5765 12.9780 5.6700 ;
      RECT 12.8440 4.5765 12.8700 5.6700 ;
      RECT 12.7360 4.5765 12.7620 5.6700 ;
      RECT 12.6280 4.5765 12.6540 5.6700 ;
      RECT 12.5200 4.5765 12.5460 5.6700 ;
      RECT 12.4120 4.5765 12.4380 5.6700 ;
      RECT 12.3040 4.5765 12.3300 5.6700 ;
      RECT 12.1960 4.5765 12.2220 5.6700 ;
      RECT 12.0880 4.5765 12.1140 5.6700 ;
      RECT 11.9800 4.5765 12.0060 5.6700 ;
      RECT 11.8720 4.5765 11.8980 5.6700 ;
      RECT 11.7640 4.5765 11.7900 5.6700 ;
      RECT 11.6560 4.5765 11.6820 5.6700 ;
      RECT 11.5480 4.5765 11.5740 5.6700 ;
      RECT 11.4400 4.5765 11.4660 5.6700 ;
      RECT 11.3320 4.5765 11.3580 5.6700 ;
      RECT 11.2240 4.5765 11.2500 5.6700 ;
      RECT 11.1160 4.5765 11.1420 5.6700 ;
      RECT 11.0080 4.5765 11.0340 5.6700 ;
      RECT 10.9000 4.5765 10.9260 5.6700 ;
      RECT 10.7920 4.5765 10.8180 5.6700 ;
      RECT 10.6840 4.5765 10.7100 5.6700 ;
      RECT 10.5760 4.5765 10.6020 5.6700 ;
      RECT 10.4680 4.5765 10.4940 5.6700 ;
      RECT 10.3600 4.5765 10.3860 5.6700 ;
      RECT 10.2520 4.5765 10.2780 5.6700 ;
      RECT 10.1440 4.5765 10.1700 5.6700 ;
      RECT 10.0360 4.5765 10.0620 5.6700 ;
      RECT 9.9280 4.5765 9.9540 5.6700 ;
      RECT 9.8200 4.5765 9.8460 5.6700 ;
      RECT 9.7120 4.5765 9.7380 5.6700 ;
      RECT 9.6040 4.5765 9.6300 5.6700 ;
      RECT 9.4960 4.5765 9.5220 5.6700 ;
      RECT 9.3880 4.5765 9.4140 5.6700 ;
      RECT 9.2800 4.5765 9.3060 5.6700 ;
      RECT 9.1720 4.5765 9.1980 5.6700 ;
      RECT 9.0640 4.5765 9.0900 5.6700 ;
      RECT 8.9560 4.5765 8.9820 5.6700 ;
      RECT 8.8480 4.5765 8.8740 5.6700 ;
      RECT 8.7400 4.5765 8.7660 5.6700 ;
      RECT 8.6320 4.5765 8.6580 5.6700 ;
      RECT 8.5240 4.5765 8.5500 5.6700 ;
      RECT 8.4160 4.5765 8.4420 5.6700 ;
      RECT 8.3080 4.5765 8.3340 5.6700 ;
      RECT 8.2000 4.5765 8.2260 5.6700 ;
      RECT 8.0920 4.5765 8.1180 5.6700 ;
      RECT 7.9840 4.5765 8.0100 5.6700 ;
      RECT 7.8760 4.5765 7.9020 5.6700 ;
      RECT 7.7680 4.5765 7.7940 5.6700 ;
      RECT 7.6600 4.5765 7.6860 5.6700 ;
      RECT 7.5520 4.5765 7.5780 5.6700 ;
      RECT 7.4440 4.5765 7.4700 5.6700 ;
      RECT 7.3360 4.5765 7.3620 5.6700 ;
      RECT 7.2280 4.5765 7.2540 5.6700 ;
      RECT 7.1200 4.5765 7.1460 5.6700 ;
      RECT 7.0120 4.5765 7.0380 5.6700 ;
      RECT 6.9040 4.5765 6.9300 5.6700 ;
      RECT 6.7960 4.5765 6.8220 5.6700 ;
      RECT 6.6880 4.5765 6.7140 5.6700 ;
      RECT 6.5800 4.5765 6.6060 5.6700 ;
      RECT 6.4720 4.5765 6.4980 5.6700 ;
      RECT 6.3640 4.5765 6.3900 5.6700 ;
      RECT 6.2560 4.5765 6.2820 5.6700 ;
      RECT 6.1480 4.5765 6.1740 5.6700 ;
      RECT 6.0400 4.5765 6.0660 5.6700 ;
      RECT 5.9320 4.5765 5.9580 5.6700 ;
      RECT 5.8240 4.5765 5.8500 5.6700 ;
      RECT 5.7160 4.5765 5.7420 5.6700 ;
      RECT 5.6080 4.5765 5.6340 5.6700 ;
      RECT 5.5000 4.5765 5.5260 5.6700 ;
      RECT 5.3920 4.5765 5.4180 5.6700 ;
      RECT 5.2840 4.5765 5.3100 5.6700 ;
      RECT 5.1760 4.5765 5.2020 5.6700 ;
      RECT 5.0680 4.5765 5.0940 5.6700 ;
      RECT 4.9600 4.5765 4.9860 5.6700 ;
      RECT 4.8520 4.5765 4.8780 5.6700 ;
      RECT 4.7440 4.5765 4.7700 5.6700 ;
      RECT 4.6360 4.5765 4.6620 5.6700 ;
      RECT 4.5280 4.5765 4.5540 5.6700 ;
      RECT 4.4200 4.5765 4.4460 5.6700 ;
      RECT 4.3120 4.5765 4.3380 5.6700 ;
      RECT 4.2040 4.5765 4.2300 5.6700 ;
      RECT 4.0960 4.5765 4.1220 5.6700 ;
      RECT 3.9880 4.5765 4.0140 5.6700 ;
      RECT 3.8800 4.5765 3.9060 5.6700 ;
      RECT 3.7720 4.5765 3.7980 5.6700 ;
      RECT 3.6640 4.5765 3.6900 5.6700 ;
      RECT 3.5560 4.5765 3.5820 5.6700 ;
      RECT 3.4480 4.5765 3.4740 5.6700 ;
      RECT 3.3400 4.5765 3.3660 5.6700 ;
      RECT 3.2320 4.5765 3.2580 5.6700 ;
      RECT 3.1240 4.5765 3.1500 5.6700 ;
      RECT 3.0160 4.5765 3.0420 5.6700 ;
      RECT 2.9080 4.5765 2.9340 5.6700 ;
      RECT 2.8000 4.5765 2.8260 5.6700 ;
      RECT 2.6920 4.5765 2.7180 5.6700 ;
      RECT 2.5840 4.5765 2.6100 5.6700 ;
      RECT 2.4760 4.5765 2.5020 5.6700 ;
      RECT 2.3680 4.5765 2.3940 5.6700 ;
      RECT 2.2600 4.5765 2.2860 5.6700 ;
      RECT 2.1520 4.5765 2.1780 5.6700 ;
      RECT 2.0440 4.5765 2.0700 5.6700 ;
      RECT 1.9360 4.5765 1.9620 5.6700 ;
      RECT 1.8280 4.5765 1.8540 5.6700 ;
      RECT 1.7200 4.5765 1.7460 5.6700 ;
      RECT 1.6120 4.5765 1.6380 5.6700 ;
      RECT 1.5040 4.5765 1.5300 5.6700 ;
      RECT 1.3960 4.5765 1.4220 5.6700 ;
      RECT 1.2880 4.5765 1.3140 5.6700 ;
      RECT 1.1800 4.5765 1.2060 5.6700 ;
      RECT 1.0720 4.5765 1.0980 5.6700 ;
      RECT 0.9640 4.5765 0.9900 5.6700 ;
      RECT 0.8560 4.5765 0.8820 5.6700 ;
      RECT 0.7480 4.5765 0.7740 5.6700 ;
      RECT 0.6400 4.5765 0.6660 5.6700 ;
      RECT 0.5320 4.5765 0.5580 5.6700 ;
      RECT 0.4240 4.5765 0.4500 5.6700 ;
      RECT 0.3160 4.5765 0.3420 5.6700 ;
      RECT 0.2080 4.5765 0.2340 5.6700 ;
      RECT 0.0050 4.5765 0.0900 5.6700 ;
      RECT 15.5530 5.6565 15.6810 6.7500 ;
      RECT 15.5390 6.3220 15.6810 6.6445 ;
      RECT 15.3190 6.0490 15.4530 6.7500 ;
      RECT 15.2960 6.3840 15.4530 6.6420 ;
      RECT 15.3190 5.6565 15.4170 6.7500 ;
      RECT 15.3190 5.7775 15.4310 6.0170 ;
      RECT 15.3190 5.6565 15.4530 5.7455 ;
      RECT 15.0940 6.1070 15.2280 6.7500 ;
      RECT 15.0940 5.6565 15.1920 6.7500 ;
      RECT 14.6770 5.6565 14.7600 6.7500 ;
      RECT 14.6770 5.7450 14.7740 6.6805 ;
      RECT 30.2680 5.6565 30.3530 6.7500 ;
      RECT 30.1240 5.6565 30.1500 6.7500 ;
      RECT 30.0160 5.6565 30.0420 6.7500 ;
      RECT 29.9080 5.6565 29.9340 6.7500 ;
      RECT 29.8000 5.6565 29.8260 6.7500 ;
      RECT 29.6920 5.6565 29.7180 6.7500 ;
      RECT 29.5840 5.6565 29.6100 6.7500 ;
      RECT 29.4760 5.6565 29.5020 6.7500 ;
      RECT 29.3680 5.6565 29.3940 6.7500 ;
      RECT 29.2600 5.6565 29.2860 6.7500 ;
      RECT 29.1520 5.6565 29.1780 6.7500 ;
      RECT 29.0440 5.6565 29.0700 6.7500 ;
      RECT 28.9360 5.6565 28.9620 6.7500 ;
      RECT 28.8280 5.6565 28.8540 6.7500 ;
      RECT 28.7200 5.6565 28.7460 6.7500 ;
      RECT 28.6120 5.6565 28.6380 6.7500 ;
      RECT 28.5040 5.6565 28.5300 6.7500 ;
      RECT 28.3960 5.6565 28.4220 6.7500 ;
      RECT 28.2880 5.6565 28.3140 6.7500 ;
      RECT 28.1800 5.6565 28.2060 6.7500 ;
      RECT 28.0720 5.6565 28.0980 6.7500 ;
      RECT 27.9640 5.6565 27.9900 6.7500 ;
      RECT 27.8560 5.6565 27.8820 6.7500 ;
      RECT 27.7480 5.6565 27.7740 6.7500 ;
      RECT 27.6400 5.6565 27.6660 6.7500 ;
      RECT 27.5320 5.6565 27.5580 6.7500 ;
      RECT 27.4240 5.6565 27.4500 6.7500 ;
      RECT 27.3160 5.6565 27.3420 6.7500 ;
      RECT 27.2080 5.6565 27.2340 6.7500 ;
      RECT 27.1000 5.6565 27.1260 6.7500 ;
      RECT 26.9920 5.6565 27.0180 6.7500 ;
      RECT 26.8840 5.6565 26.9100 6.7500 ;
      RECT 26.7760 5.6565 26.8020 6.7500 ;
      RECT 26.6680 5.6565 26.6940 6.7500 ;
      RECT 26.5600 5.6565 26.5860 6.7500 ;
      RECT 26.4520 5.6565 26.4780 6.7500 ;
      RECT 26.3440 5.6565 26.3700 6.7500 ;
      RECT 26.2360 5.6565 26.2620 6.7500 ;
      RECT 26.1280 5.6565 26.1540 6.7500 ;
      RECT 26.0200 5.6565 26.0460 6.7500 ;
      RECT 25.9120 5.6565 25.9380 6.7500 ;
      RECT 25.8040 5.6565 25.8300 6.7500 ;
      RECT 25.6960 5.6565 25.7220 6.7500 ;
      RECT 25.5880 5.6565 25.6140 6.7500 ;
      RECT 25.4800 5.6565 25.5060 6.7500 ;
      RECT 25.3720 5.6565 25.3980 6.7500 ;
      RECT 25.2640 5.6565 25.2900 6.7500 ;
      RECT 25.1560 5.6565 25.1820 6.7500 ;
      RECT 25.0480 5.6565 25.0740 6.7500 ;
      RECT 24.9400 5.6565 24.9660 6.7500 ;
      RECT 24.8320 5.6565 24.8580 6.7500 ;
      RECT 24.7240 5.6565 24.7500 6.7500 ;
      RECT 24.6160 5.6565 24.6420 6.7500 ;
      RECT 24.5080 5.6565 24.5340 6.7500 ;
      RECT 24.4000 5.6565 24.4260 6.7500 ;
      RECT 24.2920 5.6565 24.3180 6.7500 ;
      RECT 24.1840 5.6565 24.2100 6.7500 ;
      RECT 24.0760 5.6565 24.1020 6.7500 ;
      RECT 23.9680 5.6565 23.9940 6.7500 ;
      RECT 23.8600 5.6565 23.8860 6.7500 ;
      RECT 23.7520 5.6565 23.7780 6.7500 ;
      RECT 23.6440 5.6565 23.6700 6.7500 ;
      RECT 23.5360 5.6565 23.5620 6.7500 ;
      RECT 23.4280 5.6565 23.4540 6.7500 ;
      RECT 23.3200 5.6565 23.3460 6.7500 ;
      RECT 23.2120 5.6565 23.2380 6.7500 ;
      RECT 23.1040 5.6565 23.1300 6.7500 ;
      RECT 22.9960 5.6565 23.0220 6.7500 ;
      RECT 22.8880 5.6565 22.9140 6.7500 ;
      RECT 22.7800 5.6565 22.8060 6.7500 ;
      RECT 22.6720 5.6565 22.6980 6.7500 ;
      RECT 22.5640 5.6565 22.5900 6.7500 ;
      RECT 22.4560 5.6565 22.4820 6.7500 ;
      RECT 22.3480 5.6565 22.3740 6.7500 ;
      RECT 22.2400 5.6565 22.2660 6.7500 ;
      RECT 22.1320 5.6565 22.1580 6.7500 ;
      RECT 22.0240 5.6565 22.0500 6.7500 ;
      RECT 21.9160 5.6565 21.9420 6.7500 ;
      RECT 21.8080 5.6565 21.8340 6.7500 ;
      RECT 21.7000 5.6565 21.7260 6.7500 ;
      RECT 21.5920 5.6565 21.6180 6.7500 ;
      RECT 21.4840 5.6565 21.5100 6.7500 ;
      RECT 21.3760 5.6565 21.4020 6.7500 ;
      RECT 21.2680 5.6565 21.2940 6.7500 ;
      RECT 21.1600 5.6565 21.1860 6.7500 ;
      RECT 21.0520 5.6565 21.0780 6.7500 ;
      RECT 20.9440 5.6565 20.9700 6.7500 ;
      RECT 20.8360 5.6565 20.8620 6.7500 ;
      RECT 20.7280 5.6565 20.7540 6.7500 ;
      RECT 20.6200 5.6565 20.6460 6.7500 ;
      RECT 20.5120 5.6565 20.5380 6.7500 ;
      RECT 20.4040 5.6565 20.4300 6.7500 ;
      RECT 20.2960 5.6565 20.3220 6.7500 ;
      RECT 20.1880 5.6565 20.2140 6.7500 ;
      RECT 20.0800 5.6565 20.1060 6.7500 ;
      RECT 19.9720 5.6565 19.9980 6.7500 ;
      RECT 19.8640 5.6565 19.8900 6.7500 ;
      RECT 19.7560 5.6565 19.7820 6.7500 ;
      RECT 19.6480 5.6565 19.6740 6.7500 ;
      RECT 19.5400 5.6565 19.5660 6.7500 ;
      RECT 19.4320 5.6565 19.4580 6.7500 ;
      RECT 19.3240 5.6565 19.3500 6.7500 ;
      RECT 19.2160 5.6565 19.2420 6.7500 ;
      RECT 19.1080 5.6565 19.1340 6.7500 ;
      RECT 19.0000 5.6565 19.0260 6.7500 ;
      RECT 18.8920 5.6565 18.9180 6.7500 ;
      RECT 18.7840 5.6565 18.8100 6.7500 ;
      RECT 18.6760 5.6565 18.7020 6.7500 ;
      RECT 18.5680 5.6565 18.5940 6.7500 ;
      RECT 18.4600 5.6565 18.4860 6.7500 ;
      RECT 18.3520 5.6565 18.3780 6.7500 ;
      RECT 18.2440 5.6565 18.2700 6.7500 ;
      RECT 18.1360 5.6565 18.1620 6.7500 ;
      RECT 18.0280 5.6565 18.0540 6.7500 ;
      RECT 17.9200 5.6565 17.9460 6.7500 ;
      RECT 17.8120 5.6565 17.8380 6.7500 ;
      RECT 17.7040 5.6565 17.7300 6.7500 ;
      RECT 17.5960 5.6565 17.6220 6.7500 ;
      RECT 17.4880 5.6565 17.5140 6.7500 ;
      RECT 17.3800 5.6565 17.4060 6.7500 ;
      RECT 17.2720 5.6565 17.2980 6.7500 ;
      RECT 17.1640 5.6565 17.1900 6.7500 ;
      RECT 17.0560 5.6565 17.0820 6.7500 ;
      RECT 16.9480 5.6565 16.9740 6.7500 ;
      RECT 16.8400 5.6565 16.8660 6.7500 ;
      RECT 16.7320 5.6565 16.7580 6.7500 ;
      RECT 16.6240 5.6565 16.6500 6.7500 ;
      RECT 16.5160 5.6565 16.5420 6.7500 ;
      RECT 16.4080 5.6565 16.4340 6.7500 ;
      RECT 16.3000 5.6565 16.3260 6.7500 ;
      RECT 16.0870 5.6565 16.1640 6.7500 ;
      RECT 14.1940 5.6565 14.2710 6.7500 ;
      RECT 14.0320 5.6565 14.0580 6.7500 ;
      RECT 13.9240 5.6565 13.9500 6.7500 ;
      RECT 13.8160 5.6565 13.8420 6.7500 ;
      RECT 13.7080 5.6565 13.7340 6.7500 ;
      RECT 13.6000 5.6565 13.6260 6.7500 ;
      RECT 13.4920 5.6565 13.5180 6.7500 ;
      RECT 13.3840 5.6565 13.4100 6.7500 ;
      RECT 13.2760 5.6565 13.3020 6.7500 ;
      RECT 13.1680 5.6565 13.1940 6.7500 ;
      RECT 13.0600 5.6565 13.0860 6.7500 ;
      RECT 12.9520 5.6565 12.9780 6.7500 ;
      RECT 12.8440 5.6565 12.8700 6.7500 ;
      RECT 12.7360 5.6565 12.7620 6.7500 ;
      RECT 12.6280 5.6565 12.6540 6.7500 ;
      RECT 12.5200 5.6565 12.5460 6.7500 ;
      RECT 12.4120 5.6565 12.4380 6.7500 ;
      RECT 12.3040 5.6565 12.3300 6.7500 ;
      RECT 12.1960 5.6565 12.2220 6.7500 ;
      RECT 12.0880 5.6565 12.1140 6.7500 ;
      RECT 11.9800 5.6565 12.0060 6.7500 ;
      RECT 11.8720 5.6565 11.8980 6.7500 ;
      RECT 11.7640 5.6565 11.7900 6.7500 ;
      RECT 11.6560 5.6565 11.6820 6.7500 ;
      RECT 11.5480 5.6565 11.5740 6.7500 ;
      RECT 11.4400 5.6565 11.4660 6.7500 ;
      RECT 11.3320 5.6565 11.3580 6.7500 ;
      RECT 11.2240 5.6565 11.2500 6.7500 ;
      RECT 11.1160 5.6565 11.1420 6.7500 ;
      RECT 11.0080 5.6565 11.0340 6.7500 ;
      RECT 10.9000 5.6565 10.9260 6.7500 ;
      RECT 10.7920 5.6565 10.8180 6.7500 ;
      RECT 10.6840 5.6565 10.7100 6.7500 ;
      RECT 10.5760 5.6565 10.6020 6.7500 ;
      RECT 10.4680 5.6565 10.4940 6.7500 ;
      RECT 10.3600 5.6565 10.3860 6.7500 ;
      RECT 10.2520 5.6565 10.2780 6.7500 ;
      RECT 10.1440 5.6565 10.1700 6.7500 ;
      RECT 10.0360 5.6565 10.0620 6.7500 ;
      RECT 9.9280 5.6565 9.9540 6.7500 ;
      RECT 9.8200 5.6565 9.8460 6.7500 ;
      RECT 9.7120 5.6565 9.7380 6.7500 ;
      RECT 9.6040 5.6565 9.6300 6.7500 ;
      RECT 9.4960 5.6565 9.5220 6.7500 ;
      RECT 9.3880 5.6565 9.4140 6.7500 ;
      RECT 9.2800 5.6565 9.3060 6.7500 ;
      RECT 9.1720 5.6565 9.1980 6.7500 ;
      RECT 9.0640 5.6565 9.0900 6.7500 ;
      RECT 8.9560 5.6565 8.9820 6.7500 ;
      RECT 8.8480 5.6565 8.8740 6.7500 ;
      RECT 8.7400 5.6565 8.7660 6.7500 ;
      RECT 8.6320 5.6565 8.6580 6.7500 ;
      RECT 8.5240 5.6565 8.5500 6.7500 ;
      RECT 8.4160 5.6565 8.4420 6.7500 ;
      RECT 8.3080 5.6565 8.3340 6.7500 ;
      RECT 8.2000 5.6565 8.2260 6.7500 ;
      RECT 8.0920 5.6565 8.1180 6.7500 ;
      RECT 7.9840 5.6565 8.0100 6.7500 ;
      RECT 7.8760 5.6565 7.9020 6.7500 ;
      RECT 7.7680 5.6565 7.7940 6.7500 ;
      RECT 7.6600 5.6565 7.6860 6.7500 ;
      RECT 7.5520 5.6565 7.5780 6.7500 ;
      RECT 7.4440 5.6565 7.4700 6.7500 ;
      RECT 7.3360 5.6565 7.3620 6.7500 ;
      RECT 7.2280 5.6565 7.2540 6.7500 ;
      RECT 7.1200 5.6565 7.1460 6.7500 ;
      RECT 7.0120 5.6565 7.0380 6.7500 ;
      RECT 6.9040 5.6565 6.9300 6.7500 ;
      RECT 6.7960 5.6565 6.8220 6.7500 ;
      RECT 6.6880 5.6565 6.7140 6.7500 ;
      RECT 6.5800 5.6565 6.6060 6.7500 ;
      RECT 6.4720 5.6565 6.4980 6.7500 ;
      RECT 6.3640 5.6565 6.3900 6.7500 ;
      RECT 6.2560 5.6565 6.2820 6.7500 ;
      RECT 6.1480 5.6565 6.1740 6.7500 ;
      RECT 6.0400 5.6565 6.0660 6.7500 ;
      RECT 5.9320 5.6565 5.9580 6.7500 ;
      RECT 5.8240 5.6565 5.8500 6.7500 ;
      RECT 5.7160 5.6565 5.7420 6.7500 ;
      RECT 5.6080 5.6565 5.6340 6.7500 ;
      RECT 5.5000 5.6565 5.5260 6.7500 ;
      RECT 5.3920 5.6565 5.4180 6.7500 ;
      RECT 5.2840 5.6565 5.3100 6.7500 ;
      RECT 5.1760 5.6565 5.2020 6.7500 ;
      RECT 5.0680 5.6565 5.0940 6.7500 ;
      RECT 4.9600 5.6565 4.9860 6.7500 ;
      RECT 4.8520 5.6565 4.8780 6.7500 ;
      RECT 4.7440 5.6565 4.7700 6.7500 ;
      RECT 4.6360 5.6565 4.6620 6.7500 ;
      RECT 4.5280 5.6565 4.5540 6.7500 ;
      RECT 4.4200 5.6565 4.4460 6.7500 ;
      RECT 4.3120 5.6565 4.3380 6.7500 ;
      RECT 4.2040 5.6565 4.2300 6.7500 ;
      RECT 4.0960 5.6565 4.1220 6.7500 ;
      RECT 3.9880 5.6565 4.0140 6.7500 ;
      RECT 3.8800 5.6565 3.9060 6.7500 ;
      RECT 3.7720 5.6565 3.7980 6.7500 ;
      RECT 3.6640 5.6565 3.6900 6.7500 ;
      RECT 3.5560 5.6565 3.5820 6.7500 ;
      RECT 3.4480 5.6565 3.4740 6.7500 ;
      RECT 3.3400 5.6565 3.3660 6.7500 ;
      RECT 3.2320 5.6565 3.2580 6.7500 ;
      RECT 3.1240 5.6565 3.1500 6.7500 ;
      RECT 3.0160 5.6565 3.0420 6.7500 ;
      RECT 2.9080 5.6565 2.9340 6.7500 ;
      RECT 2.8000 5.6565 2.8260 6.7500 ;
      RECT 2.6920 5.6565 2.7180 6.7500 ;
      RECT 2.5840 5.6565 2.6100 6.7500 ;
      RECT 2.4760 5.6565 2.5020 6.7500 ;
      RECT 2.3680 5.6565 2.3940 6.7500 ;
      RECT 2.2600 5.6565 2.2860 6.7500 ;
      RECT 2.1520 5.6565 2.1780 6.7500 ;
      RECT 2.0440 5.6565 2.0700 6.7500 ;
      RECT 1.9360 5.6565 1.9620 6.7500 ;
      RECT 1.8280 5.6565 1.8540 6.7500 ;
      RECT 1.7200 5.6565 1.7460 6.7500 ;
      RECT 1.6120 5.6565 1.6380 6.7500 ;
      RECT 1.5040 5.6565 1.5300 6.7500 ;
      RECT 1.3960 5.6565 1.4220 6.7500 ;
      RECT 1.2880 5.6565 1.3140 6.7500 ;
      RECT 1.1800 5.6565 1.2060 6.7500 ;
      RECT 1.0720 5.6565 1.0980 6.7500 ;
      RECT 0.9640 5.6565 0.9900 6.7500 ;
      RECT 0.8560 5.6565 0.8820 6.7500 ;
      RECT 0.7480 5.6565 0.7740 6.7500 ;
      RECT 0.6400 5.6565 0.6660 6.7500 ;
      RECT 0.5320 5.6565 0.5580 6.7500 ;
      RECT 0.4240 5.6565 0.4500 6.7500 ;
      RECT 0.3160 5.6565 0.3420 6.7500 ;
      RECT 0.2080 5.6565 0.2340 6.7500 ;
      RECT 0.0050 5.6565 0.0900 6.7500 ;
      RECT 15.5530 6.7365 15.6810 7.8300 ;
      RECT 15.5390 7.4020 15.6810 7.7245 ;
      RECT 15.3190 7.1290 15.4530 7.8300 ;
      RECT 15.2960 7.4640 15.4530 7.7220 ;
      RECT 15.3190 6.7365 15.4170 7.8300 ;
      RECT 15.3190 6.8575 15.4310 7.0970 ;
      RECT 15.3190 6.7365 15.4530 6.8255 ;
      RECT 15.0940 7.1870 15.2280 7.8300 ;
      RECT 15.0940 6.7365 15.1920 7.8300 ;
      RECT 14.6770 6.7365 14.7600 7.8300 ;
      RECT 14.6770 6.8250 14.7740 7.7605 ;
      RECT 30.2680 6.7365 30.3530 7.8300 ;
      RECT 30.1240 6.7365 30.1500 7.8300 ;
      RECT 30.0160 6.7365 30.0420 7.8300 ;
      RECT 29.9080 6.7365 29.9340 7.8300 ;
      RECT 29.8000 6.7365 29.8260 7.8300 ;
      RECT 29.6920 6.7365 29.7180 7.8300 ;
      RECT 29.5840 6.7365 29.6100 7.8300 ;
      RECT 29.4760 6.7365 29.5020 7.8300 ;
      RECT 29.3680 6.7365 29.3940 7.8300 ;
      RECT 29.2600 6.7365 29.2860 7.8300 ;
      RECT 29.1520 6.7365 29.1780 7.8300 ;
      RECT 29.0440 6.7365 29.0700 7.8300 ;
      RECT 28.9360 6.7365 28.9620 7.8300 ;
      RECT 28.8280 6.7365 28.8540 7.8300 ;
      RECT 28.7200 6.7365 28.7460 7.8300 ;
      RECT 28.6120 6.7365 28.6380 7.8300 ;
      RECT 28.5040 6.7365 28.5300 7.8300 ;
      RECT 28.3960 6.7365 28.4220 7.8300 ;
      RECT 28.2880 6.7365 28.3140 7.8300 ;
      RECT 28.1800 6.7365 28.2060 7.8300 ;
      RECT 28.0720 6.7365 28.0980 7.8300 ;
      RECT 27.9640 6.7365 27.9900 7.8300 ;
      RECT 27.8560 6.7365 27.8820 7.8300 ;
      RECT 27.7480 6.7365 27.7740 7.8300 ;
      RECT 27.6400 6.7365 27.6660 7.8300 ;
      RECT 27.5320 6.7365 27.5580 7.8300 ;
      RECT 27.4240 6.7365 27.4500 7.8300 ;
      RECT 27.3160 6.7365 27.3420 7.8300 ;
      RECT 27.2080 6.7365 27.2340 7.8300 ;
      RECT 27.1000 6.7365 27.1260 7.8300 ;
      RECT 26.9920 6.7365 27.0180 7.8300 ;
      RECT 26.8840 6.7365 26.9100 7.8300 ;
      RECT 26.7760 6.7365 26.8020 7.8300 ;
      RECT 26.6680 6.7365 26.6940 7.8300 ;
      RECT 26.5600 6.7365 26.5860 7.8300 ;
      RECT 26.4520 6.7365 26.4780 7.8300 ;
      RECT 26.3440 6.7365 26.3700 7.8300 ;
      RECT 26.2360 6.7365 26.2620 7.8300 ;
      RECT 26.1280 6.7365 26.1540 7.8300 ;
      RECT 26.0200 6.7365 26.0460 7.8300 ;
      RECT 25.9120 6.7365 25.9380 7.8300 ;
      RECT 25.8040 6.7365 25.8300 7.8300 ;
      RECT 25.6960 6.7365 25.7220 7.8300 ;
      RECT 25.5880 6.7365 25.6140 7.8300 ;
      RECT 25.4800 6.7365 25.5060 7.8300 ;
      RECT 25.3720 6.7365 25.3980 7.8300 ;
      RECT 25.2640 6.7365 25.2900 7.8300 ;
      RECT 25.1560 6.7365 25.1820 7.8300 ;
      RECT 25.0480 6.7365 25.0740 7.8300 ;
      RECT 24.9400 6.7365 24.9660 7.8300 ;
      RECT 24.8320 6.7365 24.8580 7.8300 ;
      RECT 24.7240 6.7365 24.7500 7.8300 ;
      RECT 24.6160 6.7365 24.6420 7.8300 ;
      RECT 24.5080 6.7365 24.5340 7.8300 ;
      RECT 24.4000 6.7365 24.4260 7.8300 ;
      RECT 24.2920 6.7365 24.3180 7.8300 ;
      RECT 24.1840 6.7365 24.2100 7.8300 ;
      RECT 24.0760 6.7365 24.1020 7.8300 ;
      RECT 23.9680 6.7365 23.9940 7.8300 ;
      RECT 23.8600 6.7365 23.8860 7.8300 ;
      RECT 23.7520 6.7365 23.7780 7.8300 ;
      RECT 23.6440 6.7365 23.6700 7.8300 ;
      RECT 23.5360 6.7365 23.5620 7.8300 ;
      RECT 23.4280 6.7365 23.4540 7.8300 ;
      RECT 23.3200 6.7365 23.3460 7.8300 ;
      RECT 23.2120 6.7365 23.2380 7.8300 ;
      RECT 23.1040 6.7365 23.1300 7.8300 ;
      RECT 22.9960 6.7365 23.0220 7.8300 ;
      RECT 22.8880 6.7365 22.9140 7.8300 ;
      RECT 22.7800 6.7365 22.8060 7.8300 ;
      RECT 22.6720 6.7365 22.6980 7.8300 ;
      RECT 22.5640 6.7365 22.5900 7.8300 ;
      RECT 22.4560 6.7365 22.4820 7.8300 ;
      RECT 22.3480 6.7365 22.3740 7.8300 ;
      RECT 22.2400 6.7365 22.2660 7.8300 ;
      RECT 22.1320 6.7365 22.1580 7.8300 ;
      RECT 22.0240 6.7365 22.0500 7.8300 ;
      RECT 21.9160 6.7365 21.9420 7.8300 ;
      RECT 21.8080 6.7365 21.8340 7.8300 ;
      RECT 21.7000 6.7365 21.7260 7.8300 ;
      RECT 21.5920 6.7365 21.6180 7.8300 ;
      RECT 21.4840 6.7365 21.5100 7.8300 ;
      RECT 21.3760 6.7365 21.4020 7.8300 ;
      RECT 21.2680 6.7365 21.2940 7.8300 ;
      RECT 21.1600 6.7365 21.1860 7.8300 ;
      RECT 21.0520 6.7365 21.0780 7.8300 ;
      RECT 20.9440 6.7365 20.9700 7.8300 ;
      RECT 20.8360 6.7365 20.8620 7.8300 ;
      RECT 20.7280 6.7365 20.7540 7.8300 ;
      RECT 20.6200 6.7365 20.6460 7.8300 ;
      RECT 20.5120 6.7365 20.5380 7.8300 ;
      RECT 20.4040 6.7365 20.4300 7.8300 ;
      RECT 20.2960 6.7365 20.3220 7.8300 ;
      RECT 20.1880 6.7365 20.2140 7.8300 ;
      RECT 20.0800 6.7365 20.1060 7.8300 ;
      RECT 19.9720 6.7365 19.9980 7.8300 ;
      RECT 19.8640 6.7365 19.8900 7.8300 ;
      RECT 19.7560 6.7365 19.7820 7.8300 ;
      RECT 19.6480 6.7365 19.6740 7.8300 ;
      RECT 19.5400 6.7365 19.5660 7.8300 ;
      RECT 19.4320 6.7365 19.4580 7.8300 ;
      RECT 19.3240 6.7365 19.3500 7.8300 ;
      RECT 19.2160 6.7365 19.2420 7.8300 ;
      RECT 19.1080 6.7365 19.1340 7.8300 ;
      RECT 19.0000 6.7365 19.0260 7.8300 ;
      RECT 18.8920 6.7365 18.9180 7.8300 ;
      RECT 18.7840 6.7365 18.8100 7.8300 ;
      RECT 18.6760 6.7365 18.7020 7.8300 ;
      RECT 18.5680 6.7365 18.5940 7.8300 ;
      RECT 18.4600 6.7365 18.4860 7.8300 ;
      RECT 18.3520 6.7365 18.3780 7.8300 ;
      RECT 18.2440 6.7365 18.2700 7.8300 ;
      RECT 18.1360 6.7365 18.1620 7.8300 ;
      RECT 18.0280 6.7365 18.0540 7.8300 ;
      RECT 17.9200 6.7365 17.9460 7.8300 ;
      RECT 17.8120 6.7365 17.8380 7.8300 ;
      RECT 17.7040 6.7365 17.7300 7.8300 ;
      RECT 17.5960 6.7365 17.6220 7.8300 ;
      RECT 17.4880 6.7365 17.5140 7.8300 ;
      RECT 17.3800 6.7365 17.4060 7.8300 ;
      RECT 17.2720 6.7365 17.2980 7.8300 ;
      RECT 17.1640 6.7365 17.1900 7.8300 ;
      RECT 17.0560 6.7365 17.0820 7.8300 ;
      RECT 16.9480 6.7365 16.9740 7.8300 ;
      RECT 16.8400 6.7365 16.8660 7.8300 ;
      RECT 16.7320 6.7365 16.7580 7.8300 ;
      RECT 16.6240 6.7365 16.6500 7.8300 ;
      RECT 16.5160 6.7365 16.5420 7.8300 ;
      RECT 16.4080 6.7365 16.4340 7.8300 ;
      RECT 16.3000 6.7365 16.3260 7.8300 ;
      RECT 16.0870 6.7365 16.1640 7.8300 ;
      RECT 14.1940 6.7365 14.2710 7.8300 ;
      RECT 14.0320 6.7365 14.0580 7.8300 ;
      RECT 13.9240 6.7365 13.9500 7.8300 ;
      RECT 13.8160 6.7365 13.8420 7.8300 ;
      RECT 13.7080 6.7365 13.7340 7.8300 ;
      RECT 13.6000 6.7365 13.6260 7.8300 ;
      RECT 13.4920 6.7365 13.5180 7.8300 ;
      RECT 13.3840 6.7365 13.4100 7.8300 ;
      RECT 13.2760 6.7365 13.3020 7.8300 ;
      RECT 13.1680 6.7365 13.1940 7.8300 ;
      RECT 13.0600 6.7365 13.0860 7.8300 ;
      RECT 12.9520 6.7365 12.9780 7.8300 ;
      RECT 12.8440 6.7365 12.8700 7.8300 ;
      RECT 12.7360 6.7365 12.7620 7.8300 ;
      RECT 12.6280 6.7365 12.6540 7.8300 ;
      RECT 12.5200 6.7365 12.5460 7.8300 ;
      RECT 12.4120 6.7365 12.4380 7.8300 ;
      RECT 12.3040 6.7365 12.3300 7.8300 ;
      RECT 12.1960 6.7365 12.2220 7.8300 ;
      RECT 12.0880 6.7365 12.1140 7.8300 ;
      RECT 11.9800 6.7365 12.0060 7.8300 ;
      RECT 11.8720 6.7365 11.8980 7.8300 ;
      RECT 11.7640 6.7365 11.7900 7.8300 ;
      RECT 11.6560 6.7365 11.6820 7.8300 ;
      RECT 11.5480 6.7365 11.5740 7.8300 ;
      RECT 11.4400 6.7365 11.4660 7.8300 ;
      RECT 11.3320 6.7365 11.3580 7.8300 ;
      RECT 11.2240 6.7365 11.2500 7.8300 ;
      RECT 11.1160 6.7365 11.1420 7.8300 ;
      RECT 11.0080 6.7365 11.0340 7.8300 ;
      RECT 10.9000 6.7365 10.9260 7.8300 ;
      RECT 10.7920 6.7365 10.8180 7.8300 ;
      RECT 10.6840 6.7365 10.7100 7.8300 ;
      RECT 10.5760 6.7365 10.6020 7.8300 ;
      RECT 10.4680 6.7365 10.4940 7.8300 ;
      RECT 10.3600 6.7365 10.3860 7.8300 ;
      RECT 10.2520 6.7365 10.2780 7.8300 ;
      RECT 10.1440 6.7365 10.1700 7.8300 ;
      RECT 10.0360 6.7365 10.0620 7.8300 ;
      RECT 9.9280 6.7365 9.9540 7.8300 ;
      RECT 9.8200 6.7365 9.8460 7.8300 ;
      RECT 9.7120 6.7365 9.7380 7.8300 ;
      RECT 9.6040 6.7365 9.6300 7.8300 ;
      RECT 9.4960 6.7365 9.5220 7.8300 ;
      RECT 9.3880 6.7365 9.4140 7.8300 ;
      RECT 9.2800 6.7365 9.3060 7.8300 ;
      RECT 9.1720 6.7365 9.1980 7.8300 ;
      RECT 9.0640 6.7365 9.0900 7.8300 ;
      RECT 8.9560 6.7365 8.9820 7.8300 ;
      RECT 8.8480 6.7365 8.8740 7.8300 ;
      RECT 8.7400 6.7365 8.7660 7.8300 ;
      RECT 8.6320 6.7365 8.6580 7.8300 ;
      RECT 8.5240 6.7365 8.5500 7.8300 ;
      RECT 8.4160 6.7365 8.4420 7.8300 ;
      RECT 8.3080 6.7365 8.3340 7.8300 ;
      RECT 8.2000 6.7365 8.2260 7.8300 ;
      RECT 8.0920 6.7365 8.1180 7.8300 ;
      RECT 7.9840 6.7365 8.0100 7.8300 ;
      RECT 7.8760 6.7365 7.9020 7.8300 ;
      RECT 7.7680 6.7365 7.7940 7.8300 ;
      RECT 7.6600 6.7365 7.6860 7.8300 ;
      RECT 7.5520 6.7365 7.5780 7.8300 ;
      RECT 7.4440 6.7365 7.4700 7.8300 ;
      RECT 7.3360 6.7365 7.3620 7.8300 ;
      RECT 7.2280 6.7365 7.2540 7.8300 ;
      RECT 7.1200 6.7365 7.1460 7.8300 ;
      RECT 7.0120 6.7365 7.0380 7.8300 ;
      RECT 6.9040 6.7365 6.9300 7.8300 ;
      RECT 6.7960 6.7365 6.8220 7.8300 ;
      RECT 6.6880 6.7365 6.7140 7.8300 ;
      RECT 6.5800 6.7365 6.6060 7.8300 ;
      RECT 6.4720 6.7365 6.4980 7.8300 ;
      RECT 6.3640 6.7365 6.3900 7.8300 ;
      RECT 6.2560 6.7365 6.2820 7.8300 ;
      RECT 6.1480 6.7365 6.1740 7.8300 ;
      RECT 6.0400 6.7365 6.0660 7.8300 ;
      RECT 5.9320 6.7365 5.9580 7.8300 ;
      RECT 5.8240 6.7365 5.8500 7.8300 ;
      RECT 5.7160 6.7365 5.7420 7.8300 ;
      RECT 5.6080 6.7365 5.6340 7.8300 ;
      RECT 5.5000 6.7365 5.5260 7.8300 ;
      RECT 5.3920 6.7365 5.4180 7.8300 ;
      RECT 5.2840 6.7365 5.3100 7.8300 ;
      RECT 5.1760 6.7365 5.2020 7.8300 ;
      RECT 5.0680 6.7365 5.0940 7.8300 ;
      RECT 4.9600 6.7365 4.9860 7.8300 ;
      RECT 4.8520 6.7365 4.8780 7.8300 ;
      RECT 4.7440 6.7365 4.7700 7.8300 ;
      RECT 4.6360 6.7365 4.6620 7.8300 ;
      RECT 4.5280 6.7365 4.5540 7.8300 ;
      RECT 4.4200 6.7365 4.4460 7.8300 ;
      RECT 4.3120 6.7365 4.3380 7.8300 ;
      RECT 4.2040 6.7365 4.2300 7.8300 ;
      RECT 4.0960 6.7365 4.1220 7.8300 ;
      RECT 3.9880 6.7365 4.0140 7.8300 ;
      RECT 3.8800 6.7365 3.9060 7.8300 ;
      RECT 3.7720 6.7365 3.7980 7.8300 ;
      RECT 3.6640 6.7365 3.6900 7.8300 ;
      RECT 3.5560 6.7365 3.5820 7.8300 ;
      RECT 3.4480 6.7365 3.4740 7.8300 ;
      RECT 3.3400 6.7365 3.3660 7.8300 ;
      RECT 3.2320 6.7365 3.2580 7.8300 ;
      RECT 3.1240 6.7365 3.1500 7.8300 ;
      RECT 3.0160 6.7365 3.0420 7.8300 ;
      RECT 2.9080 6.7365 2.9340 7.8300 ;
      RECT 2.8000 6.7365 2.8260 7.8300 ;
      RECT 2.6920 6.7365 2.7180 7.8300 ;
      RECT 2.5840 6.7365 2.6100 7.8300 ;
      RECT 2.4760 6.7365 2.5020 7.8300 ;
      RECT 2.3680 6.7365 2.3940 7.8300 ;
      RECT 2.2600 6.7365 2.2860 7.8300 ;
      RECT 2.1520 6.7365 2.1780 7.8300 ;
      RECT 2.0440 6.7365 2.0700 7.8300 ;
      RECT 1.9360 6.7365 1.9620 7.8300 ;
      RECT 1.8280 6.7365 1.8540 7.8300 ;
      RECT 1.7200 6.7365 1.7460 7.8300 ;
      RECT 1.6120 6.7365 1.6380 7.8300 ;
      RECT 1.5040 6.7365 1.5300 7.8300 ;
      RECT 1.3960 6.7365 1.4220 7.8300 ;
      RECT 1.2880 6.7365 1.3140 7.8300 ;
      RECT 1.1800 6.7365 1.2060 7.8300 ;
      RECT 1.0720 6.7365 1.0980 7.8300 ;
      RECT 0.9640 6.7365 0.9900 7.8300 ;
      RECT 0.8560 6.7365 0.8820 7.8300 ;
      RECT 0.7480 6.7365 0.7740 7.8300 ;
      RECT 0.6400 6.7365 0.6660 7.8300 ;
      RECT 0.5320 6.7365 0.5580 7.8300 ;
      RECT 0.4240 6.7365 0.4500 7.8300 ;
      RECT 0.3160 6.7365 0.3420 7.8300 ;
      RECT 0.2080 6.7365 0.2340 7.8300 ;
      RECT 0.0050 6.7365 0.0900 7.8300 ;
      RECT 15.5530 7.8165 15.6810 8.9100 ;
      RECT 15.5390 8.4820 15.6810 8.8045 ;
      RECT 15.3190 8.2090 15.4530 8.9100 ;
      RECT 15.2960 8.5440 15.4530 8.8020 ;
      RECT 15.3190 7.8165 15.4170 8.9100 ;
      RECT 15.3190 7.9375 15.4310 8.1770 ;
      RECT 15.3190 7.8165 15.4530 7.9055 ;
      RECT 15.0940 8.2670 15.2280 8.9100 ;
      RECT 15.0940 7.8165 15.1920 8.9100 ;
      RECT 14.6770 7.8165 14.7600 8.9100 ;
      RECT 14.6770 7.9050 14.7740 8.8405 ;
      RECT 30.2680 7.8165 30.3530 8.9100 ;
      RECT 30.1240 7.8165 30.1500 8.9100 ;
      RECT 30.0160 7.8165 30.0420 8.9100 ;
      RECT 29.9080 7.8165 29.9340 8.9100 ;
      RECT 29.8000 7.8165 29.8260 8.9100 ;
      RECT 29.6920 7.8165 29.7180 8.9100 ;
      RECT 29.5840 7.8165 29.6100 8.9100 ;
      RECT 29.4760 7.8165 29.5020 8.9100 ;
      RECT 29.3680 7.8165 29.3940 8.9100 ;
      RECT 29.2600 7.8165 29.2860 8.9100 ;
      RECT 29.1520 7.8165 29.1780 8.9100 ;
      RECT 29.0440 7.8165 29.0700 8.9100 ;
      RECT 28.9360 7.8165 28.9620 8.9100 ;
      RECT 28.8280 7.8165 28.8540 8.9100 ;
      RECT 28.7200 7.8165 28.7460 8.9100 ;
      RECT 28.6120 7.8165 28.6380 8.9100 ;
      RECT 28.5040 7.8165 28.5300 8.9100 ;
      RECT 28.3960 7.8165 28.4220 8.9100 ;
      RECT 28.2880 7.8165 28.3140 8.9100 ;
      RECT 28.1800 7.8165 28.2060 8.9100 ;
      RECT 28.0720 7.8165 28.0980 8.9100 ;
      RECT 27.9640 7.8165 27.9900 8.9100 ;
      RECT 27.8560 7.8165 27.8820 8.9100 ;
      RECT 27.7480 7.8165 27.7740 8.9100 ;
      RECT 27.6400 7.8165 27.6660 8.9100 ;
      RECT 27.5320 7.8165 27.5580 8.9100 ;
      RECT 27.4240 7.8165 27.4500 8.9100 ;
      RECT 27.3160 7.8165 27.3420 8.9100 ;
      RECT 27.2080 7.8165 27.2340 8.9100 ;
      RECT 27.1000 7.8165 27.1260 8.9100 ;
      RECT 26.9920 7.8165 27.0180 8.9100 ;
      RECT 26.8840 7.8165 26.9100 8.9100 ;
      RECT 26.7760 7.8165 26.8020 8.9100 ;
      RECT 26.6680 7.8165 26.6940 8.9100 ;
      RECT 26.5600 7.8165 26.5860 8.9100 ;
      RECT 26.4520 7.8165 26.4780 8.9100 ;
      RECT 26.3440 7.8165 26.3700 8.9100 ;
      RECT 26.2360 7.8165 26.2620 8.9100 ;
      RECT 26.1280 7.8165 26.1540 8.9100 ;
      RECT 26.0200 7.8165 26.0460 8.9100 ;
      RECT 25.9120 7.8165 25.9380 8.9100 ;
      RECT 25.8040 7.8165 25.8300 8.9100 ;
      RECT 25.6960 7.8165 25.7220 8.9100 ;
      RECT 25.5880 7.8165 25.6140 8.9100 ;
      RECT 25.4800 7.8165 25.5060 8.9100 ;
      RECT 25.3720 7.8165 25.3980 8.9100 ;
      RECT 25.2640 7.8165 25.2900 8.9100 ;
      RECT 25.1560 7.8165 25.1820 8.9100 ;
      RECT 25.0480 7.8165 25.0740 8.9100 ;
      RECT 24.9400 7.8165 24.9660 8.9100 ;
      RECT 24.8320 7.8165 24.8580 8.9100 ;
      RECT 24.7240 7.8165 24.7500 8.9100 ;
      RECT 24.6160 7.8165 24.6420 8.9100 ;
      RECT 24.5080 7.8165 24.5340 8.9100 ;
      RECT 24.4000 7.8165 24.4260 8.9100 ;
      RECT 24.2920 7.8165 24.3180 8.9100 ;
      RECT 24.1840 7.8165 24.2100 8.9100 ;
      RECT 24.0760 7.8165 24.1020 8.9100 ;
      RECT 23.9680 7.8165 23.9940 8.9100 ;
      RECT 23.8600 7.8165 23.8860 8.9100 ;
      RECT 23.7520 7.8165 23.7780 8.9100 ;
      RECT 23.6440 7.8165 23.6700 8.9100 ;
      RECT 23.5360 7.8165 23.5620 8.9100 ;
      RECT 23.4280 7.8165 23.4540 8.9100 ;
      RECT 23.3200 7.8165 23.3460 8.9100 ;
      RECT 23.2120 7.8165 23.2380 8.9100 ;
      RECT 23.1040 7.8165 23.1300 8.9100 ;
      RECT 22.9960 7.8165 23.0220 8.9100 ;
      RECT 22.8880 7.8165 22.9140 8.9100 ;
      RECT 22.7800 7.8165 22.8060 8.9100 ;
      RECT 22.6720 7.8165 22.6980 8.9100 ;
      RECT 22.5640 7.8165 22.5900 8.9100 ;
      RECT 22.4560 7.8165 22.4820 8.9100 ;
      RECT 22.3480 7.8165 22.3740 8.9100 ;
      RECT 22.2400 7.8165 22.2660 8.9100 ;
      RECT 22.1320 7.8165 22.1580 8.9100 ;
      RECT 22.0240 7.8165 22.0500 8.9100 ;
      RECT 21.9160 7.8165 21.9420 8.9100 ;
      RECT 21.8080 7.8165 21.8340 8.9100 ;
      RECT 21.7000 7.8165 21.7260 8.9100 ;
      RECT 21.5920 7.8165 21.6180 8.9100 ;
      RECT 21.4840 7.8165 21.5100 8.9100 ;
      RECT 21.3760 7.8165 21.4020 8.9100 ;
      RECT 21.2680 7.8165 21.2940 8.9100 ;
      RECT 21.1600 7.8165 21.1860 8.9100 ;
      RECT 21.0520 7.8165 21.0780 8.9100 ;
      RECT 20.9440 7.8165 20.9700 8.9100 ;
      RECT 20.8360 7.8165 20.8620 8.9100 ;
      RECT 20.7280 7.8165 20.7540 8.9100 ;
      RECT 20.6200 7.8165 20.6460 8.9100 ;
      RECT 20.5120 7.8165 20.5380 8.9100 ;
      RECT 20.4040 7.8165 20.4300 8.9100 ;
      RECT 20.2960 7.8165 20.3220 8.9100 ;
      RECT 20.1880 7.8165 20.2140 8.9100 ;
      RECT 20.0800 7.8165 20.1060 8.9100 ;
      RECT 19.9720 7.8165 19.9980 8.9100 ;
      RECT 19.8640 7.8165 19.8900 8.9100 ;
      RECT 19.7560 7.8165 19.7820 8.9100 ;
      RECT 19.6480 7.8165 19.6740 8.9100 ;
      RECT 19.5400 7.8165 19.5660 8.9100 ;
      RECT 19.4320 7.8165 19.4580 8.9100 ;
      RECT 19.3240 7.8165 19.3500 8.9100 ;
      RECT 19.2160 7.8165 19.2420 8.9100 ;
      RECT 19.1080 7.8165 19.1340 8.9100 ;
      RECT 19.0000 7.8165 19.0260 8.9100 ;
      RECT 18.8920 7.8165 18.9180 8.9100 ;
      RECT 18.7840 7.8165 18.8100 8.9100 ;
      RECT 18.6760 7.8165 18.7020 8.9100 ;
      RECT 18.5680 7.8165 18.5940 8.9100 ;
      RECT 18.4600 7.8165 18.4860 8.9100 ;
      RECT 18.3520 7.8165 18.3780 8.9100 ;
      RECT 18.2440 7.8165 18.2700 8.9100 ;
      RECT 18.1360 7.8165 18.1620 8.9100 ;
      RECT 18.0280 7.8165 18.0540 8.9100 ;
      RECT 17.9200 7.8165 17.9460 8.9100 ;
      RECT 17.8120 7.8165 17.8380 8.9100 ;
      RECT 17.7040 7.8165 17.7300 8.9100 ;
      RECT 17.5960 7.8165 17.6220 8.9100 ;
      RECT 17.4880 7.8165 17.5140 8.9100 ;
      RECT 17.3800 7.8165 17.4060 8.9100 ;
      RECT 17.2720 7.8165 17.2980 8.9100 ;
      RECT 17.1640 7.8165 17.1900 8.9100 ;
      RECT 17.0560 7.8165 17.0820 8.9100 ;
      RECT 16.9480 7.8165 16.9740 8.9100 ;
      RECT 16.8400 7.8165 16.8660 8.9100 ;
      RECT 16.7320 7.8165 16.7580 8.9100 ;
      RECT 16.6240 7.8165 16.6500 8.9100 ;
      RECT 16.5160 7.8165 16.5420 8.9100 ;
      RECT 16.4080 7.8165 16.4340 8.9100 ;
      RECT 16.3000 7.8165 16.3260 8.9100 ;
      RECT 16.0870 7.8165 16.1640 8.9100 ;
      RECT 14.1940 7.8165 14.2710 8.9100 ;
      RECT 14.0320 7.8165 14.0580 8.9100 ;
      RECT 13.9240 7.8165 13.9500 8.9100 ;
      RECT 13.8160 7.8165 13.8420 8.9100 ;
      RECT 13.7080 7.8165 13.7340 8.9100 ;
      RECT 13.6000 7.8165 13.6260 8.9100 ;
      RECT 13.4920 7.8165 13.5180 8.9100 ;
      RECT 13.3840 7.8165 13.4100 8.9100 ;
      RECT 13.2760 7.8165 13.3020 8.9100 ;
      RECT 13.1680 7.8165 13.1940 8.9100 ;
      RECT 13.0600 7.8165 13.0860 8.9100 ;
      RECT 12.9520 7.8165 12.9780 8.9100 ;
      RECT 12.8440 7.8165 12.8700 8.9100 ;
      RECT 12.7360 7.8165 12.7620 8.9100 ;
      RECT 12.6280 7.8165 12.6540 8.9100 ;
      RECT 12.5200 7.8165 12.5460 8.9100 ;
      RECT 12.4120 7.8165 12.4380 8.9100 ;
      RECT 12.3040 7.8165 12.3300 8.9100 ;
      RECT 12.1960 7.8165 12.2220 8.9100 ;
      RECT 12.0880 7.8165 12.1140 8.9100 ;
      RECT 11.9800 7.8165 12.0060 8.9100 ;
      RECT 11.8720 7.8165 11.8980 8.9100 ;
      RECT 11.7640 7.8165 11.7900 8.9100 ;
      RECT 11.6560 7.8165 11.6820 8.9100 ;
      RECT 11.5480 7.8165 11.5740 8.9100 ;
      RECT 11.4400 7.8165 11.4660 8.9100 ;
      RECT 11.3320 7.8165 11.3580 8.9100 ;
      RECT 11.2240 7.8165 11.2500 8.9100 ;
      RECT 11.1160 7.8165 11.1420 8.9100 ;
      RECT 11.0080 7.8165 11.0340 8.9100 ;
      RECT 10.9000 7.8165 10.9260 8.9100 ;
      RECT 10.7920 7.8165 10.8180 8.9100 ;
      RECT 10.6840 7.8165 10.7100 8.9100 ;
      RECT 10.5760 7.8165 10.6020 8.9100 ;
      RECT 10.4680 7.8165 10.4940 8.9100 ;
      RECT 10.3600 7.8165 10.3860 8.9100 ;
      RECT 10.2520 7.8165 10.2780 8.9100 ;
      RECT 10.1440 7.8165 10.1700 8.9100 ;
      RECT 10.0360 7.8165 10.0620 8.9100 ;
      RECT 9.9280 7.8165 9.9540 8.9100 ;
      RECT 9.8200 7.8165 9.8460 8.9100 ;
      RECT 9.7120 7.8165 9.7380 8.9100 ;
      RECT 9.6040 7.8165 9.6300 8.9100 ;
      RECT 9.4960 7.8165 9.5220 8.9100 ;
      RECT 9.3880 7.8165 9.4140 8.9100 ;
      RECT 9.2800 7.8165 9.3060 8.9100 ;
      RECT 9.1720 7.8165 9.1980 8.9100 ;
      RECT 9.0640 7.8165 9.0900 8.9100 ;
      RECT 8.9560 7.8165 8.9820 8.9100 ;
      RECT 8.8480 7.8165 8.8740 8.9100 ;
      RECT 8.7400 7.8165 8.7660 8.9100 ;
      RECT 8.6320 7.8165 8.6580 8.9100 ;
      RECT 8.5240 7.8165 8.5500 8.9100 ;
      RECT 8.4160 7.8165 8.4420 8.9100 ;
      RECT 8.3080 7.8165 8.3340 8.9100 ;
      RECT 8.2000 7.8165 8.2260 8.9100 ;
      RECT 8.0920 7.8165 8.1180 8.9100 ;
      RECT 7.9840 7.8165 8.0100 8.9100 ;
      RECT 7.8760 7.8165 7.9020 8.9100 ;
      RECT 7.7680 7.8165 7.7940 8.9100 ;
      RECT 7.6600 7.8165 7.6860 8.9100 ;
      RECT 7.5520 7.8165 7.5780 8.9100 ;
      RECT 7.4440 7.8165 7.4700 8.9100 ;
      RECT 7.3360 7.8165 7.3620 8.9100 ;
      RECT 7.2280 7.8165 7.2540 8.9100 ;
      RECT 7.1200 7.8165 7.1460 8.9100 ;
      RECT 7.0120 7.8165 7.0380 8.9100 ;
      RECT 6.9040 7.8165 6.9300 8.9100 ;
      RECT 6.7960 7.8165 6.8220 8.9100 ;
      RECT 6.6880 7.8165 6.7140 8.9100 ;
      RECT 6.5800 7.8165 6.6060 8.9100 ;
      RECT 6.4720 7.8165 6.4980 8.9100 ;
      RECT 6.3640 7.8165 6.3900 8.9100 ;
      RECT 6.2560 7.8165 6.2820 8.9100 ;
      RECT 6.1480 7.8165 6.1740 8.9100 ;
      RECT 6.0400 7.8165 6.0660 8.9100 ;
      RECT 5.9320 7.8165 5.9580 8.9100 ;
      RECT 5.8240 7.8165 5.8500 8.9100 ;
      RECT 5.7160 7.8165 5.7420 8.9100 ;
      RECT 5.6080 7.8165 5.6340 8.9100 ;
      RECT 5.5000 7.8165 5.5260 8.9100 ;
      RECT 5.3920 7.8165 5.4180 8.9100 ;
      RECT 5.2840 7.8165 5.3100 8.9100 ;
      RECT 5.1760 7.8165 5.2020 8.9100 ;
      RECT 5.0680 7.8165 5.0940 8.9100 ;
      RECT 4.9600 7.8165 4.9860 8.9100 ;
      RECT 4.8520 7.8165 4.8780 8.9100 ;
      RECT 4.7440 7.8165 4.7700 8.9100 ;
      RECT 4.6360 7.8165 4.6620 8.9100 ;
      RECT 4.5280 7.8165 4.5540 8.9100 ;
      RECT 4.4200 7.8165 4.4460 8.9100 ;
      RECT 4.3120 7.8165 4.3380 8.9100 ;
      RECT 4.2040 7.8165 4.2300 8.9100 ;
      RECT 4.0960 7.8165 4.1220 8.9100 ;
      RECT 3.9880 7.8165 4.0140 8.9100 ;
      RECT 3.8800 7.8165 3.9060 8.9100 ;
      RECT 3.7720 7.8165 3.7980 8.9100 ;
      RECT 3.6640 7.8165 3.6900 8.9100 ;
      RECT 3.5560 7.8165 3.5820 8.9100 ;
      RECT 3.4480 7.8165 3.4740 8.9100 ;
      RECT 3.3400 7.8165 3.3660 8.9100 ;
      RECT 3.2320 7.8165 3.2580 8.9100 ;
      RECT 3.1240 7.8165 3.1500 8.9100 ;
      RECT 3.0160 7.8165 3.0420 8.9100 ;
      RECT 2.9080 7.8165 2.9340 8.9100 ;
      RECT 2.8000 7.8165 2.8260 8.9100 ;
      RECT 2.6920 7.8165 2.7180 8.9100 ;
      RECT 2.5840 7.8165 2.6100 8.9100 ;
      RECT 2.4760 7.8165 2.5020 8.9100 ;
      RECT 2.3680 7.8165 2.3940 8.9100 ;
      RECT 2.2600 7.8165 2.2860 8.9100 ;
      RECT 2.1520 7.8165 2.1780 8.9100 ;
      RECT 2.0440 7.8165 2.0700 8.9100 ;
      RECT 1.9360 7.8165 1.9620 8.9100 ;
      RECT 1.8280 7.8165 1.8540 8.9100 ;
      RECT 1.7200 7.8165 1.7460 8.9100 ;
      RECT 1.6120 7.8165 1.6380 8.9100 ;
      RECT 1.5040 7.8165 1.5300 8.9100 ;
      RECT 1.3960 7.8165 1.4220 8.9100 ;
      RECT 1.2880 7.8165 1.3140 8.9100 ;
      RECT 1.1800 7.8165 1.2060 8.9100 ;
      RECT 1.0720 7.8165 1.0980 8.9100 ;
      RECT 0.9640 7.8165 0.9900 8.9100 ;
      RECT 0.8560 7.8165 0.8820 8.9100 ;
      RECT 0.7480 7.8165 0.7740 8.9100 ;
      RECT 0.6400 7.8165 0.6660 8.9100 ;
      RECT 0.5320 7.8165 0.5580 8.9100 ;
      RECT 0.4240 7.8165 0.4500 8.9100 ;
      RECT 0.3160 7.8165 0.3420 8.9100 ;
      RECT 0.2080 7.8165 0.2340 8.9100 ;
      RECT 0.0050 7.8165 0.0900 8.9100 ;
      RECT 15.5530 8.8965 15.6810 9.9900 ;
      RECT 15.5390 9.5620 15.6810 9.8845 ;
      RECT 15.3190 9.2890 15.4530 9.9900 ;
      RECT 15.2960 9.6240 15.4530 9.8820 ;
      RECT 15.3190 8.8965 15.4170 9.9900 ;
      RECT 15.3190 9.0175 15.4310 9.2570 ;
      RECT 15.3190 8.8965 15.4530 8.9855 ;
      RECT 15.0940 9.3470 15.2280 9.9900 ;
      RECT 15.0940 8.8965 15.1920 9.9900 ;
      RECT 14.6770 8.8965 14.7600 9.9900 ;
      RECT 14.6770 8.9850 14.7740 9.9205 ;
      RECT 30.2680 8.8965 30.3530 9.9900 ;
      RECT 30.1240 8.8965 30.1500 9.9900 ;
      RECT 30.0160 8.8965 30.0420 9.9900 ;
      RECT 29.9080 8.8965 29.9340 9.9900 ;
      RECT 29.8000 8.8965 29.8260 9.9900 ;
      RECT 29.6920 8.8965 29.7180 9.9900 ;
      RECT 29.5840 8.8965 29.6100 9.9900 ;
      RECT 29.4760 8.8965 29.5020 9.9900 ;
      RECT 29.3680 8.8965 29.3940 9.9900 ;
      RECT 29.2600 8.8965 29.2860 9.9900 ;
      RECT 29.1520 8.8965 29.1780 9.9900 ;
      RECT 29.0440 8.8965 29.0700 9.9900 ;
      RECT 28.9360 8.8965 28.9620 9.9900 ;
      RECT 28.8280 8.8965 28.8540 9.9900 ;
      RECT 28.7200 8.8965 28.7460 9.9900 ;
      RECT 28.6120 8.8965 28.6380 9.9900 ;
      RECT 28.5040 8.8965 28.5300 9.9900 ;
      RECT 28.3960 8.8965 28.4220 9.9900 ;
      RECT 28.2880 8.8965 28.3140 9.9900 ;
      RECT 28.1800 8.8965 28.2060 9.9900 ;
      RECT 28.0720 8.8965 28.0980 9.9900 ;
      RECT 27.9640 8.8965 27.9900 9.9900 ;
      RECT 27.8560 8.8965 27.8820 9.9900 ;
      RECT 27.7480 8.8965 27.7740 9.9900 ;
      RECT 27.6400 8.8965 27.6660 9.9900 ;
      RECT 27.5320 8.8965 27.5580 9.9900 ;
      RECT 27.4240 8.8965 27.4500 9.9900 ;
      RECT 27.3160 8.8965 27.3420 9.9900 ;
      RECT 27.2080 8.8965 27.2340 9.9900 ;
      RECT 27.1000 8.8965 27.1260 9.9900 ;
      RECT 26.9920 8.8965 27.0180 9.9900 ;
      RECT 26.8840 8.8965 26.9100 9.9900 ;
      RECT 26.7760 8.8965 26.8020 9.9900 ;
      RECT 26.6680 8.8965 26.6940 9.9900 ;
      RECT 26.5600 8.8965 26.5860 9.9900 ;
      RECT 26.4520 8.8965 26.4780 9.9900 ;
      RECT 26.3440 8.8965 26.3700 9.9900 ;
      RECT 26.2360 8.8965 26.2620 9.9900 ;
      RECT 26.1280 8.8965 26.1540 9.9900 ;
      RECT 26.0200 8.8965 26.0460 9.9900 ;
      RECT 25.9120 8.8965 25.9380 9.9900 ;
      RECT 25.8040 8.8965 25.8300 9.9900 ;
      RECT 25.6960 8.8965 25.7220 9.9900 ;
      RECT 25.5880 8.8965 25.6140 9.9900 ;
      RECT 25.4800 8.8965 25.5060 9.9900 ;
      RECT 25.3720 8.8965 25.3980 9.9900 ;
      RECT 25.2640 8.8965 25.2900 9.9900 ;
      RECT 25.1560 8.8965 25.1820 9.9900 ;
      RECT 25.0480 8.8965 25.0740 9.9900 ;
      RECT 24.9400 8.8965 24.9660 9.9900 ;
      RECT 24.8320 8.8965 24.8580 9.9900 ;
      RECT 24.7240 8.8965 24.7500 9.9900 ;
      RECT 24.6160 8.8965 24.6420 9.9900 ;
      RECT 24.5080 8.8965 24.5340 9.9900 ;
      RECT 24.4000 8.8965 24.4260 9.9900 ;
      RECT 24.2920 8.8965 24.3180 9.9900 ;
      RECT 24.1840 8.8965 24.2100 9.9900 ;
      RECT 24.0760 8.8965 24.1020 9.9900 ;
      RECT 23.9680 8.8965 23.9940 9.9900 ;
      RECT 23.8600 8.8965 23.8860 9.9900 ;
      RECT 23.7520 8.8965 23.7780 9.9900 ;
      RECT 23.6440 8.8965 23.6700 9.9900 ;
      RECT 23.5360 8.8965 23.5620 9.9900 ;
      RECT 23.4280 8.8965 23.4540 9.9900 ;
      RECT 23.3200 8.8965 23.3460 9.9900 ;
      RECT 23.2120 8.8965 23.2380 9.9900 ;
      RECT 23.1040 8.8965 23.1300 9.9900 ;
      RECT 22.9960 8.8965 23.0220 9.9900 ;
      RECT 22.8880 8.8965 22.9140 9.9900 ;
      RECT 22.7800 8.8965 22.8060 9.9900 ;
      RECT 22.6720 8.8965 22.6980 9.9900 ;
      RECT 22.5640 8.8965 22.5900 9.9900 ;
      RECT 22.4560 8.8965 22.4820 9.9900 ;
      RECT 22.3480 8.8965 22.3740 9.9900 ;
      RECT 22.2400 8.8965 22.2660 9.9900 ;
      RECT 22.1320 8.8965 22.1580 9.9900 ;
      RECT 22.0240 8.8965 22.0500 9.9900 ;
      RECT 21.9160 8.8965 21.9420 9.9900 ;
      RECT 21.8080 8.8965 21.8340 9.9900 ;
      RECT 21.7000 8.8965 21.7260 9.9900 ;
      RECT 21.5920 8.8965 21.6180 9.9900 ;
      RECT 21.4840 8.8965 21.5100 9.9900 ;
      RECT 21.3760 8.8965 21.4020 9.9900 ;
      RECT 21.2680 8.8965 21.2940 9.9900 ;
      RECT 21.1600 8.8965 21.1860 9.9900 ;
      RECT 21.0520 8.8965 21.0780 9.9900 ;
      RECT 20.9440 8.8965 20.9700 9.9900 ;
      RECT 20.8360 8.8965 20.8620 9.9900 ;
      RECT 20.7280 8.8965 20.7540 9.9900 ;
      RECT 20.6200 8.8965 20.6460 9.9900 ;
      RECT 20.5120 8.8965 20.5380 9.9900 ;
      RECT 20.4040 8.8965 20.4300 9.9900 ;
      RECT 20.2960 8.8965 20.3220 9.9900 ;
      RECT 20.1880 8.8965 20.2140 9.9900 ;
      RECT 20.0800 8.8965 20.1060 9.9900 ;
      RECT 19.9720 8.8965 19.9980 9.9900 ;
      RECT 19.8640 8.8965 19.8900 9.9900 ;
      RECT 19.7560 8.8965 19.7820 9.9900 ;
      RECT 19.6480 8.8965 19.6740 9.9900 ;
      RECT 19.5400 8.8965 19.5660 9.9900 ;
      RECT 19.4320 8.8965 19.4580 9.9900 ;
      RECT 19.3240 8.8965 19.3500 9.9900 ;
      RECT 19.2160 8.8965 19.2420 9.9900 ;
      RECT 19.1080 8.8965 19.1340 9.9900 ;
      RECT 19.0000 8.8965 19.0260 9.9900 ;
      RECT 18.8920 8.8965 18.9180 9.9900 ;
      RECT 18.7840 8.8965 18.8100 9.9900 ;
      RECT 18.6760 8.8965 18.7020 9.9900 ;
      RECT 18.5680 8.8965 18.5940 9.9900 ;
      RECT 18.4600 8.8965 18.4860 9.9900 ;
      RECT 18.3520 8.8965 18.3780 9.9900 ;
      RECT 18.2440 8.8965 18.2700 9.9900 ;
      RECT 18.1360 8.8965 18.1620 9.9900 ;
      RECT 18.0280 8.8965 18.0540 9.9900 ;
      RECT 17.9200 8.8965 17.9460 9.9900 ;
      RECT 17.8120 8.8965 17.8380 9.9900 ;
      RECT 17.7040 8.8965 17.7300 9.9900 ;
      RECT 17.5960 8.8965 17.6220 9.9900 ;
      RECT 17.4880 8.8965 17.5140 9.9900 ;
      RECT 17.3800 8.8965 17.4060 9.9900 ;
      RECT 17.2720 8.8965 17.2980 9.9900 ;
      RECT 17.1640 8.8965 17.1900 9.9900 ;
      RECT 17.0560 8.8965 17.0820 9.9900 ;
      RECT 16.9480 8.8965 16.9740 9.9900 ;
      RECT 16.8400 8.8965 16.8660 9.9900 ;
      RECT 16.7320 8.8965 16.7580 9.9900 ;
      RECT 16.6240 8.8965 16.6500 9.9900 ;
      RECT 16.5160 8.8965 16.5420 9.9900 ;
      RECT 16.4080 8.8965 16.4340 9.9900 ;
      RECT 16.3000 8.8965 16.3260 9.9900 ;
      RECT 16.0870 8.8965 16.1640 9.9900 ;
      RECT 14.1940 8.8965 14.2710 9.9900 ;
      RECT 14.0320 8.8965 14.0580 9.9900 ;
      RECT 13.9240 8.8965 13.9500 9.9900 ;
      RECT 13.8160 8.8965 13.8420 9.9900 ;
      RECT 13.7080 8.8965 13.7340 9.9900 ;
      RECT 13.6000 8.8965 13.6260 9.9900 ;
      RECT 13.4920 8.8965 13.5180 9.9900 ;
      RECT 13.3840 8.8965 13.4100 9.9900 ;
      RECT 13.2760 8.8965 13.3020 9.9900 ;
      RECT 13.1680 8.8965 13.1940 9.9900 ;
      RECT 13.0600 8.8965 13.0860 9.9900 ;
      RECT 12.9520 8.8965 12.9780 9.9900 ;
      RECT 12.8440 8.8965 12.8700 9.9900 ;
      RECT 12.7360 8.8965 12.7620 9.9900 ;
      RECT 12.6280 8.8965 12.6540 9.9900 ;
      RECT 12.5200 8.8965 12.5460 9.9900 ;
      RECT 12.4120 8.8965 12.4380 9.9900 ;
      RECT 12.3040 8.8965 12.3300 9.9900 ;
      RECT 12.1960 8.8965 12.2220 9.9900 ;
      RECT 12.0880 8.8965 12.1140 9.9900 ;
      RECT 11.9800 8.8965 12.0060 9.9900 ;
      RECT 11.8720 8.8965 11.8980 9.9900 ;
      RECT 11.7640 8.8965 11.7900 9.9900 ;
      RECT 11.6560 8.8965 11.6820 9.9900 ;
      RECT 11.5480 8.8965 11.5740 9.9900 ;
      RECT 11.4400 8.8965 11.4660 9.9900 ;
      RECT 11.3320 8.8965 11.3580 9.9900 ;
      RECT 11.2240 8.8965 11.2500 9.9900 ;
      RECT 11.1160 8.8965 11.1420 9.9900 ;
      RECT 11.0080 8.8965 11.0340 9.9900 ;
      RECT 10.9000 8.8965 10.9260 9.9900 ;
      RECT 10.7920 8.8965 10.8180 9.9900 ;
      RECT 10.6840 8.8965 10.7100 9.9900 ;
      RECT 10.5760 8.8965 10.6020 9.9900 ;
      RECT 10.4680 8.8965 10.4940 9.9900 ;
      RECT 10.3600 8.8965 10.3860 9.9900 ;
      RECT 10.2520 8.8965 10.2780 9.9900 ;
      RECT 10.1440 8.8965 10.1700 9.9900 ;
      RECT 10.0360 8.8965 10.0620 9.9900 ;
      RECT 9.9280 8.8965 9.9540 9.9900 ;
      RECT 9.8200 8.8965 9.8460 9.9900 ;
      RECT 9.7120 8.8965 9.7380 9.9900 ;
      RECT 9.6040 8.8965 9.6300 9.9900 ;
      RECT 9.4960 8.8965 9.5220 9.9900 ;
      RECT 9.3880 8.8965 9.4140 9.9900 ;
      RECT 9.2800 8.8965 9.3060 9.9900 ;
      RECT 9.1720 8.8965 9.1980 9.9900 ;
      RECT 9.0640 8.8965 9.0900 9.9900 ;
      RECT 8.9560 8.8965 8.9820 9.9900 ;
      RECT 8.8480 8.8965 8.8740 9.9900 ;
      RECT 8.7400 8.8965 8.7660 9.9900 ;
      RECT 8.6320 8.8965 8.6580 9.9900 ;
      RECT 8.5240 8.8965 8.5500 9.9900 ;
      RECT 8.4160 8.8965 8.4420 9.9900 ;
      RECT 8.3080 8.8965 8.3340 9.9900 ;
      RECT 8.2000 8.8965 8.2260 9.9900 ;
      RECT 8.0920 8.8965 8.1180 9.9900 ;
      RECT 7.9840 8.8965 8.0100 9.9900 ;
      RECT 7.8760 8.8965 7.9020 9.9900 ;
      RECT 7.7680 8.8965 7.7940 9.9900 ;
      RECT 7.6600 8.8965 7.6860 9.9900 ;
      RECT 7.5520 8.8965 7.5780 9.9900 ;
      RECT 7.4440 8.8965 7.4700 9.9900 ;
      RECT 7.3360 8.8965 7.3620 9.9900 ;
      RECT 7.2280 8.8965 7.2540 9.9900 ;
      RECT 7.1200 8.8965 7.1460 9.9900 ;
      RECT 7.0120 8.8965 7.0380 9.9900 ;
      RECT 6.9040 8.8965 6.9300 9.9900 ;
      RECT 6.7960 8.8965 6.8220 9.9900 ;
      RECT 6.6880 8.8965 6.7140 9.9900 ;
      RECT 6.5800 8.8965 6.6060 9.9900 ;
      RECT 6.4720 8.8965 6.4980 9.9900 ;
      RECT 6.3640 8.8965 6.3900 9.9900 ;
      RECT 6.2560 8.8965 6.2820 9.9900 ;
      RECT 6.1480 8.8965 6.1740 9.9900 ;
      RECT 6.0400 8.8965 6.0660 9.9900 ;
      RECT 5.9320 8.8965 5.9580 9.9900 ;
      RECT 5.8240 8.8965 5.8500 9.9900 ;
      RECT 5.7160 8.8965 5.7420 9.9900 ;
      RECT 5.6080 8.8965 5.6340 9.9900 ;
      RECT 5.5000 8.8965 5.5260 9.9900 ;
      RECT 5.3920 8.8965 5.4180 9.9900 ;
      RECT 5.2840 8.8965 5.3100 9.9900 ;
      RECT 5.1760 8.8965 5.2020 9.9900 ;
      RECT 5.0680 8.8965 5.0940 9.9900 ;
      RECT 4.9600 8.8965 4.9860 9.9900 ;
      RECT 4.8520 8.8965 4.8780 9.9900 ;
      RECT 4.7440 8.8965 4.7700 9.9900 ;
      RECT 4.6360 8.8965 4.6620 9.9900 ;
      RECT 4.5280 8.8965 4.5540 9.9900 ;
      RECT 4.4200 8.8965 4.4460 9.9900 ;
      RECT 4.3120 8.8965 4.3380 9.9900 ;
      RECT 4.2040 8.8965 4.2300 9.9900 ;
      RECT 4.0960 8.8965 4.1220 9.9900 ;
      RECT 3.9880 8.8965 4.0140 9.9900 ;
      RECT 3.8800 8.8965 3.9060 9.9900 ;
      RECT 3.7720 8.8965 3.7980 9.9900 ;
      RECT 3.6640 8.8965 3.6900 9.9900 ;
      RECT 3.5560 8.8965 3.5820 9.9900 ;
      RECT 3.4480 8.8965 3.4740 9.9900 ;
      RECT 3.3400 8.8965 3.3660 9.9900 ;
      RECT 3.2320 8.8965 3.2580 9.9900 ;
      RECT 3.1240 8.8965 3.1500 9.9900 ;
      RECT 3.0160 8.8965 3.0420 9.9900 ;
      RECT 2.9080 8.8965 2.9340 9.9900 ;
      RECT 2.8000 8.8965 2.8260 9.9900 ;
      RECT 2.6920 8.8965 2.7180 9.9900 ;
      RECT 2.5840 8.8965 2.6100 9.9900 ;
      RECT 2.4760 8.8965 2.5020 9.9900 ;
      RECT 2.3680 8.8965 2.3940 9.9900 ;
      RECT 2.2600 8.8965 2.2860 9.9900 ;
      RECT 2.1520 8.8965 2.1780 9.9900 ;
      RECT 2.0440 8.8965 2.0700 9.9900 ;
      RECT 1.9360 8.8965 1.9620 9.9900 ;
      RECT 1.8280 8.8965 1.8540 9.9900 ;
      RECT 1.7200 8.8965 1.7460 9.9900 ;
      RECT 1.6120 8.8965 1.6380 9.9900 ;
      RECT 1.5040 8.8965 1.5300 9.9900 ;
      RECT 1.3960 8.8965 1.4220 9.9900 ;
      RECT 1.2880 8.8965 1.3140 9.9900 ;
      RECT 1.1800 8.8965 1.2060 9.9900 ;
      RECT 1.0720 8.8965 1.0980 9.9900 ;
      RECT 0.9640 8.8965 0.9900 9.9900 ;
      RECT 0.8560 8.8965 0.8820 9.9900 ;
      RECT 0.7480 8.8965 0.7740 9.9900 ;
      RECT 0.6400 8.8965 0.6660 9.9900 ;
      RECT 0.5320 8.8965 0.5580 9.9900 ;
      RECT 0.4240 8.8965 0.4500 9.9900 ;
      RECT 0.3160 8.8965 0.3420 9.9900 ;
      RECT 0.2080 8.8965 0.2340 9.9900 ;
      RECT 0.0050 8.8965 0.0900 9.9900 ;
      RECT 15.5530 9.9765 15.6810 11.0700 ;
      RECT 15.5390 10.6420 15.6810 10.9645 ;
      RECT 15.3190 10.3690 15.4530 11.0700 ;
      RECT 15.2960 10.7040 15.4530 10.9620 ;
      RECT 15.3190 9.9765 15.4170 11.0700 ;
      RECT 15.3190 10.0975 15.4310 10.3370 ;
      RECT 15.3190 9.9765 15.4530 10.0655 ;
      RECT 15.0940 10.4270 15.2280 11.0700 ;
      RECT 15.0940 9.9765 15.1920 11.0700 ;
      RECT 14.6770 9.9765 14.7600 11.0700 ;
      RECT 14.6770 10.0650 14.7740 11.0005 ;
      RECT 30.2680 9.9765 30.3530 11.0700 ;
      RECT 30.1240 9.9765 30.1500 11.0700 ;
      RECT 30.0160 9.9765 30.0420 11.0700 ;
      RECT 29.9080 9.9765 29.9340 11.0700 ;
      RECT 29.8000 9.9765 29.8260 11.0700 ;
      RECT 29.6920 9.9765 29.7180 11.0700 ;
      RECT 29.5840 9.9765 29.6100 11.0700 ;
      RECT 29.4760 9.9765 29.5020 11.0700 ;
      RECT 29.3680 9.9765 29.3940 11.0700 ;
      RECT 29.2600 9.9765 29.2860 11.0700 ;
      RECT 29.1520 9.9765 29.1780 11.0700 ;
      RECT 29.0440 9.9765 29.0700 11.0700 ;
      RECT 28.9360 9.9765 28.9620 11.0700 ;
      RECT 28.8280 9.9765 28.8540 11.0700 ;
      RECT 28.7200 9.9765 28.7460 11.0700 ;
      RECT 28.6120 9.9765 28.6380 11.0700 ;
      RECT 28.5040 9.9765 28.5300 11.0700 ;
      RECT 28.3960 9.9765 28.4220 11.0700 ;
      RECT 28.2880 9.9765 28.3140 11.0700 ;
      RECT 28.1800 9.9765 28.2060 11.0700 ;
      RECT 28.0720 9.9765 28.0980 11.0700 ;
      RECT 27.9640 9.9765 27.9900 11.0700 ;
      RECT 27.8560 9.9765 27.8820 11.0700 ;
      RECT 27.7480 9.9765 27.7740 11.0700 ;
      RECT 27.6400 9.9765 27.6660 11.0700 ;
      RECT 27.5320 9.9765 27.5580 11.0700 ;
      RECT 27.4240 9.9765 27.4500 11.0700 ;
      RECT 27.3160 9.9765 27.3420 11.0700 ;
      RECT 27.2080 9.9765 27.2340 11.0700 ;
      RECT 27.1000 9.9765 27.1260 11.0700 ;
      RECT 26.9920 9.9765 27.0180 11.0700 ;
      RECT 26.8840 9.9765 26.9100 11.0700 ;
      RECT 26.7760 9.9765 26.8020 11.0700 ;
      RECT 26.6680 9.9765 26.6940 11.0700 ;
      RECT 26.5600 9.9765 26.5860 11.0700 ;
      RECT 26.4520 9.9765 26.4780 11.0700 ;
      RECT 26.3440 9.9765 26.3700 11.0700 ;
      RECT 26.2360 9.9765 26.2620 11.0700 ;
      RECT 26.1280 9.9765 26.1540 11.0700 ;
      RECT 26.0200 9.9765 26.0460 11.0700 ;
      RECT 25.9120 9.9765 25.9380 11.0700 ;
      RECT 25.8040 9.9765 25.8300 11.0700 ;
      RECT 25.6960 9.9765 25.7220 11.0700 ;
      RECT 25.5880 9.9765 25.6140 11.0700 ;
      RECT 25.4800 9.9765 25.5060 11.0700 ;
      RECT 25.3720 9.9765 25.3980 11.0700 ;
      RECT 25.2640 9.9765 25.2900 11.0700 ;
      RECT 25.1560 9.9765 25.1820 11.0700 ;
      RECT 25.0480 9.9765 25.0740 11.0700 ;
      RECT 24.9400 9.9765 24.9660 11.0700 ;
      RECT 24.8320 9.9765 24.8580 11.0700 ;
      RECT 24.7240 9.9765 24.7500 11.0700 ;
      RECT 24.6160 9.9765 24.6420 11.0700 ;
      RECT 24.5080 9.9765 24.5340 11.0700 ;
      RECT 24.4000 9.9765 24.4260 11.0700 ;
      RECT 24.2920 9.9765 24.3180 11.0700 ;
      RECT 24.1840 9.9765 24.2100 11.0700 ;
      RECT 24.0760 9.9765 24.1020 11.0700 ;
      RECT 23.9680 9.9765 23.9940 11.0700 ;
      RECT 23.8600 9.9765 23.8860 11.0700 ;
      RECT 23.7520 9.9765 23.7780 11.0700 ;
      RECT 23.6440 9.9765 23.6700 11.0700 ;
      RECT 23.5360 9.9765 23.5620 11.0700 ;
      RECT 23.4280 9.9765 23.4540 11.0700 ;
      RECT 23.3200 9.9765 23.3460 11.0700 ;
      RECT 23.2120 9.9765 23.2380 11.0700 ;
      RECT 23.1040 9.9765 23.1300 11.0700 ;
      RECT 22.9960 9.9765 23.0220 11.0700 ;
      RECT 22.8880 9.9765 22.9140 11.0700 ;
      RECT 22.7800 9.9765 22.8060 11.0700 ;
      RECT 22.6720 9.9765 22.6980 11.0700 ;
      RECT 22.5640 9.9765 22.5900 11.0700 ;
      RECT 22.4560 9.9765 22.4820 11.0700 ;
      RECT 22.3480 9.9765 22.3740 11.0700 ;
      RECT 22.2400 9.9765 22.2660 11.0700 ;
      RECT 22.1320 9.9765 22.1580 11.0700 ;
      RECT 22.0240 9.9765 22.0500 11.0700 ;
      RECT 21.9160 9.9765 21.9420 11.0700 ;
      RECT 21.8080 9.9765 21.8340 11.0700 ;
      RECT 21.7000 9.9765 21.7260 11.0700 ;
      RECT 21.5920 9.9765 21.6180 11.0700 ;
      RECT 21.4840 9.9765 21.5100 11.0700 ;
      RECT 21.3760 9.9765 21.4020 11.0700 ;
      RECT 21.2680 9.9765 21.2940 11.0700 ;
      RECT 21.1600 9.9765 21.1860 11.0700 ;
      RECT 21.0520 9.9765 21.0780 11.0700 ;
      RECT 20.9440 9.9765 20.9700 11.0700 ;
      RECT 20.8360 9.9765 20.8620 11.0700 ;
      RECT 20.7280 9.9765 20.7540 11.0700 ;
      RECT 20.6200 9.9765 20.6460 11.0700 ;
      RECT 20.5120 9.9765 20.5380 11.0700 ;
      RECT 20.4040 9.9765 20.4300 11.0700 ;
      RECT 20.2960 9.9765 20.3220 11.0700 ;
      RECT 20.1880 9.9765 20.2140 11.0700 ;
      RECT 20.0800 9.9765 20.1060 11.0700 ;
      RECT 19.9720 9.9765 19.9980 11.0700 ;
      RECT 19.8640 9.9765 19.8900 11.0700 ;
      RECT 19.7560 9.9765 19.7820 11.0700 ;
      RECT 19.6480 9.9765 19.6740 11.0700 ;
      RECT 19.5400 9.9765 19.5660 11.0700 ;
      RECT 19.4320 9.9765 19.4580 11.0700 ;
      RECT 19.3240 9.9765 19.3500 11.0700 ;
      RECT 19.2160 9.9765 19.2420 11.0700 ;
      RECT 19.1080 9.9765 19.1340 11.0700 ;
      RECT 19.0000 9.9765 19.0260 11.0700 ;
      RECT 18.8920 9.9765 18.9180 11.0700 ;
      RECT 18.7840 9.9765 18.8100 11.0700 ;
      RECT 18.6760 9.9765 18.7020 11.0700 ;
      RECT 18.5680 9.9765 18.5940 11.0700 ;
      RECT 18.4600 9.9765 18.4860 11.0700 ;
      RECT 18.3520 9.9765 18.3780 11.0700 ;
      RECT 18.2440 9.9765 18.2700 11.0700 ;
      RECT 18.1360 9.9765 18.1620 11.0700 ;
      RECT 18.0280 9.9765 18.0540 11.0700 ;
      RECT 17.9200 9.9765 17.9460 11.0700 ;
      RECT 17.8120 9.9765 17.8380 11.0700 ;
      RECT 17.7040 9.9765 17.7300 11.0700 ;
      RECT 17.5960 9.9765 17.6220 11.0700 ;
      RECT 17.4880 9.9765 17.5140 11.0700 ;
      RECT 17.3800 9.9765 17.4060 11.0700 ;
      RECT 17.2720 9.9765 17.2980 11.0700 ;
      RECT 17.1640 9.9765 17.1900 11.0700 ;
      RECT 17.0560 9.9765 17.0820 11.0700 ;
      RECT 16.9480 9.9765 16.9740 11.0700 ;
      RECT 16.8400 9.9765 16.8660 11.0700 ;
      RECT 16.7320 9.9765 16.7580 11.0700 ;
      RECT 16.6240 9.9765 16.6500 11.0700 ;
      RECT 16.5160 9.9765 16.5420 11.0700 ;
      RECT 16.4080 9.9765 16.4340 11.0700 ;
      RECT 16.3000 9.9765 16.3260 11.0700 ;
      RECT 16.0870 9.9765 16.1640 11.0700 ;
      RECT 14.1940 9.9765 14.2710 11.0700 ;
      RECT 14.0320 9.9765 14.0580 11.0700 ;
      RECT 13.9240 9.9765 13.9500 11.0700 ;
      RECT 13.8160 9.9765 13.8420 11.0700 ;
      RECT 13.7080 9.9765 13.7340 11.0700 ;
      RECT 13.6000 9.9765 13.6260 11.0700 ;
      RECT 13.4920 9.9765 13.5180 11.0700 ;
      RECT 13.3840 9.9765 13.4100 11.0700 ;
      RECT 13.2760 9.9765 13.3020 11.0700 ;
      RECT 13.1680 9.9765 13.1940 11.0700 ;
      RECT 13.0600 9.9765 13.0860 11.0700 ;
      RECT 12.9520 9.9765 12.9780 11.0700 ;
      RECT 12.8440 9.9765 12.8700 11.0700 ;
      RECT 12.7360 9.9765 12.7620 11.0700 ;
      RECT 12.6280 9.9765 12.6540 11.0700 ;
      RECT 12.5200 9.9765 12.5460 11.0700 ;
      RECT 12.4120 9.9765 12.4380 11.0700 ;
      RECT 12.3040 9.9765 12.3300 11.0700 ;
      RECT 12.1960 9.9765 12.2220 11.0700 ;
      RECT 12.0880 9.9765 12.1140 11.0700 ;
      RECT 11.9800 9.9765 12.0060 11.0700 ;
      RECT 11.8720 9.9765 11.8980 11.0700 ;
      RECT 11.7640 9.9765 11.7900 11.0700 ;
      RECT 11.6560 9.9765 11.6820 11.0700 ;
      RECT 11.5480 9.9765 11.5740 11.0700 ;
      RECT 11.4400 9.9765 11.4660 11.0700 ;
      RECT 11.3320 9.9765 11.3580 11.0700 ;
      RECT 11.2240 9.9765 11.2500 11.0700 ;
      RECT 11.1160 9.9765 11.1420 11.0700 ;
      RECT 11.0080 9.9765 11.0340 11.0700 ;
      RECT 10.9000 9.9765 10.9260 11.0700 ;
      RECT 10.7920 9.9765 10.8180 11.0700 ;
      RECT 10.6840 9.9765 10.7100 11.0700 ;
      RECT 10.5760 9.9765 10.6020 11.0700 ;
      RECT 10.4680 9.9765 10.4940 11.0700 ;
      RECT 10.3600 9.9765 10.3860 11.0700 ;
      RECT 10.2520 9.9765 10.2780 11.0700 ;
      RECT 10.1440 9.9765 10.1700 11.0700 ;
      RECT 10.0360 9.9765 10.0620 11.0700 ;
      RECT 9.9280 9.9765 9.9540 11.0700 ;
      RECT 9.8200 9.9765 9.8460 11.0700 ;
      RECT 9.7120 9.9765 9.7380 11.0700 ;
      RECT 9.6040 9.9765 9.6300 11.0700 ;
      RECT 9.4960 9.9765 9.5220 11.0700 ;
      RECT 9.3880 9.9765 9.4140 11.0700 ;
      RECT 9.2800 9.9765 9.3060 11.0700 ;
      RECT 9.1720 9.9765 9.1980 11.0700 ;
      RECT 9.0640 9.9765 9.0900 11.0700 ;
      RECT 8.9560 9.9765 8.9820 11.0700 ;
      RECT 8.8480 9.9765 8.8740 11.0700 ;
      RECT 8.7400 9.9765 8.7660 11.0700 ;
      RECT 8.6320 9.9765 8.6580 11.0700 ;
      RECT 8.5240 9.9765 8.5500 11.0700 ;
      RECT 8.4160 9.9765 8.4420 11.0700 ;
      RECT 8.3080 9.9765 8.3340 11.0700 ;
      RECT 8.2000 9.9765 8.2260 11.0700 ;
      RECT 8.0920 9.9765 8.1180 11.0700 ;
      RECT 7.9840 9.9765 8.0100 11.0700 ;
      RECT 7.8760 9.9765 7.9020 11.0700 ;
      RECT 7.7680 9.9765 7.7940 11.0700 ;
      RECT 7.6600 9.9765 7.6860 11.0700 ;
      RECT 7.5520 9.9765 7.5780 11.0700 ;
      RECT 7.4440 9.9765 7.4700 11.0700 ;
      RECT 7.3360 9.9765 7.3620 11.0700 ;
      RECT 7.2280 9.9765 7.2540 11.0700 ;
      RECT 7.1200 9.9765 7.1460 11.0700 ;
      RECT 7.0120 9.9765 7.0380 11.0700 ;
      RECT 6.9040 9.9765 6.9300 11.0700 ;
      RECT 6.7960 9.9765 6.8220 11.0700 ;
      RECT 6.6880 9.9765 6.7140 11.0700 ;
      RECT 6.5800 9.9765 6.6060 11.0700 ;
      RECT 6.4720 9.9765 6.4980 11.0700 ;
      RECT 6.3640 9.9765 6.3900 11.0700 ;
      RECT 6.2560 9.9765 6.2820 11.0700 ;
      RECT 6.1480 9.9765 6.1740 11.0700 ;
      RECT 6.0400 9.9765 6.0660 11.0700 ;
      RECT 5.9320 9.9765 5.9580 11.0700 ;
      RECT 5.8240 9.9765 5.8500 11.0700 ;
      RECT 5.7160 9.9765 5.7420 11.0700 ;
      RECT 5.6080 9.9765 5.6340 11.0700 ;
      RECT 5.5000 9.9765 5.5260 11.0700 ;
      RECT 5.3920 9.9765 5.4180 11.0700 ;
      RECT 5.2840 9.9765 5.3100 11.0700 ;
      RECT 5.1760 9.9765 5.2020 11.0700 ;
      RECT 5.0680 9.9765 5.0940 11.0700 ;
      RECT 4.9600 9.9765 4.9860 11.0700 ;
      RECT 4.8520 9.9765 4.8780 11.0700 ;
      RECT 4.7440 9.9765 4.7700 11.0700 ;
      RECT 4.6360 9.9765 4.6620 11.0700 ;
      RECT 4.5280 9.9765 4.5540 11.0700 ;
      RECT 4.4200 9.9765 4.4460 11.0700 ;
      RECT 4.3120 9.9765 4.3380 11.0700 ;
      RECT 4.2040 9.9765 4.2300 11.0700 ;
      RECT 4.0960 9.9765 4.1220 11.0700 ;
      RECT 3.9880 9.9765 4.0140 11.0700 ;
      RECT 3.8800 9.9765 3.9060 11.0700 ;
      RECT 3.7720 9.9765 3.7980 11.0700 ;
      RECT 3.6640 9.9765 3.6900 11.0700 ;
      RECT 3.5560 9.9765 3.5820 11.0700 ;
      RECT 3.4480 9.9765 3.4740 11.0700 ;
      RECT 3.3400 9.9765 3.3660 11.0700 ;
      RECT 3.2320 9.9765 3.2580 11.0700 ;
      RECT 3.1240 9.9765 3.1500 11.0700 ;
      RECT 3.0160 9.9765 3.0420 11.0700 ;
      RECT 2.9080 9.9765 2.9340 11.0700 ;
      RECT 2.8000 9.9765 2.8260 11.0700 ;
      RECT 2.6920 9.9765 2.7180 11.0700 ;
      RECT 2.5840 9.9765 2.6100 11.0700 ;
      RECT 2.4760 9.9765 2.5020 11.0700 ;
      RECT 2.3680 9.9765 2.3940 11.0700 ;
      RECT 2.2600 9.9765 2.2860 11.0700 ;
      RECT 2.1520 9.9765 2.1780 11.0700 ;
      RECT 2.0440 9.9765 2.0700 11.0700 ;
      RECT 1.9360 9.9765 1.9620 11.0700 ;
      RECT 1.8280 9.9765 1.8540 11.0700 ;
      RECT 1.7200 9.9765 1.7460 11.0700 ;
      RECT 1.6120 9.9765 1.6380 11.0700 ;
      RECT 1.5040 9.9765 1.5300 11.0700 ;
      RECT 1.3960 9.9765 1.4220 11.0700 ;
      RECT 1.2880 9.9765 1.3140 11.0700 ;
      RECT 1.1800 9.9765 1.2060 11.0700 ;
      RECT 1.0720 9.9765 1.0980 11.0700 ;
      RECT 0.9640 9.9765 0.9900 11.0700 ;
      RECT 0.8560 9.9765 0.8820 11.0700 ;
      RECT 0.7480 9.9765 0.7740 11.0700 ;
      RECT 0.6400 9.9765 0.6660 11.0700 ;
      RECT 0.5320 9.9765 0.5580 11.0700 ;
      RECT 0.4240 9.9765 0.4500 11.0700 ;
      RECT 0.3160 9.9765 0.3420 11.0700 ;
      RECT 0.2080 9.9765 0.2340 11.0700 ;
      RECT 0.0050 9.9765 0.0900 11.0700 ;
      RECT 14.1350 19.3060 30.3480 19.7470 ;
      RECT 17.7530 11.0935 30.3480 19.7470 ;
      RECT 16.2950 12.5975 30.3480 19.7470 ;
      RECT 17.5370 12.4025 30.3480 19.7470 ;
      RECT 14.1350 19.0055 16.2130 19.7470 ;
      RECT 15.5570 12.4985 16.2130 19.7470 ;
      RECT 14.1350 12.7055 15.2590 19.7470 ;
      RECT 15.1970 11.0935 15.2590 19.7470 ;
      RECT 15.5430 17.7395 16.2130 18.8475 ;
      RECT 16.2810 14.8865 30.3480 18.4795 ;
      RECT 14.1350 17.9735 15.2730 18.2355 ;
      RECT 15.5430 15.2015 16.2130 17.5335 ;
      RECT 14.1350 15.5795 15.2730 16.8855 ;
      RECT 14.1350 12.9155 15.2730 15.5355 ;
      RECT 15.5430 12.3755 16.1590 14.1615 ;
      RECT 14.1890 12.6455 15.2730 12.8355 ;
      RECT 14.1890 11.8595 15.2590 19.7470 ;
      RECT 14.4050 11.7785 15.2590 19.7470 ;
      RECT 14.1890 12.3755 15.2730 12.6015 ;
      RECT 16.4570 12.4055 30.3480 19.7470 ;
      RECT 16.2950 11.0935 16.3750 19.7470 ;
      RECT 14.1350 11.7785 14.3230 12.5925 ;
      RECT 16.2950 11.0935 16.5910 12.4965 ;
      RECT 16.2950 12.2105 17.4550 12.4965 ;
      RECT 17.5370 11.0935 17.6710 19.7470 ;
      RECT 15.5570 12.2105 16.1590 19.7470 ;
      RECT 15.8810 11.0935 16.2130 12.3435 ;
      RECT 16.2950 12.2105 17.6710 12.3045 ;
      RECT 17.3210 11.0935 30.3480 12.3015 ;
      RECT 14.1350 12.2315 15.2730 12.2955 ;
      RECT 17.1050 11.8265 30.3480 12.3015 ;
      RECT 16.2950 11.8595 17.0230 12.4965 ;
      RECT 15.5570 11.8595 15.7990 19.7470 ;
      RECT 14.4050 11.8355 15.2730 12.0975 ;
      RECT 15.5930 11.0935 16.2130 12.0015 ;
      RECT 16.8890 11.0935 17.2390 11.9655 ;
      RECT 16.2950 11.7785 16.8070 12.4965 ;
      RECT 16.6730 11.0935 16.8070 19.7470 ;
      RECT 14.4050 11.0935 15.1150 19.7470 ;
      RECT 14.2250 11.0935 14.3230 19.7470 ;
      RECT 16.6730 11.0935 17.2390 11.7285 ;
      RECT 15.5570 11.0935 16.2130 11.7285 ;
      RECT 14.2250 11.0935 15.1150 11.7285 ;
      RECT 16.6730 11.0935 30.3480 11.7255 ;
      RECT 15.5430 11.5655 16.2130 11.7195 ;
      RECT 16.2950 11.0935 30.3480 11.4615 ;
      RECT 14.1350 11.0935 15.2590 11.4615 ;
      RECT 14.1350 11.0935 16.2130 11.2585 ;
      RECT 17.7570 10.9035 17.7750 19.7470 ;
      RECT 17.6490 10.9035 17.6670 19.7470 ;
      RECT 17.5410 10.9035 17.5590 19.7470 ;
      RECT 17.4330 10.9035 17.4510 19.7470 ;
      RECT 17.3250 10.9035 17.3430 19.7470 ;
      RECT 17.2170 10.9035 17.2350 19.7470 ;
      RECT 17.1090 10.9035 17.1270 19.7470 ;
      RECT 17.0010 10.9035 17.0190 19.7470 ;
      RECT 16.8930 10.9035 16.9110 19.7470 ;
      RECT 16.7850 10.9035 16.8030 19.7470 ;
      RECT 16.6770 10.9035 16.6950 19.7470 ;
      RECT 16.5690 10.9035 16.5870 19.7470 ;
      RECT 16.4610 10.9035 16.4790 19.7470 ;
      RECT 16.3530 10.9035 16.3710 19.7470 ;
      RECT 0.0000 12.4025 14.0170 19.7470 ;
      RECT 0.0000 15.1915 14.0310 15.2745 ;
      RECT 13.7570 11.0935 14.0530 14.8530 ;
      RECT 12.8930 12.0215 13.6750 19.7470 ;
      RECT 0.0000 11.0935 12.8110 19.7470 ;
      RECT 13.5410 11.0935 14.0530 12.3015 ;
      RECT 0.0000 11.8265 13.4590 12.3015 ;
      RECT 13.3250 11.0935 13.4590 19.7470 ;
      RECT 13.1090 11.7785 13.4590 19.7470 ;
      RECT 0.0000 11.0935 13.0270 12.3015 ;
      RECT 13.1090 11.0935 13.2430 19.7470 ;
      RECT 13.3250 11.0935 14.0530 11.7285 ;
      RECT 0.0000 11.0935 13.2430 11.7255 ;
      RECT 0.0000 11.0935 14.0530 11.4615 ;
      RECT 13.3290 11.0670 13.3470 19.7470 ;
      RECT 13.2210 11.0670 13.2390 19.7470 ;
        RECT 15.5530 19.1835 15.6810 20.2770 ;
        RECT 15.5390 19.8490 15.6810 20.1715 ;
        RECT 15.3190 19.5760 15.4530 20.2770 ;
        RECT 15.2960 19.9110 15.4530 20.1690 ;
        RECT 15.3190 19.1835 15.4170 20.2770 ;
        RECT 15.3190 19.3045 15.4310 19.5440 ;
        RECT 15.3190 19.1835 15.4530 19.2725 ;
        RECT 15.0940 19.6340 15.2280 20.2770 ;
        RECT 15.0940 19.1835 15.1920 20.2770 ;
        RECT 14.6770 19.1835 14.7600 20.2770 ;
        RECT 14.6770 19.2720 14.7740 20.2075 ;
        RECT 30.2680 19.1835 30.3530 20.2770 ;
        RECT 30.1240 19.1835 30.1500 20.2770 ;
        RECT 30.0160 19.1835 30.0420 20.2770 ;
        RECT 29.9080 19.1835 29.9340 20.2770 ;
        RECT 29.8000 19.1835 29.8260 20.2770 ;
        RECT 29.6920 19.1835 29.7180 20.2770 ;
        RECT 29.5840 19.1835 29.6100 20.2770 ;
        RECT 29.4760 19.1835 29.5020 20.2770 ;
        RECT 29.3680 19.1835 29.3940 20.2770 ;
        RECT 29.2600 19.1835 29.2860 20.2770 ;
        RECT 29.1520 19.1835 29.1780 20.2770 ;
        RECT 29.0440 19.1835 29.0700 20.2770 ;
        RECT 28.9360 19.1835 28.9620 20.2770 ;
        RECT 28.8280 19.1835 28.8540 20.2770 ;
        RECT 28.7200 19.1835 28.7460 20.2770 ;
        RECT 28.6120 19.1835 28.6380 20.2770 ;
        RECT 28.5040 19.1835 28.5300 20.2770 ;
        RECT 28.3960 19.1835 28.4220 20.2770 ;
        RECT 28.2880 19.1835 28.3140 20.2770 ;
        RECT 28.1800 19.1835 28.2060 20.2770 ;
        RECT 28.0720 19.1835 28.0980 20.2770 ;
        RECT 27.9640 19.1835 27.9900 20.2770 ;
        RECT 27.8560 19.1835 27.8820 20.2770 ;
        RECT 27.7480 19.1835 27.7740 20.2770 ;
        RECT 27.6400 19.1835 27.6660 20.2770 ;
        RECT 27.5320 19.1835 27.5580 20.2770 ;
        RECT 27.4240 19.1835 27.4500 20.2770 ;
        RECT 27.3160 19.1835 27.3420 20.2770 ;
        RECT 27.2080 19.1835 27.2340 20.2770 ;
        RECT 27.1000 19.1835 27.1260 20.2770 ;
        RECT 26.9920 19.1835 27.0180 20.2770 ;
        RECT 26.8840 19.1835 26.9100 20.2770 ;
        RECT 26.7760 19.1835 26.8020 20.2770 ;
        RECT 26.6680 19.1835 26.6940 20.2770 ;
        RECT 26.5600 19.1835 26.5860 20.2770 ;
        RECT 26.4520 19.1835 26.4780 20.2770 ;
        RECT 26.3440 19.1835 26.3700 20.2770 ;
        RECT 26.2360 19.1835 26.2620 20.2770 ;
        RECT 26.1280 19.1835 26.1540 20.2770 ;
        RECT 26.0200 19.1835 26.0460 20.2770 ;
        RECT 25.9120 19.1835 25.9380 20.2770 ;
        RECT 25.8040 19.1835 25.8300 20.2770 ;
        RECT 25.6960 19.1835 25.7220 20.2770 ;
        RECT 25.5880 19.1835 25.6140 20.2770 ;
        RECT 25.4800 19.1835 25.5060 20.2770 ;
        RECT 25.3720 19.1835 25.3980 20.2770 ;
        RECT 25.2640 19.1835 25.2900 20.2770 ;
        RECT 25.1560 19.1835 25.1820 20.2770 ;
        RECT 25.0480 19.1835 25.0740 20.2770 ;
        RECT 24.9400 19.1835 24.9660 20.2770 ;
        RECT 24.8320 19.1835 24.8580 20.2770 ;
        RECT 24.7240 19.1835 24.7500 20.2770 ;
        RECT 24.6160 19.1835 24.6420 20.2770 ;
        RECT 24.5080 19.1835 24.5340 20.2770 ;
        RECT 24.4000 19.1835 24.4260 20.2770 ;
        RECT 24.2920 19.1835 24.3180 20.2770 ;
        RECT 24.1840 19.1835 24.2100 20.2770 ;
        RECT 24.0760 19.1835 24.1020 20.2770 ;
        RECT 23.9680 19.1835 23.9940 20.2770 ;
        RECT 23.8600 19.1835 23.8860 20.2770 ;
        RECT 23.7520 19.1835 23.7780 20.2770 ;
        RECT 23.6440 19.1835 23.6700 20.2770 ;
        RECT 23.5360 19.1835 23.5620 20.2770 ;
        RECT 23.4280 19.1835 23.4540 20.2770 ;
        RECT 23.3200 19.1835 23.3460 20.2770 ;
        RECT 23.2120 19.1835 23.2380 20.2770 ;
        RECT 23.1040 19.1835 23.1300 20.2770 ;
        RECT 22.9960 19.1835 23.0220 20.2770 ;
        RECT 22.8880 19.1835 22.9140 20.2770 ;
        RECT 22.7800 19.1835 22.8060 20.2770 ;
        RECT 22.6720 19.1835 22.6980 20.2770 ;
        RECT 22.5640 19.1835 22.5900 20.2770 ;
        RECT 22.4560 19.1835 22.4820 20.2770 ;
        RECT 22.3480 19.1835 22.3740 20.2770 ;
        RECT 22.2400 19.1835 22.2660 20.2770 ;
        RECT 22.1320 19.1835 22.1580 20.2770 ;
        RECT 22.0240 19.1835 22.0500 20.2770 ;
        RECT 21.9160 19.1835 21.9420 20.2770 ;
        RECT 21.8080 19.1835 21.8340 20.2770 ;
        RECT 21.7000 19.1835 21.7260 20.2770 ;
        RECT 21.5920 19.1835 21.6180 20.2770 ;
        RECT 21.4840 19.1835 21.5100 20.2770 ;
        RECT 21.3760 19.1835 21.4020 20.2770 ;
        RECT 21.2680 19.1835 21.2940 20.2770 ;
        RECT 21.1600 19.1835 21.1860 20.2770 ;
        RECT 21.0520 19.1835 21.0780 20.2770 ;
        RECT 20.9440 19.1835 20.9700 20.2770 ;
        RECT 20.8360 19.1835 20.8620 20.2770 ;
        RECT 20.7280 19.1835 20.7540 20.2770 ;
        RECT 20.6200 19.1835 20.6460 20.2770 ;
        RECT 20.5120 19.1835 20.5380 20.2770 ;
        RECT 20.4040 19.1835 20.4300 20.2770 ;
        RECT 20.2960 19.1835 20.3220 20.2770 ;
        RECT 20.1880 19.1835 20.2140 20.2770 ;
        RECT 20.0800 19.1835 20.1060 20.2770 ;
        RECT 19.9720 19.1835 19.9980 20.2770 ;
        RECT 19.8640 19.1835 19.8900 20.2770 ;
        RECT 19.7560 19.1835 19.7820 20.2770 ;
        RECT 19.6480 19.1835 19.6740 20.2770 ;
        RECT 19.5400 19.1835 19.5660 20.2770 ;
        RECT 19.4320 19.1835 19.4580 20.2770 ;
        RECT 19.3240 19.1835 19.3500 20.2770 ;
        RECT 19.2160 19.1835 19.2420 20.2770 ;
        RECT 19.1080 19.1835 19.1340 20.2770 ;
        RECT 19.0000 19.1835 19.0260 20.2770 ;
        RECT 18.8920 19.1835 18.9180 20.2770 ;
        RECT 18.7840 19.1835 18.8100 20.2770 ;
        RECT 18.6760 19.1835 18.7020 20.2770 ;
        RECT 18.5680 19.1835 18.5940 20.2770 ;
        RECT 18.4600 19.1835 18.4860 20.2770 ;
        RECT 18.3520 19.1835 18.3780 20.2770 ;
        RECT 18.2440 19.1835 18.2700 20.2770 ;
        RECT 18.1360 19.1835 18.1620 20.2770 ;
        RECT 18.0280 19.1835 18.0540 20.2770 ;
        RECT 17.9200 19.1835 17.9460 20.2770 ;
        RECT 17.8120 19.1835 17.8380 20.2770 ;
        RECT 17.7040 19.1835 17.7300 20.2770 ;
        RECT 17.5960 19.1835 17.6220 20.2770 ;
        RECT 17.4880 19.1835 17.5140 20.2770 ;
        RECT 17.3800 19.1835 17.4060 20.2770 ;
        RECT 17.2720 19.1835 17.2980 20.2770 ;
        RECT 17.1640 19.1835 17.1900 20.2770 ;
        RECT 17.0560 19.1835 17.0820 20.2770 ;
        RECT 16.9480 19.1835 16.9740 20.2770 ;
        RECT 16.8400 19.1835 16.8660 20.2770 ;
        RECT 16.7320 19.1835 16.7580 20.2770 ;
        RECT 16.6240 19.1835 16.6500 20.2770 ;
        RECT 16.5160 19.1835 16.5420 20.2770 ;
        RECT 16.4080 19.1835 16.4340 20.2770 ;
        RECT 16.3000 19.1835 16.3260 20.2770 ;
        RECT 16.0870 19.1835 16.1640 20.2770 ;
        RECT 14.1940 19.1835 14.2710 20.2770 ;
        RECT 14.0320 19.1835 14.0580 20.2770 ;
        RECT 13.9240 19.1835 13.9500 20.2770 ;
        RECT 13.8160 19.1835 13.8420 20.2770 ;
        RECT 13.7080 19.1835 13.7340 20.2770 ;
        RECT 13.6000 19.1835 13.6260 20.2770 ;
        RECT 13.4920 19.1835 13.5180 20.2770 ;
        RECT 13.3840 19.1835 13.4100 20.2770 ;
        RECT 13.2760 19.1835 13.3020 20.2770 ;
        RECT 13.1680 19.1835 13.1940 20.2770 ;
        RECT 13.0600 19.1835 13.0860 20.2770 ;
        RECT 12.9520 19.1835 12.9780 20.2770 ;
        RECT 12.8440 19.1835 12.8700 20.2770 ;
        RECT 12.7360 19.1835 12.7620 20.2770 ;
        RECT 12.6280 19.1835 12.6540 20.2770 ;
        RECT 12.5200 19.1835 12.5460 20.2770 ;
        RECT 12.4120 19.1835 12.4380 20.2770 ;
        RECT 12.3040 19.1835 12.3300 20.2770 ;
        RECT 12.1960 19.1835 12.2220 20.2770 ;
        RECT 12.0880 19.1835 12.1140 20.2770 ;
        RECT 11.9800 19.1835 12.0060 20.2770 ;
        RECT 11.8720 19.1835 11.8980 20.2770 ;
        RECT 11.7640 19.1835 11.7900 20.2770 ;
        RECT 11.6560 19.1835 11.6820 20.2770 ;
        RECT 11.5480 19.1835 11.5740 20.2770 ;
        RECT 11.4400 19.1835 11.4660 20.2770 ;
        RECT 11.3320 19.1835 11.3580 20.2770 ;
        RECT 11.2240 19.1835 11.2500 20.2770 ;
        RECT 11.1160 19.1835 11.1420 20.2770 ;
        RECT 11.0080 19.1835 11.0340 20.2770 ;
        RECT 10.9000 19.1835 10.9260 20.2770 ;
        RECT 10.7920 19.1835 10.8180 20.2770 ;
        RECT 10.6840 19.1835 10.7100 20.2770 ;
        RECT 10.5760 19.1835 10.6020 20.2770 ;
        RECT 10.4680 19.1835 10.4940 20.2770 ;
        RECT 10.3600 19.1835 10.3860 20.2770 ;
        RECT 10.2520 19.1835 10.2780 20.2770 ;
        RECT 10.1440 19.1835 10.1700 20.2770 ;
        RECT 10.0360 19.1835 10.0620 20.2770 ;
        RECT 9.9280 19.1835 9.9540 20.2770 ;
        RECT 9.8200 19.1835 9.8460 20.2770 ;
        RECT 9.7120 19.1835 9.7380 20.2770 ;
        RECT 9.6040 19.1835 9.6300 20.2770 ;
        RECT 9.4960 19.1835 9.5220 20.2770 ;
        RECT 9.3880 19.1835 9.4140 20.2770 ;
        RECT 9.2800 19.1835 9.3060 20.2770 ;
        RECT 9.1720 19.1835 9.1980 20.2770 ;
        RECT 9.0640 19.1835 9.0900 20.2770 ;
        RECT 8.9560 19.1835 8.9820 20.2770 ;
        RECT 8.8480 19.1835 8.8740 20.2770 ;
        RECT 8.7400 19.1835 8.7660 20.2770 ;
        RECT 8.6320 19.1835 8.6580 20.2770 ;
        RECT 8.5240 19.1835 8.5500 20.2770 ;
        RECT 8.4160 19.1835 8.4420 20.2770 ;
        RECT 8.3080 19.1835 8.3340 20.2770 ;
        RECT 8.2000 19.1835 8.2260 20.2770 ;
        RECT 8.0920 19.1835 8.1180 20.2770 ;
        RECT 7.9840 19.1835 8.0100 20.2770 ;
        RECT 7.8760 19.1835 7.9020 20.2770 ;
        RECT 7.7680 19.1835 7.7940 20.2770 ;
        RECT 7.6600 19.1835 7.6860 20.2770 ;
        RECT 7.5520 19.1835 7.5780 20.2770 ;
        RECT 7.4440 19.1835 7.4700 20.2770 ;
        RECT 7.3360 19.1835 7.3620 20.2770 ;
        RECT 7.2280 19.1835 7.2540 20.2770 ;
        RECT 7.1200 19.1835 7.1460 20.2770 ;
        RECT 7.0120 19.1835 7.0380 20.2770 ;
        RECT 6.9040 19.1835 6.9300 20.2770 ;
        RECT 6.7960 19.1835 6.8220 20.2770 ;
        RECT 6.6880 19.1835 6.7140 20.2770 ;
        RECT 6.5800 19.1835 6.6060 20.2770 ;
        RECT 6.4720 19.1835 6.4980 20.2770 ;
        RECT 6.3640 19.1835 6.3900 20.2770 ;
        RECT 6.2560 19.1835 6.2820 20.2770 ;
        RECT 6.1480 19.1835 6.1740 20.2770 ;
        RECT 6.0400 19.1835 6.0660 20.2770 ;
        RECT 5.9320 19.1835 5.9580 20.2770 ;
        RECT 5.8240 19.1835 5.8500 20.2770 ;
        RECT 5.7160 19.1835 5.7420 20.2770 ;
        RECT 5.6080 19.1835 5.6340 20.2770 ;
        RECT 5.5000 19.1835 5.5260 20.2770 ;
        RECT 5.3920 19.1835 5.4180 20.2770 ;
        RECT 5.2840 19.1835 5.3100 20.2770 ;
        RECT 5.1760 19.1835 5.2020 20.2770 ;
        RECT 5.0680 19.1835 5.0940 20.2770 ;
        RECT 4.9600 19.1835 4.9860 20.2770 ;
        RECT 4.8520 19.1835 4.8780 20.2770 ;
        RECT 4.7440 19.1835 4.7700 20.2770 ;
        RECT 4.6360 19.1835 4.6620 20.2770 ;
        RECT 4.5280 19.1835 4.5540 20.2770 ;
        RECT 4.4200 19.1835 4.4460 20.2770 ;
        RECT 4.3120 19.1835 4.3380 20.2770 ;
        RECT 4.2040 19.1835 4.2300 20.2770 ;
        RECT 4.0960 19.1835 4.1220 20.2770 ;
        RECT 3.9880 19.1835 4.0140 20.2770 ;
        RECT 3.8800 19.1835 3.9060 20.2770 ;
        RECT 3.7720 19.1835 3.7980 20.2770 ;
        RECT 3.6640 19.1835 3.6900 20.2770 ;
        RECT 3.5560 19.1835 3.5820 20.2770 ;
        RECT 3.4480 19.1835 3.4740 20.2770 ;
        RECT 3.3400 19.1835 3.3660 20.2770 ;
        RECT 3.2320 19.1835 3.2580 20.2770 ;
        RECT 3.1240 19.1835 3.1500 20.2770 ;
        RECT 3.0160 19.1835 3.0420 20.2770 ;
        RECT 2.9080 19.1835 2.9340 20.2770 ;
        RECT 2.8000 19.1835 2.8260 20.2770 ;
        RECT 2.6920 19.1835 2.7180 20.2770 ;
        RECT 2.5840 19.1835 2.6100 20.2770 ;
        RECT 2.4760 19.1835 2.5020 20.2770 ;
        RECT 2.3680 19.1835 2.3940 20.2770 ;
        RECT 2.2600 19.1835 2.2860 20.2770 ;
        RECT 2.1520 19.1835 2.1780 20.2770 ;
        RECT 2.0440 19.1835 2.0700 20.2770 ;
        RECT 1.9360 19.1835 1.9620 20.2770 ;
        RECT 1.8280 19.1835 1.8540 20.2770 ;
        RECT 1.7200 19.1835 1.7460 20.2770 ;
        RECT 1.6120 19.1835 1.6380 20.2770 ;
        RECT 1.5040 19.1835 1.5300 20.2770 ;
        RECT 1.3960 19.1835 1.4220 20.2770 ;
        RECT 1.2880 19.1835 1.3140 20.2770 ;
        RECT 1.1800 19.1835 1.2060 20.2770 ;
        RECT 1.0720 19.1835 1.0980 20.2770 ;
        RECT 0.9640 19.1835 0.9900 20.2770 ;
        RECT 0.8560 19.1835 0.8820 20.2770 ;
        RECT 0.7480 19.1835 0.7740 20.2770 ;
        RECT 0.6400 19.1835 0.6660 20.2770 ;
        RECT 0.5320 19.1835 0.5580 20.2770 ;
        RECT 0.4240 19.1835 0.4500 20.2770 ;
        RECT 0.3160 19.1835 0.3420 20.2770 ;
        RECT 0.2080 19.1835 0.2340 20.2770 ;
        RECT 0.0050 19.1835 0.0900 20.2770 ;
        RECT 15.5530 20.2635 15.6810 21.3570 ;
        RECT 15.5390 20.9290 15.6810 21.2515 ;
        RECT 15.3190 20.6560 15.4530 21.3570 ;
        RECT 15.2960 20.9910 15.4530 21.2490 ;
        RECT 15.3190 20.2635 15.4170 21.3570 ;
        RECT 15.3190 20.3845 15.4310 20.6240 ;
        RECT 15.3190 20.2635 15.4530 20.3525 ;
        RECT 15.0940 20.7140 15.2280 21.3570 ;
        RECT 15.0940 20.2635 15.1920 21.3570 ;
        RECT 14.6770 20.2635 14.7600 21.3570 ;
        RECT 14.6770 20.3520 14.7740 21.2875 ;
        RECT 30.2680 20.2635 30.3530 21.3570 ;
        RECT 30.1240 20.2635 30.1500 21.3570 ;
        RECT 30.0160 20.2635 30.0420 21.3570 ;
        RECT 29.9080 20.2635 29.9340 21.3570 ;
        RECT 29.8000 20.2635 29.8260 21.3570 ;
        RECT 29.6920 20.2635 29.7180 21.3570 ;
        RECT 29.5840 20.2635 29.6100 21.3570 ;
        RECT 29.4760 20.2635 29.5020 21.3570 ;
        RECT 29.3680 20.2635 29.3940 21.3570 ;
        RECT 29.2600 20.2635 29.2860 21.3570 ;
        RECT 29.1520 20.2635 29.1780 21.3570 ;
        RECT 29.0440 20.2635 29.0700 21.3570 ;
        RECT 28.9360 20.2635 28.9620 21.3570 ;
        RECT 28.8280 20.2635 28.8540 21.3570 ;
        RECT 28.7200 20.2635 28.7460 21.3570 ;
        RECT 28.6120 20.2635 28.6380 21.3570 ;
        RECT 28.5040 20.2635 28.5300 21.3570 ;
        RECT 28.3960 20.2635 28.4220 21.3570 ;
        RECT 28.2880 20.2635 28.3140 21.3570 ;
        RECT 28.1800 20.2635 28.2060 21.3570 ;
        RECT 28.0720 20.2635 28.0980 21.3570 ;
        RECT 27.9640 20.2635 27.9900 21.3570 ;
        RECT 27.8560 20.2635 27.8820 21.3570 ;
        RECT 27.7480 20.2635 27.7740 21.3570 ;
        RECT 27.6400 20.2635 27.6660 21.3570 ;
        RECT 27.5320 20.2635 27.5580 21.3570 ;
        RECT 27.4240 20.2635 27.4500 21.3570 ;
        RECT 27.3160 20.2635 27.3420 21.3570 ;
        RECT 27.2080 20.2635 27.2340 21.3570 ;
        RECT 27.1000 20.2635 27.1260 21.3570 ;
        RECT 26.9920 20.2635 27.0180 21.3570 ;
        RECT 26.8840 20.2635 26.9100 21.3570 ;
        RECT 26.7760 20.2635 26.8020 21.3570 ;
        RECT 26.6680 20.2635 26.6940 21.3570 ;
        RECT 26.5600 20.2635 26.5860 21.3570 ;
        RECT 26.4520 20.2635 26.4780 21.3570 ;
        RECT 26.3440 20.2635 26.3700 21.3570 ;
        RECT 26.2360 20.2635 26.2620 21.3570 ;
        RECT 26.1280 20.2635 26.1540 21.3570 ;
        RECT 26.0200 20.2635 26.0460 21.3570 ;
        RECT 25.9120 20.2635 25.9380 21.3570 ;
        RECT 25.8040 20.2635 25.8300 21.3570 ;
        RECT 25.6960 20.2635 25.7220 21.3570 ;
        RECT 25.5880 20.2635 25.6140 21.3570 ;
        RECT 25.4800 20.2635 25.5060 21.3570 ;
        RECT 25.3720 20.2635 25.3980 21.3570 ;
        RECT 25.2640 20.2635 25.2900 21.3570 ;
        RECT 25.1560 20.2635 25.1820 21.3570 ;
        RECT 25.0480 20.2635 25.0740 21.3570 ;
        RECT 24.9400 20.2635 24.9660 21.3570 ;
        RECT 24.8320 20.2635 24.8580 21.3570 ;
        RECT 24.7240 20.2635 24.7500 21.3570 ;
        RECT 24.6160 20.2635 24.6420 21.3570 ;
        RECT 24.5080 20.2635 24.5340 21.3570 ;
        RECT 24.4000 20.2635 24.4260 21.3570 ;
        RECT 24.2920 20.2635 24.3180 21.3570 ;
        RECT 24.1840 20.2635 24.2100 21.3570 ;
        RECT 24.0760 20.2635 24.1020 21.3570 ;
        RECT 23.9680 20.2635 23.9940 21.3570 ;
        RECT 23.8600 20.2635 23.8860 21.3570 ;
        RECT 23.7520 20.2635 23.7780 21.3570 ;
        RECT 23.6440 20.2635 23.6700 21.3570 ;
        RECT 23.5360 20.2635 23.5620 21.3570 ;
        RECT 23.4280 20.2635 23.4540 21.3570 ;
        RECT 23.3200 20.2635 23.3460 21.3570 ;
        RECT 23.2120 20.2635 23.2380 21.3570 ;
        RECT 23.1040 20.2635 23.1300 21.3570 ;
        RECT 22.9960 20.2635 23.0220 21.3570 ;
        RECT 22.8880 20.2635 22.9140 21.3570 ;
        RECT 22.7800 20.2635 22.8060 21.3570 ;
        RECT 22.6720 20.2635 22.6980 21.3570 ;
        RECT 22.5640 20.2635 22.5900 21.3570 ;
        RECT 22.4560 20.2635 22.4820 21.3570 ;
        RECT 22.3480 20.2635 22.3740 21.3570 ;
        RECT 22.2400 20.2635 22.2660 21.3570 ;
        RECT 22.1320 20.2635 22.1580 21.3570 ;
        RECT 22.0240 20.2635 22.0500 21.3570 ;
        RECT 21.9160 20.2635 21.9420 21.3570 ;
        RECT 21.8080 20.2635 21.8340 21.3570 ;
        RECT 21.7000 20.2635 21.7260 21.3570 ;
        RECT 21.5920 20.2635 21.6180 21.3570 ;
        RECT 21.4840 20.2635 21.5100 21.3570 ;
        RECT 21.3760 20.2635 21.4020 21.3570 ;
        RECT 21.2680 20.2635 21.2940 21.3570 ;
        RECT 21.1600 20.2635 21.1860 21.3570 ;
        RECT 21.0520 20.2635 21.0780 21.3570 ;
        RECT 20.9440 20.2635 20.9700 21.3570 ;
        RECT 20.8360 20.2635 20.8620 21.3570 ;
        RECT 20.7280 20.2635 20.7540 21.3570 ;
        RECT 20.6200 20.2635 20.6460 21.3570 ;
        RECT 20.5120 20.2635 20.5380 21.3570 ;
        RECT 20.4040 20.2635 20.4300 21.3570 ;
        RECT 20.2960 20.2635 20.3220 21.3570 ;
        RECT 20.1880 20.2635 20.2140 21.3570 ;
        RECT 20.0800 20.2635 20.1060 21.3570 ;
        RECT 19.9720 20.2635 19.9980 21.3570 ;
        RECT 19.8640 20.2635 19.8900 21.3570 ;
        RECT 19.7560 20.2635 19.7820 21.3570 ;
        RECT 19.6480 20.2635 19.6740 21.3570 ;
        RECT 19.5400 20.2635 19.5660 21.3570 ;
        RECT 19.4320 20.2635 19.4580 21.3570 ;
        RECT 19.3240 20.2635 19.3500 21.3570 ;
        RECT 19.2160 20.2635 19.2420 21.3570 ;
        RECT 19.1080 20.2635 19.1340 21.3570 ;
        RECT 19.0000 20.2635 19.0260 21.3570 ;
        RECT 18.8920 20.2635 18.9180 21.3570 ;
        RECT 18.7840 20.2635 18.8100 21.3570 ;
        RECT 18.6760 20.2635 18.7020 21.3570 ;
        RECT 18.5680 20.2635 18.5940 21.3570 ;
        RECT 18.4600 20.2635 18.4860 21.3570 ;
        RECT 18.3520 20.2635 18.3780 21.3570 ;
        RECT 18.2440 20.2635 18.2700 21.3570 ;
        RECT 18.1360 20.2635 18.1620 21.3570 ;
        RECT 18.0280 20.2635 18.0540 21.3570 ;
        RECT 17.9200 20.2635 17.9460 21.3570 ;
        RECT 17.8120 20.2635 17.8380 21.3570 ;
        RECT 17.7040 20.2635 17.7300 21.3570 ;
        RECT 17.5960 20.2635 17.6220 21.3570 ;
        RECT 17.4880 20.2635 17.5140 21.3570 ;
        RECT 17.3800 20.2635 17.4060 21.3570 ;
        RECT 17.2720 20.2635 17.2980 21.3570 ;
        RECT 17.1640 20.2635 17.1900 21.3570 ;
        RECT 17.0560 20.2635 17.0820 21.3570 ;
        RECT 16.9480 20.2635 16.9740 21.3570 ;
        RECT 16.8400 20.2635 16.8660 21.3570 ;
        RECT 16.7320 20.2635 16.7580 21.3570 ;
        RECT 16.6240 20.2635 16.6500 21.3570 ;
        RECT 16.5160 20.2635 16.5420 21.3570 ;
        RECT 16.4080 20.2635 16.4340 21.3570 ;
        RECT 16.3000 20.2635 16.3260 21.3570 ;
        RECT 16.0870 20.2635 16.1640 21.3570 ;
        RECT 14.1940 20.2635 14.2710 21.3570 ;
        RECT 14.0320 20.2635 14.0580 21.3570 ;
        RECT 13.9240 20.2635 13.9500 21.3570 ;
        RECT 13.8160 20.2635 13.8420 21.3570 ;
        RECT 13.7080 20.2635 13.7340 21.3570 ;
        RECT 13.6000 20.2635 13.6260 21.3570 ;
        RECT 13.4920 20.2635 13.5180 21.3570 ;
        RECT 13.3840 20.2635 13.4100 21.3570 ;
        RECT 13.2760 20.2635 13.3020 21.3570 ;
        RECT 13.1680 20.2635 13.1940 21.3570 ;
        RECT 13.0600 20.2635 13.0860 21.3570 ;
        RECT 12.9520 20.2635 12.9780 21.3570 ;
        RECT 12.8440 20.2635 12.8700 21.3570 ;
        RECT 12.7360 20.2635 12.7620 21.3570 ;
        RECT 12.6280 20.2635 12.6540 21.3570 ;
        RECT 12.5200 20.2635 12.5460 21.3570 ;
        RECT 12.4120 20.2635 12.4380 21.3570 ;
        RECT 12.3040 20.2635 12.3300 21.3570 ;
        RECT 12.1960 20.2635 12.2220 21.3570 ;
        RECT 12.0880 20.2635 12.1140 21.3570 ;
        RECT 11.9800 20.2635 12.0060 21.3570 ;
        RECT 11.8720 20.2635 11.8980 21.3570 ;
        RECT 11.7640 20.2635 11.7900 21.3570 ;
        RECT 11.6560 20.2635 11.6820 21.3570 ;
        RECT 11.5480 20.2635 11.5740 21.3570 ;
        RECT 11.4400 20.2635 11.4660 21.3570 ;
        RECT 11.3320 20.2635 11.3580 21.3570 ;
        RECT 11.2240 20.2635 11.2500 21.3570 ;
        RECT 11.1160 20.2635 11.1420 21.3570 ;
        RECT 11.0080 20.2635 11.0340 21.3570 ;
        RECT 10.9000 20.2635 10.9260 21.3570 ;
        RECT 10.7920 20.2635 10.8180 21.3570 ;
        RECT 10.6840 20.2635 10.7100 21.3570 ;
        RECT 10.5760 20.2635 10.6020 21.3570 ;
        RECT 10.4680 20.2635 10.4940 21.3570 ;
        RECT 10.3600 20.2635 10.3860 21.3570 ;
        RECT 10.2520 20.2635 10.2780 21.3570 ;
        RECT 10.1440 20.2635 10.1700 21.3570 ;
        RECT 10.0360 20.2635 10.0620 21.3570 ;
        RECT 9.9280 20.2635 9.9540 21.3570 ;
        RECT 9.8200 20.2635 9.8460 21.3570 ;
        RECT 9.7120 20.2635 9.7380 21.3570 ;
        RECT 9.6040 20.2635 9.6300 21.3570 ;
        RECT 9.4960 20.2635 9.5220 21.3570 ;
        RECT 9.3880 20.2635 9.4140 21.3570 ;
        RECT 9.2800 20.2635 9.3060 21.3570 ;
        RECT 9.1720 20.2635 9.1980 21.3570 ;
        RECT 9.0640 20.2635 9.0900 21.3570 ;
        RECT 8.9560 20.2635 8.9820 21.3570 ;
        RECT 8.8480 20.2635 8.8740 21.3570 ;
        RECT 8.7400 20.2635 8.7660 21.3570 ;
        RECT 8.6320 20.2635 8.6580 21.3570 ;
        RECT 8.5240 20.2635 8.5500 21.3570 ;
        RECT 8.4160 20.2635 8.4420 21.3570 ;
        RECT 8.3080 20.2635 8.3340 21.3570 ;
        RECT 8.2000 20.2635 8.2260 21.3570 ;
        RECT 8.0920 20.2635 8.1180 21.3570 ;
        RECT 7.9840 20.2635 8.0100 21.3570 ;
        RECT 7.8760 20.2635 7.9020 21.3570 ;
        RECT 7.7680 20.2635 7.7940 21.3570 ;
        RECT 7.6600 20.2635 7.6860 21.3570 ;
        RECT 7.5520 20.2635 7.5780 21.3570 ;
        RECT 7.4440 20.2635 7.4700 21.3570 ;
        RECT 7.3360 20.2635 7.3620 21.3570 ;
        RECT 7.2280 20.2635 7.2540 21.3570 ;
        RECT 7.1200 20.2635 7.1460 21.3570 ;
        RECT 7.0120 20.2635 7.0380 21.3570 ;
        RECT 6.9040 20.2635 6.9300 21.3570 ;
        RECT 6.7960 20.2635 6.8220 21.3570 ;
        RECT 6.6880 20.2635 6.7140 21.3570 ;
        RECT 6.5800 20.2635 6.6060 21.3570 ;
        RECT 6.4720 20.2635 6.4980 21.3570 ;
        RECT 6.3640 20.2635 6.3900 21.3570 ;
        RECT 6.2560 20.2635 6.2820 21.3570 ;
        RECT 6.1480 20.2635 6.1740 21.3570 ;
        RECT 6.0400 20.2635 6.0660 21.3570 ;
        RECT 5.9320 20.2635 5.9580 21.3570 ;
        RECT 5.8240 20.2635 5.8500 21.3570 ;
        RECT 5.7160 20.2635 5.7420 21.3570 ;
        RECT 5.6080 20.2635 5.6340 21.3570 ;
        RECT 5.5000 20.2635 5.5260 21.3570 ;
        RECT 5.3920 20.2635 5.4180 21.3570 ;
        RECT 5.2840 20.2635 5.3100 21.3570 ;
        RECT 5.1760 20.2635 5.2020 21.3570 ;
        RECT 5.0680 20.2635 5.0940 21.3570 ;
        RECT 4.9600 20.2635 4.9860 21.3570 ;
        RECT 4.8520 20.2635 4.8780 21.3570 ;
        RECT 4.7440 20.2635 4.7700 21.3570 ;
        RECT 4.6360 20.2635 4.6620 21.3570 ;
        RECT 4.5280 20.2635 4.5540 21.3570 ;
        RECT 4.4200 20.2635 4.4460 21.3570 ;
        RECT 4.3120 20.2635 4.3380 21.3570 ;
        RECT 4.2040 20.2635 4.2300 21.3570 ;
        RECT 4.0960 20.2635 4.1220 21.3570 ;
        RECT 3.9880 20.2635 4.0140 21.3570 ;
        RECT 3.8800 20.2635 3.9060 21.3570 ;
        RECT 3.7720 20.2635 3.7980 21.3570 ;
        RECT 3.6640 20.2635 3.6900 21.3570 ;
        RECT 3.5560 20.2635 3.5820 21.3570 ;
        RECT 3.4480 20.2635 3.4740 21.3570 ;
        RECT 3.3400 20.2635 3.3660 21.3570 ;
        RECT 3.2320 20.2635 3.2580 21.3570 ;
        RECT 3.1240 20.2635 3.1500 21.3570 ;
        RECT 3.0160 20.2635 3.0420 21.3570 ;
        RECT 2.9080 20.2635 2.9340 21.3570 ;
        RECT 2.8000 20.2635 2.8260 21.3570 ;
        RECT 2.6920 20.2635 2.7180 21.3570 ;
        RECT 2.5840 20.2635 2.6100 21.3570 ;
        RECT 2.4760 20.2635 2.5020 21.3570 ;
        RECT 2.3680 20.2635 2.3940 21.3570 ;
        RECT 2.2600 20.2635 2.2860 21.3570 ;
        RECT 2.1520 20.2635 2.1780 21.3570 ;
        RECT 2.0440 20.2635 2.0700 21.3570 ;
        RECT 1.9360 20.2635 1.9620 21.3570 ;
        RECT 1.8280 20.2635 1.8540 21.3570 ;
        RECT 1.7200 20.2635 1.7460 21.3570 ;
        RECT 1.6120 20.2635 1.6380 21.3570 ;
        RECT 1.5040 20.2635 1.5300 21.3570 ;
        RECT 1.3960 20.2635 1.4220 21.3570 ;
        RECT 1.2880 20.2635 1.3140 21.3570 ;
        RECT 1.1800 20.2635 1.2060 21.3570 ;
        RECT 1.0720 20.2635 1.0980 21.3570 ;
        RECT 0.9640 20.2635 0.9900 21.3570 ;
        RECT 0.8560 20.2635 0.8820 21.3570 ;
        RECT 0.7480 20.2635 0.7740 21.3570 ;
        RECT 0.6400 20.2635 0.6660 21.3570 ;
        RECT 0.5320 20.2635 0.5580 21.3570 ;
        RECT 0.4240 20.2635 0.4500 21.3570 ;
        RECT 0.3160 20.2635 0.3420 21.3570 ;
        RECT 0.2080 20.2635 0.2340 21.3570 ;
        RECT 0.0050 20.2635 0.0900 21.3570 ;
        RECT 15.5530 21.3435 15.6810 22.4370 ;
        RECT 15.5390 22.0090 15.6810 22.3315 ;
        RECT 15.3190 21.7360 15.4530 22.4370 ;
        RECT 15.2960 22.0710 15.4530 22.3290 ;
        RECT 15.3190 21.3435 15.4170 22.4370 ;
        RECT 15.3190 21.4645 15.4310 21.7040 ;
        RECT 15.3190 21.3435 15.4530 21.4325 ;
        RECT 15.0940 21.7940 15.2280 22.4370 ;
        RECT 15.0940 21.3435 15.1920 22.4370 ;
        RECT 14.6770 21.3435 14.7600 22.4370 ;
        RECT 14.6770 21.4320 14.7740 22.3675 ;
        RECT 30.2680 21.3435 30.3530 22.4370 ;
        RECT 30.1240 21.3435 30.1500 22.4370 ;
        RECT 30.0160 21.3435 30.0420 22.4370 ;
        RECT 29.9080 21.3435 29.9340 22.4370 ;
        RECT 29.8000 21.3435 29.8260 22.4370 ;
        RECT 29.6920 21.3435 29.7180 22.4370 ;
        RECT 29.5840 21.3435 29.6100 22.4370 ;
        RECT 29.4760 21.3435 29.5020 22.4370 ;
        RECT 29.3680 21.3435 29.3940 22.4370 ;
        RECT 29.2600 21.3435 29.2860 22.4370 ;
        RECT 29.1520 21.3435 29.1780 22.4370 ;
        RECT 29.0440 21.3435 29.0700 22.4370 ;
        RECT 28.9360 21.3435 28.9620 22.4370 ;
        RECT 28.8280 21.3435 28.8540 22.4370 ;
        RECT 28.7200 21.3435 28.7460 22.4370 ;
        RECT 28.6120 21.3435 28.6380 22.4370 ;
        RECT 28.5040 21.3435 28.5300 22.4370 ;
        RECT 28.3960 21.3435 28.4220 22.4370 ;
        RECT 28.2880 21.3435 28.3140 22.4370 ;
        RECT 28.1800 21.3435 28.2060 22.4370 ;
        RECT 28.0720 21.3435 28.0980 22.4370 ;
        RECT 27.9640 21.3435 27.9900 22.4370 ;
        RECT 27.8560 21.3435 27.8820 22.4370 ;
        RECT 27.7480 21.3435 27.7740 22.4370 ;
        RECT 27.6400 21.3435 27.6660 22.4370 ;
        RECT 27.5320 21.3435 27.5580 22.4370 ;
        RECT 27.4240 21.3435 27.4500 22.4370 ;
        RECT 27.3160 21.3435 27.3420 22.4370 ;
        RECT 27.2080 21.3435 27.2340 22.4370 ;
        RECT 27.1000 21.3435 27.1260 22.4370 ;
        RECT 26.9920 21.3435 27.0180 22.4370 ;
        RECT 26.8840 21.3435 26.9100 22.4370 ;
        RECT 26.7760 21.3435 26.8020 22.4370 ;
        RECT 26.6680 21.3435 26.6940 22.4370 ;
        RECT 26.5600 21.3435 26.5860 22.4370 ;
        RECT 26.4520 21.3435 26.4780 22.4370 ;
        RECT 26.3440 21.3435 26.3700 22.4370 ;
        RECT 26.2360 21.3435 26.2620 22.4370 ;
        RECT 26.1280 21.3435 26.1540 22.4370 ;
        RECT 26.0200 21.3435 26.0460 22.4370 ;
        RECT 25.9120 21.3435 25.9380 22.4370 ;
        RECT 25.8040 21.3435 25.8300 22.4370 ;
        RECT 25.6960 21.3435 25.7220 22.4370 ;
        RECT 25.5880 21.3435 25.6140 22.4370 ;
        RECT 25.4800 21.3435 25.5060 22.4370 ;
        RECT 25.3720 21.3435 25.3980 22.4370 ;
        RECT 25.2640 21.3435 25.2900 22.4370 ;
        RECT 25.1560 21.3435 25.1820 22.4370 ;
        RECT 25.0480 21.3435 25.0740 22.4370 ;
        RECT 24.9400 21.3435 24.9660 22.4370 ;
        RECT 24.8320 21.3435 24.8580 22.4370 ;
        RECT 24.7240 21.3435 24.7500 22.4370 ;
        RECT 24.6160 21.3435 24.6420 22.4370 ;
        RECT 24.5080 21.3435 24.5340 22.4370 ;
        RECT 24.4000 21.3435 24.4260 22.4370 ;
        RECT 24.2920 21.3435 24.3180 22.4370 ;
        RECT 24.1840 21.3435 24.2100 22.4370 ;
        RECT 24.0760 21.3435 24.1020 22.4370 ;
        RECT 23.9680 21.3435 23.9940 22.4370 ;
        RECT 23.8600 21.3435 23.8860 22.4370 ;
        RECT 23.7520 21.3435 23.7780 22.4370 ;
        RECT 23.6440 21.3435 23.6700 22.4370 ;
        RECT 23.5360 21.3435 23.5620 22.4370 ;
        RECT 23.4280 21.3435 23.4540 22.4370 ;
        RECT 23.3200 21.3435 23.3460 22.4370 ;
        RECT 23.2120 21.3435 23.2380 22.4370 ;
        RECT 23.1040 21.3435 23.1300 22.4370 ;
        RECT 22.9960 21.3435 23.0220 22.4370 ;
        RECT 22.8880 21.3435 22.9140 22.4370 ;
        RECT 22.7800 21.3435 22.8060 22.4370 ;
        RECT 22.6720 21.3435 22.6980 22.4370 ;
        RECT 22.5640 21.3435 22.5900 22.4370 ;
        RECT 22.4560 21.3435 22.4820 22.4370 ;
        RECT 22.3480 21.3435 22.3740 22.4370 ;
        RECT 22.2400 21.3435 22.2660 22.4370 ;
        RECT 22.1320 21.3435 22.1580 22.4370 ;
        RECT 22.0240 21.3435 22.0500 22.4370 ;
        RECT 21.9160 21.3435 21.9420 22.4370 ;
        RECT 21.8080 21.3435 21.8340 22.4370 ;
        RECT 21.7000 21.3435 21.7260 22.4370 ;
        RECT 21.5920 21.3435 21.6180 22.4370 ;
        RECT 21.4840 21.3435 21.5100 22.4370 ;
        RECT 21.3760 21.3435 21.4020 22.4370 ;
        RECT 21.2680 21.3435 21.2940 22.4370 ;
        RECT 21.1600 21.3435 21.1860 22.4370 ;
        RECT 21.0520 21.3435 21.0780 22.4370 ;
        RECT 20.9440 21.3435 20.9700 22.4370 ;
        RECT 20.8360 21.3435 20.8620 22.4370 ;
        RECT 20.7280 21.3435 20.7540 22.4370 ;
        RECT 20.6200 21.3435 20.6460 22.4370 ;
        RECT 20.5120 21.3435 20.5380 22.4370 ;
        RECT 20.4040 21.3435 20.4300 22.4370 ;
        RECT 20.2960 21.3435 20.3220 22.4370 ;
        RECT 20.1880 21.3435 20.2140 22.4370 ;
        RECT 20.0800 21.3435 20.1060 22.4370 ;
        RECT 19.9720 21.3435 19.9980 22.4370 ;
        RECT 19.8640 21.3435 19.8900 22.4370 ;
        RECT 19.7560 21.3435 19.7820 22.4370 ;
        RECT 19.6480 21.3435 19.6740 22.4370 ;
        RECT 19.5400 21.3435 19.5660 22.4370 ;
        RECT 19.4320 21.3435 19.4580 22.4370 ;
        RECT 19.3240 21.3435 19.3500 22.4370 ;
        RECT 19.2160 21.3435 19.2420 22.4370 ;
        RECT 19.1080 21.3435 19.1340 22.4370 ;
        RECT 19.0000 21.3435 19.0260 22.4370 ;
        RECT 18.8920 21.3435 18.9180 22.4370 ;
        RECT 18.7840 21.3435 18.8100 22.4370 ;
        RECT 18.6760 21.3435 18.7020 22.4370 ;
        RECT 18.5680 21.3435 18.5940 22.4370 ;
        RECT 18.4600 21.3435 18.4860 22.4370 ;
        RECT 18.3520 21.3435 18.3780 22.4370 ;
        RECT 18.2440 21.3435 18.2700 22.4370 ;
        RECT 18.1360 21.3435 18.1620 22.4370 ;
        RECT 18.0280 21.3435 18.0540 22.4370 ;
        RECT 17.9200 21.3435 17.9460 22.4370 ;
        RECT 17.8120 21.3435 17.8380 22.4370 ;
        RECT 17.7040 21.3435 17.7300 22.4370 ;
        RECT 17.5960 21.3435 17.6220 22.4370 ;
        RECT 17.4880 21.3435 17.5140 22.4370 ;
        RECT 17.3800 21.3435 17.4060 22.4370 ;
        RECT 17.2720 21.3435 17.2980 22.4370 ;
        RECT 17.1640 21.3435 17.1900 22.4370 ;
        RECT 17.0560 21.3435 17.0820 22.4370 ;
        RECT 16.9480 21.3435 16.9740 22.4370 ;
        RECT 16.8400 21.3435 16.8660 22.4370 ;
        RECT 16.7320 21.3435 16.7580 22.4370 ;
        RECT 16.6240 21.3435 16.6500 22.4370 ;
        RECT 16.5160 21.3435 16.5420 22.4370 ;
        RECT 16.4080 21.3435 16.4340 22.4370 ;
        RECT 16.3000 21.3435 16.3260 22.4370 ;
        RECT 16.0870 21.3435 16.1640 22.4370 ;
        RECT 14.1940 21.3435 14.2710 22.4370 ;
        RECT 14.0320 21.3435 14.0580 22.4370 ;
        RECT 13.9240 21.3435 13.9500 22.4370 ;
        RECT 13.8160 21.3435 13.8420 22.4370 ;
        RECT 13.7080 21.3435 13.7340 22.4370 ;
        RECT 13.6000 21.3435 13.6260 22.4370 ;
        RECT 13.4920 21.3435 13.5180 22.4370 ;
        RECT 13.3840 21.3435 13.4100 22.4370 ;
        RECT 13.2760 21.3435 13.3020 22.4370 ;
        RECT 13.1680 21.3435 13.1940 22.4370 ;
        RECT 13.0600 21.3435 13.0860 22.4370 ;
        RECT 12.9520 21.3435 12.9780 22.4370 ;
        RECT 12.8440 21.3435 12.8700 22.4370 ;
        RECT 12.7360 21.3435 12.7620 22.4370 ;
        RECT 12.6280 21.3435 12.6540 22.4370 ;
        RECT 12.5200 21.3435 12.5460 22.4370 ;
        RECT 12.4120 21.3435 12.4380 22.4370 ;
        RECT 12.3040 21.3435 12.3300 22.4370 ;
        RECT 12.1960 21.3435 12.2220 22.4370 ;
        RECT 12.0880 21.3435 12.1140 22.4370 ;
        RECT 11.9800 21.3435 12.0060 22.4370 ;
        RECT 11.8720 21.3435 11.8980 22.4370 ;
        RECT 11.7640 21.3435 11.7900 22.4370 ;
        RECT 11.6560 21.3435 11.6820 22.4370 ;
        RECT 11.5480 21.3435 11.5740 22.4370 ;
        RECT 11.4400 21.3435 11.4660 22.4370 ;
        RECT 11.3320 21.3435 11.3580 22.4370 ;
        RECT 11.2240 21.3435 11.2500 22.4370 ;
        RECT 11.1160 21.3435 11.1420 22.4370 ;
        RECT 11.0080 21.3435 11.0340 22.4370 ;
        RECT 10.9000 21.3435 10.9260 22.4370 ;
        RECT 10.7920 21.3435 10.8180 22.4370 ;
        RECT 10.6840 21.3435 10.7100 22.4370 ;
        RECT 10.5760 21.3435 10.6020 22.4370 ;
        RECT 10.4680 21.3435 10.4940 22.4370 ;
        RECT 10.3600 21.3435 10.3860 22.4370 ;
        RECT 10.2520 21.3435 10.2780 22.4370 ;
        RECT 10.1440 21.3435 10.1700 22.4370 ;
        RECT 10.0360 21.3435 10.0620 22.4370 ;
        RECT 9.9280 21.3435 9.9540 22.4370 ;
        RECT 9.8200 21.3435 9.8460 22.4370 ;
        RECT 9.7120 21.3435 9.7380 22.4370 ;
        RECT 9.6040 21.3435 9.6300 22.4370 ;
        RECT 9.4960 21.3435 9.5220 22.4370 ;
        RECT 9.3880 21.3435 9.4140 22.4370 ;
        RECT 9.2800 21.3435 9.3060 22.4370 ;
        RECT 9.1720 21.3435 9.1980 22.4370 ;
        RECT 9.0640 21.3435 9.0900 22.4370 ;
        RECT 8.9560 21.3435 8.9820 22.4370 ;
        RECT 8.8480 21.3435 8.8740 22.4370 ;
        RECT 8.7400 21.3435 8.7660 22.4370 ;
        RECT 8.6320 21.3435 8.6580 22.4370 ;
        RECT 8.5240 21.3435 8.5500 22.4370 ;
        RECT 8.4160 21.3435 8.4420 22.4370 ;
        RECT 8.3080 21.3435 8.3340 22.4370 ;
        RECT 8.2000 21.3435 8.2260 22.4370 ;
        RECT 8.0920 21.3435 8.1180 22.4370 ;
        RECT 7.9840 21.3435 8.0100 22.4370 ;
        RECT 7.8760 21.3435 7.9020 22.4370 ;
        RECT 7.7680 21.3435 7.7940 22.4370 ;
        RECT 7.6600 21.3435 7.6860 22.4370 ;
        RECT 7.5520 21.3435 7.5780 22.4370 ;
        RECT 7.4440 21.3435 7.4700 22.4370 ;
        RECT 7.3360 21.3435 7.3620 22.4370 ;
        RECT 7.2280 21.3435 7.2540 22.4370 ;
        RECT 7.1200 21.3435 7.1460 22.4370 ;
        RECT 7.0120 21.3435 7.0380 22.4370 ;
        RECT 6.9040 21.3435 6.9300 22.4370 ;
        RECT 6.7960 21.3435 6.8220 22.4370 ;
        RECT 6.6880 21.3435 6.7140 22.4370 ;
        RECT 6.5800 21.3435 6.6060 22.4370 ;
        RECT 6.4720 21.3435 6.4980 22.4370 ;
        RECT 6.3640 21.3435 6.3900 22.4370 ;
        RECT 6.2560 21.3435 6.2820 22.4370 ;
        RECT 6.1480 21.3435 6.1740 22.4370 ;
        RECT 6.0400 21.3435 6.0660 22.4370 ;
        RECT 5.9320 21.3435 5.9580 22.4370 ;
        RECT 5.8240 21.3435 5.8500 22.4370 ;
        RECT 5.7160 21.3435 5.7420 22.4370 ;
        RECT 5.6080 21.3435 5.6340 22.4370 ;
        RECT 5.5000 21.3435 5.5260 22.4370 ;
        RECT 5.3920 21.3435 5.4180 22.4370 ;
        RECT 5.2840 21.3435 5.3100 22.4370 ;
        RECT 5.1760 21.3435 5.2020 22.4370 ;
        RECT 5.0680 21.3435 5.0940 22.4370 ;
        RECT 4.9600 21.3435 4.9860 22.4370 ;
        RECT 4.8520 21.3435 4.8780 22.4370 ;
        RECT 4.7440 21.3435 4.7700 22.4370 ;
        RECT 4.6360 21.3435 4.6620 22.4370 ;
        RECT 4.5280 21.3435 4.5540 22.4370 ;
        RECT 4.4200 21.3435 4.4460 22.4370 ;
        RECT 4.3120 21.3435 4.3380 22.4370 ;
        RECT 4.2040 21.3435 4.2300 22.4370 ;
        RECT 4.0960 21.3435 4.1220 22.4370 ;
        RECT 3.9880 21.3435 4.0140 22.4370 ;
        RECT 3.8800 21.3435 3.9060 22.4370 ;
        RECT 3.7720 21.3435 3.7980 22.4370 ;
        RECT 3.6640 21.3435 3.6900 22.4370 ;
        RECT 3.5560 21.3435 3.5820 22.4370 ;
        RECT 3.4480 21.3435 3.4740 22.4370 ;
        RECT 3.3400 21.3435 3.3660 22.4370 ;
        RECT 3.2320 21.3435 3.2580 22.4370 ;
        RECT 3.1240 21.3435 3.1500 22.4370 ;
        RECT 3.0160 21.3435 3.0420 22.4370 ;
        RECT 2.9080 21.3435 2.9340 22.4370 ;
        RECT 2.8000 21.3435 2.8260 22.4370 ;
        RECT 2.6920 21.3435 2.7180 22.4370 ;
        RECT 2.5840 21.3435 2.6100 22.4370 ;
        RECT 2.4760 21.3435 2.5020 22.4370 ;
        RECT 2.3680 21.3435 2.3940 22.4370 ;
        RECT 2.2600 21.3435 2.2860 22.4370 ;
        RECT 2.1520 21.3435 2.1780 22.4370 ;
        RECT 2.0440 21.3435 2.0700 22.4370 ;
        RECT 1.9360 21.3435 1.9620 22.4370 ;
        RECT 1.8280 21.3435 1.8540 22.4370 ;
        RECT 1.7200 21.3435 1.7460 22.4370 ;
        RECT 1.6120 21.3435 1.6380 22.4370 ;
        RECT 1.5040 21.3435 1.5300 22.4370 ;
        RECT 1.3960 21.3435 1.4220 22.4370 ;
        RECT 1.2880 21.3435 1.3140 22.4370 ;
        RECT 1.1800 21.3435 1.2060 22.4370 ;
        RECT 1.0720 21.3435 1.0980 22.4370 ;
        RECT 0.9640 21.3435 0.9900 22.4370 ;
        RECT 0.8560 21.3435 0.8820 22.4370 ;
        RECT 0.7480 21.3435 0.7740 22.4370 ;
        RECT 0.6400 21.3435 0.6660 22.4370 ;
        RECT 0.5320 21.3435 0.5580 22.4370 ;
        RECT 0.4240 21.3435 0.4500 22.4370 ;
        RECT 0.3160 21.3435 0.3420 22.4370 ;
        RECT 0.2080 21.3435 0.2340 22.4370 ;
        RECT 0.0050 21.3435 0.0900 22.4370 ;
        RECT 15.5530 22.4235 15.6810 23.5170 ;
        RECT 15.5390 23.0890 15.6810 23.4115 ;
        RECT 15.3190 22.8160 15.4530 23.5170 ;
        RECT 15.2960 23.1510 15.4530 23.4090 ;
        RECT 15.3190 22.4235 15.4170 23.5170 ;
        RECT 15.3190 22.5445 15.4310 22.7840 ;
        RECT 15.3190 22.4235 15.4530 22.5125 ;
        RECT 15.0940 22.8740 15.2280 23.5170 ;
        RECT 15.0940 22.4235 15.1920 23.5170 ;
        RECT 14.6770 22.4235 14.7600 23.5170 ;
        RECT 14.6770 22.5120 14.7740 23.4475 ;
        RECT 30.2680 22.4235 30.3530 23.5170 ;
        RECT 30.1240 22.4235 30.1500 23.5170 ;
        RECT 30.0160 22.4235 30.0420 23.5170 ;
        RECT 29.9080 22.4235 29.9340 23.5170 ;
        RECT 29.8000 22.4235 29.8260 23.5170 ;
        RECT 29.6920 22.4235 29.7180 23.5170 ;
        RECT 29.5840 22.4235 29.6100 23.5170 ;
        RECT 29.4760 22.4235 29.5020 23.5170 ;
        RECT 29.3680 22.4235 29.3940 23.5170 ;
        RECT 29.2600 22.4235 29.2860 23.5170 ;
        RECT 29.1520 22.4235 29.1780 23.5170 ;
        RECT 29.0440 22.4235 29.0700 23.5170 ;
        RECT 28.9360 22.4235 28.9620 23.5170 ;
        RECT 28.8280 22.4235 28.8540 23.5170 ;
        RECT 28.7200 22.4235 28.7460 23.5170 ;
        RECT 28.6120 22.4235 28.6380 23.5170 ;
        RECT 28.5040 22.4235 28.5300 23.5170 ;
        RECT 28.3960 22.4235 28.4220 23.5170 ;
        RECT 28.2880 22.4235 28.3140 23.5170 ;
        RECT 28.1800 22.4235 28.2060 23.5170 ;
        RECT 28.0720 22.4235 28.0980 23.5170 ;
        RECT 27.9640 22.4235 27.9900 23.5170 ;
        RECT 27.8560 22.4235 27.8820 23.5170 ;
        RECT 27.7480 22.4235 27.7740 23.5170 ;
        RECT 27.6400 22.4235 27.6660 23.5170 ;
        RECT 27.5320 22.4235 27.5580 23.5170 ;
        RECT 27.4240 22.4235 27.4500 23.5170 ;
        RECT 27.3160 22.4235 27.3420 23.5170 ;
        RECT 27.2080 22.4235 27.2340 23.5170 ;
        RECT 27.1000 22.4235 27.1260 23.5170 ;
        RECT 26.9920 22.4235 27.0180 23.5170 ;
        RECT 26.8840 22.4235 26.9100 23.5170 ;
        RECT 26.7760 22.4235 26.8020 23.5170 ;
        RECT 26.6680 22.4235 26.6940 23.5170 ;
        RECT 26.5600 22.4235 26.5860 23.5170 ;
        RECT 26.4520 22.4235 26.4780 23.5170 ;
        RECT 26.3440 22.4235 26.3700 23.5170 ;
        RECT 26.2360 22.4235 26.2620 23.5170 ;
        RECT 26.1280 22.4235 26.1540 23.5170 ;
        RECT 26.0200 22.4235 26.0460 23.5170 ;
        RECT 25.9120 22.4235 25.9380 23.5170 ;
        RECT 25.8040 22.4235 25.8300 23.5170 ;
        RECT 25.6960 22.4235 25.7220 23.5170 ;
        RECT 25.5880 22.4235 25.6140 23.5170 ;
        RECT 25.4800 22.4235 25.5060 23.5170 ;
        RECT 25.3720 22.4235 25.3980 23.5170 ;
        RECT 25.2640 22.4235 25.2900 23.5170 ;
        RECT 25.1560 22.4235 25.1820 23.5170 ;
        RECT 25.0480 22.4235 25.0740 23.5170 ;
        RECT 24.9400 22.4235 24.9660 23.5170 ;
        RECT 24.8320 22.4235 24.8580 23.5170 ;
        RECT 24.7240 22.4235 24.7500 23.5170 ;
        RECT 24.6160 22.4235 24.6420 23.5170 ;
        RECT 24.5080 22.4235 24.5340 23.5170 ;
        RECT 24.4000 22.4235 24.4260 23.5170 ;
        RECT 24.2920 22.4235 24.3180 23.5170 ;
        RECT 24.1840 22.4235 24.2100 23.5170 ;
        RECT 24.0760 22.4235 24.1020 23.5170 ;
        RECT 23.9680 22.4235 23.9940 23.5170 ;
        RECT 23.8600 22.4235 23.8860 23.5170 ;
        RECT 23.7520 22.4235 23.7780 23.5170 ;
        RECT 23.6440 22.4235 23.6700 23.5170 ;
        RECT 23.5360 22.4235 23.5620 23.5170 ;
        RECT 23.4280 22.4235 23.4540 23.5170 ;
        RECT 23.3200 22.4235 23.3460 23.5170 ;
        RECT 23.2120 22.4235 23.2380 23.5170 ;
        RECT 23.1040 22.4235 23.1300 23.5170 ;
        RECT 22.9960 22.4235 23.0220 23.5170 ;
        RECT 22.8880 22.4235 22.9140 23.5170 ;
        RECT 22.7800 22.4235 22.8060 23.5170 ;
        RECT 22.6720 22.4235 22.6980 23.5170 ;
        RECT 22.5640 22.4235 22.5900 23.5170 ;
        RECT 22.4560 22.4235 22.4820 23.5170 ;
        RECT 22.3480 22.4235 22.3740 23.5170 ;
        RECT 22.2400 22.4235 22.2660 23.5170 ;
        RECT 22.1320 22.4235 22.1580 23.5170 ;
        RECT 22.0240 22.4235 22.0500 23.5170 ;
        RECT 21.9160 22.4235 21.9420 23.5170 ;
        RECT 21.8080 22.4235 21.8340 23.5170 ;
        RECT 21.7000 22.4235 21.7260 23.5170 ;
        RECT 21.5920 22.4235 21.6180 23.5170 ;
        RECT 21.4840 22.4235 21.5100 23.5170 ;
        RECT 21.3760 22.4235 21.4020 23.5170 ;
        RECT 21.2680 22.4235 21.2940 23.5170 ;
        RECT 21.1600 22.4235 21.1860 23.5170 ;
        RECT 21.0520 22.4235 21.0780 23.5170 ;
        RECT 20.9440 22.4235 20.9700 23.5170 ;
        RECT 20.8360 22.4235 20.8620 23.5170 ;
        RECT 20.7280 22.4235 20.7540 23.5170 ;
        RECT 20.6200 22.4235 20.6460 23.5170 ;
        RECT 20.5120 22.4235 20.5380 23.5170 ;
        RECT 20.4040 22.4235 20.4300 23.5170 ;
        RECT 20.2960 22.4235 20.3220 23.5170 ;
        RECT 20.1880 22.4235 20.2140 23.5170 ;
        RECT 20.0800 22.4235 20.1060 23.5170 ;
        RECT 19.9720 22.4235 19.9980 23.5170 ;
        RECT 19.8640 22.4235 19.8900 23.5170 ;
        RECT 19.7560 22.4235 19.7820 23.5170 ;
        RECT 19.6480 22.4235 19.6740 23.5170 ;
        RECT 19.5400 22.4235 19.5660 23.5170 ;
        RECT 19.4320 22.4235 19.4580 23.5170 ;
        RECT 19.3240 22.4235 19.3500 23.5170 ;
        RECT 19.2160 22.4235 19.2420 23.5170 ;
        RECT 19.1080 22.4235 19.1340 23.5170 ;
        RECT 19.0000 22.4235 19.0260 23.5170 ;
        RECT 18.8920 22.4235 18.9180 23.5170 ;
        RECT 18.7840 22.4235 18.8100 23.5170 ;
        RECT 18.6760 22.4235 18.7020 23.5170 ;
        RECT 18.5680 22.4235 18.5940 23.5170 ;
        RECT 18.4600 22.4235 18.4860 23.5170 ;
        RECT 18.3520 22.4235 18.3780 23.5170 ;
        RECT 18.2440 22.4235 18.2700 23.5170 ;
        RECT 18.1360 22.4235 18.1620 23.5170 ;
        RECT 18.0280 22.4235 18.0540 23.5170 ;
        RECT 17.9200 22.4235 17.9460 23.5170 ;
        RECT 17.8120 22.4235 17.8380 23.5170 ;
        RECT 17.7040 22.4235 17.7300 23.5170 ;
        RECT 17.5960 22.4235 17.6220 23.5170 ;
        RECT 17.4880 22.4235 17.5140 23.5170 ;
        RECT 17.3800 22.4235 17.4060 23.5170 ;
        RECT 17.2720 22.4235 17.2980 23.5170 ;
        RECT 17.1640 22.4235 17.1900 23.5170 ;
        RECT 17.0560 22.4235 17.0820 23.5170 ;
        RECT 16.9480 22.4235 16.9740 23.5170 ;
        RECT 16.8400 22.4235 16.8660 23.5170 ;
        RECT 16.7320 22.4235 16.7580 23.5170 ;
        RECT 16.6240 22.4235 16.6500 23.5170 ;
        RECT 16.5160 22.4235 16.5420 23.5170 ;
        RECT 16.4080 22.4235 16.4340 23.5170 ;
        RECT 16.3000 22.4235 16.3260 23.5170 ;
        RECT 16.0870 22.4235 16.1640 23.5170 ;
        RECT 14.1940 22.4235 14.2710 23.5170 ;
        RECT 14.0320 22.4235 14.0580 23.5170 ;
        RECT 13.9240 22.4235 13.9500 23.5170 ;
        RECT 13.8160 22.4235 13.8420 23.5170 ;
        RECT 13.7080 22.4235 13.7340 23.5170 ;
        RECT 13.6000 22.4235 13.6260 23.5170 ;
        RECT 13.4920 22.4235 13.5180 23.5170 ;
        RECT 13.3840 22.4235 13.4100 23.5170 ;
        RECT 13.2760 22.4235 13.3020 23.5170 ;
        RECT 13.1680 22.4235 13.1940 23.5170 ;
        RECT 13.0600 22.4235 13.0860 23.5170 ;
        RECT 12.9520 22.4235 12.9780 23.5170 ;
        RECT 12.8440 22.4235 12.8700 23.5170 ;
        RECT 12.7360 22.4235 12.7620 23.5170 ;
        RECT 12.6280 22.4235 12.6540 23.5170 ;
        RECT 12.5200 22.4235 12.5460 23.5170 ;
        RECT 12.4120 22.4235 12.4380 23.5170 ;
        RECT 12.3040 22.4235 12.3300 23.5170 ;
        RECT 12.1960 22.4235 12.2220 23.5170 ;
        RECT 12.0880 22.4235 12.1140 23.5170 ;
        RECT 11.9800 22.4235 12.0060 23.5170 ;
        RECT 11.8720 22.4235 11.8980 23.5170 ;
        RECT 11.7640 22.4235 11.7900 23.5170 ;
        RECT 11.6560 22.4235 11.6820 23.5170 ;
        RECT 11.5480 22.4235 11.5740 23.5170 ;
        RECT 11.4400 22.4235 11.4660 23.5170 ;
        RECT 11.3320 22.4235 11.3580 23.5170 ;
        RECT 11.2240 22.4235 11.2500 23.5170 ;
        RECT 11.1160 22.4235 11.1420 23.5170 ;
        RECT 11.0080 22.4235 11.0340 23.5170 ;
        RECT 10.9000 22.4235 10.9260 23.5170 ;
        RECT 10.7920 22.4235 10.8180 23.5170 ;
        RECT 10.6840 22.4235 10.7100 23.5170 ;
        RECT 10.5760 22.4235 10.6020 23.5170 ;
        RECT 10.4680 22.4235 10.4940 23.5170 ;
        RECT 10.3600 22.4235 10.3860 23.5170 ;
        RECT 10.2520 22.4235 10.2780 23.5170 ;
        RECT 10.1440 22.4235 10.1700 23.5170 ;
        RECT 10.0360 22.4235 10.0620 23.5170 ;
        RECT 9.9280 22.4235 9.9540 23.5170 ;
        RECT 9.8200 22.4235 9.8460 23.5170 ;
        RECT 9.7120 22.4235 9.7380 23.5170 ;
        RECT 9.6040 22.4235 9.6300 23.5170 ;
        RECT 9.4960 22.4235 9.5220 23.5170 ;
        RECT 9.3880 22.4235 9.4140 23.5170 ;
        RECT 9.2800 22.4235 9.3060 23.5170 ;
        RECT 9.1720 22.4235 9.1980 23.5170 ;
        RECT 9.0640 22.4235 9.0900 23.5170 ;
        RECT 8.9560 22.4235 8.9820 23.5170 ;
        RECT 8.8480 22.4235 8.8740 23.5170 ;
        RECT 8.7400 22.4235 8.7660 23.5170 ;
        RECT 8.6320 22.4235 8.6580 23.5170 ;
        RECT 8.5240 22.4235 8.5500 23.5170 ;
        RECT 8.4160 22.4235 8.4420 23.5170 ;
        RECT 8.3080 22.4235 8.3340 23.5170 ;
        RECT 8.2000 22.4235 8.2260 23.5170 ;
        RECT 8.0920 22.4235 8.1180 23.5170 ;
        RECT 7.9840 22.4235 8.0100 23.5170 ;
        RECT 7.8760 22.4235 7.9020 23.5170 ;
        RECT 7.7680 22.4235 7.7940 23.5170 ;
        RECT 7.6600 22.4235 7.6860 23.5170 ;
        RECT 7.5520 22.4235 7.5780 23.5170 ;
        RECT 7.4440 22.4235 7.4700 23.5170 ;
        RECT 7.3360 22.4235 7.3620 23.5170 ;
        RECT 7.2280 22.4235 7.2540 23.5170 ;
        RECT 7.1200 22.4235 7.1460 23.5170 ;
        RECT 7.0120 22.4235 7.0380 23.5170 ;
        RECT 6.9040 22.4235 6.9300 23.5170 ;
        RECT 6.7960 22.4235 6.8220 23.5170 ;
        RECT 6.6880 22.4235 6.7140 23.5170 ;
        RECT 6.5800 22.4235 6.6060 23.5170 ;
        RECT 6.4720 22.4235 6.4980 23.5170 ;
        RECT 6.3640 22.4235 6.3900 23.5170 ;
        RECT 6.2560 22.4235 6.2820 23.5170 ;
        RECT 6.1480 22.4235 6.1740 23.5170 ;
        RECT 6.0400 22.4235 6.0660 23.5170 ;
        RECT 5.9320 22.4235 5.9580 23.5170 ;
        RECT 5.8240 22.4235 5.8500 23.5170 ;
        RECT 5.7160 22.4235 5.7420 23.5170 ;
        RECT 5.6080 22.4235 5.6340 23.5170 ;
        RECT 5.5000 22.4235 5.5260 23.5170 ;
        RECT 5.3920 22.4235 5.4180 23.5170 ;
        RECT 5.2840 22.4235 5.3100 23.5170 ;
        RECT 5.1760 22.4235 5.2020 23.5170 ;
        RECT 5.0680 22.4235 5.0940 23.5170 ;
        RECT 4.9600 22.4235 4.9860 23.5170 ;
        RECT 4.8520 22.4235 4.8780 23.5170 ;
        RECT 4.7440 22.4235 4.7700 23.5170 ;
        RECT 4.6360 22.4235 4.6620 23.5170 ;
        RECT 4.5280 22.4235 4.5540 23.5170 ;
        RECT 4.4200 22.4235 4.4460 23.5170 ;
        RECT 4.3120 22.4235 4.3380 23.5170 ;
        RECT 4.2040 22.4235 4.2300 23.5170 ;
        RECT 4.0960 22.4235 4.1220 23.5170 ;
        RECT 3.9880 22.4235 4.0140 23.5170 ;
        RECT 3.8800 22.4235 3.9060 23.5170 ;
        RECT 3.7720 22.4235 3.7980 23.5170 ;
        RECT 3.6640 22.4235 3.6900 23.5170 ;
        RECT 3.5560 22.4235 3.5820 23.5170 ;
        RECT 3.4480 22.4235 3.4740 23.5170 ;
        RECT 3.3400 22.4235 3.3660 23.5170 ;
        RECT 3.2320 22.4235 3.2580 23.5170 ;
        RECT 3.1240 22.4235 3.1500 23.5170 ;
        RECT 3.0160 22.4235 3.0420 23.5170 ;
        RECT 2.9080 22.4235 2.9340 23.5170 ;
        RECT 2.8000 22.4235 2.8260 23.5170 ;
        RECT 2.6920 22.4235 2.7180 23.5170 ;
        RECT 2.5840 22.4235 2.6100 23.5170 ;
        RECT 2.4760 22.4235 2.5020 23.5170 ;
        RECT 2.3680 22.4235 2.3940 23.5170 ;
        RECT 2.2600 22.4235 2.2860 23.5170 ;
        RECT 2.1520 22.4235 2.1780 23.5170 ;
        RECT 2.0440 22.4235 2.0700 23.5170 ;
        RECT 1.9360 22.4235 1.9620 23.5170 ;
        RECT 1.8280 22.4235 1.8540 23.5170 ;
        RECT 1.7200 22.4235 1.7460 23.5170 ;
        RECT 1.6120 22.4235 1.6380 23.5170 ;
        RECT 1.5040 22.4235 1.5300 23.5170 ;
        RECT 1.3960 22.4235 1.4220 23.5170 ;
        RECT 1.2880 22.4235 1.3140 23.5170 ;
        RECT 1.1800 22.4235 1.2060 23.5170 ;
        RECT 1.0720 22.4235 1.0980 23.5170 ;
        RECT 0.9640 22.4235 0.9900 23.5170 ;
        RECT 0.8560 22.4235 0.8820 23.5170 ;
        RECT 0.7480 22.4235 0.7740 23.5170 ;
        RECT 0.6400 22.4235 0.6660 23.5170 ;
        RECT 0.5320 22.4235 0.5580 23.5170 ;
        RECT 0.4240 22.4235 0.4500 23.5170 ;
        RECT 0.3160 22.4235 0.3420 23.5170 ;
        RECT 0.2080 22.4235 0.2340 23.5170 ;
        RECT 0.0050 22.4235 0.0900 23.5170 ;
        RECT 15.5530 23.5035 15.6810 24.5970 ;
        RECT 15.5390 24.1690 15.6810 24.4915 ;
        RECT 15.3190 23.8960 15.4530 24.5970 ;
        RECT 15.2960 24.2310 15.4530 24.4890 ;
        RECT 15.3190 23.5035 15.4170 24.5970 ;
        RECT 15.3190 23.6245 15.4310 23.8640 ;
        RECT 15.3190 23.5035 15.4530 23.5925 ;
        RECT 15.0940 23.9540 15.2280 24.5970 ;
        RECT 15.0940 23.5035 15.1920 24.5970 ;
        RECT 14.6770 23.5035 14.7600 24.5970 ;
        RECT 14.6770 23.5920 14.7740 24.5275 ;
        RECT 30.2680 23.5035 30.3530 24.5970 ;
        RECT 30.1240 23.5035 30.1500 24.5970 ;
        RECT 30.0160 23.5035 30.0420 24.5970 ;
        RECT 29.9080 23.5035 29.9340 24.5970 ;
        RECT 29.8000 23.5035 29.8260 24.5970 ;
        RECT 29.6920 23.5035 29.7180 24.5970 ;
        RECT 29.5840 23.5035 29.6100 24.5970 ;
        RECT 29.4760 23.5035 29.5020 24.5970 ;
        RECT 29.3680 23.5035 29.3940 24.5970 ;
        RECT 29.2600 23.5035 29.2860 24.5970 ;
        RECT 29.1520 23.5035 29.1780 24.5970 ;
        RECT 29.0440 23.5035 29.0700 24.5970 ;
        RECT 28.9360 23.5035 28.9620 24.5970 ;
        RECT 28.8280 23.5035 28.8540 24.5970 ;
        RECT 28.7200 23.5035 28.7460 24.5970 ;
        RECT 28.6120 23.5035 28.6380 24.5970 ;
        RECT 28.5040 23.5035 28.5300 24.5970 ;
        RECT 28.3960 23.5035 28.4220 24.5970 ;
        RECT 28.2880 23.5035 28.3140 24.5970 ;
        RECT 28.1800 23.5035 28.2060 24.5970 ;
        RECT 28.0720 23.5035 28.0980 24.5970 ;
        RECT 27.9640 23.5035 27.9900 24.5970 ;
        RECT 27.8560 23.5035 27.8820 24.5970 ;
        RECT 27.7480 23.5035 27.7740 24.5970 ;
        RECT 27.6400 23.5035 27.6660 24.5970 ;
        RECT 27.5320 23.5035 27.5580 24.5970 ;
        RECT 27.4240 23.5035 27.4500 24.5970 ;
        RECT 27.3160 23.5035 27.3420 24.5970 ;
        RECT 27.2080 23.5035 27.2340 24.5970 ;
        RECT 27.1000 23.5035 27.1260 24.5970 ;
        RECT 26.9920 23.5035 27.0180 24.5970 ;
        RECT 26.8840 23.5035 26.9100 24.5970 ;
        RECT 26.7760 23.5035 26.8020 24.5970 ;
        RECT 26.6680 23.5035 26.6940 24.5970 ;
        RECT 26.5600 23.5035 26.5860 24.5970 ;
        RECT 26.4520 23.5035 26.4780 24.5970 ;
        RECT 26.3440 23.5035 26.3700 24.5970 ;
        RECT 26.2360 23.5035 26.2620 24.5970 ;
        RECT 26.1280 23.5035 26.1540 24.5970 ;
        RECT 26.0200 23.5035 26.0460 24.5970 ;
        RECT 25.9120 23.5035 25.9380 24.5970 ;
        RECT 25.8040 23.5035 25.8300 24.5970 ;
        RECT 25.6960 23.5035 25.7220 24.5970 ;
        RECT 25.5880 23.5035 25.6140 24.5970 ;
        RECT 25.4800 23.5035 25.5060 24.5970 ;
        RECT 25.3720 23.5035 25.3980 24.5970 ;
        RECT 25.2640 23.5035 25.2900 24.5970 ;
        RECT 25.1560 23.5035 25.1820 24.5970 ;
        RECT 25.0480 23.5035 25.0740 24.5970 ;
        RECT 24.9400 23.5035 24.9660 24.5970 ;
        RECT 24.8320 23.5035 24.8580 24.5970 ;
        RECT 24.7240 23.5035 24.7500 24.5970 ;
        RECT 24.6160 23.5035 24.6420 24.5970 ;
        RECT 24.5080 23.5035 24.5340 24.5970 ;
        RECT 24.4000 23.5035 24.4260 24.5970 ;
        RECT 24.2920 23.5035 24.3180 24.5970 ;
        RECT 24.1840 23.5035 24.2100 24.5970 ;
        RECT 24.0760 23.5035 24.1020 24.5970 ;
        RECT 23.9680 23.5035 23.9940 24.5970 ;
        RECT 23.8600 23.5035 23.8860 24.5970 ;
        RECT 23.7520 23.5035 23.7780 24.5970 ;
        RECT 23.6440 23.5035 23.6700 24.5970 ;
        RECT 23.5360 23.5035 23.5620 24.5970 ;
        RECT 23.4280 23.5035 23.4540 24.5970 ;
        RECT 23.3200 23.5035 23.3460 24.5970 ;
        RECT 23.2120 23.5035 23.2380 24.5970 ;
        RECT 23.1040 23.5035 23.1300 24.5970 ;
        RECT 22.9960 23.5035 23.0220 24.5970 ;
        RECT 22.8880 23.5035 22.9140 24.5970 ;
        RECT 22.7800 23.5035 22.8060 24.5970 ;
        RECT 22.6720 23.5035 22.6980 24.5970 ;
        RECT 22.5640 23.5035 22.5900 24.5970 ;
        RECT 22.4560 23.5035 22.4820 24.5970 ;
        RECT 22.3480 23.5035 22.3740 24.5970 ;
        RECT 22.2400 23.5035 22.2660 24.5970 ;
        RECT 22.1320 23.5035 22.1580 24.5970 ;
        RECT 22.0240 23.5035 22.0500 24.5970 ;
        RECT 21.9160 23.5035 21.9420 24.5970 ;
        RECT 21.8080 23.5035 21.8340 24.5970 ;
        RECT 21.7000 23.5035 21.7260 24.5970 ;
        RECT 21.5920 23.5035 21.6180 24.5970 ;
        RECT 21.4840 23.5035 21.5100 24.5970 ;
        RECT 21.3760 23.5035 21.4020 24.5970 ;
        RECT 21.2680 23.5035 21.2940 24.5970 ;
        RECT 21.1600 23.5035 21.1860 24.5970 ;
        RECT 21.0520 23.5035 21.0780 24.5970 ;
        RECT 20.9440 23.5035 20.9700 24.5970 ;
        RECT 20.8360 23.5035 20.8620 24.5970 ;
        RECT 20.7280 23.5035 20.7540 24.5970 ;
        RECT 20.6200 23.5035 20.6460 24.5970 ;
        RECT 20.5120 23.5035 20.5380 24.5970 ;
        RECT 20.4040 23.5035 20.4300 24.5970 ;
        RECT 20.2960 23.5035 20.3220 24.5970 ;
        RECT 20.1880 23.5035 20.2140 24.5970 ;
        RECT 20.0800 23.5035 20.1060 24.5970 ;
        RECT 19.9720 23.5035 19.9980 24.5970 ;
        RECT 19.8640 23.5035 19.8900 24.5970 ;
        RECT 19.7560 23.5035 19.7820 24.5970 ;
        RECT 19.6480 23.5035 19.6740 24.5970 ;
        RECT 19.5400 23.5035 19.5660 24.5970 ;
        RECT 19.4320 23.5035 19.4580 24.5970 ;
        RECT 19.3240 23.5035 19.3500 24.5970 ;
        RECT 19.2160 23.5035 19.2420 24.5970 ;
        RECT 19.1080 23.5035 19.1340 24.5970 ;
        RECT 19.0000 23.5035 19.0260 24.5970 ;
        RECT 18.8920 23.5035 18.9180 24.5970 ;
        RECT 18.7840 23.5035 18.8100 24.5970 ;
        RECT 18.6760 23.5035 18.7020 24.5970 ;
        RECT 18.5680 23.5035 18.5940 24.5970 ;
        RECT 18.4600 23.5035 18.4860 24.5970 ;
        RECT 18.3520 23.5035 18.3780 24.5970 ;
        RECT 18.2440 23.5035 18.2700 24.5970 ;
        RECT 18.1360 23.5035 18.1620 24.5970 ;
        RECT 18.0280 23.5035 18.0540 24.5970 ;
        RECT 17.9200 23.5035 17.9460 24.5970 ;
        RECT 17.8120 23.5035 17.8380 24.5970 ;
        RECT 17.7040 23.5035 17.7300 24.5970 ;
        RECT 17.5960 23.5035 17.6220 24.5970 ;
        RECT 17.4880 23.5035 17.5140 24.5970 ;
        RECT 17.3800 23.5035 17.4060 24.5970 ;
        RECT 17.2720 23.5035 17.2980 24.5970 ;
        RECT 17.1640 23.5035 17.1900 24.5970 ;
        RECT 17.0560 23.5035 17.0820 24.5970 ;
        RECT 16.9480 23.5035 16.9740 24.5970 ;
        RECT 16.8400 23.5035 16.8660 24.5970 ;
        RECT 16.7320 23.5035 16.7580 24.5970 ;
        RECT 16.6240 23.5035 16.6500 24.5970 ;
        RECT 16.5160 23.5035 16.5420 24.5970 ;
        RECT 16.4080 23.5035 16.4340 24.5970 ;
        RECT 16.3000 23.5035 16.3260 24.5970 ;
        RECT 16.0870 23.5035 16.1640 24.5970 ;
        RECT 14.1940 23.5035 14.2710 24.5970 ;
        RECT 14.0320 23.5035 14.0580 24.5970 ;
        RECT 13.9240 23.5035 13.9500 24.5970 ;
        RECT 13.8160 23.5035 13.8420 24.5970 ;
        RECT 13.7080 23.5035 13.7340 24.5970 ;
        RECT 13.6000 23.5035 13.6260 24.5970 ;
        RECT 13.4920 23.5035 13.5180 24.5970 ;
        RECT 13.3840 23.5035 13.4100 24.5970 ;
        RECT 13.2760 23.5035 13.3020 24.5970 ;
        RECT 13.1680 23.5035 13.1940 24.5970 ;
        RECT 13.0600 23.5035 13.0860 24.5970 ;
        RECT 12.9520 23.5035 12.9780 24.5970 ;
        RECT 12.8440 23.5035 12.8700 24.5970 ;
        RECT 12.7360 23.5035 12.7620 24.5970 ;
        RECT 12.6280 23.5035 12.6540 24.5970 ;
        RECT 12.5200 23.5035 12.5460 24.5970 ;
        RECT 12.4120 23.5035 12.4380 24.5970 ;
        RECT 12.3040 23.5035 12.3300 24.5970 ;
        RECT 12.1960 23.5035 12.2220 24.5970 ;
        RECT 12.0880 23.5035 12.1140 24.5970 ;
        RECT 11.9800 23.5035 12.0060 24.5970 ;
        RECT 11.8720 23.5035 11.8980 24.5970 ;
        RECT 11.7640 23.5035 11.7900 24.5970 ;
        RECT 11.6560 23.5035 11.6820 24.5970 ;
        RECT 11.5480 23.5035 11.5740 24.5970 ;
        RECT 11.4400 23.5035 11.4660 24.5970 ;
        RECT 11.3320 23.5035 11.3580 24.5970 ;
        RECT 11.2240 23.5035 11.2500 24.5970 ;
        RECT 11.1160 23.5035 11.1420 24.5970 ;
        RECT 11.0080 23.5035 11.0340 24.5970 ;
        RECT 10.9000 23.5035 10.9260 24.5970 ;
        RECT 10.7920 23.5035 10.8180 24.5970 ;
        RECT 10.6840 23.5035 10.7100 24.5970 ;
        RECT 10.5760 23.5035 10.6020 24.5970 ;
        RECT 10.4680 23.5035 10.4940 24.5970 ;
        RECT 10.3600 23.5035 10.3860 24.5970 ;
        RECT 10.2520 23.5035 10.2780 24.5970 ;
        RECT 10.1440 23.5035 10.1700 24.5970 ;
        RECT 10.0360 23.5035 10.0620 24.5970 ;
        RECT 9.9280 23.5035 9.9540 24.5970 ;
        RECT 9.8200 23.5035 9.8460 24.5970 ;
        RECT 9.7120 23.5035 9.7380 24.5970 ;
        RECT 9.6040 23.5035 9.6300 24.5970 ;
        RECT 9.4960 23.5035 9.5220 24.5970 ;
        RECT 9.3880 23.5035 9.4140 24.5970 ;
        RECT 9.2800 23.5035 9.3060 24.5970 ;
        RECT 9.1720 23.5035 9.1980 24.5970 ;
        RECT 9.0640 23.5035 9.0900 24.5970 ;
        RECT 8.9560 23.5035 8.9820 24.5970 ;
        RECT 8.8480 23.5035 8.8740 24.5970 ;
        RECT 8.7400 23.5035 8.7660 24.5970 ;
        RECT 8.6320 23.5035 8.6580 24.5970 ;
        RECT 8.5240 23.5035 8.5500 24.5970 ;
        RECT 8.4160 23.5035 8.4420 24.5970 ;
        RECT 8.3080 23.5035 8.3340 24.5970 ;
        RECT 8.2000 23.5035 8.2260 24.5970 ;
        RECT 8.0920 23.5035 8.1180 24.5970 ;
        RECT 7.9840 23.5035 8.0100 24.5970 ;
        RECT 7.8760 23.5035 7.9020 24.5970 ;
        RECT 7.7680 23.5035 7.7940 24.5970 ;
        RECT 7.6600 23.5035 7.6860 24.5970 ;
        RECT 7.5520 23.5035 7.5780 24.5970 ;
        RECT 7.4440 23.5035 7.4700 24.5970 ;
        RECT 7.3360 23.5035 7.3620 24.5970 ;
        RECT 7.2280 23.5035 7.2540 24.5970 ;
        RECT 7.1200 23.5035 7.1460 24.5970 ;
        RECT 7.0120 23.5035 7.0380 24.5970 ;
        RECT 6.9040 23.5035 6.9300 24.5970 ;
        RECT 6.7960 23.5035 6.8220 24.5970 ;
        RECT 6.6880 23.5035 6.7140 24.5970 ;
        RECT 6.5800 23.5035 6.6060 24.5970 ;
        RECT 6.4720 23.5035 6.4980 24.5970 ;
        RECT 6.3640 23.5035 6.3900 24.5970 ;
        RECT 6.2560 23.5035 6.2820 24.5970 ;
        RECT 6.1480 23.5035 6.1740 24.5970 ;
        RECT 6.0400 23.5035 6.0660 24.5970 ;
        RECT 5.9320 23.5035 5.9580 24.5970 ;
        RECT 5.8240 23.5035 5.8500 24.5970 ;
        RECT 5.7160 23.5035 5.7420 24.5970 ;
        RECT 5.6080 23.5035 5.6340 24.5970 ;
        RECT 5.5000 23.5035 5.5260 24.5970 ;
        RECT 5.3920 23.5035 5.4180 24.5970 ;
        RECT 5.2840 23.5035 5.3100 24.5970 ;
        RECT 5.1760 23.5035 5.2020 24.5970 ;
        RECT 5.0680 23.5035 5.0940 24.5970 ;
        RECT 4.9600 23.5035 4.9860 24.5970 ;
        RECT 4.8520 23.5035 4.8780 24.5970 ;
        RECT 4.7440 23.5035 4.7700 24.5970 ;
        RECT 4.6360 23.5035 4.6620 24.5970 ;
        RECT 4.5280 23.5035 4.5540 24.5970 ;
        RECT 4.4200 23.5035 4.4460 24.5970 ;
        RECT 4.3120 23.5035 4.3380 24.5970 ;
        RECT 4.2040 23.5035 4.2300 24.5970 ;
        RECT 4.0960 23.5035 4.1220 24.5970 ;
        RECT 3.9880 23.5035 4.0140 24.5970 ;
        RECT 3.8800 23.5035 3.9060 24.5970 ;
        RECT 3.7720 23.5035 3.7980 24.5970 ;
        RECT 3.6640 23.5035 3.6900 24.5970 ;
        RECT 3.5560 23.5035 3.5820 24.5970 ;
        RECT 3.4480 23.5035 3.4740 24.5970 ;
        RECT 3.3400 23.5035 3.3660 24.5970 ;
        RECT 3.2320 23.5035 3.2580 24.5970 ;
        RECT 3.1240 23.5035 3.1500 24.5970 ;
        RECT 3.0160 23.5035 3.0420 24.5970 ;
        RECT 2.9080 23.5035 2.9340 24.5970 ;
        RECT 2.8000 23.5035 2.8260 24.5970 ;
        RECT 2.6920 23.5035 2.7180 24.5970 ;
        RECT 2.5840 23.5035 2.6100 24.5970 ;
        RECT 2.4760 23.5035 2.5020 24.5970 ;
        RECT 2.3680 23.5035 2.3940 24.5970 ;
        RECT 2.2600 23.5035 2.2860 24.5970 ;
        RECT 2.1520 23.5035 2.1780 24.5970 ;
        RECT 2.0440 23.5035 2.0700 24.5970 ;
        RECT 1.9360 23.5035 1.9620 24.5970 ;
        RECT 1.8280 23.5035 1.8540 24.5970 ;
        RECT 1.7200 23.5035 1.7460 24.5970 ;
        RECT 1.6120 23.5035 1.6380 24.5970 ;
        RECT 1.5040 23.5035 1.5300 24.5970 ;
        RECT 1.3960 23.5035 1.4220 24.5970 ;
        RECT 1.2880 23.5035 1.3140 24.5970 ;
        RECT 1.1800 23.5035 1.2060 24.5970 ;
        RECT 1.0720 23.5035 1.0980 24.5970 ;
        RECT 0.9640 23.5035 0.9900 24.5970 ;
        RECT 0.8560 23.5035 0.8820 24.5970 ;
        RECT 0.7480 23.5035 0.7740 24.5970 ;
        RECT 0.6400 23.5035 0.6660 24.5970 ;
        RECT 0.5320 23.5035 0.5580 24.5970 ;
        RECT 0.4240 23.5035 0.4500 24.5970 ;
        RECT 0.3160 23.5035 0.3420 24.5970 ;
        RECT 0.2080 23.5035 0.2340 24.5970 ;
        RECT 0.0050 23.5035 0.0900 24.5970 ;
        RECT 15.5530 24.5835 15.6810 25.6770 ;
        RECT 15.5390 25.2490 15.6810 25.5715 ;
        RECT 15.3190 24.9760 15.4530 25.6770 ;
        RECT 15.2960 25.3110 15.4530 25.5690 ;
        RECT 15.3190 24.5835 15.4170 25.6770 ;
        RECT 15.3190 24.7045 15.4310 24.9440 ;
        RECT 15.3190 24.5835 15.4530 24.6725 ;
        RECT 15.0940 25.0340 15.2280 25.6770 ;
        RECT 15.0940 24.5835 15.1920 25.6770 ;
        RECT 14.6770 24.5835 14.7600 25.6770 ;
        RECT 14.6770 24.6720 14.7740 25.6075 ;
        RECT 30.2680 24.5835 30.3530 25.6770 ;
        RECT 30.1240 24.5835 30.1500 25.6770 ;
        RECT 30.0160 24.5835 30.0420 25.6770 ;
        RECT 29.9080 24.5835 29.9340 25.6770 ;
        RECT 29.8000 24.5835 29.8260 25.6770 ;
        RECT 29.6920 24.5835 29.7180 25.6770 ;
        RECT 29.5840 24.5835 29.6100 25.6770 ;
        RECT 29.4760 24.5835 29.5020 25.6770 ;
        RECT 29.3680 24.5835 29.3940 25.6770 ;
        RECT 29.2600 24.5835 29.2860 25.6770 ;
        RECT 29.1520 24.5835 29.1780 25.6770 ;
        RECT 29.0440 24.5835 29.0700 25.6770 ;
        RECT 28.9360 24.5835 28.9620 25.6770 ;
        RECT 28.8280 24.5835 28.8540 25.6770 ;
        RECT 28.7200 24.5835 28.7460 25.6770 ;
        RECT 28.6120 24.5835 28.6380 25.6770 ;
        RECT 28.5040 24.5835 28.5300 25.6770 ;
        RECT 28.3960 24.5835 28.4220 25.6770 ;
        RECT 28.2880 24.5835 28.3140 25.6770 ;
        RECT 28.1800 24.5835 28.2060 25.6770 ;
        RECT 28.0720 24.5835 28.0980 25.6770 ;
        RECT 27.9640 24.5835 27.9900 25.6770 ;
        RECT 27.8560 24.5835 27.8820 25.6770 ;
        RECT 27.7480 24.5835 27.7740 25.6770 ;
        RECT 27.6400 24.5835 27.6660 25.6770 ;
        RECT 27.5320 24.5835 27.5580 25.6770 ;
        RECT 27.4240 24.5835 27.4500 25.6770 ;
        RECT 27.3160 24.5835 27.3420 25.6770 ;
        RECT 27.2080 24.5835 27.2340 25.6770 ;
        RECT 27.1000 24.5835 27.1260 25.6770 ;
        RECT 26.9920 24.5835 27.0180 25.6770 ;
        RECT 26.8840 24.5835 26.9100 25.6770 ;
        RECT 26.7760 24.5835 26.8020 25.6770 ;
        RECT 26.6680 24.5835 26.6940 25.6770 ;
        RECT 26.5600 24.5835 26.5860 25.6770 ;
        RECT 26.4520 24.5835 26.4780 25.6770 ;
        RECT 26.3440 24.5835 26.3700 25.6770 ;
        RECT 26.2360 24.5835 26.2620 25.6770 ;
        RECT 26.1280 24.5835 26.1540 25.6770 ;
        RECT 26.0200 24.5835 26.0460 25.6770 ;
        RECT 25.9120 24.5835 25.9380 25.6770 ;
        RECT 25.8040 24.5835 25.8300 25.6770 ;
        RECT 25.6960 24.5835 25.7220 25.6770 ;
        RECT 25.5880 24.5835 25.6140 25.6770 ;
        RECT 25.4800 24.5835 25.5060 25.6770 ;
        RECT 25.3720 24.5835 25.3980 25.6770 ;
        RECT 25.2640 24.5835 25.2900 25.6770 ;
        RECT 25.1560 24.5835 25.1820 25.6770 ;
        RECT 25.0480 24.5835 25.0740 25.6770 ;
        RECT 24.9400 24.5835 24.9660 25.6770 ;
        RECT 24.8320 24.5835 24.8580 25.6770 ;
        RECT 24.7240 24.5835 24.7500 25.6770 ;
        RECT 24.6160 24.5835 24.6420 25.6770 ;
        RECT 24.5080 24.5835 24.5340 25.6770 ;
        RECT 24.4000 24.5835 24.4260 25.6770 ;
        RECT 24.2920 24.5835 24.3180 25.6770 ;
        RECT 24.1840 24.5835 24.2100 25.6770 ;
        RECT 24.0760 24.5835 24.1020 25.6770 ;
        RECT 23.9680 24.5835 23.9940 25.6770 ;
        RECT 23.8600 24.5835 23.8860 25.6770 ;
        RECT 23.7520 24.5835 23.7780 25.6770 ;
        RECT 23.6440 24.5835 23.6700 25.6770 ;
        RECT 23.5360 24.5835 23.5620 25.6770 ;
        RECT 23.4280 24.5835 23.4540 25.6770 ;
        RECT 23.3200 24.5835 23.3460 25.6770 ;
        RECT 23.2120 24.5835 23.2380 25.6770 ;
        RECT 23.1040 24.5835 23.1300 25.6770 ;
        RECT 22.9960 24.5835 23.0220 25.6770 ;
        RECT 22.8880 24.5835 22.9140 25.6770 ;
        RECT 22.7800 24.5835 22.8060 25.6770 ;
        RECT 22.6720 24.5835 22.6980 25.6770 ;
        RECT 22.5640 24.5835 22.5900 25.6770 ;
        RECT 22.4560 24.5835 22.4820 25.6770 ;
        RECT 22.3480 24.5835 22.3740 25.6770 ;
        RECT 22.2400 24.5835 22.2660 25.6770 ;
        RECT 22.1320 24.5835 22.1580 25.6770 ;
        RECT 22.0240 24.5835 22.0500 25.6770 ;
        RECT 21.9160 24.5835 21.9420 25.6770 ;
        RECT 21.8080 24.5835 21.8340 25.6770 ;
        RECT 21.7000 24.5835 21.7260 25.6770 ;
        RECT 21.5920 24.5835 21.6180 25.6770 ;
        RECT 21.4840 24.5835 21.5100 25.6770 ;
        RECT 21.3760 24.5835 21.4020 25.6770 ;
        RECT 21.2680 24.5835 21.2940 25.6770 ;
        RECT 21.1600 24.5835 21.1860 25.6770 ;
        RECT 21.0520 24.5835 21.0780 25.6770 ;
        RECT 20.9440 24.5835 20.9700 25.6770 ;
        RECT 20.8360 24.5835 20.8620 25.6770 ;
        RECT 20.7280 24.5835 20.7540 25.6770 ;
        RECT 20.6200 24.5835 20.6460 25.6770 ;
        RECT 20.5120 24.5835 20.5380 25.6770 ;
        RECT 20.4040 24.5835 20.4300 25.6770 ;
        RECT 20.2960 24.5835 20.3220 25.6770 ;
        RECT 20.1880 24.5835 20.2140 25.6770 ;
        RECT 20.0800 24.5835 20.1060 25.6770 ;
        RECT 19.9720 24.5835 19.9980 25.6770 ;
        RECT 19.8640 24.5835 19.8900 25.6770 ;
        RECT 19.7560 24.5835 19.7820 25.6770 ;
        RECT 19.6480 24.5835 19.6740 25.6770 ;
        RECT 19.5400 24.5835 19.5660 25.6770 ;
        RECT 19.4320 24.5835 19.4580 25.6770 ;
        RECT 19.3240 24.5835 19.3500 25.6770 ;
        RECT 19.2160 24.5835 19.2420 25.6770 ;
        RECT 19.1080 24.5835 19.1340 25.6770 ;
        RECT 19.0000 24.5835 19.0260 25.6770 ;
        RECT 18.8920 24.5835 18.9180 25.6770 ;
        RECT 18.7840 24.5835 18.8100 25.6770 ;
        RECT 18.6760 24.5835 18.7020 25.6770 ;
        RECT 18.5680 24.5835 18.5940 25.6770 ;
        RECT 18.4600 24.5835 18.4860 25.6770 ;
        RECT 18.3520 24.5835 18.3780 25.6770 ;
        RECT 18.2440 24.5835 18.2700 25.6770 ;
        RECT 18.1360 24.5835 18.1620 25.6770 ;
        RECT 18.0280 24.5835 18.0540 25.6770 ;
        RECT 17.9200 24.5835 17.9460 25.6770 ;
        RECT 17.8120 24.5835 17.8380 25.6770 ;
        RECT 17.7040 24.5835 17.7300 25.6770 ;
        RECT 17.5960 24.5835 17.6220 25.6770 ;
        RECT 17.4880 24.5835 17.5140 25.6770 ;
        RECT 17.3800 24.5835 17.4060 25.6770 ;
        RECT 17.2720 24.5835 17.2980 25.6770 ;
        RECT 17.1640 24.5835 17.1900 25.6770 ;
        RECT 17.0560 24.5835 17.0820 25.6770 ;
        RECT 16.9480 24.5835 16.9740 25.6770 ;
        RECT 16.8400 24.5835 16.8660 25.6770 ;
        RECT 16.7320 24.5835 16.7580 25.6770 ;
        RECT 16.6240 24.5835 16.6500 25.6770 ;
        RECT 16.5160 24.5835 16.5420 25.6770 ;
        RECT 16.4080 24.5835 16.4340 25.6770 ;
        RECT 16.3000 24.5835 16.3260 25.6770 ;
        RECT 16.0870 24.5835 16.1640 25.6770 ;
        RECT 14.1940 24.5835 14.2710 25.6770 ;
        RECT 14.0320 24.5835 14.0580 25.6770 ;
        RECT 13.9240 24.5835 13.9500 25.6770 ;
        RECT 13.8160 24.5835 13.8420 25.6770 ;
        RECT 13.7080 24.5835 13.7340 25.6770 ;
        RECT 13.6000 24.5835 13.6260 25.6770 ;
        RECT 13.4920 24.5835 13.5180 25.6770 ;
        RECT 13.3840 24.5835 13.4100 25.6770 ;
        RECT 13.2760 24.5835 13.3020 25.6770 ;
        RECT 13.1680 24.5835 13.1940 25.6770 ;
        RECT 13.0600 24.5835 13.0860 25.6770 ;
        RECT 12.9520 24.5835 12.9780 25.6770 ;
        RECT 12.8440 24.5835 12.8700 25.6770 ;
        RECT 12.7360 24.5835 12.7620 25.6770 ;
        RECT 12.6280 24.5835 12.6540 25.6770 ;
        RECT 12.5200 24.5835 12.5460 25.6770 ;
        RECT 12.4120 24.5835 12.4380 25.6770 ;
        RECT 12.3040 24.5835 12.3300 25.6770 ;
        RECT 12.1960 24.5835 12.2220 25.6770 ;
        RECT 12.0880 24.5835 12.1140 25.6770 ;
        RECT 11.9800 24.5835 12.0060 25.6770 ;
        RECT 11.8720 24.5835 11.8980 25.6770 ;
        RECT 11.7640 24.5835 11.7900 25.6770 ;
        RECT 11.6560 24.5835 11.6820 25.6770 ;
        RECT 11.5480 24.5835 11.5740 25.6770 ;
        RECT 11.4400 24.5835 11.4660 25.6770 ;
        RECT 11.3320 24.5835 11.3580 25.6770 ;
        RECT 11.2240 24.5835 11.2500 25.6770 ;
        RECT 11.1160 24.5835 11.1420 25.6770 ;
        RECT 11.0080 24.5835 11.0340 25.6770 ;
        RECT 10.9000 24.5835 10.9260 25.6770 ;
        RECT 10.7920 24.5835 10.8180 25.6770 ;
        RECT 10.6840 24.5835 10.7100 25.6770 ;
        RECT 10.5760 24.5835 10.6020 25.6770 ;
        RECT 10.4680 24.5835 10.4940 25.6770 ;
        RECT 10.3600 24.5835 10.3860 25.6770 ;
        RECT 10.2520 24.5835 10.2780 25.6770 ;
        RECT 10.1440 24.5835 10.1700 25.6770 ;
        RECT 10.0360 24.5835 10.0620 25.6770 ;
        RECT 9.9280 24.5835 9.9540 25.6770 ;
        RECT 9.8200 24.5835 9.8460 25.6770 ;
        RECT 9.7120 24.5835 9.7380 25.6770 ;
        RECT 9.6040 24.5835 9.6300 25.6770 ;
        RECT 9.4960 24.5835 9.5220 25.6770 ;
        RECT 9.3880 24.5835 9.4140 25.6770 ;
        RECT 9.2800 24.5835 9.3060 25.6770 ;
        RECT 9.1720 24.5835 9.1980 25.6770 ;
        RECT 9.0640 24.5835 9.0900 25.6770 ;
        RECT 8.9560 24.5835 8.9820 25.6770 ;
        RECT 8.8480 24.5835 8.8740 25.6770 ;
        RECT 8.7400 24.5835 8.7660 25.6770 ;
        RECT 8.6320 24.5835 8.6580 25.6770 ;
        RECT 8.5240 24.5835 8.5500 25.6770 ;
        RECT 8.4160 24.5835 8.4420 25.6770 ;
        RECT 8.3080 24.5835 8.3340 25.6770 ;
        RECT 8.2000 24.5835 8.2260 25.6770 ;
        RECT 8.0920 24.5835 8.1180 25.6770 ;
        RECT 7.9840 24.5835 8.0100 25.6770 ;
        RECT 7.8760 24.5835 7.9020 25.6770 ;
        RECT 7.7680 24.5835 7.7940 25.6770 ;
        RECT 7.6600 24.5835 7.6860 25.6770 ;
        RECT 7.5520 24.5835 7.5780 25.6770 ;
        RECT 7.4440 24.5835 7.4700 25.6770 ;
        RECT 7.3360 24.5835 7.3620 25.6770 ;
        RECT 7.2280 24.5835 7.2540 25.6770 ;
        RECT 7.1200 24.5835 7.1460 25.6770 ;
        RECT 7.0120 24.5835 7.0380 25.6770 ;
        RECT 6.9040 24.5835 6.9300 25.6770 ;
        RECT 6.7960 24.5835 6.8220 25.6770 ;
        RECT 6.6880 24.5835 6.7140 25.6770 ;
        RECT 6.5800 24.5835 6.6060 25.6770 ;
        RECT 6.4720 24.5835 6.4980 25.6770 ;
        RECT 6.3640 24.5835 6.3900 25.6770 ;
        RECT 6.2560 24.5835 6.2820 25.6770 ;
        RECT 6.1480 24.5835 6.1740 25.6770 ;
        RECT 6.0400 24.5835 6.0660 25.6770 ;
        RECT 5.9320 24.5835 5.9580 25.6770 ;
        RECT 5.8240 24.5835 5.8500 25.6770 ;
        RECT 5.7160 24.5835 5.7420 25.6770 ;
        RECT 5.6080 24.5835 5.6340 25.6770 ;
        RECT 5.5000 24.5835 5.5260 25.6770 ;
        RECT 5.3920 24.5835 5.4180 25.6770 ;
        RECT 5.2840 24.5835 5.3100 25.6770 ;
        RECT 5.1760 24.5835 5.2020 25.6770 ;
        RECT 5.0680 24.5835 5.0940 25.6770 ;
        RECT 4.9600 24.5835 4.9860 25.6770 ;
        RECT 4.8520 24.5835 4.8780 25.6770 ;
        RECT 4.7440 24.5835 4.7700 25.6770 ;
        RECT 4.6360 24.5835 4.6620 25.6770 ;
        RECT 4.5280 24.5835 4.5540 25.6770 ;
        RECT 4.4200 24.5835 4.4460 25.6770 ;
        RECT 4.3120 24.5835 4.3380 25.6770 ;
        RECT 4.2040 24.5835 4.2300 25.6770 ;
        RECT 4.0960 24.5835 4.1220 25.6770 ;
        RECT 3.9880 24.5835 4.0140 25.6770 ;
        RECT 3.8800 24.5835 3.9060 25.6770 ;
        RECT 3.7720 24.5835 3.7980 25.6770 ;
        RECT 3.6640 24.5835 3.6900 25.6770 ;
        RECT 3.5560 24.5835 3.5820 25.6770 ;
        RECT 3.4480 24.5835 3.4740 25.6770 ;
        RECT 3.3400 24.5835 3.3660 25.6770 ;
        RECT 3.2320 24.5835 3.2580 25.6770 ;
        RECT 3.1240 24.5835 3.1500 25.6770 ;
        RECT 3.0160 24.5835 3.0420 25.6770 ;
        RECT 2.9080 24.5835 2.9340 25.6770 ;
        RECT 2.8000 24.5835 2.8260 25.6770 ;
        RECT 2.6920 24.5835 2.7180 25.6770 ;
        RECT 2.5840 24.5835 2.6100 25.6770 ;
        RECT 2.4760 24.5835 2.5020 25.6770 ;
        RECT 2.3680 24.5835 2.3940 25.6770 ;
        RECT 2.2600 24.5835 2.2860 25.6770 ;
        RECT 2.1520 24.5835 2.1780 25.6770 ;
        RECT 2.0440 24.5835 2.0700 25.6770 ;
        RECT 1.9360 24.5835 1.9620 25.6770 ;
        RECT 1.8280 24.5835 1.8540 25.6770 ;
        RECT 1.7200 24.5835 1.7460 25.6770 ;
        RECT 1.6120 24.5835 1.6380 25.6770 ;
        RECT 1.5040 24.5835 1.5300 25.6770 ;
        RECT 1.3960 24.5835 1.4220 25.6770 ;
        RECT 1.2880 24.5835 1.3140 25.6770 ;
        RECT 1.1800 24.5835 1.2060 25.6770 ;
        RECT 1.0720 24.5835 1.0980 25.6770 ;
        RECT 0.9640 24.5835 0.9900 25.6770 ;
        RECT 0.8560 24.5835 0.8820 25.6770 ;
        RECT 0.7480 24.5835 0.7740 25.6770 ;
        RECT 0.6400 24.5835 0.6660 25.6770 ;
        RECT 0.5320 24.5835 0.5580 25.6770 ;
        RECT 0.4240 24.5835 0.4500 25.6770 ;
        RECT 0.3160 24.5835 0.3420 25.6770 ;
        RECT 0.2080 24.5835 0.2340 25.6770 ;
        RECT 0.0050 24.5835 0.0900 25.6770 ;
        RECT 15.5530 25.6635 15.6810 26.7570 ;
        RECT 15.5390 26.3290 15.6810 26.6515 ;
        RECT 15.3190 26.0560 15.4530 26.7570 ;
        RECT 15.2960 26.3910 15.4530 26.6490 ;
        RECT 15.3190 25.6635 15.4170 26.7570 ;
        RECT 15.3190 25.7845 15.4310 26.0240 ;
        RECT 15.3190 25.6635 15.4530 25.7525 ;
        RECT 15.0940 26.1140 15.2280 26.7570 ;
        RECT 15.0940 25.6635 15.1920 26.7570 ;
        RECT 14.6770 25.6635 14.7600 26.7570 ;
        RECT 14.6770 25.7520 14.7740 26.6875 ;
        RECT 30.2680 25.6635 30.3530 26.7570 ;
        RECT 30.1240 25.6635 30.1500 26.7570 ;
        RECT 30.0160 25.6635 30.0420 26.7570 ;
        RECT 29.9080 25.6635 29.9340 26.7570 ;
        RECT 29.8000 25.6635 29.8260 26.7570 ;
        RECT 29.6920 25.6635 29.7180 26.7570 ;
        RECT 29.5840 25.6635 29.6100 26.7570 ;
        RECT 29.4760 25.6635 29.5020 26.7570 ;
        RECT 29.3680 25.6635 29.3940 26.7570 ;
        RECT 29.2600 25.6635 29.2860 26.7570 ;
        RECT 29.1520 25.6635 29.1780 26.7570 ;
        RECT 29.0440 25.6635 29.0700 26.7570 ;
        RECT 28.9360 25.6635 28.9620 26.7570 ;
        RECT 28.8280 25.6635 28.8540 26.7570 ;
        RECT 28.7200 25.6635 28.7460 26.7570 ;
        RECT 28.6120 25.6635 28.6380 26.7570 ;
        RECT 28.5040 25.6635 28.5300 26.7570 ;
        RECT 28.3960 25.6635 28.4220 26.7570 ;
        RECT 28.2880 25.6635 28.3140 26.7570 ;
        RECT 28.1800 25.6635 28.2060 26.7570 ;
        RECT 28.0720 25.6635 28.0980 26.7570 ;
        RECT 27.9640 25.6635 27.9900 26.7570 ;
        RECT 27.8560 25.6635 27.8820 26.7570 ;
        RECT 27.7480 25.6635 27.7740 26.7570 ;
        RECT 27.6400 25.6635 27.6660 26.7570 ;
        RECT 27.5320 25.6635 27.5580 26.7570 ;
        RECT 27.4240 25.6635 27.4500 26.7570 ;
        RECT 27.3160 25.6635 27.3420 26.7570 ;
        RECT 27.2080 25.6635 27.2340 26.7570 ;
        RECT 27.1000 25.6635 27.1260 26.7570 ;
        RECT 26.9920 25.6635 27.0180 26.7570 ;
        RECT 26.8840 25.6635 26.9100 26.7570 ;
        RECT 26.7760 25.6635 26.8020 26.7570 ;
        RECT 26.6680 25.6635 26.6940 26.7570 ;
        RECT 26.5600 25.6635 26.5860 26.7570 ;
        RECT 26.4520 25.6635 26.4780 26.7570 ;
        RECT 26.3440 25.6635 26.3700 26.7570 ;
        RECT 26.2360 25.6635 26.2620 26.7570 ;
        RECT 26.1280 25.6635 26.1540 26.7570 ;
        RECT 26.0200 25.6635 26.0460 26.7570 ;
        RECT 25.9120 25.6635 25.9380 26.7570 ;
        RECT 25.8040 25.6635 25.8300 26.7570 ;
        RECT 25.6960 25.6635 25.7220 26.7570 ;
        RECT 25.5880 25.6635 25.6140 26.7570 ;
        RECT 25.4800 25.6635 25.5060 26.7570 ;
        RECT 25.3720 25.6635 25.3980 26.7570 ;
        RECT 25.2640 25.6635 25.2900 26.7570 ;
        RECT 25.1560 25.6635 25.1820 26.7570 ;
        RECT 25.0480 25.6635 25.0740 26.7570 ;
        RECT 24.9400 25.6635 24.9660 26.7570 ;
        RECT 24.8320 25.6635 24.8580 26.7570 ;
        RECT 24.7240 25.6635 24.7500 26.7570 ;
        RECT 24.6160 25.6635 24.6420 26.7570 ;
        RECT 24.5080 25.6635 24.5340 26.7570 ;
        RECT 24.4000 25.6635 24.4260 26.7570 ;
        RECT 24.2920 25.6635 24.3180 26.7570 ;
        RECT 24.1840 25.6635 24.2100 26.7570 ;
        RECT 24.0760 25.6635 24.1020 26.7570 ;
        RECT 23.9680 25.6635 23.9940 26.7570 ;
        RECT 23.8600 25.6635 23.8860 26.7570 ;
        RECT 23.7520 25.6635 23.7780 26.7570 ;
        RECT 23.6440 25.6635 23.6700 26.7570 ;
        RECT 23.5360 25.6635 23.5620 26.7570 ;
        RECT 23.4280 25.6635 23.4540 26.7570 ;
        RECT 23.3200 25.6635 23.3460 26.7570 ;
        RECT 23.2120 25.6635 23.2380 26.7570 ;
        RECT 23.1040 25.6635 23.1300 26.7570 ;
        RECT 22.9960 25.6635 23.0220 26.7570 ;
        RECT 22.8880 25.6635 22.9140 26.7570 ;
        RECT 22.7800 25.6635 22.8060 26.7570 ;
        RECT 22.6720 25.6635 22.6980 26.7570 ;
        RECT 22.5640 25.6635 22.5900 26.7570 ;
        RECT 22.4560 25.6635 22.4820 26.7570 ;
        RECT 22.3480 25.6635 22.3740 26.7570 ;
        RECT 22.2400 25.6635 22.2660 26.7570 ;
        RECT 22.1320 25.6635 22.1580 26.7570 ;
        RECT 22.0240 25.6635 22.0500 26.7570 ;
        RECT 21.9160 25.6635 21.9420 26.7570 ;
        RECT 21.8080 25.6635 21.8340 26.7570 ;
        RECT 21.7000 25.6635 21.7260 26.7570 ;
        RECT 21.5920 25.6635 21.6180 26.7570 ;
        RECT 21.4840 25.6635 21.5100 26.7570 ;
        RECT 21.3760 25.6635 21.4020 26.7570 ;
        RECT 21.2680 25.6635 21.2940 26.7570 ;
        RECT 21.1600 25.6635 21.1860 26.7570 ;
        RECT 21.0520 25.6635 21.0780 26.7570 ;
        RECT 20.9440 25.6635 20.9700 26.7570 ;
        RECT 20.8360 25.6635 20.8620 26.7570 ;
        RECT 20.7280 25.6635 20.7540 26.7570 ;
        RECT 20.6200 25.6635 20.6460 26.7570 ;
        RECT 20.5120 25.6635 20.5380 26.7570 ;
        RECT 20.4040 25.6635 20.4300 26.7570 ;
        RECT 20.2960 25.6635 20.3220 26.7570 ;
        RECT 20.1880 25.6635 20.2140 26.7570 ;
        RECT 20.0800 25.6635 20.1060 26.7570 ;
        RECT 19.9720 25.6635 19.9980 26.7570 ;
        RECT 19.8640 25.6635 19.8900 26.7570 ;
        RECT 19.7560 25.6635 19.7820 26.7570 ;
        RECT 19.6480 25.6635 19.6740 26.7570 ;
        RECT 19.5400 25.6635 19.5660 26.7570 ;
        RECT 19.4320 25.6635 19.4580 26.7570 ;
        RECT 19.3240 25.6635 19.3500 26.7570 ;
        RECT 19.2160 25.6635 19.2420 26.7570 ;
        RECT 19.1080 25.6635 19.1340 26.7570 ;
        RECT 19.0000 25.6635 19.0260 26.7570 ;
        RECT 18.8920 25.6635 18.9180 26.7570 ;
        RECT 18.7840 25.6635 18.8100 26.7570 ;
        RECT 18.6760 25.6635 18.7020 26.7570 ;
        RECT 18.5680 25.6635 18.5940 26.7570 ;
        RECT 18.4600 25.6635 18.4860 26.7570 ;
        RECT 18.3520 25.6635 18.3780 26.7570 ;
        RECT 18.2440 25.6635 18.2700 26.7570 ;
        RECT 18.1360 25.6635 18.1620 26.7570 ;
        RECT 18.0280 25.6635 18.0540 26.7570 ;
        RECT 17.9200 25.6635 17.9460 26.7570 ;
        RECT 17.8120 25.6635 17.8380 26.7570 ;
        RECT 17.7040 25.6635 17.7300 26.7570 ;
        RECT 17.5960 25.6635 17.6220 26.7570 ;
        RECT 17.4880 25.6635 17.5140 26.7570 ;
        RECT 17.3800 25.6635 17.4060 26.7570 ;
        RECT 17.2720 25.6635 17.2980 26.7570 ;
        RECT 17.1640 25.6635 17.1900 26.7570 ;
        RECT 17.0560 25.6635 17.0820 26.7570 ;
        RECT 16.9480 25.6635 16.9740 26.7570 ;
        RECT 16.8400 25.6635 16.8660 26.7570 ;
        RECT 16.7320 25.6635 16.7580 26.7570 ;
        RECT 16.6240 25.6635 16.6500 26.7570 ;
        RECT 16.5160 25.6635 16.5420 26.7570 ;
        RECT 16.4080 25.6635 16.4340 26.7570 ;
        RECT 16.3000 25.6635 16.3260 26.7570 ;
        RECT 16.0870 25.6635 16.1640 26.7570 ;
        RECT 14.1940 25.6635 14.2710 26.7570 ;
        RECT 14.0320 25.6635 14.0580 26.7570 ;
        RECT 13.9240 25.6635 13.9500 26.7570 ;
        RECT 13.8160 25.6635 13.8420 26.7570 ;
        RECT 13.7080 25.6635 13.7340 26.7570 ;
        RECT 13.6000 25.6635 13.6260 26.7570 ;
        RECT 13.4920 25.6635 13.5180 26.7570 ;
        RECT 13.3840 25.6635 13.4100 26.7570 ;
        RECT 13.2760 25.6635 13.3020 26.7570 ;
        RECT 13.1680 25.6635 13.1940 26.7570 ;
        RECT 13.0600 25.6635 13.0860 26.7570 ;
        RECT 12.9520 25.6635 12.9780 26.7570 ;
        RECT 12.8440 25.6635 12.8700 26.7570 ;
        RECT 12.7360 25.6635 12.7620 26.7570 ;
        RECT 12.6280 25.6635 12.6540 26.7570 ;
        RECT 12.5200 25.6635 12.5460 26.7570 ;
        RECT 12.4120 25.6635 12.4380 26.7570 ;
        RECT 12.3040 25.6635 12.3300 26.7570 ;
        RECT 12.1960 25.6635 12.2220 26.7570 ;
        RECT 12.0880 25.6635 12.1140 26.7570 ;
        RECT 11.9800 25.6635 12.0060 26.7570 ;
        RECT 11.8720 25.6635 11.8980 26.7570 ;
        RECT 11.7640 25.6635 11.7900 26.7570 ;
        RECT 11.6560 25.6635 11.6820 26.7570 ;
        RECT 11.5480 25.6635 11.5740 26.7570 ;
        RECT 11.4400 25.6635 11.4660 26.7570 ;
        RECT 11.3320 25.6635 11.3580 26.7570 ;
        RECT 11.2240 25.6635 11.2500 26.7570 ;
        RECT 11.1160 25.6635 11.1420 26.7570 ;
        RECT 11.0080 25.6635 11.0340 26.7570 ;
        RECT 10.9000 25.6635 10.9260 26.7570 ;
        RECT 10.7920 25.6635 10.8180 26.7570 ;
        RECT 10.6840 25.6635 10.7100 26.7570 ;
        RECT 10.5760 25.6635 10.6020 26.7570 ;
        RECT 10.4680 25.6635 10.4940 26.7570 ;
        RECT 10.3600 25.6635 10.3860 26.7570 ;
        RECT 10.2520 25.6635 10.2780 26.7570 ;
        RECT 10.1440 25.6635 10.1700 26.7570 ;
        RECT 10.0360 25.6635 10.0620 26.7570 ;
        RECT 9.9280 25.6635 9.9540 26.7570 ;
        RECT 9.8200 25.6635 9.8460 26.7570 ;
        RECT 9.7120 25.6635 9.7380 26.7570 ;
        RECT 9.6040 25.6635 9.6300 26.7570 ;
        RECT 9.4960 25.6635 9.5220 26.7570 ;
        RECT 9.3880 25.6635 9.4140 26.7570 ;
        RECT 9.2800 25.6635 9.3060 26.7570 ;
        RECT 9.1720 25.6635 9.1980 26.7570 ;
        RECT 9.0640 25.6635 9.0900 26.7570 ;
        RECT 8.9560 25.6635 8.9820 26.7570 ;
        RECT 8.8480 25.6635 8.8740 26.7570 ;
        RECT 8.7400 25.6635 8.7660 26.7570 ;
        RECT 8.6320 25.6635 8.6580 26.7570 ;
        RECT 8.5240 25.6635 8.5500 26.7570 ;
        RECT 8.4160 25.6635 8.4420 26.7570 ;
        RECT 8.3080 25.6635 8.3340 26.7570 ;
        RECT 8.2000 25.6635 8.2260 26.7570 ;
        RECT 8.0920 25.6635 8.1180 26.7570 ;
        RECT 7.9840 25.6635 8.0100 26.7570 ;
        RECT 7.8760 25.6635 7.9020 26.7570 ;
        RECT 7.7680 25.6635 7.7940 26.7570 ;
        RECT 7.6600 25.6635 7.6860 26.7570 ;
        RECT 7.5520 25.6635 7.5780 26.7570 ;
        RECT 7.4440 25.6635 7.4700 26.7570 ;
        RECT 7.3360 25.6635 7.3620 26.7570 ;
        RECT 7.2280 25.6635 7.2540 26.7570 ;
        RECT 7.1200 25.6635 7.1460 26.7570 ;
        RECT 7.0120 25.6635 7.0380 26.7570 ;
        RECT 6.9040 25.6635 6.9300 26.7570 ;
        RECT 6.7960 25.6635 6.8220 26.7570 ;
        RECT 6.6880 25.6635 6.7140 26.7570 ;
        RECT 6.5800 25.6635 6.6060 26.7570 ;
        RECT 6.4720 25.6635 6.4980 26.7570 ;
        RECT 6.3640 25.6635 6.3900 26.7570 ;
        RECT 6.2560 25.6635 6.2820 26.7570 ;
        RECT 6.1480 25.6635 6.1740 26.7570 ;
        RECT 6.0400 25.6635 6.0660 26.7570 ;
        RECT 5.9320 25.6635 5.9580 26.7570 ;
        RECT 5.8240 25.6635 5.8500 26.7570 ;
        RECT 5.7160 25.6635 5.7420 26.7570 ;
        RECT 5.6080 25.6635 5.6340 26.7570 ;
        RECT 5.5000 25.6635 5.5260 26.7570 ;
        RECT 5.3920 25.6635 5.4180 26.7570 ;
        RECT 5.2840 25.6635 5.3100 26.7570 ;
        RECT 5.1760 25.6635 5.2020 26.7570 ;
        RECT 5.0680 25.6635 5.0940 26.7570 ;
        RECT 4.9600 25.6635 4.9860 26.7570 ;
        RECT 4.8520 25.6635 4.8780 26.7570 ;
        RECT 4.7440 25.6635 4.7700 26.7570 ;
        RECT 4.6360 25.6635 4.6620 26.7570 ;
        RECT 4.5280 25.6635 4.5540 26.7570 ;
        RECT 4.4200 25.6635 4.4460 26.7570 ;
        RECT 4.3120 25.6635 4.3380 26.7570 ;
        RECT 4.2040 25.6635 4.2300 26.7570 ;
        RECT 4.0960 25.6635 4.1220 26.7570 ;
        RECT 3.9880 25.6635 4.0140 26.7570 ;
        RECT 3.8800 25.6635 3.9060 26.7570 ;
        RECT 3.7720 25.6635 3.7980 26.7570 ;
        RECT 3.6640 25.6635 3.6900 26.7570 ;
        RECT 3.5560 25.6635 3.5820 26.7570 ;
        RECT 3.4480 25.6635 3.4740 26.7570 ;
        RECT 3.3400 25.6635 3.3660 26.7570 ;
        RECT 3.2320 25.6635 3.2580 26.7570 ;
        RECT 3.1240 25.6635 3.1500 26.7570 ;
        RECT 3.0160 25.6635 3.0420 26.7570 ;
        RECT 2.9080 25.6635 2.9340 26.7570 ;
        RECT 2.8000 25.6635 2.8260 26.7570 ;
        RECT 2.6920 25.6635 2.7180 26.7570 ;
        RECT 2.5840 25.6635 2.6100 26.7570 ;
        RECT 2.4760 25.6635 2.5020 26.7570 ;
        RECT 2.3680 25.6635 2.3940 26.7570 ;
        RECT 2.2600 25.6635 2.2860 26.7570 ;
        RECT 2.1520 25.6635 2.1780 26.7570 ;
        RECT 2.0440 25.6635 2.0700 26.7570 ;
        RECT 1.9360 25.6635 1.9620 26.7570 ;
        RECT 1.8280 25.6635 1.8540 26.7570 ;
        RECT 1.7200 25.6635 1.7460 26.7570 ;
        RECT 1.6120 25.6635 1.6380 26.7570 ;
        RECT 1.5040 25.6635 1.5300 26.7570 ;
        RECT 1.3960 25.6635 1.4220 26.7570 ;
        RECT 1.2880 25.6635 1.3140 26.7570 ;
        RECT 1.1800 25.6635 1.2060 26.7570 ;
        RECT 1.0720 25.6635 1.0980 26.7570 ;
        RECT 0.9640 25.6635 0.9900 26.7570 ;
        RECT 0.8560 25.6635 0.8820 26.7570 ;
        RECT 0.7480 25.6635 0.7740 26.7570 ;
        RECT 0.6400 25.6635 0.6660 26.7570 ;
        RECT 0.5320 25.6635 0.5580 26.7570 ;
        RECT 0.4240 25.6635 0.4500 26.7570 ;
        RECT 0.3160 25.6635 0.3420 26.7570 ;
        RECT 0.2080 25.6635 0.2340 26.7570 ;
        RECT 0.0050 25.6635 0.0900 26.7570 ;
        RECT 15.5530 26.7435 15.6810 27.8370 ;
        RECT 15.5390 27.4090 15.6810 27.7315 ;
        RECT 15.3190 27.1360 15.4530 27.8370 ;
        RECT 15.2960 27.4710 15.4530 27.7290 ;
        RECT 15.3190 26.7435 15.4170 27.8370 ;
        RECT 15.3190 26.8645 15.4310 27.1040 ;
        RECT 15.3190 26.7435 15.4530 26.8325 ;
        RECT 15.0940 27.1940 15.2280 27.8370 ;
        RECT 15.0940 26.7435 15.1920 27.8370 ;
        RECT 14.6770 26.7435 14.7600 27.8370 ;
        RECT 14.6770 26.8320 14.7740 27.7675 ;
        RECT 30.2680 26.7435 30.3530 27.8370 ;
        RECT 30.1240 26.7435 30.1500 27.8370 ;
        RECT 30.0160 26.7435 30.0420 27.8370 ;
        RECT 29.9080 26.7435 29.9340 27.8370 ;
        RECT 29.8000 26.7435 29.8260 27.8370 ;
        RECT 29.6920 26.7435 29.7180 27.8370 ;
        RECT 29.5840 26.7435 29.6100 27.8370 ;
        RECT 29.4760 26.7435 29.5020 27.8370 ;
        RECT 29.3680 26.7435 29.3940 27.8370 ;
        RECT 29.2600 26.7435 29.2860 27.8370 ;
        RECT 29.1520 26.7435 29.1780 27.8370 ;
        RECT 29.0440 26.7435 29.0700 27.8370 ;
        RECT 28.9360 26.7435 28.9620 27.8370 ;
        RECT 28.8280 26.7435 28.8540 27.8370 ;
        RECT 28.7200 26.7435 28.7460 27.8370 ;
        RECT 28.6120 26.7435 28.6380 27.8370 ;
        RECT 28.5040 26.7435 28.5300 27.8370 ;
        RECT 28.3960 26.7435 28.4220 27.8370 ;
        RECT 28.2880 26.7435 28.3140 27.8370 ;
        RECT 28.1800 26.7435 28.2060 27.8370 ;
        RECT 28.0720 26.7435 28.0980 27.8370 ;
        RECT 27.9640 26.7435 27.9900 27.8370 ;
        RECT 27.8560 26.7435 27.8820 27.8370 ;
        RECT 27.7480 26.7435 27.7740 27.8370 ;
        RECT 27.6400 26.7435 27.6660 27.8370 ;
        RECT 27.5320 26.7435 27.5580 27.8370 ;
        RECT 27.4240 26.7435 27.4500 27.8370 ;
        RECT 27.3160 26.7435 27.3420 27.8370 ;
        RECT 27.2080 26.7435 27.2340 27.8370 ;
        RECT 27.1000 26.7435 27.1260 27.8370 ;
        RECT 26.9920 26.7435 27.0180 27.8370 ;
        RECT 26.8840 26.7435 26.9100 27.8370 ;
        RECT 26.7760 26.7435 26.8020 27.8370 ;
        RECT 26.6680 26.7435 26.6940 27.8370 ;
        RECT 26.5600 26.7435 26.5860 27.8370 ;
        RECT 26.4520 26.7435 26.4780 27.8370 ;
        RECT 26.3440 26.7435 26.3700 27.8370 ;
        RECT 26.2360 26.7435 26.2620 27.8370 ;
        RECT 26.1280 26.7435 26.1540 27.8370 ;
        RECT 26.0200 26.7435 26.0460 27.8370 ;
        RECT 25.9120 26.7435 25.9380 27.8370 ;
        RECT 25.8040 26.7435 25.8300 27.8370 ;
        RECT 25.6960 26.7435 25.7220 27.8370 ;
        RECT 25.5880 26.7435 25.6140 27.8370 ;
        RECT 25.4800 26.7435 25.5060 27.8370 ;
        RECT 25.3720 26.7435 25.3980 27.8370 ;
        RECT 25.2640 26.7435 25.2900 27.8370 ;
        RECT 25.1560 26.7435 25.1820 27.8370 ;
        RECT 25.0480 26.7435 25.0740 27.8370 ;
        RECT 24.9400 26.7435 24.9660 27.8370 ;
        RECT 24.8320 26.7435 24.8580 27.8370 ;
        RECT 24.7240 26.7435 24.7500 27.8370 ;
        RECT 24.6160 26.7435 24.6420 27.8370 ;
        RECT 24.5080 26.7435 24.5340 27.8370 ;
        RECT 24.4000 26.7435 24.4260 27.8370 ;
        RECT 24.2920 26.7435 24.3180 27.8370 ;
        RECT 24.1840 26.7435 24.2100 27.8370 ;
        RECT 24.0760 26.7435 24.1020 27.8370 ;
        RECT 23.9680 26.7435 23.9940 27.8370 ;
        RECT 23.8600 26.7435 23.8860 27.8370 ;
        RECT 23.7520 26.7435 23.7780 27.8370 ;
        RECT 23.6440 26.7435 23.6700 27.8370 ;
        RECT 23.5360 26.7435 23.5620 27.8370 ;
        RECT 23.4280 26.7435 23.4540 27.8370 ;
        RECT 23.3200 26.7435 23.3460 27.8370 ;
        RECT 23.2120 26.7435 23.2380 27.8370 ;
        RECT 23.1040 26.7435 23.1300 27.8370 ;
        RECT 22.9960 26.7435 23.0220 27.8370 ;
        RECT 22.8880 26.7435 22.9140 27.8370 ;
        RECT 22.7800 26.7435 22.8060 27.8370 ;
        RECT 22.6720 26.7435 22.6980 27.8370 ;
        RECT 22.5640 26.7435 22.5900 27.8370 ;
        RECT 22.4560 26.7435 22.4820 27.8370 ;
        RECT 22.3480 26.7435 22.3740 27.8370 ;
        RECT 22.2400 26.7435 22.2660 27.8370 ;
        RECT 22.1320 26.7435 22.1580 27.8370 ;
        RECT 22.0240 26.7435 22.0500 27.8370 ;
        RECT 21.9160 26.7435 21.9420 27.8370 ;
        RECT 21.8080 26.7435 21.8340 27.8370 ;
        RECT 21.7000 26.7435 21.7260 27.8370 ;
        RECT 21.5920 26.7435 21.6180 27.8370 ;
        RECT 21.4840 26.7435 21.5100 27.8370 ;
        RECT 21.3760 26.7435 21.4020 27.8370 ;
        RECT 21.2680 26.7435 21.2940 27.8370 ;
        RECT 21.1600 26.7435 21.1860 27.8370 ;
        RECT 21.0520 26.7435 21.0780 27.8370 ;
        RECT 20.9440 26.7435 20.9700 27.8370 ;
        RECT 20.8360 26.7435 20.8620 27.8370 ;
        RECT 20.7280 26.7435 20.7540 27.8370 ;
        RECT 20.6200 26.7435 20.6460 27.8370 ;
        RECT 20.5120 26.7435 20.5380 27.8370 ;
        RECT 20.4040 26.7435 20.4300 27.8370 ;
        RECT 20.2960 26.7435 20.3220 27.8370 ;
        RECT 20.1880 26.7435 20.2140 27.8370 ;
        RECT 20.0800 26.7435 20.1060 27.8370 ;
        RECT 19.9720 26.7435 19.9980 27.8370 ;
        RECT 19.8640 26.7435 19.8900 27.8370 ;
        RECT 19.7560 26.7435 19.7820 27.8370 ;
        RECT 19.6480 26.7435 19.6740 27.8370 ;
        RECT 19.5400 26.7435 19.5660 27.8370 ;
        RECT 19.4320 26.7435 19.4580 27.8370 ;
        RECT 19.3240 26.7435 19.3500 27.8370 ;
        RECT 19.2160 26.7435 19.2420 27.8370 ;
        RECT 19.1080 26.7435 19.1340 27.8370 ;
        RECT 19.0000 26.7435 19.0260 27.8370 ;
        RECT 18.8920 26.7435 18.9180 27.8370 ;
        RECT 18.7840 26.7435 18.8100 27.8370 ;
        RECT 18.6760 26.7435 18.7020 27.8370 ;
        RECT 18.5680 26.7435 18.5940 27.8370 ;
        RECT 18.4600 26.7435 18.4860 27.8370 ;
        RECT 18.3520 26.7435 18.3780 27.8370 ;
        RECT 18.2440 26.7435 18.2700 27.8370 ;
        RECT 18.1360 26.7435 18.1620 27.8370 ;
        RECT 18.0280 26.7435 18.0540 27.8370 ;
        RECT 17.9200 26.7435 17.9460 27.8370 ;
        RECT 17.8120 26.7435 17.8380 27.8370 ;
        RECT 17.7040 26.7435 17.7300 27.8370 ;
        RECT 17.5960 26.7435 17.6220 27.8370 ;
        RECT 17.4880 26.7435 17.5140 27.8370 ;
        RECT 17.3800 26.7435 17.4060 27.8370 ;
        RECT 17.2720 26.7435 17.2980 27.8370 ;
        RECT 17.1640 26.7435 17.1900 27.8370 ;
        RECT 17.0560 26.7435 17.0820 27.8370 ;
        RECT 16.9480 26.7435 16.9740 27.8370 ;
        RECT 16.8400 26.7435 16.8660 27.8370 ;
        RECT 16.7320 26.7435 16.7580 27.8370 ;
        RECT 16.6240 26.7435 16.6500 27.8370 ;
        RECT 16.5160 26.7435 16.5420 27.8370 ;
        RECT 16.4080 26.7435 16.4340 27.8370 ;
        RECT 16.3000 26.7435 16.3260 27.8370 ;
        RECT 16.0870 26.7435 16.1640 27.8370 ;
        RECT 14.1940 26.7435 14.2710 27.8370 ;
        RECT 14.0320 26.7435 14.0580 27.8370 ;
        RECT 13.9240 26.7435 13.9500 27.8370 ;
        RECT 13.8160 26.7435 13.8420 27.8370 ;
        RECT 13.7080 26.7435 13.7340 27.8370 ;
        RECT 13.6000 26.7435 13.6260 27.8370 ;
        RECT 13.4920 26.7435 13.5180 27.8370 ;
        RECT 13.3840 26.7435 13.4100 27.8370 ;
        RECT 13.2760 26.7435 13.3020 27.8370 ;
        RECT 13.1680 26.7435 13.1940 27.8370 ;
        RECT 13.0600 26.7435 13.0860 27.8370 ;
        RECT 12.9520 26.7435 12.9780 27.8370 ;
        RECT 12.8440 26.7435 12.8700 27.8370 ;
        RECT 12.7360 26.7435 12.7620 27.8370 ;
        RECT 12.6280 26.7435 12.6540 27.8370 ;
        RECT 12.5200 26.7435 12.5460 27.8370 ;
        RECT 12.4120 26.7435 12.4380 27.8370 ;
        RECT 12.3040 26.7435 12.3300 27.8370 ;
        RECT 12.1960 26.7435 12.2220 27.8370 ;
        RECT 12.0880 26.7435 12.1140 27.8370 ;
        RECT 11.9800 26.7435 12.0060 27.8370 ;
        RECT 11.8720 26.7435 11.8980 27.8370 ;
        RECT 11.7640 26.7435 11.7900 27.8370 ;
        RECT 11.6560 26.7435 11.6820 27.8370 ;
        RECT 11.5480 26.7435 11.5740 27.8370 ;
        RECT 11.4400 26.7435 11.4660 27.8370 ;
        RECT 11.3320 26.7435 11.3580 27.8370 ;
        RECT 11.2240 26.7435 11.2500 27.8370 ;
        RECT 11.1160 26.7435 11.1420 27.8370 ;
        RECT 11.0080 26.7435 11.0340 27.8370 ;
        RECT 10.9000 26.7435 10.9260 27.8370 ;
        RECT 10.7920 26.7435 10.8180 27.8370 ;
        RECT 10.6840 26.7435 10.7100 27.8370 ;
        RECT 10.5760 26.7435 10.6020 27.8370 ;
        RECT 10.4680 26.7435 10.4940 27.8370 ;
        RECT 10.3600 26.7435 10.3860 27.8370 ;
        RECT 10.2520 26.7435 10.2780 27.8370 ;
        RECT 10.1440 26.7435 10.1700 27.8370 ;
        RECT 10.0360 26.7435 10.0620 27.8370 ;
        RECT 9.9280 26.7435 9.9540 27.8370 ;
        RECT 9.8200 26.7435 9.8460 27.8370 ;
        RECT 9.7120 26.7435 9.7380 27.8370 ;
        RECT 9.6040 26.7435 9.6300 27.8370 ;
        RECT 9.4960 26.7435 9.5220 27.8370 ;
        RECT 9.3880 26.7435 9.4140 27.8370 ;
        RECT 9.2800 26.7435 9.3060 27.8370 ;
        RECT 9.1720 26.7435 9.1980 27.8370 ;
        RECT 9.0640 26.7435 9.0900 27.8370 ;
        RECT 8.9560 26.7435 8.9820 27.8370 ;
        RECT 8.8480 26.7435 8.8740 27.8370 ;
        RECT 8.7400 26.7435 8.7660 27.8370 ;
        RECT 8.6320 26.7435 8.6580 27.8370 ;
        RECT 8.5240 26.7435 8.5500 27.8370 ;
        RECT 8.4160 26.7435 8.4420 27.8370 ;
        RECT 8.3080 26.7435 8.3340 27.8370 ;
        RECT 8.2000 26.7435 8.2260 27.8370 ;
        RECT 8.0920 26.7435 8.1180 27.8370 ;
        RECT 7.9840 26.7435 8.0100 27.8370 ;
        RECT 7.8760 26.7435 7.9020 27.8370 ;
        RECT 7.7680 26.7435 7.7940 27.8370 ;
        RECT 7.6600 26.7435 7.6860 27.8370 ;
        RECT 7.5520 26.7435 7.5780 27.8370 ;
        RECT 7.4440 26.7435 7.4700 27.8370 ;
        RECT 7.3360 26.7435 7.3620 27.8370 ;
        RECT 7.2280 26.7435 7.2540 27.8370 ;
        RECT 7.1200 26.7435 7.1460 27.8370 ;
        RECT 7.0120 26.7435 7.0380 27.8370 ;
        RECT 6.9040 26.7435 6.9300 27.8370 ;
        RECT 6.7960 26.7435 6.8220 27.8370 ;
        RECT 6.6880 26.7435 6.7140 27.8370 ;
        RECT 6.5800 26.7435 6.6060 27.8370 ;
        RECT 6.4720 26.7435 6.4980 27.8370 ;
        RECT 6.3640 26.7435 6.3900 27.8370 ;
        RECT 6.2560 26.7435 6.2820 27.8370 ;
        RECT 6.1480 26.7435 6.1740 27.8370 ;
        RECT 6.0400 26.7435 6.0660 27.8370 ;
        RECT 5.9320 26.7435 5.9580 27.8370 ;
        RECT 5.8240 26.7435 5.8500 27.8370 ;
        RECT 5.7160 26.7435 5.7420 27.8370 ;
        RECT 5.6080 26.7435 5.6340 27.8370 ;
        RECT 5.5000 26.7435 5.5260 27.8370 ;
        RECT 5.3920 26.7435 5.4180 27.8370 ;
        RECT 5.2840 26.7435 5.3100 27.8370 ;
        RECT 5.1760 26.7435 5.2020 27.8370 ;
        RECT 5.0680 26.7435 5.0940 27.8370 ;
        RECT 4.9600 26.7435 4.9860 27.8370 ;
        RECT 4.8520 26.7435 4.8780 27.8370 ;
        RECT 4.7440 26.7435 4.7700 27.8370 ;
        RECT 4.6360 26.7435 4.6620 27.8370 ;
        RECT 4.5280 26.7435 4.5540 27.8370 ;
        RECT 4.4200 26.7435 4.4460 27.8370 ;
        RECT 4.3120 26.7435 4.3380 27.8370 ;
        RECT 4.2040 26.7435 4.2300 27.8370 ;
        RECT 4.0960 26.7435 4.1220 27.8370 ;
        RECT 3.9880 26.7435 4.0140 27.8370 ;
        RECT 3.8800 26.7435 3.9060 27.8370 ;
        RECT 3.7720 26.7435 3.7980 27.8370 ;
        RECT 3.6640 26.7435 3.6900 27.8370 ;
        RECT 3.5560 26.7435 3.5820 27.8370 ;
        RECT 3.4480 26.7435 3.4740 27.8370 ;
        RECT 3.3400 26.7435 3.3660 27.8370 ;
        RECT 3.2320 26.7435 3.2580 27.8370 ;
        RECT 3.1240 26.7435 3.1500 27.8370 ;
        RECT 3.0160 26.7435 3.0420 27.8370 ;
        RECT 2.9080 26.7435 2.9340 27.8370 ;
        RECT 2.8000 26.7435 2.8260 27.8370 ;
        RECT 2.6920 26.7435 2.7180 27.8370 ;
        RECT 2.5840 26.7435 2.6100 27.8370 ;
        RECT 2.4760 26.7435 2.5020 27.8370 ;
        RECT 2.3680 26.7435 2.3940 27.8370 ;
        RECT 2.2600 26.7435 2.2860 27.8370 ;
        RECT 2.1520 26.7435 2.1780 27.8370 ;
        RECT 2.0440 26.7435 2.0700 27.8370 ;
        RECT 1.9360 26.7435 1.9620 27.8370 ;
        RECT 1.8280 26.7435 1.8540 27.8370 ;
        RECT 1.7200 26.7435 1.7460 27.8370 ;
        RECT 1.6120 26.7435 1.6380 27.8370 ;
        RECT 1.5040 26.7435 1.5300 27.8370 ;
        RECT 1.3960 26.7435 1.4220 27.8370 ;
        RECT 1.2880 26.7435 1.3140 27.8370 ;
        RECT 1.1800 26.7435 1.2060 27.8370 ;
        RECT 1.0720 26.7435 1.0980 27.8370 ;
        RECT 0.9640 26.7435 0.9900 27.8370 ;
        RECT 0.8560 26.7435 0.8820 27.8370 ;
        RECT 0.7480 26.7435 0.7740 27.8370 ;
        RECT 0.6400 26.7435 0.6660 27.8370 ;
        RECT 0.5320 26.7435 0.5580 27.8370 ;
        RECT 0.4240 26.7435 0.4500 27.8370 ;
        RECT 0.3160 26.7435 0.3420 27.8370 ;
        RECT 0.2080 26.7435 0.2340 27.8370 ;
        RECT 0.0050 26.7435 0.0900 27.8370 ;
        RECT 15.5530 27.8235 15.6810 28.9170 ;
        RECT 15.5390 28.4890 15.6810 28.8115 ;
        RECT 15.3190 28.2160 15.4530 28.9170 ;
        RECT 15.2960 28.5510 15.4530 28.8090 ;
        RECT 15.3190 27.8235 15.4170 28.9170 ;
        RECT 15.3190 27.9445 15.4310 28.1840 ;
        RECT 15.3190 27.8235 15.4530 27.9125 ;
        RECT 15.0940 28.2740 15.2280 28.9170 ;
        RECT 15.0940 27.8235 15.1920 28.9170 ;
        RECT 14.6770 27.8235 14.7600 28.9170 ;
        RECT 14.6770 27.9120 14.7740 28.8475 ;
        RECT 30.2680 27.8235 30.3530 28.9170 ;
        RECT 30.1240 27.8235 30.1500 28.9170 ;
        RECT 30.0160 27.8235 30.0420 28.9170 ;
        RECT 29.9080 27.8235 29.9340 28.9170 ;
        RECT 29.8000 27.8235 29.8260 28.9170 ;
        RECT 29.6920 27.8235 29.7180 28.9170 ;
        RECT 29.5840 27.8235 29.6100 28.9170 ;
        RECT 29.4760 27.8235 29.5020 28.9170 ;
        RECT 29.3680 27.8235 29.3940 28.9170 ;
        RECT 29.2600 27.8235 29.2860 28.9170 ;
        RECT 29.1520 27.8235 29.1780 28.9170 ;
        RECT 29.0440 27.8235 29.0700 28.9170 ;
        RECT 28.9360 27.8235 28.9620 28.9170 ;
        RECT 28.8280 27.8235 28.8540 28.9170 ;
        RECT 28.7200 27.8235 28.7460 28.9170 ;
        RECT 28.6120 27.8235 28.6380 28.9170 ;
        RECT 28.5040 27.8235 28.5300 28.9170 ;
        RECT 28.3960 27.8235 28.4220 28.9170 ;
        RECT 28.2880 27.8235 28.3140 28.9170 ;
        RECT 28.1800 27.8235 28.2060 28.9170 ;
        RECT 28.0720 27.8235 28.0980 28.9170 ;
        RECT 27.9640 27.8235 27.9900 28.9170 ;
        RECT 27.8560 27.8235 27.8820 28.9170 ;
        RECT 27.7480 27.8235 27.7740 28.9170 ;
        RECT 27.6400 27.8235 27.6660 28.9170 ;
        RECT 27.5320 27.8235 27.5580 28.9170 ;
        RECT 27.4240 27.8235 27.4500 28.9170 ;
        RECT 27.3160 27.8235 27.3420 28.9170 ;
        RECT 27.2080 27.8235 27.2340 28.9170 ;
        RECT 27.1000 27.8235 27.1260 28.9170 ;
        RECT 26.9920 27.8235 27.0180 28.9170 ;
        RECT 26.8840 27.8235 26.9100 28.9170 ;
        RECT 26.7760 27.8235 26.8020 28.9170 ;
        RECT 26.6680 27.8235 26.6940 28.9170 ;
        RECT 26.5600 27.8235 26.5860 28.9170 ;
        RECT 26.4520 27.8235 26.4780 28.9170 ;
        RECT 26.3440 27.8235 26.3700 28.9170 ;
        RECT 26.2360 27.8235 26.2620 28.9170 ;
        RECT 26.1280 27.8235 26.1540 28.9170 ;
        RECT 26.0200 27.8235 26.0460 28.9170 ;
        RECT 25.9120 27.8235 25.9380 28.9170 ;
        RECT 25.8040 27.8235 25.8300 28.9170 ;
        RECT 25.6960 27.8235 25.7220 28.9170 ;
        RECT 25.5880 27.8235 25.6140 28.9170 ;
        RECT 25.4800 27.8235 25.5060 28.9170 ;
        RECT 25.3720 27.8235 25.3980 28.9170 ;
        RECT 25.2640 27.8235 25.2900 28.9170 ;
        RECT 25.1560 27.8235 25.1820 28.9170 ;
        RECT 25.0480 27.8235 25.0740 28.9170 ;
        RECT 24.9400 27.8235 24.9660 28.9170 ;
        RECT 24.8320 27.8235 24.8580 28.9170 ;
        RECT 24.7240 27.8235 24.7500 28.9170 ;
        RECT 24.6160 27.8235 24.6420 28.9170 ;
        RECT 24.5080 27.8235 24.5340 28.9170 ;
        RECT 24.4000 27.8235 24.4260 28.9170 ;
        RECT 24.2920 27.8235 24.3180 28.9170 ;
        RECT 24.1840 27.8235 24.2100 28.9170 ;
        RECT 24.0760 27.8235 24.1020 28.9170 ;
        RECT 23.9680 27.8235 23.9940 28.9170 ;
        RECT 23.8600 27.8235 23.8860 28.9170 ;
        RECT 23.7520 27.8235 23.7780 28.9170 ;
        RECT 23.6440 27.8235 23.6700 28.9170 ;
        RECT 23.5360 27.8235 23.5620 28.9170 ;
        RECT 23.4280 27.8235 23.4540 28.9170 ;
        RECT 23.3200 27.8235 23.3460 28.9170 ;
        RECT 23.2120 27.8235 23.2380 28.9170 ;
        RECT 23.1040 27.8235 23.1300 28.9170 ;
        RECT 22.9960 27.8235 23.0220 28.9170 ;
        RECT 22.8880 27.8235 22.9140 28.9170 ;
        RECT 22.7800 27.8235 22.8060 28.9170 ;
        RECT 22.6720 27.8235 22.6980 28.9170 ;
        RECT 22.5640 27.8235 22.5900 28.9170 ;
        RECT 22.4560 27.8235 22.4820 28.9170 ;
        RECT 22.3480 27.8235 22.3740 28.9170 ;
        RECT 22.2400 27.8235 22.2660 28.9170 ;
        RECT 22.1320 27.8235 22.1580 28.9170 ;
        RECT 22.0240 27.8235 22.0500 28.9170 ;
        RECT 21.9160 27.8235 21.9420 28.9170 ;
        RECT 21.8080 27.8235 21.8340 28.9170 ;
        RECT 21.7000 27.8235 21.7260 28.9170 ;
        RECT 21.5920 27.8235 21.6180 28.9170 ;
        RECT 21.4840 27.8235 21.5100 28.9170 ;
        RECT 21.3760 27.8235 21.4020 28.9170 ;
        RECT 21.2680 27.8235 21.2940 28.9170 ;
        RECT 21.1600 27.8235 21.1860 28.9170 ;
        RECT 21.0520 27.8235 21.0780 28.9170 ;
        RECT 20.9440 27.8235 20.9700 28.9170 ;
        RECT 20.8360 27.8235 20.8620 28.9170 ;
        RECT 20.7280 27.8235 20.7540 28.9170 ;
        RECT 20.6200 27.8235 20.6460 28.9170 ;
        RECT 20.5120 27.8235 20.5380 28.9170 ;
        RECT 20.4040 27.8235 20.4300 28.9170 ;
        RECT 20.2960 27.8235 20.3220 28.9170 ;
        RECT 20.1880 27.8235 20.2140 28.9170 ;
        RECT 20.0800 27.8235 20.1060 28.9170 ;
        RECT 19.9720 27.8235 19.9980 28.9170 ;
        RECT 19.8640 27.8235 19.8900 28.9170 ;
        RECT 19.7560 27.8235 19.7820 28.9170 ;
        RECT 19.6480 27.8235 19.6740 28.9170 ;
        RECT 19.5400 27.8235 19.5660 28.9170 ;
        RECT 19.4320 27.8235 19.4580 28.9170 ;
        RECT 19.3240 27.8235 19.3500 28.9170 ;
        RECT 19.2160 27.8235 19.2420 28.9170 ;
        RECT 19.1080 27.8235 19.1340 28.9170 ;
        RECT 19.0000 27.8235 19.0260 28.9170 ;
        RECT 18.8920 27.8235 18.9180 28.9170 ;
        RECT 18.7840 27.8235 18.8100 28.9170 ;
        RECT 18.6760 27.8235 18.7020 28.9170 ;
        RECT 18.5680 27.8235 18.5940 28.9170 ;
        RECT 18.4600 27.8235 18.4860 28.9170 ;
        RECT 18.3520 27.8235 18.3780 28.9170 ;
        RECT 18.2440 27.8235 18.2700 28.9170 ;
        RECT 18.1360 27.8235 18.1620 28.9170 ;
        RECT 18.0280 27.8235 18.0540 28.9170 ;
        RECT 17.9200 27.8235 17.9460 28.9170 ;
        RECT 17.8120 27.8235 17.8380 28.9170 ;
        RECT 17.7040 27.8235 17.7300 28.9170 ;
        RECT 17.5960 27.8235 17.6220 28.9170 ;
        RECT 17.4880 27.8235 17.5140 28.9170 ;
        RECT 17.3800 27.8235 17.4060 28.9170 ;
        RECT 17.2720 27.8235 17.2980 28.9170 ;
        RECT 17.1640 27.8235 17.1900 28.9170 ;
        RECT 17.0560 27.8235 17.0820 28.9170 ;
        RECT 16.9480 27.8235 16.9740 28.9170 ;
        RECT 16.8400 27.8235 16.8660 28.9170 ;
        RECT 16.7320 27.8235 16.7580 28.9170 ;
        RECT 16.6240 27.8235 16.6500 28.9170 ;
        RECT 16.5160 27.8235 16.5420 28.9170 ;
        RECT 16.4080 27.8235 16.4340 28.9170 ;
        RECT 16.3000 27.8235 16.3260 28.9170 ;
        RECT 16.0870 27.8235 16.1640 28.9170 ;
        RECT 14.1940 27.8235 14.2710 28.9170 ;
        RECT 14.0320 27.8235 14.0580 28.9170 ;
        RECT 13.9240 27.8235 13.9500 28.9170 ;
        RECT 13.8160 27.8235 13.8420 28.9170 ;
        RECT 13.7080 27.8235 13.7340 28.9170 ;
        RECT 13.6000 27.8235 13.6260 28.9170 ;
        RECT 13.4920 27.8235 13.5180 28.9170 ;
        RECT 13.3840 27.8235 13.4100 28.9170 ;
        RECT 13.2760 27.8235 13.3020 28.9170 ;
        RECT 13.1680 27.8235 13.1940 28.9170 ;
        RECT 13.0600 27.8235 13.0860 28.9170 ;
        RECT 12.9520 27.8235 12.9780 28.9170 ;
        RECT 12.8440 27.8235 12.8700 28.9170 ;
        RECT 12.7360 27.8235 12.7620 28.9170 ;
        RECT 12.6280 27.8235 12.6540 28.9170 ;
        RECT 12.5200 27.8235 12.5460 28.9170 ;
        RECT 12.4120 27.8235 12.4380 28.9170 ;
        RECT 12.3040 27.8235 12.3300 28.9170 ;
        RECT 12.1960 27.8235 12.2220 28.9170 ;
        RECT 12.0880 27.8235 12.1140 28.9170 ;
        RECT 11.9800 27.8235 12.0060 28.9170 ;
        RECT 11.8720 27.8235 11.8980 28.9170 ;
        RECT 11.7640 27.8235 11.7900 28.9170 ;
        RECT 11.6560 27.8235 11.6820 28.9170 ;
        RECT 11.5480 27.8235 11.5740 28.9170 ;
        RECT 11.4400 27.8235 11.4660 28.9170 ;
        RECT 11.3320 27.8235 11.3580 28.9170 ;
        RECT 11.2240 27.8235 11.2500 28.9170 ;
        RECT 11.1160 27.8235 11.1420 28.9170 ;
        RECT 11.0080 27.8235 11.0340 28.9170 ;
        RECT 10.9000 27.8235 10.9260 28.9170 ;
        RECT 10.7920 27.8235 10.8180 28.9170 ;
        RECT 10.6840 27.8235 10.7100 28.9170 ;
        RECT 10.5760 27.8235 10.6020 28.9170 ;
        RECT 10.4680 27.8235 10.4940 28.9170 ;
        RECT 10.3600 27.8235 10.3860 28.9170 ;
        RECT 10.2520 27.8235 10.2780 28.9170 ;
        RECT 10.1440 27.8235 10.1700 28.9170 ;
        RECT 10.0360 27.8235 10.0620 28.9170 ;
        RECT 9.9280 27.8235 9.9540 28.9170 ;
        RECT 9.8200 27.8235 9.8460 28.9170 ;
        RECT 9.7120 27.8235 9.7380 28.9170 ;
        RECT 9.6040 27.8235 9.6300 28.9170 ;
        RECT 9.4960 27.8235 9.5220 28.9170 ;
        RECT 9.3880 27.8235 9.4140 28.9170 ;
        RECT 9.2800 27.8235 9.3060 28.9170 ;
        RECT 9.1720 27.8235 9.1980 28.9170 ;
        RECT 9.0640 27.8235 9.0900 28.9170 ;
        RECT 8.9560 27.8235 8.9820 28.9170 ;
        RECT 8.8480 27.8235 8.8740 28.9170 ;
        RECT 8.7400 27.8235 8.7660 28.9170 ;
        RECT 8.6320 27.8235 8.6580 28.9170 ;
        RECT 8.5240 27.8235 8.5500 28.9170 ;
        RECT 8.4160 27.8235 8.4420 28.9170 ;
        RECT 8.3080 27.8235 8.3340 28.9170 ;
        RECT 8.2000 27.8235 8.2260 28.9170 ;
        RECT 8.0920 27.8235 8.1180 28.9170 ;
        RECT 7.9840 27.8235 8.0100 28.9170 ;
        RECT 7.8760 27.8235 7.9020 28.9170 ;
        RECT 7.7680 27.8235 7.7940 28.9170 ;
        RECT 7.6600 27.8235 7.6860 28.9170 ;
        RECT 7.5520 27.8235 7.5780 28.9170 ;
        RECT 7.4440 27.8235 7.4700 28.9170 ;
        RECT 7.3360 27.8235 7.3620 28.9170 ;
        RECT 7.2280 27.8235 7.2540 28.9170 ;
        RECT 7.1200 27.8235 7.1460 28.9170 ;
        RECT 7.0120 27.8235 7.0380 28.9170 ;
        RECT 6.9040 27.8235 6.9300 28.9170 ;
        RECT 6.7960 27.8235 6.8220 28.9170 ;
        RECT 6.6880 27.8235 6.7140 28.9170 ;
        RECT 6.5800 27.8235 6.6060 28.9170 ;
        RECT 6.4720 27.8235 6.4980 28.9170 ;
        RECT 6.3640 27.8235 6.3900 28.9170 ;
        RECT 6.2560 27.8235 6.2820 28.9170 ;
        RECT 6.1480 27.8235 6.1740 28.9170 ;
        RECT 6.0400 27.8235 6.0660 28.9170 ;
        RECT 5.9320 27.8235 5.9580 28.9170 ;
        RECT 5.8240 27.8235 5.8500 28.9170 ;
        RECT 5.7160 27.8235 5.7420 28.9170 ;
        RECT 5.6080 27.8235 5.6340 28.9170 ;
        RECT 5.5000 27.8235 5.5260 28.9170 ;
        RECT 5.3920 27.8235 5.4180 28.9170 ;
        RECT 5.2840 27.8235 5.3100 28.9170 ;
        RECT 5.1760 27.8235 5.2020 28.9170 ;
        RECT 5.0680 27.8235 5.0940 28.9170 ;
        RECT 4.9600 27.8235 4.9860 28.9170 ;
        RECT 4.8520 27.8235 4.8780 28.9170 ;
        RECT 4.7440 27.8235 4.7700 28.9170 ;
        RECT 4.6360 27.8235 4.6620 28.9170 ;
        RECT 4.5280 27.8235 4.5540 28.9170 ;
        RECT 4.4200 27.8235 4.4460 28.9170 ;
        RECT 4.3120 27.8235 4.3380 28.9170 ;
        RECT 4.2040 27.8235 4.2300 28.9170 ;
        RECT 4.0960 27.8235 4.1220 28.9170 ;
        RECT 3.9880 27.8235 4.0140 28.9170 ;
        RECT 3.8800 27.8235 3.9060 28.9170 ;
        RECT 3.7720 27.8235 3.7980 28.9170 ;
        RECT 3.6640 27.8235 3.6900 28.9170 ;
        RECT 3.5560 27.8235 3.5820 28.9170 ;
        RECT 3.4480 27.8235 3.4740 28.9170 ;
        RECT 3.3400 27.8235 3.3660 28.9170 ;
        RECT 3.2320 27.8235 3.2580 28.9170 ;
        RECT 3.1240 27.8235 3.1500 28.9170 ;
        RECT 3.0160 27.8235 3.0420 28.9170 ;
        RECT 2.9080 27.8235 2.9340 28.9170 ;
        RECT 2.8000 27.8235 2.8260 28.9170 ;
        RECT 2.6920 27.8235 2.7180 28.9170 ;
        RECT 2.5840 27.8235 2.6100 28.9170 ;
        RECT 2.4760 27.8235 2.5020 28.9170 ;
        RECT 2.3680 27.8235 2.3940 28.9170 ;
        RECT 2.2600 27.8235 2.2860 28.9170 ;
        RECT 2.1520 27.8235 2.1780 28.9170 ;
        RECT 2.0440 27.8235 2.0700 28.9170 ;
        RECT 1.9360 27.8235 1.9620 28.9170 ;
        RECT 1.8280 27.8235 1.8540 28.9170 ;
        RECT 1.7200 27.8235 1.7460 28.9170 ;
        RECT 1.6120 27.8235 1.6380 28.9170 ;
        RECT 1.5040 27.8235 1.5300 28.9170 ;
        RECT 1.3960 27.8235 1.4220 28.9170 ;
        RECT 1.2880 27.8235 1.3140 28.9170 ;
        RECT 1.1800 27.8235 1.2060 28.9170 ;
        RECT 1.0720 27.8235 1.0980 28.9170 ;
        RECT 0.9640 27.8235 0.9900 28.9170 ;
        RECT 0.8560 27.8235 0.8820 28.9170 ;
        RECT 0.7480 27.8235 0.7740 28.9170 ;
        RECT 0.6400 27.8235 0.6660 28.9170 ;
        RECT 0.5320 27.8235 0.5580 28.9170 ;
        RECT 0.4240 27.8235 0.4500 28.9170 ;
        RECT 0.3160 27.8235 0.3420 28.9170 ;
        RECT 0.2080 27.8235 0.2340 28.9170 ;
        RECT 0.0050 27.8235 0.0900 28.9170 ;
        RECT 15.5530 28.9035 15.6810 29.9970 ;
        RECT 15.5390 29.5690 15.6810 29.8915 ;
        RECT 15.3190 29.2960 15.4530 29.9970 ;
        RECT 15.2960 29.6310 15.4530 29.8890 ;
        RECT 15.3190 28.9035 15.4170 29.9970 ;
        RECT 15.3190 29.0245 15.4310 29.2640 ;
        RECT 15.3190 28.9035 15.4530 28.9925 ;
        RECT 15.0940 29.3540 15.2280 29.9970 ;
        RECT 15.0940 28.9035 15.1920 29.9970 ;
        RECT 14.6770 28.9035 14.7600 29.9970 ;
        RECT 14.6770 28.9920 14.7740 29.9275 ;
        RECT 30.2680 28.9035 30.3530 29.9970 ;
        RECT 30.1240 28.9035 30.1500 29.9970 ;
        RECT 30.0160 28.9035 30.0420 29.9970 ;
        RECT 29.9080 28.9035 29.9340 29.9970 ;
        RECT 29.8000 28.9035 29.8260 29.9970 ;
        RECT 29.6920 28.9035 29.7180 29.9970 ;
        RECT 29.5840 28.9035 29.6100 29.9970 ;
        RECT 29.4760 28.9035 29.5020 29.9970 ;
        RECT 29.3680 28.9035 29.3940 29.9970 ;
        RECT 29.2600 28.9035 29.2860 29.9970 ;
        RECT 29.1520 28.9035 29.1780 29.9970 ;
        RECT 29.0440 28.9035 29.0700 29.9970 ;
        RECT 28.9360 28.9035 28.9620 29.9970 ;
        RECT 28.8280 28.9035 28.8540 29.9970 ;
        RECT 28.7200 28.9035 28.7460 29.9970 ;
        RECT 28.6120 28.9035 28.6380 29.9970 ;
        RECT 28.5040 28.9035 28.5300 29.9970 ;
        RECT 28.3960 28.9035 28.4220 29.9970 ;
        RECT 28.2880 28.9035 28.3140 29.9970 ;
        RECT 28.1800 28.9035 28.2060 29.9970 ;
        RECT 28.0720 28.9035 28.0980 29.9970 ;
        RECT 27.9640 28.9035 27.9900 29.9970 ;
        RECT 27.8560 28.9035 27.8820 29.9970 ;
        RECT 27.7480 28.9035 27.7740 29.9970 ;
        RECT 27.6400 28.9035 27.6660 29.9970 ;
        RECT 27.5320 28.9035 27.5580 29.9970 ;
        RECT 27.4240 28.9035 27.4500 29.9970 ;
        RECT 27.3160 28.9035 27.3420 29.9970 ;
        RECT 27.2080 28.9035 27.2340 29.9970 ;
        RECT 27.1000 28.9035 27.1260 29.9970 ;
        RECT 26.9920 28.9035 27.0180 29.9970 ;
        RECT 26.8840 28.9035 26.9100 29.9970 ;
        RECT 26.7760 28.9035 26.8020 29.9970 ;
        RECT 26.6680 28.9035 26.6940 29.9970 ;
        RECT 26.5600 28.9035 26.5860 29.9970 ;
        RECT 26.4520 28.9035 26.4780 29.9970 ;
        RECT 26.3440 28.9035 26.3700 29.9970 ;
        RECT 26.2360 28.9035 26.2620 29.9970 ;
        RECT 26.1280 28.9035 26.1540 29.9970 ;
        RECT 26.0200 28.9035 26.0460 29.9970 ;
        RECT 25.9120 28.9035 25.9380 29.9970 ;
        RECT 25.8040 28.9035 25.8300 29.9970 ;
        RECT 25.6960 28.9035 25.7220 29.9970 ;
        RECT 25.5880 28.9035 25.6140 29.9970 ;
        RECT 25.4800 28.9035 25.5060 29.9970 ;
        RECT 25.3720 28.9035 25.3980 29.9970 ;
        RECT 25.2640 28.9035 25.2900 29.9970 ;
        RECT 25.1560 28.9035 25.1820 29.9970 ;
        RECT 25.0480 28.9035 25.0740 29.9970 ;
        RECT 24.9400 28.9035 24.9660 29.9970 ;
        RECT 24.8320 28.9035 24.8580 29.9970 ;
        RECT 24.7240 28.9035 24.7500 29.9970 ;
        RECT 24.6160 28.9035 24.6420 29.9970 ;
        RECT 24.5080 28.9035 24.5340 29.9970 ;
        RECT 24.4000 28.9035 24.4260 29.9970 ;
        RECT 24.2920 28.9035 24.3180 29.9970 ;
        RECT 24.1840 28.9035 24.2100 29.9970 ;
        RECT 24.0760 28.9035 24.1020 29.9970 ;
        RECT 23.9680 28.9035 23.9940 29.9970 ;
        RECT 23.8600 28.9035 23.8860 29.9970 ;
        RECT 23.7520 28.9035 23.7780 29.9970 ;
        RECT 23.6440 28.9035 23.6700 29.9970 ;
        RECT 23.5360 28.9035 23.5620 29.9970 ;
        RECT 23.4280 28.9035 23.4540 29.9970 ;
        RECT 23.3200 28.9035 23.3460 29.9970 ;
        RECT 23.2120 28.9035 23.2380 29.9970 ;
        RECT 23.1040 28.9035 23.1300 29.9970 ;
        RECT 22.9960 28.9035 23.0220 29.9970 ;
        RECT 22.8880 28.9035 22.9140 29.9970 ;
        RECT 22.7800 28.9035 22.8060 29.9970 ;
        RECT 22.6720 28.9035 22.6980 29.9970 ;
        RECT 22.5640 28.9035 22.5900 29.9970 ;
        RECT 22.4560 28.9035 22.4820 29.9970 ;
        RECT 22.3480 28.9035 22.3740 29.9970 ;
        RECT 22.2400 28.9035 22.2660 29.9970 ;
        RECT 22.1320 28.9035 22.1580 29.9970 ;
        RECT 22.0240 28.9035 22.0500 29.9970 ;
        RECT 21.9160 28.9035 21.9420 29.9970 ;
        RECT 21.8080 28.9035 21.8340 29.9970 ;
        RECT 21.7000 28.9035 21.7260 29.9970 ;
        RECT 21.5920 28.9035 21.6180 29.9970 ;
        RECT 21.4840 28.9035 21.5100 29.9970 ;
        RECT 21.3760 28.9035 21.4020 29.9970 ;
        RECT 21.2680 28.9035 21.2940 29.9970 ;
        RECT 21.1600 28.9035 21.1860 29.9970 ;
        RECT 21.0520 28.9035 21.0780 29.9970 ;
        RECT 20.9440 28.9035 20.9700 29.9970 ;
        RECT 20.8360 28.9035 20.8620 29.9970 ;
        RECT 20.7280 28.9035 20.7540 29.9970 ;
        RECT 20.6200 28.9035 20.6460 29.9970 ;
        RECT 20.5120 28.9035 20.5380 29.9970 ;
        RECT 20.4040 28.9035 20.4300 29.9970 ;
        RECT 20.2960 28.9035 20.3220 29.9970 ;
        RECT 20.1880 28.9035 20.2140 29.9970 ;
        RECT 20.0800 28.9035 20.1060 29.9970 ;
        RECT 19.9720 28.9035 19.9980 29.9970 ;
        RECT 19.8640 28.9035 19.8900 29.9970 ;
        RECT 19.7560 28.9035 19.7820 29.9970 ;
        RECT 19.6480 28.9035 19.6740 29.9970 ;
        RECT 19.5400 28.9035 19.5660 29.9970 ;
        RECT 19.4320 28.9035 19.4580 29.9970 ;
        RECT 19.3240 28.9035 19.3500 29.9970 ;
        RECT 19.2160 28.9035 19.2420 29.9970 ;
        RECT 19.1080 28.9035 19.1340 29.9970 ;
        RECT 19.0000 28.9035 19.0260 29.9970 ;
        RECT 18.8920 28.9035 18.9180 29.9970 ;
        RECT 18.7840 28.9035 18.8100 29.9970 ;
        RECT 18.6760 28.9035 18.7020 29.9970 ;
        RECT 18.5680 28.9035 18.5940 29.9970 ;
        RECT 18.4600 28.9035 18.4860 29.9970 ;
        RECT 18.3520 28.9035 18.3780 29.9970 ;
        RECT 18.2440 28.9035 18.2700 29.9970 ;
        RECT 18.1360 28.9035 18.1620 29.9970 ;
        RECT 18.0280 28.9035 18.0540 29.9970 ;
        RECT 17.9200 28.9035 17.9460 29.9970 ;
        RECT 17.8120 28.9035 17.8380 29.9970 ;
        RECT 17.7040 28.9035 17.7300 29.9970 ;
        RECT 17.5960 28.9035 17.6220 29.9970 ;
        RECT 17.4880 28.9035 17.5140 29.9970 ;
        RECT 17.3800 28.9035 17.4060 29.9970 ;
        RECT 17.2720 28.9035 17.2980 29.9970 ;
        RECT 17.1640 28.9035 17.1900 29.9970 ;
        RECT 17.0560 28.9035 17.0820 29.9970 ;
        RECT 16.9480 28.9035 16.9740 29.9970 ;
        RECT 16.8400 28.9035 16.8660 29.9970 ;
        RECT 16.7320 28.9035 16.7580 29.9970 ;
        RECT 16.6240 28.9035 16.6500 29.9970 ;
        RECT 16.5160 28.9035 16.5420 29.9970 ;
        RECT 16.4080 28.9035 16.4340 29.9970 ;
        RECT 16.3000 28.9035 16.3260 29.9970 ;
        RECT 16.0870 28.9035 16.1640 29.9970 ;
        RECT 14.1940 28.9035 14.2710 29.9970 ;
        RECT 14.0320 28.9035 14.0580 29.9970 ;
        RECT 13.9240 28.9035 13.9500 29.9970 ;
        RECT 13.8160 28.9035 13.8420 29.9970 ;
        RECT 13.7080 28.9035 13.7340 29.9970 ;
        RECT 13.6000 28.9035 13.6260 29.9970 ;
        RECT 13.4920 28.9035 13.5180 29.9970 ;
        RECT 13.3840 28.9035 13.4100 29.9970 ;
        RECT 13.2760 28.9035 13.3020 29.9970 ;
        RECT 13.1680 28.9035 13.1940 29.9970 ;
        RECT 13.0600 28.9035 13.0860 29.9970 ;
        RECT 12.9520 28.9035 12.9780 29.9970 ;
        RECT 12.8440 28.9035 12.8700 29.9970 ;
        RECT 12.7360 28.9035 12.7620 29.9970 ;
        RECT 12.6280 28.9035 12.6540 29.9970 ;
        RECT 12.5200 28.9035 12.5460 29.9970 ;
        RECT 12.4120 28.9035 12.4380 29.9970 ;
        RECT 12.3040 28.9035 12.3300 29.9970 ;
        RECT 12.1960 28.9035 12.2220 29.9970 ;
        RECT 12.0880 28.9035 12.1140 29.9970 ;
        RECT 11.9800 28.9035 12.0060 29.9970 ;
        RECT 11.8720 28.9035 11.8980 29.9970 ;
        RECT 11.7640 28.9035 11.7900 29.9970 ;
        RECT 11.6560 28.9035 11.6820 29.9970 ;
        RECT 11.5480 28.9035 11.5740 29.9970 ;
        RECT 11.4400 28.9035 11.4660 29.9970 ;
        RECT 11.3320 28.9035 11.3580 29.9970 ;
        RECT 11.2240 28.9035 11.2500 29.9970 ;
        RECT 11.1160 28.9035 11.1420 29.9970 ;
        RECT 11.0080 28.9035 11.0340 29.9970 ;
        RECT 10.9000 28.9035 10.9260 29.9970 ;
        RECT 10.7920 28.9035 10.8180 29.9970 ;
        RECT 10.6840 28.9035 10.7100 29.9970 ;
        RECT 10.5760 28.9035 10.6020 29.9970 ;
        RECT 10.4680 28.9035 10.4940 29.9970 ;
        RECT 10.3600 28.9035 10.3860 29.9970 ;
        RECT 10.2520 28.9035 10.2780 29.9970 ;
        RECT 10.1440 28.9035 10.1700 29.9970 ;
        RECT 10.0360 28.9035 10.0620 29.9970 ;
        RECT 9.9280 28.9035 9.9540 29.9970 ;
        RECT 9.8200 28.9035 9.8460 29.9970 ;
        RECT 9.7120 28.9035 9.7380 29.9970 ;
        RECT 9.6040 28.9035 9.6300 29.9970 ;
        RECT 9.4960 28.9035 9.5220 29.9970 ;
        RECT 9.3880 28.9035 9.4140 29.9970 ;
        RECT 9.2800 28.9035 9.3060 29.9970 ;
        RECT 9.1720 28.9035 9.1980 29.9970 ;
        RECT 9.0640 28.9035 9.0900 29.9970 ;
        RECT 8.9560 28.9035 8.9820 29.9970 ;
        RECT 8.8480 28.9035 8.8740 29.9970 ;
        RECT 8.7400 28.9035 8.7660 29.9970 ;
        RECT 8.6320 28.9035 8.6580 29.9970 ;
        RECT 8.5240 28.9035 8.5500 29.9970 ;
        RECT 8.4160 28.9035 8.4420 29.9970 ;
        RECT 8.3080 28.9035 8.3340 29.9970 ;
        RECT 8.2000 28.9035 8.2260 29.9970 ;
        RECT 8.0920 28.9035 8.1180 29.9970 ;
        RECT 7.9840 28.9035 8.0100 29.9970 ;
        RECT 7.8760 28.9035 7.9020 29.9970 ;
        RECT 7.7680 28.9035 7.7940 29.9970 ;
        RECT 7.6600 28.9035 7.6860 29.9970 ;
        RECT 7.5520 28.9035 7.5780 29.9970 ;
        RECT 7.4440 28.9035 7.4700 29.9970 ;
        RECT 7.3360 28.9035 7.3620 29.9970 ;
        RECT 7.2280 28.9035 7.2540 29.9970 ;
        RECT 7.1200 28.9035 7.1460 29.9970 ;
        RECT 7.0120 28.9035 7.0380 29.9970 ;
        RECT 6.9040 28.9035 6.9300 29.9970 ;
        RECT 6.7960 28.9035 6.8220 29.9970 ;
        RECT 6.6880 28.9035 6.7140 29.9970 ;
        RECT 6.5800 28.9035 6.6060 29.9970 ;
        RECT 6.4720 28.9035 6.4980 29.9970 ;
        RECT 6.3640 28.9035 6.3900 29.9970 ;
        RECT 6.2560 28.9035 6.2820 29.9970 ;
        RECT 6.1480 28.9035 6.1740 29.9970 ;
        RECT 6.0400 28.9035 6.0660 29.9970 ;
        RECT 5.9320 28.9035 5.9580 29.9970 ;
        RECT 5.8240 28.9035 5.8500 29.9970 ;
        RECT 5.7160 28.9035 5.7420 29.9970 ;
        RECT 5.6080 28.9035 5.6340 29.9970 ;
        RECT 5.5000 28.9035 5.5260 29.9970 ;
        RECT 5.3920 28.9035 5.4180 29.9970 ;
        RECT 5.2840 28.9035 5.3100 29.9970 ;
        RECT 5.1760 28.9035 5.2020 29.9970 ;
        RECT 5.0680 28.9035 5.0940 29.9970 ;
        RECT 4.9600 28.9035 4.9860 29.9970 ;
        RECT 4.8520 28.9035 4.8780 29.9970 ;
        RECT 4.7440 28.9035 4.7700 29.9970 ;
        RECT 4.6360 28.9035 4.6620 29.9970 ;
        RECT 4.5280 28.9035 4.5540 29.9970 ;
        RECT 4.4200 28.9035 4.4460 29.9970 ;
        RECT 4.3120 28.9035 4.3380 29.9970 ;
        RECT 4.2040 28.9035 4.2300 29.9970 ;
        RECT 4.0960 28.9035 4.1220 29.9970 ;
        RECT 3.9880 28.9035 4.0140 29.9970 ;
        RECT 3.8800 28.9035 3.9060 29.9970 ;
        RECT 3.7720 28.9035 3.7980 29.9970 ;
        RECT 3.6640 28.9035 3.6900 29.9970 ;
        RECT 3.5560 28.9035 3.5820 29.9970 ;
        RECT 3.4480 28.9035 3.4740 29.9970 ;
        RECT 3.3400 28.9035 3.3660 29.9970 ;
        RECT 3.2320 28.9035 3.2580 29.9970 ;
        RECT 3.1240 28.9035 3.1500 29.9970 ;
        RECT 3.0160 28.9035 3.0420 29.9970 ;
        RECT 2.9080 28.9035 2.9340 29.9970 ;
        RECT 2.8000 28.9035 2.8260 29.9970 ;
        RECT 2.6920 28.9035 2.7180 29.9970 ;
        RECT 2.5840 28.9035 2.6100 29.9970 ;
        RECT 2.4760 28.9035 2.5020 29.9970 ;
        RECT 2.3680 28.9035 2.3940 29.9970 ;
        RECT 2.2600 28.9035 2.2860 29.9970 ;
        RECT 2.1520 28.9035 2.1780 29.9970 ;
        RECT 2.0440 28.9035 2.0700 29.9970 ;
        RECT 1.9360 28.9035 1.9620 29.9970 ;
        RECT 1.8280 28.9035 1.8540 29.9970 ;
        RECT 1.7200 28.9035 1.7460 29.9970 ;
        RECT 1.6120 28.9035 1.6380 29.9970 ;
        RECT 1.5040 28.9035 1.5300 29.9970 ;
        RECT 1.3960 28.9035 1.4220 29.9970 ;
        RECT 1.2880 28.9035 1.3140 29.9970 ;
        RECT 1.1800 28.9035 1.2060 29.9970 ;
        RECT 1.0720 28.9035 1.0980 29.9970 ;
        RECT 0.9640 28.9035 0.9900 29.9970 ;
        RECT 0.8560 28.9035 0.8820 29.9970 ;
        RECT 0.7480 28.9035 0.7740 29.9970 ;
        RECT 0.6400 28.9035 0.6660 29.9970 ;
        RECT 0.5320 28.9035 0.5580 29.9970 ;
        RECT 0.4240 28.9035 0.4500 29.9970 ;
        RECT 0.3160 28.9035 0.3420 29.9970 ;
        RECT 0.2080 28.9035 0.2340 29.9970 ;
        RECT 0.0050 28.9035 0.0900 29.9970 ;
  LAYER V3 SPACING 0.018  ;
      RECT 0.0050 1.2200 30.3530 1.3500 ;
      RECT 30.2360 0.2565 30.3530 1.3500 ;
      RECT 16.2140 1.1240 30.2180 1.3500 ;
      RECT 14.8820 1.1240 16.1960 1.3500 ;
      RECT 14.1620 0.2565 14.7920 1.3500 ;
      RECT 0.1400 1.1240 14.1440 1.3500 ;
      RECT 0.0050 0.2565 0.1220 1.3500 ;
      RECT 30.2000 0.2565 30.3530 1.1720 ;
      RECT 16.2680 0.2565 30.1820 1.3500 ;
      RECT 15.5210 0.2565 16.2500 1.1720 ;
      RECT 15.2870 0.4520 15.4850 1.3500 ;
      RECT 14.1080 0.3560 15.2600 1.1720 ;
      RECT 0.1760 0.2565 14.0900 1.3500 ;
      RECT 0.0050 0.2565 0.1580 1.1720 ;
      RECT 15.4670 0.2565 30.3530 1.0760 ;
      RECT 0.0050 0.3560 15.4490 1.0760 ;
      RECT 15.2420 0.2565 30.3530 0.4280 ;
      RECT 0.0050 0.2565 15.2240 1.0760 ;
      RECT 0.0050 0.2565 30.3530 0.3320 ;
      RECT 0.0050 2.3000 30.3530 2.4300 ;
      RECT 30.2360 1.3365 30.3530 2.4300 ;
      RECT 16.2140 2.2040 30.2180 2.4300 ;
      RECT 14.8820 2.2040 16.1960 2.4300 ;
      RECT 14.1620 1.3365 14.7920 2.4300 ;
      RECT 0.1400 2.2040 14.1440 2.4300 ;
      RECT 0.0050 1.3365 0.1220 2.4300 ;
      RECT 30.2000 1.3365 30.3530 2.2520 ;
      RECT 16.2680 1.3365 30.1820 2.4300 ;
      RECT 15.5210 1.3365 16.2500 2.2520 ;
      RECT 15.2870 1.5320 15.4850 2.4300 ;
      RECT 14.1080 1.4360 15.2600 2.2520 ;
      RECT 0.1760 1.3365 14.0900 2.4300 ;
      RECT 0.0050 1.3365 0.1580 2.2520 ;
      RECT 15.4670 1.3365 30.3530 2.1560 ;
      RECT 0.0050 1.4360 15.4490 2.1560 ;
      RECT 15.2420 1.3365 30.3530 1.5080 ;
      RECT 0.0050 1.3365 15.2240 2.1560 ;
      RECT 0.0050 1.3365 30.3530 1.4120 ;
      RECT 0.0050 3.3800 30.3530 3.5100 ;
      RECT 30.2360 2.4165 30.3530 3.5100 ;
      RECT 16.2140 3.2840 30.2180 3.5100 ;
      RECT 14.8820 3.2840 16.1960 3.5100 ;
      RECT 14.1620 2.4165 14.7920 3.5100 ;
      RECT 0.1400 3.2840 14.1440 3.5100 ;
      RECT 0.0050 2.4165 0.1220 3.5100 ;
      RECT 30.2000 2.4165 30.3530 3.3320 ;
      RECT 16.2680 2.4165 30.1820 3.5100 ;
      RECT 15.5210 2.4165 16.2500 3.3320 ;
      RECT 15.2870 2.6120 15.4850 3.5100 ;
      RECT 14.1080 2.5160 15.2600 3.3320 ;
      RECT 0.1760 2.4165 14.0900 3.5100 ;
      RECT 0.0050 2.4165 0.1580 3.3320 ;
      RECT 15.4670 2.4165 30.3530 3.2360 ;
      RECT 0.0050 2.5160 15.4490 3.2360 ;
      RECT 15.2420 2.4165 30.3530 2.5880 ;
      RECT 0.0050 2.4165 15.2240 3.2360 ;
      RECT 0.0050 2.4165 30.3530 2.4920 ;
      RECT 0.0050 4.4600 30.3530 4.5900 ;
      RECT 30.2360 3.4965 30.3530 4.5900 ;
      RECT 16.2140 4.3640 30.2180 4.5900 ;
      RECT 14.8820 4.3640 16.1960 4.5900 ;
      RECT 14.1620 3.4965 14.7920 4.5900 ;
      RECT 0.1400 4.3640 14.1440 4.5900 ;
      RECT 0.0050 3.4965 0.1220 4.5900 ;
      RECT 30.2000 3.4965 30.3530 4.4120 ;
      RECT 16.2680 3.4965 30.1820 4.5900 ;
      RECT 15.5210 3.4965 16.2500 4.4120 ;
      RECT 15.2870 3.6920 15.4850 4.5900 ;
      RECT 14.1080 3.5960 15.2600 4.4120 ;
      RECT 0.1760 3.4965 14.0900 4.5900 ;
      RECT 0.0050 3.4965 0.1580 4.4120 ;
      RECT 15.4670 3.4965 30.3530 4.3160 ;
      RECT 0.0050 3.5960 15.4490 4.3160 ;
      RECT 15.2420 3.4965 30.3530 3.6680 ;
      RECT 0.0050 3.4965 15.2240 4.3160 ;
      RECT 0.0050 3.4965 30.3530 3.5720 ;
      RECT 0.0050 5.5400 30.3530 5.6700 ;
      RECT 30.2360 4.5765 30.3530 5.6700 ;
      RECT 16.2140 5.4440 30.2180 5.6700 ;
      RECT 14.8820 5.4440 16.1960 5.6700 ;
      RECT 14.1620 4.5765 14.7920 5.6700 ;
      RECT 0.1400 5.4440 14.1440 5.6700 ;
      RECT 0.0050 4.5765 0.1220 5.6700 ;
      RECT 30.2000 4.5765 30.3530 5.4920 ;
      RECT 16.2680 4.5765 30.1820 5.6700 ;
      RECT 15.5210 4.5765 16.2500 5.4920 ;
      RECT 15.2870 4.7720 15.4850 5.6700 ;
      RECT 14.1080 4.6760 15.2600 5.4920 ;
      RECT 0.1760 4.5765 14.0900 5.6700 ;
      RECT 0.0050 4.5765 0.1580 5.4920 ;
      RECT 15.4670 4.5765 30.3530 5.3960 ;
      RECT 0.0050 4.6760 15.4490 5.3960 ;
      RECT 15.2420 4.5765 30.3530 4.7480 ;
      RECT 0.0050 4.5765 15.2240 5.3960 ;
      RECT 0.0050 4.5765 30.3530 4.6520 ;
      RECT 0.0050 6.6200 30.3530 6.7500 ;
      RECT 30.2360 5.6565 30.3530 6.7500 ;
      RECT 16.2140 6.5240 30.2180 6.7500 ;
      RECT 14.8820 6.5240 16.1960 6.7500 ;
      RECT 14.1620 5.6565 14.7920 6.7500 ;
      RECT 0.1400 6.5240 14.1440 6.7500 ;
      RECT 0.0050 5.6565 0.1220 6.7500 ;
      RECT 30.2000 5.6565 30.3530 6.5720 ;
      RECT 16.2680 5.6565 30.1820 6.7500 ;
      RECT 15.5210 5.6565 16.2500 6.5720 ;
      RECT 15.2870 5.8520 15.4850 6.7500 ;
      RECT 14.1080 5.7560 15.2600 6.5720 ;
      RECT 0.1760 5.6565 14.0900 6.7500 ;
      RECT 0.0050 5.6565 0.1580 6.5720 ;
      RECT 15.4670 5.6565 30.3530 6.4760 ;
      RECT 0.0050 5.7560 15.4490 6.4760 ;
      RECT 15.2420 5.6565 30.3530 5.8280 ;
      RECT 0.0050 5.6565 15.2240 6.4760 ;
      RECT 0.0050 5.6565 30.3530 5.7320 ;
      RECT 0.0050 7.7000 30.3530 7.8300 ;
      RECT 30.2360 6.7365 30.3530 7.8300 ;
      RECT 16.2140 7.6040 30.2180 7.8300 ;
      RECT 14.8820 7.6040 16.1960 7.8300 ;
      RECT 14.1620 6.7365 14.7920 7.8300 ;
      RECT 0.1400 7.6040 14.1440 7.8300 ;
      RECT 0.0050 6.7365 0.1220 7.8300 ;
      RECT 30.2000 6.7365 30.3530 7.6520 ;
      RECT 16.2680 6.7365 30.1820 7.8300 ;
      RECT 15.5210 6.7365 16.2500 7.6520 ;
      RECT 15.2870 6.9320 15.4850 7.8300 ;
      RECT 14.1080 6.8360 15.2600 7.6520 ;
      RECT 0.1760 6.7365 14.0900 7.8300 ;
      RECT 0.0050 6.7365 0.1580 7.6520 ;
      RECT 15.4670 6.7365 30.3530 7.5560 ;
      RECT 0.0050 6.8360 15.4490 7.5560 ;
      RECT 15.2420 6.7365 30.3530 6.9080 ;
      RECT 0.0050 6.7365 15.2240 7.5560 ;
      RECT 0.0050 6.7365 30.3530 6.8120 ;
      RECT 0.0050 8.7800 30.3530 8.9100 ;
      RECT 30.2360 7.8165 30.3530 8.9100 ;
      RECT 16.2140 8.6840 30.2180 8.9100 ;
      RECT 14.8820 8.6840 16.1960 8.9100 ;
      RECT 14.1620 7.8165 14.7920 8.9100 ;
      RECT 0.1400 8.6840 14.1440 8.9100 ;
      RECT 0.0050 7.8165 0.1220 8.9100 ;
      RECT 30.2000 7.8165 30.3530 8.7320 ;
      RECT 16.2680 7.8165 30.1820 8.9100 ;
      RECT 15.5210 7.8165 16.2500 8.7320 ;
      RECT 15.2870 8.0120 15.4850 8.9100 ;
      RECT 14.1080 7.9160 15.2600 8.7320 ;
      RECT 0.1760 7.8165 14.0900 8.9100 ;
      RECT 0.0050 7.8165 0.1580 8.7320 ;
      RECT 15.4670 7.8165 30.3530 8.6360 ;
      RECT 0.0050 7.9160 15.4490 8.6360 ;
      RECT 15.2420 7.8165 30.3530 7.9880 ;
      RECT 0.0050 7.8165 15.2240 8.6360 ;
      RECT 0.0050 7.8165 30.3530 7.8920 ;
      RECT 0.0050 9.8600 30.3530 9.9900 ;
      RECT 30.2360 8.8965 30.3530 9.9900 ;
      RECT 16.2140 9.7640 30.2180 9.9900 ;
      RECT 14.8820 9.7640 16.1960 9.9900 ;
      RECT 14.1620 8.8965 14.7920 9.9900 ;
      RECT 0.1400 9.7640 14.1440 9.9900 ;
      RECT 0.0050 8.8965 0.1220 9.9900 ;
      RECT 30.2000 8.8965 30.3530 9.8120 ;
      RECT 16.2680 8.8965 30.1820 9.9900 ;
      RECT 15.5210 8.8965 16.2500 9.8120 ;
      RECT 15.2870 9.0920 15.4850 9.9900 ;
      RECT 14.1080 8.9960 15.2600 9.8120 ;
      RECT 0.1760 8.8965 14.0900 9.9900 ;
      RECT 0.0050 8.8965 0.1580 9.8120 ;
      RECT 15.4670 8.8965 30.3530 9.7160 ;
      RECT 0.0050 8.9960 15.4490 9.7160 ;
      RECT 15.2420 8.8965 30.3530 9.0680 ;
      RECT 0.0050 8.8965 15.2240 9.7160 ;
      RECT 0.0050 8.8965 30.3530 8.9720 ;
      RECT 0.0050 10.9400 30.3530 11.0700 ;
      RECT 30.2360 9.9765 30.3530 11.0700 ;
      RECT 16.2140 10.8440 30.2180 11.0700 ;
      RECT 14.8820 10.8440 16.1960 11.0700 ;
      RECT 14.1620 9.9765 14.7920 11.0700 ;
      RECT 0.1400 10.8440 14.1440 11.0700 ;
      RECT 0.0050 9.9765 0.1220 11.0700 ;
      RECT 30.2000 9.9765 30.3530 10.8920 ;
      RECT 16.2680 9.9765 30.1820 11.0700 ;
      RECT 15.5210 9.9765 16.2500 10.8920 ;
      RECT 15.2870 10.1720 15.4850 11.0700 ;
      RECT 14.1080 10.0760 15.2600 10.8920 ;
      RECT 0.1760 9.9765 14.0900 11.0700 ;
      RECT 0.0050 9.9765 0.1580 10.8920 ;
      RECT 15.4670 9.9765 30.3530 10.7960 ;
      RECT 0.0050 10.0760 15.4490 10.7960 ;
      RECT 15.2420 9.9765 30.3530 10.1480 ;
      RECT 0.0050 9.9765 15.2240 10.7960 ;
      RECT 0.0050 9.9765 30.3530 10.0520 ;
      RECT 0.0000 18.4135 30.3480 19.7470 ;
      RECT 17.7210 11.0935 30.3480 19.7470 ;
      RECT 15.5210 12.5575 30.3480 19.7470 ;
      RECT 16.4250 12.3655 30.3480 19.7470 ;
      RECT 15.4690 11.0935 15.5030 19.7470 ;
      RECT 15.4170 11.0935 15.4510 19.7470 ;
      RECT 15.3650 11.0935 15.3990 19.7470 ;
      RECT 15.3130 11.0935 15.3470 19.7470 ;
      RECT 0.0000 12.6535 15.2950 19.7470 ;
      RECT 0.0000 15.2455 30.3480 18.1975 ;
      RECT 14.1570 12.0775 15.8310 15.0295 ;
      RECT 0.0000 12.3655 14.1390 19.7470 ;
      RECT 0.0000 12.4615 16.4070 12.6295 ;
      RECT 16.2090 12.3655 30.3480 12.5335 ;
      RECT 0.0000 12.3655 16.1910 12.6295 ;
      RECT 17.5050 11.0935 17.7030 19.7470 ;
      RECT 13.7250 12.1735 17.4870 12.4375 ;
      RECT 12.8610 11.7895 13.7070 19.7470 ;
      RECT 0.0000 11.0935 12.8430 19.7470 ;
      RECT 17.2890 11.0935 30.3480 12.3415 ;
      RECT 17.0730 11.7895 30.3480 12.3415 ;
      RECT 15.8490 12.0775 17.0550 12.4375 ;
      RECT 0.0000 12.0775 15.8310 12.3415 ;
      RECT 16.8570 11.0935 17.2710 12.1495 ;
      RECT 16.2630 11.7895 30.3480 12.1495 ;
      RECT 15.5210 11.7895 16.2450 12.1495 ;
      RECT 14.1030 11.7895 15.2950 12.6295 ;
      RECT 0.0000 11.7895 14.0850 12.3415 ;
      RECT 15.5610 11.7415 16.8390 11.8615 ;
      RECT 14.3730 11.7415 15.5430 11.8615 ;
      RECT 13.5090 11.7415 14.3550 11.8615 ;
      RECT 13.0770 11.7415 13.4910 19.7470 ;
      RECT 0.0000 11.0935 13.0590 12.3415 ;
      RECT 16.6410 11.0935 30.3480 11.7655 ;
      RECT 15.1650 11.0935 16.6230 11.7655 ;
      RECT 14.1930 11.0935 15.1470 11.7655 ;
      RECT 13.2930 11.0935 14.1750 11.7655 ;
      RECT 0.0000 11.0935 13.2750 11.7655 ;
      RECT 0.0000 11.0935 30.3480 11.7175 ;
        RECT 0.0050 20.1470 30.3530 20.2770 ;
        RECT 30.2360 19.1835 30.3530 20.2770 ;
        RECT 16.2140 20.0510 30.2180 20.2770 ;
        RECT 14.8820 20.0510 16.1960 20.2770 ;
        RECT 14.1620 19.1835 14.7920 20.2770 ;
        RECT 0.1400 20.0510 14.1440 20.2770 ;
        RECT 0.0050 19.1835 0.1220 20.2770 ;
        RECT 30.2000 19.1835 30.3530 20.0990 ;
        RECT 16.2680 19.1835 30.1820 20.2770 ;
        RECT 15.5210 19.1835 16.2500 20.0990 ;
        RECT 15.2870 19.3790 15.4850 20.2770 ;
        RECT 14.1080 19.2830 15.2600 20.0990 ;
        RECT 0.1760 19.1835 14.0900 20.2770 ;
        RECT 0.0050 19.1835 0.1580 20.0990 ;
        RECT 15.4670 19.1835 30.3530 20.0030 ;
        RECT 0.0050 19.2830 15.4490 20.0030 ;
        RECT 15.2420 19.1835 30.3530 19.3550 ;
        RECT 0.0050 19.1835 15.2240 20.0030 ;
        RECT 0.0050 19.1835 30.3530 19.2590 ;
        RECT 0.0050 21.2270 30.3530 21.3570 ;
        RECT 30.2360 20.2635 30.3530 21.3570 ;
        RECT 16.2140 21.1310 30.2180 21.3570 ;
        RECT 14.8820 21.1310 16.1960 21.3570 ;
        RECT 14.1620 20.2635 14.7920 21.3570 ;
        RECT 0.1400 21.1310 14.1440 21.3570 ;
        RECT 0.0050 20.2635 0.1220 21.3570 ;
        RECT 30.2000 20.2635 30.3530 21.1790 ;
        RECT 16.2680 20.2635 30.1820 21.3570 ;
        RECT 15.5210 20.2635 16.2500 21.1790 ;
        RECT 15.2870 20.4590 15.4850 21.3570 ;
        RECT 14.1080 20.3630 15.2600 21.1790 ;
        RECT 0.1760 20.2635 14.0900 21.3570 ;
        RECT 0.0050 20.2635 0.1580 21.1790 ;
        RECT 15.4670 20.2635 30.3530 21.0830 ;
        RECT 0.0050 20.3630 15.4490 21.0830 ;
        RECT 15.2420 20.2635 30.3530 20.4350 ;
        RECT 0.0050 20.2635 15.2240 21.0830 ;
        RECT 0.0050 20.2635 30.3530 20.3390 ;
        RECT 0.0050 22.3070 30.3530 22.4370 ;
        RECT 30.2360 21.3435 30.3530 22.4370 ;
        RECT 16.2140 22.2110 30.2180 22.4370 ;
        RECT 14.8820 22.2110 16.1960 22.4370 ;
        RECT 14.1620 21.3435 14.7920 22.4370 ;
        RECT 0.1400 22.2110 14.1440 22.4370 ;
        RECT 0.0050 21.3435 0.1220 22.4370 ;
        RECT 30.2000 21.3435 30.3530 22.2590 ;
        RECT 16.2680 21.3435 30.1820 22.4370 ;
        RECT 15.5210 21.3435 16.2500 22.2590 ;
        RECT 15.2870 21.5390 15.4850 22.4370 ;
        RECT 14.1080 21.4430 15.2600 22.2590 ;
        RECT 0.1760 21.3435 14.0900 22.4370 ;
        RECT 0.0050 21.3435 0.1580 22.2590 ;
        RECT 15.4670 21.3435 30.3530 22.1630 ;
        RECT 0.0050 21.4430 15.4490 22.1630 ;
        RECT 15.2420 21.3435 30.3530 21.5150 ;
        RECT 0.0050 21.3435 15.2240 22.1630 ;
        RECT 0.0050 21.3435 30.3530 21.4190 ;
        RECT 0.0050 23.3870 30.3530 23.5170 ;
        RECT 30.2360 22.4235 30.3530 23.5170 ;
        RECT 16.2140 23.2910 30.2180 23.5170 ;
        RECT 14.8820 23.2910 16.1960 23.5170 ;
        RECT 14.1620 22.4235 14.7920 23.5170 ;
        RECT 0.1400 23.2910 14.1440 23.5170 ;
        RECT 0.0050 22.4235 0.1220 23.5170 ;
        RECT 30.2000 22.4235 30.3530 23.3390 ;
        RECT 16.2680 22.4235 30.1820 23.5170 ;
        RECT 15.5210 22.4235 16.2500 23.3390 ;
        RECT 15.2870 22.6190 15.4850 23.5170 ;
        RECT 14.1080 22.5230 15.2600 23.3390 ;
        RECT 0.1760 22.4235 14.0900 23.5170 ;
        RECT 0.0050 22.4235 0.1580 23.3390 ;
        RECT 15.4670 22.4235 30.3530 23.2430 ;
        RECT 0.0050 22.5230 15.4490 23.2430 ;
        RECT 15.2420 22.4235 30.3530 22.5950 ;
        RECT 0.0050 22.4235 15.2240 23.2430 ;
        RECT 0.0050 22.4235 30.3530 22.4990 ;
        RECT 0.0050 24.4670 30.3530 24.5970 ;
        RECT 30.2360 23.5035 30.3530 24.5970 ;
        RECT 16.2140 24.3710 30.2180 24.5970 ;
        RECT 14.8820 24.3710 16.1960 24.5970 ;
        RECT 14.1620 23.5035 14.7920 24.5970 ;
        RECT 0.1400 24.3710 14.1440 24.5970 ;
        RECT 0.0050 23.5035 0.1220 24.5970 ;
        RECT 30.2000 23.5035 30.3530 24.4190 ;
        RECT 16.2680 23.5035 30.1820 24.5970 ;
        RECT 15.5210 23.5035 16.2500 24.4190 ;
        RECT 15.2870 23.6990 15.4850 24.5970 ;
        RECT 14.1080 23.6030 15.2600 24.4190 ;
        RECT 0.1760 23.5035 14.0900 24.5970 ;
        RECT 0.0050 23.5035 0.1580 24.4190 ;
        RECT 15.4670 23.5035 30.3530 24.3230 ;
        RECT 0.0050 23.6030 15.4490 24.3230 ;
        RECT 15.2420 23.5035 30.3530 23.6750 ;
        RECT 0.0050 23.5035 15.2240 24.3230 ;
        RECT 0.0050 23.5035 30.3530 23.5790 ;
        RECT 0.0050 25.5470 30.3530 25.6770 ;
        RECT 30.2360 24.5835 30.3530 25.6770 ;
        RECT 16.2140 25.4510 30.2180 25.6770 ;
        RECT 14.8820 25.4510 16.1960 25.6770 ;
        RECT 14.1620 24.5835 14.7920 25.6770 ;
        RECT 0.1400 25.4510 14.1440 25.6770 ;
        RECT 0.0050 24.5835 0.1220 25.6770 ;
        RECT 30.2000 24.5835 30.3530 25.4990 ;
        RECT 16.2680 24.5835 30.1820 25.6770 ;
        RECT 15.5210 24.5835 16.2500 25.4990 ;
        RECT 15.2870 24.7790 15.4850 25.6770 ;
        RECT 14.1080 24.6830 15.2600 25.4990 ;
        RECT 0.1760 24.5835 14.0900 25.6770 ;
        RECT 0.0050 24.5835 0.1580 25.4990 ;
        RECT 15.4670 24.5835 30.3530 25.4030 ;
        RECT 0.0050 24.6830 15.4490 25.4030 ;
        RECT 15.2420 24.5835 30.3530 24.7550 ;
        RECT 0.0050 24.5835 15.2240 25.4030 ;
        RECT 0.0050 24.5835 30.3530 24.6590 ;
        RECT 0.0050 26.6270 30.3530 26.7570 ;
        RECT 30.2360 25.6635 30.3530 26.7570 ;
        RECT 16.2140 26.5310 30.2180 26.7570 ;
        RECT 14.8820 26.5310 16.1960 26.7570 ;
        RECT 14.1620 25.6635 14.7920 26.7570 ;
        RECT 0.1400 26.5310 14.1440 26.7570 ;
        RECT 0.0050 25.6635 0.1220 26.7570 ;
        RECT 30.2000 25.6635 30.3530 26.5790 ;
        RECT 16.2680 25.6635 30.1820 26.7570 ;
        RECT 15.5210 25.6635 16.2500 26.5790 ;
        RECT 15.2870 25.8590 15.4850 26.7570 ;
        RECT 14.1080 25.7630 15.2600 26.5790 ;
        RECT 0.1760 25.6635 14.0900 26.7570 ;
        RECT 0.0050 25.6635 0.1580 26.5790 ;
        RECT 15.4670 25.6635 30.3530 26.4830 ;
        RECT 0.0050 25.7630 15.4490 26.4830 ;
        RECT 15.2420 25.6635 30.3530 25.8350 ;
        RECT 0.0050 25.6635 15.2240 26.4830 ;
        RECT 0.0050 25.6635 30.3530 25.7390 ;
        RECT 0.0050 27.7070 30.3530 27.8370 ;
        RECT 30.2360 26.7435 30.3530 27.8370 ;
        RECT 16.2140 27.6110 30.2180 27.8370 ;
        RECT 14.8820 27.6110 16.1960 27.8370 ;
        RECT 14.1620 26.7435 14.7920 27.8370 ;
        RECT 0.1400 27.6110 14.1440 27.8370 ;
        RECT 0.0050 26.7435 0.1220 27.8370 ;
        RECT 30.2000 26.7435 30.3530 27.6590 ;
        RECT 16.2680 26.7435 30.1820 27.8370 ;
        RECT 15.5210 26.7435 16.2500 27.6590 ;
        RECT 15.2870 26.9390 15.4850 27.8370 ;
        RECT 14.1080 26.8430 15.2600 27.6590 ;
        RECT 0.1760 26.7435 14.0900 27.8370 ;
        RECT 0.0050 26.7435 0.1580 27.6590 ;
        RECT 15.4670 26.7435 30.3530 27.5630 ;
        RECT 0.0050 26.8430 15.4490 27.5630 ;
        RECT 15.2420 26.7435 30.3530 26.9150 ;
        RECT 0.0050 26.7435 15.2240 27.5630 ;
        RECT 0.0050 26.7435 30.3530 26.8190 ;
        RECT 0.0050 28.7870 30.3530 28.9170 ;
        RECT 30.2360 27.8235 30.3530 28.9170 ;
        RECT 16.2140 28.6910 30.2180 28.9170 ;
        RECT 14.8820 28.6910 16.1960 28.9170 ;
        RECT 14.1620 27.8235 14.7920 28.9170 ;
        RECT 0.1400 28.6910 14.1440 28.9170 ;
        RECT 0.0050 27.8235 0.1220 28.9170 ;
        RECT 30.2000 27.8235 30.3530 28.7390 ;
        RECT 16.2680 27.8235 30.1820 28.9170 ;
        RECT 15.5210 27.8235 16.2500 28.7390 ;
        RECT 15.2870 28.0190 15.4850 28.9170 ;
        RECT 14.1080 27.9230 15.2600 28.7390 ;
        RECT 0.1760 27.8235 14.0900 28.9170 ;
        RECT 0.0050 27.8235 0.1580 28.7390 ;
        RECT 15.4670 27.8235 30.3530 28.6430 ;
        RECT 0.0050 27.9230 15.4490 28.6430 ;
        RECT 15.2420 27.8235 30.3530 27.9950 ;
        RECT 0.0050 27.8235 15.2240 28.6430 ;
        RECT 0.0050 27.8235 30.3530 27.8990 ;
        RECT 0.0050 29.8670 30.3530 29.9970 ;
        RECT 30.2360 28.9035 30.3530 29.9970 ;
        RECT 16.2140 29.7710 30.2180 29.9970 ;
        RECT 14.8820 29.7710 16.1960 29.9970 ;
        RECT 14.1620 28.9035 14.7920 29.9970 ;
        RECT 0.1400 29.7710 14.1440 29.9970 ;
        RECT 0.0050 28.9035 0.1220 29.9970 ;
        RECT 30.2000 28.9035 30.3530 29.8190 ;
        RECT 16.2680 28.9035 30.1820 29.9970 ;
        RECT 15.5210 28.9035 16.2500 29.8190 ;
        RECT 15.2870 29.0990 15.4850 29.9970 ;
        RECT 14.1080 29.0030 15.2600 29.8190 ;
        RECT 0.1760 28.9035 14.0900 29.9970 ;
        RECT 0.0050 28.9035 0.1580 29.8190 ;
        RECT 15.4670 28.9035 30.3530 29.7230 ;
        RECT 0.0050 29.0030 15.4490 29.7230 ;
        RECT 15.2420 28.9035 30.3530 29.0750 ;
        RECT 0.0050 28.9035 15.2240 29.7230 ;
        RECT 0.0050 28.9035 30.3530 28.9790 ;
  LAYER M4  ;
      RECT 1.6000 12.8065 28.8355 12.8305 ;
      RECT 1.6000 13.0945 28.8355 13.1185 ;
      RECT 1.6000 13.4785 28.8355 13.5025 ;
      RECT 1.6000 13.5745 28.8355 13.5985 ;
      RECT 1.6000 13.9105 28.8355 13.9345 ;
      RECT 1.6000 14.2945 28.8355 14.3185 ;
      RECT 1.6000 14.3905 28.8355 14.4145 ;
      RECT 10.4760 11.4295 19.8720 11.6455 ;
      RECT 17.8670 11.7655 17.9510 11.7895 ;
      RECT 17.6785 12.1975 17.8085 12.2215 ;
      RECT 17.6870 13.1425 17.8040 13.1665 ;
      RECT 17.6865 12.8550 17.8035 12.8790 ;
      RECT 17.0375 12.1975 17.6085 12.2215 ;
      RECT 17.0975 12.9625 17.2055 12.9865 ;
      RECT 15.7750 13.3495 16.8680 13.3735 ;
      RECT 16.4630 12.9175 16.5470 12.9415 ;
      RECT 15.6790 14.1175 16.5470 14.1415 ;
      RECT 16.4630 14.2135 16.5470 14.2375 ;
      RECT 16.2850 12.4375 16.3690 12.4615 ;
      RECT 16.2470 13.7815 16.3310 13.8055 ;
      RECT 16.2470 14.5015 16.3310 14.5255 ;
      RECT 15.9780 11.1495 16.2410 11.1735 ;
      RECT 16.1090 14.9335 16.2210 14.9575 ;
      RECT 16.0690 12.3415 16.1530 12.3655 ;
      RECT 15.8550 11.0535 16.1180 11.0775 ;
      RECT 15.8550 19.6585 16.1180 19.6825 ;
      RECT 15.8710 13.8295 16.1150 13.8535 ;
      RECT 16.0310 13.9735 16.1150 13.9975 ;
      RECT 14.5750 14.2135 16.1150 14.2375 ;
      RECT 16.0310 14.5015 16.1150 14.5255 ;
      RECT 15.7970 19.5625 16.0600 19.5865 ;
      RECT 15.7960 10.9575 16.0590 10.9815 ;
      RECT 14.3100 14.5975 16.0380 14.8135 ;
      RECT 14.3100 17.7655 16.0380 17.9815 ;
      RECT 15.7580 10.8615 16.0210 10.8855 ;
      RECT 15.7580 19.3705 16.0210 19.3945 ;
      RECT 15.9230 14.9335 16.0070 14.9575 ;
      RECT 15.1510 15.3175 16.0070 15.3415 ;
      RECT 15.5350 17.5735 16.0070 17.5975 ;
      RECT 15.9230 17.6695 16.0070 17.6935 ;
      RECT 15.7100 10.7655 15.9730 10.7895 ;
      RECT 15.7100 19.2745 15.9730 19.2985 ;
      RECT 15.4870 16.6615 15.9320 16.6855 ;
      RECT 15.6660 10.6695 15.9290 10.6935 ;
      RECT 15.6660 19.6105 15.9290 19.6345 ;
      RECT 15.6170 11.0055 15.8800 11.0295 ;
      RECT 15.6170 19.5145 15.8800 19.5385 ;
      RECT 15.7480 13.9735 15.8690 13.9975 ;
      RECT 15.7270 16.0855 15.8600 16.1095 ;
      RECT 15.5700 10.9095 15.8330 10.9335 ;
      RECT 15.5700 19.4185 15.8330 19.4425 ;
      RECT 15.5350 10.6215 15.7980 10.6455 ;
      RECT 15.5350 19.3225 15.7980 19.3465 ;
      RECT 14.7190 17.6695 15.7880 17.6935 ;
      RECT 15.7040 18.8215 15.7880 18.8455 ;
      RECT 15.4790 10.4775 15.7420 10.5015 ;
      RECT 15.4790 19.2265 15.7420 19.2505 ;
      RECT 15.6310 14.9335 15.7160 14.9575 ;
      RECT 14.5270 15.5095 15.6440 15.5335 ;
      RECT 15.1720 13.3495 15.6290 13.3735 ;
      RECT 14.9990 11.1975 15.2660 11.2215 ;
      RECT 14.9990 19.0825 15.2660 19.1065 ;
      RECT 15.1360 14.8855 15.2450 14.9095 ;
      RECT 14.9760 11.1015 15.2180 11.1255 ;
      RECT 14.9760 19.7065 15.2180 19.7305 ;
      RECT 14.9200 10.6215 15.1620 10.6455 ;
      RECT 14.9490 19.8025 15.1620 19.8265 ;
      RECT 15.0650 14.5015 15.1490 14.5255 ;
      RECT 14.8660 10.7175 15.1140 10.7415 ;
      RECT 14.8660 19.6585 15.1140 19.6825 ;
      RECT 14.6320 17.0935 15.0530 17.1175 ;
      RECT 14.6000 11.0535 14.8670 11.0775 ;
      RECT 14.6000 19.8025 14.8670 19.8265 ;
      RECT 14.7400 15.6535 14.8610 15.6775 ;
      RECT 14.7320 18.8215 14.8160 18.8455 ;
      RECT 14.5660 10.9575 14.8130 10.9815 ;
      RECT 14.4990 19.3705 14.8130 19.3945 ;
      RECT 14.5400 10.8615 14.7700 10.8855 ;
      RECT 14.5280 19.7065 14.7700 19.7305 ;
      RECT 14.4870 10.7655 14.7170 10.7895 ;
      RECT 14.6330 17.2375 14.7170 17.2615 ;
      RECT 14.4370 19.2745 14.7170 19.2985 ;
      RECT 14.4420 10.6695 14.6720 10.6935 ;
      RECT 14.4420 19.6105 14.6720 19.6345 ;
      RECT 13.4800 14.5015 14.6690 14.5255 ;
      RECT 14.4040 10.9095 14.6340 10.9335 ;
      RECT 14.4040 19.5145 14.6340 19.5385 ;
      RECT 14.3860 10.8135 14.5790 10.8375 ;
      RECT 14.3860 19.4185 14.5790 19.4425 ;
      RECT 14.3370 10.7175 14.5300 10.7415 ;
      RECT 14.3370 19.3225 14.5300 19.3465 ;
      RECT 14.3410 15.4135 14.5250 15.4375 ;
      RECT 14.2850 10.6215 14.4780 10.6455 ;
      RECT 14.2850 19.2265 14.4780 19.2505 ;
      RECT 13.8010 12.7255 14.4770 12.7495 ;
      RECT 14.3410 15.5095 14.4250 15.5335 ;
      RECT 14.0720 11.1495 14.3350 11.1735 ;
      RECT 14.1950 13.3495 14.2790 13.3735 ;
      RECT 14.1260 14.9335 14.2380 14.9575 ;
      RECT 13.7630 12.9175 13.8470 12.9415 ;
  LAYER V4  ;
      RECT 17.9160 11.7655 17.9400 11.7895 ;
      RECT 17.9160 12.8065 17.9400 12.8305 ;
      RECT 17.7480 12.8550 17.7720 12.8790 ;
      RECT 17.7480 13.1425 17.7720 13.1665 ;
      RECT 17.7475 12.1975 17.7715 12.2215 ;
      RECT 17.1135 12.1975 17.1375 12.2215 ;
      RECT 17.1135 12.9625 17.1375 12.9865 ;
      RECT 16.5120 12.9175 16.5360 12.9415 ;
      RECT 16.5120 13.0945 16.5360 13.1185 ;
      RECT 16.5120 14.1175 16.5360 14.1415 ;
      RECT 16.5120 14.2135 16.5360 14.2375 ;
      RECT 16.2960 12.4375 16.3200 12.4615 ;
      RECT 16.2960 13.4785 16.3200 13.5025 ;
      RECT 16.2960 13.7815 16.3200 13.8055 ;
      RECT 16.2960 13.9105 16.3200 13.9345 ;
      RECT 16.2960 14.2945 16.3200 14.3185 ;
      RECT 16.2960 14.5015 16.3200 14.5255 ;
      RECT 16.1270 11.1495 16.1510 11.1735 ;
      RECT 16.1280 11.4295 16.1510 11.6455 ;
      RECT 16.1270 14.9335 16.1510 14.9575 ;
      RECT 16.0800 12.3415 16.1040 12.3655 ;
      RECT 16.0800 13.5745 16.1040 13.5985 ;
      RECT 16.0800 13.8295 16.1040 13.8535 ;
      RECT 16.0800 13.9735 16.1040 13.9975 ;
      RECT 16.0800 14.2135 16.1040 14.2375 ;
      RECT 16.0800 14.5015 16.1040 14.5255 ;
      RECT 15.9720 14.9335 15.9960 14.9575 ;
      RECT 15.9720 15.3175 15.9960 15.3415 ;
      RECT 15.9720 17.5735 15.9960 17.5975 ;
      RECT 15.9720 17.6695 15.9960 17.6935 ;
      RECT 15.8820 11.0535 15.9060 11.0775 ;
      RECT 15.8820 13.8295 15.9060 13.8535 ;
      RECT 15.8820 19.6585 15.9060 19.6825 ;
      RECT 15.8340 10.9575 15.8580 10.9815 ;
      RECT 15.8340 13.9735 15.8580 13.9975 ;
      RECT 15.8340 19.5625 15.8580 19.5865 ;
      RECT 15.7860 10.8615 15.8100 10.8855 ;
      RECT 15.7860 13.3495 15.8100 13.3735 ;
      RECT 15.7860 19.3705 15.8100 19.3945 ;
      RECT 15.7380 10.7655 15.7620 10.7895 ;
      RECT 15.7380 16.0855 15.7620 16.1095 ;
      RECT 15.7380 18.8215 15.7620 18.8455 ;
      RECT 15.7380 19.2745 15.7620 19.2985 ;
      RECT 15.6900 10.6695 15.7140 10.6935 ;
      RECT 15.6900 14.1175 15.7140 14.1415 ;
      RECT 15.6900 19.6105 15.7140 19.6345 ;
      RECT 15.6420 11.0055 15.6660 11.0295 ;
      RECT 15.6420 14.9335 15.6660 14.9575 ;
      RECT 15.6420 19.5145 15.6660 19.5385 ;
      RECT 15.5940 10.9095 15.6180 10.9335 ;
      RECT 15.5940 13.3495 15.6180 13.3735 ;
      RECT 15.5940 19.4185 15.6180 19.4425 ;
      RECT 15.5460 10.6215 15.5700 10.6455 ;
      RECT 15.5460 17.5735 15.5700 17.5975 ;
      RECT 15.5460 19.3225 15.5700 19.3465 ;
      RECT 15.4980 10.4775 15.5220 10.5015 ;
      RECT 15.4980 16.6615 15.5220 16.6855 ;
      RECT 15.4980 19.2265 15.5220 19.2505 ;
      RECT 15.2100 11.1975 15.2340 11.2215 ;
      RECT 15.2100 14.8855 15.2340 14.9095 ;
      RECT 15.2100 19.0825 15.2340 19.1065 ;
      RECT 15.1620 11.1015 15.1860 11.1255 ;
      RECT 15.1620 15.3175 15.1860 15.3415 ;
      RECT 15.1620 19.7065 15.1860 19.7305 ;
      RECT 15.1140 10.6215 15.1380 10.6455 ;
      RECT 15.1140 14.5015 15.1380 14.5255 ;
      RECT 15.1140 19.8025 15.1380 19.8265 ;
      RECT 15.0180 10.7175 15.0420 10.7415 ;
      RECT 15.0180 17.0935 15.0420 17.1175 ;
      RECT 15.0180 19.6585 15.0420 19.6825 ;
      RECT 14.8260 11.0535 14.8500 11.0775 ;
      RECT 14.8260 15.6535 14.8500 15.6775 ;
      RECT 14.8260 19.8025 14.8500 19.8265 ;
      RECT 14.7780 10.9575 14.8020 10.9815 ;
      RECT 14.7780 18.8215 14.8020 18.8455 ;
      RECT 14.7780 19.3705 14.8020 19.3945 ;
      RECT 14.7300 10.8615 14.7540 10.8855 ;
      RECT 14.7300 17.6695 14.7540 17.6935 ;
      RECT 14.7300 19.7065 14.7540 19.7305 ;
      RECT 14.6820 10.7655 14.7060 10.7895 ;
      RECT 14.6820 17.2375 14.7060 17.2615 ;
      RECT 14.6820 19.2745 14.7060 19.2985 ;
      RECT 14.6340 10.6695 14.6580 10.6935 ;
      RECT 14.6340 14.5015 14.6580 14.5255 ;
      RECT 14.6340 19.6105 14.6580 19.6345 ;
      RECT 14.5860 10.9095 14.6100 10.9335 ;
      RECT 14.5860 14.2135 14.6100 14.2375 ;
      RECT 14.5860 19.5145 14.6100 19.5385 ;
      RECT 14.5380 10.8135 14.5620 10.8375 ;
      RECT 14.5380 15.5095 14.5620 15.5335 ;
      RECT 14.5380 19.4185 14.5620 19.4425 ;
      RECT 14.4900 10.7175 14.5140 10.7415 ;
      RECT 14.4900 15.4135 14.5140 15.4375 ;
      RECT 14.4900 19.3225 14.5140 19.3465 ;
      RECT 14.4420 10.6215 14.4660 10.6455 ;
      RECT 14.4420 12.7255 14.4660 12.7495 ;
      RECT 14.4420 19.2265 14.4660 19.2505 ;
      RECT 14.3520 15.4135 14.3760 15.4375 ;
      RECT 14.3520 15.5095 14.3760 15.5335 ;
      RECT 14.2440 13.3495 14.2680 13.3735 ;
      RECT 14.2440 14.3905 14.2680 14.4145 ;
      RECT 14.1840 11.1495 14.2080 11.1735 ;
      RECT 14.1850 11.4295 14.2080 11.6455 ;
      RECT 14.1840 14.9335 14.2080 14.9575 ;
      RECT 13.8120 12.7255 13.8360 12.7495 ;
      RECT 13.8120 12.9175 13.8360 12.9415 ;
  LAYER M5  ;
      RECT 17.9160 11.7545 17.9400 12.8415 ;
      RECT 17.7475 12.1520 17.7715 13.2125 ;
      RECT 17.1135 12.1560 17.1375 13.0270 ;
      RECT 16.5120 12.9065 16.5360 13.1295 ;
      RECT 16.5120 14.1065 16.5360 14.2485 ;
      RECT 16.2960 12.4265 16.3200 13.5135 ;
      RECT 16.2960 13.7705 16.3200 13.9455 ;
      RECT 16.2960 14.2835 16.3200 14.5365 ;
      RECT 16.1270 11.1315 16.1510 14.9755 ;
      RECT 16.0800 12.3305 16.1040 13.6095 ;
      RECT 16.0800 13.8185 16.1040 14.0085 ;
      RECT 16.0800 14.2025 16.1040 14.5365 ;
      RECT 15.9720 14.9225 15.9960 15.3525 ;
      RECT 15.9720 17.5625 15.9960 17.7045 ;
      RECT 15.8820 10.4010 15.9060 19.9025 ;
      RECT 15.8340 10.4010 15.8580 19.9015 ;
      RECT 15.7860 10.4010 15.8100 19.9015 ;
      RECT 15.7380 10.4010 15.7620 19.8725 ;
      RECT 15.6900 10.4010 15.7140 19.8695 ;
      RECT 15.6420 10.4010 15.6660 19.8715 ;
      RECT 15.5940 10.4010 15.6180 19.8645 ;
      RECT 15.5460 10.4010 15.5700 19.8805 ;
      RECT 15.4980 10.4010 15.5220 19.8795 ;
      RECT 15.2100 10.6065 15.2340 19.9355 ;
      RECT 15.1620 10.6075 15.1860 19.9365 ;
      RECT 15.1140 10.6065 15.1380 19.9355 ;
      RECT 15.0180 10.6225 15.0420 19.9365 ;
      RECT 14.8260 10.6215 14.8500 19.8895 ;
      RECT 14.7780 10.6215 14.8020 19.8895 ;
      RECT 14.7300 10.6215 14.7540 19.8895 ;
      RECT 14.6820 10.6215 14.7060 19.8895 ;
      RECT 14.6340 10.6215 14.6580 19.8895 ;
      RECT 14.5860 10.5925 14.6100 19.8895 ;
      RECT 14.5380 10.5485 14.5620 19.6035 ;
      RECT 14.4900 10.5115 14.5140 19.5575 ;
      RECT 14.4420 10.4575 14.4660 19.5035 ;
      RECT 14.3520 15.4025 14.3760 15.5445 ;
      RECT 14.2440 13.3385 14.2680 14.4255 ;
      RECT 14.1840 11.1315 14.2080 14.9755 ;
      RECT 13.8120 12.7145 13.8360 12.9525 ;
  LAYER M2  ;
    RECT 0.108 0.036 30.2400 30.2040 ;
  LAYER M1  ;
    RECT 0.108 0.036 30.2400 30.2040 ;
  END
END srambank_256x4x20_6t122 
